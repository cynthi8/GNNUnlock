//key=0010100101011010
// Main module
module c7552_AntiSAT_16(1, 5, 9, 12, 15, 18, 23, 26, 29, 32, 35, 38, 41, 44, 47, 50, 53, 54, 55, 56, 57, 58, 59, 60, 61, 62, 63, 64, 65, 66, 69, 70, 73, 74, 75, 76, 77, 78, 79, 80, 81, 82, 83, 84, 85, 86, 87, 88, 89, 94, 97, 100, 103, 106, 109, 110, 111, 112, 113, 114, 115, 118, 121, 124, 127, 130, 133, 134, 135, 138, 141, 144, 147, 150, 151, 152, 153, 154, 155, 156, 157, 158, 159, 160, 161, 162, 163, 164, 165, 166, 167, 168, 169, 170, 171, 172, 173, 174, 175, 176, 177, 178, 179, 180, 181, 182, 183, 184, 185, 186, 187, 188, 189, 190, 191, 192, 193, 194, 195, 196, 197, 198, 199, 200, 201, 202, 203, 204, 205, 206, 207, 208, 209, 210, 211, 212, 213, 214, 215, 216, 217, 218, 219, 220, 221, 222, 223, 224, 225, 226, 227, 228, 229, 230, 231, 232, 233, 234, 235, 236, 237, 238, 239, 240, 241, 242, 245, 248, 251, 254, 257, 260, 263, 267, 271, 274, 277, 280, 283, 286, 289, 293, 296, 299, 303, 307, 310, 313, 316, 319, 322, 325, 328, 331, 334, 337, 340, 343, 346, 349, 352, 355, 358, 361, 364, 367, 382, keyinput0, keyinput1, keyinput2, keyinput3, keyinput4, keyinput5, keyinput6, keyinput7, keyinput8, keyinput9, keyinput10, keyinput11, keyinput12, keyinput13, keyinput14, keyinput15, 241, 387, 388, 478, 482, 484, 486, 489, 492, 501, 505, 507, 509, 511, 513, 515, 517, 519, 535, 537, 539, 541, 543, 545, 547, 549, 551, 553, 556, 559, 561, 563, 565, 567, 569, 571, 573, 582, 643, 707, 813, 881, 882, 883, 884, 885, 889, 945, 1110, 1111, 1112, 1113, 1114, 1489, 1490, 1781, 10025, 10101, 10102, 10103, 10104, 10109, 10110, 10111, 10112, 10350, 10351, 10352, 10353, 10574, 10575, 10576, 10628, 10632, 10641, 10704, 10706, 10711, 10712, 10713, 10714, 10715, 10716, 10717, 10718, 10729, 10759, 10760, 10761, 10762, 10763, 10827, 10837, 10838, 10839, 10840, 10868, 10869, 10870, 10871, 10905, 10906, 10907, 10908, 11333, 11334, 11340, 11342);

  input 1, 5, 9, 12, 15, 18, 23, 26, 29, 32, 35, 38, 41, 44, 47, 50, 53, 54, 55, 56, 57, 58, 59, 60, 61, 62, 63, 64, 65, 66, 69, 70, 73, 74, 75, 76, 77, 78, 79, 80, 81, 82, 83, 84, 85, 86, 87, 88, 89, 94, 97, 100, 103, 106, 109, 110, 111, 112, 113, 114, 115, 118, 121, 124, 127, 130, 133, 134, 135, 138, 141, 144, 147, 150, 151, 152, 153, 154, 155, 156, 157, 158, 159, 160, 161, 162, 163, 164, 165, 166, 167, 168, 169, 170, 171, 172, 173, 174, 175, 176, 177, 178, 179, 180, 181, 182, 183, 184, 185, 186, 187, 188, 189, 190, 191, 192, 193, 194, 195, 196, 197, 198, 199, 200, 201, 202, 203, 204, 205, 206, 207, 208, 209, 210, 211, 212, 213, 214, 215, 216, 217, 218, 219, 220, 221, 222, 223, 224, 225, 226, 227, 228, 229, 230, 231, 232, 233, 234, 235, 236, 237, 238, 239, 240, 241, 242, 245, 248, 251, 254, 257, 260, 263, 267, 271, 274, 277, 280, 283, 286, 289, 293, 296, 299, 303, 307, 310, 313, 316, 319, 322, 325, 328, 331, 334, 337, 340, 343, 346, 349, 352, 355, 358, 361, 364, 367, 382, keyinput0, keyinput1, keyinput2, keyinput3, keyinput4, keyinput5, keyinput6, keyinput7, keyinput8, keyinput9, keyinput10, keyinput11, keyinput12, keyinput13, keyinput14, keyinput15;
  output 241, 387, 388, 478, 482, 484, 486, 489, 492, 501, 505, 507, 509, 511, 513, 515, 517, 519, 535, 537, 539, 541, 543, 545, 547, 549, 551, 553, 556, 559, 561, 563, 565, 567, 569, 571, 573, 582, 643, 707, 813, 881, 882, 883, 884, 885, 889, 945, 1110, 1111, 1112, 1113, 1114, 1489, 1490, 1781, 10025, 10101, 10102, 10103, 10104, 10109, 10110, 10111, 10112, 10350, 10351, 10352, 10353, 10574, 10575, 10576, 10628, 10632, 10641, 10704, 10706, 10711, 10712, 10713, 10714, 10715, 10716, 10717, 10718, 10729, 10759, 10760, 10761, 10762, 10763, 10827, 10837, 10838, 10839, 10840, 10868, 10869, 10870, 10871, 10905, 10906, 10907, 10908, 11333, 11334, 11340, 11342;
  wire 10002, 10003, 10006, 10007, 10010, 10013, 10014, 10015, 10016, 10017, 10018, 10019, 10020, 10021, 10022, 10023, 10024, 10026, 10028, 10032, 10033, 10034, 10035, 10036, 10037, 10038, 10039, 10040, 10041, 10042, 10043, 10050, 10053, 10054, 10055, 10056, 10057, 10058, 10059, 10060, 10061, 10062, 10067, 10070, 10073, 10076, 10077, 10082, 10083, 10084, 10085, 10086, 10093, 10094, 10105, 10106, 10107, 10108, 10113, 10114, 10115, 10116, 10119, 10124, 10130, 10131, 10132, 10133, 10134, 10135, 10136, 10137, 10138, 10139, 10140, 10141, 10148, 10155, 10156, 10157, 10158, 10159, 10160, 10161, 10162, 10163, 10164, 10165, 10170, 10173, 10176, 10177, 10178, 10179, 10180, 10183, 10186, 10189, 10192, 10195, 10196, 10197, 10200, 10203, 10204, 10205, 10206, 10212, 10213, 10230, 10231, 10232, 10233, 10234, 10237, 10238, 10239, 10240, 10241, 10242, 10247, 10248, 10259, 10264, 10265, 10266, 10267, 10268, 10269, 10270, 10271, 10272, 10273, 10278, 10279, 1028, 10280, 10281, 10282, 10283, 10287, 10288, 10289, 1029, 10290, 10291, 10292, 10293, 10294, 10295, 10296, 10299, 10300, 10301, 10306, 10307, 10308, 10311, 10314, 10315, 10316, 10317, 10318, 10321, 10324, 10325, 10326, 10327, 10328, 10329, 10330, 10331, 10332, 10333, 10334, 10337, 10338, 10339, 10340, 10341, 10344, 10354, 10357, 10360, 10367, 10375, 10381, 10388, 10391, 10399, 10402, 10406, 10409, 10412, 10415, 10419, 10422, 10425, 10428, 10431, 10432, 10437, 10438, 10439, 10440, 10441, 10444, 10445, 10450, 10451, 10455, 10456, 10465, 10466, 10479, 10497, 10509, 10512, 10515, 10516, 10517, 10518, 10519, 10522, 10525, 10528, 10531, 10534, 10535, 10536, 10539, 10542, 10543, 10544, 10545, 10546, 10547, 10548, 10549, 10550, 10551, 10552, 10553, 10554, 10555, 10556, 10557, 10558, 10559, 10560, 10561, 10562, 10563, 10564, 10565, 10566, 10567, 10568, 10569, 10570, 10571, 10572, 10573, 10577, 10581, 10582, 10583, 10587, 10588, 10589, 10594, 10595, 10596, 10597, 10598, 10602, 10609, 10610, 10621, 10626, 10627, 10629, 10631, 10637, 10638, 10639, 10640, 10642, 10643, 10644, 10645, 10647, 10648, 10649, 10652, 10659, 10662, 10665, 10668, 10671, 10672, 10673, 10674, 10675, 10678, 10681, 10682, 10683, 10684, 10685, 10686, 10687, 10688, 10689, 10690, 10691, 10694, 10695, 10696, 10697, 10698, 10701, 10705, 10707, 10708, 10709, 10710, 10719, 10720, 10730, 10731, 10737, 10738, 10739, 10746, 10747, 10748, 10749, 10750, 10753, 10754, 10764, 10765, 10766, 10767, 10768, 10769, 10770, 10771, 10772, 10773, 10774, 10775, 10776, 10778, 10781, 10784, 10789, 10792, 10796, 10797, 10798, 10799, 10800, 10803, 10806, 10809, 10812, 10815, 10816, 10817, 10820, 10823, 10824, 10825, 10826, 10832, 10833, 10834, 10835, 10836, 10845, 10846, 10857, 10862, 10863, 10864, 10865, 10866, 10867, 10872, 10873, 10874, 10875, 10876, 10879, 10882, 10883, 10884, 10885, 10886, 10887, 10888, 10889, 10890, 10891, 10892, 10895, 10896, 10897, 10898, 10899, 10902, 10909, 10910, 10915, 10916, 10917, 10918, 10919, 10922, 10923, 10928, 10931, 10934, 10935, 10936, 10937, 10938, 10941, 10944, 10947, 10950, 10953, 10954, 10955, 10958, 10961, 10962, 10963, 10964, 10969, 10970, 10981, 10986, 10987, 10988, 10989, 10990, 10991, 10992, 10995, 10998, 10999, 11000, 11001, 11002, 11003, 11004, 11005, 11006, 11007, 11008, 11011, 11012, 11013, 11014, 11015, 11018, 11023, 11024, 11027, 11028, 11029, 11030, 11031, 11034, 11035, 11040, 11041, 11042, 11043, 11044, 11047, 11050, 11053, 11056, 11059, 11062, 11065, 11066, 11067, 11070, 11073, 11074, 11075, 11076, 11077, 11078, 1109, 11095, 11098, 11099, 11100, 11103, 11106, 11107, 11108, 11109, 11110, 11111, 11112, 11113, 11114, 11115, 11116, 11117, 11118, 11119, 11120, 11121, 11122, 11123, 11124, 11127, 11130, 11137, 11138, 11139, 11140, 11141, 11142, 11143, 11144, 11145, 1115, 11152, 11153, 11154, 11155, 11156, 11159, 1116, 11162, 11165, 11168, 11171, 11174, 11177, 11180, 11183, 11184, 11185, 11186, 11187, 11188, 1119, 11205, 11210, 11211, 11212, 11213, 11214, 11215, 11216, 11217, 11218, 11219, 11220, 11222, 11223, 11224, 11225, 11226, 11227, 11228, 11229, 11231, 11232, 11233, 11236, 11239, 11242, 11243, 11244, 11245, 11246, 1125, 11250, 11252, 11257, 11260, 11261, 11262, 11263, 11264, 11265, 11267, 11268, 11269, 11270, 11272, 11277, 11278, 11279, 11280, 11282, 11283, 11284, 11285, 11286, 11288, 11289, 11290, 11291, 11292, 11293, 11294, 11295, 11296, 11297, 11298, 11299, 11302, 11307, 11308, 11309, 11312, 11313, 11314, 11315, 11316, 11317, 1132, 11320, 11321, 11323, 11327, 11328, 11329, 11331, 11335, 11336, 11337, 11338, 11339, 11341, 1136, 1141, 1147, 1154, 1160, 1167, 1174, 1175, 1182, 1189, 1194, 1199, 1206, 1211, 1218, 1222, 1227, 1233, 1240, 1244, 1249, 1256, 1263, 1270, 1277, 1284, 1287, 1290, 1293, 1296, 1299, 1302, 1305, 1308, 1311, 1314, 1317, 1320, 1323, 1326, 1329, 1332, 1335, 1338, 1341, 1344, 1347, 1350, 1353, 1356, 1359, 1362, 1365, 1368, 1371, 1374, 1377, 1380, 1383, 1386, 1389, 1392, 1395, 1398, 1401, 1404, 1407, 1410, 1413, 1416, 1419, 1422, 1425, 1428, 1431, 1434, 1437, 1440, 1443, 1446, 1449, 1452, 1455, 1458, 1461, 1464, 1467, 1470, 1473, 1476, 1479, 1482, 1485, 1537, 1551, 1649, 1703, 1708, 1713, 1721, 1758, 1782, 1783, 1789, 1793, 1794, 1795, 1796, 1797, 1798, 1799, 1805, 1811, 1812, 1813, 1814, 1815, 1816, 1817, 1818, 1819, 1820, 1821, 1822, 1828, 1829, 1830, 1832, 1833, 1834, 1835, 1839, 1840, 1841, 1842, 1843, 1845, 1851, 1857, 1858, 1859, 1860, 1861, 1862, 1863, 1864, 1865, 1866, 1867, 1868, 1869, 1870, 1871, 1872, 1873, 1874, 1875, 1876, 1877, 1878, 1879, 1880, 1881, 1882, 1883, 1884, 1885, 1892, 1899, 1906, 1913, 1919, 1926, 1927, 1928, 1929, 1930, 1931, 1932, 1933, 1934, 1935, 1936, 1937, 1938, 1939, 1940, 1941, 1942, 1943, 1944, 1945, 1946, 1947, 1953, 1957, 1958, 1959, 1960, 1961, 1962, 1963, 1965, 1966, 1967, 1968, 1969, 1970, 1971, 1972, 1973, 1974, 1975, 1976, 1977, 1983, 1989, 1990, 1991, 1992, 1993, 1994, 1995, 1996, 1997, 2003, 2010, 2011, 2012, 2013, 2014, 2015, 2016, 2017, 2018, 2019, 2020, 2021, 2022, 2023, 2024, 2031, 2038, 2045, 2052, 2058, 2064, 2065, 2066, 2067, 2068, 2069, 2070, 2071, 2072, 2073, 2074, 2081, 2086, 2107, 2108, 2110, 2111, 2112, 2113, 2114, 2115, 2117, 2171, 2172, 2230, 2231, 2235, 2239, 2240, 2241, 2242, 2243, 2244, 2245, 2246, 2247, 2248, 2249, 2250, 2251, 2252, 2253, 2254, 2255, 2256, 2257, 2267, 2268, 2269, 2274, 2275, 2277, 2278, 2279, 2280, 2281, 2282, 2283, 2284, 2285, 2286, 2287, 2293, 2299, 2300, 2301, 2302, 2303, 2304, 2305, 2306, 2307, 2308, 2309, 2315, 2321, 2322, 2323, 2324, 2325, 2326, 2327, 2328, 2329, 2330, 2331, 2337, 2338, 2339, 2340, 2341, 2342, 2343, 2344, 2345, 2346, 2347, 2348, 2349, 2350, 2351, 2352, 2353, 2354, 2355, 2356, 2357, 2358, 2359, 2360, 2361, 2362, 2363, 2364, 2365, 2366, 2367, 2368, 2374, 2375, 2376, 2377, 2378, 2379, 2380, 2381, 2382, 2383, 2384, 2390, 2396, 2397, 2398, 2399, 2400, 2401, 2402, 2403, 2404, 2405, 2406, 2412, 2418, 2419, 2420, 2421, 2422, 2423, 2424, 2425, 2426, 2427, 2428, 2429, 2430, 2431, 2432, 2433, 2434, 2435, 2436, 2437, 2441, 2442, 2446, 2450, 2454, 2458, 2462, 2466, 2470, 2474, 2478, 2482, 2488, 2496, 2502, 2508, 2523, 2533, 2537, 2538, 2542, 2546, 2550, 2554, 2561, 2567, 2573, 2604, 2607, 2611, 2615, 2619, 2626, 2632, 2638, 2644, 2650, 2653, 2654, 2658, 2662, 2666, 2670, 2674, 2680, 2688, 2692, 2696, 2700, 2704, 2728, 2729, 2733, 2737, 2741, 2745, 2749, 2753, 2757, 2761, 2765, 2766, 2769, 2772, 2775, 2778, 2781, 2784, 2787, 2790, 2793, 2796, 2866, 2867, 2868, 2869, 2878, 2913, 2914, 2915, 2916, 2917, 2918, 2919, 2920, 2921, 2922, 2923, 2924, 2925, 2926, 2927, 2928, 2929, 2930, 2931, 2932, 2933, 2934, 2935, 2936, 2937, 2988, 3005, 3006, 3007, 3008, 3009, 3020, 3021, 3022, 3023, 3024, 3025, 3026, 3027, 3028, 3029, 3032, 3033, 3034, 3035, 3036, 3037, 3038, 3039, 3040, 3041, 3061, 3064, 3067, 3070, 3073, 3080, 3096, 3097, 3101, 3107, 3114, 3122, 3126, 3130, 3131, 3134, 3135, 3136, 3137, 3140, 3144, 3149, 3155, 3159, 3167, 3168, 3169, 3173, 3178, 3184, 3185, 3189, 3195, 3202, 3210, 3211, 3215, 3221, 3228, 3229, 3232, 3236, 3241, 3247, 3251, 3255, 3259, 3263, 3267, 3273, 3281, 3287, 3293, 3299, 3303, 3307, 3311, 3315, 3322, 3328, 3334, 3340, 3343, 3349, 3355, 3361, 3362, 3363, 3364, 3365, 3366, 3367, 3368, 3369, 3370, 3371, 3372, 3373, 3374, 3375, 3379, 3380, 3381, 3384, 3390, 3398, 3404, 3410, 3416, 3420, 3424, 3428, 3432, 3436, 3440, 3444, 3448, 3452, 3453, 3454, 3458, 3462, 3466, 3470, 3474, 3478, 3482, 3486, 3487, 3490, 3493, 3496, 3499, 3502, 3507, 3510, 3515, 3518, 3521, 3524, 3527, 3530, 3535, 3539, 3542, 3545, 3548, 3551, 3552, 3553, 3557, 3560, 3563, 3566, 3569, 3570, 3571, 3574, 3577, 3580, 3583, 3586, 3589, 3592, 3595, 3598, 3601, 3604, 3607, 3610, 3613, 3616, 3619, 3622, 3625, 3628, 3631, 3634, 3637, 3640, 3643, 3646, 3649, 3652, 3655, 3658, 3661, 3664, 3667, 3670, 3673, 3676, 3679, 3682, 3685, 3688, 3691, 3694, 3697, 3700, 3703, 3706, 3709, 3712, 3715, 3718, 3721, 3724, 3727, 3730, 3733, 3736, 3739, 3742, 3745, 3748, 3751, 3754, 3757, 3760, 3763, 3766, 3769, 3772, 3775, 3778, 3781, 3782, 3783, 3786, 3789, 3792, 3795, 3798, 3801, 3804, 3807, 3810, 3813, 3816, 3819, 3822, 3825, 3828, 3831, 3834, 3837, 3840, 3843, 3846, 3849, 3852, 3855, 3858, 3861, 3864, 3867, 3870, 3873, 3876, 3879, 3882, 3885, 3888, 3891, 3953, 3954, 3955, 3956, 3958, 3964, 4193, 4303, 4308, 4313, 4326, 4327, 4333, 4334, 4411, 4412, 4463, 4464, 4465, 4466, 4467, 4468, 4469, 4470, 4471, 4472, 4473, 4474, 4475, 4476, 4477, 4478, 4479, 4480, 4481, 4482, 4483, 4484, 4485, 4486, 4487, 4488, 4489, 4490, 4491, 4492, 4493, 4494, 4495, 4496, 4497, 4498, 4499, 4500, 4501, 4502, 4503, 4504, 4505, 4506, 4507, 4508, 4509, 4510, 4511, 4512, 4513, 4514, 4515, 4516, 4517, 4518, 4519, 4520, 4521, 4522, 4523, 4524, 4525, 4526, 4527, 4528, 4529, 4530, 4531, 4532, 4533, 4534, 4535, 4536, 4537, 4538, 4539, 4540, 4541, 4542, 4543, 4544, 4545, 4549, 4555, 4562, 4563, 4566, 4570, 4575, 4576, 4577, 4581, 4586, 4592, 4593, 4597, 4603, 4610, 4611, 4612, 4613, 4614, 4615, 4616, 4617, 4618, 4619, 4620, 4621, 4622, 4623, 4624, 4625, 4626, 4627, 4628, 4629, 4630, 4631, 4632, 4633, 4634, 4635, 4636, 4637, 4638, 4639, 4640, 4641, 4642, 4643, 4644, 4645, 4646, 4647, 4648, 4649, 4650, 4651, 4652, 4653, 4656, 4657, 4661, 4667, 467, 4674, 4675, 4678, 4682, 4687, 469, 4693, 4694, 4695, 4696, 4697, 4698, 4699, 4700, 4701, 4702, 4706, 4711, 4717, 4718, 4722, 4728, 4735, 4743, 4744, 4745, 4746, 4747, 4748, 4749, 4750, 4751, 4752, 4753, 4754, 4755, 4756, 4757, 4758, 4759, 4760, 4761, 4762, 4763, 4764, 4765, 4766, 4767, 4768, 4769, 4775, 4776, 4777, 4778, 4779, 4780, 4781, 4782, 4783, 4784, 4789, 4790, 4793, 4794, 4795, 4796, 4799, 4800, 4801, 4802, 4803, 4806, 4809, 4810, 4813, 4814, 4817, 4820, 4823, 4826, 4829, 4832, 4835, 4838, 4841, 4844, 4847, 4850, 4853, 4856, 4859, 4862, 4865, 4868, 4871, 4874, 4877, 4880, 4883, 4886, 4889, 4892, 4895, 4898, 4901, 4904, 4907, 4910, 4913, 4916, 4919, 4922, 4925, 4928, 4931, 4934, 4937, 494, 4940, 4943, 4946, 4949, 4952, 4955, 4958, 4961, 4964, 4967, 4970, 4973, 4976, 4979, 4982, 4985, 4988, 4991, 4994, 4997, 5000, 5003, 5006, 5009, 5012, 5015, 5018, 5021, 5024, 5027, 5030, 5033, 5036, 5039, 5042, 5045, 5046, 5047, 5048, 5049, 5052, 5055, 5058, 5061, 5064, 5065, 5066, 5067, 5068, 5071, 5074, 5077, 5080, 5083, 5086, 5089, 5092, 5095, 5098, 5101, 5104, 5107, 5110, 5111, 5112, 5113, 5114, 5117, 5120, 5123, 5126, 5129, 5132, 5135, 5138, 5141, 5144, 5147, 5150, 5153, 5156, 5159, 5162, 5165, 5166, 5167, 5168, 5169, 5170, 5171, 5172, 5173, 5174, 5175, 5176, 5177, 5178, 5179, 5180, 5181, 5182, 5183, 5184, 5185, 5186, 5187, 5188, 5189, 5190, 5191, 5192, 5193, 5196, 5197, 5198, 5199, 5200, 5201, 5202, 5203, 5204, 5205, 5206, 5207, 5208, 5209, 5210, 5211, 5212, 5213, 528, 5283, 5284, 5285, 5286, 5287, 5288, 5289, 5290, 5291, 5292, 5293, 5294, 5295, 5296, 5297, 5298, 5299, 5300, 5314, 5315, 5316, 5317, 5318, 5319, 5320, 5321, 5322, 5323, 5324, 5363, 5364, 5365, 5366, 5367, 5425, 5426, 5427, 5429, 5430, 5431, 5432, 5433, 5451, 5452, 5453, 5454, 5455, 5456, 5457, 5469, 5474, 5475, 5476, 5477, 5571, 5572, 5573, 5574, 5584, 5585, 5586, 5587, 5602, 5603, 5604, 5605, 5631, 5632, 5640, 5654, 5670, 5683, 5690, 5697, 5707, 5718, 5728, 5735, 5736, 5740, 5744, 5747, 575, 5751, 5755, 5758, 5762, 5766, 5769, 5770, 5771, 5778, 578, 5789, 5799, 5807, 5821, 5837, 585, 5850, 5856, 5863, 5870, 5881, 5892, 5898, 590, 5905, 5915, 5926, 593, 5936, 5943, 5944, 5945, 5946, 5947, 5948, 5949, 5950, 5951, 5952, 5953, 5954, 5955, 5956, 5957, 5958, 5959, 596, 5960, 5966, 5967, 5968, 5969, 5970, 5971, 5972, 5973, 5974, 5975, 5976, 5977, 5978, 5979, 5980, 5981, 5989, 599, 5990, 5991, 5996, 6000, 6003, 6009, 6014, 6018, 6021, 6022, 6023, 6024, 6025, 6026, 6027, 6028, 6029, 6030, 6031, 6032, 6033, 6034, 6035, 6036, 6037, 6038, 6039, 604, 6040, 6041, 6047, 6052, 6056, 6059, 6060, 6061, 6062, 6063, 6064, 6065, 6066, 6067, 6068, 6069, 6070, 6071, 6072, 6073, 6074, 6075, 6076, 6077, 6078, 6079, 6083, 6087, 609, 6090, 6091, 6092, 6093, 6094, 6095, 6096, 6097, 6098, 6099, 6100, 6101, 6102, 6103, 6104, 6105, 6106, 6107, 6108, 6109, 6110, 6111, 6112, 6113, 6114, 6115, 6116, 6117, 6118, 6119, 6120, 6121, 6122, 6123, 6124, 6125, 6126, 6127, 6131, 6135, 6136, 6137, 614, 6141, 6145, 6148, 6149, 6150, 6151, 6152, 6153, 6154, 6155, 6156, 6157, 6158, 6159, 6160, 6161, 6162, 6163, 6164, 6165, 6166, 6170, 6174, 6177, 6181, 6182, 6183, 6184, 6185, 6186, 6187, 6188, 6189, 6190, 6191, 6192, 6193, 6194, 6195, 6196, 6199, 6202, 6203, 6204, 6207, 6210, 6213, 6214, 6217, 6220, 6223, 6224, 6225, 6226, 6227, 6228, 6229, 6230, 6231, 6232, 6235, 6236, 6239, 6240, 6241, 6242, 6243, 6246, 6249, 625, 6252, 6255, 6256, 6257, 6258, 6259, 6260, 6261, 6262, 6263, 6266, 628, 632, 636, 641, 642, 644, 651, 6540, 6541, 6542, 6543, 6544, 6545, 6546, 6547, 6555, 6556, 6557, 6558, 6559, 6560, 6561, 6569, 657, 6594, 6595, 6596, 6597, 6598, 6599, 660, 6600, 6601, 6602, 6603, 6604, 6605, 6606, 6621, 6622, 6623, 6624, 6625, 6626, 6627, 6628, 6629, 6639, 6640, 6641, 6642, 6643, 6644, 6645, 6646, 6647, 6648, 6649, 6650, 6651, 6652, 6653, 6654, 6655, 6656, 6657, 6658, 6659, 666, 6660, 6661, 6668, 6677, 6678, 6679, 6680, 6681, 6682, 6683, 6684, 6685, 6686, 6687, 6688, 6689, 6690, 6702, 6703, 6704, 6705, 6706, 6707, 6708, 6709, 6710, 6711, 6712, 672, 6729, 673, 6730, 6731, 6732, 6733, 6734, 6735, 6736, 674, 6741, 6742, 6743, 6744, 6751, 6752, 6753, 6754, 6755, 6756, 6757, 6758, 676, 6761, 6762, 6766, 6767, 6768, 6769, 6770, 6771, 6772, 6773, 6774, 6775, 6776, 6777, 6778, 6779, 6780, 6781, 6782, 6783, 6784, 6787, 6788, 6789, 6790, 6791, 6792, 6793, 6794, 6795, 6796, 6797, 6800, 6803, 6806, 6809, 6812, 6815, 6818, 682, 6821, 6824, 6827, 6830, 6833, 6836, 6837, 6838, 6839, 6840, 6841, 6842, 6843, 6844, 6845, 6848, 6849, 6850, 6851, 6852, 6853, 6854, 6855, 6856, 6857, 6858, 6859, 6860, 6861, 6862, 6863, 6864, 6865, 6866, 6867, 6870, 6871, 6872, 6873, 6874, 6875, 6876, 6877, 6878, 6879, 688, 6880, 6881, 6884, 6885, 6886, 6887, 6888, 6889, 689, 6890, 6891, 6892, 6893, 6894, 6901, 6912, 6923, 6929, 6936, 6946, 695, 6957, 6967, 6968, 6969, 6970, 6977, 6988, 6998, 700, 7006, 7020, 7036, 7049, 705, 7055, 7056, 7057, 706, 7060, 7061, 7062, 7063, 7064, 7065, 7066, 7067, 7068, 7073, 7077, 708, 7080, 7086, 7091, 7095, 7098, 7099, 7100, 7103, 7104, 7105, 7106, 7107, 7114, 7125, 7136, 7142, 7149, 715, 7159, 7170, 7180, 7187, 7188, 7191, 7194, 7198, 7202, 7205, 7209, 721, 7213, 7216, 7219, 7222, 7229, 7240, 7250, 7258, 727, 7272, 7288, 7301, 7307, 7314, 7318, 7322, 7325, 7328, 733, 7331, 7334, 7337, 734, 7340, 7343, 7346, 7351, 7355, 7358, 7364, 7369, 7373, 7376, 7377, 7378, 7381, 7384, 7387, 7391, 7394, 7398, 7402, 7405, 7408, 7411, 7414, 7417, 742, 7420, 7423, 7426, 7429, 7432, 7435, 7438, 7441, 7444, 7447, 7450, 7453, 7456, 7459, 7462, 7465, 7468, 7471, 7474, 7477, 7478, 7479, 748, 7482, 7485, 7488, 749, 7491, 7494, 7497, 750, 7500, 7503, 7506, 7509, 7512, 7515, 7518, 7521, 7524, 7527, 7530, 7533, 7536, 7539, 7542, 7545, 7548, 7551, 7552, 7553, 7556, 7557, 7558, 7559, 7560, 7563, 7566, 7569, 7572, 7573, 7574, 7577, 758, 7580, 7581, 7582, 7585, 7588, 759, 7591, 7609, 7613, 762, 7620, 7649, 7650, 7655, 7659, 7668, 7671, 768, 774, 7744, 780, 7822, 7825, 7826, 7852, 786, 794, 800, 806, 8114, 8117, 812, 8131, 8134, 814, 8144, 8145, 8146, 8156, 8166, 8169, 8183, 8186, 8196, 8200, 8204, 8208, 821, 8216, 8217, 8218, 8219, 8232, 8233, 8242, 8243, 8244, 8245, 8246, 8247, 8248, 8249, 8250, 8251, 8252, 8253, 8254, 8260, 8261, 8262, 8269, 827, 8274, 8275, 8276, 8277, 8278, 8279, 8280, 8281, 8282, 8283, 8284, 8285, 8288, 8294, 8295, 8296, 8297, 8298, 8307, 8315, 8317, 8319, 8321, 8322, 8323, 8324, 8325, 8326, 833, 8333, 8337, 8338, 8339, 8340, 8341, 8342, 8343, 8344, 8345, 8346, 8347, 8348, 8349, 8350, 8351, 8352, 8353, 8354, 8355, 8356, 8357, 8358, 8365, 8369, 8370, 8371, 8372, 8373, 8374, 8375, 8376, 8377, 8378, 8379, 8380, 8381, 8382, 8383, 8384, 8385, 8386, 8387, 8388, 8389, 839, 8390, 8391, 8392, 8393, 8394, 8404, 8405, 8409, 8410, 8411, 8412, 8415, 8416, 8417, 8418, 8421, 8430, 8433, 8434, 8435, 8436, 8437, 8438, 8439, 8440, 8441, 8442, 8443, 8444, 8447, 8448, 8449, 845, 8450, 8451, 8452, 8453, 8454, 8455, 8456, 8457, 8460, 8463, 8466, 8469, 8470, 8471, 8474, 8477, 8480, 8483, 8484, 8485, 8488, 8489, 8490, 8491, 8492, 8493, 8494, 8495, 8496, 8497, 8500, 8501, 8502, 8503, 8504, 8505, 8506, 8507, 8508, 8509, 8510, 8511, 8512, 8513, 8514, 8515, 8516, 8517, 8518, 8519, 8522, 8525, 8528, 853, 8531, 8534, 8537, 8538, 8539, 8540, 8541, 8545, 8546, 8547, 8548, 8551, 8552, 8553, 8554, 8555, 8558, 8561, 8564, 8565, 8566, 8569, 8572, 8575, 8578, 8579, 8580, 8583, 8586, 8589, 859, 8592, 8595, 8598, 8601, 8604, 8607, 8608, 8609, 8610, 8615, 8616, 8617, 8618, 8619, 8624, 8625, 8626, 8627, 8632, 8633, 8634, 8637, 8638, 8639, 8644, 8645, 8646, 8647, 8648, 865, 8653, 8654, 8655, 8660, 8663, 8666, 8669, 8672, 8675, 8678, 8681, 8684, 8687, 8690, 8693, 8696, 8699, 8702, 8705, 8708, 871, 8711, 8714, 8717, 8718, 8721, 8724, 8727, 8730, 8733, 8734, 8735, 8738, 8741, 8744, 8747, 8750, 8753, 8754, 8755, 8756, 8757, 8760, 8763, 8766, 8769, 8772, 8775, 8778, 8781, 8784, 8787, 8790, 8793, 8796, 8799, 8802, 8805, 8808, 8811, 8814, 8815, 8816, 8817, 8818, 8840, 8857, 886, 8861, 8862, 8863, 8864, 8865, 8866, 887, 8871, 8874, 8878, 8879, 8880, 8881, 8882, 8883, 8884, 8885, 8886, 8887, 8888, 8898, 8902, 8920, 8924, 8927, 8931, 8943, 8950, 8956, 8959, 8960, 8963, 8966, 8991, 8992, 8995, 8996, 9001, 9005, 9024, 9025, 9029, 9035, 9053, 9054, 9064, 9065, 9066, 9067, 9068, 9071, 9072, 9073, 9074, 9077, 9079, 9082, 9083, 9086, 9087, 9088, 9089, 9092, 9093, 9094, 9095, 9098, 9099, 9103, 9107, 9111, 9117, 9127, 9146, 9149, 9159, 9160, 9161, 9165, 9169, 9173, 9179, 9180, 9181, 9182, 9183, 9193, 9203, 9206, 9220, 9223, 9234, 9235, 9236, 9237, 9238, 9242, 9243, 9244, 9245, 9246, 9247, 9248, 9249, 9250, 9251, 9252, 9256, 9257, 9258, 9259, 9260, 9261, 9262, 9265, 9268, 9271, 9272, 9273, 9274, 9275, 9276, 9280, 9285, 9286, 9287, 9288, 9290, 9292, 9294, 9296, 9297, 9298, 9299, 9300, 9301, 9307, 9314, 9315, 9318, 9319, 9320, 9321, 9322, 9323, 9324, 9326, 9332, 9339, 9344, 9352, 9354, 9356, 9358, 9359, 9360, 9361, 9362, 9363, 9364, 9365, 9366, 9367, 9368, 9369, 9370, 9371, 9372, 9375, 9381, 9382, 9383, 9384, 9385, 9392, 9393, 9394, 9395, 9396, 9397, 9398, 9399, 9400, 9401, 9402, 9407, 9408, 9412, 9413, 9414, 9415, 9416, 9417, 9418, 9419, 9420, 9421, 9422, 9423, 9426, 9429, 9432, 9435, 9442, 9445, 9454, 9455, 9456, 9459, 9460, 9461, 9462, 9465, 9466, 9467, 9468, 9473, 9476, 9477, 9478, 9485, 9488, 9493, 9494, 9495, 9498, 9499, 9500, 9505, 9506, 9507, 9508, 9509, 9514, 9515, 9516, 9517, 9520, 9526, 9531, 9539, 9540, 9541, 9543, 9551, 9555, 9556, 9557, 9560, 9561, 9562, 9563, 9564, 9565, 9566, 9567, 9568, 9569, 957, 9570, 9571, 9575, 9579, 9581, 9582, 9585, 9591, 9592, 9593, 9594, 9595, 9596, 9597, 9598, 9599, 9600, 9601, 9602, 9603, 9604, 9605, 9608, 9611, 9612, 9613, 9614, 9615, 9616, 9617, 9618, 9621, 9622, 9623, 9624, 9626, 9629, 9632, 9635, 9642, 9645, 9646, 9649, 9650, 9653, 9656, 9659, 9660, 9661, 9662, 9663, 9666, 9667, 9670, 9671, 9674, 9675, 9678, 9679, 9682, 9685, 9690, 9691, 9692, 9695, 9698, 9702, 9707, 9710, 9711, 9714, 9715, 9716, 9717, 9720, 9721, 9722, 9723, 9726, 9727, 9732, 9733, 9734, 9735, 9736, 9737, 9738, 9739, 9740, 9741, 9742, 9754, 9758, 9762, 9763, 9764, 9765, 9766, 9767, 9768, 9769, 9773, 9774, 9775, 9779, 9784, 9785, 9786, 9790, 9791, 9795, 9796, 9797, 9798, 9799, 9800, 9801, 9802, 9803, 9805, 9806, 9809, 9813, 9814, 9815, 9816, 9817, 9820, 9825, 9826, 9827, 9828, 9829, 9830, 9835, 9836, 9837, 9838, 9846, 9847, 9862, 9863, 9866, 9873, 9876, 9890, 9891, 9892, 9893, 9894, 9895, 9896, 9897, 9898, 9899, 9900, 9901, 9902, 9903, 9904, 9905, 9906, 9907, 9908, 9909, 9910, 9911, 9917, 9923, 9924, 9925, 9932, 9935, 9938, 9939, 9945, 9946, 9947, 9948, 9949, 9953, 9954, 9955, 9956, 9957, 9958, 9959, 9960, 9961, 9964, 9967, 9968, 9969, 9970, 9971, 9972, 9973, 9974, 9975, 9976, 9977, 9978, 9979, 9982, 9983, 9986, 9989, 9992, 9995, 9996, 9997, 9998, 9999, 10711_in, flip_signal;

  not ginst1 (10002, 9717);
  nand ginst2 (10003, 9722, 9876);
  not ginst3 (10006, 9723);
  nand ginst4 (10007, 9830, 9829);
  nand ginst5 (10010, 9828, 9827);
  and ginst6 (10013, 9791, 8307, 8269);
  and ginst7 (10014, 9758, 9344, 8307, 8269);
  and ginst8 (10015, 367, 9754, 9344, 8307, 8269);
  and ginst9 (10016, 9786, 8394, 8421);
  and ginst10 (10017, 9820, 9332, 8394, 8421);
  and ginst11 (10018, 9786, 8394, 8421);
  and ginst12 (10019, 9820, 9332, 8394, 8421);
  and ginst13 (10020, 9809, 8298, 8262);
  and ginst14 (10021, 9779, 9385, 8298, 8262);
  and ginst15 (10022, 367, 9775, 9385, 8298, 8262);
  not ginst16 (10023, 9945);
  not ginst17 (10024, 9946);
  nand ginst18 (10025, 9740, 9893);
  not ginst19 (10026, 9923);
  not ginst20 (10028, 9924);
  nand ginst21 (10032, 8595, 9897);
  nand ginst22 (10033, 8598, 9899);
  nand ginst23 (10034, 8601, 9901);
  nand ginst24 (10035, 8604, 9903);
  nand ginst25 (10036, 4803, 9906);
  nand ginst26 (10037, 4806, 9908);
  nand ginst27 (10038, 8627, 9910);
  and ginst28 (10039, 9809, 8298);
  and ginst29 (10040, 9779, 9385, 8298);
  and ginst30 (10041, 367, 9775, 9385, 8298);
  and ginst31 (10042, 9779, 9385);
  and ginst32 (10043, 367, 9775, 9385);
  nand ginst33 (10050, 8727, 9938);
  not ginst34 (10053, 9817);
  and ginst35 (10054, 9817, 9029);
  and ginst36 (10055, 9786, 8394);
  and ginst37 (10056, 9820, 9332, 8394);
  and ginst38 (10057, 9791, 8307);
  and ginst39 (10058, 9758, 9344, 8307);
  and ginst40 (10059, 367, 9754, 9344, 8307);
  and ginst41 (10060, 9758, 9344);
  and ginst42 (10061, 367, 9754, 9344);
  nand ginst43 (10062, 4997, 9947);
  nand ginst44 (10067, 8811, 9953);
  nand ginst45 (10070, 9955, 9836);
  nand ginst46 (10073, 9956, 9838);
  nand ginst47 (10076, 9068, 9957);
  nand ginst48 (10077, 9074, 9959);
  nand ginst49 (10082, 9089, 9967);
  nand ginst50 (10083, 9095, 9969);
  nand ginst51 (10084, 4871, 9971);
  nand ginst52 (10085, 6214, 9973);
  nand ginst53 (10086, 6217, 9975);
  nand ginst54 (10093, 5027, 9995);
  nand ginst55 (10094, 6232, 9997);
  or ginst56 (10101, 9238, 9732, 10013, 10014, 10015);
  or ginst57 (10102, 9339, 9526, 10016, 10017, 9734);
  or ginst58 (10103, 9339, 9531, 10018, 10019, 9735);
  or ginst59 (10104, 9242, 9736, 10020, 10021, 10022);
  and ginst60 (10105, 9925, 9894);
  and ginst61 (10106, 9925, 9895);
  and ginst62 (10107, 9925, 9896);
  and ginst63 (10108, 9925, 8253);
  nand ginst64 (10109, 10032, 9898);
  nand ginst65 (10110, 10033, 9900);
  nand ginst66 (10111, 10034, 9902);
  nand ginst67 (10112, 10035, 9904);
  nand ginst68 (10113, 10036, 9907);
  nand ginst69 (10114, 10037, 9909);
  nand ginst70 (10115, 10038, 9911);
  or ginst71 (10116, 9265, 10039, 10040, 10041);
  or ginst72 (10119, 9809, 10042, 10043);
  not ginst73 (10124, 9925);
  and ginst74 (10130, 9768, 9925);
  not ginst75 (10131, 9932);
  not ginst76 (10132, 9935);
  and ginst77 (10133, 9932, 8920);
  nand ginst78 (10134, 10050, 9939);
  not ginst79 (10135, 9983);
  nand ginst80 (10136, 9983, 9324);
  not ginst81 (10137, 9986);
  nand ginst82 (10138, 9986, 9784);
  and ginst83 (10139, 9785, 10053);
  or ginst84 (10140, 8943, 10055, 10056, 9790);
  or ginst85 (10141, 9268, 10057, 10058, 10059);
  or ginst86 (10148, 9791, 10060, 10061);
  nand ginst87 (10155, 10062, 9948);
  not ginst88 (10156, 9989);
  nand ginst89 (10157, 9989, 9805);
  not ginst90 (10158, 9992);
  nand ginst91 (10159, 9992, 9806);
  not ginst92 (10160, 9949);
  nand ginst93 (10161, 10067, 9954);
  not ginst94 (10162, 10007);
  nand ginst95 (10163, 10007, 9825);
  not ginst96 (10164, 10010);
  nand ginst97 (10165, 10010, 9826);
  nand ginst98 (10170, 10076, 9958);
  nand ginst99 (10173, 10077, 9960);
  not ginst100 (10176, 9961);
  nand ginst101 (10177, 9961, 9082);
  not ginst102 (10178, 9964);
  nand ginst103 (10179, 9964, 9086);
  nand ginst104 (10180, 10082, 9968);
  nand ginst105 (10183, 10083, 9970);
  nand ginst106 (10186, 9972, 10084);
  nand ginst107 (10189, 9974, 10085);
  nand ginst108 (10192, 9976, 10086);
  not ginst109 (10195, 9979);
  nand ginst110 (10196, 9979, 9982);
  nand ginst111 (10197, 9996, 10093);
  nand ginst112 (10200, 9998, 10094);
  not ginst113 (10203, 9999);
  nand ginst114 (10204, 9999, 10002);
  not ginst115 (10205, 10003);
  nand ginst116 (10206, 10003, 10006);
  nand ginst117 (10212, 10070, 4308);
  nand ginst118 (10213, 10073, 4313);
  and ginst119 (10230, 9774, 10131);
  nand ginst120 (10231, 8730, 10135);
  nand ginst121 (10232, 9478, 10137);
  or ginst122 (10233, 10139, 10054);
  nand ginst123 (10234, 7100, 10140);
  nand ginst124 (10237, 9485, 10156);
  nand ginst125 (10238, 9488, 10158);
  nand ginst126 (10239, 9517, 10162);
  nand ginst127 (10240, 9520, 10164);
  not ginst128 (10241, 10070);
  not ginst129 (10242, 10073);
  nand ginst130 (10247, 8146, 10176);
  nand ginst131 (10248, 8156, 10178);
  nand ginst132 (10259, 9692, 10195);
  nand ginst133 (10264, 9717, 10203);
  nand ginst134 (10265, 9723, 10205);
  and ginst135 (10266, 10026, 10124);
  and ginst136 (10267, 10028, 10124);
  and ginst137 (10268, 9742, 10124);
  and ginst138 (10269, 6923, 10124);
  nand ginst139 (10270, 6762, 10116);
  nand ginst140 (10271, 3061, 10241);
  nand ginst141 (10272, 3064, 10242);
  not ginst142 (10273, 10116);
  and ginst143 (10278, 10141, 5728, 5707, 5718, 5697);
  and ginst144 (10279, 10141, 5728, 5707, 5718);
  and ginst145 (1028, 382, 641);
  and ginst146 (10280, 10141, 5728, 5718);
  and ginst147 (10281, 10141, 5728);
  and ginst148 (10282, 6784, 10141);
  not ginst149 (10283, 10119);
  and ginst150 (10287, 10148, 5936, 5915, 5926, 5905);
  and ginst151 (10288, 10148, 5936, 5915, 5926);
  and ginst152 (10289, 10148, 5936, 5926);
  nand ginst153 (1029, 382, 705);
  and ginst154 (10290, 10148, 5936);
  and ginst155 (10291, 6881, 10148);
  and ginst156 (10292, 8898, 10124);
  nand ginst157 (10293, 10231, 10136);
  nand ginst158 (10294, 10232, 10138);
  nand ginst159 (10295, 8412, 10233);
  and ginst160 (10296, 8959, 10234);
  nand ginst161 (10299, 10237, 10157);
  nand ginst162 (10300, 10238, 10159);
  or ginst163 (10301, 10230, 10133);
  nand ginst164 (10306, 10239, 10163);
  nand ginst165 (10307, 10240, 10165);
  not ginst166 (10308, 10148);
  not ginst167 (10311, 10141);
  not ginst168 (10314, 10170);
  nand ginst169 (10315, 10170, 9071);
  not ginst170 (10316, 10173);
  nand ginst171 (10317, 10173, 9077);
  nand ginst172 (10318, 10247, 10177);
  nand ginst173 (10321, 10248, 10179);
  not ginst174 (10324, 10180);
  nand ginst175 (10325, 10180, 9092);
  not ginst176 (10326, 10183);
  nand ginst177 (10327, 10183, 9098);
  not ginst178 (10328, 10186);
  nand ginst179 (10329, 10186, 9674);
  not ginst180 (10330, 10189);
  nand ginst181 (10331, 10189, 9678);
  not ginst182 (10332, 10192);
  nand ginst183 (10333, 10192, 9977);
  nand ginst184 (10334, 10259, 10196);
  not ginst185 (10337, 10197);
  nand ginst186 (10338, 10197, 9710);
  not ginst187 (10339, 10200);
  nand ginst188 (10340, 10200, 9714);
  nand ginst189 (10341, 10264, 10204);
  nand ginst190 (10344, 10265, 10206);
  or ginst191 (10350, 10266, 10105);
  or ginst192 (10351, 10267, 10106);
  or ginst193 (10352, 10268, 10107);
  or ginst194 (10353, 10269, 10108);
  and ginst195 (10354, 8857, 10270);
  nand ginst196 (10357, 10271, 10212);
  nand ginst197 (10360, 10272, 10213);
  or ginst198 (10367, 7620, 10282);
  or ginst199 (10375, 7671, 10291);
  or ginst200 (10381, 10292, 10130);
  and ginst201 (10388, 10114, 10134, 10293, 10294);
  and ginst202 (10391, 9582, 10295);
  and ginst203 (10399, 10113, 10115, 10299, 10300);
  and ginst204 (10402, 10155, 10161, 10306, 10307);
  or ginst205 (10406, 3229, 6888, 6889, 6890, 10287);
  or ginst206 (10409, 3232, 6891, 6892, 10288);
  or ginst207 (10412, 3236, 6893, 10289);
  or ginst208 (10415, 3241, 10290);
  or ginst209 (10419, 3137, 6791, 6792, 6793, 10278);
  or ginst210 (10422, 3140, 6794, 6795, 10279);
  or ginst211 (10425, 3144, 6796, 10280);
  or ginst212 (10428, 3149, 10281);
  nand ginst213 (10431, 8117, 10314);
  nand ginst214 (10432, 8134, 10316);
  nand ginst215 (10437, 8169, 10324);
  nand ginst216 (10438, 8186, 10326);
  nand ginst217 (10439, 9117, 10328);
  nand ginst218 (10440, 9127, 10330);
  nand ginst219 (10441, 9682, 10332);
  nand ginst220 (10444, 9183, 10337);
  nand ginst221 (10445, 9193, 10339);
  not ginst222 (10450, 10296);
  and ginst223 (10451, 10296, 4193);
  not ginst224 (10455, 10308);
  nand ginst225 (10456, 10308, 8242);
  not ginst226 (10465, 10311);
  nand ginst227 (10466, 10311, 8247);
  not ginst228 (10479, 10273);
  not ginst229 (10497, 10301);
  nand ginst230 (10509, 10431, 10315);
  nand ginst231 (10512, 10432, 10317);
  not ginst232 (10515, 10318);
  nand ginst233 (10516, 10318, 8632);
  not ginst234 (10517, 10321);
  nand ginst235 (10518, 10321, 8637);
  nand ginst236 (10519, 10437, 10325);
  nand ginst237 (10522, 10438, 10327);
  nand ginst238 (10525, 10439, 10329);
  nand ginst239 (10528, 10440, 10331);
  nand ginst240 (10531, 10441, 10333);
  not ginst241 (10534, 10334);
  nand ginst242 (10535, 10334, 9695);
  nand ginst243 (10536, 10444, 10338);
  nand ginst244 (10539, 10445, 10340);
  not ginst245 (10542, 10341);
  nand ginst246 (10543, 10341, 9720);
  not ginst247 (10544, 10344);
  nand ginst248 (10545, 10344, 9726);
  and ginst249 (10546, 5631, 10450);
  not ginst250 (10547, 10391);
  and ginst251 (10548, 10391, 8950);
  and ginst252 (10549, 5165, 10367);
  not ginst253 (10550, 10354);
  and ginst254 (10551, 10354, 3126);
  nand ginst255 (10552, 7411, 10455);
  and ginst256 (10553, 10375, 9539);
  and ginst257 (10554, 10375, 9540);
  and ginst258 (10555, 10375, 9541);
  and ginst259 (10556, 10375, 6761);
  not ginst260 (10557, 10406);
  nand ginst261 (10558, 10406, 8243);
  not ginst262 (10559, 10409);
  nand ginst263 (10560, 10409, 8244);
  not ginst264 (10561, 10412);
  nand ginst265 (10562, 10412, 8245);
  not ginst266 (10563, 10415);
  nand ginst267 (10564, 10415, 8246);
  nand ginst268 (10565, 7426, 10465);
  not ginst269 (10566, 10419);
  nand ginst270 (10567, 10419, 8248);
  not ginst271 (10568, 10422);
  nand ginst272 (10569, 10422, 8249);
  not ginst273 (10570, 10425);
  nand ginst274 (10571, 10425, 8250);
  not ginst275 (10572, 10428);
  nand ginst276 (10573, 10428, 8251);
  not ginst277 (10574, 10399);
  not ginst278 (10575, 10402);
  not ginst279 (10576, 10388);
  and ginst280 (10577, 10399, 10402, 10388);
  and ginst281 (10581, 10360, 9543, 10273);
  and ginst282 (10582, 10357, 9905, 10273);
  not ginst283 (10583, 10367);
  and ginst284 (10587, 10367, 5735);
  and ginst285 (10588, 10367, 3135);
  not ginst286 (10589, 10375);
  and ginst287 (10594, 10381, 7180, 7159, 7170, 7149);
  and ginst288 (10595, 10381, 7180, 7159, 7170);
  and ginst289 (10596, 10381, 7180, 7170);
  and ginst290 (10597, 10381, 7180);
  and ginst291 (10598, 8444, 10381);
  not ginst292 (10602, 10381);
  nand ginst293 (10609, 7479, 10515);
  nand ginst294 (10610, 7491, 10517);
  nand ginst295 (10621, 9149, 10534);
  nand ginst296 (10626, 9206, 10542);
  nand ginst297 (10627, 9223, 10544);
  or ginst298 (10628, 10546, 10451);
  and ginst299 (10629, 9733, 10547);
  and ginst300 (10631, 5166, 10550);
  nand ginst301 (10632, 10552, 10456);
  nand ginst302 (10637, 7414, 10557);
  nand ginst303 (10638, 7417, 10559);
  nand ginst304 (10639, 7420, 10561);
  nand ginst305 (10640, 7423, 10563);
  nand ginst306 (10641, 10565, 10466);
  nand ginst307 (10642, 7429, 10566);
  nand ginst308 (10643, 7432, 10568);
  nand ginst309 (10644, 7435, 10570);
  nand ginst310 (10645, 7438, 10572);
  and ginst311 (10647, 886, 887, 10577);
  and ginst312 (10648, 10360, 8857, 10479);
  and ginst313 (10649, 10357, 7609, 10479);
  or ginst314 (10652, 8966, 10598);
  or ginst315 (10659, 4675, 8451, 8452, 8453, 10594);
  or ginst316 (10662, 4678, 8454, 8455, 10595);
  or ginst317 (10665, 4682, 8456, 10596);
  or ginst318 (10668, 4687, 10597);
  not ginst319 (10671, 10509);
  nand ginst320 (10672, 10509, 8615);
  not ginst321 (10673, 10512);
  nand ginst322 (10674, 10512, 8624);
  nand ginst323 (10675, 10609, 10516);
  nand ginst324 (10678, 10610, 10518);
  not ginst325 (10681, 10519);
  nand ginst326 (10682, 10519, 8644);
  not ginst327 (10683, 10522);
  nand ginst328 (10684, 10522, 8653);
  not ginst329 (10685, 10525);
  nand ginst330 (10686, 10525, 9454);
  not ginst331 (10687, 10528);
  nand ginst332 (10688, 10528, 9459);
  not ginst333 (10689, 10531);
  nand ginst334 (10690, 10531, 9978);
  nand ginst335 (10691, 10621, 10535);
  not ginst336 (10694, 10536);
  nand ginst337 (10695, 10536, 9493);
  not ginst338 (10696, 10539);
  nand ginst339 (10697, 10539, 9498);
  nand ginst340 (10698, 10626, 10543);
  nand ginst341 (10701, 10627, 10545);
  or ginst342 (10704, 10629, 10548);
  and ginst343 (10705, 3159, 10583);
  or ginst344 (10706, 10631, 10551);
  and ginst345 (10707, 9737, 10589);
  and ginst346 (10708, 9738, 10589);
  and ginst347 (10709, 9243, 10589);
  and ginst348 (10710, 5892, 10589);
  xor ginst349 (10711, 10711_in, flip_signal);
  nand ginst350 (10711_in, 10637, 10558);
  nand ginst351 (10712, 10638, 10560);
  nand ginst352 (10713, 10639, 10562);
  nand ginst353 (10714, 10640, 10564);
  nand ginst354 (10715, 10642, 10567);
  nand ginst355 (10716, 10643, 10569);
  nand ginst356 (10717, 10644, 10571);
  nand ginst357 (10718, 10645, 10573);
  not ginst358 (10719, 10602);
  nand ginst359 (10720, 10602, 9244);
  not ginst360 (10729, 10647);
  and ginst361 (10730, 5178, 10583);
  and ginst362 (10731, 2533, 10583);
  nand ginst363 (10737, 7447, 10671);
  nand ginst364 (10738, 7465, 10673);
  or ginst365 (10739, 10648, 10649, 10581, 10582);
  nand ginst366 (10746, 7503, 10681);
  nand ginst367 (10747, 7521, 10683);
  nand ginst368 (10748, 8678, 10685);
  nand ginst369 (10749, 8690, 10687);
  nand ginst370 (10750, 9685, 10689);
  nand ginst371 (10753, 8757, 10694);
  nand ginst372 (10754, 8769, 10696);
  or ginst373 (10759, 10705, 10549);
  or ginst374 (10760, 10707, 10553);
  or ginst375 (10761, 10708, 10554);
  or ginst376 (10762, 10709, 10555);
  or ginst377 (10763, 10710, 10556);
  nand ginst378 (10764, 8580, 10719);
  and ginst379 (10765, 10652, 9890);
  and ginst380 (10766, 10652, 9891);
  and ginst381 (10767, 10652, 9892);
  and ginst382 (10768, 10652, 8252);
  not ginst383 (10769, 10659);
  nand ginst384 (10770, 10659, 9245);
  not ginst385 (10771, 10662);
  nand ginst386 (10772, 10662, 9246);
  not ginst387 (10773, 10665);
  nand ginst388 (10774, 10665, 9247);
  not ginst389 (10775, 10668);
  nand ginst390 (10776, 10668, 9248);
  or ginst391 (10778, 10730, 10587);
  or ginst392 (10781, 10731, 10588);
  not ginst393 (10784, 10652);
  nand ginst394 (10789, 10737, 10672);
  nand ginst395 (10792, 10738, 10674);
  not ginst396 (10796, 10675);
  nand ginst397 (10797, 10675, 8633);
  not ginst398 (10798, 10678);
  nand ginst399 (10799, 10678, 8638);
  nand ginst400 (10800, 10746, 10682);
  nand ginst401 (10803, 10747, 10684);
  nand ginst402 (10806, 10748, 10686);
  nand ginst403 (10809, 10749, 10688);
  nand ginst404 (10812, 10750, 10690);
  not ginst405 (10815, 10691);
  nand ginst406 (10816, 10691, 9866);
  nand ginst407 (10817, 10753, 10695);
  nand ginst408 (10820, 10754, 10697);
  not ginst409 (10823, 10698);
  nand ginst410 (10824, 10698, 9505);
  not ginst411 (10825, 10701);
  nand ginst412 (10826, 10701, 9514);
  nand ginst413 (10827, 10764, 10720);
  nand ginst414 (10832, 8583, 10769);
  nand ginst415 (10833, 8586, 10771);
  nand ginst416 (10834, 8589, 10773);
  nand ginst417 (10835, 8592, 10775);
  not ginst418 (10836, 10739);
  not ginst419 (10837, 10778);
  not ginst420 (10838, 10778);
  not ginst421 (10839, 10781);
  not ginst422 (10840, 10781);
  nand ginst423 (10845, 7482, 10796);
  nand ginst424 (10846, 7494, 10798);
  nand ginst425 (10857, 9473, 10815);
  nand ginst426 (10862, 8781, 10823);
  nand ginst427 (10863, 8799, 10825);
  and ginst428 (10864, 10023, 10784);
  and ginst429 (10865, 10024, 10784);
  and ginst430 (10866, 9739, 10784);
  and ginst431 (10867, 7136, 10784);
  nand ginst432 (10868, 10832, 10770);
  nand ginst433 (10869, 10833, 10772);
  nand ginst434 (10870, 10834, 10774);
  nand ginst435 (10871, 10835, 10776);
  not ginst436 (10872, 10789);
  nand ginst437 (10873, 10789, 8616);
  not ginst438 (10874, 10792);
  nand ginst439 (10875, 10792, 8625);
  nand ginst440 (10876, 10845, 10797);
  nand ginst441 (10879, 10846, 10799);
  not ginst442 (10882, 10800);
  nand ginst443 (10883, 10800, 8645);
  not ginst444 (10884, 10803);
  nand ginst445 (10885, 10803, 8654);
  not ginst446 (10886, 10806);
  nand ginst447 (10887, 10806, 9455);
  not ginst448 (10888, 10809);
  nand ginst449 (10889, 10809, 9460);
  not ginst450 (10890, 10812);
  nand ginst451 (10891, 10812, 9862);
  nand ginst452 (10892, 10857, 10816);
  not ginst453 (10895, 10817);
  nand ginst454 (10896, 10817, 9494);
  not ginst455 (10897, 10820);
  nand ginst456 (10898, 10820, 9499);
  nand ginst457 (10899, 10862, 10824);
  nand ginst458 (10902, 10863, 10826);
  or ginst459 (10905, 10864, 10765);
  or ginst460 (10906, 10865, 10766);
  or ginst461 (10907, 10866, 10767);
  or ginst462 (10908, 10867, 10768);
  nand ginst463 (10909, 7450, 10872);
  nand ginst464 (10910, 7468, 10874);
  nand ginst465 (10915, 7506, 10882);
  nand ginst466 (10916, 7524, 10884);
  nand ginst467 (10917, 8681, 10886);
  nand ginst468 (10918, 8693, 10888);
  nand ginst469 (10919, 9462, 10890);
  nand ginst470 (10922, 8760, 10895);
  nand ginst471 (10923, 8772, 10897);
  nand ginst472 (10928, 10909, 10873);
  nand ginst473 (10931, 10910, 10875);
  not ginst474 (10934, 10876);
  nand ginst475 (10935, 10876, 8634);
  not ginst476 (10936, 10879);
  nand ginst477 (10937, 10879, 8639);
  nand ginst478 (10938, 10915, 10883);
  nand ginst479 (10941, 10916, 10885);
  nand ginst480 (10944, 10917, 10887);
  nand ginst481 (10947, 10918, 10889);
  nand ginst482 (10950, 10919, 10891);
  not ginst483 (10953, 10892);
  nand ginst484 (10954, 10892, 9476);
  nand ginst485 (10955, 10922, 10896);
  nand ginst486 (10958, 10923, 10898);
  not ginst487 (10961, 10899);
  nand ginst488 (10962, 10899, 9506);
  not ginst489 (10963, 10902);
  nand ginst490 (10964, 10902, 9515);
  nand ginst491 (10969, 7485, 10934);
  nand ginst492 (10970, 7497, 10936);
  nand ginst493 (10981, 8718, 10953);
  nand ginst494 (10986, 8784, 10961);
  nand ginst495 (10987, 8802, 10963);
  not ginst496 (10988, 10928);
  nand ginst497 (10989, 10928, 8617);
  not ginst498 (10990, 10931);
  nand ginst499 (10991, 10931, 8626);
  nand ginst500 (10992, 10969, 10935);
  nand ginst501 (10995, 10970, 10937);
  not ginst502 (10998, 10938);
  nand ginst503 (10999, 10938, 8646);
  not ginst504 (11000, 10941);
  nand ginst505 (11001, 10941, 8655);
  not ginst506 (11002, 10944);
  nand ginst507 (11003, 10944, 9456);
  not ginst508 (11004, 10947);
  nand ginst509 (11005, 10947, 9461);
  not ginst510 (11006, 10950);
  nand ginst511 (11007, 10950, 9465);
  nand ginst512 (11008, 10981, 10954);
  not ginst513 (11011, 10955);
  nand ginst514 (11012, 10955, 9495);
  not ginst515 (11013, 10958);
  nand ginst516 (11014, 10958, 9500);
  nand ginst517 (11015, 10986, 10962);
  nand ginst518 (11018, 10987, 10964);
  nand ginst519 (11023, 7453, 10988);
  nand ginst520 (11024, 7471, 10990);
  nand ginst521 (11027, 7509, 10998);
  nand ginst522 (11028, 7527, 11000);
  nand ginst523 (11029, 8684, 11002);
  nand ginst524 (11030, 8696, 11004);
  nand ginst525 (11031, 8702, 11006);
  nand ginst526 (11034, 8763, 11011);
  nand ginst527 (11035, 8775, 11013);
  not ginst528 (11040, 10992);
  nand ginst529 (11041, 10992, 8294);
  not ginst530 (11042, 10995);
  nand ginst531 (11043, 10995, 8295);
  nand ginst532 (11044, 11023, 10989);
  nand ginst533 (11047, 11024, 10991);
  nand ginst534 (11050, 11027, 10999);
  nand ginst535 (11053, 11028, 11001);
  nand ginst536 (11056, 11029, 11003);
  nand ginst537 (11059, 11030, 11005);
  nand ginst538 (11062, 11031, 11007);
  not ginst539 (11065, 11008);
  nand ginst540 (11066, 11008, 9477);
  nand ginst541 (11067, 11034, 11012);
  nand ginst542 (11070, 11035, 11014);
  not ginst543 (11073, 11015);
  nand ginst544 (11074, 11015, 9507);
  not ginst545 (11075, 11018);
  nand ginst546 (11076, 11018, 9516);
  nand ginst547 (11077, 7488, 11040);
  nand ginst548 (11078, 7500, 11042);
  and ginst549 (1109, 469, 596);
  nand ginst550 (11095, 8721, 11065);
  nand ginst551 (11098, 8787, 11073);
  nand ginst552 (11099, 8805, 11075);
  nand ginst553 (1110, 242, 593);
  nand ginst554 (11100, 11077, 11041);
  nand ginst555 (11103, 11078, 11043);
  not ginst556 (11106, 11056);
  nand ginst557 (11107, 11056, 9319);
  not ginst558 (11108, 11059);
  nand ginst559 (11109, 11059, 9320);
  not ginst560 (1111, 625);
  not ginst561 (11110, 11067);
  nand ginst562 (11111, 11067, 9381);
  not ginst563 (11112, 11070);
  nand ginst564 (11113, 11070, 9382);
  not ginst565 (11114, 11044);
  nand ginst566 (11115, 11044, 8618);
  not ginst567 (11116, 11047);
  nand ginst568 (11117, 11047, 8619);
  not ginst569 (11118, 11050);
  nand ginst570 (11119, 11050, 8647);
  nand ginst571 (1112, 242, 593);
  not ginst572 (11120, 11053);
  nand ginst573 (11121, 11053, 8648);
  not ginst574 (11122, 11062);
  nand ginst575 (11123, 11062, 9466);
  nand ginst576 (11124, 11095, 11066);
  nand ginst577 (11127, 11098, 11074);
  nand ginst578 (1113, 469, 596);
  nand ginst579 (11130, 11099, 11076);
  nand ginst580 (11137, 8687, 11106);
  nand ginst581 (11138, 8699, 11108);
  nand ginst582 (11139, 8766, 11110);
  not ginst583 (1114, 625);
  nand ginst584 (11140, 8778, 11112);
  nand ginst585 (11141, 7456, 11114);
  nand ginst586 (11142, 7474, 11116);
  nand ginst587 (11143, 7512, 11118);
  nand ginst588 (11144, 7530, 11120);
  nand ginst589 (11145, 8705, 11122);
  not ginst590 (1115, 871);
  and ginst591 (11152, 11103, 8871, 10283);
  and ginst592 (11153, 11100, 7655, 10283);
  and ginst593 (11154, 11103, 9551, 10119);
  and ginst594 (11155, 11100, 9917, 10119);
  nand ginst595 (11156, 11137, 11107);
  nand ginst596 (11159, 11138, 11109);
  not ginst597 (1116, 590);
  nand ginst598 (11162, 11139, 11111);
  nand ginst599 (11165, 11140, 11113);
  nand ginst600 (11168, 11141, 11115);
  nand ginst601 (11171, 11142, 11117);
  nand ginst602 (11174, 11143, 11119);
  nand ginst603 (11177, 11144, 11121);
  nand ginst604 (11180, 11145, 11123);
  not ginst605 (11183, 11124);
  nand ginst606 (11184, 11124, 9468);
  not ginst607 (11185, 11127);
  nand ginst608 (11186, 11127, 9508);
  not ginst609 (11187, 11130);
  nand ginst610 (11188, 11130, 9509);
  not ginst611 (1119, 628);
  or ginst612 (11205, 11152, 11153, 11154, 11155);
  nand ginst613 (11210, 8724, 11183);
  nand ginst614 (11211, 8790, 11185);
  nand ginst615 (11212, 8808, 11187);
  not ginst616 (11213, 11168);
  nand ginst617 (11214, 11168, 8260);
  not ginst618 (11215, 11171);
  nand ginst619 (11216, 11171, 8261);
  not ginst620 (11217, 11174);
  nand ginst621 (11218, 11174, 8296);
  not ginst622 (11219, 11177);
  nand ginst623 (11220, 11177, 8297);
  and ginst624 (11222, 11159, 9575, 1218);
  and ginst625 (11223, 11156, 8927, 1218);
  and ginst626 (11224, 11159, 9935, 750);
  and ginst627 (11225, 11156, 10132, 750);
  and ginst628 (11226, 11165, 9608, 10497);
  and ginst629 (11227, 11162, 9001, 10497);
  and ginst630 (11228, 11165, 9949, 10301);
  and ginst631 (11229, 11162, 10160, 10301);
  not ginst632 (11231, 11180);
  nand ginst633 (11232, 11180, 9467);
  nand ginst634 (11233, 11210, 11184);
  nand ginst635 (11236, 11211, 11186);
  nand ginst636 (11239, 11212, 11188);
  nand ginst637 (11242, 7459, 11213);
  nand ginst638 (11243, 7462, 11215);
  nand ginst639 (11244, 7515, 11217);
  nand ginst640 (11245, 7518, 11219);
  not ginst641 (11246, 11205);
  not ginst642 (1125, 682);
  nand ginst643 (11250, 8708, 11231);
  or ginst644 (11252, 11222, 11223, 11224, 11225);
  or ginst645 (11257, 11226, 11227, 11228, 11229);
  nand ginst646 (11260, 11242, 11214);
  nand ginst647 (11261, 11243, 11216);
  nand ginst648 (11262, 11244, 11218);
  nand ginst649 (11263, 11245, 11220);
  not ginst650 (11264, 11233);
  nand ginst651 (11265, 11233, 9322);
  not ginst652 (11267, 11236);
  nand ginst653 (11268, 11236, 9383);
  not ginst654 (11269, 11239);
  nand ginst655 (11270, 11239, 9384);
  nand ginst656 (11272, 11250, 11232);
  not ginst657 (11277, 11261);
  and ginst658 (11278, 10273, 11260);
  not ginst659 (11279, 11263);
  and ginst660 (11280, 10119, 11262);
  nand ginst661 (11282, 8714, 11264);
  not ginst662 (11283, 11252);
  nand ginst663 (11284, 8793, 11267);
  nand ginst664 (11285, 8796, 11269);
  not ginst665 (11286, 11257);
  and ginst666 (11288, 11277, 10479);
  and ginst667 (11289, 11279, 10283);
  not ginst668 (11290, 11272);
  nand ginst669 (11291, 11272, 9321);
  nand ginst670 (11292, 11282, 11265);
  nand ginst671 (11293, 11284, 11268);
  nand ginst672 (11294, 11285, 11270);
  nand ginst673 (11295, 8711, 11290);
  not ginst674 (11296, 11292);
  not ginst675 (11297, 11294);
  and ginst676 (11298, 10301, 11293);
  or ginst677 (11299, 11288, 11278);
  or ginst678 (11302, 11289, 11280);
  nand ginst679 (11307, 11295, 11291);
  and ginst680 (11308, 11296, 1218);
  and ginst681 (11309, 11297, 10497);
  nand ginst682 (11312, 11302, 11246);
  nand ginst683 (11313, 11299, 10836);
  not ginst684 (11314, 11299);
  not ginst685 (11315, 11302);
  and ginst686 (11316, 750, 11307);
  or ginst687 (11317, 11309, 11298);
  not ginst688 (1132, 628);
  nand ginst689 (11320, 11205, 11315);
  nand ginst690 (11321, 10739, 11314);
  or ginst691 (11323, 11308, 11316);
  nand ginst692 (11327, 11312, 11320);
  nand ginst693 (11328, 11313, 11321);
  nand ginst694 (11329, 11317, 11286);
  not ginst695 (11331, 11317);
  not ginst696 (11333, 11327);
  not ginst697 (11334, 11328);
  nand ginst698 (11335, 11257, 11331);
  nand ginst699 (11336, 11323, 11283);
  not ginst700 (11337, 11323);
  nand ginst701 (11338, 11329, 11335);
  nand ginst702 (11339, 11252, 11337);
  not ginst703 (11340, 11338);
  nand ginst704 (11341, 11336, 11339);
  not ginst705 (11342, 11341);
  not ginst706 (1136, 682);
  not ginst707 (1141, 628);
  not ginst708 (1147, 682);
  not ginst709 (1154, 632);
  not ginst710 (1160, 676);
  and ginst711 (1167, 700, 614);
  and ginst712 (1174, 700, 614);
  not ginst713 (1175, 682);
  not ginst714 (1182, 676);
  not ginst715 (1189, 657);
  not ginst716 (1194, 676);
  not ginst717 (1199, 682);
  not ginst718 (1206, 689);
  not ginst719 (1211, 695);
  not ginst720 (1218, 750);
  not ginst721 (1222, 1028);
  not ginst722 (1227, 632);
  not ginst723 (1233, 676);
  not ginst724 (1240, 632);
  not ginst725 (1244, 676);
  not ginst726 (1249, 689);
  not ginst727 (1256, 689);
  not ginst728 (1263, 695);
  not ginst729 (1270, 689);
  not ginst730 (1277, 689);
  not ginst731 (1284, 700);
  not ginst732 (1287, 614);
  not ginst733 (1290, 666);
  not ginst734 (1293, 660);
  not ginst735 (1296, 651);
  not ginst736 (1299, 614);
  not ginst737 (1302, 644);
  not ginst738 (1305, 700);
  not ginst739 (1308, 614);
  not ginst740 (1311, 614);
  not ginst741 (1314, 666);
  not ginst742 (1317, 660);
  not ginst743 (1320, 651);
  not ginst744 (1323, 644);
  not ginst745 (1326, 609);
  not ginst746 (1329, 604);
  not ginst747 (1332, 742);
  not ginst748 (1335, 599);
  not ginst749 (1338, 727);
  not ginst750 (1341, 721);
  not ginst751 (1344, 715);
  not ginst752 (1347, 734);
  not ginst753 (1350, 708);
  not ginst754 (1353, 609);
  not ginst755 (1356, 604);
  not ginst756 (1359, 742);
  not ginst757 (1362, 734);
  not ginst758 (1365, 599);
  not ginst759 (1368, 727);
  not ginst760 (1371, 721);
  not ginst761 (1374, 715);
  not ginst762 (1377, 708);
  not ginst763 (1380, 806);
  not ginst764 (1383, 800);
  not ginst765 (1386, 794);
  not ginst766 (1389, 786);
  not ginst767 (1392, 780);
  not ginst768 (1395, 774);
  not ginst769 (1398, 768);
  not ginst770 (1401, 762);
  not ginst771 (1404, 806);
  not ginst772 (1407, 800);
  not ginst773 (1410, 794);
  not ginst774 (1413, 780);
  not ginst775 (1416, 774);
  not ginst776 (1419, 768);
  not ginst777 (1422, 762);
  not ginst778 (1425, 786);
  not ginst779 (1428, 636);
  not ginst780 (1431, 636);
  not ginst781 (1434, 865);
  not ginst782 (1437, 859);
  not ginst783 (1440, 853);
  not ginst784 (1443, 845);
  not ginst785 (1446, 839);
  not ginst786 (1449, 833);
  not ginst787 (1452, 827);
  not ginst788 (1455, 821);
  not ginst789 (1458, 814);
  not ginst790 (1461, 865);
  not ginst791 (1464, 859);
  not ginst792 (1467, 853);
  not ginst793 (1470, 839);
  not ginst794 (1473, 833);
  not ginst795 (1476, 827);
  not ginst796 (1479, 821);
  not ginst797 (1482, 845);
  not ginst798 (1485, 814);
  not ginst799 (1489, 1109);
  not ginst800 (1490, 1116);
  and ginst801 (1537, 957, 614);
  and ginst802 (1551, 614, 957);
  and ginst803 (1649, 1029, 636);
  not ginst804 (1703, 957);
  nor ginst805 (1708, 957, 614);
  not ginst806 (1713, 957);
  nor ginst807 (1721, 614, 957);
  not ginst808 (1758, 1029);
  and ginst809 (1781, 163, 1116);
  and ginst810 (1782, 170, 1125);
  not ginst811 (1783, 1125);
  not ginst812 (1789, 1136);
  and ginst813 (1793, 169, 1125);
  and ginst814 (1794, 168, 1125);
  and ginst815 (1795, 167, 1125);
  and ginst816 (1796, 166, 1136);
  and ginst817 (1797, 165, 1136);
  and ginst818 (1798, 164, 1136);
  not ginst819 (1799, 1147);
  not ginst820 (1805, 1160);
  and ginst821 (1811, 177, 1147);
  and ginst822 (1812, 176, 1147);
  and ginst823 (1813, 175, 1147);
  and ginst824 (1814, 174, 1147);
  and ginst825 (1815, 173, 1147);
  and ginst826 (1816, 157, 1160);
  and ginst827 (1817, 156, 1160);
  and ginst828 (1818, 155, 1160);
  and ginst829 (1819, 154, 1160);
  and ginst830 (1820, 153, 1160);
  not ginst831 (1821, 1284);
  not ginst832 (1822, 1287);
  not ginst833 (1828, 1290);
  not ginst834 (1829, 1293);
  not ginst835 (1830, 1296);
  not ginst836 (1832, 1299);
  not ginst837 (1833, 1302);
  not ginst838 (1834, 1305);
  not ginst839 (1835, 1308);
  not ginst840 (1839, 1311);
  not ginst841 (1840, 1314);
  not ginst842 (1841, 1317);
  not ginst843 (1842, 1320);
  not ginst844 (1843, 1323);
  not ginst845 (1845, 1175);
  not ginst846 (1851, 1182);
  and ginst847 (1857, 181, 1175);
  and ginst848 (1858, 171, 1175);
  and ginst849 (1859, 180, 1175);
  and ginst850 (1860, 179, 1175);
  and ginst851 (1861, 178, 1175);
  and ginst852 (1862, 161, 1182);
  and ginst853 (1863, 151, 1182);
  and ginst854 (1864, 160, 1182);
  and ginst855 (1865, 159, 1182);
  and ginst856 (1866, 158, 1182);
  not ginst857 (1867, 1326);
  not ginst858 (1868, 1329);
  not ginst859 (1869, 1332);
  not ginst860 (1870, 1335);
  not ginst861 (1871, 1338);
  not ginst862 (1872, 1341);
  not ginst863 (1873, 1344);
  not ginst864 (1874, 1347);
  not ginst865 (1875, 1350);
  not ginst866 (1876, 1353);
  not ginst867 (1877, 1356);
  not ginst868 (1878, 1359);
  not ginst869 (1879, 1362);
  not ginst870 (1880, 1365);
  not ginst871 (1881, 1368);
  not ginst872 (1882, 1371);
  not ginst873 (1883, 1374);
  not ginst874 (1884, 1377);
  not ginst875 (1885, 1199);
  not ginst876 (1892, 1194);
  not ginst877 (1899, 1199);
  not ginst878 (1906, 1194);
  not ginst879 (1913, 1211);
  not ginst880 (1919, 1194);
  and ginst881 (1926, 44, 1211);
  and ginst882 (1927, 41, 1211);
  and ginst883 (1928, 29, 1211);
  and ginst884 (1929, 26, 1211);
  and ginst885 (1930, 23, 1211);
  not ginst886 (1931, 1380);
  not ginst887 (1932, 1383);
  not ginst888 (1933, 1386);
  not ginst889 (1934, 1389);
  not ginst890 (1935, 1392);
  not ginst891 (1936, 1395);
  not ginst892 (1937, 1398);
  not ginst893 (1938, 1401);
  not ginst894 (1939, 1404);
  not ginst895 (1940, 1407);
  not ginst896 (1941, 1410);
  not ginst897 (1942, 1413);
  not ginst898 (1943, 1416);
  not ginst899 (1944, 1419);
  not ginst900 (1945, 1422);
  not ginst901 (1946, 1425);
  not ginst902 (1947, 1233);
  not ginst903 (1953, 1244);
  and ginst904 (1957, 209, 1233);
  and ginst905 (1958, 216, 1233);
  and ginst906 (1959, 215, 1233);
  and ginst907 (1960, 214, 1233);
  and ginst908 (1961, 213, 1244);
  and ginst909 (1962, 212, 1244);
  and ginst910 (1963, 211, 1244);
  not ginst911 (1965, 1428);
  and ginst912 (1966, 1222, 636);
  not ginst913 (1967, 1431);
  not ginst914 (1968, 1434);
  not ginst915 (1969, 1437);
  not ginst916 (1970, 1440);
  not ginst917 (1971, 1443);
  not ginst918 (1972, 1446);
  not ginst919 (1973, 1449);
  not ginst920 (1974, 1452);
  not ginst921 (1975, 1455);
  not ginst922 (1976, 1458);
  not ginst923 (1977, 1249);
  not ginst924 (1983, 1256);
  and ginst925 (1989, 642, 1249);
  and ginst926 (1990, 644, 1249);
  and ginst927 (1991, 651, 1249);
  and ginst928 (1992, 674, 1249);
  and ginst929 (1993, 660, 1249);
  and ginst930 (1994, 666, 1256);
  and ginst931 (1995, 672, 1256);
  and ginst932 (1996, 673, 1256);
  not ginst933 (1997, 1263);
  not ginst934 (2003, 1194);
  and ginst935 (2010, 47, 1263);
  and ginst936 (2011, 35, 1263);
  and ginst937 (2012, 32, 1263);
  and ginst938 (2013, 50, 1263);
  and ginst939 (2014, 66, 1263);
  not ginst940 (2015, 1461);
  not ginst941 (2016, 1464);
  not ginst942 (2017, 1467);
  not ginst943 (2018, 1470);
  not ginst944 (2019, 1473);
  not ginst945 (2020, 1476);
  not ginst946 (2021, 1479);
  not ginst947 (2022, 1482);
  not ginst948 (2023, 1485);
  not ginst949 (2024, 1206);
  not ginst950 (2031, 1206);
  not ginst951 (2038, 1206);
  not ginst952 (2045, 1206);
  not ginst953 (2052, 1270);
  not ginst954 (2058, 1277);
  and ginst955 (2064, 706, 1270);
  and ginst956 (2065, 708, 1270);
  and ginst957 (2066, 715, 1270);
  and ginst958 (2067, 721, 1270);
  and ginst959 (2068, 727, 1270);
  and ginst960 (2069, 733, 1277);
  and ginst961 (2070, 734, 1277);
  and ginst962 (2071, 742, 1277);
  and ginst963 (2072, 748, 1277);
  and ginst964 (2073, 749, 1277);
  not ginst965 (2074, 1189);
  not ginst966 (2081, 1189);
  not ginst967 (2086, 1222);
  nand ginst968 (2107, 1287, 1821);
  nand ginst969 (2108, 1284, 1822);
  not ginst970 (2110, 1703);
  nand ginst971 (2111, 1703, 1832);
  nand ginst972 (2112, 1308, 1834);
  nand ginst973 (2113, 1305, 1835);
  not ginst974 (2114, 1713);
  nand ginst975 (2115, 1713, 1839);
  not ginst976 (2117, 1721);
  not ginst977 (2171, 1758);
  nand ginst978 (2172, 1758, 1965);
  not ginst979 (2230, 1708);
  not ginst980 (2231, 1537);
  not ginst981 (2235, 1551);
  or ginst982 (2239, 1783, 1782);
  or ginst983 (2240, 1783, 1125);
  or ginst984 (2241, 1783, 1793);
  or ginst985 (2242, 1783, 1794);
  or ginst986 (2243, 1783, 1795);
  or ginst987 (2244, 1789, 1796);
  or ginst988 (2245, 1789, 1797);
  or ginst989 (2246, 1789, 1798);
  or ginst990 (2247, 1799, 1811);
  or ginst991 (2248, 1799, 1812);
  or ginst992 (2249, 1799, 1813);
  or ginst993 (2250, 1799, 1814);
  or ginst994 (2251, 1799, 1815);
  or ginst995 (2252, 1805, 1816);
  or ginst996 (2253, 1805, 1817);
  or ginst997 (2254, 1805, 1818);
  or ginst998 (2255, 1805, 1819);
  or ginst999 (2256, 1805, 1820);
  nand ginst1000 (2257, 2107, 2108);
  not ginst1001 (2267, 2074);
  nand ginst1002 (2268, 1299, 2110);
  nand ginst1003 (2269, 2112, 2113);
  nand ginst1004 (2274, 1311, 2114);
  not ginst1005 (2275, 2081);
  and ginst1006 (2277, 141, 1845);
  and ginst1007 (2278, 147, 1845);
  and ginst1008 (2279, 138, 1845);
  and ginst1009 (2280, 144, 1845);
  and ginst1010 (2281, 135, 1845);
  and ginst1011 (2282, 141, 1851);
  and ginst1012 (2283, 147, 1851);
  and ginst1013 (2284, 138, 1851);
  and ginst1014 (2285, 144, 1851);
  and ginst1015 (2286, 135, 1851);
  not ginst1016 (2287, 1885);
  not ginst1017 (2293, 1892);
  and ginst1018 (2299, 103, 1885);
  and ginst1019 (2300, 130, 1885);
  and ginst1020 (2301, 127, 1885);
  and ginst1021 (2302, 124, 1885);
  and ginst1022 (2303, 100, 1885);
  and ginst1023 (2304, 103, 1892);
  and ginst1024 (2305, 130, 1892);
  and ginst1025 (2306, 127, 1892);
  and ginst1026 (2307, 124, 1892);
  and ginst1027 (2308, 100, 1892);
  not ginst1028 (2309, 1899);
  not ginst1029 (2315, 1906);
  and ginst1030 (2321, 115, 1899);
  and ginst1031 (2322, 118, 1899);
  and ginst1032 (2323, 97, 1899);
  and ginst1033 (2324, 94, 1899);
  and ginst1034 (2325, 121, 1899);
  and ginst1035 (2326, 115, 1906);
  and ginst1036 (2327, 118, 1906);
  and ginst1037 (2328, 97, 1906);
  and ginst1038 (2329, 94, 1906);
  and ginst1039 (2330, 121, 1906);
  not ginst1040 (2331, 1919);
  and ginst1041 (2337, 208, 1913);
  and ginst1042 (2338, 198, 1913);
  and ginst1043 (2339, 207, 1913);
  and ginst1044 (2340, 206, 1913);
  and ginst1045 (2341, 205, 1913);
  and ginst1046 (2342, 44, 1919);
  and ginst1047 (2343, 41, 1919);
  and ginst1048 (2344, 29, 1919);
  and ginst1049 (2345, 26, 1919);
  and ginst1050 (2346, 23, 1919);
  or ginst1051 (2347, 1947, 1233);
  or ginst1052 (2348, 1947, 1957);
  or ginst1053 (2349, 1947, 1958);
  or ginst1054 (2350, 1947, 1959);
  or ginst1055 (2351, 1947, 1960);
  or ginst1056 (2352, 1953, 1961);
  or ginst1057 (2353, 1953, 1962);
  or ginst1058 (2354, 1953, 1963);
  nand ginst1059 (2355, 1428, 2171);
  not ginst1060 (2356, 2086);
  nand ginst1061 (2357, 2086, 1967);
  and ginst1062 (2358, 114, 1977);
  and ginst1063 (2359, 113, 1977);
  and ginst1064 (2360, 111, 1977);
  and ginst1065 (2361, 87, 1977);
  and ginst1066 (2362, 112, 1977);
  and ginst1067 (2363, 88, 1983);
  and ginst1068 (2364, 245, 1983);
  and ginst1069 (2365, 271, 1983);
  and ginst1070 (2366, 759, 1983);
  and ginst1071 (2367, 70, 1983);
  not ginst1072 (2368, 2003);
  and ginst1073 (2374, 193, 1997);
  and ginst1074 (2375, 192, 1997);
  and ginst1075 (2376, 191, 1997);
  and ginst1076 (2377, 190, 1997);
  and ginst1077 (2378, 189, 1997);
  and ginst1078 (2379, 47, 2003);
  and ginst1079 (2380, 35, 2003);
  and ginst1080 (2381, 32, 2003);
  and ginst1081 (2382, 50, 2003);
  and ginst1082 (2383, 66, 2003);
  not ginst1083 (2384, 2024);
  not ginst1084 (2390, 2031);
  and ginst1085 (2396, 58, 2024);
  and ginst1086 (2397, 77, 2024);
  and ginst1087 (2398, 78, 2024);
  and ginst1088 (2399, 59, 2024);
  and ginst1089 (2400, 81, 2024);
  and ginst1090 (2401, 80, 2031);
  and ginst1091 (2402, 79, 2031);
  and ginst1092 (2403, 60, 2031);
  and ginst1093 (2404, 61, 2031);
  and ginst1094 (2405, 62, 2031);
  not ginst1095 (2406, 2038);
  not ginst1096 (2412, 2045);
  and ginst1097 (2418, 69, 2038);
  and ginst1098 (2419, 70, 2038);
  and ginst1099 (2420, 74, 2038);
  and ginst1100 (2421, 76, 2038);
  and ginst1101 (2422, 75, 2038);
  and ginst1102 (2423, 73, 2045);
  and ginst1103 (2424, 53, 2045);
  and ginst1104 (2425, 54, 2045);
  and ginst1105 (2426, 55, 2045);
  and ginst1106 (2427, 56, 2045);
  and ginst1107 (2428, 82, 2052);
  and ginst1108 (2429, 65, 2052);
  and ginst1109 (2430, 83, 2052);
  and ginst1110 (2431, 84, 2052);
  and ginst1111 (2432, 85, 2052);
  and ginst1112 (2433, 64, 2058);
  and ginst1113 (2434, 63, 2058);
  and ginst1114 (2435, 86, 2058);
  and ginst1115 (2436, 109, 2058);
  and ginst1116 (2437, 110, 2058);
  and ginst1117 (2441, 2239, 1119);
  and ginst1118 (2442, 2240, 1119);
  and ginst1119 (2446, 2241, 1119);
  and ginst1120 (2450, 2242, 1119);
  and ginst1121 (2454, 2243, 1119);
  and ginst1122 (2458, 2244, 1132);
  and ginst1123 (2462, 2247, 1141);
  and ginst1124 (2466, 2248, 1141);
  and ginst1125 (2470, 2249, 1141);
  and ginst1126 (2474, 2250, 1141);
  and ginst1127 (2478, 2251, 1141);
  and ginst1128 (2482, 2252, 1154);
  and ginst1129 (2488, 2253, 1154);
  and ginst1130 (2496, 2254, 1154);
  and ginst1131 (2502, 2255, 1154);
  and ginst1132 (2508, 2256, 1154);
  nand ginst1133 (2523, 2268, 2111);
  nand ginst1134 (2533, 2274, 2115);
  not ginst1135 (2537, 2235);
  or ginst1136 (2538, 2278, 1858);
  or ginst1137 (2542, 2279, 1859);
  or ginst1138 (2546, 2280, 1860);
  or ginst1139 (2550, 2281, 1861);
  or ginst1140 (2554, 2283, 1863);
  or ginst1141 (2561, 2284, 1864);
  or ginst1142 (2567, 2285, 1865);
  or ginst1143 (2573, 2286, 1866);
  or ginst1144 (2604, 2338, 1927);
  or ginst1145 (2607, 2339, 1928);
  or ginst1146 (2611, 2340, 1929);
  or ginst1147 (2615, 2341, 1930);
  and ginst1148 (2619, 2348, 1227);
  and ginst1149 (2626, 2349, 1227);
  and ginst1150 (2632, 2350, 1227);
  and ginst1151 (2638, 2351, 1227);
  and ginst1152 (2644, 2352, 1240);
  nand ginst1153 (2650, 2355, 2172);
  nand ginst1154 (2653, 1431, 2356);
  or ginst1155 (2654, 2359, 1990);
  or ginst1156 (2658, 2360, 1991);
  or ginst1157 (2662, 2361, 1992);
  or ginst1158 (2666, 2362, 1993);
  or ginst1159 (2670, 2363, 1994);
  or ginst1160 (2674, 2366, 1256);
  or ginst1161 (2680, 2367, 1256);
  or ginst1162 (2688, 2374, 2010);
  or ginst1163 (2692, 2375, 2011);
  or ginst1164 (2696, 2376, 2012);
  or ginst1165 (2700, 2377, 2013);
  or ginst1166 (2704, 2378, 2014);
  and ginst1167 (2728, 2347, 1227);
  or ginst1168 (2729, 2429, 2065);
  or ginst1169 (2733, 2430, 2066);
  or ginst1170 (2737, 2431, 2067);
  or ginst1171 (2741, 2432, 2068);
  or ginst1172 (2745, 2433, 2069);
  or ginst1173 (2749, 2434, 2070);
  or ginst1174 (2753, 2435, 2071);
  or ginst1175 (2757, 2436, 2072);
  or ginst1176 (2761, 2437, 2073);
  not ginst1177 (2765, 2231);
  and ginst1178 (2766, 2354, 1240);
  and ginst1179 (2769, 2353, 1240);
  and ginst1180 (2772, 2246, 1132);
  and ginst1181 (2775, 2245, 1132);
  or ginst1182 (2778, 2282, 1862);
  or ginst1183 (2781, 2358, 1989);
  or ginst1184 (2784, 2365, 1996);
  or ginst1185 (2787, 2364, 1995);
  or ginst1186 (2790, 2337, 1926);
  or ginst1187 (2793, 2277, 1857);
  or ginst1188 (2796, 2428, 2064);
  and ginst1189 (2866, 2257, 1537);
  and ginst1190 (2867, 2257, 1537);
  and ginst1191 (2868, 2257, 1537);
  and ginst1192 (2869, 2257, 1537);
  and ginst1193 (2878, 2269, 1551);
  and ginst1194 (2913, 204, 2287);
  and ginst1195 (2914, 203, 2287);
  and ginst1196 (2915, 202, 2287);
  and ginst1197 (2916, 201, 2287);
  and ginst1198 (2917, 200, 2287);
  and ginst1199 (2918, 235, 2293);
  and ginst1200 (2919, 234, 2293);
  and ginst1201 (2920, 233, 2293);
  and ginst1202 (2921, 232, 2293);
  and ginst1203 (2922, 231, 2293);
  and ginst1204 (2923, 197, 2309);
  and ginst1205 (2924, 187, 2309);
  and ginst1206 (2925, 196, 2309);
  and ginst1207 (2926, 195, 2309);
  and ginst1208 (2927, 194, 2309);
  and ginst1209 (2928, 227, 2315);
  and ginst1210 (2929, 217, 2315);
  and ginst1211 (2930, 226, 2315);
  and ginst1212 (2931, 225, 2315);
  and ginst1213 (2932, 224, 2315);
  and ginst1214 (2933, 239, 2331);
  and ginst1215 (2934, 229, 2331);
  and ginst1216 (2935, 238, 2331);
  and ginst1217 (2936, 237, 2331);
  and ginst1218 (2937, 236, 2331);
  nand ginst1219 (2988, 2653, 2357);
  and ginst1220 (3005, 223, 2368);
  and ginst1221 (3006, 222, 2368);
  and ginst1222 (3007, 221, 2368);
  and ginst1223 (3008, 220, 2368);
  and ginst1224 (3009, 219, 2368);
  and ginst1225 (3020, 812, 2384);
  and ginst1226 (3021, 814, 2384);
  and ginst1227 (3022, 821, 2384);
  and ginst1228 (3023, 827, 2384);
  and ginst1229 (3024, 833, 2384);
  and ginst1230 (3025, 839, 2390);
  and ginst1231 (3026, 845, 2390);
  and ginst1232 (3027, 853, 2390);
  and ginst1233 (3028, 859, 2390);
  and ginst1234 (3029, 865, 2390);
  and ginst1235 (3032, 758, 2406);
  and ginst1236 (3033, 759, 2406);
  and ginst1237 (3034, 762, 2406);
  and ginst1238 (3035, 768, 2406);
  and ginst1239 (3036, 774, 2406);
  and ginst1240 (3037, 780, 2412);
  and ginst1241 (3038, 786, 2412);
  and ginst1242 (3039, 794, 2412);
  and ginst1243 (3040, 800, 2412);
  and ginst1244 (3041, 806, 2412);
  not ginst1245 (3061, 2257);
  not ginst1246 (3064, 2257);
  not ginst1247 (3067, 2269);
  not ginst1248 (3070, 2269);
  not ginst1249 (3073, 2728);
  not ginst1250 (3080, 2441);
  and ginst1251 (3096, 666, 2644);
  and ginst1252 (3097, 660, 2638);
  and ginst1253 (3101, 1189, 2632);
  and ginst1254 (3107, 651, 2626);
  and ginst1255 (3114, 644, 2619);
  and ginst1256 (3122, 2523, 2257);
  or ginst1257 (3126, 1167, 2866);
  and ginst1258 (3130, 2523, 2257);
  or ginst1259 (3131, 1167, 2869);
  and ginst1260 (3134, 2523, 2257);
  not ginst1261 (3135, 2533);
  and ginst1262 (3136, 666, 2644);
  and ginst1263 (3137, 660, 2638);
  and ginst1264 (3140, 1189, 2632);
  and ginst1265 (3144, 651, 2626);
  and ginst1266 (3149, 644, 2619);
  and ginst1267 (3155, 2533, 2269);
  or ginst1268 (3159, 1174, 2878);
  not ginst1269 (3167, 2778);
  and ginst1270 (3168, 609, 2508);
  and ginst1271 (3169, 604, 2502);
  and ginst1272 (3173, 742, 2496);
  and ginst1273 (3178, 734, 2488);
  and ginst1274 (3184, 599, 2482);
  and ginst1275 (3185, 727, 2573);
  and ginst1276 (3189, 721, 2567);
  and ginst1277 (3195, 715, 2561);
  and ginst1278 (3202, 708, 2554);
  and ginst1279 (3210, 609, 2508);
  and ginst1280 (3211, 604, 2502);
  and ginst1281 (3215, 742, 2496);
  and ginst1282 (3221, 2488, 734);
  and ginst1283 (3228, 599, 2482);
  and ginst1284 (3229, 727, 2573);
  and ginst1285 (3232, 721, 2567);
  and ginst1286 (3236, 715, 2561);
  and ginst1287 (3241, 708, 2554);
  or ginst1288 (3247, 2913, 2299);
  or ginst1289 (3251, 2914, 2300);
  or ginst1290 (3255, 2915, 2301);
  or ginst1291 (3259, 2916, 2302);
  or ginst1292 (3263, 2917, 2303);
  or ginst1293 (3267, 2918, 2304);
  or ginst1294 (3273, 2919, 2305);
  or ginst1295 (3281, 2920, 2306);
  or ginst1296 (3287, 2921, 2307);
  or ginst1297 (3293, 2922, 2308);
  or ginst1298 (3299, 2924, 2322);
  or ginst1299 (3303, 2925, 2323);
  or ginst1300 (3307, 2926, 2324);
  or ginst1301 (3311, 2927, 2325);
  or ginst1302 (3315, 2929, 2327);
  or ginst1303 (3322, 2930, 2328);
  or ginst1304 (3328, 2931, 2329);
  or ginst1305 (3334, 2932, 2330);
  or ginst1306 (3340, 2934, 2343);
  or ginst1307 (3343, 2935, 2344);
  or ginst1308 (3349, 2936, 2345);
  or ginst1309 (3355, 2937, 2346);
  and ginst1310 (3361, 2761, 2478);
  and ginst1311 (3362, 2757, 2474);
  and ginst1312 (3363, 2753, 2470);
  and ginst1313 (3364, 2749, 2466);
  and ginst1314 (3365, 2745, 2462);
  and ginst1315 (3366, 2741, 2550);
  and ginst1316 (3367, 2737, 2546);
  and ginst1317 (3368, 2733, 2542);
  and ginst1318 (3369, 2729, 2538);
  and ginst1319 (3370, 2670, 2458);
  and ginst1320 (3371, 2666, 2454);
  and ginst1321 (3372, 2662, 2450);
  and ginst1322 (3373, 2658, 2446);
  and ginst1323 (3374, 2654, 2442);
  and ginst1324 (3375, 2988, 2650);
  and ginst1325 (3379, 2650, 1966);
  not ginst1326 (3380, 2781);
  and ginst1327 (3381, 695, 2604);
  or ginst1328 (3384, 3005, 2379);
  or ginst1329 (3390, 3006, 2380);
  or ginst1330 (3398, 3007, 2381);
  or ginst1331 (3404, 3008, 2382);
  or ginst1332 (3410, 3009, 2383);
  or ginst1333 (3416, 3021, 2397);
  or ginst1334 (3420, 3022, 2398);
  or ginst1335 (3424, 3023, 2399);
  or ginst1336 (3428, 3024, 2400);
  or ginst1337 (3432, 3025, 2401);
  or ginst1338 (3436, 3026, 2402);
  or ginst1339 (3440, 3027, 2403);
  or ginst1340 (3444, 3028, 2404);
  or ginst1341 (3448, 3029, 2405);
  not ginst1342 (3452, 2790);
  not ginst1343 (3453, 2793);
  or ginst1344 (3454, 3034, 2420);
  or ginst1345 (3458, 3035, 2421);
  or ginst1346 (3462, 3036, 2422);
  or ginst1347 (3466, 3037, 2423);
  or ginst1348 (3470, 3038, 2424);
  or ginst1349 (3474, 3039, 2425);
  or ginst1350 (3478, 3040, 2426);
  or ginst1351 (3482, 3041, 2427);
  not ginst1352 (3486, 2796);
  not ginst1353 (3487, 2644);
  not ginst1354 (3490, 2638);
  not ginst1355 (3493, 2632);
  not ginst1356 (3496, 2626);
  not ginst1357 (3499, 2619);
  not ginst1358 (3502, 2523);
  nor ginst1359 (3507, 1167, 2868);
  not ginst1360 (3510, 2523);
  nor ginst1361 (3515, 644, 2619);
  not ginst1362 (3518, 2644);
  not ginst1363 (3521, 2638);
  not ginst1364 (3524, 2632);
  not ginst1365 (3527, 2626);
  not ginst1366 (3530, 2619);
  not ginst1367 (3535, 2619);
  not ginst1368 (3539, 2632);
  not ginst1369 (3542, 2626);
  not ginst1370 (3545, 2644);
  not ginst1371 (3548, 2638);
  not ginst1372 (3551, 2766);
  not ginst1373 (3552, 2769);
  not ginst1374 (3553, 2442);
  not ginst1375 (3557, 2450);
  not ginst1376 (3560, 2446);
  not ginst1377 (3563, 2458);
  not ginst1378 (3566, 2454);
  not ginst1379 (3569, 2772);
  not ginst1380 (3570, 2775);
  not ginst1381 (3571, 2554);
  not ginst1382 (3574, 2567);
  not ginst1383 (3577, 2561);
  not ginst1384 (3580, 2482);
  not ginst1385 (3583, 2573);
  not ginst1386 (3586, 2496);
  not ginst1387 (3589, 2488);
  not ginst1388 (3592, 2508);
  not ginst1389 (3595, 2502);
  not ginst1390 (3598, 2508);
  not ginst1391 (3601, 2502);
  not ginst1392 (3604, 2496);
  not ginst1393 (3607, 2482);
  not ginst1394 (3610, 2573);
  not ginst1395 (3613, 2567);
  not ginst1396 (3616, 2561);
  not ginst1397 (3619, 2488);
  not ginst1398 (3622, 2554);
  nor ginst1399 (3625, 734, 2488);
  nor ginst1400 (3628, 708, 2554);
  not ginst1401 (3631, 2508);
  not ginst1402 (3634, 2502);
  not ginst1403 (3637, 2496);
  not ginst1404 (3640, 2488);
  not ginst1405 (3643, 2482);
  not ginst1406 (3646, 2573);
  not ginst1407 (3649, 2567);
  not ginst1408 (3652, 2561);
  not ginst1409 (3655, 2554);
  nor ginst1410 (3658, 2488, 734);
  not ginst1411 (3661, 2674);
  not ginst1412 (3664, 2674);
  not ginst1413 (3667, 2761);
  not ginst1414 (3670, 2478);
  not ginst1415 (3673, 2757);
  not ginst1416 (3676, 2474);
  not ginst1417 (3679, 2753);
  not ginst1418 (3682, 2470);
  not ginst1419 (3685, 2745);
  not ginst1420 (3688, 2462);
  not ginst1421 (3691, 2741);
  not ginst1422 (3694, 2550);
  not ginst1423 (3697, 2737);
  not ginst1424 (3700, 2546);
  not ginst1425 (3703, 2733);
  not ginst1426 (3706, 2542);
  not ginst1427 (3709, 2749);
  not ginst1428 (3712, 2466);
  not ginst1429 (3715, 2729);
  not ginst1430 (3718, 2538);
  not ginst1431 (3721, 2704);
  not ginst1432 (3724, 2700);
  not ginst1433 (3727, 2696);
  not ginst1434 (3730, 2688);
  not ginst1435 (3733, 2692);
  not ginst1436 (3736, 2670);
  not ginst1437 (3739, 2458);
  not ginst1438 (3742, 2666);
  not ginst1439 (3745, 2454);
  not ginst1440 (3748, 2662);
  not ginst1441 (3751, 2450);
  not ginst1442 (3754, 2658);
  not ginst1443 (3757, 2446);
  not ginst1444 (3760, 2654);
  not ginst1445 (3763, 2442);
  not ginst1446 (3766, 2654);
  not ginst1447 (3769, 2662);
  not ginst1448 (3772, 2658);
  not ginst1449 (3775, 2670);
  not ginst1450 (3778, 2666);
  not ginst1451 (3781, 2784);
  not ginst1452 (3782, 2787);
  or ginst1453 (3783, 2928, 2326);
  or ginst1454 (3786, 2933, 2342);
  or ginst1455 (3789, 2923, 2321);
  not ginst1456 (3792, 2688);
  not ginst1457 (3795, 2696);
  not ginst1458 (3798, 2692);
  not ginst1459 (3801, 2704);
  not ginst1460 (3804, 2700);
  not ginst1461 (3807, 2604);
  not ginst1462 (3810, 2611);
  not ginst1463 (3813, 2607);
  not ginst1464 (3816, 2615);
  not ginst1465 (3819, 2538);
  not ginst1466 (3822, 2546);
  not ginst1467 (3825, 2542);
  not ginst1468 (3828, 2462);
  not ginst1469 (3831, 2550);
  not ginst1470 (3834, 2470);
  not ginst1471 (3837, 2466);
  not ginst1472 (3840, 2478);
  not ginst1473 (3843, 2474);
  not ginst1474 (3846, 2615);
  not ginst1475 (3849, 2611);
  not ginst1476 (3852, 2607);
  not ginst1477 (3855, 2680);
  not ginst1478 (3858, 2729);
  not ginst1479 (3861, 2737);
  not ginst1480 (3864, 2733);
  not ginst1481 (3867, 2745);
  not ginst1482 (387, 1);
  not ginst1483 (3870, 2741);
  not ginst1484 (3873, 2753);
  not ginst1485 (3876, 2749);
  not ginst1486 (3879, 2761);
  not ginst1487 (388, 1);
  not ginst1488 (3882, 2757);
  or ginst1489 (3885, 3033, 2419);
  or ginst1490 (3888, 3032, 2418);
  or ginst1491 (3891, 3020, 2396);
  nand ginst1492 (3953, 3067, 2117);
  not ginst1493 (3954, 3067);
  nand ginst1494 (3955, 3070, 2537);
  not ginst1495 (3956, 3070);
  not ginst1496 (3958, 3073);
  not ginst1497 (3964, 3080);
  or ginst1498 (4193, 1649, 3379);
  or ginst1499 (4303, 1167, 2867, 3130);
  not ginst1500 (4308, 3061);
  not ginst1501 (4313, 3064);
  nand ginst1502 (4326, 2769, 3551);
  nand ginst1503 (4327, 2766, 3552);
  nand ginst1504 (4333, 2775, 3569);
  nand ginst1505 (4334, 2772, 3570);
  nand ginst1506 (4411, 2787, 3781);
  nand ginst1507 (4412, 2784, 3782);
  nand ginst1508 (4463, 3487, 1828);
  not ginst1509 (4464, 3487);
  nand ginst1510 (4465, 3490, 1829);
  not ginst1511 (4466, 3490);
  nand ginst1512 (4467, 3493, 2267);
  not ginst1513 (4468, 3493);
  nand ginst1514 (4469, 3496, 1830);
  not ginst1515 (4470, 3496);
  nand ginst1516 (4471, 3499, 1833);
  not ginst1517 (4472, 3499);
  not ginst1518 (4473, 3122);
  not ginst1519 (4474, 3126);
  nand ginst1520 (4475, 3518, 1840);
  not ginst1521 (4476, 3518);
  nand ginst1522 (4477, 3521, 1841);
  not ginst1523 (4478, 3521);
  nand ginst1524 (4479, 3524, 2275);
  not ginst1525 (4480, 3524);
  nand ginst1526 (4481, 3527, 1842);
  not ginst1527 (4482, 3527);
  nand ginst1528 (4483, 3530, 1843);
  not ginst1529 (4484, 3530);
  not ginst1530 (4485, 3155);
  not ginst1531 (4486, 3159);
  nand ginst1532 (4487, 1721, 3954);
  nand ginst1533 (4488, 2235, 3956);
  not ginst1534 (4489, 3535);
  nand ginst1535 (4490, 3535, 3958);
  not ginst1536 (4491, 3539);
  not ginst1537 (4492, 3542);
  not ginst1538 (4493, 3545);
  not ginst1539 (4494, 3548);
  not ginst1540 (4495, 3553);
  nand ginst1541 (4496, 3553, 3964);
  not ginst1542 (4497, 3557);
  not ginst1543 (4498, 3560);
  not ginst1544 (4499, 3563);
  not ginst1545 (4500, 3566);
  not ginst1546 (4501, 3571);
  nand ginst1547 (4502, 3571, 3167);
  not ginst1548 (4503, 3574);
  not ginst1549 (4504, 3577);
  not ginst1550 (4505, 3580);
  not ginst1551 (4506, 3583);
  nand ginst1552 (4507, 3598, 1867);
  not ginst1553 (4508, 3598);
  nand ginst1554 (4509, 3601, 1868);
  not ginst1555 (4510, 3601);
  nand ginst1556 (4511, 3604, 1869);
  not ginst1557 (4512, 3604);
  nand ginst1558 (4513, 3607, 1870);
  not ginst1559 (4514, 3607);
  nand ginst1560 (4515, 3610, 1871);
  not ginst1561 (4516, 3610);
  nand ginst1562 (4517, 3613, 1872);
  not ginst1563 (4518, 3613);
  nand ginst1564 (4519, 3616, 1873);
  not ginst1565 (4520, 3616);
  nand ginst1566 (4521, 3619, 1874);
  not ginst1567 (4522, 3619);
  nand ginst1568 (4523, 3622, 1875);
  not ginst1569 (4524, 3622);
  nand ginst1570 (4525, 3631, 1876);
  not ginst1571 (4526, 3631);
  nand ginst1572 (4527, 3634, 1877);
  not ginst1573 (4528, 3634);
  nand ginst1574 (4529, 3637, 1878);
  not ginst1575 (4530, 3637);
  nand ginst1576 (4531, 3640, 1879);
  not ginst1577 (4532, 3640);
  nand ginst1578 (4533, 3643, 1880);
  not ginst1579 (4534, 3643);
  nand ginst1580 (4535, 3646, 1881);
  not ginst1581 (4536, 3646);
  nand ginst1582 (4537, 3649, 1882);
  not ginst1583 (4538, 3649);
  nand ginst1584 (4539, 3652, 1883);
  not ginst1585 (4540, 3652);
  nand ginst1586 (4541, 3655, 1884);
  not ginst1587 (4542, 3655);
  not ginst1588 (4543, 3658);
  and ginst1589 (4544, 806, 3293);
  and ginst1590 (4545, 800, 3287);
  and ginst1591 (4549, 794, 3281);
  and ginst1592 (4555, 3273, 786);
  and ginst1593 (4562, 780, 3267);
  and ginst1594 (4563, 774, 3355);
  and ginst1595 (4566, 768, 3349);
  and ginst1596 (4570, 762, 3343);
  not ginst1597 (4575, 3661);
  and ginst1598 (4576, 806, 3293);
  and ginst1599 (4577, 800, 3287);
  and ginst1600 (4581, 794, 3281);
  and ginst1601 (4586, 786, 3273);
  and ginst1602 (4592, 780, 3267);
  and ginst1603 (4593, 774, 3355);
  and ginst1604 (4597, 768, 3349);
  and ginst1605 (4603, 762, 3343);
  not ginst1606 (4610, 3664);
  not ginst1607 (4611, 3667);
  not ginst1608 (4612, 3670);
  not ginst1609 (4613, 3673);
  not ginst1610 (4614, 3676);
  not ginst1611 (4615, 3679);
  not ginst1612 (4616, 3682);
  not ginst1613 (4617, 3685);
  not ginst1614 (4618, 3688);
  not ginst1615 (4619, 3691);
  not ginst1616 (4620, 3694);
  not ginst1617 (4621, 3697);
  not ginst1618 (4622, 3700);
  not ginst1619 (4623, 3703);
  not ginst1620 (4624, 3706);
  not ginst1621 (4625, 3709);
  not ginst1622 (4626, 3712);
  not ginst1623 (4627, 3715);
  not ginst1624 (4628, 3718);
  not ginst1625 (4629, 3721);
  and ginst1626 (4630, 3448, 2704);
  not ginst1627 (4631, 3724);
  and ginst1628 (4632, 3444, 2700);
  not ginst1629 (4633, 3727);
  and ginst1630 (4634, 3440, 2696);
  and ginst1631 (4635, 3436, 2692);
  not ginst1632 (4636, 3730);
  and ginst1633 (4637, 3432, 2688);
  and ginst1634 (4638, 3428, 3311);
  and ginst1635 (4639, 3424, 3307);
  and ginst1636 (4640, 3420, 3303);
  and ginst1637 (4641, 3416, 3299);
  not ginst1638 (4642, 3733);
  not ginst1639 (4643, 3736);
  not ginst1640 (4644, 3739);
  not ginst1641 (4645, 3742);
  not ginst1642 (4646, 3745);
  not ginst1643 (4647, 3748);
  not ginst1644 (4648, 3751);
  not ginst1645 (4649, 3754);
  not ginst1646 (4650, 3757);
  not ginst1647 (4651, 3760);
  not ginst1648 (4652, 3763);
  not ginst1649 (4653, 3375);
  and ginst1650 (4656, 865, 3410);
  and ginst1651 (4657, 859, 3404);
  and ginst1652 (4661, 853, 3398);
  and ginst1653 (4667, 3390, 845);
  not ginst1654 (467, 57);
  and ginst1655 (4674, 839, 3384);
  and ginst1656 (4675, 833, 3334);
  and ginst1657 (4678, 827, 3328);
  and ginst1658 (4682, 821, 3322);
  and ginst1659 (4687, 814, 3315);
  and ginst1660 (469, 134, 133);
  not ginst1661 (4693, 3766);
  nand ginst1662 (4694, 3766, 3380);
  not ginst1663 (4695, 3769);
  not ginst1664 (4696, 3772);
  not ginst1665 (4697, 3775);
  not ginst1666 (4698, 3778);
  not ginst1667 (4699, 3783);
  not ginst1668 (4700, 3786);
  and ginst1669 (4701, 865, 3410);
  and ginst1670 (4702, 859, 3404);
  and ginst1671 (4706, 853, 3398);
  and ginst1672 (4711, 845, 3390);
  and ginst1673 (4717, 839, 3384);
  and ginst1674 (4718, 833, 3334);
  and ginst1675 (4722, 827, 3328);
  and ginst1676 (4728, 821, 3322);
  and ginst1677 (4735, 814, 3315);
  not ginst1678 (4743, 3789);
  not ginst1679 (4744, 3792);
  not ginst1680 (4745, 3807);
  nand ginst1681 (4746, 3807, 3452);
  not ginst1682 (4747, 3810);
  not ginst1683 (4748, 3813);
  not ginst1684 (4749, 3816);
  not ginst1685 (4750, 3819);
  nand ginst1686 (4751, 3819, 3453);
  not ginst1687 (4752, 3822);
  not ginst1688 (4753, 3825);
  not ginst1689 (4754, 3828);
  not ginst1690 (4755, 3831);
  and ginst1691 (4756, 3482, 3263);
  and ginst1692 (4757, 3478, 3259);
  and ginst1693 (4758, 3474, 3255);
  and ginst1694 (4759, 3470, 3251);
  and ginst1695 (4760, 3466, 3247);
  not ginst1696 (4761, 3846);
  and ginst1697 (4762, 3462, 2615);
  not ginst1698 (4763, 3849);
  and ginst1699 (4764, 3458, 2611);
  not ginst1700 (4765, 3852);
  and ginst1701 (4766, 3454, 2607);
  and ginst1702 (4767, 2680, 3381);
  not ginst1703 (4768, 3855);
  and ginst1704 (4769, 3340, 695);
  not ginst1705 (4775, 3858);
  nand ginst1706 (4776, 3858, 3486);
  not ginst1707 (4777, 3861);
  not ginst1708 (4778, 3864);
  not ginst1709 (4779, 3867);
  not ginst1710 (478, 248);
  not ginst1711 (4780, 3870);
  not ginst1712 (4781, 3885);
  not ginst1713 (4782, 3888);
  not ginst1714 (4783, 3891);
  or ginst1715 (4784, 3131, 3134);
  not ginst1716 (4789, 3502);
  not ginst1717 (4790, 3131);
  not ginst1718 (4793, 3507);
  not ginst1719 (4794, 3510);
  not ginst1720 (4795, 3515);
  not ginst1721 (4796, 3114);
  not ginst1722 (4799, 3586);
  not ginst1723 (4800, 3589);
  not ginst1724 (4801, 3592);
  not ginst1725 (4802, 3595);
  nand ginst1726 (4803, 4326, 4327);
  nand ginst1727 (4806, 4333, 4334);
  not ginst1728 (4809, 3625);
  not ginst1729 (4810, 3178);
  not ginst1730 (4813, 3628);
  not ginst1731 (4814, 3202);
  not ginst1732 (4817, 3221);
  not ginst1733 (482, 254);
  not ginst1734 (4820, 3293);
  not ginst1735 (4823, 3287);
  not ginst1736 (4826, 3281);
  not ginst1737 (4829, 3273);
  not ginst1738 (4832, 3267);
  not ginst1739 (4835, 3355);
  not ginst1740 (4838, 3349);
  not ginst1741 (484, 257);
  not ginst1742 (4841, 3343);
  nor ginst1743 (4844, 3273, 786);
  not ginst1744 (4847, 3293);
  not ginst1745 (4850, 3287);
  not ginst1746 (4853, 3281);
  not ginst1747 (4856, 3267);
  not ginst1748 (4859, 3355);
  not ginst1749 (486, 260);
  not ginst1750 (4862, 3349);
  not ginst1751 (4865, 3343);
  not ginst1752 (4868, 3273);
  nor ginst1753 (4871, 786, 3273);
  not ginst1754 (4874, 3448);
  not ginst1755 (4877, 3444);
  not ginst1756 (4880, 3440);
  not ginst1757 (4883, 3432);
  not ginst1758 (4886, 3428);
  not ginst1759 (4889, 3311);
  not ginst1760 (489, 263);
  not ginst1761 (4892, 3424);
  not ginst1762 (4895, 3307);
  not ginst1763 (4898, 3420);
  not ginst1764 (4901, 3303);
  not ginst1765 (4904, 3436);
  not ginst1766 (4907, 3416);
  not ginst1767 (4910, 3299);
  not ginst1768 (4913, 3410);
  not ginst1769 (4916, 3404);
  not ginst1770 (4919, 3398);
  not ginst1771 (492, 267);
  not ginst1772 (4922, 3390);
  not ginst1773 (4925, 3384);
  not ginst1774 (4928, 3334);
  not ginst1775 (4931, 3328);
  not ginst1776 (4934, 3322);
  not ginst1777 (4937, 3315);
  and ginst1778 (494, 162, 172, 188, 199);
  nor ginst1779 (4940, 3390, 845);
  not ginst1780 (4943, 3315);
  not ginst1781 (4946, 3328);
  not ginst1782 (4949, 3322);
  not ginst1783 (4952, 3384);
  not ginst1784 (4955, 3334);
  not ginst1785 (4958, 3398);
  not ginst1786 (4961, 3390);
  not ginst1787 (4964, 3410);
  not ginst1788 (4967, 3404);
  not ginst1789 (4970, 3340);
  not ginst1790 (4973, 3349);
  not ginst1791 (4976, 3343);
  not ginst1792 (4979, 3267);
  not ginst1793 (4982, 3355);
  not ginst1794 (4985, 3281);
  not ginst1795 (4988, 3273);
  not ginst1796 (4991, 3293);
  not ginst1797 (4994, 3287);
  nand ginst1798 (4997, 4411, 4412);
  not ginst1799 (5000, 3410);
  not ginst1800 (5003, 3404);
  not ginst1801 (5006, 3398);
  not ginst1802 (5009, 3384);
  not ginst1803 (501, 274);
  not ginst1804 (5012, 3334);
  not ginst1805 (5015, 3328);
  not ginst1806 (5018, 3322);
  not ginst1807 (5021, 3390);
  not ginst1808 (5024, 3315);
  nor ginst1809 (5027, 845, 3390);
  nor ginst1810 (5030, 814, 3315);
  not ginst1811 (5033, 3299);
  not ginst1812 (5036, 3307);
  not ginst1813 (5039, 3303);
  not ginst1814 (5042, 3311);
  not ginst1815 (5045, 3795);
  not ginst1816 (5046, 3798);
  not ginst1817 (5047, 3801);
  not ginst1818 (5048, 3804);
  not ginst1819 (5049, 3247);
  not ginst1820 (505, 280);
  not ginst1821 (5052, 3255);
  not ginst1822 (5055, 3251);
  not ginst1823 (5058, 3263);
  not ginst1824 (5061, 3259);
  not ginst1825 (5064, 3834);
  not ginst1826 (5065, 3837);
  not ginst1827 (5066, 3840);
  not ginst1828 (5067, 3843);
  not ginst1829 (5068, 3482);
  not ginst1830 (507, 283);
  not ginst1831 (5071, 3263);
  not ginst1832 (5074, 3478);
  not ginst1833 (5077, 3259);
  not ginst1834 (5080, 3474);
  not ginst1835 (5083, 3255);
  not ginst1836 (5086, 3466);
  not ginst1837 (5089, 3247);
  not ginst1838 (509, 286);
  not ginst1839 (5092, 3462);
  not ginst1840 (5095, 3458);
  not ginst1841 (5098, 3454);
  not ginst1842 (5101, 3470);
  not ginst1843 (5104, 3251);
  not ginst1844 (5107, 3381);
  not ginst1845 (511, 289);
  not ginst1846 (5110, 3873);
  not ginst1847 (5111, 3876);
  not ginst1848 (5112, 3879);
  not ginst1849 (5113, 3882);
  not ginst1850 (5114, 3458);
  not ginst1851 (5117, 3454);
  not ginst1852 (5120, 3466);
  not ginst1853 (5123, 3462);
  not ginst1854 (5126, 3474);
  not ginst1855 (5129, 3470);
  not ginst1856 (513, 293);
  not ginst1857 (5132, 3482);
  not ginst1858 (5135, 3478);
  not ginst1859 (5138, 3416);
  not ginst1860 (5141, 3424);
  not ginst1861 (5144, 3420);
  not ginst1862 (5147, 3432);
  not ginst1863 (515, 296);
  not ginst1864 (5150, 3428);
  not ginst1865 (5153, 3440);
  not ginst1866 (5156, 3436);
  not ginst1867 (5159, 3448);
  not ginst1868 (5162, 3444);
  nand ginst1869 (5165, 4486, 4485);
  nand ginst1870 (5166, 4474, 4473);
  nand ginst1871 (5167, 1290, 4464);
  nand ginst1872 (5168, 1293, 4466);
  nand ginst1873 (5169, 2074, 4468);
  not ginst1874 (517, 299);
  nand ginst1875 (5170, 1296, 4470);
  nand ginst1876 (5171, 1302, 4472);
  nand ginst1877 (5172, 1314, 4476);
  nand ginst1878 (5173, 1317, 4478);
  nand ginst1879 (5174, 2081, 4480);
  nand ginst1880 (5175, 1320, 4482);
  nand ginst1881 (5176, 1323, 4484);
  nand ginst1882 (5177, 3953, 4487);
  nand ginst1883 (5178, 3955, 4488);
  nand ginst1884 (5179, 3073, 4489);
  nand ginst1885 (5180, 3542, 4491);
  nand ginst1886 (5181, 3539, 4492);
  nand ginst1887 (5182, 3548, 4493);
  nand ginst1888 (5183, 3545, 4494);
  nand ginst1889 (5184, 3080, 4495);
  nand ginst1890 (5185, 3560, 4497);
  nand ginst1891 (5186, 3557, 4498);
  nand ginst1892 (5187, 3566, 4499);
  nand ginst1893 (5188, 3563, 4500);
  nand ginst1894 (5189, 2778, 4501);
  not ginst1895 (519, 303);
  nand ginst1896 (5190, 3577, 4503);
  nand ginst1897 (5191, 3574, 4504);
  nand ginst1898 (5192, 3583, 4505);
  nand ginst1899 (5193, 3580, 4506);
  nand ginst1900 (5196, 1326, 4508);
  nand ginst1901 (5197, 1329, 4510);
  nand ginst1902 (5198, 1332, 4512);
  nand ginst1903 (5199, 1335, 4514);
  nand ginst1904 (5200, 1338, 4516);
  nand ginst1905 (5201, 1341, 4518);
  nand ginst1906 (5202, 1344, 4520);
  nand ginst1907 (5203, 1347, 4522);
  nand ginst1908 (5204, 1350, 4524);
  nand ginst1909 (5205, 1353, 4526);
  nand ginst1910 (5206, 1356, 4528);
  nand ginst1911 (5207, 1359, 4530);
  nand ginst1912 (5208, 1362, 4532);
  nand ginst1913 (5209, 1365, 4534);
  nand ginst1914 (5210, 1368, 4536);
  nand ginst1915 (5211, 1371, 4538);
  nand ginst1916 (5212, 1374, 4540);
  nand ginst1917 (5213, 1377, 4542);
  and ginst1918 (528, 150, 184, 228, 240);
  nand ginst1919 (5283, 3670, 4611);
  nand ginst1920 (5284, 3667, 4612);
  nand ginst1921 (5285, 3676, 4613);
  nand ginst1922 (5286, 3673, 4614);
  nand ginst1923 (5287, 3682, 4615);
  nand ginst1924 (5288, 3679, 4616);
  nand ginst1925 (5289, 3688, 4617);
  nand ginst1926 (5290, 3685, 4618);
  nand ginst1927 (5291, 3694, 4619);
  nand ginst1928 (5292, 3691, 4620);
  nand ginst1929 (5293, 3700, 4621);
  nand ginst1930 (5294, 3697, 4622);
  nand ginst1931 (5295, 3706, 4623);
  nand ginst1932 (5296, 3703, 4624);
  nand ginst1933 (5297, 3712, 4625);
  nand ginst1934 (5298, 3709, 4626);
  nand ginst1935 (5299, 3718, 4627);
  nand ginst1936 (5300, 3715, 4628);
  nand ginst1937 (5314, 3739, 4643);
  nand ginst1938 (5315, 3736, 4644);
  nand ginst1939 (5316, 3745, 4645);
  nand ginst1940 (5317, 3742, 4646);
  nand ginst1941 (5318, 3751, 4647);
  nand ginst1942 (5319, 3748, 4648);
  nand ginst1943 (5320, 3757, 4649);
  nand ginst1944 (5321, 3754, 4650);
  nand ginst1945 (5322, 3763, 4651);
  nand ginst1946 (5323, 3760, 4652);
  not ginst1947 (5324, 4193);
  not ginst1948 (535, 307);
  nand ginst1949 (5363, 2781, 4693);
  nand ginst1950 (5364, 3772, 4695);
  nand ginst1951 (5365, 3769, 4696);
  nand ginst1952 (5366, 3778, 4697);
  nand ginst1953 (5367, 3775, 4698);
  not ginst1954 (537, 310);
  not ginst1955 (539, 313);
  not ginst1956 (541, 316);
  nand ginst1957 (5425, 2790, 4745);
  nand ginst1958 (5426, 3813, 4747);
  nand ginst1959 (5427, 3810, 4748);
  nand ginst1960 (5429, 2793, 4750);
  not ginst1961 (543, 319);
  nand ginst1962 (5430, 3825, 4752);
  nand ginst1963 (5431, 3822, 4753);
  nand ginst1964 (5432, 3831, 4754);
  nand ginst1965 (5433, 3828, 4755);
  not ginst1966 (545, 322);
  nand ginst1967 (5451, 2796, 4775);
  nand ginst1968 (5452, 3864, 4777);
  nand ginst1969 (5453, 3861, 4778);
  nand ginst1970 (5454, 3870, 4779);
  nand ginst1971 (5455, 3867, 4780);
  nand ginst1972 (5456, 3888, 4781);
  nand ginst1973 (5457, 3885, 4782);
  not ginst1974 (5469, 4303);
  not ginst1975 (547, 325);
  nand ginst1976 (5474, 3589, 4799);
  nand ginst1977 (5475, 3586, 4800);
  nand ginst1978 (5476, 3595, 4801);
  nand ginst1979 (5477, 3592, 4802);
  not ginst1980 (549, 328);
  not ginst1981 (551, 331);
  not ginst1982 (553, 334);
  not ginst1983 (556, 337);
  nand ginst1984 (5571, 3798, 5045);
  nand ginst1985 (5572, 3795, 5046);
  nand ginst1986 (5573, 3804, 5047);
  nand ginst1987 (5574, 3801, 5048);
  nand ginst1988 (5584, 3837, 5064);
  nand ginst1989 (5585, 3834, 5065);
  nand ginst1990 (5586, 3843, 5066);
  nand ginst1991 (5587, 3840, 5067);
  not ginst1992 (559, 343);
  nand ginst1993 (5602, 3876, 5110);
  nand ginst1994 (5603, 3873, 5111);
  nand ginst1995 (5604, 3882, 5112);
  nand ginst1996 (5605, 3879, 5113);
  not ginst1997 (561, 346);
  not ginst1998 (563, 349);
  nand ginst1999 (5631, 5324, 4653);
  nand ginst2000 (5632, 4463, 5167);
  nand ginst2001 (5640, 4465, 5168);
  not ginst2002 (565, 352);
  nand ginst2003 (5654, 4467, 5169);
  not ginst2004 (567, 355);
  nand ginst2005 (5670, 4469, 5170);
  nand ginst2006 (5683, 4471, 5171);
  not ginst2007 (569, 358);
  nand ginst2008 (5690, 4475, 5172);
  nand ginst2009 (5697, 4477, 5173);
  nand ginst2010 (5707, 4479, 5174);
  not ginst2011 (571, 361);
  nand ginst2012 (5718, 4481, 5175);
  nand ginst2013 (5728, 4483, 5176);
  not ginst2014 (573, 364);
  not ginst2015 (5735, 5177);
  nand ginst2016 (5736, 5179, 4490);
  nand ginst2017 (5740, 5180, 5181);
  nand ginst2018 (5744, 5182, 5183);
  nand ginst2019 (5747, 5184, 4496);
  and ginst2020 (575, 183, 182, 185, 186);
  nand ginst2021 (5751, 5185, 5186);
  nand ginst2022 (5755, 5187, 5188);
  nand ginst2023 (5758, 5189, 4502);
  nand ginst2024 (5762, 5190, 5191);
  nand ginst2025 (5766, 5192, 5193);
  not ginst2026 (5769, 4803);
  not ginst2027 (5770, 4806);
  nand ginst2028 (5771, 4507, 5196);
  nand ginst2029 (5778, 4509, 5197);
  and ginst2030 (578, 210, 152, 218, 230);
  nand ginst2031 (5789, 4511, 5198);
  nand ginst2032 (5799, 4513, 5199);
  nand ginst2033 (5807, 4515, 5200);
  not ginst2034 (582, 15);
  nand ginst2035 (5821, 4517, 5201);
  nand ginst2036 (5837, 4519, 5202);
  not ginst2037 (585, 5);
  nand ginst2038 (5850, 4521, 5203);
  nand ginst2039 (5856, 4523, 5204);
  nand ginst2040 (5863, 4525, 5205);
  nand ginst2041 (5870, 4527, 5206);
  nand ginst2042 (5881, 4529, 5207);
  nand ginst2043 (5892, 4531, 5208);
  nand ginst2044 (5898, 4533, 5209);
  not ginst2045 (590, 1);
  nand ginst2046 (5905, 4535, 5210);
  nand ginst2047 (5915, 4537, 5211);
  nand ginst2048 (5926, 4539, 5212);
  not ginst2049 (593, 5);
  nand ginst2050 (5936, 4541, 5213);
  not ginst2051 (5943, 4817);
  nand ginst2052 (5944, 4820, 1931);
  not ginst2053 (5945, 4820);
  nand ginst2054 (5946, 4823, 1932);
  not ginst2055 (5947, 4823);
  nand ginst2056 (5948, 4826, 1933);
  not ginst2057 (5949, 4826);
  nand ginst2058 (5950, 4829, 1934);
  not ginst2059 (5951, 4829);
  nand ginst2060 (5952, 4832, 1935);
  not ginst2061 (5953, 4832);
  nand ginst2062 (5954, 4835, 1936);
  not ginst2063 (5955, 4835);
  nand ginst2064 (5956, 4838, 1937);
  not ginst2065 (5957, 4838);
  nand ginst2066 (5958, 4841, 1938);
  not ginst2067 (5959, 4841);
  not ginst2068 (596, 5);
  and ginst2069 (5960, 2674, 4769);
  not ginst2070 (5966, 4844);
  nand ginst2071 (5967, 4847, 1939);
  not ginst2072 (5968, 4847);
  nand ginst2073 (5969, 4850, 1940);
  not ginst2074 (5970, 4850);
  nand ginst2075 (5971, 4853, 1941);
  not ginst2076 (5972, 4853);
  nand ginst2077 (5973, 4856, 1942);
  not ginst2078 (5974, 4856);
  nand ginst2079 (5975, 4859, 1943);
  not ginst2080 (5976, 4859);
  nand ginst2081 (5977, 4862, 1944);
  not ginst2082 (5978, 4862);
  nand ginst2083 (5979, 4865, 1945);
  not ginst2084 (5980, 4865);
  and ginst2085 (5981, 2674, 4769);
  nand ginst2086 (5989, 4868, 1946);
  not ginst2087 (599, 289);
  not ginst2088 (5990, 4868);
  nand ginst2089 (5991, 5283, 5284);
  nand ginst2090 (5996, 5285, 5286);
  nand ginst2091 (6000, 5287, 5288);
  nand ginst2092 (6003, 5289, 5290);
  nand ginst2093 (6009, 5291, 5292);
  nand ginst2094 (6014, 5293, 5294);
  nand ginst2095 (6018, 5295, 5296);
  nand ginst2096 (6021, 5297, 5298);
  nand ginst2097 (6022, 5299, 5300);
  not ginst2098 (6023, 4874);
  nand ginst2099 (6024, 4874, 4629);
  not ginst2100 (6025, 4877);
  nand ginst2101 (6026, 4877, 4631);
  not ginst2102 (6027, 4880);
  nand ginst2103 (6028, 4880, 4633);
  not ginst2104 (6029, 4883);
  nand ginst2105 (6030, 4883, 4636);
  not ginst2106 (6031, 4886);
  not ginst2107 (6032, 4889);
  not ginst2108 (6033, 4892);
  not ginst2109 (6034, 4895);
  not ginst2110 (6035, 4898);
  not ginst2111 (6036, 4901);
  not ginst2112 (6037, 4904);
  nand ginst2113 (6038, 4904, 4642);
  not ginst2114 (6039, 4907);
  not ginst2115 (604, 299);
  not ginst2116 (6040, 4910);
  nand ginst2117 (6041, 5314, 5315);
  nand ginst2118 (6047, 5316, 5317);
  nand ginst2119 (6052, 5318, 5319);
  nand ginst2120 (6056, 5320, 5321);
  nand ginst2121 (6059, 5322, 5323);
  nand ginst2122 (6060, 4913, 1968);
  not ginst2123 (6061, 4913);
  nand ginst2124 (6062, 4916, 1969);
  not ginst2125 (6063, 4916);
  nand ginst2126 (6064, 4919, 1970);
  not ginst2127 (6065, 4919);
  nand ginst2128 (6066, 4922, 1971);
  not ginst2129 (6067, 4922);
  nand ginst2130 (6068, 4925, 1972);
  not ginst2131 (6069, 4925);
  nand ginst2132 (6070, 4928, 1973);
  not ginst2133 (6071, 4928);
  nand ginst2134 (6072, 4931, 1974);
  not ginst2135 (6073, 4931);
  nand ginst2136 (6074, 4934, 1975);
  not ginst2137 (6075, 4934);
  nand ginst2138 (6076, 4937, 1976);
  not ginst2139 (6077, 4937);
  not ginst2140 (6078, 4940);
  nand ginst2141 (6079, 5363, 4694);
  nand ginst2142 (6083, 5364, 5365);
  nand ginst2143 (6087, 5366, 5367);
  not ginst2144 (609, 303);
  not ginst2145 (6090, 4943);
  nand ginst2146 (6091, 4943, 4699);
  not ginst2147 (6092, 4946);
  not ginst2148 (6093, 4949);
  not ginst2149 (6094, 4952);
  not ginst2150 (6095, 4955);
  not ginst2151 (6096, 4970);
  nand ginst2152 (6097, 4970, 4700);
  not ginst2153 (6098, 4973);
  not ginst2154 (6099, 4976);
  not ginst2155 (6100, 4979);
  not ginst2156 (6101, 4982);
  not ginst2157 (6102, 4997);
  nand ginst2158 (6103, 5000, 2015);
  not ginst2159 (6104, 5000);
  nand ginst2160 (6105, 5003, 2016);
  not ginst2161 (6106, 5003);
  nand ginst2162 (6107, 5006, 2017);
  not ginst2163 (6108, 5006);
  nand ginst2164 (6109, 5009, 2018);
  not ginst2165 (6110, 5009);
  nand ginst2166 (6111, 5012, 2019);
  not ginst2167 (6112, 5012);
  nand ginst2168 (6113, 5015, 2020);
  not ginst2169 (6114, 5015);
  nand ginst2170 (6115, 5018, 2021);
  not ginst2171 (6116, 5018);
  nand ginst2172 (6117, 5021, 2022);
  not ginst2173 (6118, 5021);
  nand ginst2174 (6119, 5024, 2023);
  not ginst2175 (6120, 5024);
  not ginst2176 (6121, 5033);
  nand ginst2177 (6122, 5033, 4743);
  not ginst2178 (6123, 5036);
  not ginst2179 (6124, 5039);
  nand ginst2180 (6125, 5042, 4744);
  not ginst2181 (6126, 5042);
  nand ginst2182 (6127, 5425, 4746);
  nand ginst2183 (6131, 5426, 5427);
  not ginst2184 (6135, 5049);
  nand ginst2185 (6136, 5049, 4749);
  nand ginst2186 (6137, 5429, 4751);
  not ginst2187 (614, 38);
  nand ginst2188 (6141, 5430, 5431);
  nand ginst2189 (6145, 5432, 5433);
  not ginst2190 (6148, 5068);
  not ginst2191 (6149, 5071);
  not ginst2192 (6150, 5074);
  not ginst2193 (6151, 5077);
  not ginst2194 (6152, 5080);
  not ginst2195 (6153, 5083);
  not ginst2196 (6154, 5086);
  not ginst2197 (6155, 5089);
  not ginst2198 (6156, 5092);
  nand ginst2199 (6157, 5092, 4761);
  not ginst2200 (6158, 5095);
  nand ginst2201 (6159, 5095, 4763);
  not ginst2202 (6160, 5098);
  nand ginst2203 (6161, 5098, 4765);
  not ginst2204 (6162, 5101);
  not ginst2205 (6163, 5104);
  nand ginst2206 (6164, 5107, 4768);
  not ginst2207 (6165, 5107);
  nand ginst2208 (6166, 5451, 4776);
  nand ginst2209 (6170, 5452, 5453);
  nand ginst2210 (6174, 5454, 5455);
  nand ginst2211 (6177, 5456, 5457);
  not ginst2212 (6181, 5114);
  not ginst2213 (6182, 5117);
  not ginst2214 (6183, 5120);
  not ginst2215 (6184, 5123);
  not ginst2216 (6185, 5138);
  nand ginst2217 (6186, 5138, 4783);
  not ginst2218 (6187, 5141);
  not ginst2219 (6188, 5144);
  not ginst2220 (6189, 5147);
  not ginst2221 (6190, 5150);
  not ginst2222 (6191, 4784);
  nand ginst2223 (6192, 4784, 2230);
  not ginst2224 (6193, 4790);
  nand ginst2225 (6194, 4790, 2765);
  not ginst2226 (6195, 4796);
  nand ginst2227 (6196, 5476, 5477);
  nand ginst2228 (6199, 5474, 5475);
  not ginst2229 (6202, 4810);
  not ginst2230 (6203, 4814);
  not ginst2231 (6204, 4769);
  not ginst2232 (6207, 4555);
  not ginst2233 (6210, 4769);
  not ginst2234 (6213, 4871);
  not ginst2235 (6214, 4586);
  nor ginst2236 (6217, 2674, 4769);
  not ginst2237 (6220, 4667);
  not ginst2238 (6223, 4958);
  not ginst2239 (6224, 4961);
  not ginst2240 (6225, 4964);
  not ginst2241 (6226, 4967);
  not ginst2242 (6227, 4985);
  not ginst2243 (6228, 4988);
  not ginst2244 (6229, 4991);
  not ginst2245 (6230, 4994);
  not ginst2246 (6231, 5027);
  not ginst2247 (6232, 4711);
  not ginst2248 (6235, 5030);
  not ginst2249 (6236, 4735);
  not ginst2250 (6239, 5052);
  not ginst2251 (6240, 5055);
  not ginst2252 (6241, 5058);
  not ginst2253 (6242, 5061);
  nand ginst2254 (6243, 5573, 5574);
  nand ginst2255 (6246, 5571, 5572);
  nand ginst2256 (6249, 5586, 5587);
  not ginst2257 (625, 15);
  nand ginst2258 (6252, 5584, 5585);
  not ginst2259 (6255, 5126);
  not ginst2260 (6256, 5129);
  not ginst2261 (6257, 5132);
  not ginst2262 (6258, 5135);
  not ginst2263 (6259, 5153);
  not ginst2264 (6260, 5156);
  not ginst2265 (6261, 5159);
  not ginst2266 (6262, 5162);
  nand ginst2267 (6263, 5604, 5605);
  nand ginst2268 (6266, 5602, 5603);
  nand ginst2269 (628, 12, 9);
  nand ginst2270 (632, 12, 9);
  not ginst2271 (636, 38);
  not ginst2272 (641, 245);
  not ginst2273 (642, 248);
  not ginst2274 (643, 251);
  not ginst2275 (644, 251);
  not ginst2276 (651, 254);
  nand ginst2277 (6540, 1380, 5945);
  nand ginst2278 (6541, 1383, 5947);
  nand ginst2279 (6542, 1386, 5949);
  nand ginst2280 (6543, 1389, 5951);
  nand ginst2281 (6544, 1392, 5953);
  nand ginst2282 (6545, 1395, 5955);
  nand ginst2283 (6546, 1398, 5957);
  nand ginst2284 (6547, 1401, 5959);
  nand ginst2285 (6555, 1404, 5968);
  nand ginst2286 (6556, 1407, 5970);
  nand ginst2287 (6557, 1410, 5972);
  nand ginst2288 (6558, 1413, 5974);
  nand ginst2289 (6559, 1416, 5976);
  nand ginst2290 (6560, 1419, 5978);
  nand ginst2291 (6561, 1422, 5980);
  nand ginst2292 (6569, 1425, 5990);
  not ginst2293 (657, 106);
  nand ginst2294 (6594, 3721, 6023);
  nand ginst2295 (6595, 3724, 6025);
  nand ginst2296 (6596, 3727, 6027);
  nand ginst2297 (6597, 3730, 6029);
  nand ginst2298 (6598, 4889, 6031);
  nand ginst2299 (6599, 4886, 6032);
  not ginst2300 (660, 257);
  nand ginst2301 (6600, 4895, 6033);
  nand ginst2302 (6601, 4892, 6034);
  nand ginst2303 (6602, 4901, 6035);
  nand ginst2304 (6603, 4898, 6036);
  nand ginst2305 (6604, 3733, 6037);
  nand ginst2306 (6605, 4910, 6039);
  nand ginst2307 (6606, 4907, 6040);
  nand ginst2308 (6621, 1434, 6061);
  nand ginst2309 (6622, 1437, 6063);
  nand ginst2310 (6623, 1440, 6065);
  nand ginst2311 (6624, 1443, 6067);
  nand ginst2312 (6625, 1446, 6069);
  nand ginst2313 (6626, 1449, 6071);
  nand ginst2314 (6627, 1452, 6073);
  nand ginst2315 (6628, 1455, 6075);
  nand ginst2316 (6629, 1458, 6077);
  nand ginst2317 (6639, 3783, 6090);
  nand ginst2318 (6640, 4949, 6092);
  nand ginst2319 (6641, 4946, 6093);
  nand ginst2320 (6642, 4955, 6094);
  nand ginst2321 (6643, 4952, 6095);
  nand ginst2322 (6644, 3786, 6096);
  nand ginst2323 (6645, 4976, 6098);
  nand ginst2324 (6646, 4973, 6099);
  nand ginst2325 (6647, 4982, 6100);
  nand ginst2326 (6648, 4979, 6101);
  nand ginst2327 (6649, 1461, 6104);
  nand ginst2328 (6650, 1464, 6106);
  nand ginst2329 (6651, 1467, 6108);
  nand ginst2330 (6652, 1470, 6110);
  nand ginst2331 (6653, 1473, 6112);
  nand ginst2332 (6654, 1476, 6114);
  nand ginst2333 (6655, 1479, 6116);
  nand ginst2334 (6656, 1482, 6118);
  nand ginst2335 (6657, 1485, 6120);
  nand ginst2336 (6658, 3789, 6121);
  nand ginst2337 (6659, 5039, 6123);
  not ginst2338 (666, 260);
  nand ginst2339 (6660, 5036, 6124);
  nand ginst2340 (6661, 3792, 6126);
  nand ginst2341 (6668, 3816, 6135);
  nand ginst2342 (6677, 5071, 6148);
  nand ginst2343 (6678, 5068, 6149);
  nand ginst2344 (6679, 5077, 6150);
  nand ginst2345 (6680, 5074, 6151);
  nand ginst2346 (6681, 5083, 6152);
  nand ginst2347 (6682, 5080, 6153);
  nand ginst2348 (6683, 5089, 6154);
  nand ginst2349 (6684, 5086, 6155);
  nand ginst2350 (6685, 3846, 6156);
  nand ginst2351 (6686, 3849, 6158);
  nand ginst2352 (6687, 3852, 6160);
  nand ginst2353 (6688, 5104, 6162);
  nand ginst2354 (6689, 5101, 6163);
  nand ginst2355 (6690, 3855, 6165);
  nand ginst2356 (6702, 5117, 6181);
  nand ginst2357 (6703, 5114, 6182);
  nand ginst2358 (6704, 5123, 6183);
  nand ginst2359 (6705, 5120, 6184);
  nand ginst2360 (6706, 3891, 6185);
  nand ginst2361 (6707, 5144, 6187);
  nand ginst2362 (6708, 5141, 6188);
  nand ginst2363 (6709, 5150, 6189);
  nand ginst2364 (6710, 5147, 6190);
  nand ginst2365 (6711, 1708, 6191);
  nand ginst2366 (6712, 2231, 6193);
  not ginst2367 (672, 263);
  nand ginst2368 (6729, 4961, 6223);
  not ginst2369 (673, 267);
  nand ginst2370 (6730, 4958, 6224);
  nand ginst2371 (6731, 4967, 6225);
  nand ginst2372 (6732, 4964, 6226);
  nand ginst2373 (6733, 4988, 6227);
  nand ginst2374 (6734, 4985, 6228);
  nand ginst2375 (6735, 4994, 6229);
  nand ginst2376 (6736, 4991, 6230);
  not ginst2377 (674, 106);
  nand ginst2378 (6741, 5055, 6239);
  nand ginst2379 (6742, 5052, 6240);
  nand ginst2380 (6743, 5061, 6241);
  nand ginst2381 (6744, 5058, 6242);
  nand ginst2382 (6751, 5129, 6255);
  nand ginst2383 (6752, 5126, 6256);
  nand ginst2384 (6753, 5135, 6257);
  nand ginst2385 (6754, 5132, 6258);
  nand ginst2386 (6755, 5156, 6259);
  nand ginst2387 (6756, 5153, 6260);
  nand ginst2388 (6757, 5162, 6261);
  nand ginst2389 (6758, 5159, 6262);
  not ginst2390 (676, 18);
  not ginst2391 (6761, 5892);
  and ginst2392 (6762, 5683, 5670, 5654, 5640, 5632);
  and ginst2393 (6766, 5632, 3097);
  and ginst2394 (6767, 5640, 5632, 3101);
  and ginst2395 (6768, 5654, 5632, 3107, 5640);
  and ginst2396 (6769, 5670, 5654, 5632, 3114, 5640);
  and ginst2397 (6770, 5640, 3101);
  and ginst2398 (6771, 5654, 3107, 5640);
  and ginst2399 (6772, 5670, 5654, 3114, 5640);
  and ginst2400 (6773, 5683, 5654, 5640, 5670);
  and ginst2401 (6774, 5640, 3101);
  and ginst2402 (6775, 5654, 3107, 5640);
  and ginst2403 (6776, 5670, 5654, 3114, 5640);
  and ginst2404 (6777, 5654, 3107);
  and ginst2405 (6778, 5670, 5654, 3114);
  and ginst2406 (6779, 5683, 5654, 5670);
  and ginst2407 (6780, 5654, 3107);
  and ginst2408 (6781, 5670, 5654, 3114);
  and ginst2409 (6782, 5670, 3114);
  and ginst2410 (6783, 5683, 5670);
  and ginst2411 (6784, 5697, 5728, 5707, 5690, 5718);
  and ginst2412 (6787, 5690, 3137);
  and ginst2413 (6788, 5697, 5690, 3140);
  and ginst2414 (6789, 5707, 5690, 3144, 5697);
  and ginst2415 (6790, 5718, 5707, 5690, 3149, 5697);
  and ginst2416 (6791, 5697, 3140);
  and ginst2417 (6792, 5707, 3144, 5697);
  and ginst2418 (6793, 5718, 5707, 3149, 5697);
  and ginst2419 (6794, 3144, 5707);
  and ginst2420 (6795, 5718, 5707, 3149);
  and ginst2421 (6796, 5718, 3149);
  not ginst2422 (6797, 5736);
  not ginst2423 (6800, 5740);
  not ginst2424 (6803, 5747);
  not ginst2425 (6806, 5751);
  not ginst2426 (6809, 5758);
  not ginst2427 (6812, 5762);
  not ginst2428 (6815, 5744);
  not ginst2429 (6818, 5744);
  not ginst2430 (682, 18);
  not ginst2431 (6821, 5755);
  not ginst2432 (6824, 5755);
  not ginst2433 (6827, 5766);
  not ginst2434 (6830, 5766);
  and ginst2435 (6833, 5850, 5789, 5778, 5771);
  and ginst2436 (6836, 5771, 3169);
  and ginst2437 (6837, 5778, 5771, 3173);
  and ginst2438 (6838, 5789, 5771, 3178, 5778);
  and ginst2439 (6839, 5778, 3173);
  and ginst2440 (6840, 5789, 3178, 5778);
  and ginst2441 (6841, 5850, 5789, 5778);
  and ginst2442 (6842, 5778, 3173);
  and ginst2443 (6843, 5789, 3178, 5778);
  and ginst2444 (6844, 5789, 3178);
  and ginst2445 (6845, 5856, 5837, 5821, 5807, 5799);
  and ginst2446 (6848, 5799, 3185);
  and ginst2447 (6849, 5807, 5799, 3189);
  and ginst2448 (6850, 5821, 5799, 3195, 5807);
  and ginst2449 (6851, 5837, 5821, 5799, 3202, 5807);
  and ginst2450 (6852, 5807, 3189);
  and ginst2451 (6853, 5821, 3195, 5807);
  and ginst2452 (6854, 5837, 5821, 3202, 5807);
  and ginst2453 (6855, 5856, 5821, 5807, 5837);
  and ginst2454 (6856, 5807, 3189);
  and ginst2455 (6857, 5821, 3195, 5807);
  and ginst2456 (6858, 5837, 5821, 3202, 5807);
  and ginst2457 (6859, 5821, 3195);
  and ginst2458 (6860, 5837, 5821, 3202);
  and ginst2459 (6861, 5856, 5821, 5837);
  and ginst2460 (6862, 5821, 3195);
  and ginst2461 (6863, 5837, 5821, 3202);
  and ginst2462 (6864, 5837, 3202);
  and ginst2463 (6865, 5850, 5789);
  and ginst2464 (6866, 5856, 5837);
  and ginst2465 (6867, 5870, 5892, 5881, 5863);
  and ginst2466 (6870, 5863, 3211);
  and ginst2467 (6871, 5870, 5863, 3215);
  and ginst2468 (6872, 5881, 5863, 3221, 5870);
  and ginst2469 (6873, 5870, 3215);
  and ginst2470 (6874, 5881, 3221, 5870);
  and ginst2471 (6875, 5892, 5881, 5870);
  and ginst2472 (6876, 5870, 3215);
  and ginst2473 (6877, 3221, 5881, 5870);
  and ginst2474 (6878, 5881, 3221);
  and ginst2475 (6879, 5892, 5881);
  and ginst2476 (688, 382, 263);
  and ginst2477 (6880, 5881, 3221);
  and ginst2478 (6881, 5905, 5936, 5915, 5898, 5926);
  and ginst2479 (6884, 5898, 3229);
  and ginst2480 (6885, 5905, 5898, 3232);
  and ginst2481 (6886, 5915, 5898, 3236, 5905);
  and ginst2482 (6887, 5926, 5915, 5898, 3241, 5905);
  and ginst2483 (6888, 5905, 3232);
  and ginst2484 (6889, 5915, 3236, 5905);
  not ginst2485 (689, 18);
  and ginst2486 (6890, 5926, 5915, 3241, 5905);
  and ginst2487 (6891, 3236, 5915);
  and ginst2488 (6892, 5926, 5915, 3241);
  and ginst2489 (6893, 5926, 3241);
  nand ginst2490 (6894, 5944, 6540);
  nand ginst2491 (6901, 5946, 6541);
  nand ginst2492 (6912, 5948, 6542);
  nand ginst2493 (6923, 5950, 6543);
  nand ginst2494 (6929, 5952, 6544);
  nand ginst2495 (6936, 5954, 6545);
  nand ginst2496 (6946, 5956, 6546);
  not ginst2497 (695, 18);
  nand ginst2498 (6957, 5958, 6547);
  nand ginst2499 (6967, 6204, 4575);
  not ginst2500 (6968, 6204);
  not ginst2501 (6969, 6207);
  nand ginst2502 (6970, 5967, 6555);
  nand ginst2503 (6977, 5969, 6556);
  nand ginst2504 (6988, 5971, 6557);
  nand ginst2505 (6998, 5973, 6558);
  nand ginst2506 (700, 382, 267);
  nand ginst2507 (7006, 5975, 6559);
  nand ginst2508 (7020, 5977, 6560);
  nand ginst2509 (7036, 5979, 6561);
  nand ginst2510 (7049, 5989, 6569);
  not ginst2511 (705, 271);
  nand ginst2512 (7055, 6210, 4610);
  not ginst2513 (7056, 6210);
  and ginst2514 (7057, 6021, 6000, 5996, 5991);
  not ginst2515 (706, 274);
  and ginst2516 (7060, 5991, 3362);
  and ginst2517 (7061, 5996, 5991, 3363);
  and ginst2518 (7062, 6000, 5991, 3364, 5996);
  and ginst2519 (7063, 6022, 6018, 6014, 6009, 6003);
  and ginst2520 (7064, 6003, 3366);
  and ginst2521 (7065, 6009, 6003, 3367);
  and ginst2522 (7066, 6014, 6003, 3368, 6009);
  and ginst2523 (7067, 6018, 6014, 6003, 3369, 6009);
  nand ginst2524 (7068, 6594, 6024);
  not ginst2525 (707, 277);
  nand ginst2526 (7073, 6595, 6026);
  nand ginst2527 (7077, 6596, 6028);
  not ginst2528 (708, 277);
  nand ginst2529 (7080, 6597, 6030);
  nand ginst2530 (7086, 6598, 6599);
  nand ginst2531 (7091, 6600, 6601);
  nand ginst2532 (7095, 6602, 6603);
  nand ginst2533 (7098, 6604, 6038);
  nand ginst2534 (7099, 6605, 6606);
  and ginst2535 (7100, 6059, 6056, 6052, 6047, 6041);
  and ginst2536 (7103, 6041, 3371);
  and ginst2537 (7104, 6047, 6041, 3372);
  and ginst2538 (7105, 6052, 6041, 3373, 6047);
  and ginst2539 (7106, 6056, 6052, 6041, 3374, 6047);
  nand ginst2540 (7107, 6060, 6621);
  nand ginst2541 (7114, 6062, 6622);
  nand ginst2542 (7125, 6064, 6623);
  nand ginst2543 (7136, 6066, 6624);
  nand ginst2544 (7142, 6068, 6625);
  nand ginst2545 (7149, 6070, 6626);
  not ginst2546 (715, 280);
  nand ginst2547 (7159, 6072, 6627);
  nand ginst2548 (7170, 6074, 6628);
  nand ginst2549 (7180, 6076, 6629);
  not ginst2550 (7187, 6220);
  not ginst2551 (7188, 6079);
  not ginst2552 (7191, 6083);
  nand ginst2553 (7194, 6639, 6091);
  nand ginst2554 (7198, 6640, 6641);
  nand ginst2555 (7202, 6642, 6643);
  nand ginst2556 (7205, 6644, 6097);
  nand ginst2557 (7209, 6645, 6646);
  not ginst2558 (721, 283);
  nand ginst2559 (7213, 6647, 6648);
  not ginst2560 (7216, 6087);
  not ginst2561 (7219, 6087);
  nand ginst2562 (7222, 6103, 6649);
  nand ginst2563 (7229, 6105, 6650);
  nand ginst2564 (7240, 6107, 6651);
  nand ginst2565 (7250, 6109, 6652);
  nand ginst2566 (7258, 6111, 6653);
  not ginst2567 (727, 286);
  nand ginst2568 (7272, 6113, 6654);
  nand ginst2569 (7288, 6115, 6655);
  nand ginst2570 (7301, 6117, 6656);
  nand ginst2571 (7307, 6119, 6657);
  nand ginst2572 (7314, 6658, 6122);
  nand ginst2573 (7318, 6659, 6660);
  nand ginst2574 (7322, 6125, 6661);
  not ginst2575 (7325, 6127);
  not ginst2576 (7328, 6131);
  not ginst2577 (733, 289);
  nand ginst2578 (7331, 6668, 6136);
  not ginst2579 (7334, 6137);
  not ginst2580 (7337, 6141);
  not ginst2581 (734, 293);
  not ginst2582 (7340, 6145);
  not ginst2583 (7343, 6145);
  nand ginst2584 (7346, 6677, 6678);
  nand ginst2585 (7351, 6679, 6680);
  nand ginst2586 (7355, 6681, 6682);
  nand ginst2587 (7358, 6683, 6684);
  nand ginst2588 (7364, 6685, 6157);
  nand ginst2589 (7369, 6686, 6159);
  nand ginst2590 (7373, 6687, 6161);
  nand ginst2591 (7376, 6688, 6689);
  nand ginst2592 (7377, 6164, 6690);
  not ginst2593 (7378, 6166);
  not ginst2594 (7381, 6170);
  not ginst2595 (7384, 6177);
  nand ginst2596 (7387, 6702, 6703);
  nand ginst2597 (7391, 6704, 6705);
  nand ginst2598 (7394, 6706, 6186);
  nand ginst2599 (7398, 6707, 6708);
  nand ginst2600 (7402, 6709, 6710);
  not ginst2601 (7405, 6174);
  not ginst2602 (7408, 6174);
  not ginst2603 (7411, 5936);
  not ginst2604 (7414, 5898);
  not ginst2605 (7417, 5905);
  not ginst2606 (742, 296);
  not ginst2607 (7420, 5915);
  not ginst2608 (7423, 5926);
  not ginst2609 (7426, 5728);
  not ginst2610 (7429, 5690);
  not ginst2611 (7432, 5697);
  not ginst2612 (7435, 5707);
  not ginst2613 (7438, 5718);
  nand ginst2614 (7441, 6192, 6711);
  nand ginst2615 (7444, 6194, 6712);
  not ginst2616 (7447, 5683);
  not ginst2617 (7450, 5670);
  not ginst2618 (7453, 5632);
  not ginst2619 (7456, 5654);
  not ginst2620 (7459, 5640);
  not ginst2621 (7462, 5640);
  not ginst2622 (7465, 5683);
  not ginst2623 (7468, 5670);
  not ginst2624 (7471, 5632);
  not ginst2625 (7474, 5654);
  not ginst2626 (7477, 6196);
  not ginst2627 (7478, 6199);
  not ginst2628 (7479, 5850);
  not ginst2629 (748, 299);
  not ginst2630 (7482, 5789);
  not ginst2631 (7485, 5771);
  not ginst2632 (7488, 5778);
  not ginst2633 (749, 303);
  not ginst2634 (7491, 5850);
  not ginst2635 (7494, 5789);
  not ginst2636 (7497, 5771);
  not ginst2637 (750, 367);
  not ginst2638 (7500, 5778);
  not ginst2639 (7503, 5856);
  not ginst2640 (7506, 5837);
  not ginst2641 (7509, 5799);
  not ginst2642 (7512, 5821);
  not ginst2643 (7515, 5807);
  not ginst2644 (7518, 5807);
  not ginst2645 (7521, 5856);
  not ginst2646 (7524, 5837);
  not ginst2647 (7527, 5799);
  not ginst2648 (7530, 5821);
  not ginst2649 (7533, 5863);
  not ginst2650 (7536, 5863);
  not ginst2651 (7539, 5870);
  not ginst2652 (7542, 5870);
  not ginst2653 (7545, 5881);
  not ginst2654 (7548, 5881);
  not ginst2655 (7551, 6214);
  not ginst2656 (7552, 6217);
  not ginst2657 (7553, 5981);
  not ginst2658 (7556, 6249);
  not ginst2659 (7557, 6252);
  not ginst2660 (7558, 6243);
  not ginst2661 (7559, 6246);
  nand ginst2662 (7560, 6731, 6732);
  nand ginst2663 (7563, 6729, 6730);
  nand ginst2664 (7566, 6735, 6736);
  nand ginst2665 (7569, 6733, 6734);
  not ginst2666 (7572, 6232);
  not ginst2667 (7573, 6236);
  nand ginst2668 (7574, 6743, 6744);
  nand ginst2669 (7577, 6741, 6742);
  not ginst2670 (758, 307);
  not ginst2671 (7580, 6263);
  not ginst2672 (7581, 6266);
  nand ginst2673 (7582, 6753, 6754);
  nand ginst2674 (7585, 6751, 6752);
  nand ginst2675 (7588, 6757, 6758);
  not ginst2676 (759, 310);
  nand ginst2677 (7591, 6755, 6756);
  or ginst2678 (7609, 3096, 6766, 6767, 6768, 6769);
  or ginst2679 (7613, 3107, 6782);
  not ginst2680 (762, 313);
  or ginst2681 (7620, 3136, 6787, 6788, 6789, 6790);
  or ginst2682 (7649, 3168, 6836, 6837, 6838);
  or ginst2683 (7650, 3173, 6844);
  or ginst2684 (7655, 3184, 6848, 6849, 6850, 6851);
  or ginst2685 (7659, 3195, 6864);
  or ginst2686 (7668, 3210, 6870, 6871, 6872);
  or ginst2687 (7671, 3228, 6884, 6885, 6886, 6887);
  not ginst2688 (768, 316);
  not ginst2689 (774, 319);
  nand ginst2690 (7744, 3661, 6968);
  not ginst2691 (780, 322);
  nand ginst2692 (7822, 3664, 7056);
  or ginst2693 (7825, 3361, 7060, 7061, 7062);
  or ginst2694 (7826, 3365, 7064, 7065, 7066, 7067);
  or ginst2695 (7852, 3370, 7103, 7104, 7105, 7106);
  not ginst2696 (786, 325);
  not ginst2697 (794, 328);
  not ginst2698 (800, 331);
  not ginst2699 (806, 334);
  or ginst2700 (8114, 3101, 6777, 6778, 6779);
  or ginst2701 (8117, 3097, 6770, 6771, 6772, 6773);
  not ginst2702 (812, 337);
  not ginst2703 (813, 340);
  nor ginst2704 (8131, 3101, 6780, 6781);
  nor ginst2705 (8134, 3097, 6774, 6775, 6776);
  not ginst2706 (814, 340);
  nand ginst2707 (8144, 6199, 7477);
  nand ginst2708 (8145, 6196, 7478);
  or ginst2709 (8146, 3169, 6839, 6840, 6841);
  nor ginst2710 (8156, 3169, 6842, 6843);
  or ginst2711 (8166, 3189, 6859, 6860, 6861);
  or ginst2712 (8169, 3185, 6852, 6853, 6854, 6855);
  nor ginst2713 (8183, 3189, 6862, 6863);
  nor ginst2714 (8186, 3185, 6856, 6857, 6858);
  or ginst2715 (8196, 3211, 6873, 6874, 6875);
  nor ginst2716 (8200, 3211, 6876, 6877);
  or ginst2717 (8204, 3215, 6878, 6879);
  nor ginst2718 (8208, 3215, 6880);
  not ginst2719 (821, 343);
  nand ginst2720 (8216, 6252, 7556);
  nand ginst2721 (8217, 6249, 7557);
  nand ginst2722 (8218, 6246, 7558);
  nand ginst2723 (8219, 6243, 7559);
  nand ginst2724 (8232, 6266, 7580);
  nand ginst2725 (8233, 6263, 7581);
  not ginst2726 (8242, 7411);
  not ginst2727 (8243, 7414);
  not ginst2728 (8244, 7417);
  not ginst2729 (8245, 7420);
  not ginst2730 (8246, 7423);
  not ginst2731 (8247, 7426);
  not ginst2732 (8248, 7429);
  not ginst2733 (8249, 7432);
  not ginst2734 (8250, 7435);
  not ginst2735 (8251, 7438);
  not ginst2736 (8252, 7136);
  not ginst2737 (8253, 6923);
  not ginst2738 (8254, 6762);
  not ginst2739 (8260, 7459);
  not ginst2740 (8261, 7462);
  and ginst2741 (8262, 3122, 6762);
  and ginst2742 (8269, 3155, 6784);
  not ginst2743 (827, 346);
  not ginst2744 (8274, 6815);
  not ginst2745 (8275, 6818);
  not ginst2746 (8276, 6821);
  not ginst2747 (8277, 6824);
  not ginst2748 (8278, 6827);
  not ginst2749 (8279, 6830);
  and ginst2750 (8280, 5740, 5736, 6815);
  and ginst2751 (8281, 6800, 6797, 6818);
  and ginst2752 (8282, 5751, 5747, 6821);
  and ginst2753 (8283, 6806, 6803, 6824);
  and ginst2754 (8284, 5762, 5758, 6827);
  and ginst2755 (8285, 6812, 6809, 6830);
  not ginst2756 (8288, 6845);
  not ginst2757 (8294, 7488);
  not ginst2758 (8295, 7500);
  not ginst2759 (8296, 7515);
  not ginst2760 (8297, 7518);
  and ginst2761 (8298, 6833, 6845);
  and ginst2762 (8307, 6867, 6881);
  not ginst2763 (8315, 7533);
  not ginst2764 (8317, 7536);
  not ginst2765 (8319, 7539);
  not ginst2766 (8321, 7542);
  nand ginst2767 (8322, 7545, 4543);
  not ginst2768 (8323, 7545);
  nand ginst2769 (8324, 7548, 5943);
  not ginst2770 (8325, 7548);
  nand ginst2771 (8326, 6967, 7744);
  not ginst2772 (833, 349);
  and ginst2773 (8333, 6901, 6923, 6912, 6894);
  and ginst2774 (8337, 6894, 4545);
  and ginst2775 (8338, 6901, 6894, 4549);
  and ginst2776 (8339, 6912, 6894, 4555, 6901);
  and ginst2777 (8340, 6901, 4549);
  and ginst2778 (8341, 6912, 4555, 6901);
  and ginst2779 (8342, 6923, 6912, 6901);
  and ginst2780 (8343, 6901, 4549);
  and ginst2781 (8344, 4555, 6912, 6901);
  and ginst2782 (8345, 6912, 4555);
  and ginst2783 (8346, 6923, 6912);
  and ginst2784 (8347, 6912, 4555);
  and ginst2785 (8348, 6929, 4563);
  and ginst2786 (8349, 6936, 6929, 4566);
  and ginst2787 (8350, 6946, 6929, 4570, 6936);
  and ginst2788 (8351, 6957, 6946, 6929, 5960, 6936);
  and ginst2789 (8352, 6936, 4566);
  and ginst2790 (8353, 6946, 4570, 6936);
  and ginst2791 (8354, 6957, 6946, 5960, 6936);
  and ginst2792 (8355, 4570, 6946);
  and ginst2793 (8356, 6957, 6946, 5960);
  and ginst2794 (8357, 6957, 5960);
  nand ginst2795 (8358, 7055, 7822);
  and ginst2796 (8365, 7049, 6988, 6977, 6970);
  and ginst2797 (8369, 6970, 4577);
  and ginst2798 (8370, 6977, 6970, 4581);
  and ginst2799 (8371, 6988, 6970, 4586, 6977);
  and ginst2800 (8372, 6977, 4581);
  and ginst2801 (8373, 6988, 4586, 6977);
  and ginst2802 (8374, 7049, 6988, 6977);
  and ginst2803 (8375, 6977, 4581);
  and ginst2804 (8376, 6988, 4586, 6977);
  and ginst2805 (8377, 6988, 4586);
  and ginst2806 (8378, 6998, 4593);
  and ginst2807 (8379, 7006, 6998, 4597);
  and ginst2808 (8380, 7020, 6998, 4603, 7006);
  and ginst2809 (8381, 7036, 7020, 6998, 5981, 7006);
  and ginst2810 (8382, 7006, 4597);
  and ginst2811 (8383, 7020, 4603, 7006);
  and ginst2812 (8384, 7036, 7020, 5981, 7006);
  and ginst2813 (8385, 7006, 4597);
  and ginst2814 (8386, 7020, 4603, 7006);
  and ginst2815 (8387, 7036, 7020, 5981, 7006);
  and ginst2816 (8388, 7020, 4603);
  and ginst2817 (8389, 7036, 7020, 5981);
  not ginst2818 (839, 352);
  and ginst2819 (8390, 7020, 4603);
  and ginst2820 (8391, 7036, 7020, 5981);
  and ginst2821 (8392, 7036, 5981);
  and ginst2822 (8393, 7049, 6988);
  and ginst2823 (8394, 7057, 7063);
  and ginst2824 (8404, 7057, 7826);
  and ginst2825 (8405, 7098, 7077, 7073, 7068);
  and ginst2826 (8409, 7068, 4632);
  and ginst2827 (8410, 7073, 7068, 4634);
  and ginst2828 (8411, 7077, 7068, 4635, 7073);
  and ginst2829 (8412, 7099, 7095, 7091, 7086, 7080);
  and ginst2830 (8415, 7080, 4638);
  and ginst2831 (8416, 7086, 7080, 4639);
  and ginst2832 (8417, 7091, 7080, 4640, 7086);
  and ginst2833 (8418, 7095, 7091, 7080, 4641, 7086);
  and ginst2834 (8421, 3375, 7100);
  and ginst2835 (8430, 7114, 7136, 7125, 7107);
  and ginst2836 (8433, 7107, 4657);
  and ginst2837 (8434, 7114, 7107, 4661);
  and ginst2838 (8435, 7125, 7107, 4667, 7114);
  and ginst2839 (8436, 7114, 4661);
  and ginst2840 (8437, 7125, 4667, 7114);
  and ginst2841 (8438, 7136, 7125, 7114);
  and ginst2842 (8439, 7114, 4661);
  and ginst2843 (8440, 4667, 7125, 7114);
  and ginst2844 (8441, 7125, 4667);
  and ginst2845 (8442, 7136, 7125);
  and ginst2846 (8443, 7125, 4667);
  and ginst2847 (8444, 7149, 7180, 7159, 7142, 7170);
  and ginst2848 (8447, 7142, 4675);
  and ginst2849 (8448, 7149, 7142, 4678);
  and ginst2850 (8449, 7159, 7142, 4682, 7149);
  not ginst2851 (845, 355);
  and ginst2852 (8450, 7170, 7159, 7142, 4687, 7149);
  and ginst2853 (8451, 7149, 4678);
  and ginst2854 (8452, 7159, 4682, 7149);
  and ginst2855 (8453, 7170, 7159, 4687, 7149);
  and ginst2856 (8454, 4682, 7159);
  and ginst2857 (8455, 7170, 7159, 4687);
  and ginst2858 (8456, 7170, 4687);
  not ginst2859 (8457, 7194);
  not ginst2860 (8460, 7198);
  not ginst2861 (8463, 7205);
  not ginst2862 (8466, 7209);
  not ginst2863 (8469, 7216);
  not ginst2864 (8470, 7219);
  not ginst2865 (8471, 7202);
  not ginst2866 (8474, 7202);
  not ginst2867 (8477, 7213);
  not ginst2868 (8480, 7213);
  and ginst2869 (8483, 6083, 6079, 7216);
  and ginst2870 (8484, 7191, 7188, 7219);
  and ginst2871 (8485, 7301, 7240, 7229, 7222);
  and ginst2872 (8488, 7222, 4702);
  and ginst2873 (8489, 7229, 7222, 4706);
  and ginst2874 (8490, 7240, 7222, 4711, 7229);
  and ginst2875 (8491, 7229, 4706);
  and ginst2876 (8492, 7240, 4711, 7229);
  and ginst2877 (8493, 7301, 7240, 7229);
  and ginst2878 (8494, 7229, 4706);
  and ginst2879 (8495, 7240, 4711, 7229);
  and ginst2880 (8496, 7240, 4711);
  and ginst2881 (8497, 7307, 7288, 7272, 7258, 7250);
  and ginst2882 (8500, 7250, 4718);
  and ginst2883 (8501, 7258, 7250, 4722);
  and ginst2884 (8502, 7272, 7250, 4728, 7258);
  and ginst2885 (8503, 7288, 7272, 7250, 4735, 7258);
  and ginst2886 (8504, 7258, 4722);
  and ginst2887 (8505, 7272, 4728, 7258);
  and ginst2888 (8506, 7288, 7272, 4735, 7258);
  and ginst2889 (8507, 7307, 7272, 7258, 7288);
  and ginst2890 (8508, 7258, 4722);
  and ginst2891 (8509, 7272, 4728, 7258);
  and ginst2892 (8510, 7288, 7272, 4735, 7258);
  and ginst2893 (8511, 7272, 4728);
  and ginst2894 (8512, 7288, 7272, 4735);
  and ginst2895 (8513, 7307, 7272, 7288);
  and ginst2896 (8514, 7272, 4728);
  and ginst2897 (8515, 7288, 7272, 4735);
  and ginst2898 (8516, 7288, 4735);
  and ginst2899 (8517, 7301, 7240);
  and ginst2900 (8518, 7307, 7288);
  not ginst2901 (8519, 7314);
  not ginst2902 (8522, 7318);
  not ginst2903 (8525, 7322);
  not ginst2904 (8528, 7322);
  not ginst2905 (853, 358);
  not ginst2906 (8531, 7331);
  not ginst2907 (8534, 7331);
  not ginst2908 (8537, 7340);
  not ginst2909 (8538, 7343);
  and ginst2910 (8539, 6141, 6137, 7340);
  and ginst2911 (8540, 7337, 7334, 7343);
  and ginst2912 (8541, 7376, 7355, 7351, 7346);
  and ginst2913 (8545, 7346, 4757);
  and ginst2914 (8546, 7351, 7346, 4758);
  and ginst2915 (8547, 7355, 7346, 4759, 7351);
  and ginst2916 (8548, 7377, 7373, 7369, 7364, 7358);
  and ginst2917 (8551, 7358, 4762);
  and ginst2918 (8552, 7364, 7358, 4764);
  and ginst2919 (8553, 7369, 7358, 4766, 7364);
  and ginst2920 (8554, 7373, 7369, 7358, 4767, 7364);
  not ginst2921 (8555, 7387);
  not ginst2922 (8558, 7394);
  not ginst2923 (8561, 7398);
  not ginst2924 (8564, 7405);
  not ginst2925 (8565, 7408);
  not ginst2926 (8566, 7391);
  not ginst2927 (8569, 7391);
  not ginst2928 (8572, 7402);
  not ginst2929 (8575, 7402);
  and ginst2930 (8578, 6170, 6166, 7405);
  and ginst2931 (8579, 7381, 7378, 7408);
  not ginst2932 (8580, 7180);
  not ginst2933 (8583, 7142);
  not ginst2934 (8586, 7149);
  not ginst2935 (8589, 7159);
  not ginst2936 (859, 361);
  not ginst2937 (8592, 7170);
  not ginst2938 (8595, 6929);
  not ginst2939 (8598, 6936);
  not ginst2940 (8601, 6946);
  not ginst2941 (8604, 6957);
  not ginst2942 (8607, 7441);
  nand ginst2943 (8608, 7441, 5469);
  not ginst2944 (8609, 7444);
  nand ginst2945 (8610, 7444, 4793);
  not ginst2946 (8615, 7447);
  not ginst2947 (8616, 7450);
  not ginst2948 (8617, 7453);
  not ginst2949 (8618, 7456);
  not ginst2950 (8619, 7474);
  not ginst2951 (8624, 7465);
  not ginst2952 (8625, 7468);
  not ginst2953 (8626, 7471);
  nand ginst2954 (8627, 8144, 8145);
  not ginst2955 (8632, 7479);
  not ginst2956 (8633, 7482);
  not ginst2957 (8634, 7485);
  not ginst2958 (8637, 7491);
  not ginst2959 (8638, 7494);
  not ginst2960 (8639, 7497);
  not ginst2961 (8644, 7503);
  not ginst2962 (8645, 7506);
  not ginst2963 (8646, 7509);
  not ginst2964 (8647, 7512);
  not ginst2965 (8648, 7530);
  not ginst2966 (865, 364);
  not ginst2967 (8653, 7521);
  not ginst2968 (8654, 7524);
  not ginst2969 (8655, 7527);
  not ginst2970 (8660, 6894);
  not ginst2971 (8663, 6894);
  not ginst2972 (8666, 6901);
  not ginst2973 (8669, 6901);
  not ginst2974 (8672, 6912);
  not ginst2975 (8675, 6912);
  not ginst2976 (8678, 7049);
  not ginst2977 (8681, 6988);
  not ginst2978 (8684, 6970);
  not ginst2979 (8687, 6977);
  not ginst2980 (8690, 7049);
  not ginst2981 (8693, 6988);
  not ginst2982 (8696, 6970);
  not ginst2983 (8699, 6977);
  not ginst2984 (8702, 7036);
  not ginst2985 (8705, 6998);
  not ginst2986 (8708, 7020);
  not ginst2987 (871, 367);
  not ginst2988 (8711, 7006);
  not ginst2989 (8714, 7006);
  not ginst2990 (8717, 7553);
  not ginst2991 (8718, 7036);
  not ginst2992 (8721, 6998);
  not ginst2993 (8724, 7020);
  nand ginst2994 (8727, 8216, 8217);
  nand ginst2995 (8730, 8218, 8219);
  not ginst2996 (8733, 7574);
  not ginst2997 (8734, 7577);
  not ginst2998 (8735, 7107);
  not ginst2999 (8738, 7107);
  not ginst3000 (8741, 7114);
  not ginst3001 (8744, 7114);
  not ginst3002 (8747, 7125);
  not ginst3003 (8750, 7125);
  not ginst3004 (8753, 7560);
  not ginst3005 (8754, 7563);
  not ginst3006 (8755, 7566);
  not ginst3007 (8756, 7569);
  not ginst3008 (8757, 7301);
  not ginst3009 (8760, 7240);
  not ginst3010 (8763, 7222);
  not ginst3011 (8766, 7229);
  not ginst3012 (8769, 7301);
  not ginst3013 (8772, 7240);
  not ginst3014 (8775, 7222);
  not ginst3015 (8778, 7229);
  not ginst3016 (8781, 7307);
  not ginst3017 (8784, 7288);
  not ginst3018 (8787, 7250);
  not ginst3019 (8790, 7272);
  not ginst3020 (8793, 7258);
  not ginst3021 (8796, 7258);
  not ginst3022 (8799, 7307);
  not ginst3023 (8802, 7288);
  not ginst3024 (8805, 7250);
  not ginst3025 (8808, 7272);
  nand ginst3026 (881, 467, 585);
  nand ginst3027 (8811, 8232, 8233);
  not ginst3028 (8814, 7588);
  not ginst3029 (8815, 7591);
  not ginst3030 (8816, 7582);
  not ginst3031 (8817, 7585);
  and ginst3032 (8818, 7620, 3155);
  not ginst3033 (882, 528);
  not ginst3034 (883, 578);
  not ginst3035 (884, 575);
  and ginst3036 (8840, 3122, 7609);
  not ginst3037 (885, 494);
  not ginst3038 (8857, 7609);
  and ginst3039 (886, 528, 578);
  and ginst3040 (8861, 6797, 5740, 8274);
  and ginst3041 (8862, 5736, 6800, 8275);
  and ginst3042 (8863, 6803, 5751, 8276);
  and ginst3043 (8864, 5747, 6806, 8277);
  and ginst3044 (8865, 6809, 5762, 8278);
  and ginst3045 (8866, 5758, 6812, 8279);
  and ginst3046 (887, 575, 494);
  not ginst3047 (8871, 7655);
  and ginst3048 (8874, 6833, 7655);
  and ginst3049 (8878, 7671, 6867);
  not ginst3050 (8879, 8196);
  nand ginst3051 (8880, 8196, 8315);
  not ginst3052 (8881, 8200);
  nand ginst3053 (8882, 8200, 8317);
  not ginst3054 (8883, 8204);
  nand ginst3055 (8884, 8204, 8319);
  not ginst3056 (8885, 8208);
  nand ginst3057 (8886, 8208, 8321);
  nand ginst3058 (8887, 3658, 8323);
  nand ginst3059 (8888, 4817, 8325);
  not ginst3060 (889, 590);
  or ginst3061 (8898, 4544, 8337, 8338, 8339);
  or ginst3062 (8902, 4562, 8348, 8349, 8350, 8351);
  or ginst3063 (8920, 4576, 8369, 8370, 8371);
  or ginst3064 (8924, 4581, 8377);
  or ginst3065 (8927, 4592, 8378, 8379, 8380, 8381);
  or ginst3066 (8931, 4603, 8392);
  or ginst3067 (8943, 7825, 8404);
  or ginst3068 (8950, 4630, 8409, 8410, 8411);
  or ginst3069 (8956, 4637, 8415, 8416, 8417, 8418);
  not ginst3070 (8959, 7852);
  and ginst3071 (8960, 3375, 7852);
  or ginst3072 (8963, 4656, 8433, 8434, 8435);
  or ginst3073 (8966, 4674, 8447, 8448, 8449, 8450);
  and ginst3074 (8991, 7188, 6083, 8469);
  and ginst3075 (8992, 6079, 7191, 8470);
  or ginst3076 (8995, 4701, 8488, 8489, 8490);
  or ginst3077 (8996, 4706, 8496);
  or ginst3078 (9001, 4717, 8500, 8501, 8502, 8503);
  or ginst3079 (9005, 4728, 8516);
  and ginst3080 (9024, 7334, 6141, 8537);
  and ginst3081 (9025, 6137, 7337, 8538);
  or ginst3082 (9029, 4756, 8545, 8546, 8547);
  or ginst3083 (9035, 4760, 8551, 8552, 8553, 8554);
  and ginst3084 (9053, 7378, 6170, 8564);
  and ginst3085 (9054, 6166, 7381, 8565);
  nand ginst3086 (9064, 4303, 8607);
  nand ginst3087 (9065, 3507, 8609);
  not ginst3088 (9066, 8114);
  nand ginst3089 (9067, 8114, 4795);
  or ginst3090 (9068, 7613, 6783);
  not ginst3091 (9071, 8117);
  not ginst3092 (9072, 8131);
  nand ginst3093 (9073, 8131, 6195);
  not ginst3094 (9074, 7613);
  not ginst3095 (9077, 8134);
  or ginst3096 (9079, 7650, 6865);
  not ginst3097 (9082, 8146);
  not ginst3098 (9083, 7650);
  not ginst3099 (9086, 8156);
  not ginst3100 (9087, 8166);
  nand ginst3101 (9088, 8166, 4813);
  or ginst3102 (9089, 7659, 6866);
  not ginst3103 (9092, 8169);
  not ginst3104 (9093, 8183);
  nand ginst3105 (9094, 8183, 6203);
  not ginst3106 (9095, 7659);
  not ginst3107 (9098, 8186);
  or ginst3108 (9099, 4545, 8340, 8341, 8342);
  nor ginst3109 (9103, 4545, 8343, 8344);
  or ginst3110 (9107, 4549, 8345, 8346);
  nor ginst3111 (9111, 4549, 8347);
  or ginst3112 (9117, 4577, 8372, 8373, 8374);
  nor ginst3113 (9127, 4577, 8375, 8376);
  nor ginst3114 (9146, 4597, 8390, 8391);
  nor ginst3115 (9149, 4593, 8385, 8386, 8387);
  nand ginst3116 (9159, 7577, 8733);
  nand ginst3117 (9160, 7574, 8734);
  or ginst3118 (9161, 4657, 8436, 8437, 8438);
  nor ginst3119 (9165, 4657, 8439, 8440);
  or ginst3120 (9169, 4661, 8441, 8442);
  nor ginst3121 (9173, 4661, 8443);
  nand ginst3122 (9179, 7563, 8753);
  nand ginst3123 (9180, 7560, 8754);
  nand ginst3124 (9181, 7569, 8755);
  nand ginst3125 (9182, 7566, 8756);
  or ginst3126 (9183, 4702, 8491, 8492, 8493);
  nor ginst3127 (9193, 4702, 8494, 8495);
  or ginst3128 (9203, 4722, 8511, 8512, 8513);
  or ginst3129 (9206, 4718, 8504, 8505, 8506, 8507);
  nor ginst3130 (9220, 4722, 8514, 8515);
  nor ginst3131 (9223, 4718, 8508, 8509, 8510);
  nand ginst3132 (9234, 7591, 8814);
  nand ginst3133 (9235, 7588, 8815);
  nand ginst3134 (9236, 7585, 8816);
  nand ginst3135 (9237, 7582, 8817);
  or ginst3136 (9238, 3159, 8818);
  or ginst3137 (9242, 3126, 8840);
  nand ginst3138 (9243, 8324, 8888);
  not ginst3139 (9244, 8580);
  not ginst3140 (9245, 8583);
  not ginst3141 (9246, 8586);
  not ginst3142 (9247, 8589);
  not ginst3143 (9248, 8592);
  not ginst3144 (9249, 8595);
  not ginst3145 (9250, 8598);
  not ginst3146 (9251, 8601);
  not ginst3147 (9252, 8604);
  nor ginst3148 (9256, 8861, 8280);
  nor ginst3149 (9257, 8862, 8281);
  nor ginst3150 (9258, 8863, 8282);
  nor ginst3151 (9259, 8864, 8283);
  nor ginst3152 (9260, 8865, 8284);
  nor ginst3153 (9261, 8866, 8285);
  not ginst3154 (9262, 8627);
  or ginst3155 (9265, 7649, 8874);
  or ginst3156 (9268, 7668, 8878);
  nand ginst3157 (9271, 7533, 8879);
  nand ginst3158 (9272, 7536, 8881);
  nand ginst3159 (9273, 7539, 8883);
  nand ginst3160 (9274, 7542, 8885);
  nand ginst3161 (9275, 8322, 8887);
  not ginst3162 (9276, 8333);
  and ginst3163 (9280, 6936, 8326, 6946, 6929, 6957);
  and ginst3164 (9285, 367, 8326, 6946, 6957, 6936);
  and ginst3165 (9286, 367, 8326, 6946, 6957);
  and ginst3166 (9287, 367, 8326, 6957);
  and ginst3167 (9288, 367, 8326);
  not ginst3168 (9290, 8660);
  not ginst3169 (9292, 8663);
  not ginst3170 (9294, 8666);
  not ginst3171 (9296, 8669);
  nand ginst3172 (9297, 8672, 5966);
  not ginst3173 (9298, 8672);
  nand ginst3174 (9299, 8675, 6969);
  not ginst3175 (9300, 8675);
  not ginst3176 (9301, 8365);
  and ginst3177 (9307, 8358, 7036, 7020, 7006, 6998);
  and ginst3178 (9314, 8358, 7020, 7006, 7036);
  and ginst3179 (9315, 8358, 7020, 7036);
  and ginst3180 (9318, 8358, 7036);
  not ginst3181 (9319, 8687);
  not ginst3182 (9320, 8699);
  not ginst3183 (9321, 8711);
  not ginst3184 (9322, 8714);
  not ginst3185 (9323, 8727);
  not ginst3186 (9324, 8730);
  not ginst3187 (9326, 8405);
  and ginst3188 (9332, 8405, 8412);
  or ginst3189 (9339, 4193, 8960);
  and ginst3190 (9344, 8430, 8444);
  not ginst3191 (9352, 8735);
  not ginst3192 (9354, 8738);
  not ginst3193 (9356, 8741);
  not ginst3194 (9358, 8744);
  nand ginst3195 (9359, 8747, 6078);
  not ginst3196 (9360, 8747);
  nand ginst3197 (9361, 8750, 7187);
  not ginst3198 (9362, 8750);
  not ginst3199 (9363, 8471);
  not ginst3200 (9364, 8474);
  not ginst3201 (9365, 8477);
  not ginst3202 (9366, 8480);
  nor ginst3203 (9367, 8991, 8483);
  nor ginst3204 (9368, 8992, 8484);
  and ginst3205 (9369, 7198, 7194, 8471);
  and ginst3206 (9370, 8460, 8457, 8474);
  and ginst3207 (9371, 7209, 7205, 8477);
  and ginst3208 (9372, 8466, 8463, 8480);
  not ginst3209 (9375, 8497);
  not ginst3210 (9381, 8766);
  not ginst3211 (9382, 8778);
  not ginst3212 (9383, 8793);
  not ginst3213 (9384, 8796);
  and ginst3214 (9385, 8485, 8497);
  not ginst3215 (9392, 8525);
  not ginst3216 (9393, 8528);
  not ginst3217 (9394, 8531);
  not ginst3218 (9395, 8534);
  and ginst3219 (9396, 7318, 7314, 8525);
  and ginst3220 (9397, 8522, 8519, 8528);
  and ginst3221 (9398, 6131, 6127, 8531);
  and ginst3222 (9399, 7328, 7325, 8534);
  nor ginst3223 (9400, 9024, 8539);
  nor ginst3224 (9401, 9025, 8540);
  not ginst3225 (9402, 8541);
  nand ginst3226 (9407, 8548, 89);
  and ginst3227 (9408, 8541, 8548);
  not ginst3228 (9412, 8811);
  not ginst3229 (9413, 8566);
  not ginst3230 (9414, 8569);
  not ginst3231 (9415, 8572);
  not ginst3232 (9416, 8575);
  nor ginst3233 (9417, 9053, 8578);
  nor ginst3234 (9418, 9054, 8579);
  and ginst3235 (9419, 7387, 6177, 8566);
  and ginst3236 (9420, 8555, 7384, 8569);
  and ginst3237 (9421, 7398, 7394, 8572);
  and ginst3238 (9422, 8561, 8558, 8575);
  not ginst3239 (9423, 8326);
  nand ginst3240 (9426, 9064, 8608);
  nand ginst3241 (9429, 9065, 8610);
  nand ginst3242 (9432, 3515, 9066);
  nand ginst3243 (9435, 4796, 9072);
  nand ginst3244 (9442, 3628, 9087);
  nand ginst3245 (9445, 4814, 9093);
  not ginst3246 (945, 657);
  not ginst3247 (9454, 8678);
  not ginst3248 (9455, 8681);
  not ginst3249 (9456, 8684);
  not ginst3250 (9459, 8690);
  not ginst3251 (9460, 8693);
  not ginst3252 (9461, 8696);
  not ginst3253 (9462, 8358);
  not ginst3254 (9465, 8702);
  not ginst3255 (9466, 8705);
  not ginst3256 (9467, 8708);
  not ginst3257 (9468, 8724);
  not ginst3258 (9473, 8358);
  not ginst3259 (9476, 8718);
  not ginst3260 (9477, 8721);
  nand ginst3261 (9478, 9159, 9160);
  nand ginst3262 (9485, 9179, 9180);
  nand ginst3263 (9488, 9181, 9182);
  not ginst3264 (9493, 8757);
  not ginst3265 (9494, 8760);
  not ginst3266 (9495, 8763);
  not ginst3267 (9498, 8769);
  not ginst3268 (9499, 8772);
  not ginst3269 (9500, 8775);
  not ginst3270 (9505, 8781);
  not ginst3271 (9506, 8784);
  not ginst3272 (9507, 8787);
  not ginst3273 (9508, 8790);
  not ginst3274 (9509, 8808);
  not ginst3275 (9514, 8799);
  not ginst3276 (9515, 8802);
  not ginst3277 (9516, 8805);
  nand ginst3278 (9517, 9234, 9235);
  nand ginst3279 (9520, 9236, 9237);
  and ginst3280 (9526, 8943, 8421);
  and ginst3281 (9531, 8943, 8421);
  nand ginst3282 (9539, 9271, 8880);
  nand ginst3283 (9540, 9273, 8884);
  not ginst3284 (9541, 9275);
  and ginst3285 (9543, 8857, 8254);
  and ginst3286 (9551, 8871, 8288);
  nand ginst3287 (9555, 9272, 8882);
  nand ginst3288 (9556, 9274, 8886);
  not ginst3289 (9557, 8898);
  and ginst3290 (9560, 8902, 8333);
  not ginst3291 (9561, 9099);
  nand ginst3292 (9562, 9099, 9290);
  not ginst3293 (9563, 9103);
  nand ginst3294 (9564, 9103, 9292);
  not ginst3295 (9565, 9107);
  nand ginst3296 (9566, 9107, 9294);
  not ginst3297 (9567, 9111);
  nand ginst3298 (9568, 9111, 9296);
  nand ginst3299 (9569, 4844, 9298);
  not ginst3300 (957, 688);
  nand ginst3301 (9570, 6207, 9300);
  not ginst3302 (9571, 8920);
  not ginst3303 (9575, 8927);
  and ginst3304 (9579, 8365, 8927);
  not ginst3305 (9581, 8950);
  not ginst3306 (9582, 8956);
  and ginst3307 (9585, 8405, 8956);
  and ginst3308 (9591, 8966, 8430);
  not ginst3309 (9592, 9161);
  nand ginst3310 (9593, 9161, 9352);
  not ginst3311 (9594, 9165);
  nand ginst3312 (9595, 9165, 9354);
  not ginst3313 (9596, 9169);
  nand ginst3314 (9597, 9169, 9356);
  not ginst3315 (9598, 9173);
  nand ginst3316 (9599, 9173, 9358);
  nand ginst3317 (9600, 4940, 9360);
  nand ginst3318 (9601, 6220, 9362);
  and ginst3319 (9602, 8457, 7198, 9363);
  and ginst3320 (9603, 7194, 8460, 9364);
  and ginst3321 (9604, 8463, 7209, 9365);
  and ginst3322 (9605, 7205, 8466, 9366);
  not ginst3323 (9608, 9001);
  and ginst3324 (9611, 8485, 9001);
  and ginst3325 (9612, 8519, 7318, 9392);
  and ginst3326 (9613, 7314, 8522, 9393);
  and ginst3327 (9614, 7325, 6131, 9394);
  and ginst3328 (9615, 6127, 7328, 9395);
  not ginst3329 (9616, 9029);
  not ginst3330 (9617, 9035);
  and ginst3331 (9618, 8541, 9035);
  and ginst3332 (9621, 7384, 7387, 9413);
  and ginst3333 (9622, 6177, 8555, 9414);
  and ginst3334 (9623, 8558, 7398, 9415);
  and ginst3335 (9624, 7394, 8561, 9416);
  or ginst3336 (9626, 4563, 8352, 8353, 8354, 9285);
  or ginst3337 (9629, 4566, 8355, 8356, 9286);
  or ginst3338 (9632, 4570, 8357, 9287);
  or ginst3339 (9635, 5960, 9288);
  nand ginst3340 (9642, 9067, 9432);
  not ginst3341 (9645, 9068);
  nand ginst3342 (9646, 9073, 9435);
  not ginst3343 (9649, 9074);
  nand ginst3344 (9650, 9257, 9256);
  nand ginst3345 (9653, 9259, 9258);
  nand ginst3346 (9656, 9261, 9260);
  not ginst3347 (9659, 9079);
  nand ginst3348 (9660, 9079, 4809);
  not ginst3349 (9661, 9083);
  nand ginst3350 (9662, 9083, 6202);
  nand ginst3351 (9663, 9088, 9442);
  not ginst3352 (9666, 9089);
  nand ginst3353 (9667, 9094, 9445);
  not ginst3354 (9670, 9095);
  or ginst3355 (9671, 8924, 8393);
  not ginst3356 (9674, 9117);
  not ginst3357 (9675, 8924);
  not ginst3358 (9678, 9127);
  or ginst3359 (9679, 4597, 8388, 8389, 9315);
  or ginst3360 (9682, 8931, 9318);
  or ginst3361 (9685, 4593, 8382, 8383, 8384, 9314);
  not ginst3362 (9690, 9146);
  nand ginst3363 (9691, 9146, 8717);
  not ginst3364 (9692, 8931);
  not ginst3365 (9695, 9149);
  nand ginst3366 (9698, 9401, 9400);
  nand ginst3367 (9702, 9368, 9367);
  or ginst3368 (9707, 8996, 8517);
  not ginst3369 (9710, 9183);
  not ginst3370 (9711, 8996);
  not ginst3371 (9714, 9193);
  not ginst3372 (9715, 9203);
  nand ginst3373 (9716, 9203, 6235);
  or ginst3374 (9717, 9005, 8518);
  not ginst3375 (9720, 9206);
  not ginst3376 (9721, 9220);
  nand ginst3377 (9722, 9220, 7573);
  not ginst3378 (9723, 9005);
  not ginst3379 (9726, 9223);
  nand ginst3380 (9727, 9418, 9417);
  and ginst3381 (9732, 9268, 8269);
  nand ginst3382 (9733, 9581, 9326);
  and ginst3383 (9734, 89, 9408, 9332, 8394, 8421);
  and ginst3384 (9735, 89, 9408, 9332, 8394, 8421);
  and ginst3385 (9736, 9265, 8262);
  not ginst3386 (9737, 9555);
  not ginst3387 (9738, 9556);
  nand ginst3388 (9739, 9361, 9601);
  nand ginst3389 (9740, 9423, 1115);
  not ginst3390 (9741, 9423);
  nand ginst3391 (9742, 9299, 9570);
  and ginst3392 (9754, 8333, 9280);
  or ginst3393 (9758, 8898, 9560);
  nand ginst3394 (9762, 8660, 9561);
  nand ginst3395 (9763, 8663, 9563);
  nand ginst3396 (9764, 8666, 9565);
  nand ginst3397 (9765, 8669, 9567);
  nand ginst3398 (9766, 9297, 9569);
  and ginst3399 (9767, 9280, 367);
  nand ginst3400 (9768, 9557, 9276);
  not ginst3401 (9769, 9307);
  nand ginst3402 (9773, 9307, 367);
  nand ginst3403 (9774, 9571, 9301);
  and ginst3404 (9775, 8365, 9307);
  or ginst3405 (9779, 8920, 9579);
  not ginst3406 (9784, 9478);
  nand ginst3407 (9785, 9616, 9402);
  or ginst3408 (9786, 8950, 9585);
  and ginst3409 (9790, 89, 9408, 9332, 8394);
  or ginst3410 (9791, 8963, 9591);
  nand ginst3411 (9795, 8735, 9592);
  nand ginst3412 (9796, 8738, 9594);
  nand ginst3413 (9797, 8741, 9596);
  nand ginst3414 (9798, 8744, 9598);
  nand ginst3415 (9799, 9359, 9600);
  nor ginst3416 (9800, 9602, 9369);
  nor ginst3417 (9801, 9603, 9370);
  nor ginst3418 (9802, 9604, 9371);
  nor ginst3419 (9803, 9605, 9372);
  not ginst3420 (9805, 9485);
  not ginst3421 (9806, 9488);
  or ginst3422 (9809, 8995, 9611);
  nor ginst3423 (9813, 9612, 9396);
  nor ginst3424 (9814, 9613, 9397);
  nor ginst3425 (9815, 9614, 9398);
  nor ginst3426 (9816, 9615, 9399);
  and ginst3427 (9817, 9617, 9407);
  or ginst3428 (9820, 9029, 9618);
  not ginst3429 (9825, 9517);
  not ginst3430 (9826, 9520);
  nor ginst3431 (9827, 9621, 9419);
  nor ginst3432 (9828, 9622, 9420);
  nor ginst3433 (9829, 9623, 9421);
  nor ginst3434 (9830, 9624, 9422);
  not ginst3435 (9835, 9426);
  nand ginst3436 (9836, 9426, 4789);
  not ginst3437 (9837, 9429);
  nand ginst3438 (9838, 9429, 4794);
  nand ginst3439 (9846, 3625, 9659);
  nand ginst3440 (9847, 4810, 9661);
  not ginst3441 (9862, 9462);
  nand ginst3442 (9863, 7553, 9690);
  not ginst3443 (9866, 9473);
  nand ginst3444 (9873, 5030, 9715);
  nand ginst3445 (9876, 6236, 9721);
  nand ginst3446 (9890, 9795, 9593);
  nand ginst3447 (9891, 9797, 9597);
  not ginst3448 (9892, 9799);
  nand ginst3449 (9893, 871, 9741);
  nand ginst3450 (9894, 9762, 9562);
  nand ginst3451 (9895, 9764, 9566);
  not ginst3452 (9896, 9766);
  not ginst3453 (9897, 9626);
  nand ginst3454 (9898, 9626, 9249);
  not ginst3455 (9899, 9629);
  nand ginst3456 (9900, 9629, 9250);
  not ginst3457 (9901, 9632);
  nand ginst3458 (9902, 9632, 9251);
  not ginst3459 (9903, 9635);
  nand ginst3460 (9904, 9635, 9252);
  not ginst3461 (9905, 9543);
  not ginst3462 (9906, 9650);
  nand ginst3463 (9907, 9650, 5769);
  not ginst3464 (9908, 9653);
  nand ginst3465 (9909, 9653, 5770);
  not ginst3466 (9910, 9656);
  nand ginst3467 (9911, 9656, 9262);
  not ginst3468 (9917, 9551);
  nand ginst3469 (9923, 9763, 9564);
  nand ginst3470 (9924, 9765, 9568);
  or ginst3471 (9925, 8902, 9767);
  and ginst3472 (9932, 9575, 9773);
  and ginst3473 (9935, 9575, 9769);
  not ginst3474 (9938, 9698);
  nand ginst3475 (9939, 9698, 9323);
  nand ginst3476 (9945, 9796, 9595);
  nand ginst3477 (9946, 9798, 9599);
  not ginst3478 (9947, 9702);
  nand ginst3479 (9948, 9702, 6102);
  and ginst3480 (9949, 9608, 9375);
  not ginst3481 (9953, 9727);
  nand ginst3482 (9954, 9727, 9412);
  nand ginst3483 (9955, 3502, 9835);
  nand ginst3484 (9956, 3510, 9837);
  not ginst3485 (9957, 9642);
  nand ginst3486 (9958, 9642, 9645);
  not ginst3487 (9959, 9646);
  nand ginst3488 (9960, 9646, 9649);
  nand ginst3489 (9961, 9660, 9846);
  nand ginst3490 (9964, 9662, 9847);
  not ginst3491 (9967, 9663);
  nand ginst3492 (9968, 9663, 9666);
  not ginst3493 (9969, 9667);
  nand ginst3494 (9970, 9667, 9670);
  not ginst3495 (9971, 9671);
  nand ginst3496 (9972, 9671, 6213);
  not ginst3497 (9973, 9675);
  nand ginst3498 (9974, 9675, 7551);
  not ginst3499 (9975, 9679);
  nand ginst3500 (9976, 9679, 7552);
  not ginst3501 (9977, 9682);
  not ginst3502 (9978, 9685);
  nand ginst3503 (9979, 9691, 9863);
  not ginst3504 (9982, 9692);
  nand ginst3505 (9983, 9814, 9813);
  nand ginst3506 (9986, 9816, 9815);
  nand ginst3507 (9989, 9801, 9800);
  nand ginst3508 (9992, 9803, 9802);
  not ginst3509 (9995, 9707);
  nand ginst3510 (9996, 9707, 6231);
  not ginst3511 (9997, 9711);
  nand ginst3512 (9998, 9711, 7572);
  nand ginst3513 (9999, 9716, 9873);

  SatHard block1 (flip_signal, 3390, 4538, 1863, 5944, 6540, 2315, 1395, 6067, keyinput0, keyinput1, keyinput2, keyinput3, keyinput4, keyinput5, keyinput6, keyinput7, keyinput8, keyinput9, keyinput10, keyinput11, keyinput12, keyinput13, keyinput14, keyinput15);

endmodule

/*************** SatHard block ***************/
module SatHard (flip_signal, 3390, 4538, 1863, 5944, 6540, 2315, 1395, 6067, keyinput0, keyinput1, keyinput2, keyinput3, keyinput4, keyinput5, keyinput6, keyinput7, keyinput8, keyinput9, keyinput10, keyinput11, keyinput12, keyinput13, keyinput14, keyinput15);

  input 3390, 4538, 1863, 5944, 6540, 2315, 1395, 6067;
  input keyinput0, keyinput1, keyinput2, keyinput3, keyinput4, keyinput5, keyinput6, keyinput7, keyinput8, keyinput9, keyinput10, keyinput11, keyinput12, keyinput13, keyinput14, keyinput15;
  output flip_signal;
  wire newWire0, newWire1, newWire2, newWire3, newWire4, newWire5, newWire6, newWire7, newWire8, newWire9, newWire10, newWire11, newWire12, newWire13, newWire14, newWire15, newWire16, newWire17;

  //SatHard key=0010100101011010
  wire [7:0] sat_res_inputs;
  assign sat_res_inputs[7:0] = {3390, 4538, 1863, 5944, 6540, 2315, 1395, 6067};
  wire [15:0] keyinputs, keyvalue;
  assign keyinputs[15:0] = {keyinput0, keyinput1, keyinput2, keyinput3, keyinput4, keyinput5, keyinput6, keyinput7, keyinput8, keyinput9, keyinput10, keyinput11, keyinput12, keyinput13, keyinput14, keyinput15};
  assign keyvalue[15:0] = 16'b0010100101011010;

  assign flip_signal = ( (keyinputs!=keyvalue) & (sat_res_inputs[7:0]==~keyinputs[7:0]) & (sat_res_inputs[7:0]==keyinputs[15:8]) ) ? 'b1 : 'b0;

endmodule
/*************** SatHard block ***************/
