//key=0100000100110000111101110000000101100111101101101001111010100001
// Main module
module c3540_SFLL-HD(2)_64(1, 13, 20, 33, 41, 45, 50, 58, 68, 77, 87, 97, 107, 116, 124, 125, 128, 132, 137, 143, 150, 159, 169, 179, 190, 200, 213, 222, 223, 226, 232, 238, 244, 250, 257, 264, 270, 274, 283, 294, 303, 311, 317, 322, 326, 329, 330, 343, 349, 350, keyinput0, keyinput1, keyinput2, keyinput3, keyinput4, keyinput5, keyinput6, keyinput7, keyinput8, keyinput9, keyinput10, keyinput11, keyinput12, keyinput13, keyinput14, keyinput15, keyinput16, keyinput17, keyinput18, keyinput19, keyinput20, keyinput21, keyinput22, keyinput23, keyinput24, keyinput25, keyinput26, keyinput27, keyinput28, keyinput29, keyinput30, keyinput31, keyinput32, keyinput33, keyinput34, keyinput35, keyinput36, keyinput37, keyinput38, keyinput39, keyinput40, keyinput41, keyinput42, keyinput43, keyinput44, keyinput45, keyinput46, keyinput47, keyinput48, keyinput49, keyinput50, keyinput51, keyinput52, keyinput53, keyinput54, keyinput55, keyinput56, keyinput57, keyinput58, keyinput59, keyinput60, keyinput61, keyinput62, keyinput63, 1713, 1947, 3195, 3833, 3987, 4028, 4145, 4589, 4667, 4815, 4944, 5002, 5045, 5047, 5078, 5102, 5120, 5121, 5192, 5231, 5360, 5361);

  input 1, 13, 20, 33, 41, 45, 50, 58, 68, 77, 87, 97, 107, 116, 124, 125, 128, 132, 137, 143, 150, 159, 169, 179, 190, 200, 213, 222, 223, 226, 232, 238, 244, 250, 257, 264, 270, 274, 283, 294, 303, 311, 317, 322, 326, 329, 330, 343, 349, 350, keyinput0, keyinput1, keyinput2, keyinput3, keyinput4, keyinput5, keyinput6, keyinput7, keyinput8, keyinput9, keyinput10, keyinput11, keyinput12, keyinput13, keyinput14, keyinput15, keyinput16, keyinput17, keyinput18, keyinput19, keyinput20, keyinput21, keyinput22, keyinput23, keyinput24, keyinput25, keyinput26, keyinput27, keyinput28, keyinput29, keyinput30, keyinput31, keyinput32, keyinput33, keyinput34, keyinput35, keyinput36, keyinput37, keyinput38, keyinput39, keyinput40, keyinput41, keyinput42, keyinput43, keyinput44, keyinput45, keyinput46, keyinput47, keyinput48, keyinput49, keyinput50, keyinput51, keyinput52, keyinput53, keyinput54, keyinput55, keyinput56, keyinput57, keyinput58, keyinput59, keyinput60, keyinput61, keyinput62, keyinput63;
  output 1713, 1947, 3195, 3833, 3987, 4028, 4145, 4589, 4667, 4815, 4944, 5002, 5045, 5047, 5078, 5102, 5120, 5121, 5192, 5231, 5360, 5361;
  wire 1067, 1117, 1179, 1196, 1197, 1202, 1219, 1250, 1251, 1252, 1253, 1254, 1255, 1256, 1257, 1258, 1259, 1260, 1261, 1262, 1263, 1264, 1267, 1268, 1271, 1272, 1273, 1276, 1279, 1298, 1302, 1306, 1315, 1322, 1325, 1328, 1331, 1334, 1337, 1338, 1339, 1340, 1343, 1344, 1345, 1346, 1347, 1348, 1349, 1350, 1351, 1352, 1353, 1358, 1363, 1366, 1369, 1384, 1401, 1402, 1403, 1404, 1405, 1406, 1407, 1408, 1409, 1426, 1427, 1452, 1459, 1460, 1461, 1464, 1467, 1468, 1469, 1470, 1471, 1474, 1475, 1478, 1481, 1484, 1487, 1490, 1493, 1496, 1499, 1502, 1505, 1507, 1508, 1509, 1510, 1511, 1512, 1520, 1562, 1579, 1580, 1581, 1582, 1583, 1584, 1585, 1586, 1587, 1588, 1589, 1590, 1591, 1592, 1593, 1594, 1595, 1596, 1597, 1598, 1599, 1600, 1643, 1644, 1645, 1646, 1647, 1648, 1649, 1650, 1667, 1670, 1673, 1674, 1675, 1676, 1677, 1678, 1679, 1680, 1691, 1692, 1693, 1694, 1714, 1715, 1718, 1721, 1722, 1725, 1726, 1727, 1728, 1729, 1730, 1731, 1735, 1736, 1737, 1738, 1747, 1756, 1761, 1764, 1765, 1766, 1767, 1768, 1769, 1770, 1787, 1788, 1789, 1790, 1791, 1792, 1793, 1794, 1795, 1796, 1797, 1798, 1799, 1800, 1801, 1802, 1803, 1806, 1809, 1812, 1815, 1818, 1821, 1824, 1833, 1842, 1843, 1844, 1845, 1846, 1847, 1848, 1849, 1850, 1851, 1852, 1853, 1854, 1855, 1856, 1857, 1858, 1859, 1860, 1861, 1862, 1863, 1864, 1869, 1870, 1873, 1874, 1875, 1878, 1879, 1880, 1883, 1884, 1885, 1888, 1889, 1890, 1893, 1894, 1895, 1898, 1899, 1900, 1903, 1904, 1905, 1908, 1909, 1912, 1913, 1917, 1922, 1926, 1930, 1933, 1936, 1939, 1940, 1941, 1942, 1943, 1944, 1945, 1946, 1960, 1961, 1966, 1981, 1982, 1983, 1986, 1987, 1988, 1989, 1990, 1991, 2022, 2023, 2024, 2025, 2026, 2027, 2028, 2029, 2030, 2031, 2032, 2033, 2034, 2035, 2036, 2037, 2038, 2043, 2052, 2057, 2068, 2073, 2078, 2083, 2088, 2093, 2098, 2103, 2121, 2122, 2123, 2124, 2125, 2126, 2127, 2128, 2133, 2134, 2135, 2136, 2137, 2138, 2139, 2141, 2142, 2143, 2144, 2145, 2146, 2147, 2148, 2149, 2150, 2151, 2152, 2153, 2154, 2155, 2156, 2157, 2158, 2175, 2178, 2179, 2180, 2181, 2183, 2184, 2185, 2188, 2191, 2194, 2197, 2200, 2203, 2206, 2209, 2210, 2211, 2212, 2221, 2230, 2231, 2232, 2233, 2234, 2235, 2236, 2237, 2238, 2239, 2240, 2241, 2242, 2243, 2244, 2245, 2270, 2277, 2282, 2287, 2294, 2299, 2304, 2307, 2310, 2313, 2316, 2319, 2322, 2325, 2328, 2331, 2334, 2341, 2342, 2347, 2348, 2349, 2350, 2351, 2352, 2353, 2354, 2355, 2374, 2375, 2376, 2379, 2398, 2417, 2418, 2419, 2420, 2421, 2422, 2425, 2426, 2427, 2430, 2431, 2432, 2435, 2436, 2437, 2438, 2439, 2440, 2443, 2444, 2445, 2448, 2449, 2450, 2467, 2468, 2469, 2470, 2471, 2474, 2475, 2476, 2477, 2478, 2481, 2482, 2483, 2486, 2487, 2488, 2497, 2506, 2515, 2524, 2533, 2542, 2551, 2560, 2569, 2578, 2587, 2596, 2605, 2614, 2623, 2632, 2633, 2634, 2635, 2636, 2637, 2638, 2639, 2640, 2641, 2642, 2643, 2644, 2645, 2646, 2647, 2648, 2652, 2656, 2659, 2662, 2666, 2670, 2673, 2677, 2681, 2684, 2688, 2692, 2697, 2702, 2706, 2710, 2715, 2719, 2723, 2728, 2729, 2730, 2731, 2732, 2733, 2734, 2735, 2736, 2737, 2738, 2739, 2740, 2741, 2742, 2743, 2744, 2745, 2746, 2748, 2749, 2750, 2751, 2754, 2755, 2756, 2757, 2758, 2761, 2764, 2768, 2769, 2898, 2899, 2900, 2901, 2962, 2966, 2967, 2970, 2973, 2977, 2980, 2984, 2985, 2986, 2987, 2988, 2989, 2990, 2991, 2992, 2993, 2994, 2995, 2996, 2997, 2998, 2999, 3000, 3001, 3002, 3003, 3004, 3005, 3006, 3007, 3008, 3009, 3010, 3011, 3012, 3013, 3014, 3015, 3016, 3017, 3018, 3019, 3020, 3021, 3022, 3023, 3024, 3025, 3026, 3027, 3028, 3029, 3030, 3031, 3032, 3033, 3034, 3035, 3036, 3037, 3038, 3039, 3040, 3041, 3042, 3043, 3044, 3045, 3046, 3047, 3048, 3049, 3050, 3051, 3052, 3053, 3054, 3055, 3056, 3057, 3058, 3059, 3060, 3061, 3062, 3063, 3064, 3065, 3066, 3067, 3068, 3069, 3070, 3071, 3072, 3073, 3074, 3075, 3076, 3077, 3078, 3079, 3080, 3081, 3082, 3083, 3084, 3085, 3086, 3087, 3088, 3089, 3090, 3091, 3092, 3093, 3094, 3095, 3096, 3097, 3098, 3099, 3100, 3101, 3102, 3103, 3104, 3105, 3106, 3107, 3108, 3109, 3110, 3111, 3112, 3115, 3118, 3119, 3122, 3125, 3128, 3131, 3134, 3135, 3138, 3141, 3142, 3145, 3148, 3149, 3152, 3155, 3158, 3161, 3164, 3165, 3168, 3171, 3172, 3175, 3178, 3181, 3184, 3187, 3190, 3191, 3192, 3193, 3194, 3196, 3206, 3207, 3208, 3209, 3210, 3211, 3212, 3213, 3214, 3215, 3216, 3217, 3218, 3219, 3220, 3221, 3222, 3223, 3224, 3225, 3226, 3227, 3228, 3229, 3230, 3231, 3232, 3233, 3234, 3235, 3236, 3237, 3238, 3239, 3240, 3241, 3242, 3243, 3244, 3245, 3246, 3247, 3248, 3249, 3250, 3251, 3252, 3253, 3254, 3255, 3256, 3257, 3258, 3259, 3260, 3261, 3262, 3263, 3264, 3265, 3266, 3267, 3268, 3269, 3270, 3271, 3272, 3273, 3274, 3275, 3276, 3277, 3278, 3279, 3280, 3281, 3282, 3283, 3284, 3285, 3286, 3287, 3288, 3289, 3290, 3291, 3292, 3293, 3294, 3295, 3296, 3297, 3298, 3299, 3300, 3301, 3302, 3303, 3304, 3305, 3306, 3307, 3308, 3309, 3310, 3311, 3312, 3313, 3314, 3315, 3316, 3317, 3318, 3319, 3320, 3321, 3322, 3323, 3324, 3325, 3326, 3327, 3328, 3329, 3330, 3331, 3332, 3333, 3334, 3383, 3384, 3387, 3388, 3389, 3390, 3391, 3392, 3393, 3394, 3395, 3396, 3397, 3398, 3399, 3400, 3401, 3402, 3403, 3404, 3405, 3406, 3407, 3410, 3413, 3414, 3415, 3419, 3423, 3426, 3429, 3430, 3431, 3434, 3437, 3438, 3439, 3442, 3445, 3446, 3447, 3451, 3455, 3458, 3461, 3462, 3463, 3466, 3469, 3470, 3471, 3472, 3475, 3478, 3481, 3484, 3487, 3490, 3493, 3496, 3499, 3502, 3505, 3508, 3511, 3514, 3517, 3520, 3523, 3534, 3535, 3536, 3537, 3538, 3539, 3540, 3541, 3542, 3543, 3544, 3545, 3546, 3547, 3548, 3549, 3550, 3551, 3552, 3557, 3568, 3573, 3578, 3589, 3594, 3605, 3626, 3627, 3628, 3629, 3630, 3631, 3632, 3633, 3634, 3635, 3636, 3637, 3638, 3639, 3640, 3641, 3642, 3643, 3644, 3645, 3648, 3651, 3652, 3653, 3654, 3657, 3658, 3661, 3662, 3663, 3664, 3667, 3670, 3671, 3672, 3673, 3676, 3677, 3680, 3681, 3682, 3685, 3686, 3687, 3688, 3689, 3690, 3693, 3694, 3695, 3696, 3697, 3700, 3703, 3704, 3705, 3706, 3707, 3708, 3711, 3712, 3713, 3714, 3715, 3716, 3717, 3718, 3719, 3720, 3721, 3731, 3734, 3740, 3743, 3753, 3756, 3762, 3765, 3766, 3773, 3774, 3775, 3776, 3777, 3778, 3779, 3780, 3786, 3789, 3800, 3803, 3809, 3812, 3815, 3818, 3821, 3824, 3827, 3830, 3834, 3835, 3838, 3845, 3850, 3855, 3858, 3861, 3865, 3868, 3884, 3885, 3894, 3895, 3898, 3899, 3906, 3911, 3912, 3913, 3916, 3917, 3920, 3921, 3924, 3925, 3926, 3930, 3931, 3932, 3935, 3936, 3937, 3940, 3947, 3948, 3950, 3953, 3956, 3959, 3962, 3965, 3968, 3971, 3974, 3977, 3980, 3983, 3992, 3996, 4013, 4029, 4030, 4031, 4032, 4033, 4034, 4035, 4042, 4043, 4044, 4045, 4046, 4047, 4048, 4049, 4050, 4051, 4052, 4053, 4054, 4055, 4056, 4057, 4058, 4059, 4062, 4065, 4066, 4067, 4070, 4073, 4074, 4075, 4076, 4077, 4078, 4079, 4080, 4085, 4086, 4088, 4090, 4091, 4094, 4098, 4101, 4104, 4105, 4106, 4107, 4108, 4109, 4110, 4111, 4112, 4113, 4114, 4115, 4116, 4119, 4122, 4123, 4126, 4127, 4128, 4139, 4142, 4146, 4147, 4148, 4149, 4150, 4151, 4152, 4153, 4154, 4161, 4167, 4174, 4182, 4186, 4189, 4190, 4191, 4192, 4193, 4194, 4195, 4196, 4197, 4200, 4203, 4209, 4213, 4218, 4223, 4238, 4239, 4241, 4242, 4247, 4251, 4252, 4253, 4254, 4255, 4256, 4257, 4258, 4283, 4284, 4287, 4291, 4295, 4296, 4299, 4303, 4304, 4305, 4310, 4316, 4317, 4318, 4319, 4322, 4325, 4326, 4327, 4328, 4329, 4330, 4331, 4335, 4338, 4341, 4344, 4347, 4350, 4353, 4356, 4359, 4362, 4365, 4368, 4371, 4376, 4377, 4387, 4390, 4393, 4398, 4413, 4416, 4421, 4427, 4430, 4435, 4442, 4443, 4446, 4447, 4448, 4452, 4458, 4461, 4462, 4463, 4464, 4465, 4468, 4472, 4475, 4479, 4484, 4486, 4487, 4491, 4493, 4496, 4497, 4498, 4503, 4506, 4507, 4508, 4509, 4510, 4511, 4515, 4526, 4527, 4528, 4529, 4530, 4531, 4534, 4537, 4540, 4545, 4549, 4552, 4555, 4558, 4559, 4562, 4563, 4564, 4568, 4569, 4572, 4573, 4576, 4581, 4584, 4587, 4588, 4593, 4596, 4597, 4599, 4602, 4603, 4608, 4613, 4616, 4619, 4623, 4628, 4629, 4630, 4635, 4636, 4640, 4641, 4642, 4643, 4644, 4647, 4650, 4656, 4659, 4664, 4668, 4669, 4670, 4673, 4674, 4675, 4676, 4677, 4678, 4679, 4687, 4688, 4691, 4694, 4697, 4700, 4704, 4705, 4706, 4707, 4708, 4711, 4716, 4717, 4721, 4722, 4726, 4727, 4730, 4733, 4740, 4743, 4747, 4748, 4749, 4750, 4753, 4754, 4755, 4756, 4757, 4769, 4772, 4775, 4778, 4786, 4787, 4788, 4789, 4794, 4797, 4800, 4805, 4808, 4812, 4816, 4817, 4818, 4822, 4823, 4826, 4829, 4830, 4831, 4838, 4844, 4847, 4850, 4854, 4859, 4860, 4868, 4870, 4872, 4873, 4876, 4880, 4885, 4889, 4895, 4896, 4897, 4898, 4899, 4900, 4901, 4902, 4904, 4905, 4906, 4907, 4913, 4916, 4920, 4921, 4924, 4925, 4926, 4928, 4929, 4930, 4931, 4937, 4940, 4946, 4949, 4950, 4951, 4952, 4953, 4954, 4957, 4964, 4965, 4968, 4969, 4970, 4973, 4978, 4979, 4980, 4981, 4982, 4983, 4984, 4985, 4988, 4991, 4996, 4999, 5007, 5010, 5013, 5018, 5021, 5026, 5029, 5030, 5039, 5042, 5046, 5050, 5055, 5058, 5061, 5066, 5070, 5080, 5085, 5094, 5095, 5097, 5103, 5108, 5109, 5110, 5111, 5114, 5117, 5122, 5125, 5128, 5133, 5136, 5139, 5145, 5151, 5154, 5159, 5160, 5163, 5166, 5173, 5174, 5177, 5182, 5183, 5184, 5188, 5193, 5196, 5197, 5198, 5199, 5201, 5203, 5205, 5209, 5212, 5215, 5217, 5219, 5220, 5221, 5222, 5223, 5224, 5225, 5228, 5232, 5233, 5234, 5235, 5236, 5240, 5242, 5243, 5245, 5246, 5250, 5253, 5254, 5257, 5258, 5261, 5266, 5269, 5277, 5278, 5279, 5283, 5284, 5285, 5286, 5289, 5292, 5295, 5298, 5303, 5306, 5309, 5312, 5313, 5322, 5323, 5324, 5327, 5332, 5335, 5340, 5341, 5344, 5345, 5348, 5349, 5350, 5351, 5352, 5353, 5354, 5355, 5356, 5357, 5358, 5359, 655, 665, 670, 679, 683, 686, 690, 699, 702, 706, 715, 724, 727, 736, 740, 749, 753, 763, 768, 769, 772, 779, 782, 786, 793, 794, 798, 803, 820, 821, 825, 829, 832, 835, 836, 839, 842, 845, 848, 851, 854, 858, 861, 864, 867, 870, 874, 877, 880, 883, 886, 889, 890, 891, 892, 895, 896, 913, 914, 915, 916, 917, 920, 923, 926, 929, 932, 935, 938, 941, 944, 947, 950, 953, 956, 959, 962, 965, 5102_in, flip_signal;

  and ginst1 (1067, 250, 768);
  or ginst2 (1117, 820, 20);
  or ginst3 (1179, 895, 169);
  not ginst4 (1196, 793);
  or ginst5 (1197, 915, 1);
  and ginst6 (1202, 913, 914);
  or ginst7 (1219, 916, 1);
  and ginst8 (1250, 842, 848, 854);
  nand ginst9 (1251, 226, 655);
  nand ginst10 (1252, 232, 670);
  nand ginst11 (1253, 238, 690);
  nand ginst12 (1254, 244, 706);
  nand ginst13 (1255, 250, 715);
  nand ginst14 (1256, 257, 727);
  nand ginst15 (1257, 264, 740);
  nand ginst16 (1258, 270, 753);
  not ginst17 (1259, 926);
  not ginst18 (1260, 929);
  not ginst19 (1261, 932);
  not ginst20 (1262, 935);
  nand ginst21 (1263, 679, 686);
  nand ginst22 (1264, 736, 749);
  nand ginst23 (1267, 683, 699);
  not ginst24 (1268, 665);
  not ginst25 (1271, 953);
  not ginst26 (1272, 959);
  not ginst27 (1273, 839);
  not ginst28 (1276, 839);
  not ginst29 (1279, 782);
  not ginst30 (1298, 825);
  not ginst31 (1302, 832);
  and ginst32 (1306, 779, 835);
  and ginst33 (1315, 779, 836, 832);
  and ginst34 (1322, 769, 836);
  and ginst35 (1325, 772, 786, 798);
  nand ginst36 (1328, 772, 786, 798);
  nand ginst37 (1331, 772, 786);
  not ginst38 (1334, 874);
  nand ginst39 (1337, 782, 794, 45);
  nand ginst40 (1338, 842, 848, 854);
  not ginst41 (1339, 956);
  and ginst42 (1340, 861, 867, 870);
  nand ginst43 (1343, 861, 867, 870);
  not ginst44 (1344, 962);
  not ginst45 (1345, 803);
  not ginst46 (1346, 803);
  not ginst47 (1347, 803);
  not ginst48 (1348, 803);
  not ginst49 (1349, 803);
  not ginst50 (1350, 803);
  not ginst51 (1351, 803);
  not ginst52 (1352, 803);
  or ginst53 (1353, 883, 886);
  nor ginst54 (1358, 883, 886);
  not ginst55 (1363, 892);
  not ginst56 (1366, 892);
  not ginst57 (1369, 821);
  not ginst58 (1384, 825);
  not ginst59 (1401, 896);
  not ginst60 (1402, 896);
  not ginst61 (1403, 896);
  not ginst62 (1404, 896);
  not ginst63 (1405, 896);
  not ginst64 (1406, 896);
  not ginst65 (1407, 896);
  not ginst66 (1408, 896);
  or ginst67 (1409, 1, 1196);
  not ginst68 (1426, 829);
  not ginst69 (1427, 829);
  and ginst70 (1452, 769, 782, 794);
  not ginst71 (1459, 917);
  not ginst72 (1460, 965);
  or ginst73 (1461, 920, 923);
  nor ginst74 (1464, 920, 923);
  not ginst75 (1467, 938);
  not ginst76 (1468, 941);
  not ginst77 (1469, 944);
  not ginst78 (1470, 947);
  not ginst79 (1471, 679);
  not ginst80 (1474, 950);
  not ginst81 (1475, 686);
  not ginst82 (1478, 702);
  not ginst83 (1481, 724);
  not ginst84 (1484, 736);
  not ginst85 (1487, 749);
  not ginst86 (1490, 763);
  not ginst87 (1493, 877);
  not ginst88 (1496, 877);
  not ginst89 (1499, 880);
  not ginst90 (1502, 880);
  nand ginst91 (1505, 702, 1250);
  and ginst92 (1507, 1251, 1252, 1253, 1254);
  and ginst93 (1508, 1255, 1256, 1257, 1258);
  nand ginst94 (1509, 929, 1259);
  nand ginst95 (1510, 926, 1260);
  nand ginst96 (1511, 935, 1261);
  nand ginst97 (1512, 932, 1262);
  and ginst98 (1520, 655, 1263);
  and ginst99 (1562, 874, 1337);
  not ginst100 (1579, 1117);
  and ginst101 (1580, 803, 1117);
  and ginst102 (1581, 1338, 1345);
  not ginst103 (1582, 1117);
  and ginst104 (1583, 803, 1117);
  not ginst105 (1584, 1117);
  and ginst106 (1585, 803, 1117);
  and ginst107 (1586, 854, 1347);
  not ginst108 (1587, 1117);
  and ginst109 (1588, 803, 1117);
  and ginst110 (1589, 77, 1348);
  not ginst111 (1590, 1117);
  and ginst112 (1591, 803, 1117);
  and ginst113 (1592, 1343, 1349);
  not ginst114 (1593, 1117);
  and ginst115 (1594, 803, 1117);
  not ginst116 (1595, 1117);
  and ginst117 (1596, 803, 1117);
  and ginst118 (1597, 870, 1351);
  not ginst119 (1598, 1117);
  and ginst120 (1599, 803, 1117);
  and ginst121 (1600, 116, 1352);
  and ginst122 (1643, 222, 1401);
  and ginst123 (1644, 223, 1402);
  and ginst124 (1645, 226, 1403);
  and ginst125 (1646, 232, 1404);
  and ginst126 (1647, 238, 1405);
  and ginst127 (1648, 244, 1406);
  and ginst128 (1649, 250, 1407);
  and ginst129 (1650, 257, 1408);
  and ginst130 (1667, 1, 13, 1426);
  and ginst131 (1670, 1, 13, 1427);
  not ginst132 (1673, 1202);
  not ginst133 (1674, 1202);
  not ginst134 (1675, 1202);
  not ginst135 (1676, 1202);
  not ginst136 (1677, 1202);
  not ginst137 (1678, 1202);
  not ginst138 (1679, 1202);
  not ginst139 (1680, 1202);
  nand ginst140 (1691, 941, 1467);
  nand ginst141 (1692, 938, 1468);
  nand ginst142 (1693, 947, 1469);
  nand ginst143 (1694, 944, 1470);
  not ginst144 (1713, 1505);
  and ginst145 (1714, 87, 1264);
  nand ginst146 (1715, 1509, 1510);
  nand ginst147 (1718, 1511, 1512);
  nand ginst148 (1721, 1507, 1508);
  and ginst149 (1722, 763, 1340);
  nand ginst150 (1725, 763, 1340);
  not ginst151 (1726, 1268);
  nand ginst152 (1727, 1493, 1271);
  not ginst153 (1728, 1493);
  and ginst154 (1729, 683, 1268);
  nand ginst155 (1730, 1499, 1272);
  not ginst156 (1731, 1499);
  nand ginst157 (1735, 87, 1264);
  not ginst158 (1736, 1273);
  not ginst159 (1737, 1276);
  nand ginst160 (1738, 1325, 821);
  nand ginst161 (1747, 1325, 825);
  nand ginst162 (1756, 772, 1279, 798);
  nand ginst163 (1761, 772, 786, 798, 1302);
  nand ginst164 (1764, 1496, 1339);
  not ginst165 (1765, 1496);
  nand ginst166 (1766, 1502, 1344);
  not ginst167 (1767, 1502);
  not ginst168 (1768, 1328);
  not ginst169 (1769, 1334);
  not ginst170 (1770, 1331);
  and ginst171 (1787, 845, 1579);
  and ginst172 (1788, 150, 1580);
  and ginst173 (1789, 851, 1582);
  and ginst174 (1790, 159, 1583);
  and ginst175 (1791, 77, 1584);
  and ginst176 (1792, 50, 1585);
  and ginst177 (1793, 858, 1587);
  and ginst178 (1794, 845, 1588);
  and ginst179 (1795, 864, 1590);
  and ginst180 (1796, 851, 1591);
  and ginst181 (1797, 107, 1593);
  and ginst182 (1798, 77, 1594);
  and ginst183 (1799, 116, 1595);
  and ginst184 (1800, 858, 1596);
  and ginst185 (1801, 283, 1598);
  and ginst186 (1802, 864, 1599);
  and ginst187 (1803, 200, 1363);
  and ginst188 (1806, 889, 1363);
  and ginst189 (1809, 890, 1366);
  and ginst190 (1812, 891, 1366);
  nand ginst191 (1815, 1298, 1302);
  nand ginst192 (1818, 821, 1302);
  nand ginst193 (1821, 772, 1279, 1179);
  nand ginst194 (1824, 786, 794, 1298);
  nand ginst195 (1833, 786, 1298);
  not ginst196 (1842, 1369);
  not ginst197 (1843, 1369);
  not ginst198 (1844, 1369);
  not ginst199 (1845, 1369);
  not ginst200 (1846, 1369);
  not ginst201 (1847, 1369);
  not ginst202 (1848, 1369);
  not ginst203 (1849, 1384);
  and ginst204 (1850, 1384, 896);
  not ginst205 (1851, 1384);
  and ginst206 (1852, 1384, 896);
  not ginst207 (1853, 1384);
  and ginst208 (1854, 1384, 896);
  not ginst209 (1855, 1384);
  and ginst210 (1856, 1384, 896);
  not ginst211 (1857, 1384);
  and ginst212 (1858, 1384, 896);
  not ginst213 (1859, 1384);
  and ginst214 (1860, 1384, 896);
  not ginst215 (1861, 1384);
  and ginst216 (1862, 1384, 896);
  not ginst217 (1863, 1384);
  and ginst218 (1864, 1384, 896);
  and ginst219 (1869, 1202, 1409);
  nor ginst220 (1870, 50, 1409);
  not ginst221 (1873, 1306);
  and ginst222 (1874, 1202, 1409);
  nor ginst223 (1875, 58, 1409);
  not ginst224 (1878, 1306);
  and ginst225 (1879, 1202, 1409);
  nor ginst226 (1880, 68, 1409);
  not ginst227 (1883, 1306);
  and ginst228 (1884, 1202, 1409);
  nor ginst229 (1885, 77, 1409);
  not ginst230 (1888, 1306);
  and ginst231 (1889, 1202, 1409);
  nor ginst232 (1890, 87, 1409);
  not ginst233 (1893, 1322);
  and ginst234 (1894, 1202, 1409);
  nor ginst235 (1895, 97, 1409);
  not ginst236 (1898, 1315);
  and ginst237 (1899, 1202, 1409);
  nor ginst238 (1900, 107, 1409);
  not ginst239 (1903, 1315);
  and ginst240 (1904, 1202, 1409);
  nor ginst241 (1905, 116, 1409);
  not ginst242 (1908, 1315);
  and ginst243 (1909, 1452, 213);
  nand ginst244 (1912, 1452, 213);
  and ginst245 (1913, 1452, 213, 343);
  nand ginst246 (1917, 1452, 213, 343);
  and ginst247 (1922, 1452, 213, 343);
  nand ginst248 (1926, 1452, 213, 343);
  not ginst249 (1930, 1464);
  nand ginst250 (1933, 1691, 1692);
  nand ginst251 (1936, 1693, 1694);
  not ginst252 (1939, 1471);
  nand ginst253 (1940, 1471, 1474);
  not ginst254 (1941, 1475);
  not ginst255 (1942, 1478);
  not ginst256 (1943, 1481);
  not ginst257 (1944, 1484);
  not ginst258 (1945, 1487);
  not ginst259 (1946, 1490);
  not ginst260 (1947, 1714);
  nand ginst261 (1960, 953, 1728);
  nand ginst262 (1961, 959, 1731);
  and ginst263 (1966, 1520, 1276);
  nand ginst264 (1981, 956, 1765);
  nand ginst265 (1982, 962, 1767);
  and ginst266 (1983, 1067, 1768);
  or ginst267 (1986, 1581, 1787, 1788);
  or ginst268 (1987, 1586, 1791, 1792);
  or ginst269 (1988, 1589, 1793, 1794);
  or ginst270 (1989, 1592, 1795, 1796);
  or ginst271 (1990, 1597, 1799, 1800);
  or ginst272 (1991, 1600, 1801, 1802);
  and ginst273 (2022, 77, 1849);
  and ginst274 (2023, 223, 1850);
  and ginst275 (2024, 87, 1851);
  and ginst276 (2025, 226, 1852);
  and ginst277 (2026, 97, 1853);
  and ginst278 (2027, 232, 1854);
  and ginst279 (2028, 107, 1855);
  and ginst280 (2029, 238, 1856);
  and ginst281 (2030, 116, 1857);
  and ginst282 (2031, 244, 1858);
  and ginst283 (2032, 283, 1859);
  and ginst284 (2033, 250, 1860);
  and ginst285 (2034, 294, 1861);
  and ginst286 (2035, 257, 1862);
  and ginst287 (2036, 303, 1863);
  and ginst288 (2037, 264, 1864);
  not ginst289 (2038, 1667);
  not ginst290 (2043, 1667);
  not ginst291 (2052, 1670);
  not ginst292 (2057, 1670);
  and ginst293 (2068, 50, 1197, 1869);
  and ginst294 (2073, 58, 1197, 1874);
  and ginst295 (2078, 68, 1197, 1879);
  and ginst296 (2083, 77, 1197, 1884);
  and ginst297 (2088, 87, 1219, 1889);
  and ginst298 (2093, 97, 1219, 1894);
  and ginst299 (2098, 107, 1219, 1899);
  and ginst300 (2103, 116, 1219, 1904);
  not ginst301 (2121, 1562);
  not ginst302 (2122, 1562);
  not ginst303 (2123, 1562);
  not ginst304 (2124, 1562);
  not ginst305 (2125, 1562);
  not ginst306 (2126, 1562);
  not ginst307 (2127, 1562);
  not ginst308 (2128, 1562);
  nand ginst309 (2133, 950, 1939);
  nand ginst310 (2134, 1478, 1941);
  nand ginst311 (2135, 1475, 1942);
  nand ginst312 (2136, 1484, 1943);
  nand ginst313 (2137, 1481, 1944);
  nand ginst314 (2138, 1490, 1945);
  nand ginst315 (2139, 1487, 1946);
  not ginst316 (2141, 1933);
  not ginst317 (2142, 1936);
  not ginst318 (2143, 1738);
  and ginst319 (2144, 1738, 1747);
  not ginst320 (2145, 1747);
  nand ginst321 (2146, 1727, 1960);
  nand ginst322 (2147, 1730, 1961);
  and ginst323 (2148, 1722, 1267, 665, 58);
  not ginst324 (2149, 1738);
  and ginst325 (2150, 1738, 1747);
  not ginst326 (2151, 1747);
  not ginst327 (2152, 1738);
  not ginst328 (2153, 1747);
  and ginst329 (2154, 1738, 1747);
  not ginst330 (2155, 1738);
  not ginst331 (2156, 1747);
  and ginst332 (2157, 1738, 1747);
  not ginst333 (2158, 1761);
  not ginst334 (2175, 1761);
  nand ginst335 (2178, 1764, 1981);
  nand ginst336 (2179, 1766, 1982);
  not ginst337 (2180, 1756);
  and ginst338 (2181, 1756, 1328);
  not ginst339 (2183, 1756);
  and ginst340 (2184, 1331, 1756);
  nand ginst341 (2185, 1358, 1812);
  nand ginst342 (2188, 1358, 1809);
  nand ginst343 (2191, 1353, 1812);
  nand ginst344 (2194, 1353, 1809);
  nand ginst345 (2197, 1358, 1806);
  nand ginst346 (2200, 1358, 1803);
  nand ginst347 (2203, 1353, 1806);
  nand ginst348 (2206, 1353, 1803);
  not ginst349 (2209, 1815);
  not ginst350 (2210, 1818);
  and ginst351 (2211, 1815, 1818);
  not ginst352 (2212, 1821);
  not ginst353 (2221, 1821);
  not ginst354 (2230, 1833);
  not ginst355 (2231, 1833);
  not ginst356 (2232, 1833);
  not ginst357 (2233, 1833);
  not ginst358 (2234, 1824);
  not ginst359 (2235, 1824);
  not ginst360 (2236, 1824);
  not ginst361 (2237, 1824);
  or ginst362 (2238, 2022, 1643, 2023);
  or ginst363 (2239, 2024, 1644, 2025);
  or ginst364 (2240, 2026, 1645, 2027);
  or ginst365 (2241, 2028, 1646, 2029);
  or ginst366 (2242, 2030, 1647, 2031);
  or ginst367 (2243, 2032, 1648, 2033);
  or ginst368 (2244, 2034, 1649, 2035);
  or ginst369 (2245, 2036, 1650, 2037);
  and ginst370 (2270, 1986, 1673);
  and ginst371 (2277, 1987, 1675);
  and ginst372 (2282, 1988, 1676);
  and ginst373 (2287, 1989, 1677);
  and ginst374 (2294, 1990, 1679);
  and ginst375 (2299, 1991, 1680);
  not ginst376 (2304, 1917);
  and ginst377 (2307, 1930, 350);
  nand ginst378 (2310, 1930, 350);
  not ginst379 (2313, 1715);
  not ginst380 (2316, 1718);
  not ginst381 (2319, 1715);
  not ginst382 (2322, 1718);
  nand ginst383 (2325, 1940, 2133);
  nand ginst384 (2328, 2134, 2135);
  nand ginst385 (2331, 2136, 2137);
  nand ginst386 (2334, 2138, 2139);
  nand ginst387 (2341, 1936, 2141);
  nand ginst388 (2342, 1933, 2142);
  and ginst389 (2347, 724, 2144);
  and ginst390 (2348, 2146, 699, 1726);
  and ginst391 (2349, 753, 2147);
  and ginst392 (2350, 2148, 1273);
  and ginst393 (2351, 736, 2150);
  and ginst394 (2352, 1735, 2153);
  and ginst395 (2353, 763, 2154);
  and ginst396 (2354, 1725, 2156);
  and ginst397 (2355, 749, 2157);
  not ginst398 (2374, 2178);
  not ginst399 (2375, 2179);
  and ginst400 (2376, 1520, 2180);
  and ginst401 (2379, 1721, 2181);
  and ginst402 (2398, 665, 2211);
  and ginst403 (2417, 2057, 226, 1873);
  and ginst404 (2418, 2057, 274, 1306);
  and ginst405 (2419, 2052, 2238);
  and ginst406 (2420, 2057, 232, 1878);
  and ginst407 (2421, 2057, 274, 1306);
  and ginst408 (2422, 2052, 2239);
  and ginst409 (2425, 2057, 238, 1883);
  and ginst410 (2426, 2057, 274, 1306);
  and ginst411 (2427, 2052, 2240);
  and ginst412 (2430, 2057, 244, 1888);
  and ginst413 (2431, 2057, 274, 1306);
  and ginst414 (2432, 2052, 2241);
  and ginst415 (2435, 2043, 250, 1893);
  and ginst416 (2436, 2043, 274, 1322);
  and ginst417 (2437, 2038, 2242);
  and ginst418 (2438, 2043, 257, 1898);
  and ginst419 (2439, 2043, 274, 1315);
  and ginst420 (2440, 2038, 2243);
  and ginst421 (2443, 2043, 264, 1903);
  and ginst422 (2444, 2043, 274, 1315);
  and ginst423 (2445, 2038, 2244);
  and ginst424 (2448, 2043, 270, 1908);
  and ginst425 (2449, 2043, 274, 1315);
  and ginst426 (2450, 2038, 2245);
  not ginst427 (2467, 2313);
  not ginst428 (2468, 2316);
  not ginst429 (2469, 2319);
  not ginst430 (2470, 2322);
  nand ginst431 (2471, 2341, 2342);
  not ginst432 (2474, 2325);
  not ginst433 (2475, 2328);
  not ginst434 (2476, 2331);
  not ginst435 (2477, 2334);
  or ginst436 (2478, 2348, 1729);
  not ginst437 (2481, 2175);
  and ginst438 (2482, 2175, 1334);
  and ginst439 (2483, 2349, 2183);
  and ginst440 (2486, 2374, 1346);
  and ginst441 (2487, 2375, 1350);
  not ginst442 (2488, 2185);
  not ginst443 (2497, 2188);
  not ginst444 (2506, 2191);
  not ginst445 (2515, 2194);
  not ginst446 (2524, 2197);
  not ginst447 (2533, 2200);
  not ginst448 (2542, 2203);
  not ginst449 (2551, 2206);
  not ginst450 (2560, 2185);
  not ginst451 (2569, 2188);
  not ginst452 (2578, 2191);
  not ginst453 (2587, 2194);
  not ginst454 (2596, 2197);
  not ginst455 (2605, 2200);
  not ginst456 (2614, 2203);
  not ginst457 (2623, 2206);
  not ginst458 (2632, 2212);
  and ginst459 (2633, 2212, 1833);
  not ginst460 (2634, 2212);
  and ginst461 (2635, 2212, 1833);
  not ginst462 (2636, 2212);
  and ginst463 (2637, 2212, 1833);
  not ginst464 (2638, 2212);
  and ginst465 (2639, 2212, 1833);
  not ginst466 (2640, 2221);
  and ginst467 (2641, 2221, 1824);
  not ginst468 (2642, 2221);
  and ginst469 (2643, 2221, 1824);
  not ginst470 (2644, 2221);
  and ginst471 (2645, 2221, 1824);
  not ginst472 (2646, 2221);
  and ginst473 (2647, 2221, 1824);
  or ginst474 (2648, 2270, 1870, 2068);
  nor ginst475 (2652, 2270, 1870, 2068);
  or ginst476 (2656, 2417, 2418, 2419);
  or ginst477 (2659, 2420, 2421, 2422);
  or ginst478 (2662, 2277, 1880, 2078);
  nor ginst479 (2666, 2277, 1880, 2078);
  or ginst480 (2670, 2425, 2426, 2427);
  or ginst481 (2673, 2282, 1885, 2083);
  nor ginst482 (2677, 2282, 1885, 2083);
  or ginst483 (2681, 2430, 2431, 2432);
  or ginst484 (2684, 2287, 1890, 2088);
  nor ginst485 (2688, 2287, 1890, 2088);
  or ginst486 (2692, 2435, 2436, 2437);
  or ginst487 (2697, 2438, 2439, 2440);
  or ginst488 (2702, 2294, 1900, 2098);
  nor ginst489 (2706, 2294, 1900, 2098);
  or ginst490 (2710, 2443, 2444, 2445);
  or ginst491 (2715, 2299, 1905, 2103);
  nor ginst492 (2719, 2299, 1905, 2103);
  or ginst493 (2723, 2448, 2449, 2450);
  not ginst494 (2728, 2304);
  not ginst495 (2729, 2158);
  and ginst496 (2730, 1562, 2158);
  not ginst497 (2731, 2158);
  and ginst498 (2732, 1562, 2158);
  not ginst499 (2733, 2158);
  and ginst500 (2734, 1562, 2158);
  not ginst501 (2735, 2158);
  and ginst502 (2736, 1562, 2158);
  not ginst503 (2737, 2158);
  and ginst504 (2738, 1562, 2158);
  not ginst505 (2739, 2158);
  and ginst506 (2740, 1562, 2158);
  not ginst507 (2741, 2158);
  and ginst508 (2742, 1562, 2158);
  not ginst509 (2743, 2158);
  and ginst510 (2744, 1562, 2158);
  or ginst511 (2745, 2376, 1983, 2379);
  nor ginst512 (2746, 2376, 1983, 2379);
  nand ginst513 (2748, 2316, 2467);
  nand ginst514 (2749, 2313, 2468);
  nand ginst515 (2750, 2322, 2469);
  nand ginst516 (2751, 2319, 2470);
  nand ginst517 (2754, 2328, 2474);
  nand ginst518 (2755, 2325, 2475);
  nand ginst519 (2756, 2334, 2476);
  nand ginst520 (2757, 2331, 2477);
  and ginst521 (2758, 1520, 2481);
  and ginst522 (2761, 1722, 2482);
  and ginst523 (2764, 2478, 1770);
  or ginst524 (2768, 2486, 1789, 1790);
  or ginst525 (2769, 2487, 1797, 1798);
  and ginst526 (2898, 665, 2633);
  and ginst527 (2899, 679, 2635);
  and ginst528 (2900, 686, 2637);
  and ginst529 (2901, 702, 2639);
  not ginst530 (2962, 2746);
  nand ginst531 (2966, 2748, 2749);
  nand ginst532 (2967, 2750, 2751);
  not ginst533 (2970, 2471);
  nand ginst534 (2973, 2754, 2755);
  nand ginst535 (2977, 2756, 2757);
  and ginst536 (2980, 2471, 2143);
  not ginst537 (2984, 2488);
  not ginst538 (2985, 2497);
  not ginst539 (2986, 2506);
  not ginst540 (2987, 2515);
  not ginst541 (2988, 2524);
  not ginst542 (2989, 2533);
  not ginst543 (2990, 2542);
  not ginst544 (2991, 2551);
  not ginst545 (2992, 2488);
  not ginst546 (2993, 2497);
  not ginst547 (2994, 2506);
  not ginst548 (2995, 2515);
  not ginst549 (2996, 2524);
  not ginst550 (2997, 2533);
  not ginst551 (2998, 2542);
  not ginst552 (2999, 2551);
  not ginst553 (3000, 2488);
  not ginst554 (3001, 2497);
  not ginst555 (3002, 2506);
  not ginst556 (3003, 2515);
  not ginst557 (3004, 2524);
  not ginst558 (3005, 2533);
  not ginst559 (3006, 2542);
  not ginst560 (3007, 2551);
  not ginst561 (3008, 2488);
  not ginst562 (3009, 2497);
  not ginst563 (3010, 2506);
  not ginst564 (3011, 2515);
  not ginst565 (3012, 2524);
  not ginst566 (3013, 2533);
  not ginst567 (3014, 2542);
  not ginst568 (3015, 2551);
  not ginst569 (3016, 2488);
  not ginst570 (3017, 2497);
  not ginst571 (3018, 2506);
  not ginst572 (3019, 2515);
  not ginst573 (3020, 2524);
  not ginst574 (3021, 2533);
  not ginst575 (3022, 2542);
  not ginst576 (3023, 2551);
  not ginst577 (3024, 2488);
  not ginst578 (3025, 2497);
  not ginst579 (3026, 2506);
  not ginst580 (3027, 2515);
  not ginst581 (3028, 2524);
  not ginst582 (3029, 2533);
  not ginst583 (3030, 2542);
  not ginst584 (3031, 2551);
  not ginst585 (3032, 2488);
  not ginst586 (3033, 2497);
  not ginst587 (3034, 2506);
  not ginst588 (3035, 2515);
  not ginst589 (3036, 2524);
  not ginst590 (3037, 2533);
  not ginst591 (3038, 2542);
  not ginst592 (3039, 2551);
  not ginst593 (3040, 2488);
  not ginst594 (3041, 2497);
  not ginst595 (3042, 2506);
  not ginst596 (3043, 2515);
  not ginst597 (3044, 2524);
  not ginst598 (3045, 2533);
  not ginst599 (3046, 2542);
  not ginst600 (3047, 2551);
  not ginst601 (3048, 2560);
  not ginst602 (3049, 2569);
  not ginst603 (3050, 2578);
  not ginst604 (3051, 2587);
  not ginst605 (3052, 2596);
  not ginst606 (3053, 2605);
  not ginst607 (3054, 2614);
  not ginst608 (3055, 2623);
  not ginst609 (3056, 2560);
  not ginst610 (3057, 2569);
  not ginst611 (3058, 2578);
  not ginst612 (3059, 2587);
  not ginst613 (3060, 2596);
  not ginst614 (3061, 2605);
  not ginst615 (3062, 2614);
  not ginst616 (3063, 2623);
  not ginst617 (3064, 2560);
  not ginst618 (3065, 2569);
  not ginst619 (3066, 2578);
  not ginst620 (3067, 2587);
  not ginst621 (3068, 2596);
  not ginst622 (3069, 2605);
  not ginst623 (3070, 2614);
  not ginst624 (3071, 2623);
  not ginst625 (3072, 2560);
  not ginst626 (3073, 2569);
  not ginst627 (3074, 2578);
  not ginst628 (3075, 2587);
  not ginst629 (3076, 2596);
  not ginst630 (3077, 2605);
  not ginst631 (3078, 2614);
  not ginst632 (3079, 2623);
  not ginst633 (3080, 2560);
  not ginst634 (3081, 2569);
  not ginst635 (3082, 2578);
  not ginst636 (3083, 2587);
  not ginst637 (3084, 2596);
  not ginst638 (3085, 2605);
  not ginst639 (3086, 2614);
  not ginst640 (3087, 2623);
  not ginst641 (3088, 2560);
  not ginst642 (3089, 2569);
  not ginst643 (3090, 2578);
  not ginst644 (3091, 2587);
  not ginst645 (3092, 2596);
  not ginst646 (3093, 2605);
  not ginst647 (3094, 2614);
  not ginst648 (3095, 2623);
  not ginst649 (3096, 2560);
  not ginst650 (3097, 2569);
  not ginst651 (3098, 2578);
  not ginst652 (3099, 2587);
  not ginst653 (3100, 2596);
  not ginst654 (3101, 2605);
  not ginst655 (3102, 2614);
  not ginst656 (3103, 2623);
  not ginst657 (3104, 2560);
  not ginst658 (3105, 2569);
  not ginst659 (3106, 2578);
  not ginst660 (3107, 2587);
  not ginst661 (3108, 2596);
  not ginst662 (3109, 2605);
  not ginst663 (3110, 2614);
  not ginst664 (3111, 2623);
  not ginst665 (3112, 2656);
  not ginst666 (3115, 2656);
  not ginst667 (3118, 2652);
  and ginst668 (3119, 2768, 1674);
  not ginst669 (3122, 2659);
  not ginst670 (3125, 2659);
  not ginst671 (3128, 2670);
  not ginst672 (3131, 2670);
  not ginst673 (3134, 2666);
  not ginst674 (3135, 2681);
  not ginst675 (3138, 2681);
  not ginst676 (3141, 2677);
  not ginst677 (3142, 2692);
  not ginst678 (3145, 2692);
  not ginst679 (3148, 2688);
  and ginst680 (3149, 2769, 1678);
  not ginst681 (3152, 2697);
  not ginst682 (3155, 2697);
  not ginst683 (3158, 2710);
  not ginst684 (3161, 2710);
  not ginst685 (3164, 2706);
  not ginst686 (3165, 2723);
  not ginst687 (3168, 2723);
  not ginst688 (3171, 2719);
  and ginst689 (3172, 1909, 2648);
  and ginst690 (3175, 1913, 2662);
  and ginst691 (3178, 1913, 2673);
  and ginst692 (3181, 1913, 2684);
  and ginst693 (3184, 1922, 2702);
  and ginst694 (3187, 1922, 2715);
  not ginst695 (3190, 2692);
  not ginst696 (3191, 2697);
  not ginst697 (3192, 2710);
  not ginst698 (3193, 2723);
  and ginst699 (3194, 2692, 2697, 2710, 2723, 1459);
  nand ginst700 (3195, 2745, 2962);
  not ginst701 (3196, 2966);
  or ginst702 (3206, 2980, 2145, 2347);
  and ginst703 (3207, 124, 2984);
  and ginst704 (3208, 159, 2985);
  and ginst705 (3209, 150, 2986);
  and ginst706 (3210, 143, 2987);
  and ginst707 (3211, 137, 2988);
  and ginst708 (3212, 132, 2989);
  and ginst709 (3213, 128, 2990);
  and ginst710 (3214, 125, 2991);
  and ginst711 (3215, 125, 2992);
  and ginst712 (3216, 655, 2993);
  and ginst713 (3217, 159, 2994);
  and ginst714 (3218, 150, 2995);
  and ginst715 (3219, 143, 2996);
  and ginst716 (3220, 137, 2997);
  and ginst717 (3221, 132, 2998);
  and ginst718 (3222, 128, 2999);
  and ginst719 (3223, 128, 3000);
  and ginst720 (3224, 670, 3001);
  and ginst721 (3225, 655, 3002);
  and ginst722 (3226, 159, 3003);
  and ginst723 (3227, 150, 3004);
  and ginst724 (3228, 143, 3005);
  and ginst725 (3229, 137, 3006);
  and ginst726 (3230, 132, 3007);
  and ginst727 (3231, 132, 3008);
  and ginst728 (3232, 690, 3009);
  and ginst729 (3233, 670, 3010);
  and ginst730 (3234, 655, 3011);
  and ginst731 (3235, 159, 3012);
  and ginst732 (3236, 150, 3013);
  and ginst733 (3237, 143, 3014);
  and ginst734 (3238, 137, 3015);
  and ginst735 (3239, 137, 3016);
  and ginst736 (3240, 706, 3017);
  and ginst737 (3241, 690, 3018);
  and ginst738 (3242, 670, 3019);
  and ginst739 (3243, 655, 3020);
  and ginst740 (3244, 159, 3021);
  and ginst741 (3245, 150, 3022);
  and ginst742 (3246, 143, 3023);
  and ginst743 (3247, 143, 3024);
  and ginst744 (3248, 715, 3025);
  and ginst745 (3249, 706, 3026);
  and ginst746 (3250, 690, 3027);
  and ginst747 (3251, 670, 3028);
  and ginst748 (3252, 655, 3029);
  and ginst749 (3253, 159, 3030);
  and ginst750 (3254, 150, 3031);
  and ginst751 (3255, 150, 3032);
  and ginst752 (3256, 727, 3033);
  and ginst753 (3257, 715, 3034);
  and ginst754 (3258, 706, 3035);
  and ginst755 (3259, 690, 3036);
  and ginst756 (3260, 670, 3037);
  and ginst757 (3261, 655, 3038);
  and ginst758 (3262, 159, 3039);
  and ginst759 (3263, 159, 3040);
  and ginst760 (3264, 740, 3041);
  and ginst761 (3265, 727, 3042);
  and ginst762 (3266, 715, 3043);
  and ginst763 (3267, 706, 3044);
  and ginst764 (3268, 690, 3045);
  and ginst765 (3269, 670, 3046);
  and ginst766 (3270, 655, 3047);
  and ginst767 (3271, 283, 3048);
  and ginst768 (3272, 670, 3049);
  and ginst769 (3273, 690, 3050);
  and ginst770 (3274, 706, 3051);
  and ginst771 (3275, 715, 3052);
  and ginst772 (3276, 727, 3053);
  and ginst773 (3277, 740, 3054);
  and ginst774 (3278, 753, 3055);
  and ginst775 (3279, 294, 3056);
  and ginst776 (3280, 690, 3057);
  and ginst777 (3281, 706, 3058);
  and ginst778 (3282, 715, 3059);
  and ginst779 (3283, 727, 3060);
  and ginst780 (3284, 740, 3061);
  and ginst781 (3285, 753, 3062);
  and ginst782 (3286, 283, 3063);
  and ginst783 (3287, 303, 3064);
  and ginst784 (3288, 706, 3065);
  and ginst785 (3289, 715, 3066);
  and ginst786 (3290, 727, 3067);
  and ginst787 (3291, 740, 3068);
  and ginst788 (3292, 753, 3069);
  and ginst789 (3293, 283, 3070);
  and ginst790 (3294, 294, 3071);
  and ginst791 (3295, 311, 3072);
  and ginst792 (3296, 715, 3073);
  and ginst793 (3297, 727, 3074);
  and ginst794 (3298, 740, 3075);
  and ginst795 (3299, 753, 3076);
  and ginst796 (3300, 283, 3077);
  and ginst797 (3301, 294, 3078);
  and ginst798 (3302, 303, 3079);
  and ginst799 (3303, 317, 3080);
  and ginst800 (3304, 727, 3081);
  and ginst801 (3305, 740, 3082);
  and ginst802 (3306, 753, 3083);
  and ginst803 (3307, 283, 3084);
  and ginst804 (3308, 294, 3085);
  and ginst805 (3309, 303, 3086);
  and ginst806 (3310, 311, 3087);
  and ginst807 (3311, 322, 3088);
  and ginst808 (3312, 740, 3089);
  and ginst809 (3313, 753, 3090);
  and ginst810 (3314, 283, 3091);
  and ginst811 (3315, 294, 3092);
  and ginst812 (3316, 303, 3093);
  and ginst813 (3317, 311, 3094);
  and ginst814 (3318, 317, 3095);
  and ginst815 (3319, 326, 3096);
  and ginst816 (3320, 753, 3097);
  and ginst817 (3321, 283, 3098);
  and ginst818 (3322, 294, 3099);
  and ginst819 (3323, 303, 3100);
  and ginst820 (3324, 311, 3101);
  and ginst821 (3325, 317, 3102);
  and ginst822 (3326, 322, 3103);
  and ginst823 (3327, 329, 3104);
  and ginst824 (3328, 283, 3105);
  and ginst825 (3329, 294, 3106);
  and ginst826 (3330, 303, 3107);
  and ginst827 (3331, 311, 3108);
  and ginst828 (3332, 317, 3109);
  and ginst829 (3333, 322, 3110);
  and ginst830 (3334, 326, 3111);
  and ginst831 (3383, 3190, 3191, 3192, 3193, 917);
  not ginst832 (3384, 2977);
  and ginst833 (3387, 3196, 1736);
  and ginst834 (3388, 2977, 2149);
  and ginst835 (3389, 2973, 1737);
  nor ginst836 (3390, 3207, 3208, 3209, 3210, 3211, 3212, 3213, 3214);
  nor ginst837 (3391, 3215, 3216, 3217, 3218, 3219, 3220, 3221, 3222);
  nor ginst838 (3392, 3223, 3224, 3225, 3226, 3227, 3228, 3229, 3230);
  nor ginst839 (3393, 3231, 3232, 3233, 3234, 3235, 3236, 3237, 3238);
  nor ginst840 (3394, 3239, 3240, 3241, 3242, 3243, 3244, 3245, 3246);
  nor ginst841 (3395, 3247, 3248, 3249, 3250, 3251, 3252, 3253, 3254);
  nor ginst842 (3396, 3255, 3256, 3257, 3258, 3259, 3260, 3261, 3262);
  nor ginst843 (3397, 3263, 3264, 3265, 3266, 3267, 3268, 3269, 3270);
  nor ginst844 (3398, 3271, 3272, 3273, 3274, 3275, 3276, 3277, 3278);
  nor ginst845 (3399, 3279, 3280, 3281, 3282, 3283, 3284, 3285, 3286);
  nor ginst846 (3400, 3287, 3288, 3289, 3290, 3291, 3292, 3293, 3294);
  nor ginst847 (3401, 3295, 3296, 3297, 3298, 3299, 3300, 3301, 3302);
  nor ginst848 (3402, 3303, 3304, 3305, 3306, 3307, 3308, 3309, 3310);
  nor ginst849 (3403, 3311, 3312, 3313, 3314, 3315, 3316, 3317, 3318);
  nor ginst850 (3404, 3319, 3320, 3321, 3322, 3323, 3324, 3325, 3326);
  nor ginst851 (3405, 3327, 3328, 3329, 3330, 3331, 3332, 3333, 3334);
  and ginst852 (3406, 3206, 2641);
  and ginst853 (3407, 169, 2648, 3112);
  and ginst854 (3410, 179, 2648, 3115);
  and ginst855 (3413, 190, 2652, 3115);
  and ginst856 (3414, 200, 2652, 3112);
  or ginst857 (3415, 3119, 1875, 2073);
  nor ginst858 (3419, 3119, 1875, 2073);
  and ginst859 (3423, 169, 2662, 3128);
  and ginst860 (3426, 179, 2662, 3131);
  and ginst861 (3429, 190, 2666, 3131);
  and ginst862 (3430, 200, 2666, 3128);
  and ginst863 (3431, 169, 2673, 3135);
  and ginst864 (3434, 179, 2673, 3138);
  and ginst865 (3437, 190, 2677, 3138);
  and ginst866 (3438, 200, 2677, 3135);
  and ginst867 (3439, 169, 2684, 3142);
  and ginst868 (3442, 179, 2684, 3145);
  and ginst869 (3445, 190, 2688, 3145);
  and ginst870 (3446, 200, 2688, 3142);
  or ginst871 (3447, 3149, 1895, 2093);
  nor ginst872 (3451, 3149, 1895, 2093);
  and ginst873 (3455, 169, 2702, 3158);
  and ginst874 (3458, 179, 2702, 3161);
  and ginst875 (3461, 190, 2706, 3161);
  and ginst876 (3462, 200, 2706, 3158);
  and ginst877 (3463, 169, 2715, 3165);
  and ginst878 (3466, 179, 2715, 3168);
  and ginst879 (3469, 190, 2719, 3168);
  and ginst880 (3470, 200, 2719, 3165);
  or ginst881 (3471, 3194, 3383);
  not ginst882 (3472, 2967);
  not ginst883 (3475, 2970);
  not ginst884 (3478, 2967);
  not ginst885 (3481, 2970);
  not ginst886 (3484, 2973);
  not ginst887 (3487, 2973);
  not ginst888 (3490, 3172);
  not ginst889 (3493, 3172);
  not ginst890 (3496, 3175);
  not ginst891 (3499, 3175);
  not ginst892 (3502, 3178);
  not ginst893 (3505, 3178);
  not ginst894 (3508, 3181);
  not ginst895 (3511, 3181);
  not ginst896 (3514, 3184);
  not ginst897 (3517, 3184);
  not ginst898 (3520, 3187);
  not ginst899 (3523, 3187);
  nor ginst900 (3534, 3387, 2350);
  or ginst901 (3535, 3388, 2151, 2351);
  nor ginst902 (3536, 3389, 1966);
  and ginst903 (3537, 3390, 2209);
  and ginst904 (3538, 3398, 2210);
  and ginst905 (3539, 3391, 1842);
  and ginst906 (3540, 3399, 1369);
  and ginst907 (3541, 3392, 1843);
  and ginst908 (3542, 3400, 1369);
  and ginst909 (3543, 3393, 1844);
  and ginst910 (3544, 3401, 1369);
  and ginst911 (3545, 3394, 1845);
  and ginst912 (3546, 3402, 1369);
  and ginst913 (3547, 3395, 1846);
  and ginst914 (3548, 3403, 1369);
  and ginst915 (3549, 3396, 1847);
  and ginst916 (3550, 3404, 1369);
  and ginst917 (3551, 3397, 1848);
  and ginst918 (3552, 3405, 1369);
  or ginst919 (3557, 3413, 3414, 3118);
  or ginst920 (3568, 3429, 3430, 3134);
  or ginst921 (3573, 3437, 3438, 3141);
  or ginst922 (3578, 3445, 3446, 3148);
  or ginst923 (3589, 3461, 3462, 3164);
  or ginst924 (3594, 3469, 3470, 3171);
  and ginst925 (3605, 3471, 2728);
  not ginst926 (3626, 3478);
  not ginst927 (3627, 3481);
  not ginst928 (3628, 3487);
  not ginst929 (3629, 3484);
  not ginst930 (3630, 3472);
  not ginst931 (3631, 3475);
  and ginst932 (3632, 3536, 2152);
  and ginst933 (3633, 3534, 2155);
  or ginst934 (3634, 3537, 3538, 2398);
  or ginst935 (3635, 3539, 3540);
  or ginst936 (3636, 3541, 3542);
  or ginst937 (3637, 3543, 3544);
  or ginst938 (3638, 3545, 3546);
  or ginst939 (3639, 3547, 3548);
  or ginst940 (3640, 3549, 3550);
  or ginst941 (3641, 3551, 3552);
  and ginst942 (3642, 3535, 2643);
  or ginst943 (3643, 3407, 3410);
  nor ginst944 (3644, 3407, 3410);
  and ginst945 (3645, 169, 3415, 3122);
  and ginst946 (3648, 179, 3415, 3125);
  and ginst947 (3651, 190, 3419, 3125);
  and ginst948 (3652, 200, 3419, 3122);
  not ginst949 (3653, 3419);
  or ginst950 (3654, 3423, 3426);
  nor ginst951 (3657, 3423, 3426);
  or ginst952 (3658, 3431, 3434);
  nor ginst953 (3661, 3431, 3434);
  or ginst954 (3662, 3439, 3442);
  nor ginst955 (3663, 3439, 3442);
  and ginst956 (3664, 169, 3447, 3152);
  and ginst957 (3667, 179, 3447, 3155);
  and ginst958 (3670, 190, 3451, 3155);
  and ginst959 (3671, 200, 3451, 3152);
  not ginst960 (3672, 3451);
  or ginst961 (3673, 3455, 3458);
  nor ginst962 (3676, 3455, 3458);
  or ginst963 (3677, 3463, 3466);
  nor ginst964 (3680, 3463, 3466);
  not ginst965 (3681, 3493);
  and ginst966 (3682, 1909, 3415);
  not ginst967 (3685, 3496);
  not ginst968 (3686, 3499);
  not ginst969 (3687, 3502);
  not ginst970 (3688, 3505);
  not ginst971 (3689, 3511);
  and ginst972 (3690, 1922, 3447);
  not ginst973 (3693, 3517);
  not ginst974 (3694, 3520);
  not ginst975 (3695, 3523);
  not ginst976 (3696, 3514);
  not ginst977 (3697, 3384);
  not ginst978 (3700, 3384);
  not ginst979 (3703, 3490);
  not ginst980 (3704, 3508);
  nand ginst981 (3705, 3475, 3630);
  nand ginst982 (3706, 3472, 3631);
  nand ginst983 (3707, 3481, 3626);
  nand ginst984 (3708, 3478, 3627);
  or ginst985 (3711, 3632, 2352, 2353);
  or ginst986 (3712, 3633, 2354, 2355);
  and ginst987 (3713, 3634, 2632);
  and ginst988 (3714, 3635, 2634);
  and ginst989 (3715, 3636, 2636);
  and ginst990 (3716, 3637, 2638);
  and ginst991 (3717, 3638, 2640);
  and ginst992 (3718, 3639, 2642);
  and ginst993 (3719, 3640, 2644);
  and ginst994 (3720, 3641, 2646);
  and ginst995 (3721, 3644, 3557);
  or ginst996 (3731, 3651, 3652, 3653);
  and ginst997 (3734, 3657, 3568);
  and ginst998 (3740, 3661, 3573);
  and ginst999 (3743, 3663, 3578);
  or ginst1000 (3753, 3670, 3671, 3672);
  and ginst1001 (3756, 3676, 3589);
  and ginst1002 (3762, 3680, 3594);
  not ginst1003 (3765, 3643);
  not ginst1004 (3766, 3662);
  nand ginst1005 (3773, 3705, 3706);
  nand ginst1006 (3774, 3707, 3708);
  nand ginst1007 (3775, 3700, 3628);
  not ginst1008 (3776, 3700);
  nand ginst1009 (3777, 3697, 3629);
  not ginst1010 (3778, 3697);
  and ginst1011 (3779, 3712, 2645);
  and ginst1012 (3780, 3711, 2647);
  or ginst1013 (3786, 3645, 3648);
  nor ginst1014 (3789, 3645, 3648);
  or ginst1015 (3800, 3664, 3667);
  nor ginst1016 (3803, 3664, 3667);
  and ginst1017 (3809, 3654, 1917);
  and ginst1018 (3812, 3658, 1917);
  and ginst1019 (3815, 3673, 1926);
  and ginst1020 (3818, 3677, 1926);
  not ginst1021 (3821, 3682);
  not ginst1022 (3824, 3682);
  not ginst1023 (3827, 3690);
  not ginst1024 (3830, 3690);
  nand ginst1025 (3833, 3773, 3774);
  nand ginst1026 (3834, 3487, 3776);
  nand ginst1027 (3835, 3484, 3778);
  and ginst1028 (3838, 3789, 3731);
  and ginst1029 (3845, 3803, 3753);
  not ginst1030 (3850, 3721);
  not ginst1031 (3855, 3734);
  not ginst1032 (3858, 3740);
  not ginst1033 (3861, 3743);
  not ginst1034 (3865, 3756);
  not ginst1035 (3868, 3762);
  nand ginst1036 (3884, 3775, 3834);
  nand ginst1037 (3885, 3777, 3835);
  nand ginst1038 (3894, 3721, 3786);
  nand ginst1039 (3895, 3743, 3800);
  not ginst1040 (3898, 3821);
  not ginst1041 (3899, 3824);
  not ginst1042 (3906, 3830);
  not ginst1043 (3911, 3827);
  and ginst1044 (3912, 3786, 1912);
  not ginst1045 (3913, 3812);
  and ginst1046 (3916, 3800, 1917);
  not ginst1047 (3917, 3818);
  not ginst1048 (3920, 3809);
  not ginst1049 (3921, 3818);
  not ginst1050 (3924, 3884);
  not ginst1051 (3925, 3885);
  and ginst1052 (3926, 3721, 3838, 3734, 3740);
  nand ginst1053 (3930, 3721, 3838, 3654);
  nand ginst1054 (3931, 3658, 3838, 3734, 3721);
  and ginst1055 (3932, 3743, 3845, 3756, 3762);
  nand ginst1056 (3935, 3743, 3845, 3673);
  nand ginst1057 (3936, 3677, 3845, 3756, 3743);
  not ginst1058 (3937, 3838);
  not ginst1059 (3940, 3845);
  not ginst1060 (3947, 3912);
  not ginst1061 (3948, 3916);
  not ginst1062 (3950, 3850);
  not ginst1063 (3953, 3850);
  not ginst1064 (3956, 3855);
  not ginst1065 (3959, 3855);
  not ginst1066 (3962, 3858);
  not ginst1067 (3965, 3858);
  not ginst1068 (3968, 3861);
  not ginst1069 (3971, 3861);
  not ginst1070 (3974, 3865);
  not ginst1071 (3977, 3865);
  not ginst1072 (3980, 3868);
  not ginst1073 (3983, 3868);
  nand ginst1074 (3987, 3924, 3925);
  nand ginst1075 (3992, 3765, 3894, 3930, 3931);
  nand ginst1076 (3996, 3766, 3895, 3935, 3936);
  not ginst1077 (4013, 3921);
  and ginst1078 (4028, 3932, 3926);
  nand ginst1079 (4029, 3953, 3681);
  nand ginst1080 (4030, 3959, 3686);
  nand ginst1081 (4031, 3965, 3688);
  nand ginst1082 (4032, 3971, 3689);
  nand ginst1083 (4033, 3977, 3693);
  nand ginst1084 (4034, 3983, 3695);
  not ginst1085 (4035, 3926);
  not ginst1086 (4042, 3953);
  not ginst1087 (4043, 3956);
  nand ginst1088 (4044, 3956, 3685);
  not ginst1089 (4045, 3959);
  not ginst1090 (4046, 3962);
  nand ginst1091 (4047, 3962, 3687);
  not ginst1092 (4048, 3965);
  not ginst1093 (4049, 3971);
  not ginst1094 (4050, 3977);
  not ginst1095 (4051, 3980);
  nand ginst1096 (4052, 3980, 3694);
  not ginst1097 (4053, 3983);
  not ginst1098 (4054, 3974);
  nand ginst1099 (4055, 3974, 3696);
  and ginst1100 (4056, 3932, 2304);
  not ginst1101 (4057, 3950);
  nand ginst1102 (4058, 3950, 3703);
  not ginst1103 (4059, 3937);
  not ginst1104 (4062, 3937);
  not ginst1105 (4065, 3968);
  nand ginst1106 (4066, 3968, 3704);
  not ginst1107 (4067, 3940);
  not ginst1108 (4070, 3940);
  nand ginst1109 (4073, 3926, 3996);
  not ginst1110 (4074, 3992);
  nand ginst1111 (4075, 3493, 4042);
  nand ginst1112 (4076, 3499, 4045);
  nand ginst1113 (4077, 3505, 4048);
  nand ginst1114 (4078, 3511, 4049);
  nand ginst1115 (4079, 3517, 4050);
  nand ginst1116 (4080, 3523, 4053);
  nand ginst1117 (4085, 3496, 4043);
  nand ginst1118 (4086, 3502, 4046);
  nand ginst1119 (4088, 3520, 4051);
  nand ginst1120 (4090, 3514, 4054);
  and ginst1121 (4091, 3996, 1926);
  or ginst1122 (4094, 3605, 4056);
  nand ginst1123 (4098, 3490, 4057);
  nand ginst1124 (4101, 3508, 4065);
  and ginst1125 (4104, 4073, 4074);
  nand ginst1126 (4105, 4075, 4029);
  nand ginst1127 (4106, 4062, 3899);
  nand ginst1128 (4107, 4076, 4030);
  nand ginst1129 (4108, 4077, 4031);
  nand ginst1130 (4109, 4078, 4032);
  nand ginst1131 (4110, 4070, 3906);
  nand ginst1132 (4111, 4079, 4033);
  nand ginst1133 (4112, 4080, 4034);
  not ginst1134 (4113, 4059);
  nand ginst1135 (4114, 4059, 3898);
  not ginst1136 (4115, 4062);
  nand ginst1137 (4116, 4085, 4044);
  nand ginst1138 (4119, 4086, 4047);
  not ginst1139 (4122, 4070);
  nand ginst1140 (4123, 4088, 4052);
  not ginst1141 (4126, 4067);
  nand ginst1142 (4127, 4067, 3911);
  nand ginst1143 (4128, 4090, 4055);
  nand ginst1144 (4139, 4098, 4058);
  nand ginst1145 (4142, 4101, 4066);
  not ginst1146 (4145, 4104);
  not ginst1147 (4146, 4105);
  nand ginst1148 (4147, 3824, 4115);
  not ginst1149 (4148, 4107);
  not ginst1150 (4149, 4108);
  not ginst1151 (4150, 4109);
  nand ginst1152 (4151, 3830, 4122);
  not ginst1153 (4152, 4111);
  not ginst1154 (4153, 4112);
  nand ginst1155 (4154, 3821, 4113);
  nand ginst1156 (4161, 3827, 4126);
  not ginst1157 (4167, 4091);
  not ginst1158 (4174, 4094);
  not ginst1159 (4182, 4091);
  and ginst1160 (4186, 330, 4094);
  and ginst1161 (4189, 4146, 2230);
  nand ginst1162 (4190, 4147, 4106);
  and ginst1163 (4191, 4148, 2232);
  and ginst1164 (4192, 4149, 2233);
  and ginst1165 (4193, 4150, 2234);
  nand ginst1166 (4194, 4151, 4110);
  and ginst1167 (4195, 4152, 2236);
  and ginst1168 (4196, 4153, 2237);
  nand ginst1169 (4197, 4154, 4114);
  not ginst1170 (4200, 4116);
  not ginst1171 (4203, 4116);
  not ginst1172 (4209, 4119);
  not ginst1173 (4213, 4119);
  nand ginst1174 (4218, 4161, 4127);
  not ginst1175 (4223, 4123);
  and ginst1176 (4238, 4128, 3917);
  not ginst1177 (4239, 4139);
  not ginst1178 (4241, 4142);
  and ginst1179 (4242, 330, 4123);
  not ginst1180 (4247, 4128);
  nor ginst1181 (4251, 3713, 4189, 2898);
  not ginst1182 (4252, 4190);
  nor ginst1183 (4253, 3715, 4191, 2900);
  nor ginst1184 (4254, 3716, 4192, 2901);
  nor ginst1185 (4255, 3717, 4193, 3406);
  not ginst1186 (4256, 4194);
  nor ginst1187 (4257, 3719, 4195, 3779);
  nor ginst1188 (4258, 3720, 4196, 3780);
  and ginst1189 (4283, 4167, 4035);
  and ginst1190 (4284, 4174, 4035);
  or ginst1191 (4287, 3815, 4238);
  not ginst1192 (4291, 4186);
  not ginst1193 (4295, 4167);
  not ginst1194 (4296, 4167);
  not ginst1195 (4299, 4182);
  and ginst1196 (4303, 4252, 2231);
  and ginst1197 (4304, 4256, 2235);
  not ginst1198 (4305, 4197);
  or ginst1199 (4310, 3992, 4283);
  and ginst1200 (4316, 4174, 4213, 4203);
  and ginst1201 (4317, 4174, 4209);
  and ginst1202 (4318, 4223, 4128, 4218);
  and ginst1203 (4319, 4223, 4128);
  and ginst1204 (4322, 4167, 4209);
  nand ginst1205 (4325, 4203, 3913);
  nand ginst1206 (4326, 4203, 4213, 4167);
  nand ginst1207 (4327, 4218, 3815);
  nand ginst1208 (4328, 4218, 4128, 3917);
  nand ginst1209 (4329, 4247, 4013);
  not ginst1210 (4330, 4247);
  and ginst1211 (4331, 330, 4094, 4295);
  and ginst1212 (4335, 4251, 2730);
  and ginst1213 (4338, 4253, 2734);
  and ginst1214 (4341, 4254, 2736);
  and ginst1215 (4344, 4255, 2738);
  and ginst1216 (4347, 4257, 2742);
  and ginst1217 (4350, 4258, 2744);
  not ginst1218 (4353, 4197);
  not ginst1219 (4356, 4203);
  not ginst1220 (4359, 4209);
  not ginst1221 (4362, 4218);
  not ginst1222 (4365, 4242);
  not ginst1223 (4368, 4242);
  and ginst1224 (4371, 4223, 4223);
  nor ginst1225 (4376, 3714, 4303, 2899);
  nor ginst1226 (4377, 3718, 4304, 3642);
  and ginst1227 (4387, 330, 4317);
  and ginst1228 (4390, 330, 4318);
  nand ginst1229 (4393, 3921, 4330);
  not ginst1230 (4398, 4287);
  not ginst1231 (4413, 4284);
  nand ginst1232 (4416, 3920, 4325, 4326);
  or ginst1233 (4421, 3812, 4322);
  nand ginst1234 (4427, 3948, 4327, 4328);
  not ginst1235 (4430, 4287);
  and ginst1236 (4435, 330, 4316);
  or ginst1237 (4442, 4331, 4296);
  and ginst1238 (4443, 4174, 4305, 4203, 4213);
  nand ginst1239 (4446, 4305, 3809);
  nand ginst1240 (4447, 4305, 4200, 3913);
  nand ginst1241 (4448, 4305, 4200, 4213, 4167);
  not ginst1242 (4452, 4356);
  nand ginst1243 (4458, 4329, 4393);
  not ginst1244 (4461, 4365);
  not ginst1245 (4462, 4368);
  nand ginst1246 (4463, 4371, 1460);
  not ginst1247 (4464, 4371);
  not ginst1248 (4465, 4310);
  nor ginst1249 (4468, 4331, 4296);
  and ginst1250 (4472, 4376, 2732);
  and ginst1251 (4475, 4377, 2740);
  not ginst1252 (4479, 4310);
  not ginst1253 (4484, 4353);
  not ginst1254 (4486, 4359);
  nand ginst1255 (4487, 4359, 4299);
  not ginst1256 (4491, 4362);
  and ginst1257 (4493, 330, 4319);
  not ginst1258 (4496, 4398);
  and ginst1259 (4497, 4287, 4398);
  and ginst1260 (4498, 4442, 1769);
  nand ginst1261 (4503, 3947, 4446, 4447, 4448);
  not ginst1262 (4506, 4413);
  not ginst1263 (4507, 4435);
  not ginst1264 (4508, 4421);
  nand ginst1265 (4509, 4421, 4452);
  not ginst1266 (4510, 4427);
  nand ginst1267 (4511, 4427, 4241);
  nand ginst1268 (4515, 965, 4464);
  not ginst1269 (4526, 4416);
  nand ginst1270 (4527, 4416, 4484);
  nand ginst1271 (4528, 4182, 4486);
  not ginst1272 (4529, 4430);
  nand ginst1273 (4530, 4430, 4491);
  not ginst1274 (4531, 4387);
  not ginst1275 (4534, 4387);
  not ginst1276 (4537, 4390);
  not ginst1277 (4540, 4390);
  and ginst1278 (4545, 330, 4319, 4496);
  and ginst1279 (4549, 330, 4443);
  nand ginst1280 (4552, 4356, 4508);
  nand ginst1281 (4555, 4142, 4510);
  not ginst1282 (4558, 4493);
  nand ginst1283 (4559, 4463, 4515);
  not ginst1284 (4562, 4465);
  and ginst1285 (4563, 4310, 4465);
  not ginst1286 (4564, 4468);
  not ginst1287 (4568, 4479);
  not ginst1288 (4569, 4443);
  nand ginst1289 (4572, 4353, 4526);
  nand ginst1290 (4573, 4362, 4529);
  nand ginst1291 (4576, 4487, 4528);
  not ginst1292 (4581, 4458);
  not ginst1293 (4584, 4458);
  or ginst1294 (4587, 2758, 4498, 2761);
  nor ginst1295 (4588, 2758, 4498, 2761);
  or ginst1296 (4589, 4545, 4497);
  nand ginst1297 (4593, 4552, 4509);
  not ginst1298 (4596, 4531);
  not ginst1299 (4597, 4534);
  nand ginst1300 (4599, 4555, 4511);
  not ginst1301 (4602, 4537);
  not ginst1302 (4603, 4540);
  and ginst1303 (4608, 330, 4284, 4562);
  not ginst1304 (4613, 4503);
  not ginst1305 (4616, 4503);
  nand ginst1306 (4619, 4572, 4527);
  nand ginst1307 (4623, 4573, 4530);
  not ginst1308 (4628, 4588);
  nand ginst1309 (4629, 4569, 4506);
  not ginst1310 (4630, 4569);
  not ginst1311 (4635, 4576);
  nand ginst1312 (4636, 4576, 4291);
  not ginst1313 (4640, 4581);
  nand ginst1314 (4641, 4581, 4461);
  not ginst1315 (4642, 4584);
  nand ginst1316 (4643, 4584, 4462);
  nor ginst1317 (4644, 4608, 4563);
  and ginst1318 (4647, 4559, 2128);
  and ginst1319 (4650, 4559, 2743);
  not ginst1320 (4656, 4549);
  not ginst1321 (4659, 4549);
  not ginst1322 (4664, 4564);
  and ginst1323 (4667, 4587, 4628);
  nand ginst1324 (4668, 4413, 4630);
  not ginst1325 (4669, 4616);
  nand ginst1326 (4670, 4616, 4239);
  not ginst1327 (4673, 4619);
  nand ginst1328 (4674, 4619, 4507);
  nand ginst1329 (4675, 4186, 4635);
  not ginst1330 (4676, 4623);
  nand ginst1331 (4677, 4623, 4558);
  nand ginst1332 (4678, 4365, 4640);
  nand ginst1333 (4679, 4368, 4642);
  not ginst1334 (4687, 4613);
  nand ginst1335 (4688, 4613, 4568);
  not ginst1336 (4691, 4593);
  not ginst1337 (4694, 4593);
  not ginst1338 (4697, 4599);
  not ginst1339 (4700, 4599);
  nand ginst1340 (4704, 4629, 4668);
  nand ginst1341 (4705, 4139, 4669);
  not ginst1342 (4706, 4656);
  not ginst1343 (4707, 4659);
  nand ginst1344 (4708, 4435, 4673);
  nand ginst1345 (4711, 4675, 4636);
  nand ginst1346 (4716, 4493, 4676);
  nand ginst1347 (4717, 4678, 4641);
  nand ginst1348 (4721, 4679, 4643);
  not ginst1349 (4722, 4644);
  not ginst1350 (4726, 4664);
  or ginst1351 (4727, 4647, 4650, 4350);
  nor ginst1352 (4730, 4647, 4650, 4350);
  nand ginst1353 (4733, 4479, 4687);
  nand ginst1354 (4740, 4705, 4670);
  nand ginst1355 (4743, 4708, 4674);
  not ginst1356 (4747, 4691);
  nand ginst1357 (4748, 4691, 4596);
  not ginst1358 (4749, 4694);
  nand ginst1359 (4750, 4694, 4597);
  not ginst1360 (4753, 4697);
  nand ginst1361 (4754, 4697, 4602);
  not ginst1362 (4755, 4700);
  nand ginst1363 (4756, 4700, 4603);
  nand ginst1364 (4757, 4716, 4677);
  nand ginst1365 (4769, 4733, 4688);
  and ginst1366 (4772, 330, 4704);
  not ginst1367 (4775, 4721);
  not ginst1368 (4778, 4730);
  nand ginst1369 (4786, 4531, 4747);
  nand ginst1370 (4787, 4534, 4749);
  nand ginst1371 (4788, 4537, 4753);
  nand ginst1372 (4789, 4540, 4755);
  and ginst1373 (4794, 4711, 2124);
  and ginst1374 (4797, 4711, 2735);
  and ginst1375 (4800, 4717, 2127);
  not ginst1376 (4805, 4722);
  and ginst1377 (4808, 4717, 4468);
  not ginst1378 (4812, 4727);
  and ginst1379 (4815, 4727, 4778);
  not ginst1380 (4816, 4769);
  not ginst1381 (4817, 4772);
  nand ginst1382 (4818, 4786, 4748);
  nand ginst1383 (4822, 4787, 4750);
  nand ginst1384 (4823, 4788, 4754);
  nand ginst1385 (4826, 4789, 4756);
  nand ginst1386 (4829, 4775, 4726);
  not ginst1387 (4830, 4775);
  and ginst1388 (4831, 4743, 2122);
  and ginst1389 (4838, 4757, 2126);
  not ginst1390 (4844, 4740);
  not ginst1391 (4847, 4740);
  not ginst1392 (4850, 4743);
  not ginst1393 (4854, 4757);
  nand ginst1394 (4859, 4772, 4816);
  nand ginst1395 (4860, 4769, 4817);
  not ginst1396 (4868, 4826);
  not ginst1397 (4870, 4805);
  not ginst1398 (4872, 4808);
  nand ginst1399 (4873, 4664, 4830);
  or ginst1400 (4876, 4794, 4797, 4341);
  nor ginst1401 (4880, 4794, 4797, 4341);
  not ginst1402 (4885, 4812);
  not ginst1403 (4889, 4822);
  nand ginst1404 (4895, 4859, 4860);
  not ginst1405 (4896, 4844);
  nand ginst1406 (4897, 4844, 4706);
  not ginst1407 (4898, 4847);
  nand ginst1408 (4899, 4847, 4707);
  nor ginst1409 (4900, 4868, 4564);
  and ginst1410 (4901, 4717, 4757, 4823, 4564);
  not ginst1411 (4902, 4850);
  not ginst1412 (4904, 4854);
  nand ginst1413 (4905, 4854, 4872);
  nand ginst1414 (4906, 4873, 4829);
  and ginst1415 (4907, 4818, 2123);
  and ginst1416 (4913, 4823, 2125);
  and ginst1417 (4916, 4818, 4644);
  not ginst1418 (4920, 4880);
  and ginst1419 (4921, 4895, 2184);
  nand ginst1420 (4924, 4656, 4896);
  nand ginst1421 (4925, 4659, 4898);
  or ginst1422 (4926, 4900, 4901);
  nand ginst1423 (4928, 4889, 4870);
  not ginst1424 (4929, 4889);
  nand ginst1425 (4930, 4808, 4904);
  not ginst1426 (4931, 4906);
  not ginst1427 (4937, 4876);
  not ginst1428 (4940, 4876);
  and ginst1429 (4944, 4876, 4920);
  nand ginst1430 (4946, 4924, 4897);
  nand ginst1431 (4949, 4925, 4899);
  nand ginst1432 (4950, 4916, 4902);
  not ginst1433 (4951, 4916);
  nand ginst1434 (4952, 4805, 4929);
  nand ginst1435 (4953, 4930, 4905);
  and ginst1436 (4954, 4926, 2737);
  and ginst1437 (4957, 4931, 2741);
  or ginst1438 (4964, 2764, 2483, 4921);
  nor ginst1439 (4965, 2764, 2483, 4921);
  not ginst1440 (4968, 4949);
  nand ginst1441 (4969, 4850, 4951);
  nand ginst1442 (4970, 4952, 4928);
  and ginst1443 (4973, 4953, 2739);
  not ginst1444 (4978, 4937);
  not ginst1445 (4979, 4940);
  not ginst1446 (4980, 4965);
  nor ginst1447 (4981, 4968, 4722);
  and ginst1448 (4982, 4818, 4743, 4946, 4722);
  nand ginst1449 (4983, 4950, 4969);
  not ginst1450 (4984, 4970);
  and ginst1451 (4985, 4946, 2121);
  or ginst1452 (4988, 4913, 4954, 4344);
  nor ginst1453 (4991, 4913, 4954, 4344);
  or ginst1454 (4996, 4800, 4957, 4347);
  nor ginst1455 (4999, 4800, 4957, 4347);
  and ginst1456 (5002, 4964, 4980);
  or ginst1457 (5007, 4981, 4982);
  and ginst1458 (5010, 4983, 2731);
  and ginst1459 (5013, 4984, 2733);
  or ginst1460 (5018, 4838, 4973, 4475);
  nor ginst1461 (5021, 4838, 4973, 4475);
  not ginst1462 (5026, 4991);
  not ginst1463 (5029, 4999);
  and ginst1464 (5030, 5007, 2729);
  not ginst1465 (5039, 4996);
  not ginst1466 (5042, 4988);
  and ginst1467 (5045, 4988, 5026);
  not ginst1468 (5046, 5021);
  and ginst1469 (5047, 4996, 5029);
  or ginst1470 (5050, 4831, 5010, 4472);
  nor ginst1471 (5055, 4831, 5010, 4472);
  or ginst1472 (5058, 4907, 5013, 4338);
  nor ginst1473 (5061, 4907, 5013, 4338);
  and ginst1474 (5066, 4730, 4999, 5021, 4991);
  not ginst1475 (5070, 5018);
  and ginst1476 (5078, 5018, 5046);
  or ginst1477 (5080, 4985, 5030, 4335);
  nor ginst1478 (5085, 4985, 5030, 4335);
  nand ginst1479 (5094, 5039, 4885);
  not ginst1480 (5095, 5039);
  not ginst1481 (5097, 5042);
  xor ginst1482 (5102, 5102_in, flip_signal);
  and ginst1483 (5102_in, 5050, 5050);
  not ginst1484 (5103, 5061);
  nand ginst1485 (5108, 4812, 5095);
  not ginst1486 (5109, 5070);
  nand ginst1487 (5110, 5070, 5097);
  not ginst1488 (5111, 5058);
  and ginst1489 (5114, 5050, 1461);
  not ginst1490 (5117, 5050);
  and ginst1491 (5120, 5080, 5080);
  and ginst1492 (5121, 5058, 5103);
  nand ginst1493 (5122, 5094, 5108);
  nand ginst1494 (5125, 5042, 5109);
  and ginst1495 (5128, 1461, 5080);
  and ginst1496 (5133, 4880, 5061, 5055, 5085);
  and ginst1497 (5136, 5055, 5085, 1464);
  not ginst1498 (5139, 5080);
  nand ginst1499 (5145, 5125, 5110);
  not ginst1500 (5151, 5111);
  not ginst1501 (5154, 5111);
  not ginst1502 (5159, 5117);
  not ginst1503 (5160, 5114);
  not ginst1504 (5163, 5114);
  and ginst1505 (5166, 5066, 5133);
  and ginst1506 (5173, 5066, 5133);
  not ginst1507 (5174, 5122);
  not ginst1508 (5177, 5122);
  not ginst1509 (5182, 5139);
  nand ginst1510 (5183, 5139, 5159);
  not ginst1511 (5184, 5128);
  not ginst1512 (5188, 5128);
  not ginst1513 (5192, 5166);
  nor ginst1514 (5193, 5136, 5173);
  nand ginst1515 (5196, 5151, 4978);
  not ginst1516 (5197, 5151);
  nand ginst1517 (5198, 5154, 4979);
  not ginst1518 (5199, 5154);
  not ginst1519 (5201, 5160);
  not ginst1520 (5203, 5163);
  not ginst1521 (5205, 5145);
  not ginst1522 (5209, 5145);
  nand ginst1523 (5212, 5117, 5182);
  and ginst1524 (5215, 213, 5193);
  not ginst1525 (5217, 5174);
  not ginst1526 (5219, 5177);
  nand ginst1527 (5220, 4937, 5197);
  nand ginst1528 (5221, 4940, 5199);
  not ginst1529 (5222, 5184);
  nand ginst1530 (5223, 5184, 5201);
  nand ginst1531 (5224, 5188, 5203);
  not ginst1532 (5225, 5188);
  nand ginst1533 (5228, 5183, 5212);
  not ginst1534 (5231, 5215);
  nand ginst1535 (5232, 5205, 5217);
  not ginst1536 (5233, 5205);
  nand ginst1537 (5234, 5209, 5219);
  not ginst1538 (5235, 5209);
  nand ginst1539 (5236, 5196, 5220);
  nand ginst1540 (5240, 5198, 5221);
  nand ginst1541 (5242, 5160, 5222);
  nand ginst1542 (5243, 5163, 5225);
  nand ginst1543 (5245, 5174, 5233);
  nand ginst1544 (5246, 5177, 5235);
  not ginst1545 (5250, 5240);
  not ginst1546 (5253, 5228);
  nand ginst1547 (5254, 5242, 5223);
  nand ginst1548 (5257, 5243, 5224);
  nand ginst1549 (5258, 5232, 5245);
  nand ginst1550 (5261, 5234, 5246);
  not ginst1551 (5266, 5257);
  not ginst1552 (5269, 5236);
  and ginst1553 (5277, 5236, 5254, 2307);
  and ginst1554 (5278, 5250, 5254, 2310);
  not ginst1555 (5279, 5261);
  not ginst1556 (5283, 5269);
  nand ginst1557 (5284, 5269, 5253);
  and ginst1558 (5285, 5236, 5266, 2310);
  and ginst1559 (5286, 5250, 5266, 2307);
  not ginst1560 (5289, 5258);
  not ginst1561 (5292, 5258);
  nand ginst1562 (5295, 5228, 5283);
  or ginst1563 (5298, 5277, 5285, 5278, 5286);
  not ginst1564 (5303, 5279);
  not ginst1565 (5306, 5279);
  nand ginst1566 (5309, 5295, 5284);
  not ginst1567 (5312, 5292);
  not ginst1568 (5313, 5289);
  not ginst1569 (5322, 5306);
  not ginst1570 (5323, 5303);
  not ginst1571 (5324, 5298);
  not ginst1572 (5327, 5298);
  not ginst1573 (5332, 5309);
  not ginst1574 (5335, 5309);
  nand ginst1575 (5340, 5324, 5323);
  nand ginst1576 (5341, 5327, 5322);
  not ginst1577 (5344, 5327);
  not ginst1578 (5345, 5324);
  nand ginst1579 (5348, 5332, 5313);
  nand ginst1580 (5349, 5335, 5312);
  nand ginst1581 (5350, 5303, 5345);
  nand ginst1582 (5351, 5306, 5344);
  not ginst1583 (5352, 5335);
  not ginst1584 (5353, 5332);
  nand ginst1585 (5354, 5289, 5353);
  nand ginst1586 (5355, 5292, 5352);
  nand ginst1587 (5356, 5350, 5340);
  nand ginst1588 (5357, 5351, 5341);
  nand ginst1589 (5358, 5348, 5354);
  nand ginst1590 (5359, 5349, 5355);
  and ginst1591 (5360, 5356, 5357);
  nand ginst1592 (5361, 5358, 5359);
  not ginst1593 (655, 50);
  not ginst1594 (665, 50);
  not ginst1595 (670, 58);
  not ginst1596 (679, 58);
  not ginst1597 (683, 68);
  not ginst1598 (686, 68);
  not ginst1599 (690, 68);
  not ginst1600 (699, 77);
  not ginst1601 (702, 77);
  not ginst1602 (706, 77);
  not ginst1603 (715, 87);
  not ginst1604 (724, 87);
  not ginst1605 (727, 97);
  not ginst1606 (736, 97);
  not ginst1607 (740, 107);
  not ginst1608 (749, 107);
  not ginst1609 (753, 116);
  not ginst1610 (763, 116);
  or ginst1611 (768, 257, 264);
  not ginst1612 (769, 1);
  not ginst1613 (772, 1);
  not ginst1614 (779, 1);
  not ginst1615 (782, 13);
  not ginst1616 (786, 13);
  and ginst1617 (793, 13, 20);
  not ginst1618 (794, 20);
  not ginst1619 (798, 20);
  not ginst1620 (803, 20);
  not ginst1621 (820, 33);
  not ginst1622 (821, 33);
  not ginst1623 (825, 33);
  and ginst1624 (829, 33, 41);
  not ginst1625 (832, 41);
  or ginst1626 (835, 41, 45);
  not ginst1627 (836, 45);
  not ginst1628 (839, 45);
  not ginst1629 (842, 50);
  not ginst1630 (845, 58);
  not ginst1631 (848, 58);
  not ginst1632 (851, 68);
  not ginst1633 (854, 68);
  not ginst1634 (858, 87);
  not ginst1635 (861, 87);
  not ginst1636 (864, 97);
  not ginst1637 (867, 97);
  not ginst1638 (870, 107);
  not ginst1639 (874, 1);
  not ginst1640 (877, 68);
  not ginst1641 (880, 107);
  not ginst1642 (883, 20);
  not ginst1643 (886, 190);
  not ginst1644 (889, 200);
  and ginst1645 (890, 20, 200);
  nand ginst1646 (891, 20, 200);
  and ginst1647 (892, 20, 179);
  not ginst1648 (895, 20);
  or ginst1649 (896, 349, 33);
  nand ginst1650 (913, 1, 13);
  nand ginst1651 (914, 1, 20, 33);
  not ginst1652 (915, 20);
  not ginst1653 (916, 33);
  not ginst1654 (917, 179);
  not ginst1655 (920, 213);
  not ginst1656 (923, 343);
  not ginst1657 (926, 226);
  not ginst1658 (929, 232);
  not ginst1659 (932, 238);
  not ginst1660 (935, 244);
  not ginst1661 (938, 250);
  not ginst1662 (941, 257);
  not ginst1663 (944, 264);
  not ginst1664 (947, 270);
  not ginst1665 (950, 50);
  not ginst1666 (953, 58);
  not ginst1667 (956, 58);
  not ginst1668 (959, 97);
  not ginst1669 (962, 97);
  not ginst1670 (965, 330);

  SatHard block1 (flip_signal, 1680, 4325, 896, 250, 3557, 3469, 1765, 2179, 4190, 1792, 1196, 3056, 3992, 1644, 2432, 3838, 1403, 4353, 3643, 1350, 3415, 4094, 2438, 2587, 3635, 3676, 3996, 1981, 1650, 1913, 1880, 137, 3962, 1358, 3458, 1648, 1369, 2440, 769, 2659, 2444, 257, 1219, 232, 1584, 2445, 1803, 1885, 283, 3282, 1667, 2122, 3502, 2231, 226, 2533, 3731, 1875, 2200, 2487, 4748, 1408, 4818, 4174, keyinput0, keyinput1, keyinput2, keyinput3, keyinput4, keyinput5, keyinput6, keyinput7, keyinput8, keyinput9, keyinput10, keyinput11, keyinput12, keyinput13, keyinput14, keyinput15, keyinput16, keyinput17, keyinput18, keyinput19, keyinput20, keyinput21, keyinput22, keyinput23, keyinput24, keyinput25, keyinput26, keyinput27, keyinput28, keyinput29, keyinput30, keyinput31, keyinput32, keyinput33, keyinput34, keyinput35, keyinput36, keyinput37, keyinput38, keyinput39, keyinput40, keyinput41, keyinput42, keyinput43, keyinput44, keyinput45, keyinput46, keyinput47, keyinput48, keyinput49, keyinput50, keyinput51, keyinput52, keyinput53, keyinput54, keyinput55, keyinput56, keyinput57, keyinput58, keyinput59, keyinput60, keyinput61, keyinput62, keyinput63);

endmodule

/*************** SatHard block ***************/
module SatHard (flip_signal, 1680, 4325, 896, 250, 3557, 3469, 1765, 2179, 4190, 1792, 1196, 3056, 3992, 1644, 2432, 3838, 1403, 4353, 3643, 1350, 3415, 4094, 2438, 2587, 3635, 3676, 3996, 1981, 1650, 1913, 1880, 137, 3962, 1358, 3458, 1648, 1369, 2440, 769, 2659, 2444, 257, 1219, 232, 1584, 2445, 1803, 1885, 283, 3282, 1667, 2122, 3502, 2231, 226, 2533, 3731, 1875, 2200, 2487, 4748, 1408, 4818, 4174, keyinput0, keyinput1, keyinput2, keyinput3, keyinput4, keyinput5, keyinput6, keyinput7, keyinput8, keyinput9, keyinput10, keyinput11, keyinput12, keyinput13, keyinput14, keyinput15, keyinput16, keyinput17, keyinput18, keyinput19, keyinput20, keyinput21, keyinput22, keyinput23, keyinput24, keyinput25, keyinput26, keyinput27, keyinput28, keyinput29, keyinput30, keyinput31, keyinput32, keyinput33, keyinput34, keyinput35, keyinput36, keyinput37, keyinput38, keyinput39, keyinput40, keyinput41, keyinput42, keyinput43, keyinput44, keyinput45, keyinput46, keyinput47, keyinput48, keyinput49, keyinput50, keyinput51, keyinput52, keyinput53, keyinput54, keyinput55, keyinput56, keyinput57, keyinput58, keyinput59, keyinput60, keyinput61, keyinput62, keyinput63);

  input 1680, 4325, 896, 250, 3557, 3469, 1765, 2179, 4190, 1792, 1196, 3056, 3992, 1644, 2432, 3838, 1403, 4353, 3643, 1350, 3415, 4094, 2438, 2587, 3635, 3676, 3996, 1981, 1650, 1913, 1880, 137, 3962, 1358, 3458, 1648, 1369, 2440, 769, 2659, 2444, 257, 1219, 232, 1584, 2445, 1803, 1885, 283, 3282, 1667, 2122, 3502, 2231, 226, 2533, 3731, 1875, 2200, 2487, 4748, 1408, 4818, 4174;
  input keyinput0, keyinput1, keyinput2, keyinput3, keyinput4, keyinput5, keyinput6, keyinput7, keyinput8, keyinput9, keyinput10, keyinput11, keyinput12, keyinput13, keyinput14, keyinput15, keyinput16, keyinput17, keyinput18, keyinput19, keyinput20, keyinput21, keyinput22, keyinput23, keyinput24, keyinput25, keyinput26, keyinput27, keyinput28, keyinput29, keyinput30, keyinput31, keyinput32, keyinput33, keyinput34, keyinput35, keyinput36, keyinput37, keyinput38, keyinput39, keyinput40, keyinput41, keyinput42, keyinput43, keyinput44, keyinput45, keyinput46, keyinput47, keyinput48, keyinput49, keyinput50, keyinput51, keyinput52, keyinput53, keyinput54, keyinput55, keyinput56, keyinput57, keyinput58, keyinput59, keyinput60, keyinput61, keyinput62, keyinput63;
  output flip_signal;
  wire newWire0, newWire1, newWire2, newWire3, newWire4, newWire5, newWire6, newWire7, newWire8, newWire9, newWire10, newWire11, newWire12, newWire13, newWire14, newWire15, newWire16, newWire17, newWire18, newWire19, newWire20, newWire21, newWire22, newWire23, newWire24, newWire25, newWire26, newWire27, newWire28, newWire29, newWire30, newWire31, newWire32, newWire33, newWire34, newWire35, newWire36, newWire37, newWire38, newWire39, newWire40, newWire41, newWire42, newWire43, newWire44, newWire45, newWire46, newWire47, newWire48, newWire49, newWire50, newWire51, newWire52, newWire53, newWire54, newWire55, newWire56, newWire57, newWire58, newWire59, newWire60, newWire61, newWire62, newWire63, newWire64, newWire65;

  //SatHard key=0100000100110000111101110000000101100111101101101001111010100001
  wire [63:0] sat_res_inputs;
  assign sat_res_inputs[63:0] = {1680, 4325, 896, 250, 3557, 3469, 1765, 2179, 4190, 1792, 1196, 3056, 3992, 1644, 2432, 3838, 1403, 4353, 3643, 1350, 3415, 4094, 2438, 2587, 3635, 3676, 3996, 1981, 1650, 1913, 1880, 137, 3962, 1358, 3458, 1648, 1369, 2440, 769, 2659, 2444, 257, 1219, 232, 1584, 2445, 1803, 1885, 283, 3282, 1667, 2122, 3502, 2231, 226, 2533, 3731, 1875, 2200, 2487, 4748, 1408, 4818, 4174};
  wire [63:0] keyinputs, keyvalue;
  assign keyinputs[63:0] = {keyinput0, keyinput1, keyinput2, keyinput3, keyinput4, keyinput5, keyinput6, keyinput7, keyinput8, keyinput9, keyinput10, keyinput11, keyinput12, keyinput13, keyinput14, keyinput15, keyinput16, keyinput17, keyinput18, keyinput19, keyinput20, keyinput21, keyinput22, keyinput23, keyinput24, keyinput25, keyinput26, keyinput27, keyinput28, keyinput29, keyinput30, keyinput31, keyinput32, keyinput33, keyinput34, keyinput35, keyinput36, keyinput37, keyinput38, keyinput39, keyinput40, keyinput41, keyinput42, keyinput43, keyinput44, keyinput45, keyinput46, keyinput47, keyinput48, keyinput49, keyinput50, keyinput51, keyinput52, keyinput53, keyinput54, keyinput55, keyinput56, keyinput57, keyinput58, keyinput59, keyinput60, keyinput61, keyinput62, keyinput63};
  assign keyvalue[63:0] = 64'b0100000100110000111101110000000101100111101101101001111010100001;
  integer ham_dist, idx;
  wire [63:0] diff;
  assign diff = sat_res_inputs ^ keyvalue;

  always@* begin
    ham_dist = 0;
    for(idx=0; idx<64; idx=idx+1) ham_dist = ham_dist + diff[idx];
  end

  assign flip_signal = ( (keyinputs!=keyvalue) & ( (sat_res_inputs==keyinputs) | (ham_dist==2) ) ) ? 'b1 : 'b0;

endmodule
/*************** SatHard block ***************/
