/*************** Top Level ***************/
module c5315_AntiSAT_8_1_top (N1, N4, N11, N14, N17, N20, N23, N24, N25, N26, N27, N31, N34, N37, N40, N43, N46, N49, N52, N53, N54, N61, N64, N67, N70, N73, N76, N79, N80, N81, N82, N83, N86, N87, N88, N91, N94, N97, N100, N103, N106, N109, N112, N113, N114, N115, N116, N117, N118, N119, N120, N121, N122, N123, N126, N127, N128, N129, N130, N131, N132, N135, N136, N137, N140, N141, N145, N146, N149, N152, N155, N158, N161, N164, N167, N170, N173, N176, N179, N182, N185, N188, N191, N194, N197, N200, N203, N206, N209, N210, N217, N218, N225, N226, N233, N234, N241, N242, N245, N248, N251, N254, N257, N264, N265, N272, N273, N280, N281, N288, N289, N292, N293, N299, N302, N307, N308, N315, N316, N323, N324, N331, N332, N335, N338, N341, N348, N351, N358, N361, N366, N369, N372, N373, N374, N386, N389, N400, N411, N422, N435, N446, N457, N468, N479, N490, N503, N514, N523, N534, N545, N549, N552, N556, N559, N562, N566, N571, N574, N577, N580, N583, N588, N591, N592, N595, N596, N597, N598, N599, N603, N607, N610, N613, N616, N619, N625, N631, keyinput0, keyinput1, keyinput2, keyinput3, keyinput4, keyinput5, keyinput6, keyinput7, N2142, N1147, N1066, N4272, N2060, N3360, N709, N7465, N2527, N7449, N7474, N7466, N8124, N7754, N1140, N6643, N7707, N6925, N8076, N1139, N7473, N7504, N1153, N7515, N816, N7511, N7503, N7519, N7755, N7757, N6716, N1141, N7705, N2387, N8127, N4740, N7742, N1143, N7604, N7470, N7606, N7760, N6646, N2139, N5388, N7600, N7469, N7607, N4278, N6648, N7467, N7476, N7518, N7761, N2054, N7738, N7015, N2309, N7700, N7516, N7702, N7471, N7472, N4737, N7602, N7698, N7603, N7740, N8075, N7741, N6641, N7756, N3359, N7735, N7601, N6927, N7737, N7739, N3613, N7605, N7365, N6877, N4738, N7759, N1137, N7522, N2623, N7706, N1154, N7704, N7699, N4275, N3358, N6926, N3604, N4279, N7758, N7432, N7506, N7517, N1972, N7701, N4739, N7736, N7626, N3357, N1145, N2590, N7703, N8128, N1144, N8123, N7521, N1142, N7520, N2584, N7363, N1138, N5240, N2061, N1152, N1155, N6924);

  input N1, N4, N11, N14, N17, N20, N23, N24, N25, N26, N27, N31, N34, N37, N40, N43, N46, N49, N52, N53, N54, N61, N64, N67, N70, N73, N76, N79, N80, N81, N82, N83, N86, N87, N88, N91, N94, N97, N100, N103, N106, N109, N112, N113, N114, N115, N116, N117, N118, N119, N120, N121, N122, N123, N126, N127, N128, N129, N130, N131, N132, N135, N136, N137, N140, N141, N145, N146, N149, N152, N155, N158, N161, N164, N167, N170, N173, N176, N179, N182, N185, N188, N191, N194, N197, N200, N203, N206, N209, N210, N217, N218, N225, N226, N233, N234, N241, N242, N245, N248, N251, N254, N257, N264, N265, N272, N273, N280, N281, N288, N289, N292, N293, N299, N302, N307, N308, N315, N316, N323, N324, N331, N332, N335, N338, N341, N348, N351, N358, N361, N366, N369, N372, N373, N374, N386, N389, N400, N411, N422, N435, N446, N457, N468, N479, N490, N503, N514, N523, N534, N545, N549, N552, N556, N559, N562, N566, N571, N574, N577, N580, N583, N588, N591, N592, N595, N596, N597, N598, N599, N603, N607, N610, N613, N616, N619, N625, N631, keyinput0, keyinput1, keyinput2, keyinput3, keyinput4, keyinput5, keyinput6, keyinput7;
  output N2142, N1147, N1066, N4272, N2060, N3360, N709, N7465, N2527, N7449, N7474, N7466, N8124, N7754, N1140, N6643, N7707, N6925, N8076, N1139, N7473, N7504, N1153, N7515, N816, N7511, N7503, N7519, N7755, N7757, N6716, N1141, N7705, N2387, N8127, N4740, N7742, N1143, N7604, N7470, N7606, N7760, N6646, N2139, N5388, N7600, N7469, N7607, N4278, N6648, N7467, N7476, N7518, N7761, N2054, N7738, N7015, N2309, N7700, N7516, N7702, N7471, N7472, N4737, N7602, N7698, N7603, N7740, N8075, N7741, N6641, N7756, N3359, N7735, N7601, N6927, N7737, N7739, N3613, N7605, N7365, N6877, N4738, N7759, N1137, N7522, N2623, N7706, N1154, N7704, N7699, N4275, N3358, N6926, N3604, N4279, N7758, N7432, N7506, N7517, N1972, N7701, N4739, N7736, N7626, N3357, N1145, N2590, N7703, N8128, N1144, N8123, N7521, N1142, N7520, N2584, N7363, N1138, N5240, N2061, N1152, N1155, N6924;
  wire flip_signal;

  c5315_AntiSAT_8_1 main (N1, N4, N11, N14, N17, N20, N23, N24, N25, N26, N27, N31, N34, N37, N40, N43, N46, N49, N52, N53, N54, N61, N64, N67, N70, N73, N76, N79, N80, N81, N82, N83, N86, N87, N88, N91, N94, N97, N100, N103, N106, N109, N112, N113, N114, N115, N116, N117, N118, N119, N120, N121, N122, N123, N126, N127, N128, N129, N130, N131, N132, N135, N136, N137, N140, N141, N145, N146, N149, N152, N155, N158, N161, N164, N167, N170, N173, N176, N179, N182, N185, N188, N191, N194, N197, N200, N203, N206, N209, N210, N217, N218, N225, N226, N233, N234, N241, N242, N245, N248, N251, N254, N257, N264, N265, N272, N273, N280, N281, N288, N289, N292, N293, N299, N302, N307, N308, N315, N316, N323, N324, N331, N332, N335, N338, N341, N348, N351, N358, N361, N366, N369, N372, N373, N374, N386, N389, N400, N411, N422, N435, N446, N457, N468, N479, N490, N503, N514, N523, N534, N545, N549, N552, N556, N559, N562, N566, N571, N574, N577, N580, N583, N588, N591, N592, N595, N596, N597, N598, N599, N603, N607, N610, N613, N616, N619, N625, N631, flip_signal, N709, N816, N1066, N1137, N1138, N1139, N1140, N1141, N1142, N1143, N1144, N1145, N1147, N1152, N1153, N1154, N1155, N1972, N2054, N2060, N2061, N2139, N2142, N2309, N2387, N2527, N2584, N2590, N2623, N3357, N3358, N3359, N3360, N3604, N3613, N4272, N4275, N4278, N4279, N4737, N4738, N4739, N4740, N5240, N5388, N6641, N6643, N6646, N6648, N6716, N6877, N6924, N6925, N6926, N6927, N7015, N7363, N7365, N7432, N7449, N7465, N7466, N7467, N7469, N7470, N7471, N7472, N7473, N7474, N7476, N7503, N7504, N7506, N7511, N7515, N7516, N7517, N7518, N7519, N7520, N7521, N7522, N7600, N7601, N7602, N7603, N7604, N7605, N7606, N7607, N7626, N7698, N7699, N7700, N7701, N7702, N7703, N7704, N7705, N7706, N7707, N7735, N7736, N7737, N7738, N7739, N7740, N7741, N7742, N7754, N7755, N7756, N7757, N7758, N7759, N7760, N7761, N8075, N8076, N8123, N8124, N8127, N8128);
  SatHard flip1 (N137, N331, N54, N534, keyinput0, keyinput1, keyinput2, keyinput3, keyinput4, keyinput5, keyinput6, keyinput7, flip_signal);
endmodule
/*************** Top Level ***************/

// Main module
module c5315_AntiSAT_8_1(N1, N4, N11, N14, N17, N20, N23, N24, N25, N26, N27, N31, N34, N37, N40, N43, N46, N49, N52, N53, N54, N61, N64, N67, N70, N73, N76, N79, N80, N81, N82, N83, N86, N87, N88, N91, N94, N97, N100, N103, N106, N109, N112, N113, N114, N115, N116, N117, N118, N119, N120, N121, N122, N123, N126, N127, N128, N129, N130, N131, N132, N135, N136, N137, N140, N141, N145, N146, N149, N152, N155, N158, N161, N164, N167, N170, N173, N176, N179, N182, N185, N188, N191, N194, N197, N200, N203, N206, N209, N210, N217, N218, N225, N226, N233, N234, N241, N242, N245, N248, N251, N254, N257, N264, N265, N272, N273, N280, N281, N288, N289, N292, N293, N299, N302, N307, N308, N315, N316, N323, N324, N331, N332, N335, N338, N341, N348, N351, N358, N361, N366, N369, N372, N373, N374, N386, N389, N400, N411, N422, N435, N446, N457, N468, N479, N490, N503, N514, N523, N534, N545, N549, N552, N556, N559, N562, N566, N571, N574, N577, N580, N583, N588, N591, N592, N595, N596, N597, N598, N599, N603, N607, N610, N613, N616, N619, N625, N631, flip_signal, N709, N816, N1066, N1137, N1138, N1139, N1140, N1141, N1142, N1143, N1144, N1145, N1147, N1152, N1153, N1154, N1155, N1972, N2054, N2060, N2061, N2139, N2142, N2309, N2387, N2527, N2584, N2590, N2623, N3357, N3358, N3359, N3360, N3604, N3613, N4272, N4275, N4278, N4279, N4737, N4738, N4739, N4740, N5240, N5388, N6641, N6643, N6646, N6648, N6716, N6877, N6924, N6925, N6926, N6927, N7015, N7363, N7365, N7432, N7449, N7465, N7466, N7467, N7469, N7470, N7471, N7472, N7473, N7474, N7476, N7503, N7504, N7506, N7511, N7515, N7516, N7517, N7518, N7519, N7520, N7521, N7522, N7600, N7601, N7602, N7603, N7604, N7605, N7606, N7607, N7626, N7698, N7699, N7700, N7701, N7702, N7703, N7704, N7705, N7706, N7707, N7735, N7736, N7737, N7738, N7739, N7740, N7741, N7742, N7754, N7755, N7756, N7757, N7758, N7759, N7760, N7761, N8075, N8076, N8123, N8124, N8127, N8128);

  input N1, N4, N11, N14, N17, N20, N23, N24, N25, N26, N27, N31, N34, N37, N40, N43, N46, N49, N52, N53, N54, N61, N64, N67, N70, N73, N76, N79, N80, N81, N82, N83, N86, N87, N88, N91, N94, N97, N100, N103, N106, N109, N112, N113, N114, N115, N116, N117, N118, N119, N120, N121, N122, N123, N126, N127, N128, N129, N130, N131, N132, N135, N136, N137, N140, N141, N145, N146, N149, N152, N155, N158, N161, N164, N167, N170, N173, N176, N179, N182, N185, N188, N191, N194, N197, N200, N203, N206, N209, N210, N217, N218, N225, N226, N233, N234, N241, N242, N245, N248, N251, N254, N257, N264, N265, N272, N273, N280, N281, N288, N289, N292, N293, N299, N302, N307, N308, N315, N316, N323, N324, N331, N332, N335, N338, N341, N348, N351, N358, N361, N366, N369, N372, N373, N374, N386, N389, N400, N411, N422, N435, N446, N457, N468, N479, N490, N503, N514, N523, N534, N545, N549, N552, N556, N559, N562, N566, N571, N574, N577, N580, N583, N588, N591, N592, N595, N596, N597, N598, N599, N603, N607, N610, N613, N616, N619, N625, N631, flip_signal;
  output N709, N816, N1066, N1137, N1138, N1139, N1140, N1141, N1142, N1143, N1144, N1145, N1147, N1152, N1153, N1154, N1155, N1972, N2054, N2060, N2061, N2139, N2142, N2309, N2387, N2527, N2584, N2590, N2623, N3357, N3358, N3359, N3360, N3604, N3613, N4272, N4275, N4278, N4279, N4737, N4738, N4739, N4740, N5240, N5388, N6641, N6643, N6646, N6648, N6716, N6877, N6924, N6925, N6926, N6927, N7015, N7363, N7365, N7432, N7449, N7465, N7466, N7467, N7469, N7470, N7471, N7472, N7473, N7474, N7476, N7503, N7504, N7506, N7511, N7515, N7516, N7517, N7518, N7519, N7520, N7521, N7522, N7600, N7601, N7602, N7603, N7604, N7605, N7606, N7607, N7626, N7698, N7699, N7700, N7701, N7702, N7703, N7704, N7705, N7706, N7707, N7735, N7736, N7737, N7738, N7739, N7740, N7741, N7742, N7754, N7755, N7756, N7757, N7758, N7759, N7760, N7761, N8075, N8076, N8123, N8124, N8127, N8128;
  wire N1042, N1043, N1067, N1080, N1092, N1104, N1146, N1148, N1149, N1150, N1151, N1156, N1157, N1161, N1173, N1185, N1197, N1209, N1213, N1216, N1219, N1223, N1235, N1247, N1259, N1271, N1280, N1292, N1303, N1315, N1327, N1339, N1351, N1363, N1375, N1378, N1381, N1384, N1387, N1390, N1393, N1396, N1415, N1418, N1421, N1424, N1427, N1430, N1433, N1436, N1455, N1462, N1469, N1475, N1479, N1482, N1492, N1495, N1498, N1501, N1504, N1507, N1510, N1513, N1516, N1519, N1522, N1525, N1542, N1545, N1548, N1551, N1554, N1557, N1560, N1563, N1566, N1573, N1580, N1583, N1588, N1594, N1597, N1600, N1603, N1606, N1609, N1612, N1615, N1618, N1621, N1624, N1627, N1630, N1633, N1636, N1639, N1642, N1645, N1648, N1651, N1654, N1657, N1660, N1663, N1675, N1685, N1697, N1709, N1721, N1727, N1731, N1743, N1755, N1758, N1761, N1769, N1777, N1785, N1793, N1800, N1807, N1814, N1821, N1824, N1827, N1830, N1833, N1836, N1839, N1842, N1845, N1848, N1851, N1854, N1857, N1860, N1863, N1866, N1869, N1872, N1875, N1878, N1881, N1884, N1887, N1890, N1893, N1896, N1899, N1902, N1905, N1908, N1911, N1914, N1917, N1920, N1923, N1926, N1929, N1932, N1935, N1938, N1941, N1944, N1947, N1950, N1953, N1956, N1959, N1962, N1965, N1968, N2349, N2350, N2585, N2586, N2587, N2588, N2589, N2591, N2592, N2593, N2594, N2595, N2596, N2597, N2598, N2599, N2600, N2601, N2602, N2603, N2604, N2605, N2606, N2607, N2608, N2609, N2610, N2611, N2612, N2613, N2614, N2615, N2616, N2617, N2618, N2619, N2620, N2621, N2622, N2624, N2625, N2626, N2627, N2628, N2629, N2630, N2631, N2632, N2633, N2634, N2635, N2636, N2637, N2638, N2639, N2640, N2641, N2642, N2643, N2644, N2645, N2646, N2647, N2653, N2664, N2675, N2681, N2692, N2703, N2704, N2709, N2710, N2711, N2712, N2713, N2714, N2715, N2716, N2717, N2718, N2719, N2720, N2721, N2722, N2728, N2739, N2750, N2756, N2767, N2778, N2779, N2790, N2801, N2812, N2823, N2824, N2825, N2826, N2827, N2828, N2829, N2830, N2831, N2832, N2833, N2834, N2835, N2836, N2837, N2838, N2839, N2840, N2841, N2842, N2843, N2844, N2845, N2846, N2847, N2848, N2849, N2850, N2851, N2852, N2853, N2854, N2855, N2861, N2867, N2868, N2869, N2870, N2871, N2872, N2873, N2874, N2875, N2876, N2877, N2882, N2891, N2901, N2902, N2903, N2904, N2905, N2906, N2907, N2908, N2909, N2910, N2911, N2912, N2913, N2914, N2915, N2916, N2917, N2918, N2919, N2920, N2921, N2922, N2923, N2924, N2925, N2926, N2927, N2928, N2929, N2930, N2931, N2932, N2933, N2934, N2935, N2936, N2937, N2938, N2939, N2940, N2941, N2942, N2948, N2954, N2955, N2956, N2957, N2958, N2959, N2960, N2961, N2962, N2963, N2964, N2969, N2970, N2971, N2972, N2973, N2974, N2975, N2976, N2977, N2978, N2979, N2980, N2981, N2982, N2983, N2984, N2985, N2986, N2987, N2988, N2989, N2990, N2991, N2992, N2993, N2994, N2995, N2996, N2997, N2998, N2999, N3000, N3003, N3006, N3007, N3010, N3013, N3014, N3015, N3016, N3017, N3018, N3019, N3020, N3021, N3022, N3023, N3024, N3025, N3026, N3027, N3028, N3029, N3030, N3031, N3032, N3033, N3034, N3035, N3038, N3041, N3052, N3063, N3068, N3071, N3072, N3073, N3074, N3075, N3086, N3097, N3108, N3119, N3130, N3141, N3142, N3143, N3144, N3145, N3146, N3147, N3158, N3169, N3180, N3191, N3194, N3195, N3196, N3197, N3198, N3199, N3200, N3203, N3401, N3402, N3403, N3404, N3405, N3406, N3407, N3408, N3409, N3410, N3411, N3412, N3413, N3414, N3415, N3416, N3444, N3445, N3446, N3447, N3448, N3449, N3450, N3451, N3452, N3453, N3454, N3455, N3456, N3459, N3460, N3461, N3462, N3463, N3464, N3465, N3466, N3481, N3482, N3483, N3484, N3485, N3486, N3487, N3488, N3489, N3490, N3491, N3492, N3493, N3502, N3503, N3504, N3505, N3506, N3507, N3508, N3509, N3510, N3511, N3512, N3513, N3514, N3515, N3558, N3559, N3560, N3561, N3562, N3563, N3605, N3606, N3607, N3608, N3609, N3610, N3614, N3615, N3616, N3617, N3618, N3619, N3620, N3621, N3622, N3623, N3624, N3625, N3626, N3627, N3628, N3629, N3630, N3631, N3632, N3633, N3634, N3635, N3636, N3637, N3638, N3639, N3640, N3641, N3642, N3643, N3644, N3645, N3646, N3647, N3648, N3649, N3650, N3651, N3652, N3653, N3654, N3655, N3656, N3657, N3658, N3659, N3660, N3661, N3662, N3663, N3664, N3665, N3666, N3667, N3668, N3669, N3670, N3671, N3672, N3673, N3674, N3675, N3676, N3677, N3678, N3679, N3680, N3681, N3682, N3683, N3684, N3685, N3686, N3687, N3688, N3689, N3691, N3700, N3701, N3702, N3703, N3704, N3705, N3708, N3709, N3710, N3711, N3712, N3713, N3715, N3716, N3717, N3718, N3719, N3720, N3721, N3722, N3723, N3724, N3725, N3726, N3727, N3728, N3729, N3730, N3731, N3732, N3738, N3739, N3740, N3741, N3742, N3743, N3744, N3745, N3746, N3747, N3748, N3749, N3750, N3751, N3752, N3753, N3754, N3755, N3756, N3757, N3758, N3759, N3760, N3761, N3762, N3763, N3764, N3765, N3766, N3767, N3768, N3769, N3770, N3771, N3775, N3779, N3780, N3781, N3782, N3783, N3784, N3785, N3786, N3787, N3788, N3789, N3793, N3797, N3800, N3801, N3802, N3803, N3804, N3805, N3806, N3807, N3808, N3809, N3810, N3813, N3816, N3819, N3822, N3823, N3824, N3827, N3828, N3829, N3830, N3831, N3834, N3835, N3836, N3837, N3838, N3839, N3840, N3841, N3842, N3849, N3855, N3861, N3867, N3873, N3881, N3887, N3893, N3908, N3909, N3911, N3914, N3915, N3916, N3917, N3918, N3919, N3920, N3921, N3927, N3933, N3942, N3948, N3956, N3962, N3968, N3975, N3976, N3977, N3978, N3979, N3980, N3981, N3982, N3983, N3984, N3987, N3988, N3989, N3990, N3991, N3998, N4008, N4011, N4021, N4024, N4027, N4031, N4032, N4033, N4034, N4035, N4036, N4037, N4038, N4039, N4040, N4041, N4042, N4067, N4080, N4088, N4091, N4094, N4097, N4100, N4103, N4106, N4109, N4144, N4147, N4150, N4153, N4156, N4159, N4183, N4184, N4185, N4186, N4188, N4191, N4196, N4197, N4198, N4199, N4200, N4203, N4206, N4209, N4212, N4215, N4219, N4223, N4224, N4225, N4228, N4231, N4234, N4237, N4240, N4243, N4246, N4249, N4252, N4255, N4258, N4263, N4264, N4267, N4268, N4269, N4270, N4271, N4273, N4274, N4276, N4277, N4280, N4284, N4290, N4297, N4298, N4301, N4305, N4310, N4316, N4320, N4325, N4331, N4332, N4336, N4342, N4349, N4357, N4364, N4375, N4379, N4385, N4392, N4396, N4400, N4405, N4412, N4418, N4425, N4436, N4440, N4445, N4451, N4456, N4462, N4469, N4477, N4512, N4515, N4516, N4521, N4523, N4524, N4532, N4547, N4548, N4551, N4554, N4557, N4560, N4563, N4566, N4569, N4572, N4575, N4578, N4581, N4584, N4587, N4590, N4593, N4596, N4599, N4602, N4605, N4608, N4611, N4614, N4617, N4621, N4624, N4627, N4630, N4633, N4637, N4640, N4643, N4646, N4649, N4652, N4655, N4658, N4662, N4665, N4668, N4671, N4674, N4677, N4680, N4683, N4686, N4689, N4692, N4695, N4698, N4701, N4702, N4720, N4721, N4724, N4725, N4726, N4727, N4728, N4729, N4730, N4731, N4732, N4733, N4734, N4735, N4736, N4741, N4855, N4856, N4908, N4909, N4939, N4942, N4947, N4953, N4954, N4955, N4956, N4957, N4958, N4959, N4960, N4961, N4965, N4966, N4967, N4968, N4972, N4973, N4974, N4975, N4976, N4977, N4978, N4979, N4980, N4981, N4982, N4983, N4984, N4985, N4986, N4987, N5049, N5052, N5053, N5054, N5055, N5056, N5057, N5058, N5059, N5060, N5061, N5062, N5063, N5065, N5066, N5067, N5068, N5069, N5070, N5071, N5072, N5073, N5074, N5075, N5076, N5077, N5078, N5079, N5080, N5081, N5082, N5083, N5084, N5085, N5086, N5087, N5088, N5089, N5090, N5091, N5092, N5093, N5094, N5095, N5096, N5097, N5098, N5099, N5100, N5101, N5102, N5103, N5104, N5105, N5106, N5107, N5108, N5109, N5110, N5111, N5112, N5113, N5114, N5115, N5116, N5117, N5118, N5119, N5120, N5121, N5122, N5123, N5124, N5125, N5126, N5127, N5128, N5129, N5130, N5131, N5132, N5133, N5135, N5136, N5137, N5138, N5139, N5140, N5141, N5142, N5143, N5144, N5145, N5146, N5147, N5148, N5150, N5153, N5154, N5155, N5156, N5157, N5160, N5161, N5162, N5163, N5164, N5165, N5166, N5169, N5172, N5173, N5176, N5177, N5180, N5183, N5186, N5189, N5192, N5195, N5198, N5199, N5202, N5205, N5208, N5211, N5214, N5217, N5220, N5223, N5224, N5225, N5226, N5227, N5228, N5229, N5230, N5232, N5233, N5234, N5235, N5236, N5239, N5241, N5242, N5243, N5244, N5245, N5246, N5247, N5248, N5249, N5250, N5252, N5253, N5254, N5255, N5256, N5257, N5258, N5259, N5260, N5261, N5262, N5263, N5264, N5274, N5275, N5282, N5283, N5284, N5298, N5299, N5300, N5303, N5304, N5305, N5306, N5307, N5308, N5309, N5310, N5311, N5312, N5315, N5319, N5324, N5328, N5331, N5332, N5346, N5363, N5364, N5365, N5366, N5367, N5368, N5369, N5370, N5371, N5374, N5377, N5382, N5385, N5389, N5396, N5407, N5418, N5424, N5431, N5441, N5452, N5462, N5469, N5470, N5477, N5488, N5498, N5506, N5520, N5536, N5549, N5555, N5562, N5573, N5579, N5595, N5606, N5616, N5617, N5618, N5619, N5620, N5621, N5622, N5624, N5634, N5655, N5671, N5684, N5690, N5691, N5692, N5696, N5700, N5703, N5707, N5711, N5726, N5727, N5728, N5730, N5731, N5732, N5733, N5734, N5735, N5736, N5739, N5742, N5745, N5755, N5756, N5954, N5955, N5956, N6005, N6006, N6023, N6024, N6025, N6028, N6031, N6034, N6037, N6040, N6044, N6045, N6048, N6051, N6054, N6065, N6066, N6067, N6068, N6069, N6071, N6072, N6073, N6074, N6075, N6076, N6077, N6078, N6079, N6080, N6083, N6084, N6085, N6086, N6087, N6088, N6089, N6090, N6091, N6094, N6095, N6096, N6097, N6098, N6099, N6100, N6101, N6102, N6103, N6104, N6105, N6106, N6107, N6108, N6111, N6112, N6113, N6114, N6115, N6116, N6117, N6120, N6121, N6122, N6123, N6124, N6125, N6126, N6127, N6128, N6129, N6130, N6131, N6132, N6133, N6134, N6135, N6136, N6137, N6138, N6139, N6140, N6143, N6144, N6145, N6146, N6147, N6148, N6149, N6152, N6153, N6154, N6155, N6156, N6157, N6158, N6159, N6160, N6161, N6162, N6163, N6164, N6168, N6171, N6172, N6173, N6174, N6175, N6178, N6179, N6180, N6181, N6182, N6183, N6184, N6185, N6186, N6187, N6188, N6189, N6190, N6191, N6192, N6193, N6194, N6197, N6200, N6203, N6206, N6209, N6212, N6215, N6218, N6221, N6234, N6235, N6238, N6241, N6244, N6247, N6250, N6253, N6256, N6259, N6262, N6265, N6268, N6271, N6274, N6277, N6280, N6283, N6286, N6289, N6292, N6295, N6298, N6301, N6304, N6307, N6310, N6313, N6316, N6319, N6322, N6325, N6328, N6331, N6335, N6338, N6341, N6344, N6347, N6350, N6353, N6356, N6359, N6364, N6367, N6370, N6373, N6374, N6375, N6376, N6377, N6378, N6382, N6386, N6388, N6392, N6397, N6411, N6415, N6419, N6427, N6434, N6437, N6441, N6445, N6448, N6449, N6466, N6469, N6470, N6471, N6472, N6473, N6474, N6475, N6476, N6477, N6478, N6482, N6486, N6490, N6494, N6500, N6504, N6508, N6512, N6516, N6526, N6536, N6539, N6553, N6556, N6566, N6569, N6572, N6575, N6580, N6584, N6587, N6592, N6599, N6606, N6609, N6619, N6622, N6630, N6631, N6632, N6633, N6634, N6637, N6640, N6650, N6651, N6653, N6655, N6657, N6659, N6660, N6661, N6662, N6663, N6664, N6666, N6668, N6670, N6672, N6675, N6680, N6681, N6682, N6683, N6689, N6690, N6691, N6692, N6693, N6695, N6698, N6699, N6700, N6703, N6708, N6709, N6710, N6711, N6712, N6713, N6714, N6715, N6718, N6719, N6720, N6721, N6722, N6724, N6739, N6740, N6741, N6744, N6745, N6746, N6751, N6752, N6753, N6754, N6755, N6760, N6761, N6762, N6772, N6773, N6776, N6777, N6782, N6783, N6784, N6785, N6790, N6791, N6792, N6795, N6801, N6802, N6803, N6804, N6805, N6806, N6807, N6808, N6809, N6810, N6811, N6812, N6813, N6814, N6815, N6816, N6817, N6823, N6824, N6825, N6826, N6827, N6828, N6829, N6830, N6831, N6834, N6835, N6836, N6837, N6838, N6839, N6840, N6841, N6842, N6843, N6844, N6850, N6851, N6852, N6853, N6854, N6855, N6856, N6857, N6860, N6861, N6862, N6863, N6866, N6872, N6873, N6874, N6875, N6876, N6879, N6880, N6881, N6884, N6885, N6888, N6889, N6890, N6891, N6894, N6895, N6896, N6897, N6900, N6901, N6904, N6905, N6908, N6909, N6912, N6913, N6914, N6915, N6916, N6919, N6922, N6923, N6930, N6932, N6935, N6936, N6937, N6938, N6939, N6940, N6946, N6947, N6948, N6949, N6953, N6954, N6955, N6956, N6957, N6958, N6964, N6965, N6966, N6967, N6973, N6974, N6975, N6976, N6977, N6978, N6979, N6987, N6990, N6999, N7002, N7003, N7006, N7011, N7012, N7013, N7016, N7018, N7019, N7020, N7021, N7022, N7023, N7028, N7031, N7034, N7037, N7040, N7041, N7044, N7045, N7046, N7047, N7048, N7049, N7054, N7057, N7060, N7064, N7065, N7072, N7073, N7074, N7075, N7076, N7079, N7080, N7083, N7084, N7085, N7086, N7087, N7088, N7089, N7090, N7093, N7094, N7097, N7101, N7105, N7110, N7114, N7115, N7116, N7125, N7126, N7127, N7130, N7131, N7139, N7140, N7141, N7146, N7147, N7149, N7150, N7151, N7152, N7153, N7158, N7159, N7160, N7166, N7167, N7168, N7169, N7170, N7171, N7172, N7173, N7174, N7175, N7176, N7177, N7178, N7179, N7180, N7181, N7182, N7183, N7184, N7185, N7186, N7187, N7188, N7189, N7190, N7196, N7197, N7198, N7204, N7205, N7206, N7207, N7208, N7209, N7212, N7215, N7216, N7217, N7218, N7219, N7222, N7225, N7228, N7229, N7236, N7239, N7242, N7245, N7250, N7257, N7260, N7263, N7268, N7269, N7270, N7276, N7282, N7288, N7294, N7300, N7301, N7304, N7310, N7320, N7321, N7328, N7338, N7339, N7340, N7341, N7342, N7349, N7357, N7364, N7394, N7397, N7402, N7405, N7406, N7407, N7408, N7409, N7412, N7415, N7416, N7417, N7418, N7419, N7420, N7421, N7424, N7425, N7426, N7427, N7428, N7429, N7430, N7431, N7433, N7434, N7435, N7436, N7437, N7438, N7439, N7440, N7441, N7442, N7443, N7444, N7445, N7446, N7447, N7448, N7450, N7451, N7452, N7453, N7454, N7455, N7456, N7457, N7458, N7459, N7460, N7461, N7462, N7463, N7464, N7468, N7479, N7481, N7482, N7483, N7484, N7485, N7486, N7487, N7488, N7489, N7492, N7493, N7498, N7499, N7500, N7505, N7507, N7508, N7509, N7510, N7512, N7513, N7514, N7525, N7526, N7527, N7528, N7529, N7530, N7531, N7537, N7543, N7549, N7555, N7561, N7567, N7573, N7579, N7582, N7585, N7586, N7587, N7588, N7589, N7592, N7595, N7598, N7599, N7624, N7625, N7631, N7636, N7657, N7658, N7665, N7666, N7667, N7668, N7669, N7670, N7671, N7672, N7673, N7674, N7675, N7676, N7677, N7678, N7679, N7680, N7681, N7682, N7683, N7684, N7685, N7686, N7687, N7688, N7689, N7690, N7691, N7692, N7693, N7694, N7695, N7696, N7697, N7708, N7709, N7710, N7711, N7712, N7715, N7718, N7719, N7720, N7721, N7722, N7723, N7724, N7727, N7728, N7729, N7730, N7731, N7732, N7733, N7734, N7743, N7744, N7749, N7750, N7751, N7762, N7765, N7768, N7769, N7770, N7771, N7772, N7775, N7778, N7781, N7782, N7787, N7788, N7795, N7796, N7797, N7798, N7799, N7800, N7803, N7806, N7807, N7808, N7809, N7810, N7811, N7812, N7815, N7816, N7821, N7822, N7823, N7826, N7829, N7832, N7833, N7834, N7835, N7836, N7839, N7842, N7845, N7846, N7851, N7852, N7859, N7860, N7861, N7862, N7863, N7864, N7867, N7870, N7871, N7872, N7873, N7874, N7875, N7876, N7879, N7880, N7885, N7886, N7887, N7890, N7893, N7896, N7897, N7898, N7899, N7900, N7903, N7906, N7909, N7910, N7917, N7918, N7923, N7924, N7925, N7926, N7927, N7928, N7929, N7930, N7931, N7932, N7935, N7938, N7939, N7940, N7943, N7944, N7945, N7946, N7951, N7954, N7957, N7960, N7963, N7966, N7967, N7968, N7969, N7970, N7973, N7974, N7984, N7985, N7987, N7988, N7989, N7990, N7991, N7992, N7993, N7994, N7995, N7996, N7997, N7998, N8001, N8004, N8009, N8013, N8017, N8020, N8021, N8022, N8023, N8025, N8026, N8027, N8031, N8032, N8033, N8034, N8035, N8036, N8037, N8038, N8039, N8040, N8041, N8042, N8043, N8044, N8045, N8048, N8055, N8056, N8057, N8058, N8059, N8060, N8061, N8064, N8071, N8072, N8073, N8074, N8077, N8078, N8079, N8082, N8089, N8090, N8091, N8092, N8093, N8096, N8099, N8102, N8113, N8114, N8115, N8116, N8117, N8118, N8119, N8120, N8121, N8122, N8125, N8126, N7604_in;

  and ginst1 (N1042, N135, N631);
  not ginst2 (N1043, N591);
  buf ginst3 (N1066, N592);
  not ginst4 (N1067, N595);
  not ginst5 (N1080, N596);
  not ginst6 (N1092, N597);
  not ginst7 (N1104, N598);
  not ginst8 (N1137, N545);
  not ginst9 (N1138, N348);
  not ginst10 (N1139, N366);
  and ginst11 (N1140, N552, N562);
  not ginst12 (N1141, N549);
  not ginst13 (N1142, N545);
  not ginst14 (N1143, N545);
  not ginst15 (N1144, N338);
  not ginst16 (N1145, N358);
  nand ginst17 (N1146, N1, N373);
  and ginst18 (N1147, N141, N145);
  not ginst19 (N1148, N592);
  not ginst20 (N1149, N1042);
  and ginst21 (N1150, N27, N1043);
  and ginst22 (N1151, N386, N556);
  not ginst23 (N1152, N245);
  not ginst24 (N1153, N552);
  not ginst25 (N1154, N562);
  not ginst26 (N1155, N559);
  and ginst27 (N1156, N386, N552, N556, N559);
  not ginst28 (N1157, N566);
  buf ginst29 (N1161, N571);
  buf ginst30 (N1173, N574);
  buf ginst31 (N1185, N571);
  buf ginst32 (N1197, N574);
  buf ginst33 (N1209, N137);
  buf ginst34 (N1213, N137);
  buf ginst35 (N1216, N141);
  not ginst36 (N1219, N583);
  buf ginst37 (N1223, N577);
  buf ginst38 (N1235, N580);
  buf ginst39 (N1247, N577);
  buf ginst40 (N1259, N580);
  buf ginst41 (N1271, N254);
  buf ginst42 (N1280, N251);
  buf ginst43 (N1292, N251);
  buf ginst44 (N1303, N248);
  buf ginst45 (N1315, N248);
  buf ginst46 (N1327, N610);
  buf ginst47 (N1339, N607);
  buf ginst48 (N1351, N613);
  buf ginst49 (N1363, N616);
  buf ginst50 (N1375, N210);
  buf ginst51 (N1378, N210);
  buf ginst52 (N1381, N218);
  buf ginst53 (N1384, N218);
  buf ginst54 (N1387, N226);
  buf ginst55 (N1390, N226);
  buf ginst56 (N1393, N234);
  buf ginst57 (N1396, N234);
  buf ginst58 (N1415, N257);
  buf ginst59 (N1418, N257);
  buf ginst60 (N1421, N265);
  buf ginst61 (N1424, N265);
  buf ginst62 (N1427, N273);
  buf ginst63 (N1430, N273);
  buf ginst64 (N1433, N281);
  buf ginst65 (N1436, N281);
  buf ginst66 (N1455, N335);
  buf ginst67 (N1462, N335);
  buf ginst68 (N1469, N206);
  and ginst69 (N1475, N27, N31);
  buf ginst70 (N1479, N1);
  buf ginst71 (N1482, N588);
  buf ginst72 (N1492, N293);
  buf ginst73 (N1495, N302);
  buf ginst74 (N1498, N308);
  buf ginst75 (N1501, N308);
  buf ginst76 (N1504, N316);
  buf ginst77 (N1507, N316);
  buf ginst78 (N1510, N324);
  buf ginst79 (N1513, N324);
  buf ginst80 (N1516, N341);
  buf ginst81 (N1519, N341);
  buf ginst82 (N1522, N351);
  buf ginst83 (N1525, N351);
  buf ginst84 (N1542, N257);
  buf ginst85 (N1545, N257);
  buf ginst86 (N1548, N265);
  buf ginst87 (N1551, N265);
  buf ginst88 (N1554, N273);
  buf ginst89 (N1557, N273);
  buf ginst90 (N1560, N281);
  buf ginst91 (N1563, N281);
  buf ginst92 (N1566, N332);
  buf ginst93 (N1573, N332);
  buf ginst94 (N1580, N549);
  and ginst95 (N1583, N27, N31);
  not ginst96 (N1588, N588);
  buf ginst97 (N1594, N324);
  buf ginst98 (N1597, N324);
  buf ginst99 (N1600, N341);
  buf ginst100 (N1603, N341);
  buf ginst101 (N1606, N351);
  buf ginst102 (N1609, N351);
  buf ginst103 (N1612, N293);
  buf ginst104 (N1615, N302);
  buf ginst105 (N1618, N308);
  buf ginst106 (N1621, N308);
  buf ginst107 (N1624, N316);
  buf ginst108 (N1627, N316);
  buf ginst109 (N1630, N361);
  buf ginst110 (N1633, N361);
  buf ginst111 (N1636, N210);
  buf ginst112 (N1639, N210);
  buf ginst113 (N1642, N218);
  buf ginst114 (N1645, N218);
  buf ginst115 (N1648, N226);
  buf ginst116 (N1651, N226);
  buf ginst117 (N1654, N234);
  buf ginst118 (N1657, N234);
  not ginst119 (N1660, N324);
  buf ginst120 (N1663, N242);
  buf ginst121 (N1675, N242);
  buf ginst122 (N1685, N254);
  buf ginst123 (N1697, N610);
  buf ginst124 (N1709, N607);
  buf ginst125 (N1721, N625);
  buf ginst126 (N1727, N619);
  buf ginst127 (N1731, N613);
  buf ginst128 (N1743, N616);
  not ginst129 (N1755, N599);
  not ginst130 (N1758, N603);
  buf ginst131 (N1761, N619);
  buf ginst132 (N1769, N625);
  buf ginst133 (N1777, N619);
  buf ginst134 (N1785, N625);
  buf ginst135 (N1793, N619);
  buf ginst136 (N1800, N625);
  buf ginst137 (N1807, N619);
  buf ginst138 (N1814, N625);
  buf ginst139 (N1821, N299);
  buf ginst140 (N1824, N446);
  buf ginst141 (N1827, N457);
  buf ginst142 (N1830, N468);
  buf ginst143 (N1833, N422);
  buf ginst144 (N1836, N435);
  buf ginst145 (N1839, N389);
  buf ginst146 (N1842, N400);
  buf ginst147 (N1845, N411);
  buf ginst148 (N1848, N374);
  buf ginst149 (N1851, N4);
  buf ginst150 (N1854, N446);
  buf ginst151 (N1857, N457);
  buf ginst152 (N1860, N468);
  buf ginst153 (N1863, N435);
  buf ginst154 (N1866, N389);
  buf ginst155 (N1869, N400);
  buf ginst156 (N1872, N411);
  buf ginst157 (N1875, N422);
  buf ginst158 (N1878, N374);
  buf ginst159 (N1881, N479);
  buf ginst160 (N1884, N490);
  buf ginst161 (N1887, N503);
  buf ginst162 (N1890, N514);
  buf ginst163 (N1893, N523);
  buf ginst164 (N1896, N534);
  buf ginst165 (N1899, N54);
  buf ginst166 (N1902, N479);
  buf ginst167 (N1905, N503);
  buf ginst168 (N1908, N514);
  buf ginst169 (N1911, N523);
  buf ginst170 (N1914, N534);
  buf ginst171 (N1917, N490);
  buf ginst172 (N1920, N361);
  buf ginst173 (N1923, N369);
  buf ginst174 (N1926, N341);
  buf ginst175 (N1929, N351);
  buf ginst176 (N1932, N308);
  buf ginst177 (N1935, N316);
  buf ginst178 (N1938, N293);
  buf ginst179 (N1941, N302);
  buf ginst180 (N1944, N281);
  buf ginst181 (N1947, N289);
  buf ginst182 (N1950, N265);
  buf ginst183 (N1953, N273);
  buf ginst184 (N1956, N234);
  buf ginst185 (N1959, N257);
  buf ginst186 (N1962, N218);
  buf ginst187 (N1965, N226);
  buf ginst188 (N1968, N210);
  not ginst189 (N1972, N1146);
  and ginst190 (N2054, N136, N1148);
  not ginst191 (N2060, N1150);
  not ginst192 (N2061, N1151);
  buf ginst193 (N2139, N1209);
  buf ginst194 (N2142, N1216);
  buf ginst195 (N2309, N1479);
  and ginst196 (N2349, N514, N1104);
  or ginst197 (N2350, N514, N1067);
  buf ginst198 (N2387, N1580);
  buf ginst199 (N2527, N1821);
  not ginst200 (N2584, N1580);
  and ginst201 (N2585, N170, N1161, N1173);
  and ginst202 (N2586, N173, N1161, N1173);
  and ginst203 (N2587, N167, N1161, N1173);
  and ginst204 (N2588, N164, N1161, N1173);
  and ginst205 (N2589, N161, N1161, N1173);
  nand ginst206 (N2590, N140, N1475);
  and ginst207 (N2591, N185, N1185, N1197);
  and ginst208 (N2592, N158, N1185, N1197);
  and ginst209 (N2593, N152, N1185, N1197);
  and ginst210 (N2594, N146, N1185, N1197);
  and ginst211 (N2595, N170, N1223, N1235);
  and ginst212 (N2596, N173, N1223, N1235);
  and ginst213 (N2597, N167, N1223, N1235);
  and ginst214 (N2598, N164, N1223, N1235);
  and ginst215 (N2599, N161, N1223, N1235);
  and ginst216 (N2600, N185, N1247, N1259);
  and ginst217 (N2601, N158, N1247, N1259);
  and ginst218 (N2602, N152, N1247, N1259);
  and ginst219 (N2603, N146, N1247, N1259);
  and ginst220 (N2604, N106, N1731, N1743);
  and ginst221 (N2605, N61, N1327, N1339);
  and ginst222 (N2606, N106, N1697, N1709);
  and ginst223 (N2607, N49, N1697, N1709);
  and ginst224 (N2608, N103, N1697, N1709);
  and ginst225 (N2609, N40, N1697, N1709);
  and ginst226 (N2610, N37, N1697, N1709);
  and ginst227 (N2611, N20, N1327, N1339);
  and ginst228 (N2612, N17, N1327, N1339);
  and ginst229 (N2613, N70, N1327, N1339);
  and ginst230 (N2614, N64, N1327, N1339);
  and ginst231 (N2615, N49, N1731, N1743);
  and ginst232 (N2616, N103, N1731, N1743);
  and ginst233 (N2617, N40, N1731, N1743);
  and ginst234 (N2618, N37, N1731, N1743);
  and ginst235 (N2619, N20, N1351, N1363);
  and ginst236 (N2620, N17, N1351, N1363);
  and ginst237 (N2621, N70, N1351, N1363);
  and ginst238 (N2622, N64, N1351, N1363);
  not ginst239 (N2623, N1475);
  and ginst240 (N2624, N123, N599, N1758);
  and ginst241 (N2625, N1777, N1785);
  and ginst242 (N2626, N61, N1351, N1363);
  and ginst243 (N2627, N1761, N1769);
  not ginst244 (N2628, N1824);
  not ginst245 (N2629, N1827);
  not ginst246 (N2630, N1830);
  not ginst247 (N2631, N1833);
  not ginst248 (N2632, N1836);
  not ginst249 (N2633, N1839);
  not ginst250 (N2634, N1842);
  not ginst251 (N2635, N1845);
  not ginst252 (N2636, N1848);
  not ginst253 (N2637, N1851);
  not ginst254 (N2638, N1854);
  not ginst255 (N2639, N1857);
  not ginst256 (N2640, N1860);
  not ginst257 (N2641, N1863);
  not ginst258 (N2642, N1866);
  not ginst259 (N2643, N1869);
  not ginst260 (N2644, N1872);
  not ginst261 (N2645, N1875);
  not ginst262 (N2646, N1878);
  buf ginst263 (N2647, N1209);
  not ginst264 (N2653, N1161);
  not ginst265 (N2664, N1173);
  buf ginst266 (N2675, N1209);
  not ginst267 (N2681, N1185);
  not ginst268 (N2692, N1197);
  and ginst269 (N2703, N179, N1185, N1197);
  buf ginst270 (N2704, N1479);
  not ginst271 (N2709, N1881);
  not ginst272 (N2710, N1884);
  not ginst273 (N2711, N1887);
  not ginst274 (N2712, N1890);
  not ginst275 (N2713, N1893);
  not ginst276 (N2714, N1896);
  not ginst277 (N2715, N1899);
  not ginst278 (N2716, N1902);
  not ginst279 (N2717, N1905);
  not ginst280 (N2718, N1908);
  not ginst281 (N2719, N1911);
  not ginst282 (N2720, N1914);
  not ginst283 (N2721, N1917);
  buf ginst284 (N2722, N1213);
  not ginst285 (N2728, N1223);
  not ginst286 (N2739, N1235);
  buf ginst287 (N2750, N1213);
  not ginst288 (N2756, N1247);
  not ginst289 (N2767, N1259);
  and ginst290 (N2778, N179, N1247, N1259);
  not ginst291 (N2779, N1327);
  not ginst292 (N2790, N1339);
  not ginst293 (N2801, N1351);
  not ginst294 (N2812, N1363);
  not ginst295 (N2823, N1375);
  not ginst296 (N2824, N1378);
  not ginst297 (N2825, N1381);
  not ginst298 (N2826, N1384);
  not ginst299 (N2827, N1387);
  not ginst300 (N2828, N1390);
  not ginst301 (N2829, N1393);
  not ginst302 (N2830, N1396);
  and ginst303 (N2831, N457, N1104, N1378);
  and ginst304 (N2832, N468, N1104, N1384);
  and ginst305 (N2833, N422, N1104, N1390);
  and ginst306 (N2834, N435, N1104, N1396);
  and ginst307 (N2835, N1067, N1375);
  and ginst308 (N2836, N1067, N1381);
  and ginst309 (N2837, N1067, N1387);
  and ginst310 (N2838, N1067, N1393);
  not ginst311 (N2839, N1415);
  not ginst312 (N2840, N1418);
  not ginst313 (N2841, N1421);
  not ginst314 (N2842, N1424);
  not ginst315 (N2843, N1427);
  not ginst316 (N2844, N1430);
  not ginst317 (N2845, N1433);
  not ginst318 (N2846, N1436);
  and ginst319 (N2847, N389, N1104, N1418);
  and ginst320 (N2848, N400, N1104, N1424);
  and ginst321 (N2849, N411, N1104, N1430);
  and ginst322 (N2850, N374, N1104, N1436);
  and ginst323 (N2851, N1067, N1415);
  and ginst324 (N2852, N1067, N1421);
  and ginst325 (N2853, N1067, N1427);
  and ginst326 (N2854, N1067, N1433);
  not ginst327 (N2855, N1455);
  not ginst328 (N2861, N1462);
  and ginst329 (N2867, N292, N1455);
  and ginst330 (N2868, N288, N1455);
  and ginst331 (N2869, N280, N1455);
  and ginst332 (N2870, N272, N1455);
  and ginst333 (N2871, N264, N1455);
  and ginst334 (N2872, N241, N1462);
  and ginst335 (N2873, N233, N1462);
  and ginst336 (N2874, N225, N1462);
  and ginst337 (N2875, N217, N1462);
  and ginst338 (N2876, N209, N1462);
  buf ginst339 (N2877, N1216);
  not ginst340 (N2882, N1482);
  not ginst341 (N2891, N1475);
  not ginst342 (N2901, N1492);
  not ginst343 (N2902, N1495);
  not ginst344 (N2903, N1498);
  not ginst345 (N2904, N1501);
  not ginst346 (N2905, N1504);
  not ginst347 (N2906, N1507);
  and ginst348 (N2907, N1303, N1495);
  and ginst349 (N2908, N479, N1303, N1501);
  and ginst350 (N2909, N490, N1303, N1507);
  and ginst351 (N2910, N1492, N1663);
  and ginst352 (N2911, N1498, N1663);
  and ginst353 (N2912, N1504, N1663);
  not ginst354 (N2913, N1510);
  not ginst355 (N2914, N1513);
  not ginst356 (N2915, N1516);
  not ginst357 (N2916, N1519);
  not ginst358 (N2917, N1522);
  not ginst359 (N2918, N1525);
  and ginst360 (N2919, N503, N1104, N1513);
  not ginst361 (N2920, N2349);
  and ginst362 (N2921, N523, N1104, N1519);
  and ginst363 (N2922, N534, N1104, N1525);
  and ginst364 (N2923, N1067, N1510);
  and ginst365 (N2924, N1067, N1516);
  and ginst366 (N2925, N1067, N1522);
  not ginst367 (N2926, N1542);
  not ginst368 (N2927, N1545);
  not ginst369 (N2928, N1548);
  not ginst370 (N2929, N1551);
  not ginst371 (N2930, N1554);
  not ginst372 (N2931, N1557);
  not ginst373 (N2932, N1560);
  not ginst374 (N2933, N1563);
  and ginst375 (N2934, N389, N1303, N1545);
  and ginst376 (N2935, N400, N1303, N1551);
  and ginst377 (N2936, N411, N1303, N1557);
  and ginst378 (N2937, N374, N1303, N1563);
  and ginst379 (N2938, N1542, N1663);
  and ginst380 (N2939, N1548, N1663);
  and ginst381 (N2940, N1554, N1663);
  and ginst382 (N2941, N1560, N1663);
  not ginst383 (N2942, N1566);
  not ginst384 (N2948, N1573);
  and ginst385 (N2954, N372, N1566);
  and ginst386 (N2955, N366, N1566);
  and ginst387 (N2956, N358, N1566);
  and ginst388 (N2957, N348, N1566);
  and ginst389 (N2958, N338, N1566);
  and ginst390 (N2959, N331, N1573);
  and ginst391 (N2960, N323, N1573);
  and ginst392 (N2961, N315, N1573);
  and ginst393 (N2962, N307, N1573);
  and ginst394 (N2963, N299, N1573);
  not ginst395 (N2964, N1588);
  and ginst396 (N2969, N83, N1588);
  and ginst397 (N2970, N86, N1588);
  and ginst398 (N2971, N88, N1588);
  and ginst399 (N2972, N88, N1588);
  not ginst400 (N2973, N1594);
  not ginst401 (N2974, N1597);
  not ginst402 (N2975, N1600);
  not ginst403 (N2976, N1603);
  not ginst404 (N2977, N1606);
  not ginst405 (N2978, N1609);
  and ginst406 (N2979, N503, N1315, N1597);
  and ginst407 (N2980, N514, N1315);
  and ginst408 (N2981, N523, N1315, N1603);
  and ginst409 (N2982, N534, N1315, N1609);
  and ginst410 (N2983, N1594, N1675);
  or ginst411 (N2984, N514, N1675);
  and ginst412 (N2985, N1600, N1675);
  and ginst413 (N2986, N1606, N1675);
  not ginst414 (N2987, N1612);
  not ginst415 (N2988, N1615);
  not ginst416 (N2989, N1618);
  not ginst417 (N2990, N1621);
  not ginst418 (N2991, N1624);
  not ginst419 (N2992, N1627);
  and ginst420 (N2993, N1315, N1615);
  and ginst421 (N2994, N479, N1315, N1621);
  and ginst422 (N2995, N490, N1315, N1627);
  and ginst423 (N2996, N1612, N1675);
  and ginst424 (N2997, N1618, N1675);
  and ginst425 (N2998, N1624, N1675);
  not ginst426 (N2999, N1630);
  buf ginst427 (N3000, N1469);
  buf ginst428 (N3003, N1469);
  not ginst429 (N3006, N1633);
  buf ginst430 (N3007, N1469);
  buf ginst431 (N3010, N1469);
  and ginst432 (N3013, N1315, N1630);
  and ginst433 (N3014, N1315, N1633);
  not ginst434 (N3015, N1636);
  not ginst435 (N3016, N1639);
  not ginst436 (N3017, N1642);
  not ginst437 (N3018, N1645);
  not ginst438 (N3019, N1648);
  not ginst439 (N3020, N1651);
  not ginst440 (N3021, N1654);
  not ginst441 (N3022, N1657);
  and ginst442 (N3023, N457, N1303, N1639);
  and ginst443 (N3024, N468, N1303, N1645);
  and ginst444 (N3025, N422, N1303, N1651);
  and ginst445 (N3026, N435, N1303, N1657);
  and ginst446 (N3027, N1636, N1663);
  and ginst447 (N3028, N1642, N1663);
  and ginst448 (N3029, N1648, N1663);
  and ginst449 (N3030, N1654, N1663);
  not ginst450 (N3031, N1920);
  not ginst451 (N3032, N1923);
  not ginst452 (N3033, N1926);
  not ginst453 (N3034, N1929);
  buf ginst454 (N3035, N1660);
  buf ginst455 (N3038, N1660);
  not ginst456 (N3041, N1697);
  not ginst457 (N3052, N1709);
  not ginst458 (N3063, N1721);
  not ginst459 (N3068, N1727);
  and ginst460 (N3071, N97, N1721);
  and ginst461 (N3072, N94, N1721);
  and ginst462 (N3073, N97, N1721);
  and ginst463 (N3074, N94, N1721);
  not ginst464 (N3075, N1731);
  not ginst465 (N3086, N1743);
  not ginst466 (N3097, N1761);
  not ginst467 (N3108, N1769);
  not ginst468 (N3119, N1777);
  not ginst469 (N3130, N1785);
  not ginst470 (N3141, N1944);
  not ginst471 (N3142, N1947);
  not ginst472 (N3143, N1950);
  not ginst473 (N3144, N1953);
  not ginst474 (N3145, N1956);
  not ginst475 (N3146, N1959);
  not ginst476 (N3147, N1793);
  not ginst477 (N3158, N1800);
  not ginst478 (N3169, N1807);
  not ginst479 (N3180, N1814);
  buf ginst480 (N3191, N1821);
  not ginst481 (N3194, N1932);
  not ginst482 (N3195, N1935);
  not ginst483 (N3196, N1938);
  not ginst484 (N3197, N1941);
  not ginst485 (N3198, N1962);
  not ginst486 (N3199, N1965);
  buf ginst487 (N3200, N1469);
  not ginst488 (N3203, N1968);
  buf ginst489 (N3357, N2704);
  buf ginst490 (N3358, N2704);
  buf ginst491 (N3359, N2704);
  buf ginst492 (N3360, N2704);
  and ginst493 (N3401, N457, N1092, N2824);
  and ginst494 (N3402, N468, N1092, N2826);
  and ginst495 (N3403, N422, N1092, N2828);
  and ginst496 (N3404, N435, N1092, N2830);
  and ginst497 (N3405, N1080, N2823);
  and ginst498 (N3406, N1080, N2825);
  and ginst499 (N3407, N1080, N2827);
  and ginst500 (N3408, N1080, N2829);
  and ginst501 (N3409, N389, N1092, N2840);
  and ginst502 (N3410, N400, N1092, N2842);
  and ginst503 (N3411, N411, N1092, N2844);
  and ginst504 (N3412, N374, N1092, N2846);
  and ginst505 (N3413, N1080, N2839);
  and ginst506 (N3414, N1080, N2841);
  and ginst507 (N3415, N1080, N2843);
  and ginst508 (N3416, N1080, N2845);
  and ginst509 (N3444, N1280, N2902);
  and ginst510 (N3445, N479, N1280, N2904);
  and ginst511 (N3446, N490, N1280, N2906);
  and ginst512 (N3447, N1685, N2901);
  and ginst513 (N3448, N1685, N2903);
  and ginst514 (N3449, N1685, N2905);
  and ginst515 (N3450, N503, N1092, N2914);
  and ginst516 (N3451, N523, N1092, N2916);
  and ginst517 (N3452, N534, N1092, N2918);
  and ginst518 (N3453, N1080, N2913);
  and ginst519 (N3454, N1080, N2915);
  and ginst520 (N3455, N1080, N2917);
  and ginst521 (N3456, N2350, N2920);
  and ginst522 (N3459, N389, N1280, N2927);
  and ginst523 (N3460, N400, N1280, N2929);
  and ginst524 (N3461, N411, N1280, N2931);
  and ginst525 (N3462, N374, N1280, N2933);
  and ginst526 (N3463, N1685, N2926);
  and ginst527 (N3464, N1685, N2928);
  and ginst528 (N3465, N1685, N2930);
  and ginst529 (N3466, N1685, N2932);
  and ginst530 (N3481, N503, N1292, N2974);
  not ginst531 (N3482, N2980);
  and ginst532 (N3483, N523, N1292, N2976);
  and ginst533 (N3484, N534, N1292, N2978);
  and ginst534 (N3485, N1271, N2973);
  and ginst535 (N3486, N1271, N2975);
  and ginst536 (N3487, N1271, N2977);
  and ginst537 (N3488, N1292, N2988);
  and ginst538 (N3489, N479, N1292, N2990);
  and ginst539 (N3490, N490, N1292, N2992);
  and ginst540 (N3491, N1271, N2987);
  and ginst541 (N3492, N1271, N2989);
  and ginst542 (N3493, N1271, N2991);
  and ginst543 (N3502, N1292, N2999);
  and ginst544 (N3503, N1292, N3006);
  and ginst545 (N3504, N457, N1280, N3016);
  and ginst546 (N3505, N468, N1280, N3018);
  and ginst547 (N3506, N422, N1280, N3020);
  and ginst548 (N3507, N435, N1280, N3022);
  and ginst549 (N3508, N1685, N3015);
  and ginst550 (N3509, N1685, N3017);
  and ginst551 (N3510, N1685, N3019);
  and ginst552 (N3511, N1685, N3021);
  nand ginst553 (N3512, N1923, N3031);
  nand ginst554 (N3513, N1920, N3032);
  nand ginst555 (N3514, N1929, N3033);
  nand ginst556 (N3515, N1926, N3034);
  nand ginst557 (N3558, N1947, N3141);
  nand ginst558 (N3559, N1944, N3142);
  nand ginst559 (N3560, N1953, N3143);
  nand ginst560 (N3561, N1950, N3144);
  nand ginst561 (N3562, N1959, N3145);
  nand ginst562 (N3563, N1956, N3146);
  buf ginst563 (N3604, N3191);
  nand ginst564 (N3605, N1935, N3194);
  nand ginst565 (N3606, N1932, N3195);
  nand ginst566 (N3607, N1941, N3196);
  nand ginst567 (N3608, N1938, N3197);
  nand ginst568 (N3609, N1965, N3198);
  nand ginst569 (N3610, N1962, N3199);
  not ginst570 (N3613, N3191);
  and ginst571 (N3614, N2882, N2891);
  and ginst572 (N3615, N1482, N2891);
  and ginst573 (N3616, N200, N1173, N2653);
  and ginst574 (N3617, N203, N1173, N2653);
  and ginst575 (N3618, N197, N1173, N2653);
  and ginst576 (N3619, N194, N1173, N2653);
  and ginst577 (N3620, N191, N1173, N2653);
  and ginst578 (N3621, N182, N1197, N2681);
  and ginst579 (N3622, N188, N1197, N2681);
  and ginst580 (N3623, N155, N1197, N2681);
  and ginst581 (N3624, N149, N1197, N2681);
  and ginst582 (N3625, N2882, N2891);
  and ginst583 (N3626, N1482, N2891);
  and ginst584 (N3627, N200, N1235, N2728);
  and ginst585 (N3628, N203, N1235, N2728);
  and ginst586 (N3629, N197, N1235, N2728);
  and ginst587 (N3630, N194, N1235, N2728);
  and ginst588 (N3631, N191, N1235, N2728);
  and ginst589 (N3632, N182, N1259, N2756);
  and ginst590 (N3633, N188, N1259, N2756);
  and ginst591 (N3634, N155, N1259, N2756);
  and ginst592 (N3635, N149, N1259, N2756);
  and ginst593 (N3636, N2882, N2891);
  and ginst594 (N3637, N1482, N2891);
  and ginst595 (N3638, N109, N1743, N3075);
  and ginst596 (N3639, N2882, N2891);
  and ginst597 (N3640, N1482, N2891);
  and ginst598 (N3641, N11, N1339, N2779);
  and ginst599 (N3642, N109, N1709, N3041);
  and ginst600 (N3643, N46, N1709, N3041);
  and ginst601 (N3644, N100, N1709, N3041);
  and ginst602 (N3645, N91, N1709, N3041);
  and ginst603 (N3646, N43, N1709, N3041);
  and ginst604 (N3647, N76, N1339, N2779);
  and ginst605 (N3648, N73, N1339, N2779);
  and ginst606 (N3649, N67, N1339, N2779);
  and ginst607 (N3650, N14, N1339, N2779);
  and ginst608 (N3651, N46, N1743, N3075);
  and ginst609 (N3652, N100, N1743, N3075);
  and ginst610 (N3653, N91, N1743, N3075);
  and ginst611 (N3654, N43, N1743, N3075);
  and ginst612 (N3655, N76, N1363, N2801);
  and ginst613 (N3656, N73, N1363, N2801);
  and ginst614 (N3657, N67, N1363, N2801);
  and ginst615 (N3658, N14, N1363, N2801);
  and ginst616 (N3659, N120, N1785, N3119);
  and ginst617 (N3660, N11, N1363, N2801);
  and ginst618 (N3661, N118, N1769, N3097);
  and ginst619 (N3662, N176, N1197, N2681);
  and ginst620 (N3663, N176, N1259, N2756);
  or ginst621 (N3664, N2831, N3401);
  or ginst622 (N3665, N2832, N3402);
  or ginst623 (N3666, N2833, N3403);
  or ginst624 (N3667, N2834, N3404);
  or ginst625 (N3668, N457, N2835, N3405);
  or ginst626 (N3669, N468, N2836, N3406);
  or ginst627 (N3670, N422, N2837, N3407);
  or ginst628 (N3671, N435, N2838, N3408);
  or ginst629 (N3672, N2847, N3409);
  or ginst630 (N3673, N2848, N3410);
  or ginst631 (N3674, N2849, N3411);
  or ginst632 (N3675, N2850, N3412);
  or ginst633 (N3676, N389, N2851, N3413);
  or ginst634 (N3677, N400, N2852, N3414);
  or ginst635 (N3678, N411, N2853, N3415);
  or ginst636 (N3679, N374, N2854, N3416);
  and ginst637 (N3680, N289, N2855);
  and ginst638 (N3681, N281, N2855);
  and ginst639 (N3682, N273, N2855);
  and ginst640 (N3683, N265, N2855);
  and ginst641 (N3684, N257, N2855);
  and ginst642 (N3685, N234, N2861);
  and ginst643 (N3686, N226, N2861);
  and ginst644 (N3687, N218, N2861);
  and ginst645 (N3688, N210, N2861);
  and ginst646 (N3689, N206, N2861);
  not ginst647 (N3691, N2891);
  or ginst648 (N3700, N2907, N3444);
  or ginst649 (N3701, N2908, N3445);
  or ginst650 (N3702, N2909, N3446);
  or ginst651 (N3703, N479, N2911, N3448);
  or ginst652 (N3704, N490, N2912, N3449);
  or ginst653 (N3705, N2910, N3447);
  or ginst654 (N3708, N2919, N3450);
  or ginst655 (N3709, N2921, N3451);
  or ginst656 (N3710, N2922, N3452);
  or ginst657 (N3711, N503, N2923, N3453);
  or ginst658 (N3712, N523, N2924, N3454);
  or ginst659 (N3713, N534, N2925, N3455);
  or ginst660 (N3715, N2934, N3459);
  or ginst661 (N3716, N2935, N3460);
  or ginst662 (N3717, N2936, N3461);
  or ginst663 (N3718, N2937, N3462);
  or ginst664 (N3719, N389, N2938, N3463);
  or ginst665 (N3720, N400, N2939, N3464);
  or ginst666 (N3721, N411, N2940, N3465);
  or ginst667 (N3722, N374, N2941, N3466);
  and ginst668 (N3723, N369, N2942);
  and ginst669 (N3724, N361, N2942);
  and ginst670 (N3725, N351, N2942);
  and ginst671 (N3726, N341, N2942);
  and ginst672 (N3727, N324, N2948);
  and ginst673 (N3728, N316, N2948);
  and ginst674 (N3729, N308, N2948);
  and ginst675 (N3730, N302, N2948);
  and ginst676 (N3731, N293, N2948);
  or ginst677 (N3732, N2942, N2958);
  and ginst678 (N3738, N83, N2964);
  and ginst679 (N3739, N87, N2964);
  and ginst680 (N3740, N34, N2964);
  and ginst681 (N3741, N34, N2964);
  or ginst682 (N3742, N2979, N3481);
  or ginst683 (N3743, N2981, N3483);
  or ginst684 (N3744, N2982, N3484);
  or ginst685 (N3745, N503, N2983, N3485);
  or ginst686 (N3746, N523, N2985, N3486);
  or ginst687 (N3747, N534, N2986, N3487);
  or ginst688 (N3748, N2993, N3488);
  or ginst689 (N3749, N2994, N3489);
  or ginst690 (N3750, N2995, N3490);
  or ginst691 (N3751, N479, N2997, N3492);
  or ginst692 (N3752, N490, N2998, N3493);
  not ginst693 (N3753, N3000);
  not ginst694 (N3754, N3003);
  not ginst695 (N3755, N3007);
  not ginst696 (N3756, N3010);
  or ginst697 (N3757, N3013, N3502);
  and ginst698 (N3758, N446, N1315, N3003);
  or ginst699 (N3759, N3014, N3503);
  and ginst700 (N3760, N446, N1315, N3010);
  and ginst701 (N3761, N1675, N3000);
  and ginst702 (N3762, N1675, N3007);
  or ginst703 (N3763, N3023, N3504);
  or ginst704 (N3764, N3024, N3505);
  or ginst705 (N3765, N3025, N3506);
  or ginst706 (N3766, N3026, N3507);
  or ginst707 (N3767, N457, N3027, N3508);
  or ginst708 (N3768, N468, N3028, N3509);
  or ginst709 (N3769, N422, N3029, N3510);
  or ginst710 (N3770, N435, N3030, N3511);
  nand ginst711 (N3771, N3512, N3513);
  nand ginst712 (N3775, N3514, N3515);
  not ginst713 (N3779, N3035);
  not ginst714 (N3780, N3038);
  and ginst715 (N3781, N117, N1769, N3097);
  and ginst716 (N3782, N126, N1769, N3097);
  and ginst717 (N3783, N127, N1769, N3097);
  and ginst718 (N3784, N128, N1769, N3097);
  and ginst719 (N3785, N131, N1785, N3119);
  and ginst720 (N3786, N129, N1785, N3119);
  and ginst721 (N3787, N119, N1785, N3119);
  and ginst722 (N3788, N130, N1785, N3119);
  nand ginst723 (N3789, N3558, N3559);
  nand ginst724 (N3793, N3560, N3561);
  nand ginst725 (N3797, N3562, N3563);
  and ginst726 (N3800, N122, N1800, N3147);
  and ginst727 (N3801, N113, N1800, N3147);
  and ginst728 (N3802, N53, N1800, N3147);
  and ginst729 (N3803, N114, N1800, N3147);
  and ginst730 (N3804, N115, N1800, N3147);
  and ginst731 (N3805, N52, N1814, N3169);
  and ginst732 (N3806, N112, N1814, N3169);
  and ginst733 (N3807, N116, N1814, N3169);
  and ginst734 (N3808, N121, N1814, N3169);
  and ginst735 (N3809, N123, N1814, N3169);
  nand ginst736 (N3810, N3607, N3608);
  nand ginst737 (N3813, N3605, N3606);
  and ginst738 (N3816, N2984, N3482);
  or ginst739 (N3819, N2996, N3491);
  not ginst740 (N3822, N3200);
  nand ginst741 (N3823, N3200, N3203);
  nand ginst742 (N3824, N3609, N3610);
  not ginst743 (N3827, N3456);
  or ginst744 (N3828, N2970, N3739);
  or ginst745 (N3829, N2971, N3740);
  or ginst746 (N3830, N2972, N3741);
  or ginst747 (N3831, N2969, N3738);
  not ginst748 (N3834, N3664);
  not ginst749 (N3835, N3665);
  not ginst750 (N3836, N3666);
  not ginst751 (N3837, N3667);
  not ginst752 (N3838, N3672);
  not ginst753 (N3839, N3673);
  not ginst754 (N3840, N3674);
  not ginst755 (N3841, N3675);
  or ginst756 (N3842, N2868, N3681);
  or ginst757 (N3849, N2869, N3682);
  or ginst758 (N3855, N2870, N3683);
  or ginst759 (N3861, N2871, N3684);
  or ginst760 (N3867, N2872, N3685);
  or ginst761 (N3873, N2873, N3686);
  or ginst762 (N3881, N2874, N3687);
  or ginst763 (N3887, N2875, N3688);
  or ginst764 (N3893, N2876, N3689);
  not ginst765 (N3908, N3701);
  not ginst766 (N3909, N3702);
  not ginst767 (N3911, N3700);
  not ginst768 (N3914, N3708);
  not ginst769 (N3915, N3709);
  not ginst770 (N3916, N3710);
  not ginst771 (N3917, N3715);
  not ginst772 (N3918, N3716);
  not ginst773 (N3919, N3717);
  not ginst774 (N3920, N3718);
  or ginst775 (N3921, N2955, N3724);
  or ginst776 (N3927, N2956, N3725);
  or ginst777 (N3933, N2957, N3726);
  or ginst778 (N3942, N2959, N3727);
  or ginst779 (N3948, N2960, N3728);
  or ginst780 (N3956, N2961, N3729);
  or ginst781 (N3962, N2962, N3730);
  or ginst782 (N3968, N2963, N3731);
  not ginst783 (N3975, N3742);
  not ginst784 (N3976, N3743);
  not ginst785 (N3977, N3744);
  not ginst786 (N3978, N3749);
  not ginst787 (N3979, N3750);
  and ginst788 (N3980, N446, N1292, N3754);
  and ginst789 (N3981, N446, N1292, N3756);
  and ginst790 (N3982, N1271, N3753);
  and ginst791 (N3983, N1271, N3755);
  not ginst792 (N3984, N3757);
  not ginst793 (N3987, N3759);
  not ginst794 (N3988, N3763);
  not ginst795 (N3989, N3764);
  not ginst796 (N3990, N3765);
  not ginst797 (N3991, N3766);
  and ginst798 (N3998, N3119, N3130, N3456);
  or ginst799 (N4008, N2954, N3723);
  or ginst800 (N4011, N2867, N3680);
  not ginst801 (N4021, N3748);
  nand ginst802 (N4024, N1968, N3822);
  not ginst803 (N4027, N3705);
  and ginst804 (N4031, N1583, N3828);
  and ginst805 (N4032, N24, N2882, N3691);
  and ginst806 (N4033, N25, N1482, N3691);
  and ginst807 (N4034, N26, N2882, N3691);
  and ginst808 (N4035, N81, N1482, N3691);
  and ginst809 (N4036, N1583, N3829);
  and ginst810 (N4037, N79, N2882, N3691);
  and ginst811 (N4038, N23, N1482, N3691);
  and ginst812 (N4039, N82, N2882, N3691);
  and ginst813 (N4040, N80, N1482, N3691);
  and ginst814 (N4041, N1583, N3830);
  and ginst815 (N4042, N1583, N3831);
  and ginst816 (N4067, N514, N3732);
  and ginst817 (N4080, N514, N3732);
  and ginst818 (N4088, N3668, N3834);
  and ginst819 (N4091, N3669, N3835);
  and ginst820 (N4094, N3670, N3836);
  and ginst821 (N4097, N3671, N3837);
  and ginst822 (N4100, N3676, N3838);
  and ginst823 (N4103, N3677, N3839);
  and ginst824 (N4106, N3678, N3840);
  and ginst825 (N4109, N3679, N3841);
  and ginst826 (N4144, N3703, N3908);
  and ginst827 (N4147, N3704, N3909);
  buf ginst828 (N4150, N3705);
  and ginst829 (N4153, N3711, N3914);
  and ginst830 (N4156, N3712, N3915);
  and ginst831 (N4159, N3713, N3916);
  or ginst832 (N4183, N3758, N3980);
  or ginst833 (N4184, N3760, N3981);
  or ginst834 (N4185, N446, N3761, N3982);
  or ginst835 (N4186, N446, N3762, N3983);
  not ginst836 (N4188, N3771);
  not ginst837 (N4191, N3775);
  and ginst838 (N4196, N3035, N3771, N3775);
  and ginst839 (N4197, N3119, N3130, N3987);
  and ginst840 (N4198, N3722, N3920);
  not ginst841 (N4199, N3816);
  not ginst842 (N4200, N3789);
  not ginst843 (N4203, N3793);
  buf ginst844 (N4206, N3797);
  buf ginst845 (N4209, N3797);
  buf ginst846 (N4212, N3732);
  buf ginst847 (N4215, N3732);
  buf ginst848 (N4219, N3732);
  not ginst849 (N4223, N3810);
  not ginst850 (N4224, N3813);
  and ginst851 (N4225, N3720, N3918);
  and ginst852 (N4228, N3721, N3919);
  and ginst853 (N4231, N3770, N3991);
  and ginst854 (N4234, N3719, N3917);
  and ginst855 (N4237, N3768, N3989);
  and ginst856 (N4240, N3769, N3990);
  and ginst857 (N4243, N3767, N3988);
  and ginst858 (N4246, N3746, N3976);
  and ginst859 (N4249, N3747, N3977);
  and ginst860 (N4252, N3745, N3975);
  and ginst861 (N4255, N3751, N3978);
  and ginst862 (N4258, N3752, N3979);
  not ginst863 (N4263, N3819);
  nand ginst864 (N4264, N3823, N4024);
  not ginst865 (N4267, N3824);
  and ginst866 (N4268, N446, N3893);
  not ginst867 (N4269, N3911);
  not ginst868 (N4270, N3984);
  and ginst869 (N4271, N446, N3893);
  not ginst870 (N4272, N4031);
  or ginst871 (N4273, N3614, N3615, N4032, N4033);
  or ginst872 (N4274, N3625, N3626, N4034, N4035);
  not ginst873 (N4275, N4036);
  or ginst874 (N4276, N3636, N3637, N4037, N4038);
  or ginst875 (N4277, N3639, N3640, N4039, N4040);
  not ginst876 (N4278, N4041);
  not ginst877 (N4279, N4042);
  and ginst878 (N4280, N457, N3887);
  and ginst879 (N4284, N468, N3881);
  and ginst880 (N4290, N422, N3873);
  and ginst881 (N4297, N435, N3867);
  and ginst882 (N4298, N389, N3861);
  and ginst883 (N4301, N400, N3855);
  and ginst884 (N4305, N411, N3849);
  and ginst885 (N4310, N374, N3842);
  and ginst886 (N4316, N457, N3887);
  and ginst887 (N4320, N468, N3881);
  and ginst888 (N4325, N422, N3873);
  and ginst889 (N4331, N435, N3867);
  and ginst890 (N4332, N389, N3861);
  and ginst891 (N4336, N400, N3855);
  and ginst892 (N4342, N411, N3849);
  and ginst893 (N4349, N374, N3842);
  not ginst894 (N4357, N3968);
  not ginst895 (N4364, N3962);
  buf ginst896 (N4375, N3962);
  and ginst897 (N4379, N479, N3956);
  and ginst898 (N4385, N490, N3948);
  and ginst899 (N4392, N503, N3942);
  and ginst900 (N4396, N523, N3933);
  and ginst901 (N4400, N534, N3927);
  not ginst902 (N4405, N3921);
  buf ginst903 (N4412, N3921);
  not ginst904 (N4418, N3968);
  not ginst905 (N4425, N3962);
  buf ginst906 (N4436, N3962);
  and ginst907 (N4440, N479, N3956);
  and ginst908 (N4445, N490, N3948);
  and ginst909 (N4451, N503, N3942);
  and ginst910 (N4456, N523, N3933);
  and ginst911 (N4462, N534, N3927);
  buf ginst912 (N4469, N3921);
  not ginst913 (N4477, N3921);
  buf ginst914 (N4512, N3968);
  not ginst915 (N4515, N4183);
  not ginst916 (N4516, N4184);
  not ginst917 (N4521, N4008);
  not ginst918 (N4523, N4011);
  not ginst919 (N4524, N4198);
  not ginst920 (N4532, N3984);
  and ginst921 (N4547, N3169, N3180, N3911);
  buf ginst922 (N4548, N3893);
  buf ginst923 (N4551, N3887);
  buf ginst924 (N4554, N3881);
  buf ginst925 (N4557, N3873);
  buf ginst926 (N4560, N3867);
  buf ginst927 (N4563, N3861);
  buf ginst928 (N4566, N3855);
  buf ginst929 (N4569, N3849);
  buf ginst930 (N4572, N3842);
  nor ginst931 (N4575, N422, N3873);
  buf ginst932 (N4578, N3893);
  buf ginst933 (N4581, N3887);
  buf ginst934 (N4584, N3881);
  buf ginst935 (N4587, N3867);
  buf ginst936 (N4590, N3861);
  buf ginst937 (N4593, N3855);
  buf ginst938 (N4596, N3849);
  buf ginst939 (N4599, N3873);
  buf ginst940 (N4602, N3842);
  nor ginst941 (N4605, N422, N3873);
  nor ginst942 (N4608, N374, N3842);
  buf ginst943 (N4611, N3956);
  buf ginst944 (N4614, N3948);
  buf ginst945 (N4617, N3942);
  buf ginst946 (N4621, N3933);
  buf ginst947 (N4624, N3927);
  nor ginst948 (N4627, N490, N3948);
  buf ginst949 (N4630, N3956);
  buf ginst950 (N4633, N3942);
  buf ginst951 (N4637, N3933);
  buf ginst952 (N4640, N3927);
  buf ginst953 (N4643, N3948);
  nor ginst954 (N4646, N490, N3948);
  buf ginst955 (N4649, N3927);
  buf ginst956 (N4652, N3933);
  buf ginst957 (N4655, N3921);
  buf ginst958 (N4658, N3942);
  buf ginst959 (N4662, N3956);
  buf ginst960 (N4665, N3948);
  buf ginst961 (N4668, N3968);
  buf ginst962 (N4671, N3962);
  buf ginst963 (N4674, N3873);
  buf ginst964 (N4677, N3867);
  buf ginst965 (N4680, N3887);
  buf ginst966 (N4683, N3881);
  buf ginst967 (N4686, N3893);
  buf ginst968 (N4689, N3849);
  buf ginst969 (N4692, N3842);
  buf ginst970 (N4695, N3861);
  buf ginst971 (N4698, N3855);
  nand ginst972 (N4701, N3813, N4223);
  nand ginst973 (N4702, N3810, N4224);
  not ginst974 (N4720, N4021);
  nand ginst975 (N4721, N4021, N4263);
  not ginst976 (N4724, N4147);
  not ginst977 (N4725, N4144);
  not ginst978 (N4726, N4159);
  not ginst979 (N4727, N4156);
  not ginst980 (N4728, N4153);
  not ginst981 (N4729, N4097);
  not ginst982 (N4730, N4094);
  not ginst983 (N4731, N4091);
  not ginst984 (N4732, N4088);
  not ginst985 (N4733, N4109);
  not ginst986 (N4734, N4106);
  not ginst987 (N4735, N4103);
  not ginst988 (N4736, N4100);
  and ginst989 (N4737, N2877, N4273);
  and ginst990 (N4738, N2877, N4274);
  and ginst991 (N4739, N2877, N4276);
  and ginst992 (N4740, N2877, N4277);
  and ginst993 (N4741, N1755, N1758, N4150);
  not ginst994 (N4855, N4212);
  nand ginst995 (N4856, N2712, N4212);
  nand ginst996 (N4908, N2718, N4215);
  not ginst997 (N4909, N4215);
  and ginst998 (N4939, N4185, N4515);
  and ginst999 (N4942, N4186, N4516);
  not ginst1000 (N4947, N4219);
  and ginst1001 (N4953, N3775, N3779, N4188);
  and ginst1002 (N4954, N3771, N3780, N4191);
  and ginst1003 (N4955, N3038, N4188, N4191);
  and ginst1004 (N4956, N3097, N3108, N4109);
  and ginst1005 (N4957, N3097, N3108, N4106);
  and ginst1006 (N4958, N3097, N3108, N4103);
  and ginst1007 (N4959, N3097, N3108, N4100);
  and ginst1008 (N4960, N3119, N3130, N4159);
  and ginst1009 (N4961, N3119, N3130, N4156);
  not ginst1010 (N4965, N4225);
  not ginst1011 (N4966, N4228);
  not ginst1012 (N4967, N4231);
  not ginst1013 (N4968, N4234);
  not ginst1014 (N4972, N4246);
  not ginst1015 (N4973, N4249);
  not ginst1016 (N4974, N4252);
  nand ginst1017 (N4975, N4199, N4252);
  not ginst1018 (N4976, N4206);
  not ginst1019 (N4977, N4209);
  and ginst1020 (N4978, N3789, N3793, N4206);
  and ginst1021 (N4979, N4200, N4203, N4209);
  and ginst1022 (N4980, N3147, N3158, N4097);
  and ginst1023 (N4981, N3147, N3158, N4094);
  and ginst1024 (N4982, N3147, N3158, N4091);
  and ginst1025 (N4983, N3147, N3158, N4088);
  and ginst1026 (N4984, N3169, N3180, N4153);
  and ginst1027 (N4985, N3169, N3180, N4147);
  and ginst1028 (N4986, N3169, N3180, N4144);
  and ginst1029 (N4987, N3169, N3180, N4150);
  nand ginst1030 (N5049, N4701, N4702);
  not ginst1031 (N5052, N4237);
  not ginst1032 (N5053, N4240);
  not ginst1033 (N5054, N4243);
  not ginst1034 (N5055, N4255);
  not ginst1035 (N5056, N4258);
  nand ginst1036 (N5057, N3819, N4720);
  not ginst1037 (N5058, N4264);
  nand ginst1038 (N5059, N4264, N4267);
  and ginst1039 (N5060, N4027, N4269, N4724, N4725);
  and ginst1040 (N5061, N3827, N4726, N4727, N4728);
  and ginst1041 (N5062, N4729, N4730, N4731, N4732);
  and ginst1042 (N5063, N4733, N4734, N4735, N4736);
  and ginst1043 (N5065, N4357, N4375);
  and ginst1044 (N5066, N4357, N4364, N4379);
  and ginst1045 (N5067, N4418, N4436);
  and ginst1046 (N5068, N4418, N4425, N4440);
  not ginst1047 (N5069, N4548);
  nand ginst1048 (N5070, N2628, N4548);
  not ginst1049 (N5071, N4551);
  nand ginst1050 (N5072, N2629, N4551);
  not ginst1051 (N5073, N4554);
  nand ginst1052 (N5074, N2630, N4554);
  not ginst1053 (N5075, N4557);
  nand ginst1054 (N5076, N2631, N4557);
  not ginst1055 (N5077, N4560);
  nand ginst1056 (N5078, N2632, N4560);
  not ginst1057 (N5079, N4563);
  nand ginst1058 (N5080, N2633, N4563);
  not ginst1059 (N5081, N4566);
  nand ginst1060 (N5082, N2634, N4566);
  not ginst1061 (N5083, N4569);
  nand ginst1062 (N5084, N2635, N4569);
  not ginst1063 (N5085, N4572);
  nand ginst1064 (N5086, N2636, N4572);
  not ginst1065 (N5087, N4575);
  nand ginst1066 (N5088, N2638, N4578);
  not ginst1067 (N5089, N4578);
  nand ginst1068 (N5090, N2639, N4581);
  not ginst1069 (N5091, N4581);
  nand ginst1070 (N5092, N2640, N4584);
  not ginst1071 (N5093, N4584);
  nand ginst1072 (N5094, N2641, N4587);
  not ginst1073 (N5095, N4587);
  nand ginst1074 (N5096, N2642, N4590);
  not ginst1075 (N5097, N4590);
  nand ginst1076 (N5098, N2643, N4593);
  not ginst1077 (N5099, N4593);
  nand ginst1078 (N5100, N2644, N4596);
  not ginst1079 (N5101, N4596);
  nand ginst1080 (N5102, N2645, N4599);
  not ginst1081 (N5103, N4599);
  nand ginst1082 (N5104, N2646, N4602);
  not ginst1083 (N5105, N4602);
  not ginst1084 (N5106, N4611);
  nand ginst1085 (N5107, N2709, N4611);
  not ginst1086 (N5108, N4614);
  nand ginst1087 (N5109, N2710, N4614);
  not ginst1088 (N5110, N4617);
  nand ginst1089 (N5111, N2711, N4617);
  nand ginst1090 (N5112, N1890, N4855);
  not ginst1091 (N5113, N4621);
  nand ginst1092 (N5114, N2713, N4621);
  not ginst1093 (N5115, N4624);
  nand ginst1094 (N5116, N2714, N4624);
  and ginst1095 (N5117, N4364, N4379);
  and ginst1096 (N5118, N4364, N4379);
  and ginst1097 (N5119, N54, N4405);
  not ginst1098 (N5120, N4627);
  nand ginst1099 (N5121, N2716, N4630);
  not ginst1100 (N5122, N4630);
  nand ginst1101 (N5123, N2717, N4633);
  not ginst1102 (N5124, N4633);
  nand ginst1103 (N5125, N1908, N4909);
  nand ginst1104 (N5126, N2719, N4637);
  not ginst1105 (N5127, N4637);
  nand ginst1106 (N5128, N2720, N4640);
  not ginst1107 (N5129, N4640);
  nand ginst1108 (N5130, N2721, N4643);
  not ginst1109 (N5131, N4643);
  and ginst1110 (N5132, N4425, N4440);
  and ginst1111 (N5133, N4425, N4440);
  not ginst1112 (N5135, N4649);
  not ginst1113 (N5136, N4652);
  nand ginst1114 (N5137, N4521, N4655);
  not ginst1115 (N5138, N4655);
  not ginst1116 (N5139, N4658);
  nand ginst1117 (N5140, N4658, N4947);
  not ginst1118 (N5141, N4674);
  not ginst1119 (N5142, N4677);
  not ginst1120 (N5143, N4680);
  not ginst1121 (N5144, N4683);
  nand ginst1122 (N5145, N4523, N4686);
  not ginst1123 (N5146, N4686);
  nor ginst1124 (N5147, N4196, N4953);
  nor ginst1125 (N5148, N4954, N4955);
  not ginst1126 (N5150, N4524);
  nand ginst1127 (N5153, N4228, N4965);
  nand ginst1128 (N5154, N4225, N4966);
  nand ginst1129 (N5155, N4234, N4967);
  nand ginst1130 (N5156, N4231, N4968);
  not ginst1131 (N5157, N4532);
  nand ginst1132 (N5160, N4249, N4972);
  nand ginst1133 (N5161, N4246, N4973);
  nand ginst1134 (N5162, N3816, N4974);
  and ginst1135 (N5163, N3793, N4200, N4976);
  and ginst1136 (N5164, N3789, N4203, N4977);
  and ginst1137 (N5165, N3147, N3158, N4942);
  not ginst1138 (N5166, N4512);
  buf ginst1139 (N5169, N4290);
  not ginst1140 (N5172, N4605);
  buf ginst1141 (N5173, N4325);
  not ginst1142 (N5176, N4608);
  buf ginst1143 (N5177, N4349);
  buf ginst1144 (N5180, N4405);
  buf ginst1145 (N5183, N4357);
  buf ginst1146 (N5186, N4357);
  buf ginst1147 (N5189, N4364);
  buf ginst1148 (N5192, N4364);
  buf ginst1149 (N5195, N4385);
  not ginst1150 (N5198, N4646);
  buf ginst1151 (N5199, N4418);
  buf ginst1152 (N5202, N4425);
  buf ginst1153 (N5205, N4445);
  buf ginst1154 (N5208, N4418);
  buf ginst1155 (N5211, N4425);
  buf ginst1156 (N5214, N4477);
  buf ginst1157 (N5217, N4469);
  buf ginst1158 (N5220, N4477);
  not ginst1159 (N5223, N4662);
  not ginst1160 (N5224, N4665);
  not ginst1161 (N5225, N4668);
  not ginst1162 (N5226, N4671);
  not ginst1163 (N5227, N4689);
  not ginst1164 (N5228, N4692);
  not ginst1165 (N5229, N4695);
  not ginst1166 (N5230, N4698);
  nand ginst1167 (N5232, N4240, N5052);
  nand ginst1168 (N5233, N4237, N5053);
  nand ginst1169 (N5234, N4258, N5055);
  nand ginst1170 (N5235, N4255, N5056);
  nand ginst1171 (N5236, N4721, N5057);
  nand ginst1172 (N5239, N3824, N5058);
  and ginst1173 (N5240, N4270, N5060, N5061);
  not ginst1174 (N5241, N4939);
  nand ginst1175 (N5242, N1824, N5069);
  nand ginst1176 (N5243, N1827, N5071);
  nand ginst1177 (N5244, N1830, N5073);
  nand ginst1178 (N5245, N1833, N5075);
  nand ginst1179 (N5246, N1836, N5077);
  nand ginst1180 (N5247, N1839, N5079);
  nand ginst1181 (N5248, N1842, N5081);
  nand ginst1182 (N5249, N1845, N5083);
  nand ginst1183 (N5250, N1848, N5085);
  nand ginst1184 (N5252, N1854, N5089);
  nand ginst1185 (N5253, N1857, N5091);
  nand ginst1186 (N5254, N1860, N5093);
  nand ginst1187 (N5255, N1863, N5095);
  nand ginst1188 (N5256, N1866, N5097);
  nand ginst1189 (N5257, N1869, N5099);
  nand ginst1190 (N5258, N1872, N5101);
  nand ginst1191 (N5259, N1875, N5103);
  nand ginst1192 (N5260, N1878, N5105);
  nand ginst1193 (N5261, N1881, N5106);
  nand ginst1194 (N5262, N1884, N5108);
  nand ginst1195 (N5263, N1887, N5110);
  nand ginst1196 (N5264, N4856, N5112);
  nand ginst1197 (N5274, N1893, N5113);
  nand ginst1198 (N5275, N1896, N5115);
  nand ginst1199 (N5282, N1902, N5122);
  nand ginst1200 (N5283, N1905, N5124);
  nand ginst1201 (N5284, N4908, N5125);
  nand ginst1202 (N5298, N1911, N5127);
  nand ginst1203 (N5299, N1914, N5129);
  nand ginst1204 (N5300, N1917, N5131);
  nand ginst1205 (N5303, N4652, N5135);
  nand ginst1206 (N5304, N4649, N5136);
  nand ginst1207 (N5305, N4008, N5138);
  nand ginst1208 (N5306, N4219, N5139);
  nand ginst1209 (N5307, N4677, N5141);
  nand ginst1210 (N5308, N4674, N5142);
  nand ginst1211 (N5309, N4683, N5143);
  nand ginst1212 (N5310, N4680, N5144);
  nand ginst1213 (N5311, N4011, N5146);
  not ginst1214 (N5312, N5049);
  nand ginst1215 (N5315, N5153, N5154);
  nand ginst1216 (N5319, N5155, N5156);
  nand ginst1217 (N5324, N5160, N5161);
  nand ginst1218 (N5328, N4975, N5162);
  nor ginst1219 (N5331, N4978, N5163);
  nor ginst1220 (N5332, N4979, N5164);
  or ginst1221 (N5346, N4412, N5119);
  nand ginst1222 (N5363, N4665, N5223);
  nand ginst1223 (N5364, N4662, N5224);
  nand ginst1224 (N5365, N4671, N5225);
  nand ginst1225 (N5366, N4668, N5226);
  nand ginst1226 (N5367, N4692, N5227);
  nand ginst1227 (N5368, N4689, N5228);
  nand ginst1228 (N5369, N4698, N5229);
  nand ginst1229 (N5370, N4695, N5230);
  nand ginst1230 (N5371, N5147, N5148);
  buf ginst1231 (N5374, N4939);
  nand ginst1232 (N5377, N5232, N5233);
  nand ginst1233 (N5382, N5234, N5235);
  nand ginst1234 (N5385, N5059, N5239);
  and ginst1235 (N5388, N5062, N5063, N5241);
  nand ginst1236 (N5389, N5070, N5242);
  nand ginst1237 (N5396, N5072, N5243);
  nand ginst1238 (N5407, N5074, N5244);
  nand ginst1239 (N5418, N5076, N5245);
  nand ginst1240 (N5424, N5078, N5246);
  nand ginst1241 (N5431, N5080, N5247);
  nand ginst1242 (N5441, N5082, N5248);
  nand ginst1243 (N5452, N5084, N5249);
  nand ginst1244 (N5462, N5086, N5250);
  not ginst1245 (N5469, N5169);
  nand ginst1246 (N5470, N5088, N5252);
  nand ginst1247 (N5477, N5090, N5253);
  nand ginst1248 (N5488, N5092, N5254);
  nand ginst1249 (N5498, N5094, N5255);
  nand ginst1250 (N5506, N5096, N5256);
  nand ginst1251 (N5520, N5098, N5257);
  nand ginst1252 (N5536, N5100, N5258);
  nand ginst1253 (N5549, N5102, N5259);
  nand ginst1254 (N5555, N5104, N5260);
  nand ginst1255 (N5562, N5107, N5261);
  nand ginst1256 (N5573, N5109, N5262);
  nand ginst1257 (N5579, N5111, N5263);
  nand ginst1258 (N5595, N5114, N5274);
  nand ginst1259 (N5606, N5116, N5275);
  nand ginst1260 (N5616, N2715, N5180);
  not ginst1261 (N5617, N5180);
  not ginst1262 (N5618, N5183);
  not ginst1263 (N5619, N5186);
  not ginst1264 (N5620, N5189);
  not ginst1265 (N5621, N5192);
  not ginst1266 (N5622, N5195);
  nand ginst1267 (N5624, N5121, N5282);
  nand ginst1268 (N5634, N5123, N5283);
  nand ginst1269 (N5655, N5126, N5298);
  nand ginst1270 (N5671, N5128, N5299);
  nand ginst1271 (N5684, N5130, N5300);
  not ginst1272 (N5690, N5202);
  not ginst1273 (N5691, N5211);
  nand ginst1274 (N5692, N5303, N5304);
  nand ginst1275 (N5696, N5137, N5305);
  nand ginst1276 (N5700, N5140, N5306);
  nand ginst1277 (N5703, N5307, N5308);
  nand ginst1278 (N5707, N5309, N5310);
  nand ginst1279 (N5711, N5145, N5311);
  and ginst1280 (N5726, N4512, N5166);
  not ginst1281 (N5727, N5173);
  not ginst1282 (N5728, N5177);
  not ginst1283 (N5730, N5199);
  not ginst1284 (N5731, N5205);
  not ginst1285 (N5732, N5208);
  not ginst1286 (N5733, N5214);
  not ginst1287 (N5734, N5217);
  not ginst1288 (N5735, N5220);
  nand ginst1289 (N5736, N5365, N5366);
  nand ginst1290 (N5739, N5363, N5364);
  nand ginst1291 (N5742, N5369, N5370);
  nand ginst1292 (N5745, N5367, N5368);
  not ginst1293 (N5755, N5236);
  nand ginst1294 (N5756, N5331, N5332);
  and ginst1295 (N5954, N4396, N5264);
  nand ginst1296 (N5955, N1899, N5617);
  not ginst1297 (N5956, N5346);
  and ginst1298 (N6005, N4456, N5284);
  and ginst1299 (N6006, N4456, N5284);
  not ginst1300 (N6023, N5371);
  nand ginst1301 (N6024, N5312, N5371);
  not ginst1302 (N6025, N5315);
  not ginst1303 (N6028, N5324);
  buf ginst1304 (N6031, N5319);
  buf ginst1305 (N6034, N5319);
  buf ginst1306 (N6037, N5328);
  buf ginst1307 (N6040, N5328);
  not ginst1308 (N6044, N5385);
  or ginst1309 (N6045, N5166, N5726);
  buf ginst1310 (N6048, N5264);
  buf ginst1311 (N6051, N5284);
  buf ginst1312 (N6054, N5284);
  not ginst1313 (N6065, N5374);
  nand ginst1314 (N6066, N5054, N5374);
  not ginst1315 (N6067, N5377);
  not ginst1316 (N6068, N5382);
  nand ginst1317 (N6069, N5382, N5755);
  and ginst1318 (N6071, N4316, N5470);
  and ginst1319 (N6072, N4320, N5470, N5477);
  and ginst1320 (N6073, N4325, N5470, N5477, N5488);
  and ginst1321 (N6074, N4357, N4364, N4385, N5562);
  and ginst1322 (N6075, N4280, N5389);
  and ginst1323 (N6076, N4284, N5389, N5396);
  and ginst1324 (N6077, N4290, N5389, N5396, N5407);
  and ginst1325 (N6078, N4418, N4425, N4445, N5624);
  not ginst1326 (N6079, N5418);
  and ginst1327 (N6080, N5389, N5396, N5407, N5418);
  and ginst1328 (N6083, N4284, N5396);
  and ginst1329 (N6084, N4290, N5396, N5407);
  and ginst1330 (N6085, N5396, N5407, N5418);
  and ginst1331 (N6086, N4284, N5396);
  and ginst1332 (N6087, N4290, N5396, N5407);
  and ginst1333 (N6088, N4290, N5407);
  and ginst1334 (N6089, N5407, N5418);
  and ginst1335 (N6090, N4290, N5407);
  and ginst1336 (N6091, N5424, N5431, N5441, N5452, N5462);
  and ginst1337 (N6094, N4298, N5424);
  and ginst1338 (N6095, N4301, N5424, N5431);
  and ginst1339 (N6096, N4305, N5424, N5431, N5441);
  and ginst1340 (N6097, N4310, N5424, N5431, N5441, N5452);
  and ginst1341 (N6098, N4301, N5431);
  and ginst1342 (N6099, N4305, N5431, N5441);
  and ginst1343 (N6100, N4310, N5431, N5441, N5452);
  and ginst1344 (N6101, N4, N5431, N5441, N5452, N5462);
  and ginst1345 (N6102, N4305, N5441);
  and ginst1346 (N6103, N4310, N5441, N5452);
  and ginst1347 (N6104, N4, N5441, N5452, N5462);
  and ginst1348 (N6105, N4310, N5452);
  and ginst1349 (N6106, N4, N5452, N5462);
  and ginst1350 (N6107, N4, N5462);
  and ginst1351 (N6108, N5470, N5477, N5488, N5549);
  and ginst1352 (N6111, N4320, N5477);
  and ginst1353 (N6112, N4325, N5477, N5488);
  and ginst1354 (N6113, N5477, N5488, N5549);
  and ginst1355 (N6114, N4320, N5477);
  and ginst1356 (N6115, N4325, N5477, N5488);
  and ginst1357 (N6116, N4325, N5488);
  and ginst1358 (N6117, N5498, N5506, N5520, N5536, N5555);
  and ginst1359 (N6120, N4332, N5498);
  and ginst1360 (N6121, N4336, N5498, N5506);
  and ginst1361 (N6122, N4342, N5498, N5506, N5520);
  and ginst1362 (N6123, N4349, N5498, N5506, N5520, N5536);
  and ginst1363 (N6124, N4336, N5506);
  and ginst1364 (N6125, N4342, N5506, N5520);
  and ginst1365 (N6126, N4349, N5506, N5520, N5536);
  and ginst1366 (N6127, N5506, N5520, N5536, N5555);
  and ginst1367 (N6128, N4336, N5506);
  and ginst1368 (N6129, N4342, N5506, N5520);
  and ginst1369 (N6130, N4349, N5506, N5520, N5536);
  and ginst1370 (N6131, N4342, N5520);
  and ginst1371 (N6132, N4349, N5520, N5536);
  and ginst1372 (N6133, N5520, N5536, N5555);
  and ginst1373 (N6134, N4342, N5520);
  and ginst1374 (N6135, N4349, N5520, N5536);
  and ginst1375 (N6136, N4349, N5536);
  and ginst1376 (N6137, N5488, N5549);
  and ginst1377 (N6138, N5536, N5555);
  not ginst1378 (N6139, N5573);
  and ginst1379 (N6140, N4357, N4364, N5562, N5573);
  and ginst1380 (N6143, N4364, N4385, N5562);
  and ginst1381 (N6144, N4364, N5562, N5573);
  and ginst1382 (N6145, N4364, N4385, N5562);
  and ginst1383 (N6146, N4385, N5562);
  and ginst1384 (N6147, N5562, N5573);
  and ginst1385 (N6148, N4385, N5562);
  and ginst1386 (N6149, N4405, N5264, N5579, N5595, N5606);
  and ginst1387 (N6152, N4067, N5579);
  and ginst1388 (N6153, N4396, N5264, N5579);
  and ginst1389 (N6154, N4400, N5264, N5579, N5595);
  and ginst1390 (N6155, N4412, N5264, N5579, N5595, N5606);
  and ginst1391 (N6156, N4400, N5264, N5595);
  and ginst1392 (N6157, N4412, N5264, N5595, N5606);
  and ginst1393 (N6158, N54, N4405, N5264, N5595, N5606);
  and ginst1394 (N6159, N4400, N5595);
  and ginst1395 (N6160, N4412, N5595, N5606);
  and ginst1396 (N6161, N54, N4405, N5595, N5606);
  and ginst1397 (N6162, N4412, N5606);
  and ginst1398 (N6163, N54, N4405, N5606);
  nand ginst1399 (N6164, N5616, N5955);
  and ginst1400 (N6168, N4418, N4425, N5624, N5684);
  and ginst1401 (N6171, N4425, N4445, N5624);
  and ginst1402 (N6172, N4425, N5624, N5684);
  and ginst1403 (N6173, N4425, N4445, N5624);
  and ginst1404 (N6174, N4445, N5624);
  and ginst1405 (N6175, N4477, N5284, N5634, N5655, N5671);
  and ginst1406 (N6178, N4080, N5634);
  and ginst1407 (N6179, N4456, N5284, N5634);
  and ginst1408 (N6180, N4462, N5284, N5634, N5655);
  and ginst1409 (N6181, N4469, N5284, N5634, N5655, N5671);
  and ginst1410 (N6182, N4462, N5284, N5655);
  and ginst1411 (N6183, N4469, N5284, N5655, N5671);
  and ginst1412 (N6184, N4477, N5284, N5655, N5671);
  and ginst1413 (N6185, N4462, N5284, N5655);
  and ginst1414 (N6186, N4469, N5284, N5655, N5671);
  and ginst1415 (N6187, N4462, N5655);
  and ginst1416 (N6188, N4469, N5655, N5671);
  and ginst1417 (N6189, N4477, N5655, N5671);
  and ginst1418 (N6190, N4462, N5655);
  and ginst1419 (N6191, N4469, N5655, N5671);
  and ginst1420 (N6192, N4469, N5671);
  and ginst1421 (N6193, N5624, N5684);
  and ginst1422 (N6194, N4477, N5671);
  not ginst1423 (N6197, N5692);
  not ginst1424 (N6200, N5696);
  not ginst1425 (N6203, N5703);
  not ginst1426 (N6206, N5707);
  buf ginst1427 (N6209, N5700);
  buf ginst1428 (N6212, N5700);
  buf ginst1429 (N6215, N5711);
  buf ginst1430 (N6218, N5711);
  nand ginst1431 (N6221, N5049, N6023);
  not ginst1432 (N6234, N5756);
  nand ginst1433 (N6235, N5756, N6044);
  buf ginst1434 (N6238, N5462);
  buf ginst1435 (N6241, N5389);
  buf ginst1436 (N6244, N5389);
  buf ginst1437 (N6247, N5396);
  buf ginst1438 (N6250, N5396);
  buf ginst1439 (N6253, N5407);
  buf ginst1440 (N6256, N5407);
  buf ginst1441 (N6259, N5424);
  buf ginst1442 (N6262, N5431);
  buf ginst1443 (N6265, N5441);
  buf ginst1444 (N6268, N5452);
  buf ginst1445 (N6271, N5549);
  buf ginst1446 (N6274, N5488);
  buf ginst1447 (N6277, N5470);
  buf ginst1448 (N6280, N5477);
  buf ginst1449 (N6283, N5549);
  buf ginst1450 (N6286, N5488);
  buf ginst1451 (N6289, N5470);
  buf ginst1452 (N6292, N5477);
  buf ginst1453 (N6295, N5555);
  buf ginst1454 (N6298, N5536);
  buf ginst1455 (N6301, N5498);
  buf ginst1456 (N6304, N5520);
  buf ginst1457 (N6307, N5506);
  buf ginst1458 (N6310, N5506);
  buf ginst1459 (N6313, N5555);
  buf ginst1460 (N6316, N5536);
  buf ginst1461 (N6319, N5498);
  buf ginst1462 (N6322, N5520);
  buf ginst1463 (N6325, N5562);
  buf ginst1464 (N6328, N5562);
  buf ginst1465 (N6331, N5579);
  buf ginst1466 (N6335, N5595);
  buf ginst1467 (N6338, N5606);
  buf ginst1468 (N6341, N5684);
  buf ginst1469 (N6344, N5624);
  buf ginst1470 (N6347, N5684);
  buf ginst1471 (N6350, N5624);
  buf ginst1472 (N6353, N5671);
  buf ginst1473 (N6356, N5634);
  buf ginst1474 (N6359, N5655);
  buf ginst1475 (N6364, N5671);
  buf ginst1476 (N6367, N5634);
  buf ginst1477 (N6370, N5655);
  not ginst1478 (N6373, N5736);
  not ginst1479 (N6374, N5739);
  not ginst1480 (N6375, N5742);
  not ginst1481 (N6376, N5745);
  nand ginst1482 (N6377, N4243, N6065);
  nand ginst1483 (N6378, N5236, N6068);
  or ginst1484 (N6382, N4268, N6071, N6072, N6073);
  or ginst1485 (N6386, N3968, N5065, N5066, N6074);
  or ginst1486 (N6388, N4271, N6075, N6076, N6077);
  or ginst1487 (N6392, N3968, N5067, N5068, N6078);
  or ginst1488 (N6397, N4297, N6094, N6095, N6096, N6097);
  or ginst1489 (N6411, N4320, N6116);
  or ginst1490 (N6415, N4331, N6120, N6121, N6122, N6123);
  or ginst1491 (N6419, N4342, N6136);
  or ginst1492 (N6427, N4392, N6152, N6153, N6154, N6155);
  not ginst1493 (N6434, N6048);
  or ginst1494 (N6437, N4440, N6174);
  or ginst1495 (N6441, N4451, N6178, N6179, N6180, N6181);
  or ginst1496 (N6445, N4462, N6192);
  not ginst1497 (N6448, N6051);
  not ginst1498 (N6449, N6054);
  nand ginst1499 (N6466, N6024, N6221);
  not ginst1500 (N6469, N6031);
  not ginst1501 (N6470, N6034);
  not ginst1502 (N6471, N6037);
  not ginst1503 (N6472, N6040);
  and ginst1504 (N6473, N4524, N5315, N6031);
  and ginst1505 (N6474, N5150, N6025, N6034);
  and ginst1506 (N6475, N4532, N5324, N6037);
  and ginst1507 (N6476, N5157, N6028, N6040);
  nand ginst1508 (N6477, N5385, N6234);
  nand ginst1509 (N6478, N132, N6045);
  or ginst1510 (N6482, N4280, N6083, N6084, N6085);
  nor ginst1511 (N6486, N4280, N6086, N6087);
  or ginst1512 (N6490, N4284, N6088, N6089);
  nor ginst1513 (N6494, N4284, N6090);
  or ginst1514 (N6500, N4298, N6098, N6099, N6100, N6101);
  or ginst1515 (N6504, N4301, N6102, N6103, N6104);
  or ginst1516 (N6508, N4305, N6105, N6106);
  or ginst1517 (N6512, N4310, N6107);
  or ginst1518 (N6516, N4316, N6111, N6112, N6113);
  nor ginst1519 (N6526, N4316, N6114, N6115);
  or ginst1520 (N6536, N4336, N6131, N6132, N6133);
  or ginst1521 (N6539, N4332, N6124, N6125, N6126, N6127);
  nor ginst1522 (N6553, N4336, N6134, N6135);
  nor ginst1523 (N6556, N4332, N6128, N6129, N6130);
  or ginst1524 (N6566, N4375, N5117, N6143, N6144);
  nor ginst1525 (N6569, N4375, N5118, N6145);
  or ginst1526 (N6572, N4379, N6146, N6147);
  nor ginst1527 (N6575, N4379, N6148);
  or ginst1528 (N6580, N4067, N5954, N6156, N6157, N6158);
  or ginst1529 (N6584, N4396, N6159, N6160, N6161);
  or ginst1530 (N6587, N4400, N6162, N6163);
  or ginst1531 (N6592, N4436, N5132, N6171, N6172);
  nor ginst1532 (N6599, N4436, N5133, N6173);
  or ginst1533 (N6606, N4456, N6187, N6188, N6189);
  or ginst1534 (N6609, N4080, N6005, N6182, N6183, N6184);
  nor ginst1535 (N6619, N4456, N6190, N6191);
  nor ginst1536 (N6622, N4080, N6006, N6185, N6186);
  nand ginst1537 (N6630, N5739, N6373);
  nand ginst1538 (N6631, N5736, N6374);
  nand ginst1539 (N6632, N5745, N6375);
  nand ginst1540 (N6633, N5742, N6376);
  nand ginst1541 (N6634, N6066, N6377);
  nand ginst1542 (N6637, N6069, N6378);
  not ginst1543 (N6640, N6164);
  and ginst1544 (N6641, N6108, N6117);
  and ginst1545 (N6643, N6140, N6149);
  and ginst1546 (N6646, N6168, N6175);
  and ginst1547 (N6648, N6080, N6091);
  nand ginst1548 (N6650, N2637, N6238);
  not ginst1549 (N6651, N6238);
  not ginst1550 (N6653, N6241);
  not ginst1551 (N6655, N6244);
  not ginst1552 (N6657, N6247);
  not ginst1553 (N6659, N6250);
  nand ginst1554 (N6660, N5087, N6253);
  not ginst1555 (N6661, N6253);
  nand ginst1556 (N6662, N5469, N6256);
  not ginst1557 (N6663, N6256);
  and ginst1558 (N6664, N4, N6091);
  not ginst1559 (N6666, N6259);
  not ginst1560 (N6668, N6262);
  not ginst1561 (N6670, N6265);
  not ginst1562 (N6672, N6268);
  not ginst1563 (N6675, N6117);
  not ginst1564 (N6680, N6280);
  not ginst1565 (N6681, N6292);
  not ginst1566 (N6682, N6307);
  not ginst1567 (N6683, N6310);
  nand ginst1568 (N6689, N5120, N6325);
  not ginst1569 (N6690, N6325);
  nand ginst1570 (N6691, N5622, N6328);
  not ginst1571 (N6692, N6328);
  and ginst1572 (N6693, N54, N6149);
  not ginst1573 (N6695, N6331);
  not ginst1574 (N6698, N6335);
  nand ginst1575 (N6699, N5956, N6338);
  not ginst1576 (N6700, N6338);
  not ginst1577 (N6703, N6175);
  not ginst1578 (N6708, N6209);
  not ginst1579 (N6709, N6212);
  not ginst1580 (N6710, N6215);
  not ginst1581 (N6711, N6218);
  and ginst1582 (N6712, N5692, N5696, N6209);
  and ginst1583 (N6713, N6197, N6200, N6212);
  and ginst1584 (N6714, N5703, N5707, N6215);
  and ginst1585 (N6715, N6203, N6206, N6218);
  buf ginst1586 (N6716, N6466);
  and ginst1587 (N6718, N1777, N3130, N6164);
  and ginst1588 (N6719, N5150, N5315, N6469);
  and ginst1589 (N6720, N4524, N6025, N6470);
  and ginst1590 (N6721, N5157, N5324, N6471);
  and ginst1591 (N6722, N4532, N6028, N6472);
  nand ginst1592 (N6724, N6235, N6477);
  not ginst1593 (N6739, N6271);
  not ginst1594 (N6740, N6274);
  not ginst1595 (N6741, N6277);
  not ginst1596 (N6744, N6283);
  not ginst1597 (N6745, N6286);
  not ginst1598 (N6746, N6289);
  not ginst1599 (N6751, N6295);
  not ginst1600 (N6752, N6298);
  not ginst1601 (N6753, N6301);
  not ginst1602 (N6754, N6304);
  not ginst1603 (N6755, N6322);
  not ginst1604 (N6760, N6313);
  not ginst1605 (N6761, N6316);
  not ginst1606 (N6762, N6319);
  not ginst1607 (N6772, N6341);
  not ginst1608 (N6773, N6344);
  not ginst1609 (N6776, N6347);
  not ginst1610 (N6777, N6350);
  not ginst1611 (N6782, N6353);
  not ginst1612 (N6783, N6356);
  not ginst1613 (N6784, N6359);
  not ginst1614 (N6785, N6370);
  not ginst1615 (N6790, N6364);
  not ginst1616 (N6791, N6367);
  nand ginst1617 (N6792, N6630, N6631);
  nand ginst1618 (N6795, N6632, N6633);
  and ginst1619 (N6801, N6108, N6415);
  and ginst1620 (N6802, N6140, N6427);
  and ginst1621 (N6803, N6080, N6397);
  and ginst1622 (N6804, N6168, N6441);
  not ginst1623 (N6805, N6466);
  nand ginst1624 (N6806, N1851, N6651);
  not ginst1625 (N6807, N6482);
  nand ginst1626 (N6808, N6482, N6653);
  not ginst1627 (N6809, N6486);
  nand ginst1628 (N6810, N6486, N6655);
  not ginst1629 (N6811, N6490);
  nand ginst1630 (N6812, N6490, N6657);
  not ginst1631 (N6813, N6494);
  nand ginst1632 (N6814, N6494, N6659);
  nand ginst1633 (N6815, N4575, N6661);
  nand ginst1634 (N6816, N5169, N6663);
  or ginst1635 (N6817, N6397, N6664);
  not ginst1636 (N6823, N6500);
  nand ginst1637 (N6824, N6500, N6666);
  not ginst1638 (N6825, N6504);
  nand ginst1639 (N6826, N6504, N6668);
  not ginst1640 (N6827, N6508);
  nand ginst1641 (N6828, N6508, N6670);
  not ginst1642 (N6829, N6512);
  nand ginst1643 (N6830, N6512, N6672);
  not ginst1644 (N6831, N6415);
  not ginst1645 (N6834, N6566);
  nand ginst1646 (N6835, N5618, N6566);
  not ginst1647 (N6836, N6569);
  nand ginst1648 (N6837, N5619, N6569);
  not ginst1649 (N6838, N6572);
  nand ginst1650 (N6839, N5620, N6572);
  not ginst1651 (N6840, N6575);
  nand ginst1652 (N6841, N5621, N6575);
  nand ginst1653 (N6842, N4627, N6690);
  nand ginst1654 (N6843, N5195, N6692);
  or ginst1655 (N6844, N6427, N6693);
  not ginst1656 (N6850, N6580);
  nand ginst1657 (N6851, N6580, N6695);
  not ginst1658 (N6852, N6584);
  nand ginst1659 (N6853, N6434, N6584);
  not ginst1660 (N6854, N6587);
  nand ginst1661 (N6855, N6587, N6698);
  nand ginst1662 (N6856, N5346, N6700);
  not ginst1663 (N6857, N6441);
  and ginst1664 (N6860, N5696, N6197, N6708);
  and ginst1665 (N6861, N5692, N6200, N6709);
  and ginst1666 (N6862, N5707, N6203, N6710);
  and ginst1667 (N6863, N5703, N6206, N6711);
  or ginst1668 (N6866, N3785, N4197, N6718);
  nor ginst1669 (N6872, N6473, N6719);
  nor ginst1670 (N6873, N6474, N6720);
  nor ginst1671 (N6874, N6475, N6721);
  nor ginst1672 (N6875, N6476, N6722);
  not ginst1673 (N6876, N6637);
  buf ginst1674 (N6877, N6724);
  and ginst1675 (N6879, N6045, N6478);
  and ginst1676 (N6880, N132, N6478);
  or ginst1677 (N6881, N6137, N6411);
  not ginst1678 (N6884, N6516);
  not ginst1679 (N6885, N6411);
  not ginst1680 (N6888, N6526);
  not ginst1681 (N6889, N6536);
  nand ginst1682 (N6890, N5176, N6536);
  or ginst1683 (N6891, N6138, N6419);
  not ginst1684 (N6894, N6539);
  not ginst1685 (N6895, N6553);
  nand ginst1686 (N6896, N5728, N6553);
  not ginst1687 (N6897, N6419);
  not ginst1688 (N6900, N6556);
  or ginst1689 (N6901, N6193, N6437);
  not ginst1690 (N6904, N6592);
  not ginst1691 (N6905, N6437);
  not ginst1692 (N6908, N6599);
  or ginst1693 (N6909, N6194, N6445);
  not ginst1694 (N6912, N6606);
  not ginst1695 (N6913, N6609);
  not ginst1696 (N6914, N6619);
  nand ginst1697 (N6915, N5734, N6619);
  not ginst1698 (N6916, N6445);
  not ginst1699 (N6919, N6622);
  not ginst1700 (N6922, N6634);
  nand ginst1701 (N6923, N6067, N6634);
  or ginst1702 (N6924, N6382, N6801);
  or ginst1703 (N6925, N6386, N6802);
  or ginst1704 (N6926, N6388, N6803);
  or ginst1705 (N6927, N6392, N6804);
  not ginst1706 (N6930, N6724);
  nand ginst1707 (N6932, N6650, N6806);
  nand ginst1708 (N6935, N6241, N6807);
  nand ginst1709 (N6936, N6244, N6809);
  nand ginst1710 (N6937, N6247, N6811);
  nand ginst1711 (N6938, N6250, N6813);
  nand ginst1712 (N6939, N6660, N6815);
  nand ginst1713 (N6940, N6662, N6816);
  nand ginst1714 (N6946, N6259, N6823);
  nand ginst1715 (N6947, N6262, N6825);
  nand ginst1716 (N6948, N6265, N6827);
  nand ginst1717 (N6949, N6268, N6829);
  nand ginst1718 (N6953, N5183, N6834);
  nand ginst1719 (N6954, N5186, N6836);
  nand ginst1720 (N6955, N5189, N6838);
  nand ginst1721 (N6956, N5192, N6840);
  nand ginst1722 (N6957, N6689, N6842);
  nand ginst1723 (N6958, N6691, N6843);
  nand ginst1724 (N6964, N6331, N6850);
  nand ginst1725 (N6965, N6048, N6852);
  nand ginst1726 (N6966, N6335, N6854);
  nand ginst1727 (N6967, N6699, N6856);
  nor ginst1728 (N6973, N6712, N6860);
  nor ginst1729 (N6974, N6713, N6861);
  nor ginst1730 (N6975, N6714, N6862);
  nor ginst1731 (N6976, N6715, N6863);
  not ginst1732 (N6977, N6792);
  not ginst1733 (N6978, N6795);
  or ginst1734 (N6979, N6879, N6880);
  nand ginst1735 (N6987, N4608, N6889);
  nand ginst1736 (N6990, N5177, N6895);
  nand ginst1737 (N6999, N5217, N6914);
  nand ginst1738 (N7002, N5377, N6922);
  nand ginst1739 (N7003, N6872, N6873);
  nand ginst1740 (N7006, N6874, N6875);
  and ginst1741 (N7011, N2681, N2692, N6866);
  and ginst1742 (N7012, N2756, N2767, N6866);
  and ginst1743 (N7013, N2779, N2790, N6866);
  not ginst1744 (N7015, N6866);
  and ginst1745 (N7016, N2801, N2812, N6866);
  nand ginst1746 (N7018, N6808, N6935);
  nand ginst1747 (N7019, N6810, N6936);
  nand ginst1748 (N7020, N6812, N6937);
  nand ginst1749 (N7021, N6814, N6938);
  not ginst1750 (N7022, N6939);
  not ginst1751 (N7023, N6817);
  nand ginst1752 (N7028, N6824, N6946);
  nand ginst1753 (N7031, N6826, N6947);
  nand ginst1754 (N7034, N6828, N6948);
  nand ginst1755 (N7037, N6830, N6949);
  and ginst1756 (N7040, N6079, N6817);
  and ginst1757 (N7041, N6675, N6831);
  nand ginst1758 (N7044, N6835, N6953);
  nand ginst1759 (N7045, N6837, N6954);
  nand ginst1760 (N7046, N6839, N6955);
  nand ginst1761 (N7047, N6841, N6956);
  not ginst1762 (N7048, N6957);
  not ginst1763 (N7049, N6844);
  nand ginst1764 (N7054, N6851, N6964);
  nand ginst1765 (N7057, N6853, N6965);
  nand ginst1766 (N7060, N6855, N6966);
  and ginst1767 (N7064, N6139, N6844);
  and ginst1768 (N7065, N6703, N6857);
  not ginst1769 (N7072, N6881);
  nand ginst1770 (N7073, N5172, N6881);
  not ginst1771 (N7074, N6885);
  nand ginst1772 (N7075, N5727, N6885);
  nand ginst1773 (N7076, N6890, N6987);
  not ginst1774 (N7079, N6891);
  nand ginst1775 (N7080, N6896, N6990);
  not ginst1776 (N7083, N6897);
  not ginst1777 (N7084, N6901);
  nand ginst1778 (N7085, N5198, N6901);
  not ginst1779 (N7086, N6905);
  nand ginst1780 (N7087, N5731, N6905);
  not ginst1781 (N7088, N6909);
  nand ginst1782 (N7089, N6909, N6912);
  buf ginst1783 (N709, N141);
  nand ginst1784 (N7090, N6915, N6999);
  not ginst1785 (N7093, N6916);
  nand ginst1786 (N7094, N6973, N6974);
  nand ginst1787 (N7097, N6975, N6976);
  nand ginst1788 (N7101, N6923, N7002);
  not ginst1789 (N7105, N6932);
  not ginst1790 (N7110, N6967);
  and ginst1791 (N7114, N603, N1755, N6979);
  not ginst1792 (N7115, N7019);
  not ginst1793 (N7116, N7021);
  and ginst1794 (N7125, N6817, N7018);
  and ginst1795 (N7126, N6817, N7020);
  and ginst1796 (N7127, N6817, N7022);
  not ginst1797 (N7130, N7045);
  not ginst1798 (N7131, N7047);
  and ginst1799 (N7139, N6844, N7044);
  and ginst1800 (N7140, N6844, N7046);
  and ginst1801 (N7141, N6844, N7048);
  and ginst1802 (N7146, N1761, N3108, N6932);
  and ginst1803 (N7147, N1777, N3130, N6967);
  not ginst1804 (N7149, N7003);
  not ginst1805 (N7150, N7006);
  nand ginst1806 (N7151, N6876, N7006);
  nand ginst1807 (N7152, N4605, N7072);
  nand ginst1808 (N7153, N5173, N7074);
  nand ginst1809 (N7158, N4646, N7084);
  nand ginst1810 (N7159, N5205, N7086);
  nand ginst1811 (N7160, N6606, N7088);
  not ginst1812 (N7166, N7037);
  not ginst1813 (N7167, N7034);
  not ginst1814 (N7168, N7031);
  not ginst1815 (N7169, N7028);
  not ginst1816 (N7170, N7060);
  not ginst1817 (N7171, N7057);
  not ginst1818 (N7172, N7054);
  and ginst1819 (N7173, N7023, N7115);
  and ginst1820 (N7174, N7023, N7116);
  and ginst1821 (N7175, N6940, N7023);
  and ginst1822 (N7176, N5418, N7023);
  not ginst1823 (N7177, N7041);
  and ginst1824 (N7178, N7049, N7130);
  and ginst1825 (N7179, N7049, N7131);
  and ginst1826 (N7180, N6958, N7049);
  and ginst1827 (N7181, N5573, N7049);
  not ginst1828 (N7182, N7065);
  not ginst1829 (N7183, N7094);
  nand ginst1830 (N7184, N6977, N7094);
  not ginst1831 (N7185, N7097);
  nand ginst1832 (N7186, N6978, N7097);
  and ginst1833 (N7187, N1761, N3108, N7037);
  and ginst1834 (N7188, N1761, N3108, N7034);
  and ginst1835 (N7189, N1761, N3108, N7031);
  or ginst1836 (N7190, N3781, N4956, N7146);
  and ginst1837 (N7196, N1777, N3130, N7060);
  and ginst1838 (N7197, N1777, N3130, N7057);
  or ginst1839 (N7198, N3786, N4960, N7147);
  nand ginst1840 (N7204, N7101, N7149);
  not ginst1841 (N7205, N7101);
  nand ginst1842 (N7206, N6637, N7150);
  and ginst1843 (N7207, N1793, N3158, N7028);
  and ginst1844 (N7208, N1807, N3180, N7054);
  nand ginst1845 (N7209, N7073, N7152);
  nand ginst1846 (N7212, N7075, N7153);
  not ginst1847 (N7215, N7076);
  nand ginst1848 (N7216, N7076, N7079);
  not ginst1849 (N7217, N7080);
  nand ginst1850 (N7218, N7080, N7083);
  nand ginst1851 (N7219, N7085, N7158);
  nand ginst1852 (N7222, N7087, N7159);
  nand ginst1853 (N7225, N7089, N7160);
  not ginst1854 (N7228, N7090);
  nand ginst1855 (N7229, N7090, N7093);
  or ginst1856 (N7236, N7125, N7173);
  or ginst1857 (N7239, N7126, N7174);
  or ginst1858 (N7242, N7127, N7175);
  or ginst1859 (N7245, N7040, N7176);
  or ginst1860 (N7250, N7139, N7178);
  or ginst1861 (N7257, N7140, N7179);
  or ginst1862 (N7260, N7141, N7180);
  or ginst1863 (N7263, N7064, N7181);
  nand ginst1864 (N7268, N6792, N7183);
  nand ginst1865 (N7269, N6795, N7185);
  or ginst1866 (N7270, N3782, N4957, N7187);
  or ginst1867 (N7276, N3783, N4958, N7188);
  or ginst1868 (N7282, N3784, N4959, N7189);
  or ginst1869 (N7288, N3787, N4961, N7196);
  or ginst1870 (N7294, N3788, N3998, N7197);
  nand ginst1871 (N7300, N7003, N7205);
  nand ginst1872 (N7301, N7151, N7206);
  or ginst1873 (N7304, N3800, N4980, N7207);
  or ginst1874 (N7310, N3805, N4984, N7208);
  nand ginst1875 (N7320, N6891, N7215);
  nand ginst1876 (N7321, N6897, N7217);
  nand ginst1877 (N7328, N6916, N7228);
  and ginst1878 (N7338, N1185, N2692, N7190);
  and ginst1879 (N7339, N2681, N2692, N7198);
  and ginst1880 (N7340, N1247, N2767, N7190);
  and ginst1881 (N7341, N2756, N2767, N7198);
  and ginst1882 (N7342, N1327, N2790, N7190);
  and ginst1883 (N7349, N2779, N2790, N7198);
  and ginst1884 (N7357, N2801, N2812, N7198);
  not ginst1885 (N7363, N7198);
  and ginst1886 (N7364, N1351, N2812, N7190);
  not ginst1887 (N7365, N7190);
  nand ginst1888 (N7394, N7184, N7268);
  nand ginst1889 (N7397, N7186, N7269);
  nand ginst1890 (N7402, N7204, N7300);
  not ginst1891 (N7405, N7209);
  nand ginst1892 (N7406, N6884, N7209);
  not ginst1893 (N7407, N7212);
  nand ginst1894 (N7408, N6888, N7212);
  nand ginst1895 (N7409, N7216, N7320);
  nand ginst1896 (N7412, N7218, N7321);
  not ginst1897 (N7415, N7219);
  nand ginst1898 (N7416, N6904, N7219);
  not ginst1899 (N7417, N7222);
  nand ginst1900 (N7418, N6908, N7222);
  not ginst1901 (N7419, N7225);
  nand ginst1902 (N7420, N6913, N7225);
  nand ginst1903 (N7421, N7229, N7328);
  not ginst1904 (N7424, N7245);
  not ginst1905 (N7425, N7242);
  not ginst1906 (N7426, N7239);
  not ginst1907 (N7427, N7236);
  not ginst1908 (N7428, N7263);
  not ginst1909 (N7429, N7260);
  not ginst1910 (N7430, N7257);
  not ginst1911 (N7431, N7250);
  not ginst1912 (N7432, N7250);
  and ginst1913 (N7433, N2653, N2664, N7310);
  and ginst1914 (N7434, N1161, N2664, N7304);
  or ginst1915 (N7435, N2591, N3621, N7011, N7338);
  and ginst1916 (N7436, N1185, N2692, N7270);
  and ginst1917 (N7437, N2681, N2692, N7288);
  and ginst1918 (N7438, N1185, N2692, N7276);
  and ginst1919 (N7439, N2681, N2692, N7294);
  and ginst1920 (N7440, N1185, N2692, N7282);
  and ginst1921 (N7441, N2728, N2739, N7310);
  and ginst1922 (N7442, N1223, N2739, N7304);
  or ginst1923 (N7443, N2600, N3632, N7012, N7340);
  and ginst1924 (N7444, N1247, N2767, N7270);
  and ginst1925 (N7445, N2756, N2767, N7288);
  and ginst1926 (N7446, N1247, N2767, N7276);
  and ginst1927 (N7447, N2756, N2767, N7294);
  and ginst1928 (N7448, N1247, N2767, N7282);
  or ginst1929 (N7449, N2605, N3641, N7013, N7342);
  and ginst1930 (N7450, N3041, N3052, N7310);
  and ginst1931 (N7451, N1697, N3052, N7304);
  and ginst1932 (N7452, N2779, N2790, N7294);
  and ginst1933 (N7453, N1327, N2790, N7282);
  and ginst1934 (N7454, N2779, N2790, N7288);
  and ginst1935 (N7455, N1327, N2790, N7276);
  and ginst1936 (N7456, N1327, N2790, N7270);
  and ginst1937 (N7457, N3075, N3086, N7310);
  and ginst1938 (N7458, N1731, N3086, N7304);
  and ginst1939 (N7459, N2801, N2812, N7294);
  and ginst1940 (N7460, N1351, N2812, N7282);
  and ginst1941 (N7461, N2801, N2812, N7288);
  and ginst1942 (N7462, N1351, N2812, N7276);
  and ginst1943 (N7463, N1351, N2812, N7270);
  and ginst1944 (N7464, N599, N603, N7250);
  not ginst1945 (N7465, N7310);
  not ginst1946 (N7466, N7294);
  not ginst1947 (N7467, N7288);
  not ginst1948 (N7468, N7301);
  or ginst1949 (N7469, N2626, N3660, N7016, N7364);
  not ginst1950 (N7470, N7304);
  not ginst1951 (N7471, N7282);
  not ginst1952 (N7472, N7276);
  not ginst1953 (N7473, N7270);
  buf ginst1954 (N7474, N7394);
  buf ginst1955 (N7476, N7397);
  and ginst1956 (N7479, N3068, N7301);
  and ginst1957 (N7481, N1793, N3158, N7245);
  and ginst1958 (N7482, N1793, N3158, N7242);
  and ginst1959 (N7483, N1793, N3158, N7239);
  and ginst1960 (N7484, N1793, N3158, N7236);
  and ginst1961 (N7485, N1807, N3180, N7263);
  and ginst1962 (N7486, N1807, N3180, N7260);
  and ginst1963 (N7487, N1807, N3180, N7257);
  and ginst1964 (N7488, N1807, N3180, N7250);
  nand ginst1965 (N7489, N6979, N7250);
  nand ginst1966 (N7492, N6516, N7405);
  nand ginst1967 (N7493, N6526, N7407);
  nand ginst1968 (N7498, N6592, N7415);
  nand ginst1969 (N7499, N6599, N7417);
  nand ginst1970 (N7500, N6609, N7419);
  and ginst1971 (N7503, N7105, N7166, N7167, N7168, N7169, N7424, N7425, N7426, N7427);
  and ginst1972 (N7504, N6640, N7110, N7170, N7171, N7172, N7428, N7429, N7430, N7431);
  or ginst1973 (N7505, N2585, N3616, N7433, N7434);
  and ginst1974 (N7506, N2675, N7435);
  or ginst1975 (N7507, N2592, N3622, N7339, N7436);
  or ginst1976 (N7508, N2593, N3623, N7437, N7438);
  or ginst1977 (N7509, N2594, N3624, N7439, N7440);
  or ginst1978 (N7510, N2595, N3627, N7441, N7442);
  and ginst1979 (N7511, N2750, N7443);
  or ginst1980 (N7512, N2601, N3633, N7341, N7444);
  or ginst1981 (N7513, N2602, N3634, N7445, N7446);
  or ginst1982 (N7514, N2603, N3635, N7447, N7448);
  or ginst1983 (N7515, N2610, N3646, N7450, N7451);
  or ginst1984 (N7516, N2611, N3647, N7452, N7453);
  or ginst1985 (N7517, N2612, N3648, N7454, N7455);
  or ginst1986 (N7518, N2613, N3649, N7349, N7456);
  or ginst1987 (N7519, N2618, N3654, N7457, N7458);
  or ginst1988 (N7520, N2619, N3655, N7459, N7460);
  or ginst1989 (N7521, N2620, N3656, N7461, N7462);
  or ginst1990 (N7522, N2621, N3657, N7357, N7463);
  or ginst1991 (N7525, N2624, N4741, N7114, N7464);
  and ginst1992 (N7526, N3119, N3130, N7468);
  not ginst1993 (N7527, N7394);
  not ginst1994 (N7528, N7397);
  not ginst1995 (N7529, N7402);
  and ginst1996 (N7530, N3068, N7402);
  or ginst1997 (N7531, N3801, N4981, N7481);
  or ginst1998 (N7537, N3802, N4982, N7482);
  or ginst1999 (N7543, N3803, N4983, N7483);
  or ginst2000 (N7549, N3804, N5165, N7484);
  or ginst2001 (N7555, N3806, N4985, N7485);
  or ginst2002 (N7561, N3807, N4986, N7486);
  or ginst2003 (N7567, N3808, N4547, N7487);
  or ginst2004 (N7573, N3809, N4987, N7488);
  nand ginst2005 (N7579, N7406, N7492);
  nand ginst2006 (N7582, N7408, N7493);
  not ginst2007 (N7585, N7409);
  nand ginst2008 (N7586, N6894, N7409);
  not ginst2009 (N7587, N7412);
  nand ginst2010 (N7588, N6900, N7412);
  nand ginst2011 (N7589, N7416, N7498);
  nand ginst2012 (N7592, N7418, N7499);
  nand ginst2013 (N7595, N7420, N7500);
  not ginst2014 (N7598, N7421);
  nand ginst2015 (N7599, N6919, N7421);
  and ginst2016 (N7600, N2647, N7505);
  and ginst2017 (N7601, N2675, N7507);
  and ginst2018 (N7602, N2675, N7508);
  and ginst2019 (N7603, N2675, N7509);
  xor ginst2020 (N7604, N7604_in, flip_signal);
  and ginst2021 (N7604_in, N2722, N7510);
  and ginst2022 (N7605, N2750, N7512);
  and ginst2023 (N7606, N2750, N7513);
  and ginst2024 (N7607, N2750, N7514);
  and ginst2025 (N7624, N6979, N7489);
  and ginst2026 (N7625, N7250, N7489);
  and ginst2027 (N7626, N1149, N7525);
  and ginst2028 (N7631, N562, N6805, N6930, N7527, N7528);
  and ginst2029 (N7636, N3097, N3108, N7529);
  nand ginst2030 (N7657, N6539, N7585);
  nand ginst2031 (N7658, N6556, N7587);
  nand ginst2032 (N7665, N6622, N7598);
  and ginst2033 (N7666, N2653, N2664, N7555);
  and ginst2034 (N7667, N1161, N2664, N7531);
  and ginst2035 (N7668, N2653, N2664, N7561);
  and ginst2036 (N7669, N1161, N2664, N7537);
  and ginst2037 (N7670, N2653, N2664, N7567);
  and ginst2038 (N7671, N1161, N2664, N7543);
  and ginst2039 (N7672, N2653, N2664, N7573);
  and ginst2040 (N7673, N1161, N2664, N7549);
  and ginst2041 (N7674, N2728, N2739, N7555);
  and ginst2042 (N7675, N1223, N2739, N7531);
  and ginst2043 (N7676, N2728, N2739, N7561);
  and ginst2044 (N7677, N1223, N2739, N7537);
  and ginst2045 (N7678, N2728, N2739, N7567);
  and ginst2046 (N7679, N1223, N2739, N7543);
  and ginst2047 (N7680, N2728, N2739, N7573);
  and ginst2048 (N7681, N1223, N2739, N7549);
  and ginst2049 (N7682, N3075, N3086, N7573);
  and ginst2050 (N7683, N1731, N3086, N7549);
  and ginst2051 (N7684, N3041, N3052, N7573);
  and ginst2052 (N7685, N1697, N3052, N7549);
  and ginst2053 (N7686, N3041, N3052, N7567);
  and ginst2054 (N7687, N1697, N3052, N7543);
  and ginst2055 (N7688, N3041, N3052, N7561);
  and ginst2056 (N7689, N1697, N3052, N7537);
  and ginst2057 (N7690, N3041, N3052, N7555);
  and ginst2058 (N7691, N1697, N3052, N7531);
  and ginst2059 (N7692, N3075, N3086, N7567);
  and ginst2060 (N7693, N1731, N3086, N7543);
  and ginst2061 (N7694, N3075, N3086, N7561);
  and ginst2062 (N7695, N1731, N3086, N7537);
  and ginst2063 (N7696, N3075, N3086, N7555);
  and ginst2064 (N7697, N1731, N3086, N7531);
  or ginst2065 (N7698, N7624, N7625);
  not ginst2066 (N7699, N7573);
  not ginst2067 (N7700, N7567);
  not ginst2068 (N7701, N7561);
  not ginst2069 (N7702, N7555);
  and ginst2070 (N7703, N245, N1156, N7631);
  not ginst2071 (N7704, N7549);
  not ginst2072 (N7705, N7543);
  not ginst2073 (N7706, N7537);
  not ginst2074 (N7707, N7531);
  not ginst2075 (N7708, N7579);
  nand ginst2076 (N7709, N6739, N7579);
  not ginst2077 (N7710, N7582);
  nand ginst2078 (N7711, N6744, N7582);
  nand ginst2079 (N7712, N7586, N7657);
  nand ginst2080 (N7715, N7588, N7658);
  not ginst2081 (N7718, N7589);
  nand ginst2082 (N7719, N6772, N7589);
  not ginst2083 (N7720, N7592);
  nand ginst2084 (N7721, N6776, N7592);
  not ginst2085 (N7722, N7595);
  nand ginst2086 (N7723, N5733, N7595);
  nand ginst2087 (N7724, N7599, N7665);
  or ginst2088 (N7727, N2586, N3617, N7666, N7667);
  or ginst2089 (N7728, N2587, N3618, N7668, N7669);
  or ginst2090 (N7729, N2588, N3619, N7670, N7671);
  or ginst2091 (N7730, N2589, N3620, N7672, N7673);
  or ginst2092 (N7731, N2596, N3628, N7674, N7675);
  or ginst2093 (N7732, N2597, N3629, N7676, N7677);
  or ginst2094 (N7733, N2598, N3630, N7678, N7679);
  or ginst2095 (N7734, N2599, N3631, N7680, N7681);
  or ginst2096 (N7735, N2604, N3638, N7682, N7683);
  or ginst2097 (N7736, N2606, N3642, N7684, N7685);
  or ginst2098 (N7737, N2607, N3643, N7686, N7687);
  or ginst2099 (N7738, N2608, N3644, N7688, N7689);
  or ginst2100 (N7739, N2609, N3645, N7690, N7691);
  or ginst2101 (N7740, N2615, N3651, N7692, N7693);
  or ginst2102 (N7741, N2616, N3652, N7694, N7695);
  or ginst2103 (N7742, N2617, N3653, N7696, N7697);
  nand ginst2104 (N7743, N6271, N7708);
  nand ginst2105 (N7744, N6283, N7710);
  nand ginst2106 (N7749, N6341, N7718);
  nand ginst2107 (N7750, N6347, N7720);
  nand ginst2108 (N7751, N5214, N7722);
  and ginst2109 (N7754, N2647, N7727);
  and ginst2110 (N7755, N2647, N7728);
  and ginst2111 (N7756, N2647, N7729);
  and ginst2112 (N7757, N2647, N7730);
  and ginst2113 (N7758, N2722, N7731);
  and ginst2114 (N7759, N2722, N7732);
  and ginst2115 (N7760, N2722, N7733);
  and ginst2116 (N7761, N2722, N7734);
  nand ginst2117 (N7762, N7709, N7743);
  nand ginst2118 (N7765, N7711, N7744);
  not ginst2119 (N7768, N7712);
  nand ginst2120 (N7769, N6751, N7712);
  not ginst2121 (N7770, N7715);
  nand ginst2122 (N7771, N6760, N7715);
  nand ginst2123 (N7772, N7719, N7749);
  nand ginst2124 (N7775, N7721, N7750);
  nand ginst2125 (N7778, N7723, N7751);
  not ginst2126 (N7781, N7724);
  nand ginst2127 (N7782, N5735, N7724);
  nand ginst2128 (N7787, N6295, N7768);
  nand ginst2129 (N7788, N6313, N7770);
  nand ginst2130 (N7795, N5220, N7781);
  not ginst2131 (N7796, N7762);
  nand ginst2132 (N7797, N6740, N7762);
  not ginst2133 (N7798, N7765);
  nand ginst2134 (N7799, N6745, N7765);
  nand ginst2135 (N7800, N7769, N7787);
  nand ginst2136 (N7803, N7771, N7788);
  not ginst2137 (N7806, N7772);
  nand ginst2138 (N7807, N6773, N7772);
  not ginst2139 (N7808, N7775);
  nand ginst2140 (N7809, N6777, N7775);
  not ginst2141 (N7810, N7778);
  nand ginst2142 (N7811, N6782, N7778);
  nand ginst2143 (N7812, N7782, N7795);
  nand ginst2144 (N7815, N6274, N7796);
  nand ginst2145 (N7816, N6286, N7798);
  nand ginst2146 (N7821, N6344, N7806);
  nand ginst2147 (N7822, N6350, N7808);
  nand ginst2148 (N7823, N6353, N7810);
  nand ginst2149 (N7826, N7797, N7815);
  nand ginst2150 (N7829, N7799, N7816);
  not ginst2151 (N7832, N7800);
  nand ginst2152 (N7833, N6752, N7800);
  not ginst2153 (N7834, N7803);
  nand ginst2154 (N7835, N6761, N7803);
  nand ginst2155 (N7836, N7807, N7821);
  nand ginst2156 (N7839, N7809, N7822);
  nand ginst2157 (N7842, N7811, N7823);
  not ginst2158 (N7845, N7812);
  nand ginst2159 (N7846, N6790, N7812);
  nand ginst2160 (N7851, N6298, N7832);
  nand ginst2161 (N7852, N6316, N7834);
  nand ginst2162 (N7859, N6364, N7845);
  not ginst2163 (N7860, N7826);
  nand ginst2164 (N7861, N6741, N7826);
  not ginst2165 (N7862, N7829);
  nand ginst2166 (N7863, N6746, N7829);
  nand ginst2167 (N7864, N7833, N7851);
  nand ginst2168 (N7867, N7835, N7852);
  not ginst2169 (N7870, N7836);
  nand ginst2170 (N7871, N5730, N7836);
  not ginst2171 (N7872, N7839);
  nand ginst2172 (N7873, N5732, N7839);
  not ginst2173 (N7874, N7842);
  nand ginst2174 (N7875, N6783, N7842);
  nand ginst2175 (N7876, N7846, N7859);
  nand ginst2176 (N7879, N6277, N7860);
  nand ginst2177 (N7880, N6289, N7862);
  nand ginst2178 (N7885, N5199, N7870);
  nand ginst2179 (N7886, N5208, N7872);
  nand ginst2180 (N7887, N6356, N7874);
  nand ginst2181 (N7890, N7861, N7879);
  nand ginst2182 (N7893, N7863, N7880);
  not ginst2183 (N7896, N7864);
  nand ginst2184 (N7897, N6753, N7864);
  not ginst2185 (N7898, N7867);
  nand ginst2186 (N7899, N6762, N7867);
  nand ginst2187 (N7900, N7871, N7885);
  nand ginst2188 (N7903, N7873, N7886);
  nand ginst2189 (N7906, N7875, N7887);
  not ginst2190 (N7909, N7876);
  nand ginst2191 (N7910, N6791, N7876);
  nand ginst2192 (N7917, N6301, N7896);
  nand ginst2193 (N7918, N6319, N7898);
  nand ginst2194 (N7923, N6367, N7909);
  not ginst2195 (N7924, N7890);
  nand ginst2196 (N7925, N6680, N7890);
  not ginst2197 (N7926, N7893);
  nand ginst2198 (N7927, N6681, N7893);
  not ginst2199 (N7928, N7900);
  nand ginst2200 (N7929, N5690, N7900);
  not ginst2201 (N7930, N7903);
  nand ginst2202 (N7931, N5691, N7903);
  nand ginst2203 (N7932, N7897, N7917);
  nand ginst2204 (N7935, N7899, N7918);
  not ginst2205 (N7938, N7906);
  nand ginst2206 (N7939, N6784, N7906);
  nand ginst2207 (N7940, N7910, N7923);
  nand ginst2208 (N7943, N6280, N7924);
  nand ginst2209 (N7944, N6292, N7926);
  nand ginst2210 (N7945, N5202, N7928);
  nand ginst2211 (N7946, N5211, N7930);
  nand ginst2212 (N7951, N6359, N7938);
  nand ginst2213 (N7954, N7925, N7943);
  nand ginst2214 (N7957, N7927, N7944);
  nand ginst2215 (N7960, N7929, N7945);
  nand ginst2216 (N7963, N7931, N7946);
  not ginst2217 (N7966, N7932);
  nand ginst2218 (N7967, N6754, N7932);
  not ginst2219 (N7968, N7935);
  nand ginst2220 (N7969, N6755, N7935);
  nand ginst2221 (N7970, N7939, N7951);
  not ginst2222 (N7973, N7940);
  nand ginst2223 (N7974, N6785, N7940);
  nand ginst2224 (N7984, N6304, N7966);
  nand ginst2225 (N7985, N6322, N7968);
  nand ginst2226 (N7987, N6370, N7973);
  and ginst2227 (N7988, N1157, N6831, N7957);
  and ginst2228 (N7989, N1157, N6415, N7954);
  and ginst2229 (N7990, N566, N7041, N7957);
  and ginst2230 (N7991, N566, N7177, N7954);
  not ginst2231 (N7992, N7970);
  nand ginst2232 (N7993, N6448, N7970);
  and ginst2233 (N7994, N1219, N6857, N7963);
  and ginst2234 (N7995, N1219, N6441, N7960);
  and ginst2235 (N7996, N583, N7065, N7963);
  and ginst2236 (N7997, N583, N7182, N7960);
  nand ginst2237 (N7998, N7967, N7984);
  nand ginst2238 (N8001, N7969, N7985);
  nand ginst2239 (N8004, N7974, N7987);
  nand ginst2240 (N8009, N6051, N7992);
  or ginst2241 (N8013, N7988, N7989, N7990, N7991);
  or ginst2242 (N8017, N7994, N7995, N7996, N7997);
  not ginst2243 (N8020, N7998);
  nand ginst2244 (N8021, N6682, N7998);
  not ginst2245 (N8022, N8001);
  nand ginst2246 (N8023, N6683, N8001);
  nand ginst2247 (N8025, N7993, N8009);
  not ginst2248 (N8026, N8004);
  nand ginst2249 (N8027, N6449, N8004);
  nand ginst2250 (N8031, N6307, N8020);
  nand ginst2251 (N8032, N6310, N8022);
  not ginst2252 (N8033, N8013);
  nand ginst2253 (N8034, N6054, N8026);
  and ginst2254 (N8035, N583, N8025);
  not ginst2255 (N8036, N8017);
  nand ginst2256 (N8037, N8021, N8031);
  nand ginst2257 (N8038, N8023, N8032);
  nand ginst2258 (N8039, N8027, N8034);
  not ginst2259 (N8040, N8038);
  and ginst2260 (N8041, N566, N8037);
  not ginst2261 (N8042, N8039);
  and ginst2262 (N8043, N1157, N8040);
  and ginst2263 (N8044, N1219, N8042);
  or ginst2264 (N8045, N8041, N8043);
  or ginst2265 (N8048, N8035, N8044);
  nand ginst2266 (N8055, N8033, N8045);
  not ginst2267 (N8056, N8045);
  nand ginst2268 (N8057, N8036, N8048);
  not ginst2269 (N8058, N8048);
  nand ginst2270 (N8059, N8013, N8056);
  nand ginst2271 (N8060, N8017, N8058);
  nand ginst2272 (N8061, N8055, N8059);
  nand ginst2273 (N8064, N8057, N8060);
  and ginst2274 (N8071, N1777, N3130, N8064);
  and ginst2275 (N8072, N1761, N3108, N8061);
  not ginst2276 (N8073, N8061);
  not ginst2277 (N8074, N8064);
  or ginst2278 (N8075, N2625, N3659, N7526, N8071);
  or ginst2279 (N8076, N2627, N3661, N7636, N8072);
  and ginst2280 (N8077, N1727, N8073);
  and ginst2281 (N8078, N1727, N8074);
  or ginst2282 (N8079, N7530, N8077);
  or ginst2283 (N8082, N7479, N8078);
  and ginst2284 (N8089, N3063, N8079);
  and ginst2285 (N8090, N3063, N8082);
  and ginst2286 (N8091, N3063, N8079);
  and ginst2287 (N8092, N3063, N8082);
  or ginst2288 (N8093, N3071, N8089);
  or ginst2289 (N8096, N3072, N8090);
  or ginst2290 (N8099, N3073, N8091);
  or ginst2291 (N8102, N3074, N8092);
  and ginst2292 (N8113, N2779, N2790, N8102);
  and ginst2293 (N8114, N1327, N2790, N8099);
  and ginst2294 (N8115, N2801, N2812, N8102);
  and ginst2295 (N8116, N1351, N2812, N8099);
  and ginst2296 (N8117, N2681, N2692, N8096);
  and ginst2297 (N8118, N1185, N2692, N8093);
  and ginst2298 (N8119, N2756, N2767, N8096);
  and ginst2299 (N8120, N1247, N2767, N8093);
  or ginst2300 (N8121, N2703, N3662, N8117, N8118);
  or ginst2301 (N8122, N2778, N3663, N8119, N8120);
  or ginst2302 (N8123, N2614, N3650, N8113, N8114);
  or ginst2303 (N8124, N2622, N3658, N8115, N8116);
  and ginst2304 (N8125, N2675, N8121);
  and ginst2305 (N8126, N2750, N8122);
  not ginst2306 (N8127, N8125);
  not ginst2307 (N8128, N8126);
  buf ginst2308 (N816, N293);

endmodule

/*************** SatHard block ***************/
module SatHard (N137, N331, N54, N534, keyinput0, keyinput1, keyinput2, keyinput3, keyinput4, keyinput5, keyinput6, keyinput7, flip_signal);

  input N137, N331, N54, N534, keyinput0, keyinput1, keyinput2, keyinput3, keyinput4, keyinput5, keyinput6, keyinput7;
  output flip_signal;
  //SatHard key=01100110
  wire [3:0] sat_res_inputs;
  wire [7:0] keyinputs, keyvalue;
  assign sat_res_inputs[3:0] = {N137, N331, N54, N534};
  assign keyinputs[7:0] = {keyinput0, keyinput1, keyinput2, keyinput3, keyinput4, keyinput5, keyinput6, keyinput7};
  assign keyvalue[7:0] = 8'b01100110;

  wire g, g_bar;
  assign g = &(keyinputs[3:0] ^ sat_res_inputs ^ keyvalue[3:0]);
  assign g_bar = ~&(keyinputs[7:4] ^ sat_res_inputs ^ keyvalue[7:4]);
  assign flip_signal = g & g_bar;

endmodule
/*************** SatHard block ***************/
