/*************** Top Level ***************/
module b15_C_SFLL_HD_4_32_1_top (DATAO_REG_25__SCAN_IN, DATAO_REG_5__SCAN_IN, DATAO_REG_28__SCAN_IN, DATAO_REG_21__SCAN_IN, BE_N_REG_0__SCAN_IN, ADDRESS_REG_23__SCAN_IN, ADDRESS_REG_17__SCAN_IN, ADDRESS_REG_2__SCAN_IN, DATAO_REG_30__SCAN_IN, BE_N_REG_1__SCAN_IN, ADDRESS_REG_1__SCAN_IN, DATAO_REG_8__SCAN_IN, DATAO_REG_23__SCAN_IN, DATAO_REG_10__SCAN_IN, ADDRESS_REG_22__SCAN_IN, ADDRESS_REG_11__SCAN_IN, ADDRESS_REG_3__SCAN_IN, BE_N_REG_3__SCAN_IN, DATAO_REG_27__SCAN_IN, ADDRESS_REG_10__SCAN_IN, ADDRESS_REG_28__SCAN_IN, DATAO_REG_12__SCAN_IN, BE_N_REG_2__SCAN_IN, ADDRESS_REG_13__SCAN_IN, DATAO_REG_13__SCAN_IN, ADDRESS_REG_20__SCAN_IN, DATAO_REG_24__SCAN_IN, DATAO_REG_9__SCAN_IN, DATAO_REG_7__SCAN_IN, DATAO_REG_11__SCAN_IN, ADDRESS_REG_19__SCAN_IN, ADDRESS_REG_27__SCAN_IN, ADDRESS_REG_25__SCAN_IN, ADDRESS_REG_29__SCAN_IN, ADDRESS_REG_5__SCAN_IN, ADDRESS_REG_7__SCAN_IN, ADDRESS_REG_8__SCAN_IN, ADDRESS_REG_21__SCAN_IN, DATAO_REG_20__SCAN_IN, DATAO_REG_17__SCAN_IN, DATAO_REG_6__SCAN_IN, ADDRESS_REG_14__SCAN_IN, DATAO_REG_19__SCAN_IN, ADS_N_REG_SCAN_IN, DATAO_REG_15__SCAN_IN, DATAO_REG_26__SCAN_IN, DATAO_REG_3__SCAN_IN, DATAO_REG_1__SCAN_IN, ADDRESS_REG_26__SCAN_IN, ADDRESS_REG_18__SCAN_IN, M_IO_N_REG_SCAN_IN, DATAO_REG_31__SCAN_IN, ADDRESS_REG_16__SCAN_IN, ADDRESS_REG_9__SCAN_IN, ADDRESS_REG_12__SCAN_IN, DATAO_REG_29__SCAN_IN, DATAO_REG_0__SCAN_IN, ADDRESS_REG_4__SCAN_IN, D_C_N_REG_SCAN_IN, DATAO_REG_4__SCAN_IN, ADDRESS_REG_6__SCAN_IN, DATAO_REG_2__SCAN_IN, ADDRESS_REG_0__SCAN_IN, DATAO_REG_18__SCAN_IN, DATAO_REG_16__SCAN_IN, ADDRESS_REG_24__SCAN_IN, DATAO_REG_14__SCAN_IN, W_R_N_REG_SCAN_IN, ADDRESS_REG_15__SCAN_IN, DATAO_REG_22__SCAN_IN, DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, DATAI_27_, DATAI_26_, DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, DATAI_21_, DATAI_20_, DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, DATAI_15_, DATAI_14_, DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, DATAI_9_, DATAI_8_, DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, DATAI_2_, DATAI_1_, DATAI_0_, MEMORYFETCH_REG_SCAN_IN, NA_N, BS16_N, READY_N, HOLD, READREQUEST_REG_SCAN_IN, CODEFETCH_REG_SCAN_IN, REQUESTPENDING_REG_SCAN_IN, STATEBS16_REG_SCAN_IN, MORE_REG_SCAN_IN, FLUSH_REG_SCAN_IN, BYTEENABLE_REG_0__SCAN_IN, BYTEENABLE_REG_1__SCAN_IN, BYTEENABLE_REG_2__SCAN_IN, BYTEENABLE_REG_3__SCAN_IN, REIP_REG_31__SCAN_IN, REIP_REG_30__SCAN_IN, REIP_REG_29__SCAN_IN, REIP_REG_28__SCAN_IN, REIP_REG_27__SCAN_IN, REIP_REG_26__SCAN_IN, REIP_REG_25__SCAN_IN, REIP_REG_24__SCAN_IN, REIP_REG_23__SCAN_IN, REIP_REG_22__SCAN_IN, REIP_REG_21__SCAN_IN, REIP_REG_20__SCAN_IN, REIP_REG_19__SCAN_IN, REIP_REG_18__SCAN_IN, REIP_REG_17__SCAN_IN, REIP_REG_16__SCAN_IN, STATE_REG_2__SCAN_IN, STATE_REG_1__SCAN_IN, STATE_REG_0__SCAN_IN, DATAWIDTH_REG_0__SCAN_IN, DATAWIDTH_REG_1__SCAN_IN, DATAWIDTH_REG_2__SCAN_IN, DATAWIDTH_REG_3__SCAN_IN, DATAWIDTH_REG_4__SCAN_IN, DATAWIDTH_REG_5__SCAN_IN, DATAWIDTH_REG_6__SCAN_IN, DATAWIDTH_REG_7__SCAN_IN, DATAWIDTH_REG_8__SCAN_IN, DATAWIDTH_REG_9__SCAN_IN, DATAWIDTH_REG_10__SCAN_IN, DATAWIDTH_REG_11__SCAN_IN, DATAWIDTH_REG_12__SCAN_IN, DATAWIDTH_REG_13__SCAN_IN, DATAWIDTH_REG_14__SCAN_IN, DATAWIDTH_REG_15__SCAN_IN, DATAWIDTH_REG_16__SCAN_IN, DATAWIDTH_REG_17__SCAN_IN, DATAWIDTH_REG_18__SCAN_IN, DATAWIDTH_REG_19__SCAN_IN, DATAWIDTH_REG_20__SCAN_IN, DATAWIDTH_REG_21__SCAN_IN, DATAWIDTH_REG_22__SCAN_IN, DATAWIDTH_REG_23__SCAN_IN, DATAWIDTH_REG_24__SCAN_IN, DATAWIDTH_REG_25__SCAN_IN, DATAWIDTH_REG_26__SCAN_IN, DATAWIDTH_REG_27__SCAN_IN, DATAWIDTH_REG_28__SCAN_IN, DATAWIDTH_REG_29__SCAN_IN, DATAWIDTH_REG_30__SCAN_IN, DATAWIDTH_REG_31__SCAN_IN, STATE2_REG_3__SCAN_IN, STATE2_REG_2__SCAN_IN, STATE2_REG_1__SCAN_IN, STATE2_REG_0__SCAN_IN, INSTQUEUE_REG_15__7__SCAN_IN, INSTQUEUE_REG_15__6__SCAN_IN, INSTQUEUE_REG_15__5__SCAN_IN, INSTQUEUE_REG_15__4__SCAN_IN, INSTQUEUE_REG_15__3__SCAN_IN, INSTQUEUE_REG_15__2__SCAN_IN, INSTQUEUE_REG_15__1__SCAN_IN, INSTQUEUE_REG_15__0__SCAN_IN, INSTQUEUE_REG_14__7__SCAN_IN, INSTQUEUE_REG_14__6__SCAN_IN, INSTQUEUE_REG_14__5__SCAN_IN, INSTQUEUE_REG_14__4__SCAN_IN, INSTQUEUE_REG_14__3__SCAN_IN, INSTQUEUE_REG_14__2__SCAN_IN, INSTQUEUE_REG_14__1__SCAN_IN, INSTQUEUE_REG_14__0__SCAN_IN, INSTQUEUE_REG_13__7__SCAN_IN, INSTQUEUE_REG_13__6__SCAN_IN, INSTQUEUE_REG_13__5__SCAN_IN, INSTQUEUE_REG_13__4__SCAN_IN, INSTQUEUE_REG_13__3__SCAN_IN, INSTQUEUE_REG_13__2__SCAN_IN, INSTQUEUE_REG_13__1__SCAN_IN, INSTQUEUE_REG_13__0__SCAN_IN, INSTQUEUE_REG_12__7__SCAN_IN, INSTQUEUE_REG_12__6__SCAN_IN, INSTQUEUE_REG_12__5__SCAN_IN, INSTQUEUE_REG_12__4__SCAN_IN, INSTQUEUE_REG_12__3__SCAN_IN, INSTQUEUE_REG_12__2__SCAN_IN, INSTQUEUE_REG_12__1__SCAN_IN, INSTQUEUE_REG_12__0__SCAN_IN, INSTQUEUE_REG_11__7__SCAN_IN, INSTQUEUE_REG_11__6__SCAN_IN, INSTQUEUE_REG_11__5__SCAN_IN, INSTQUEUE_REG_11__4__SCAN_IN, INSTQUEUE_REG_11__3__SCAN_IN, INSTQUEUE_REG_11__2__SCAN_IN, INSTQUEUE_REG_11__1__SCAN_IN, INSTQUEUE_REG_11__0__SCAN_IN, INSTQUEUE_REG_10__7__SCAN_IN, INSTQUEUE_REG_10__6__SCAN_IN, INSTQUEUE_REG_10__5__SCAN_IN, INSTQUEUE_REG_10__4__SCAN_IN, INSTQUEUE_REG_10__3__SCAN_IN, INSTQUEUE_REG_10__2__SCAN_IN, INSTQUEUE_REG_10__1__SCAN_IN, INSTQUEUE_REG_10__0__SCAN_IN, INSTQUEUE_REG_9__7__SCAN_IN, INSTQUEUE_REG_9__6__SCAN_IN, INSTQUEUE_REG_9__5__SCAN_IN, INSTQUEUE_REG_9__4__SCAN_IN, INSTQUEUE_REG_9__3__SCAN_IN, INSTQUEUE_REG_9__2__SCAN_IN, INSTQUEUE_REG_9__1__SCAN_IN, INSTQUEUE_REG_9__0__SCAN_IN, INSTQUEUE_REG_8__7__SCAN_IN, INSTQUEUE_REG_8__6__SCAN_IN, INSTQUEUE_REG_8__5__SCAN_IN, INSTQUEUE_REG_8__4__SCAN_IN, INSTQUEUE_REG_8__3__SCAN_IN, INSTQUEUE_REG_8__2__SCAN_IN, INSTQUEUE_REG_8__1__SCAN_IN, INSTQUEUE_REG_8__0__SCAN_IN, INSTQUEUE_REG_7__7__SCAN_IN, INSTQUEUE_REG_7__6__SCAN_IN, INSTQUEUE_REG_7__5__SCAN_IN, INSTQUEUE_REG_7__4__SCAN_IN, INSTQUEUE_REG_7__3__SCAN_IN, INSTQUEUE_REG_7__2__SCAN_IN, INSTQUEUE_REG_7__1__SCAN_IN, INSTQUEUE_REG_7__0__SCAN_IN, INSTQUEUE_REG_6__7__SCAN_IN, INSTQUEUE_REG_6__6__SCAN_IN, INSTQUEUE_REG_6__5__SCAN_IN, INSTQUEUE_REG_6__4__SCAN_IN, INSTQUEUE_REG_6__3__SCAN_IN, INSTQUEUE_REG_6__2__SCAN_IN, INSTQUEUE_REG_6__1__SCAN_IN, INSTQUEUE_REG_6__0__SCAN_IN, INSTQUEUE_REG_5__7__SCAN_IN, INSTQUEUE_REG_5__6__SCAN_IN, INSTQUEUE_REG_5__5__SCAN_IN, INSTQUEUE_REG_5__4__SCAN_IN, INSTQUEUE_REG_5__3__SCAN_IN, INSTQUEUE_REG_5__2__SCAN_IN, INSTQUEUE_REG_5__1__SCAN_IN, INSTQUEUE_REG_5__0__SCAN_IN, INSTQUEUE_REG_4__7__SCAN_IN, INSTQUEUE_REG_4__6__SCAN_IN, INSTQUEUE_REG_4__5__SCAN_IN, INSTQUEUE_REG_4__4__SCAN_IN, INSTQUEUE_REG_4__3__SCAN_IN, INSTQUEUE_REG_4__2__SCAN_IN, INSTQUEUE_REG_4__1__SCAN_IN, INSTQUEUE_REG_4__0__SCAN_IN, INSTQUEUE_REG_3__7__SCAN_IN, INSTQUEUE_REG_3__6__SCAN_IN, INSTQUEUE_REG_3__5__SCAN_IN, INSTQUEUE_REG_3__4__SCAN_IN, INSTQUEUE_REG_3__3__SCAN_IN, INSTQUEUE_REG_3__2__SCAN_IN, INSTQUEUE_REG_3__1__SCAN_IN, INSTQUEUE_REG_3__0__SCAN_IN, INSTQUEUE_REG_2__7__SCAN_IN, INSTQUEUE_REG_2__6__SCAN_IN, INSTQUEUE_REG_2__5__SCAN_IN, INSTQUEUE_REG_2__4__SCAN_IN, INSTQUEUE_REG_2__3__SCAN_IN, INSTQUEUE_REG_2__2__SCAN_IN, INSTQUEUE_REG_2__1__SCAN_IN, INSTQUEUE_REG_2__0__SCAN_IN, INSTQUEUE_REG_1__7__SCAN_IN, INSTQUEUE_REG_1__6__SCAN_IN, INSTQUEUE_REG_1__5__SCAN_IN, INSTQUEUE_REG_1__4__SCAN_IN, INSTQUEUE_REG_1__3__SCAN_IN, INSTQUEUE_REG_1__2__SCAN_IN, INSTQUEUE_REG_1__1__SCAN_IN, INSTQUEUE_REG_1__0__SCAN_IN, INSTQUEUE_REG_0__7__SCAN_IN, INSTQUEUE_REG_0__6__SCAN_IN, INSTQUEUE_REG_0__5__SCAN_IN, INSTQUEUE_REG_0__4__SCAN_IN, INSTQUEUE_REG_0__3__SCAN_IN, INSTQUEUE_REG_0__2__SCAN_IN, INSTQUEUE_REG_0__1__SCAN_IN, INSTQUEUE_REG_0__0__SCAN_IN, INSTQUEUERD_ADDR_REG_4__SCAN_IN, INSTQUEUERD_ADDR_REG_3__SCAN_IN, INSTQUEUERD_ADDR_REG_2__SCAN_IN, INSTQUEUERD_ADDR_REG_1__SCAN_IN, INSTQUEUERD_ADDR_REG_0__SCAN_IN, INSTQUEUEWR_ADDR_REG_4__SCAN_IN, INSTQUEUEWR_ADDR_REG_3__SCAN_IN, INSTQUEUEWR_ADDR_REG_2__SCAN_IN, INSTQUEUEWR_ADDR_REG_1__SCAN_IN, INSTQUEUEWR_ADDR_REG_0__SCAN_IN, INSTADDRPOINTER_REG_0__SCAN_IN, INSTADDRPOINTER_REG_1__SCAN_IN, INSTADDRPOINTER_REG_2__SCAN_IN, INSTADDRPOINTER_REG_3__SCAN_IN, INSTADDRPOINTER_REG_4__SCAN_IN, INSTADDRPOINTER_REG_5__SCAN_IN, INSTADDRPOINTER_REG_6__SCAN_IN, INSTADDRPOINTER_REG_7__SCAN_IN, INSTADDRPOINTER_REG_8__SCAN_IN, INSTADDRPOINTER_REG_9__SCAN_IN, INSTADDRPOINTER_REG_10__SCAN_IN, INSTADDRPOINTER_REG_11__SCAN_IN, INSTADDRPOINTER_REG_12__SCAN_IN, INSTADDRPOINTER_REG_13__SCAN_IN, INSTADDRPOINTER_REG_14__SCAN_IN, INSTADDRPOINTER_REG_15__SCAN_IN, INSTADDRPOINTER_REG_16__SCAN_IN, INSTADDRPOINTER_REG_17__SCAN_IN, INSTADDRPOINTER_REG_18__SCAN_IN, INSTADDRPOINTER_REG_19__SCAN_IN, INSTADDRPOINTER_REG_20__SCAN_IN, INSTADDRPOINTER_REG_21__SCAN_IN, INSTADDRPOINTER_REG_22__SCAN_IN, INSTADDRPOINTER_REG_23__SCAN_IN, INSTADDRPOINTER_REG_24__SCAN_IN, INSTADDRPOINTER_REG_25__SCAN_IN, INSTADDRPOINTER_REG_26__SCAN_IN, INSTADDRPOINTER_REG_27__SCAN_IN, INSTADDRPOINTER_REG_28__SCAN_IN, INSTADDRPOINTER_REG_29__SCAN_IN, INSTADDRPOINTER_REG_30__SCAN_IN, INSTADDRPOINTER_REG_31__SCAN_IN, PHYADDRPOINTER_REG_0__SCAN_IN, PHYADDRPOINTER_REG_1__SCAN_IN, PHYADDRPOINTER_REG_2__SCAN_IN, PHYADDRPOINTER_REG_3__SCAN_IN, PHYADDRPOINTER_REG_4__SCAN_IN, PHYADDRPOINTER_REG_5__SCAN_IN, PHYADDRPOINTER_REG_6__SCAN_IN, PHYADDRPOINTER_REG_7__SCAN_IN, PHYADDRPOINTER_REG_8__SCAN_IN, PHYADDRPOINTER_REG_9__SCAN_IN, PHYADDRPOINTER_REG_10__SCAN_IN, PHYADDRPOINTER_REG_11__SCAN_IN, PHYADDRPOINTER_REG_12__SCAN_IN, PHYADDRPOINTER_REG_13__SCAN_IN, PHYADDRPOINTER_REG_14__SCAN_IN, PHYADDRPOINTER_REG_15__SCAN_IN, PHYADDRPOINTER_REG_16__SCAN_IN, PHYADDRPOINTER_REG_17__SCAN_IN, PHYADDRPOINTER_REG_18__SCAN_IN, PHYADDRPOINTER_REG_19__SCAN_IN, PHYADDRPOINTER_REG_20__SCAN_IN, PHYADDRPOINTER_REG_21__SCAN_IN, PHYADDRPOINTER_REG_22__SCAN_IN, PHYADDRPOINTER_REG_23__SCAN_IN, PHYADDRPOINTER_REG_24__SCAN_IN, PHYADDRPOINTER_REG_25__SCAN_IN, PHYADDRPOINTER_REG_26__SCAN_IN, PHYADDRPOINTER_REG_27__SCAN_IN, PHYADDRPOINTER_REG_28__SCAN_IN, PHYADDRPOINTER_REG_29__SCAN_IN, PHYADDRPOINTER_REG_30__SCAN_IN, PHYADDRPOINTER_REG_31__SCAN_IN, LWORD_REG_15__SCAN_IN, LWORD_REG_14__SCAN_IN, LWORD_REG_13__SCAN_IN, LWORD_REG_12__SCAN_IN, LWORD_REG_11__SCAN_IN, LWORD_REG_10__SCAN_IN, LWORD_REG_9__SCAN_IN, LWORD_REG_8__SCAN_IN, LWORD_REG_7__SCAN_IN, LWORD_REG_6__SCAN_IN, LWORD_REG_5__SCAN_IN, LWORD_REG_4__SCAN_IN, LWORD_REG_3__SCAN_IN, LWORD_REG_2__SCAN_IN, LWORD_REG_1__SCAN_IN, LWORD_REG_0__SCAN_IN, UWORD_REG_14__SCAN_IN, UWORD_REG_13__SCAN_IN, UWORD_REG_12__SCAN_IN, UWORD_REG_11__SCAN_IN, UWORD_REG_10__SCAN_IN, UWORD_REG_9__SCAN_IN, UWORD_REG_8__SCAN_IN, UWORD_REG_7__SCAN_IN, UWORD_REG_6__SCAN_IN, UWORD_REG_5__SCAN_IN, UWORD_REG_4__SCAN_IN, UWORD_REG_3__SCAN_IN, UWORD_REG_2__SCAN_IN, UWORD_REG_1__SCAN_IN, UWORD_REG_0__SCAN_IN, EAX_REG_0__SCAN_IN, EAX_REG_1__SCAN_IN, EAX_REG_2__SCAN_IN, EAX_REG_3__SCAN_IN, EAX_REG_4__SCAN_IN, EAX_REG_5__SCAN_IN, EAX_REG_6__SCAN_IN, EAX_REG_7__SCAN_IN, EAX_REG_8__SCAN_IN, EAX_REG_9__SCAN_IN, EAX_REG_10__SCAN_IN, EAX_REG_11__SCAN_IN, EAX_REG_12__SCAN_IN, EAX_REG_13__SCAN_IN, EAX_REG_14__SCAN_IN, EAX_REG_15__SCAN_IN, EAX_REG_16__SCAN_IN, EAX_REG_17__SCAN_IN, EAX_REG_18__SCAN_IN, EAX_REG_19__SCAN_IN, EAX_REG_20__SCAN_IN, EAX_REG_21__SCAN_IN, EAX_REG_22__SCAN_IN, EAX_REG_23__SCAN_IN, EAX_REG_24__SCAN_IN, EAX_REG_25__SCAN_IN, EAX_REG_26__SCAN_IN, EAX_REG_27__SCAN_IN, EAX_REG_28__SCAN_IN, EAX_REG_29__SCAN_IN, EAX_REG_30__SCAN_IN, EAX_REG_31__SCAN_IN, EBX_REG_0__SCAN_IN, EBX_REG_1__SCAN_IN, EBX_REG_2__SCAN_IN, EBX_REG_3__SCAN_IN, EBX_REG_4__SCAN_IN, EBX_REG_5__SCAN_IN, EBX_REG_6__SCAN_IN, EBX_REG_7__SCAN_IN, EBX_REG_8__SCAN_IN, EBX_REG_9__SCAN_IN, EBX_REG_10__SCAN_IN, EBX_REG_11__SCAN_IN, EBX_REG_12__SCAN_IN, EBX_REG_13__SCAN_IN, EBX_REG_14__SCAN_IN, EBX_REG_15__SCAN_IN, EBX_REG_16__SCAN_IN, EBX_REG_17__SCAN_IN, EBX_REG_18__SCAN_IN, EBX_REG_19__SCAN_IN, EBX_REG_20__SCAN_IN, EBX_REG_21__SCAN_IN, EBX_REG_22__SCAN_IN, EBX_REG_23__SCAN_IN, EBX_REG_24__SCAN_IN, EBX_REG_25__SCAN_IN, EBX_REG_26__SCAN_IN, EBX_REG_27__SCAN_IN, EBX_REG_28__SCAN_IN, EBX_REG_29__SCAN_IN, EBX_REG_30__SCAN_IN, EBX_REG_31__SCAN_IN, REIP_REG_0__SCAN_IN, REIP_REG_1__SCAN_IN, REIP_REG_2__SCAN_IN, REIP_REG_3__SCAN_IN, REIP_REG_4__SCAN_IN, REIP_REG_5__SCAN_IN, REIP_REG_6__SCAN_IN, REIP_REG_7__SCAN_IN, REIP_REG_8__SCAN_IN, REIP_REG_9__SCAN_IN, REIP_REG_10__SCAN_IN, REIP_REG_11__SCAN_IN, REIP_REG_12__SCAN_IN, REIP_REG_13__SCAN_IN, REIP_REG_14__SCAN_IN, REIP_REG_15__SCAN_IN, keyinput0, keyinput1, keyinput2, keyinput3, keyinput4, keyinput5, keyinput6, keyinput7, keyinput8, keyinput9, keyinput10, keyinput11, keyinput12, keyinput13, keyinput14, keyinput15, keyinput16, keyinput17, keyinput18, keyinput19, keyinput20, keyinput21, keyinput22, keyinput23, keyinput24, keyinput25, keyinput26, keyinput27, keyinput28, keyinput29, keyinput30, keyinput31, DATAO_REG_2__SCAN_IN_BUFF, ADDRESS_REG_17__SCAN_IN_BUFF, DATAO_REG_22__SCAN_IN_BUFF, U3460, U3176, U2834, U3097, U2809, U3464, U3119, U2938, U3124, U2992, U2920, U2884, U3122, U3179, U2853, U3107, U3055, U3011, U2891, U2830, ADDRESS_REG_2__SCAN_IN_BUFF, U2797, U2869, U3043, U2958, U3105, U3013, U3077, U3059, BE_N_REG_0__SCAN_IN_BUFF, ADDRESS_REG_9__SCAN_IN_BUFF, ADDRESS_REG_11__SCAN_IN_BUFF, U3199, U3141, ADDRESS_REG_22__SCAN_IN_BUFF, U2789, U3149, U2917, U3169, U2981, U2941, U2892, U3093, ADDRESS_REG_0__SCAN_IN_BUFF, U3003, U2906, U2875, ADDRESS_REG_6__SCAN_IN_BUFF, U2854, U3132, U3032, DATAO_REG_24__SCAN_IN_BUFF, U2872, ADDRESS_REG_3__SCAN_IN_BUFF, U3136, U3071, U2896, U3451, U3168, U3079, U2795, U2829, U2840, U2868, U3082, U2928, U2915, U3148, U2990, U3160, ADDRESS_REG_21__SCAN_IN_BUFF, U3024, U2864, U2803, U2844, U2889, U2852, U3147, U2914, U3034, U2876, U3062, U2972, U3050, U2828, U2951, W_R_N_REG_SCAN_IN_BUFF, U3014, DATAO_REG_1__SCAN_IN_BUFF, U3064, U2819, U2961, U3015, U3085, ADDRESS_REG_5__SCAN_IN_BUFF, U3208, U3027, U2993, U2987, U3201, DATAO_REG_9__SCAN_IN_BUFF, U2960, U3049, U2825, U2979, U3028, DATAO_REG_15__SCAN_IN_BUFF, U2957, U2971, U2850, U3095, U2977, U3041, U2837, U3452, U3052, ADDRESS_REG_8__SCAN_IN_BUFF, U2926, DATAO_REG_26__SCAN_IN_BUFF, U3157, U2973, DATAO_REG_29__SCAN_IN_BUFF, U3170, U3152, U3159, U3196, U3089, U2897, U3469, U2921, U2870, U3069, U3063, U3135, U3166, U3210, U3153, U2818, U2905, U2933, U2796, U3207, U2898, U3209, U3078, U2946, U2907, BE_N_REG_3__SCAN_IN_BUFF, U2943, U2866, U2881, U2976, U2899, U3175, U3180, DATAO_REG_14__SCAN_IN_BUFF, U3113, M_IO_N_REG_SCAN_IN_BUFF, U2843, U2877, U2919, U3100, U2916, U2934, DATAO_REG_12__SCAN_IN_BUFF, U3146, U2924, U3161, U3005, U2893, U2945, U3470, U3150, U3109, U3213, U2955, U3448, U3194, U2832, U2978, U3183, U2947, DATAO_REG_3__SCAN_IN_BUFF, ADDRESS_REG_15__SCAN_IN_BUFF, U3007, U3162, U3203, U3106, U2942, ADDRESS_REG_18__SCAN_IN_BUFF, U3035, U2975, U2820, U2969, U2963, U2909, U3140, U2925, U2983, U2967, U2805, U3021, U3054, U3092, U3173, U2790, U2871, U2922, U2988, U3156, ADDRESS_REG_23__SCAN_IN_BUFF, U2932, U2822, U2878, U3155, U3010, U2935, U2794, U3033, U3030, U2835, U3186, U2824, U2956, U3163, U2831, U3026, U3083, U2814, U2953, U2890, U2882, U2791, U3000, U2998, ADDRESS_REG_26__SCAN_IN_BUFF, ADDRESS_REG_27__SCAN_IN_BUFF, U3125, U2817, U3101, U2900, U2793, DATAO_REG_25__SCAN_IN_BUFF, U2995, U2985, U3121, U3009, U3099, U2952, DATAO_REG_13__SCAN_IN_BUFF, U3133, U2806, U2962, U2948, U2888, U3456, U3462, U3115, U2801, U3158, U2865, U3185, U3110, U3145, U2940, U3167, ADDRESS_REG_29__SCAN_IN_BUFF, U2863, U3174, U3198, U2813, U3057, U3459, U3068, U2827, U3154, U2901, DATAO_REG_21__SCAN_IN_BUFF, U2903, U2855, U3098, U3025, U3205, U2838, U3211, U3067, U2841, U2959, U3463, U2800, DATAO_REG_18__SCAN_IN_BUFF, U3118, DATAO_REG_23__SCAN_IN_BUFF, U2859, U3130, U2860, U3036, U3045, U3066, U3017, U2826, U3023, U2821, U2989, ADDRESS_REG_12__SCAN_IN_BUFF, U3206, U3190, U2918, BE_N_REG_2__SCAN_IN_BUFF, U3102, DATAO_REG_28__SCAN_IN_BUFF, U3472, U3193, U3151, U2858, U2931, U2912, U3129, U3137, U2804, U2846, U3461, U3037, U3202, U3084, U3002, U3143, U2815, U2845, DATAO_REG_5__SCAN_IN_BUFF, U2902, U2930, DATAO_REG_31__SCAN_IN_BUFF, ADDRESS_REG_4__SCAN_IN_BUFF, ADDRESS_REG_25__SCAN_IN_BUFF, DATAO_REG_16__SCAN_IN_BUFF, U3172, U3038, U3018, U2910, U2883, DATAO_REG_30__SCAN_IN_BUFF, U2939, U3103, U3075, U2894, U3001, U3114, U3060, U3039, DATAO_REG_7__SCAN_IN_BUFF, DATAO_REG_19__SCAN_IN_BUFF, U2799, U3047, U2879, DATAO_REG_17__SCAN_IN_BUFF, U2857, U2911, U2880, U2937, U2812, U3008, U2839, U3111, U2904, U3445, DATAO_REG_8__SCAN_IN_BUFF, U3029, U2974, U2810, U2833, U3447, U2982, DATAO_REG_20__SCAN_IN_BUFF, ADS_N_REG_SCAN_IN_BUFF, U3204, U3184, U3200, U2851, U2798, U3019, U2885, U3104, U3065, U3164, U3070, U3453, U3061, U3087, U3108, ADDRESS_REG_10__SCAN_IN_BUFF, U3127, U2867, U3138, DATAO_REG_0__SCAN_IN_BUFF, U2856, U3046, U3139, U3051, U3465, U2811, U3073, U3474, U3116, U3086, U3016, U3126, U3446, U2923, U2816, U2970, U3004, U3006, U3081, U2788, U2842, U2874, U2802, U2886, U2964, ADDRESS_REG_28__SCAN_IN_BUFF, U3020, U2913, U2895, DATAO_REG_4__SCAN_IN_BUFF, U2836, U2823, U2849, U2862, U3088, U3044, U2848, U3177, U2873, U2966, U2861, U3187, U3117, U2984, U3191, U3074, U3212, U2887, U3076, U2929, U3182, U2927, U3195, U3178, U2986, ADDRESS_REG_7__SCAN_IN_BUFF, ADDRESS_REG_13__SCAN_IN_BUFF, U3189, U2950, U3090, U3053, U2980, U3171, U3080, U2954, U2944, U3165, U3123, U3022, U3120, DATAO_REG_6__SCAN_IN_BUFF, U3072, DATAO_REG_27__SCAN_IN_BUFF, ADDRESS_REG_20__SCAN_IN_BUFF, U2968, U3144, U3134, U2847, U2994, U2936, DATAO_REG_11__SCAN_IN_BUFF, U3192, U2991, U2908, U2965, U3131, ADDRESS_REG_24__SCAN_IN_BUFF, U3181, U3040, U3197, DATAO_REG_10__SCAN_IN_BUFF, U3091, ADDRESS_REG_1__SCAN_IN_BUFF, U3112, U3042, U3188, D_C_N_REG_SCAN_IN_BUFF, U2808, ADDRESS_REG_14__SCAN_IN_BUFF, U3094, U3142, U2792, U2996, U3473, U3012, U3468, U2999, ADDRESS_REG_19__SCAN_IN_BUFF, U3471, U3058, BE_N_REG_1__SCAN_IN_BUFF, U3031, U2807, U2949, U2997, U3455, U3128, U3048, U3096, ADDRESS_REG_16__SCAN_IN_BUFF, U3056);

  input DATAO_REG_25__SCAN_IN, DATAO_REG_5__SCAN_IN, DATAO_REG_28__SCAN_IN, DATAO_REG_21__SCAN_IN, BE_N_REG_0__SCAN_IN, ADDRESS_REG_23__SCAN_IN, ADDRESS_REG_17__SCAN_IN, ADDRESS_REG_2__SCAN_IN, DATAO_REG_30__SCAN_IN, BE_N_REG_1__SCAN_IN, ADDRESS_REG_1__SCAN_IN, DATAO_REG_8__SCAN_IN, DATAO_REG_23__SCAN_IN, DATAO_REG_10__SCAN_IN, ADDRESS_REG_22__SCAN_IN, ADDRESS_REG_11__SCAN_IN, ADDRESS_REG_3__SCAN_IN, BE_N_REG_3__SCAN_IN, DATAO_REG_27__SCAN_IN, ADDRESS_REG_10__SCAN_IN, ADDRESS_REG_28__SCAN_IN, DATAO_REG_12__SCAN_IN, BE_N_REG_2__SCAN_IN, ADDRESS_REG_13__SCAN_IN, DATAO_REG_13__SCAN_IN, ADDRESS_REG_20__SCAN_IN, DATAO_REG_24__SCAN_IN, DATAO_REG_9__SCAN_IN, DATAO_REG_7__SCAN_IN, DATAO_REG_11__SCAN_IN, ADDRESS_REG_19__SCAN_IN, ADDRESS_REG_27__SCAN_IN, ADDRESS_REG_25__SCAN_IN, ADDRESS_REG_29__SCAN_IN, ADDRESS_REG_5__SCAN_IN, ADDRESS_REG_7__SCAN_IN, ADDRESS_REG_8__SCAN_IN, ADDRESS_REG_21__SCAN_IN, DATAO_REG_20__SCAN_IN, DATAO_REG_17__SCAN_IN, DATAO_REG_6__SCAN_IN, ADDRESS_REG_14__SCAN_IN, DATAO_REG_19__SCAN_IN, ADS_N_REG_SCAN_IN, DATAO_REG_15__SCAN_IN, DATAO_REG_26__SCAN_IN, DATAO_REG_3__SCAN_IN, DATAO_REG_1__SCAN_IN, ADDRESS_REG_26__SCAN_IN, ADDRESS_REG_18__SCAN_IN, M_IO_N_REG_SCAN_IN, DATAO_REG_31__SCAN_IN, ADDRESS_REG_16__SCAN_IN, ADDRESS_REG_9__SCAN_IN, ADDRESS_REG_12__SCAN_IN, DATAO_REG_29__SCAN_IN, DATAO_REG_0__SCAN_IN, ADDRESS_REG_4__SCAN_IN, D_C_N_REG_SCAN_IN, DATAO_REG_4__SCAN_IN, ADDRESS_REG_6__SCAN_IN, DATAO_REG_2__SCAN_IN, ADDRESS_REG_0__SCAN_IN, DATAO_REG_18__SCAN_IN, DATAO_REG_16__SCAN_IN, ADDRESS_REG_24__SCAN_IN, DATAO_REG_14__SCAN_IN, W_R_N_REG_SCAN_IN, ADDRESS_REG_15__SCAN_IN, DATAO_REG_22__SCAN_IN, DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, DATAI_27_, DATAI_26_, DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, DATAI_21_, DATAI_20_, DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, DATAI_15_, DATAI_14_, DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, DATAI_9_, DATAI_8_, DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, DATAI_2_, DATAI_1_, DATAI_0_, MEMORYFETCH_REG_SCAN_IN, NA_N, BS16_N, READY_N, HOLD, READREQUEST_REG_SCAN_IN, CODEFETCH_REG_SCAN_IN, REQUESTPENDING_REG_SCAN_IN, STATEBS16_REG_SCAN_IN, MORE_REG_SCAN_IN, FLUSH_REG_SCAN_IN, BYTEENABLE_REG_0__SCAN_IN, BYTEENABLE_REG_1__SCAN_IN, BYTEENABLE_REG_2__SCAN_IN, BYTEENABLE_REG_3__SCAN_IN, REIP_REG_31__SCAN_IN, REIP_REG_30__SCAN_IN, REIP_REG_29__SCAN_IN, REIP_REG_28__SCAN_IN, REIP_REG_27__SCAN_IN, REIP_REG_26__SCAN_IN, REIP_REG_25__SCAN_IN, REIP_REG_24__SCAN_IN, REIP_REG_23__SCAN_IN, REIP_REG_22__SCAN_IN, REIP_REG_21__SCAN_IN, REIP_REG_20__SCAN_IN, REIP_REG_19__SCAN_IN, REIP_REG_18__SCAN_IN, REIP_REG_17__SCAN_IN, REIP_REG_16__SCAN_IN, STATE_REG_2__SCAN_IN, STATE_REG_1__SCAN_IN, STATE_REG_0__SCAN_IN, DATAWIDTH_REG_0__SCAN_IN, DATAWIDTH_REG_1__SCAN_IN, DATAWIDTH_REG_2__SCAN_IN, DATAWIDTH_REG_3__SCAN_IN, DATAWIDTH_REG_4__SCAN_IN, DATAWIDTH_REG_5__SCAN_IN, DATAWIDTH_REG_6__SCAN_IN, DATAWIDTH_REG_7__SCAN_IN, DATAWIDTH_REG_8__SCAN_IN, DATAWIDTH_REG_9__SCAN_IN, DATAWIDTH_REG_10__SCAN_IN, DATAWIDTH_REG_11__SCAN_IN, DATAWIDTH_REG_12__SCAN_IN, DATAWIDTH_REG_13__SCAN_IN, DATAWIDTH_REG_14__SCAN_IN, DATAWIDTH_REG_15__SCAN_IN, DATAWIDTH_REG_16__SCAN_IN, DATAWIDTH_REG_17__SCAN_IN, DATAWIDTH_REG_18__SCAN_IN, DATAWIDTH_REG_19__SCAN_IN, DATAWIDTH_REG_20__SCAN_IN, DATAWIDTH_REG_21__SCAN_IN, DATAWIDTH_REG_22__SCAN_IN, DATAWIDTH_REG_23__SCAN_IN, DATAWIDTH_REG_24__SCAN_IN, DATAWIDTH_REG_25__SCAN_IN, DATAWIDTH_REG_26__SCAN_IN, DATAWIDTH_REG_27__SCAN_IN, DATAWIDTH_REG_28__SCAN_IN, DATAWIDTH_REG_29__SCAN_IN, DATAWIDTH_REG_30__SCAN_IN, DATAWIDTH_REG_31__SCAN_IN, STATE2_REG_3__SCAN_IN, STATE2_REG_2__SCAN_IN, STATE2_REG_1__SCAN_IN, STATE2_REG_0__SCAN_IN, INSTQUEUE_REG_15__7__SCAN_IN, INSTQUEUE_REG_15__6__SCAN_IN, INSTQUEUE_REG_15__5__SCAN_IN, INSTQUEUE_REG_15__4__SCAN_IN, INSTQUEUE_REG_15__3__SCAN_IN, INSTQUEUE_REG_15__2__SCAN_IN, INSTQUEUE_REG_15__1__SCAN_IN, INSTQUEUE_REG_15__0__SCAN_IN, INSTQUEUE_REG_14__7__SCAN_IN, INSTQUEUE_REG_14__6__SCAN_IN, INSTQUEUE_REG_14__5__SCAN_IN, INSTQUEUE_REG_14__4__SCAN_IN, INSTQUEUE_REG_14__3__SCAN_IN, INSTQUEUE_REG_14__2__SCAN_IN, INSTQUEUE_REG_14__1__SCAN_IN, INSTQUEUE_REG_14__0__SCAN_IN, INSTQUEUE_REG_13__7__SCAN_IN, INSTQUEUE_REG_13__6__SCAN_IN, INSTQUEUE_REG_13__5__SCAN_IN, INSTQUEUE_REG_13__4__SCAN_IN, INSTQUEUE_REG_13__3__SCAN_IN, INSTQUEUE_REG_13__2__SCAN_IN, INSTQUEUE_REG_13__1__SCAN_IN, INSTQUEUE_REG_13__0__SCAN_IN, INSTQUEUE_REG_12__7__SCAN_IN, INSTQUEUE_REG_12__6__SCAN_IN, INSTQUEUE_REG_12__5__SCAN_IN, INSTQUEUE_REG_12__4__SCAN_IN, INSTQUEUE_REG_12__3__SCAN_IN, INSTQUEUE_REG_12__2__SCAN_IN, INSTQUEUE_REG_12__1__SCAN_IN, INSTQUEUE_REG_12__0__SCAN_IN, INSTQUEUE_REG_11__7__SCAN_IN, INSTQUEUE_REG_11__6__SCAN_IN, INSTQUEUE_REG_11__5__SCAN_IN, INSTQUEUE_REG_11__4__SCAN_IN, INSTQUEUE_REG_11__3__SCAN_IN, INSTQUEUE_REG_11__2__SCAN_IN, INSTQUEUE_REG_11__1__SCAN_IN, INSTQUEUE_REG_11__0__SCAN_IN, INSTQUEUE_REG_10__7__SCAN_IN, INSTQUEUE_REG_10__6__SCAN_IN, INSTQUEUE_REG_10__5__SCAN_IN, INSTQUEUE_REG_10__4__SCAN_IN, INSTQUEUE_REG_10__3__SCAN_IN, INSTQUEUE_REG_10__2__SCAN_IN, INSTQUEUE_REG_10__1__SCAN_IN, INSTQUEUE_REG_10__0__SCAN_IN, INSTQUEUE_REG_9__7__SCAN_IN, INSTQUEUE_REG_9__6__SCAN_IN, INSTQUEUE_REG_9__5__SCAN_IN, INSTQUEUE_REG_9__4__SCAN_IN, INSTQUEUE_REG_9__3__SCAN_IN, INSTQUEUE_REG_9__2__SCAN_IN, INSTQUEUE_REG_9__1__SCAN_IN, INSTQUEUE_REG_9__0__SCAN_IN, INSTQUEUE_REG_8__7__SCAN_IN, INSTQUEUE_REG_8__6__SCAN_IN, INSTQUEUE_REG_8__5__SCAN_IN, INSTQUEUE_REG_8__4__SCAN_IN, INSTQUEUE_REG_8__3__SCAN_IN, INSTQUEUE_REG_8__2__SCAN_IN, INSTQUEUE_REG_8__1__SCAN_IN, INSTQUEUE_REG_8__0__SCAN_IN, INSTQUEUE_REG_7__7__SCAN_IN, INSTQUEUE_REG_7__6__SCAN_IN, INSTQUEUE_REG_7__5__SCAN_IN, INSTQUEUE_REG_7__4__SCAN_IN, INSTQUEUE_REG_7__3__SCAN_IN, INSTQUEUE_REG_7__2__SCAN_IN, INSTQUEUE_REG_7__1__SCAN_IN, INSTQUEUE_REG_7__0__SCAN_IN, INSTQUEUE_REG_6__7__SCAN_IN, INSTQUEUE_REG_6__6__SCAN_IN, INSTQUEUE_REG_6__5__SCAN_IN, INSTQUEUE_REG_6__4__SCAN_IN, INSTQUEUE_REG_6__3__SCAN_IN, INSTQUEUE_REG_6__2__SCAN_IN, INSTQUEUE_REG_6__1__SCAN_IN, INSTQUEUE_REG_6__0__SCAN_IN, INSTQUEUE_REG_5__7__SCAN_IN, INSTQUEUE_REG_5__6__SCAN_IN, INSTQUEUE_REG_5__5__SCAN_IN, INSTQUEUE_REG_5__4__SCAN_IN, INSTQUEUE_REG_5__3__SCAN_IN, INSTQUEUE_REG_5__2__SCAN_IN, INSTQUEUE_REG_5__1__SCAN_IN, INSTQUEUE_REG_5__0__SCAN_IN, INSTQUEUE_REG_4__7__SCAN_IN, INSTQUEUE_REG_4__6__SCAN_IN, INSTQUEUE_REG_4__5__SCAN_IN, INSTQUEUE_REG_4__4__SCAN_IN, INSTQUEUE_REG_4__3__SCAN_IN, INSTQUEUE_REG_4__2__SCAN_IN, INSTQUEUE_REG_4__1__SCAN_IN, INSTQUEUE_REG_4__0__SCAN_IN, INSTQUEUE_REG_3__7__SCAN_IN, INSTQUEUE_REG_3__6__SCAN_IN, INSTQUEUE_REG_3__5__SCAN_IN, INSTQUEUE_REG_3__4__SCAN_IN, INSTQUEUE_REG_3__3__SCAN_IN, INSTQUEUE_REG_3__2__SCAN_IN, INSTQUEUE_REG_3__1__SCAN_IN, INSTQUEUE_REG_3__0__SCAN_IN, INSTQUEUE_REG_2__7__SCAN_IN, INSTQUEUE_REG_2__6__SCAN_IN, INSTQUEUE_REG_2__5__SCAN_IN, INSTQUEUE_REG_2__4__SCAN_IN, INSTQUEUE_REG_2__3__SCAN_IN, INSTQUEUE_REG_2__2__SCAN_IN, INSTQUEUE_REG_2__1__SCAN_IN, INSTQUEUE_REG_2__0__SCAN_IN, INSTQUEUE_REG_1__7__SCAN_IN, INSTQUEUE_REG_1__6__SCAN_IN, INSTQUEUE_REG_1__5__SCAN_IN, INSTQUEUE_REG_1__4__SCAN_IN, INSTQUEUE_REG_1__3__SCAN_IN, INSTQUEUE_REG_1__2__SCAN_IN, INSTQUEUE_REG_1__1__SCAN_IN, INSTQUEUE_REG_1__0__SCAN_IN, INSTQUEUE_REG_0__7__SCAN_IN, INSTQUEUE_REG_0__6__SCAN_IN, INSTQUEUE_REG_0__5__SCAN_IN, INSTQUEUE_REG_0__4__SCAN_IN, INSTQUEUE_REG_0__3__SCAN_IN, INSTQUEUE_REG_0__2__SCAN_IN, INSTQUEUE_REG_0__1__SCAN_IN, INSTQUEUE_REG_0__0__SCAN_IN, INSTQUEUERD_ADDR_REG_4__SCAN_IN, INSTQUEUERD_ADDR_REG_3__SCAN_IN, INSTQUEUERD_ADDR_REG_2__SCAN_IN, INSTQUEUERD_ADDR_REG_1__SCAN_IN, INSTQUEUERD_ADDR_REG_0__SCAN_IN, INSTQUEUEWR_ADDR_REG_4__SCAN_IN, INSTQUEUEWR_ADDR_REG_3__SCAN_IN, INSTQUEUEWR_ADDR_REG_2__SCAN_IN, INSTQUEUEWR_ADDR_REG_1__SCAN_IN, INSTQUEUEWR_ADDR_REG_0__SCAN_IN, INSTADDRPOINTER_REG_0__SCAN_IN, INSTADDRPOINTER_REG_1__SCAN_IN, INSTADDRPOINTER_REG_2__SCAN_IN, INSTADDRPOINTER_REG_3__SCAN_IN, INSTADDRPOINTER_REG_4__SCAN_IN, INSTADDRPOINTER_REG_5__SCAN_IN, INSTADDRPOINTER_REG_6__SCAN_IN, INSTADDRPOINTER_REG_7__SCAN_IN, INSTADDRPOINTER_REG_8__SCAN_IN, INSTADDRPOINTER_REG_9__SCAN_IN, INSTADDRPOINTER_REG_10__SCAN_IN, INSTADDRPOINTER_REG_11__SCAN_IN, INSTADDRPOINTER_REG_12__SCAN_IN, INSTADDRPOINTER_REG_13__SCAN_IN, INSTADDRPOINTER_REG_14__SCAN_IN, INSTADDRPOINTER_REG_15__SCAN_IN, INSTADDRPOINTER_REG_16__SCAN_IN, INSTADDRPOINTER_REG_17__SCAN_IN, INSTADDRPOINTER_REG_18__SCAN_IN, INSTADDRPOINTER_REG_19__SCAN_IN, INSTADDRPOINTER_REG_20__SCAN_IN, INSTADDRPOINTER_REG_21__SCAN_IN, INSTADDRPOINTER_REG_22__SCAN_IN, INSTADDRPOINTER_REG_23__SCAN_IN, INSTADDRPOINTER_REG_24__SCAN_IN, INSTADDRPOINTER_REG_25__SCAN_IN, INSTADDRPOINTER_REG_26__SCAN_IN, INSTADDRPOINTER_REG_27__SCAN_IN, INSTADDRPOINTER_REG_28__SCAN_IN, INSTADDRPOINTER_REG_29__SCAN_IN, INSTADDRPOINTER_REG_30__SCAN_IN, INSTADDRPOINTER_REG_31__SCAN_IN, PHYADDRPOINTER_REG_0__SCAN_IN, PHYADDRPOINTER_REG_1__SCAN_IN, PHYADDRPOINTER_REG_2__SCAN_IN, PHYADDRPOINTER_REG_3__SCAN_IN, PHYADDRPOINTER_REG_4__SCAN_IN, PHYADDRPOINTER_REG_5__SCAN_IN, PHYADDRPOINTER_REG_6__SCAN_IN, PHYADDRPOINTER_REG_7__SCAN_IN, PHYADDRPOINTER_REG_8__SCAN_IN, PHYADDRPOINTER_REG_9__SCAN_IN, PHYADDRPOINTER_REG_10__SCAN_IN, PHYADDRPOINTER_REG_11__SCAN_IN, PHYADDRPOINTER_REG_12__SCAN_IN, PHYADDRPOINTER_REG_13__SCAN_IN, PHYADDRPOINTER_REG_14__SCAN_IN, PHYADDRPOINTER_REG_15__SCAN_IN, PHYADDRPOINTER_REG_16__SCAN_IN, PHYADDRPOINTER_REG_17__SCAN_IN, PHYADDRPOINTER_REG_18__SCAN_IN, PHYADDRPOINTER_REG_19__SCAN_IN, PHYADDRPOINTER_REG_20__SCAN_IN, PHYADDRPOINTER_REG_21__SCAN_IN, PHYADDRPOINTER_REG_22__SCAN_IN, PHYADDRPOINTER_REG_23__SCAN_IN, PHYADDRPOINTER_REG_24__SCAN_IN, PHYADDRPOINTER_REG_25__SCAN_IN, PHYADDRPOINTER_REG_26__SCAN_IN, PHYADDRPOINTER_REG_27__SCAN_IN, PHYADDRPOINTER_REG_28__SCAN_IN, PHYADDRPOINTER_REG_29__SCAN_IN, PHYADDRPOINTER_REG_30__SCAN_IN, PHYADDRPOINTER_REG_31__SCAN_IN, LWORD_REG_15__SCAN_IN, LWORD_REG_14__SCAN_IN, LWORD_REG_13__SCAN_IN, LWORD_REG_12__SCAN_IN, LWORD_REG_11__SCAN_IN, LWORD_REG_10__SCAN_IN, LWORD_REG_9__SCAN_IN, LWORD_REG_8__SCAN_IN, LWORD_REG_7__SCAN_IN, LWORD_REG_6__SCAN_IN, LWORD_REG_5__SCAN_IN, LWORD_REG_4__SCAN_IN, LWORD_REG_3__SCAN_IN, LWORD_REG_2__SCAN_IN, LWORD_REG_1__SCAN_IN, LWORD_REG_0__SCAN_IN, UWORD_REG_14__SCAN_IN, UWORD_REG_13__SCAN_IN, UWORD_REG_12__SCAN_IN, UWORD_REG_11__SCAN_IN, UWORD_REG_10__SCAN_IN, UWORD_REG_9__SCAN_IN, UWORD_REG_8__SCAN_IN, UWORD_REG_7__SCAN_IN, UWORD_REG_6__SCAN_IN, UWORD_REG_5__SCAN_IN, UWORD_REG_4__SCAN_IN, UWORD_REG_3__SCAN_IN, UWORD_REG_2__SCAN_IN, UWORD_REG_1__SCAN_IN, UWORD_REG_0__SCAN_IN, EAX_REG_0__SCAN_IN, EAX_REG_1__SCAN_IN, EAX_REG_2__SCAN_IN, EAX_REG_3__SCAN_IN, EAX_REG_4__SCAN_IN, EAX_REG_5__SCAN_IN, EAX_REG_6__SCAN_IN, EAX_REG_7__SCAN_IN, EAX_REG_8__SCAN_IN, EAX_REG_9__SCAN_IN, EAX_REG_10__SCAN_IN, EAX_REG_11__SCAN_IN, EAX_REG_12__SCAN_IN, EAX_REG_13__SCAN_IN, EAX_REG_14__SCAN_IN, EAX_REG_15__SCAN_IN, EAX_REG_16__SCAN_IN, EAX_REG_17__SCAN_IN, EAX_REG_18__SCAN_IN, EAX_REG_19__SCAN_IN, EAX_REG_20__SCAN_IN, EAX_REG_21__SCAN_IN, EAX_REG_22__SCAN_IN, EAX_REG_23__SCAN_IN, EAX_REG_24__SCAN_IN, EAX_REG_25__SCAN_IN, EAX_REG_26__SCAN_IN, EAX_REG_27__SCAN_IN, EAX_REG_28__SCAN_IN, EAX_REG_29__SCAN_IN, EAX_REG_30__SCAN_IN, EAX_REG_31__SCAN_IN, EBX_REG_0__SCAN_IN, EBX_REG_1__SCAN_IN, EBX_REG_2__SCAN_IN, EBX_REG_3__SCAN_IN, EBX_REG_4__SCAN_IN, EBX_REG_5__SCAN_IN, EBX_REG_6__SCAN_IN, EBX_REG_7__SCAN_IN, EBX_REG_8__SCAN_IN, EBX_REG_9__SCAN_IN, EBX_REG_10__SCAN_IN, EBX_REG_11__SCAN_IN, EBX_REG_12__SCAN_IN, EBX_REG_13__SCAN_IN, EBX_REG_14__SCAN_IN, EBX_REG_15__SCAN_IN, EBX_REG_16__SCAN_IN, EBX_REG_17__SCAN_IN, EBX_REG_18__SCAN_IN, EBX_REG_19__SCAN_IN, EBX_REG_20__SCAN_IN, EBX_REG_21__SCAN_IN, EBX_REG_22__SCAN_IN, EBX_REG_23__SCAN_IN, EBX_REG_24__SCAN_IN, EBX_REG_25__SCAN_IN, EBX_REG_26__SCAN_IN, EBX_REG_27__SCAN_IN, EBX_REG_28__SCAN_IN, EBX_REG_29__SCAN_IN, EBX_REG_30__SCAN_IN, EBX_REG_31__SCAN_IN, REIP_REG_0__SCAN_IN, REIP_REG_1__SCAN_IN, REIP_REG_2__SCAN_IN, REIP_REG_3__SCAN_IN, REIP_REG_4__SCAN_IN, REIP_REG_5__SCAN_IN, REIP_REG_6__SCAN_IN, REIP_REG_7__SCAN_IN, REIP_REG_8__SCAN_IN, REIP_REG_9__SCAN_IN, REIP_REG_10__SCAN_IN, REIP_REG_11__SCAN_IN, REIP_REG_12__SCAN_IN, REIP_REG_13__SCAN_IN, REIP_REG_14__SCAN_IN, REIP_REG_15__SCAN_IN, keyinput0, keyinput1, keyinput2, keyinput3, keyinput4, keyinput5, keyinput6, keyinput7, keyinput8, keyinput9, keyinput10, keyinput11, keyinput12, keyinput13, keyinput14, keyinput15, keyinput16, keyinput17, keyinput18, keyinput19, keyinput20, keyinput21, keyinput22, keyinput23, keyinput24, keyinput25, keyinput26, keyinput27, keyinput28, keyinput29, keyinput30, keyinput31;
  output DATAO_REG_2__SCAN_IN_BUFF, ADDRESS_REG_17__SCAN_IN_BUFF, DATAO_REG_22__SCAN_IN_BUFF, U3460, U3176, U2834, U3097, U2809, U3464, U3119, U2938, U3124, U2992, U2920, U2884, U3122, U3179, U2853, U3107, U3055, U3011, U2891, U2830, ADDRESS_REG_2__SCAN_IN_BUFF, U2797, U2869, U3043, U2958, U3105, U3013, U3077, U3059, BE_N_REG_0__SCAN_IN_BUFF, ADDRESS_REG_9__SCAN_IN_BUFF, ADDRESS_REG_11__SCAN_IN_BUFF, U3199, U3141, ADDRESS_REG_22__SCAN_IN_BUFF, U2789, U3149, U2917, U3169, U2981, U2941, U2892, U3093, ADDRESS_REG_0__SCAN_IN_BUFF, U3003, U2906, U2875, ADDRESS_REG_6__SCAN_IN_BUFF, U2854, U3132, U3032, DATAO_REG_24__SCAN_IN_BUFF, U2872, ADDRESS_REG_3__SCAN_IN_BUFF, U3136, U3071, U2896, U3451, U3168, U3079, U2795, U2829, U2840, U2868, U3082, U2928, U2915, U3148, U2990, U3160, ADDRESS_REG_21__SCAN_IN_BUFF, U3024, U2864, U2803, U2844, U2889, U2852, U3147, U2914, U3034, U2876, U3062, U2972, U3050, U2828, U2951, W_R_N_REG_SCAN_IN_BUFF, U3014, DATAO_REG_1__SCAN_IN_BUFF, U3064, U2819, U2961, U3015, U3085, ADDRESS_REG_5__SCAN_IN_BUFF, U3208, U3027, U2993, U2987, U3201, DATAO_REG_9__SCAN_IN_BUFF, U2960, U3049, U2825, U2979, U3028, DATAO_REG_15__SCAN_IN_BUFF, U2957, U2971, U2850, U3095, U2977, U3041, U2837, U3452, U3052, ADDRESS_REG_8__SCAN_IN_BUFF, U2926, DATAO_REG_26__SCAN_IN_BUFF, U3157, U2973, DATAO_REG_29__SCAN_IN_BUFF, U3170, U3152, U3159, U3196, U3089, U2897, U3469, U2921, U2870, U3069, U3063, U3135, U3166, U3210, U3153, U2818, U2905, U2933, U2796, U3207, U2898, U3209, U3078, U2946, U2907, BE_N_REG_3__SCAN_IN_BUFF, U2943, U2866, U2881, U2976, U2899, U3175, U3180, DATAO_REG_14__SCAN_IN_BUFF, U3113, M_IO_N_REG_SCAN_IN_BUFF, U2843, U2877, U2919, U3100, U2916, U2934, DATAO_REG_12__SCAN_IN_BUFF, U3146, U2924, U3161, U3005, U2893, U2945, U3470, U3150, U3109, U3213, U2955, U3448, U3194, U2832, U2978, U3183, U2947, DATAO_REG_3__SCAN_IN_BUFF, ADDRESS_REG_15__SCAN_IN_BUFF, U3007, U3162, U3203, U3106, U2942, ADDRESS_REG_18__SCAN_IN_BUFF, U3035, U2975, U2820, U2969, U2963, U2909, U3140, U2925, U2983, U2967, U2805, U3021, U3054, U3092, U3173, U2790, U2871, U2922, U2988, U3156, ADDRESS_REG_23__SCAN_IN_BUFF, U2932, U2822, U2878, U3155, U3010, U2935, U2794, U3033, U3030, U2835, U3186, U2824, U2956, U3163, U2831, U3026, U3083, U2814, U2953, U2890, U2882, U2791, U3000, U2998, ADDRESS_REG_26__SCAN_IN_BUFF, ADDRESS_REG_27__SCAN_IN_BUFF, U3125, U2817, U3101, U2900, U2793, DATAO_REG_25__SCAN_IN_BUFF, U2995, U2985, U3121, U3009, U3099, U2952, DATAO_REG_13__SCAN_IN_BUFF, U3133, U2806, U2962, U2948, U2888, U3456, U3462, U3115, U2801, U3158, U2865, U3185, U3110, U3145, U2940, U3167, ADDRESS_REG_29__SCAN_IN_BUFF, U2863, U3174, U3198, U2813, U3057, U3459, U3068, U2827, U3154, U2901, DATAO_REG_21__SCAN_IN_BUFF, U2903, U2855, U3098, U3025, U3205, U2838, U3211, U3067, U2841, U2959, U3463, U2800, DATAO_REG_18__SCAN_IN_BUFF, U3118, DATAO_REG_23__SCAN_IN_BUFF, U2859, U3130, U2860, U3036, U3045, U3066, U3017, U2826, U3023, U2821, U2989, ADDRESS_REG_12__SCAN_IN_BUFF, U3206, U3190, U2918, BE_N_REG_2__SCAN_IN_BUFF, U3102, DATAO_REG_28__SCAN_IN_BUFF, U3472, U3193, U3151, U2858, U2931, U2912, U3129, U3137, U2804, U2846, U3461, U3037, U3202, U3084, U3002, U3143, U2815, U2845, DATAO_REG_5__SCAN_IN_BUFF, U2902, U2930, DATAO_REG_31__SCAN_IN_BUFF, ADDRESS_REG_4__SCAN_IN_BUFF, ADDRESS_REG_25__SCAN_IN_BUFF, DATAO_REG_16__SCAN_IN_BUFF, U3172, U3038, U3018, U2910, U2883, DATAO_REG_30__SCAN_IN_BUFF, U2939, U3103, U3075, U2894, U3001, U3114, U3060, U3039, DATAO_REG_7__SCAN_IN_BUFF, DATAO_REG_19__SCAN_IN_BUFF, U2799, U3047, U2879, DATAO_REG_17__SCAN_IN_BUFF, U2857, U2911, U2880, U2937, U2812, U3008, U2839, U3111, U2904, U3445, DATAO_REG_8__SCAN_IN_BUFF, U3029, U2974, U2810, U2833, U3447, U2982, DATAO_REG_20__SCAN_IN_BUFF, ADS_N_REG_SCAN_IN_BUFF, U3204, U3184, U3200, U2851, U2798, U3019, U2885, U3104, U3065, U3164, U3070, U3453, U3061, U3087, U3108, ADDRESS_REG_10__SCAN_IN_BUFF, U3127, U2867, U3138, DATAO_REG_0__SCAN_IN_BUFF, U2856, U3046, U3139, U3051, U3465, U2811, U3073, U3474, U3116, U3086, U3016, U3126, U3446, U2923, U2816, U2970, U3004, U3006, U3081, U2788, U2842, U2874, U2802, U2886, U2964, ADDRESS_REG_28__SCAN_IN_BUFF, U3020, U2913, U2895, DATAO_REG_4__SCAN_IN_BUFF, U2836, U2823, U2849, U2862, U3088, U3044, U2848, U3177, U2873, U2966, U2861, U3187, U3117, U2984, U3191, U3074, U3212, U2887, U3076, U2929, U3182, U2927, U3195, U3178, U2986, ADDRESS_REG_7__SCAN_IN_BUFF, ADDRESS_REG_13__SCAN_IN_BUFF, U3189, U2950, U3090, U3053, U2980, U3171, U3080, U2954, U2944, U3165, U3123, U3022, U3120, DATAO_REG_6__SCAN_IN_BUFF, U3072, DATAO_REG_27__SCAN_IN_BUFF, ADDRESS_REG_20__SCAN_IN_BUFF, U2968, U3144, U3134, U2847, U2994, U2936, DATAO_REG_11__SCAN_IN_BUFF, U3192, U2991, U2908, U2965, U3131, ADDRESS_REG_24__SCAN_IN_BUFF, U3181, U3040, U3197, DATAO_REG_10__SCAN_IN_BUFF, U3091, ADDRESS_REG_1__SCAN_IN_BUFF, U3112, U3042, U3188, D_C_N_REG_SCAN_IN_BUFF, U2808, ADDRESS_REG_14__SCAN_IN_BUFF, U3094, U3142, U2792, U2996, U3473, U3012, U3468, U2999, ADDRESS_REG_19__SCAN_IN_BUFF, U3471, U3058, BE_N_REG_1__SCAN_IN_BUFF, U3031, U2807, U2949, U2997, U3455, U3128, U3048, U3096, ADDRESS_REG_16__SCAN_IN_BUFF, U3056;
  wire perturb_signal, restore_signal;

  b15_C_SFLL_HD_4_32_1 main (DATAO_REG_25__SCAN_IN, DATAO_REG_5__SCAN_IN, DATAO_REG_28__SCAN_IN, DATAO_REG_21__SCAN_IN, BE_N_REG_0__SCAN_IN, ADDRESS_REG_23__SCAN_IN, ADDRESS_REG_17__SCAN_IN, ADDRESS_REG_2__SCAN_IN, DATAO_REG_30__SCAN_IN, BE_N_REG_1__SCAN_IN, ADDRESS_REG_1__SCAN_IN, DATAO_REG_8__SCAN_IN, DATAO_REG_23__SCAN_IN, DATAO_REG_10__SCAN_IN, ADDRESS_REG_22__SCAN_IN, ADDRESS_REG_11__SCAN_IN, ADDRESS_REG_3__SCAN_IN, BE_N_REG_3__SCAN_IN, DATAO_REG_27__SCAN_IN, ADDRESS_REG_10__SCAN_IN, ADDRESS_REG_28__SCAN_IN, DATAO_REG_12__SCAN_IN, BE_N_REG_2__SCAN_IN, ADDRESS_REG_13__SCAN_IN, DATAO_REG_13__SCAN_IN, ADDRESS_REG_20__SCAN_IN, DATAO_REG_24__SCAN_IN, DATAO_REG_9__SCAN_IN, DATAO_REG_7__SCAN_IN, DATAO_REG_11__SCAN_IN, ADDRESS_REG_19__SCAN_IN, ADDRESS_REG_27__SCAN_IN, ADDRESS_REG_25__SCAN_IN, ADDRESS_REG_29__SCAN_IN, ADDRESS_REG_5__SCAN_IN, ADDRESS_REG_7__SCAN_IN, ADDRESS_REG_8__SCAN_IN, ADDRESS_REG_21__SCAN_IN, DATAO_REG_20__SCAN_IN, DATAO_REG_17__SCAN_IN, DATAO_REG_6__SCAN_IN, ADDRESS_REG_14__SCAN_IN, DATAO_REG_19__SCAN_IN, ADS_N_REG_SCAN_IN, DATAO_REG_15__SCAN_IN, DATAO_REG_26__SCAN_IN, DATAO_REG_3__SCAN_IN, DATAO_REG_1__SCAN_IN, ADDRESS_REG_26__SCAN_IN, ADDRESS_REG_18__SCAN_IN, M_IO_N_REG_SCAN_IN, DATAO_REG_31__SCAN_IN, ADDRESS_REG_16__SCAN_IN, ADDRESS_REG_9__SCAN_IN, ADDRESS_REG_12__SCAN_IN, DATAO_REG_29__SCAN_IN, DATAO_REG_0__SCAN_IN, ADDRESS_REG_4__SCAN_IN, D_C_N_REG_SCAN_IN, DATAO_REG_4__SCAN_IN, ADDRESS_REG_6__SCAN_IN, DATAO_REG_2__SCAN_IN, ADDRESS_REG_0__SCAN_IN, DATAO_REG_18__SCAN_IN, DATAO_REG_16__SCAN_IN, ADDRESS_REG_24__SCAN_IN, DATAO_REG_14__SCAN_IN, W_R_N_REG_SCAN_IN, ADDRESS_REG_15__SCAN_IN, DATAO_REG_22__SCAN_IN, DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, DATAI_27_, DATAI_26_, DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, DATAI_21_, DATAI_20_, DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, DATAI_15_, DATAI_14_, DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, DATAI_9_, DATAI_8_, DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, DATAI_2_, DATAI_1_, DATAI_0_, MEMORYFETCH_REG_SCAN_IN, NA_N, BS16_N, READY_N, HOLD, READREQUEST_REG_SCAN_IN, CODEFETCH_REG_SCAN_IN, REQUESTPENDING_REG_SCAN_IN, STATEBS16_REG_SCAN_IN, MORE_REG_SCAN_IN, FLUSH_REG_SCAN_IN, BYTEENABLE_REG_0__SCAN_IN, BYTEENABLE_REG_1__SCAN_IN, BYTEENABLE_REG_2__SCAN_IN, BYTEENABLE_REG_3__SCAN_IN, REIP_REG_31__SCAN_IN, REIP_REG_30__SCAN_IN, REIP_REG_29__SCAN_IN, REIP_REG_28__SCAN_IN, REIP_REG_27__SCAN_IN, REIP_REG_26__SCAN_IN, REIP_REG_25__SCAN_IN, REIP_REG_24__SCAN_IN, REIP_REG_23__SCAN_IN, REIP_REG_22__SCAN_IN, REIP_REG_21__SCAN_IN, REIP_REG_20__SCAN_IN, REIP_REG_19__SCAN_IN, REIP_REG_18__SCAN_IN, REIP_REG_17__SCAN_IN, REIP_REG_16__SCAN_IN, STATE_REG_2__SCAN_IN, STATE_REG_1__SCAN_IN, STATE_REG_0__SCAN_IN, DATAWIDTH_REG_0__SCAN_IN, DATAWIDTH_REG_1__SCAN_IN, DATAWIDTH_REG_2__SCAN_IN, DATAWIDTH_REG_3__SCAN_IN, DATAWIDTH_REG_4__SCAN_IN, DATAWIDTH_REG_5__SCAN_IN, DATAWIDTH_REG_6__SCAN_IN, DATAWIDTH_REG_7__SCAN_IN, DATAWIDTH_REG_8__SCAN_IN, DATAWIDTH_REG_9__SCAN_IN, DATAWIDTH_REG_10__SCAN_IN, DATAWIDTH_REG_11__SCAN_IN, DATAWIDTH_REG_12__SCAN_IN, DATAWIDTH_REG_13__SCAN_IN, DATAWIDTH_REG_14__SCAN_IN, DATAWIDTH_REG_15__SCAN_IN, DATAWIDTH_REG_16__SCAN_IN, DATAWIDTH_REG_17__SCAN_IN, DATAWIDTH_REG_18__SCAN_IN, DATAWIDTH_REG_19__SCAN_IN, DATAWIDTH_REG_20__SCAN_IN, DATAWIDTH_REG_21__SCAN_IN, DATAWIDTH_REG_22__SCAN_IN, DATAWIDTH_REG_23__SCAN_IN, DATAWIDTH_REG_24__SCAN_IN, DATAWIDTH_REG_25__SCAN_IN, DATAWIDTH_REG_26__SCAN_IN, DATAWIDTH_REG_27__SCAN_IN, DATAWIDTH_REG_28__SCAN_IN, DATAWIDTH_REG_29__SCAN_IN, DATAWIDTH_REG_30__SCAN_IN, DATAWIDTH_REG_31__SCAN_IN, STATE2_REG_3__SCAN_IN, STATE2_REG_2__SCAN_IN, STATE2_REG_1__SCAN_IN, STATE2_REG_0__SCAN_IN, INSTQUEUE_REG_15__7__SCAN_IN, INSTQUEUE_REG_15__6__SCAN_IN, INSTQUEUE_REG_15__5__SCAN_IN, INSTQUEUE_REG_15__4__SCAN_IN, INSTQUEUE_REG_15__3__SCAN_IN, INSTQUEUE_REG_15__2__SCAN_IN, INSTQUEUE_REG_15__1__SCAN_IN, INSTQUEUE_REG_15__0__SCAN_IN, INSTQUEUE_REG_14__7__SCAN_IN, INSTQUEUE_REG_14__6__SCAN_IN, INSTQUEUE_REG_14__5__SCAN_IN, INSTQUEUE_REG_14__4__SCAN_IN, INSTQUEUE_REG_14__3__SCAN_IN, INSTQUEUE_REG_14__2__SCAN_IN, INSTQUEUE_REG_14__1__SCAN_IN, INSTQUEUE_REG_14__0__SCAN_IN, INSTQUEUE_REG_13__7__SCAN_IN, INSTQUEUE_REG_13__6__SCAN_IN, INSTQUEUE_REG_13__5__SCAN_IN, INSTQUEUE_REG_13__4__SCAN_IN, INSTQUEUE_REG_13__3__SCAN_IN, INSTQUEUE_REG_13__2__SCAN_IN, INSTQUEUE_REG_13__1__SCAN_IN, INSTQUEUE_REG_13__0__SCAN_IN, INSTQUEUE_REG_12__7__SCAN_IN, INSTQUEUE_REG_12__6__SCAN_IN, INSTQUEUE_REG_12__5__SCAN_IN, INSTQUEUE_REG_12__4__SCAN_IN, INSTQUEUE_REG_12__3__SCAN_IN, INSTQUEUE_REG_12__2__SCAN_IN, INSTQUEUE_REG_12__1__SCAN_IN, INSTQUEUE_REG_12__0__SCAN_IN, INSTQUEUE_REG_11__7__SCAN_IN, INSTQUEUE_REG_11__6__SCAN_IN, INSTQUEUE_REG_11__5__SCAN_IN, INSTQUEUE_REG_11__4__SCAN_IN, INSTQUEUE_REG_11__3__SCAN_IN, INSTQUEUE_REG_11__2__SCAN_IN, INSTQUEUE_REG_11__1__SCAN_IN, INSTQUEUE_REG_11__0__SCAN_IN, INSTQUEUE_REG_10__7__SCAN_IN, INSTQUEUE_REG_10__6__SCAN_IN, INSTQUEUE_REG_10__5__SCAN_IN, INSTQUEUE_REG_10__4__SCAN_IN, INSTQUEUE_REG_10__3__SCAN_IN, INSTQUEUE_REG_10__2__SCAN_IN, INSTQUEUE_REG_10__1__SCAN_IN, INSTQUEUE_REG_10__0__SCAN_IN, INSTQUEUE_REG_9__7__SCAN_IN, INSTQUEUE_REG_9__6__SCAN_IN, INSTQUEUE_REG_9__5__SCAN_IN, INSTQUEUE_REG_9__4__SCAN_IN, INSTQUEUE_REG_9__3__SCAN_IN, INSTQUEUE_REG_9__2__SCAN_IN, INSTQUEUE_REG_9__1__SCAN_IN, INSTQUEUE_REG_9__0__SCAN_IN, INSTQUEUE_REG_8__7__SCAN_IN, INSTQUEUE_REG_8__6__SCAN_IN, INSTQUEUE_REG_8__5__SCAN_IN, INSTQUEUE_REG_8__4__SCAN_IN, INSTQUEUE_REG_8__3__SCAN_IN, INSTQUEUE_REG_8__2__SCAN_IN, INSTQUEUE_REG_8__1__SCAN_IN, INSTQUEUE_REG_8__0__SCAN_IN, INSTQUEUE_REG_7__7__SCAN_IN, INSTQUEUE_REG_7__6__SCAN_IN, INSTQUEUE_REG_7__5__SCAN_IN, INSTQUEUE_REG_7__4__SCAN_IN, INSTQUEUE_REG_7__3__SCAN_IN, INSTQUEUE_REG_7__2__SCAN_IN, INSTQUEUE_REG_7__1__SCAN_IN, INSTQUEUE_REG_7__0__SCAN_IN, INSTQUEUE_REG_6__7__SCAN_IN, INSTQUEUE_REG_6__6__SCAN_IN, INSTQUEUE_REG_6__5__SCAN_IN, INSTQUEUE_REG_6__4__SCAN_IN, INSTQUEUE_REG_6__3__SCAN_IN, INSTQUEUE_REG_6__2__SCAN_IN, INSTQUEUE_REG_6__1__SCAN_IN, INSTQUEUE_REG_6__0__SCAN_IN, INSTQUEUE_REG_5__7__SCAN_IN, INSTQUEUE_REG_5__6__SCAN_IN, INSTQUEUE_REG_5__5__SCAN_IN, INSTQUEUE_REG_5__4__SCAN_IN, INSTQUEUE_REG_5__3__SCAN_IN, INSTQUEUE_REG_5__2__SCAN_IN, INSTQUEUE_REG_5__1__SCAN_IN, INSTQUEUE_REG_5__0__SCAN_IN, INSTQUEUE_REG_4__7__SCAN_IN, INSTQUEUE_REG_4__6__SCAN_IN, INSTQUEUE_REG_4__5__SCAN_IN, INSTQUEUE_REG_4__4__SCAN_IN, INSTQUEUE_REG_4__3__SCAN_IN, INSTQUEUE_REG_4__2__SCAN_IN, INSTQUEUE_REG_4__1__SCAN_IN, INSTQUEUE_REG_4__0__SCAN_IN, INSTQUEUE_REG_3__7__SCAN_IN, INSTQUEUE_REG_3__6__SCAN_IN, INSTQUEUE_REG_3__5__SCAN_IN, INSTQUEUE_REG_3__4__SCAN_IN, INSTQUEUE_REG_3__3__SCAN_IN, INSTQUEUE_REG_3__2__SCAN_IN, INSTQUEUE_REG_3__1__SCAN_IN, INSTQUEUE_REG_3__0__SCAN_IN, INSTQUEUE_REG_2__7__SCAN_IN, INSTQUEUE_REG_2__6__SCAN_IN, INSTQUEUE_REG_2__5__SCAN_IN, INSTQUEUE_REG_2__4__SCAN_IN, INSTQUEUE_REG_2__3__SCAN_IN, INSTQUEUE_REG_2__2__SCAN_IN, INSTQUEUE_REG_2__1__SCAN_IN, INSTQUEUE_REG_2__0__SCAN_IN, INSTQUEUE_REG_1__7__SCAN_IN, INSTQUEUE_REG_1__6__SCAN_IN, INSTQUEUE_REG_1__5__SCAN_IN, INSTQUEUE_REG_1__4__SCAN_IN, INSTQUEUE_REG_1__3__SCAN_IN, INSTQUEUE_REG_1__2__SCAN_IN, INSTQUEUE_REG_1__1__SCAN_IN, INSTQUEUE_REG_1__0__SCAN_IN, INSTQUEUE_REG_0__7__SCAN_IN, INSTQUEUE_REG_0__6__SCAN_IN, INSTQUEUE_REG_0__5__SCAN_IN, INSTQUEUE_REG_0__4__SCAN_IN, INSTQUEUE_REG_0__3__SCAN_IN, INSTQUEUE_REG_0__2__SCAN_IN, INSTQUEUE_REG_0__1__SCAN_IN, INSTQUEUE_REG_0__0__SCAN_IN, INSTQUEUERD_ADDR_REG_4__SCAN_IN, INSTQUEUERD_ADDR_REG_3__SCAN_IN, INSTQUEUERD_ADDR_REG_2__SCAN_IN, INSTQUEUERD_ADDR_REG_1__SCAN_IN, INSTQUEUERD_ADDR_REG_0__SCAN_IN, INSTQUEUEWR_ADDR_REG_4__SCAN_IN, INSTQUEUEWR_ADDR_REG_3__SCAN_IN, INSTQUEUEWR_ADDR_REG_2__SCAN_IN, INSTQUEUEWR_ADDR_REG_1__SCAN_IN, INSTQUEUEWR_ADDR_REG_0__SCAN_IN, INSTADDRPOINTER_REG_0__SCAN_IN, INSTADDRPOINTER_REG_1__SCAN_IN, INSTADDRPOINTER_REG_2__SCAN_IN, INSTADDRPOINTER_REG_3__SCAN_IN, INSTADDRPOINTER_REG_4__SCAN_IN, INSTADDRPOINTER_REG_5__SCAN_IN, INSTADDRPOINTER_REG_6__SCAN_IN, INSTADDRPOINTER_REG_7__SCAN_IN, INSTADDRPOINTER_REG_8__SCAN_IN, INSTADDRPOINTER_REG_9__SCAN_IN, INSTADDRPOINTER_REG_10__SCAN_IN, INSTADDRPOINTER_REG_11__SCAN_IN, INSTADDRPOINTER_REG_12__SCAN_IN, INSTADDRPOINTER_REG_13__SCAN_IN, INSTADDRPOINTER_REG_14__SCAN_IN, INSTADDRPOINTER_REG_15__SCAN_IN, INSTADDRPOINTER_REG_16__SCAN_IN, INSTADDRPOINTER_REG_17__SCAN_IN, INSTADDRPOINTER_REG_18__SCAN_IN, INSTADDRPOINTER_REG_19__SCAN_IN, INSTADDRPOINTER_REG_20__SCAN_IN, INSTADDRPOINTER_REG_21__SCAN_IN, INSTADDRPOINTER_REG_22__SCAN_IN, INSTADDRPOINTER_REG_23__SCAN_IN, INSTADDRPOINTER_REG_24__SCAN_IN, INSTADDRPOINTER_REG_25__SCAN_IN, INSTADDRPOINTER_REG_26__SCAN_IN, INSTADDRPOINTER_REG_27__SCAN_IN, INSTADDRPOINTER_REG_28__SCAN_IN, INSTADDRPOINTER_REG_29__SCAN_IN, INSTADDRPOINTER_REG_30__SCAN_IN, INSTADDRPOINTER_REG_31__SCAN_IN, PHYADDRPOINTER_REG_0__SCAN_IN, PHYADDRPOINTER_REG_1__SCAN_IN, PHYADDRPOINTER_REG_2__SCAN_IN, PHYADDRPOINTER_REG_3__SCAN_IN, PHYADDRPOINTER_REG_4__SCAN_IN, PHYADDRPOINTER_REG_5__SCAN_IN, PHYADDRPOINTER_REG_6__SCAN_IN, PHYADDRPOINTER_REG_7__SCAN_IN, PHYADDRPOINTER_REG_8__SCAN_IN, PHYADDRPOINTER_REG_9__SCAN_IN, PHYADDRPOINTER_REG_10__SCAN_IN, PHYADDRPOINTER_REG_11__SCAN_IN, PHYADDRPOINTER_REG_12__SCAN_IN, PHYADDRPOINTER_REG_13__SCAN_IN, PHYADDRPOINTER_REG_14__SCAN_IN, PHYADDRPOINTER_REG_15__SCAN_IN, PHYADDRPOINTER_REG_16__SCAN_IN, PHYADDRPOINTER_REG_17__SCAN_IN, PHYADDRPOINTER_REG_18__SCAN_IN, PHYADDRPOINTER_REG_19__SCAN_IN, PHYADDRPOINTER_REG_20__SCAN_IN, PHYADDRPOINTER_REG_21__SCAN_IN, PHYADDRPOINTER_REG_22__SCAN_IN, PHYADDRPOINTER_REG_23__SCAN_IN, PHYADDRPOINTER_REG_24__SCAN_IN, PHYADDRPOINTER_REG_25__SCAN_IN, PHYADDRPOINTER_REG_26__SCAN_IN, PHYADDRPOINTER_REG_27__SCAN_IN, PHYADDRPOINTER_REG_28__SCAN_IN, PHYADDRPOINTER_REG_29__SCAN_IN, PHYADDRPOINTER_REG_30__SCAN_IN, PHYADDRPOINTER_REG_31__SCAN_IN, LWORD_REG_15__SCAN_IN, LWORD_REG_14__SCAN_IN, LWORD_REG_13__SCAN_IN, LWORD_REG_12__SCAN_IN, LWORD_REG_11__SCAN_IN, LWORD_REG_10__SCAN_IN, LWORD_REG_9__SCAN_IN, LWORD_REG_8__SCAN_IN, LWORD_REG_7__SCAN_IN, LWORD_REG_6__SCAN_IN, LWORD_REG_5__SCAN_IN, LWORD_REG_4__SCAN_IN, LWORD_REG_3__SCAN_IN, LWORD_REG_2__SCAN_IN, LWORD_REG_1__SCAN_IN, LWORD_REG_0__SCAN_IN, UWORD_REG_14__SCAN_IN, UWORD_REG_13__SCAN_IN, UWORD_REG_12__SCAN_IN, UWORD_REG_11__SCAN_IN, UWORD_REG_10__SCAN_IN, UWORD_REG_9__SCAN_IN, UWORD_REG_8__SCAN_IN, UWORD_REG_7__SCAN_IN, UWORD_REG_6__SCAN_IN, UWORD_REG_5__SCAN_IN, UWORD_REG_4__SCAN_IN, UWORD_REG_3__SCAN_IN, UWORD_REG_2__SCAN_IN, UWORD_REG_1__SCAN_IN, UWORD_REG_0__SCAN_IN, EAX_REG_0__SCAN_IN, EAX_REG_1__SCAN_IN, EAX_REG_2__SCAN_IN, EAX_REG_3__SCAN_IN, EAX_REG_4__SCAN_IN, EAX_REG_5__SCAN_IN, EAX_REG_6__SCAN_IN, EAX_REG_7__SCAN_IN, EAX_REG_8__SCAN_IN, EAX_REG_9__SCAN_IN, EAX_REG_10__SCAN_IN, EAX_REG_11__SCAN_IN, EAX_REG_12__SCAN_IN, EAX_REG_13__SCAN_IN, EAX_REG_14__SCAN_IN, EAX_REG_15__SCAN_IN, EAX_REG_16__SCAN_IN, EAX_REG_17__SCAN_IN, EAX_REG_18__SCAN_IN, EAX_REG_19__SCAN_IN, EAX_REG_20__SCAN_IN, EAX_REG_21__SCAN_IN, EAX_REG_22__SCAN_IN, EAX_REG_23__SCAN_IN, EAX_REG_24__SCAN_IN, EAX_REG_25__SCAN_IN, EAX_REG_26__SCAN_IN, EAX_REG_27__SCAN_IN, EAX_REG_28__SCAN_IN, EAX_REG_29__SCAN_IN, EAX_REG_30__SCAN_IN, EAX_REG_31__SCAN_IN, EBX_REG_0__SCAN_IN, EBX_REG_1__SCAN_IN, EBX_REG_2__SCAN_IN, EBX_REG_3__SCAN_IN, EBX_REG_4__SCAN_IN, EBX_REG_5__SCAN_IN, EBX_REG_6__SCAN_IN, EBX_REG_7__SCAN_IN, EBX_REG_8__SCAN_IN, EBX_REG_9__SCAN_IN, EBX_REG_10__SCAN_IN, EBX_REG_11__SCAN_IN, EBX_REG_12__SCAN_IN, EBX_REG_13__SCAN_IN, EBX_REG_14__SCAN_IN, EBX_REG_15__SCAN_IN, EBX_REG_16__SCAN_IN, EBX_REG_17__SCAN_IN, EBX_REG_18__SCAN_IN, EBX_REG_19__SCAN_IN, EBX_REG_20__SCAN_IN, EBX_REG_21__SCAN_IN, EBX_REG_22__SCAN_IN, EBX_REG_23__SCAN_IN, EBX_REG_24__SCAN_IN, EBX_REG_25__SCAN_IN, EBX_REG_26__SCAN_IN, EBX_REG_27__SCAN_IN, EBX_REG_28__SCAN_IN, EBX_REG_29__SCAN_IN, EBX_REG_30__SCAN_IN, EBX_REG_31__SCAN_IN, REIP_REG_0__SCAN_IN, REIP_REG_1__SCAN_IN, REIP_REG_2__SCAN_IN, REIP_REG_3__SCAN_IN, REIP_REG_4__SCAN_IN, REIP_REG_5__SCAN_IN, REIP_REG_6__SCAN_IN, REIP_REG_7__SCAN_IN, REIP_REG_8__SCAN_IN, REIP_REG_9__SCAN_IN, REIP_REG_10__SCAN_IN, REIP_REG_11__SCAN_IN, REIP_REG_12__SCAN_IN, REIP_REG_13__SCAN_IN, REIP_REG_14__SCAN_IN, REIP_REG_15__SCAN_IN, perturb_signal, restore_signal, DATAO_REG_25__SCAN_IN_BUFF, DATAO_REG_5__SCAN_IN_BUFF, DATAO_REG_28__SCAN_IN_BUFF, DATAO_REG_21__SCAN_IN_BUFF, BE_N_REG_0__SCAN_IN_BUFF, ADDRESS_REG_23__SCAN_IN_BUFF, ADDRESS_REG_17__SCAN_IN_BUFF, ADDRESS_REG_2__SCAN_IN_BUFF, DATAO_REG_30__SCAN_IN_BUFF, BE_N_REG_1__SCAN_IN_BUFF, ADDRESS_REG_1__SCAN_IN_BUFF, DATAO_REG_8__SCAN_IN_BUFF, DATAO_REG_23__SCAN_IN_BUFF, DATAO_REG_10__SCAN_IN_BUFF, ADDRESS_REG_22__SCAN_IN_BUFF, ADDRESS_REG_11__SCAN_IN_BUFF, ADDRESS_REG_3__SCAN_IN_BUFF, BE_N_REG_3__SCAN_IN_BUFF, DATAO_REG_27__SCAN_IN_BUFF, ADDRESS_REG_10__SCAN_IN_BUFF, ADDRESS_REG_28__SCAN_IN_BUFF, DATAO_REG_12__SCAN_IN_BUFF, BE_N_REG_2__SCAN_IN_BUFF, ADDRESS_REG_13__SCAN_IN_BUFF, DATAO_REG_13__SCAN_IN_BUFF, ADDRESS_REG_20__SCAN_IN_BUFF, DATAO_REG_24__SCAN_IN_BUFF, DATAO_REG_9__SCAN_IN_BUFF, DATAO_REG_7__SCAN_IN_BUFF, DATAO_REG_11__SCAN_IN_BUFF, ADDRESS_REG_19__SCAN_IN_BUFF, ADDRESS_REG_27__SCAN_IN_BUFF, ADDRESS_REG_25__SCAN_IN_BUFF, ADDRESS_REG_29__SCAN_IN_BUFF, ADDRESS_REG_5__SCAN_IN_BUFF, ADDRESS_REG_7__SCAN_IN_BUFF, ADDRESS_REG_8__SCAN_IN_BUFF, ADDRESS_REG_21__SCAN_IN_BUFF, DATAO_REG_20__SCAN_IN_BUFF, DATAO_REG_17__SCAN_IN_BUFF, DATAO_REG_6__SCAN_IN_BUFF, ADDRESS_REG_14__SCAN_IN_BUFF, DATAO_REG_19__SCAN_IN_BUFF, ADS_N_REG_SCAN_IN_BUFF, DATAO_REG_15__SCAN_IN_BUFF, DATAO_REG_26__SCAN_IN_BUFF, DATAO_REG_3__SCAN_IN_BUFF, DATAO_REG_1__SCAN_IN_BUFF, ADDRESS_REG_26__SCAN_IN_BUFF, ADDRESS_REG_18__SCAN_IN_BUFF, M_IO_N_REG_SCAN_IN_BUFF, DATAO_REG_31__SCAN_IN_BUFF, ADDRESS_REG_16__SCAN_IN_BUFF, ADDRESS_REG_9__SCAN_IN_BUFF, ADDRESS_REG_12__SCAN_IN_BUFF, DATAO_REG_29__SCAN_IN_BUFF, DATAO_REG_0__SCAN_IN_BUFF, ADDRESS_REG_4__SCAN_IN_BUFF, D_C_N_REG_SCAN_IN_BUFF, DATAO_REG_4__SCAN_IN_BUFF, ADDRESS_REG_6__SCAN_IN_BUFF, DATAO_REG_2__SCAN_IN_BUFF, ADDRESS_REG_0__SCAN_IN_BUFF, DATAO_REG_18__SCAN_IN_BUFF, DATAO_REG_16__SCAN_IN_BUFF, ADDRESS_REG_24__SCAN_IN_BUFF, DATAO_REG_14__SCAN_IN_BUFF, W_R_N_REG_SCAN_IN_BUFF, ADDRESS_REG_15__SCAN_IN_BUFF, DATAO_REG_22__SCAN_IN_BUFF, U3445, U3446, U3447, U3448, U3213, U3212, U3211, U3210, U3209, U3208, U3207, U3206, U3205, U3204, U3203, U3202, U3201, U3200, U3199, U3198, U3197, U3196, U3195, U3194, U3193, U3192, U3191, U3190, U3189, U3188, U3187, U3186, U3185, U3184, U3183, U3182, U3181, U3451, U3452, U3180, U3179, U3178, U3177, U3176, U3175, U3174, U3173, U3172, U3171, U3170, U3169, U3168, U3167, U3166, U3165, U3164, U3163, U3162, U3161, U3160, U3159, U3158, U3157, U3156, U3155, U3154, U3153, U3152, U3151, U3453, U3150, U3149, U3148, U3147, U3146, U3145, U3144, U3143, U3142, U3141, U3140, U3139, U3138, U3137, U3136, U3135, U3134, U3133, U3132, U3131, U3130, U3129, U3128, U3127, U3126, U3125, U3124, U3123, U3122, U3121, U3120, U3119, U3118, U3117, U3116, U3115, U3114, U3113, U3112, U3111, U3110, U3109, U3108, U3107, U3106, U3105, U3104, U3103, U3102, U3101, U3100, U3099, U3098, U3097, U3096, U3095, U3094, U3093, U3092, U3091, U3090, U3089, U3088, U3087, U3086, U3085, U3084, U3083, U3082, U3081, U3080, U3079, U3078, U3077, U3076, U3075, U3074, U3073, U3072, U3071, U3070, U3069, U3068, U3067, U3066, U3065, U3064, U3063, U3062, U3061, U3060, U3059, U3058, U3057, U3056, U3055, U3054, U3053, U3052, U3051, U3050, U3049, U3048, U3047, U3046, U3045, U3044, U3043, U3042, U3041, U3040, U3039, U3038, U3037, U3036, U3035, U3034, U3033, U3032, U3031, U3030, U3029, U3028, U3027, U3026, U3025, U3024, U3023, U3022, U3021, U3020, U3455, U3456, U3459, U3460, U3461, U3019, U3462, U3463, U3464, U3465, U3018, U3017, U3016, U3015, U3014, U3013, U3012, U3011, U3010, U3009, U3008, U3007, U3006, U3005, U3004, U3003, U3002, U3001, U3000, U2999, U2998, U2997, U2996, U2995, U2994, U2993, U2992, U2991, U2990, U2989, U2988, U2987, U2986, U2985, U2984, U2983, U2982, U2981, U2980, U2979, U2978, U2977, U2976, U2975, U2974, U2973, U2972, U2971, U2970, U2969, U2968, U2967, U2966, U2965, U2964, U2963, U2962, U2961, U2960, U2959, U2958, U2957, U2956, U2955, U2954, U2953, U2952, U2951, U2950, U2949, U2948, U2947, U2946, U2945, U2944, U2943, U2942, U2941, U2940, U2939, U2938, U2937, U2936, U2935, U2934, U2933, U2932, U2931, U2930, U2929, U2928, U2927, U2926, U2925, U2924, U2923, U2922, U2921, U2920, U2919, U2918, U2917, U2916, U2915, U2914, U2913, U2912, U2911, U2910, U2909, U2908, U2907, U2906, U2905, U2904, U2903, U2902, U2901, U2900, U2899, U2898, U2897, U2896, U2895, U2894, U2893, U2892, U2891, U2890, U2889, U2888, U2887, U2886, U2885, U2884, U2883, U2882, U2881, U2880, U2879, U2878, U2877, U2876, U2875, U2874, U2873, U2872, U2871, U2870, U2869, U2868, U2867, U2866, U2865, U2864, U2863, U2862, U2861, U2860, U2859, U2858, U2857, U2856, U2855, U2854, U2853, U2852, U2851, U2850, U2849, U2848, U2847, U2846, U2845, U2844, U2843, U2842, U2841, U2840, U2839, U2838, U2837, U2836, U2835, U2834, U2833, U2832, U2831, U2830, U2829, U2828, U2827, U2826, U2825, U2824, U2823, U2822, U2821, U2820, U2819, U2818, U2817, U2816, U2815, U2814, U2813, U2812, U2811, U2810, U2809, U2808, U2807, U2806, U2805, U2804, U2803, U2802, U2801, U2800, U2799, U2798, U2797, U2796, U2795, U3468, U2794, U3469, U3470, U2793, U3471, U2792, U3472, U2791, U3473, U2790, U2789, U3474, U2788);
  Perturb perturb (INSTQUEUE_REG_12__2__SCAN_IN, INSTQUEUE_REG_2__5__SCAN_IN, INSTQUEUE_REG_1__0__SCAN_IN, INSTQUEUE_REG_0__4__SCAN_IN, INSTADDRPOINTER_REG_21__SCAN_IN, INSTQUEUE_REG_9__5__SCAN_IN, INSTQUEUE_REG_1__1__SCAN_IN, INSTQUEUE_REG_2__1__SCAN_IN, INSTQUEUE_REG_12__0__SCAN_IN, INSTADDRPOINTER_REG_20__SCAN_IN, INSTQUEUEWR_ADDR_REG_1__SCAN_IN, INSTQUEUE_REG_10__0__SCAN_IN, INSTADDRPOINTER_REG_11__SCAN_IN, INSTADDRPOINTER_REG_2__SCAN_IN, INSTQUEUERD_ADDR_REG_1__SCAN_IN, INSTADDRPOINTER_REG_4__SCAN_IN, INSTQUEUE_REG_14__5__SCAN_IN, INSTQUEUE_REG_0__7__SCAN_IN, INSTQUEUE_REG_6__6__SCAN_IN, INSTQUEUE_REG_9__3__SCAN_IN, INSTQUEUE_REG_2__7__SCAN_IN, INSTQUEUE_REG_1__3__SCAN_IN, INSTQUEUE_REG_3__7__SCAN_IN, INSTQUEUE_REG_5__0__SCAN_IN, STATE2_REG_2__SCAN_IN, INSTQUEUE_REG_11__3__SCAN_IN, INSTQUEUE_REG_6__2__SCAN_IN, EBX_REG_5__SCAN_IN, INSTQUEUE_REG_12__5__SCAN_IN, INSTQUEUE_REG_5__7__SCAN_IN, INSTQUEUE_REG_12__7__SCAN_IN, INSTQUEUEWR_ADDR_REG_2__SCAN_IN, perturb_signal);
  Restore restore (INSTQUEUE_REG_12__2__SCAN_IN, INSTQUEUE_REG_2__5__SCAN_IN, INSTQUEUE_REG_1__0__SCAN_IN, INSTQUEUE_REG_0__4__SCAN_IN, INSTADDRPOINTER_REG_21__SCAN_IN, INSTQUEUE_REG_9__5__SCAN_IN, INSTQUEUE_REG_1__1__SCAN_IN, INSTQUEUE_REG_2__1__SCAN_IN, INSTQUEUE_REG_12__0__SCAN_IN, INSTADDRPOINTER_REG_20__SCAN_IN, INSTQUEUEWR_ADDR_REG_1__SCAN_IN, INSTQUEUE_REG_10__0__SCAN_IN, INSTADDRPOINTER_REG_11__SCAN_IN, INSTADDRPOINTER_REG_2__SCAN_IN, INSTQUEUERD_ADDR_REG_1__SCAN_IN, INSTADDRPOINTER_REG_4__SCAN_IN, INSTQUEUE_REG_14__5__SCAN_IN, INSTQUEUE_REG_0__7__SCAN_IN, INSTQUEUE_REG_6__6__SCAN_IN, INSTQUEUE_REG_9__3__SCAN_IN, INSTQUEUE_REG_2__7__SCAN_IN, INSTQUEUE_REG_1__3__SCAN_IN, INSTQUEUE_REG_3__7__SCAN_IN, INSTQUEUE_REG_5__0__SCAN_IN, STATE2_REG_2__SCAN_IN, INSTQUEUE_REG_11__3__SCAN_IN, INSTQUEUE_REG_6__2__SCAN_IN, EBX_REG_5__SCAN_IN, INSTQUEUE_REG_12__5__SCAN_IN, INSTQUEUE_REG_5__7__SCAN_IN, INSTQUEUE_REG_12__7__SCAN_IN, INSTQUEUEWR_ADDR_REG_2__SCAN_IN, keyinput0, keyinput1, keyinput2, keyinput3, keyinput4, keyinput5, keyinput6, keyinput7, keyinput8, keyinput9, keyinput10, keyinput11, keyinput12, keyinput13, keyinput14, keyinput15, keyinput16, keyinput17, keyinput18, keyinput19, keyinput20, keyinput21, keyinput22, keyinput23, keyinput24, keyinput25, keyinput26, keyinput27, keyinput28, keyinput29, keyinput30, keyinput31, restore_signal);
endmodule
/*************** Top Level ***************/

// Main module
module b15_C_SFLL_HD_4_32_1(DATAO_REG_25__SCAN_IN, DATAO_REG_5__SCAN_IN, DATAO_REG_28__SCAN_IN, DATAO_REG_21__SCAN_IN, BE_N_REG_0__SCAN_IN, ADDRESS_REG_23__SCAN_IN, ADDRESS_REG_17__SCAN_IN, ADDRESS_REG_2__SCAN_IN, DATAO_REG_30__SCAN_IN, BE_N_REG_1__SCAN_IN, ADDRESS_REG_1__SCAN_IN, DATAO_REG_8__SCAN_IN, DATAO_REG_23__SCAN_IN, DATAO_REG_10__SCAN_IN, ADDRESS_REG_22__SCAN_IN, ADDRESS_REG_11__SCAN_IN, ADDRESS_REG_3__SCAN_IN, BE_N_REG_3__SCAN_IN, DATAO_REG_27__SCAN_IN, ADDRESS_REG_10__SCAN_IN, ADDRESS_REG_28__SCAN_IN, DATAO_REG_12__SCAN_IN, BE_N_REG_2__SCAN_IN, ADDRESS_REG_13__SCAN_IN, DATAO_REG_13__SCAN_IN, ADDRESS_REG_20__SCAN_IN, DATAO_REG_24__SCAN_IN, DATAO_REG_9__SCAN_IN, DATAO_REG_7__SCAN_IN, DATAO_REG_11__SCAN_IN, ADDRESS_REG_19__SCAN_IN, ADDRESS_REG_27__SCAN_IN, ADDRESS_REG_25__SCAN_IN, ADDRESS_REG_29__SCAN_IN, ADDRESS_REG_5__SCAN_IN, ADDRESS_REG_7__SCAN_IN, ADDRESS_REG_8__SCAN_IN, ADDRESS_REG_21__SCAN_IN, DATAO_REG_20__SCAN_IN, DATAO_REG_17__SCAN_IN, DATAO_REG_6__SCAN_IN, ADDRESS_REG_14__SCAN_IN, DATAO_REG_19__SCAN_IN, ADS_N_REG_SCAN_IN, DATAO_REG_15__SCAN_IN, DATAO_REG_26__SCAN_IN, DATAO_REG_3__SCAN_IN, DATAO_REG_1__SCAN_IN, ADDRESS_REG_26__SCAN_IN, ADDRESS_REG_18__SCAN_IN, M_IO_N_REG_SCAN_IN, DATAO_REG_31__SCAN_IN, ADDRESS_REG_16__SCAN_IN, ADDRESS_REG_9__SCAN_IN, ADDRESS_REG_12__SCAN_IN, DATAO_REG_29__SCAN_IN, DATAO_REG_0__SCAN_IN, ADDRESS_REG_4__SCAN_IN, D_C_N_REG_SCAN_IN, DATAO_REG_4__SCAN_IN, ADDRESS_REG_6__SCAN_IN, DATAO_REG_2__SCAN_IN, ADDRESS_REG_0__SCAN_IN, DATAO_REG_18__SCAN_IN, DATAO_REG_16__SCAN_IN, ADDRESS_REG_24__SCAN_IN, DATAO_REG_14__SCAN_IN, W_R_N_REG_SCAN_IN, ADDRESS_REG_15__SCAN_IN, DATAO_REG_22__SCAN_IN, DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, DATAI_27_, DATAI_26_, DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, DATAI_21_, DATAI_20_, DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, DATAI_15_, DATAI_14_, DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, DATAI_9_, DATAI_8_, DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, DATAI_2_, DATAI_1_, DATAI_0_, MEMORYFETCH_REG_SCAN_IN, NA_N, BS16_N, READY_N, HOLD, READREQUEST_REG_SCAN_IN, CODEFETCH_REG_SCAN_IN, REQUESTPENDING_REG_SCAN_IN, STATEBS16_REG_SCAN_IN, MORE_REG_SCAN_IN, FLUSH_REG_SCAN_IN, BYTEENABLE_REG_0__SCAN_IN, BYTEENABLE_REG_1__SCAN_IN, BYTEENABLE_REG_2__SCAN_IN, BYTEENABLE_REG_3__SCAN_IN, REIP_REG_31__SCAN_IN, REIP_REG_30__SCAN_IN, REIP_REG_29__SCAN_IN, REIP_REG_28__SCAN_IN, REIP_REG_27__SCAN_IN, REIP_REG_26__SCAN_IN, REIP_REG_25__SCAN_IN, REIP_REG_24__SCAN_IN, REIP_REG_23__SCAN_IN, REIP_REG_22__SCAN_IN, REIP_REG_21__SCAN_IN, REIP_REG_20__SCAN_IN, REIP_REG_19__SCAN_IN, REIP_REG_18__SCAN_IN, REIP_REG_17__SCAN_IN, REIP_REG_16__SCAN_IN, STATE_REG_2__SCAN_IN, STATE_REG_1__SCAN_IN, STATE_REG_0__SCAN_IN, DATAWIDTH_REG_0__SCAN_IN, DATAWIDTH_REG_1__SCAN_IN, DATAWIDTH_REG_2__SCAN_IN, DATAWIDTH_REG_3__SCAN_IN, DATAWIDTH_REG_4__SCAN_IN, DATAWIDTH_REG_5__SCAN_IN, DATAWIDTH_REG_6__SCAN_IN, DATAWIDTH_REG_7__SCAN_IN, DATAWIDTH_REG_8__SCAN_IN, DATAWIDTH_REG_9__SCAN_IN, DATAWIDTH_REG_10__SCAN_IN, DATAWIDTH_REG_11__SCAN_IN, DATAWIDTH_REG_12__SCAN_IN, DATAWIDTH_REG_13__SCAN_IN, DATAWIDTH_REG_14__SCAN_IN, DATAWIDTH_REG_15__SCAN_IN, DATAWIDTH_REG_16__SCAN_IN, DATAWIDTH_REG_17__SCAN_IN, DATAWIDTH_REG_18__SCAN_IN, DATAWIDTH_REG_19__SCAN_IN, DATAWIDTH_REG_20__SCAN_IN, DATAWIDTH_REG_21__SCAN_IN, DATAWIDTH_REG_22__SCAN_IN, DATAWIDTH_REG_23__SCAN_IN, DATAWIDTH_REG_24__SCAN_IN, DATAWIDTH_REG_25__SCAN_IN, DATAWIDTH_REG_26__SCAN_IN, DATAWIDTH_REG_27__SCAN_IN, DATAWIDTH_REG_28__SCAN_IN, DATAWIDTH_REG_29__SCAN_IN, DATAWIDTH_REG_30__SCAN_IN, DATAWIDTH_REG_31__SCAN_IN, STATE2_REG_3__SCAN_IN, STATE2_REG_2__SCAN_IN, STATE2_REG_1__SCAN_IN, STATE2_REG_0__SCAN_IN, INSTQUEUE_REG_15__7__SCAN_IN, INSTQUEUE_REG_15__6__SCAN_IN, INSTQUEUE_REG_15__5__SCAN_IN, INSTQUEUE_REG_15__4__SCAN_IN, INSTQUEUE_REG_15__3__SCAN_IN, INSTQUEUE_REG_15__2__SCAN_IN, INSTQUEUE_REG_15__1__SCAN_IN, INSTQUEUE_REG_15__0__SCAN_IN, INSTQUEUE_REG_14__7__SCAN_IN, INSTQUEUE_REG_14__6__SCAN_IN, INSTQUEUE_REG_14__5__SCAN_IN, INSTQUEUE_REG_14__4__SCAN_IN, INSTQUEUE_REG_14__3__SCAN_IN, INSTQUEUE_REG_14__2__SCAN_IN, INSTQUEUE_REG_14__1__SCAN_IN, INSTQUEUE_REG_14__0__SCAN_IN, INSTQUEUE_REG_13__7__SCAN_IN, INSTQUEUE_REG_13__6__SCAN_IN, INSTQUEUE_REG_13__5__SCAN_IN, INSTQUEUE_REG_13__4__SCAN_IN, INSTQUEUE_REG_13__3__SCAN_IN, INSTQUEUE_REG_13__2__SCAN_IN, INSTQUEUE_REG_13__1__SCAN_IN, INSTQUEUE_REG_13__0__SCAN_IN, INSTQUEUE_REG_12__7__SCAN_IN, INSTQUEUE_REG_12__6__SCAN_IN, INSTQUEUE_REG_12__5__SCAN_IN, INSTQUEUE_REG_12__4__SCAN_IN, INSTQUEUE_REG_12__3__SCAN_IN, INSTQUEUE_REG_12__2__SCAN_IN, INSTQUEUE_REG_12__1__SCAN_IN, INSTQUEUE_REG_12__0__SCAN_IN, INSTQUEUE_REG_11__7__SCAN_IN, INSTQUEUE_REG_11__6__SCAN_IN, INSTQUEUE_REG_11__5__SCAN_IN, INSTQUEUE_REG_11__4__SCAN_IN, INSTQUEUE_REG_11__3__SCAN_IN, INSTQUEUE_REG_11__2__SCAN_IN, INSTQUEUE_REG_11__1__SCAN_IN, INSTQUEUE_REG_11__0__SCAN_IN, INSTQUEUE_REG_10__7__SCAN_IN, INSTQUEUE_REG_10__6__SCAN_IN, INSTQUEUE_REG_10__5__SCAN_IN, INSTQUEUE_REG_10__4__SCAN_IN, INSTQUEUE_REG_10__3__SCAN_IN, INSTQUEUE_REG_10__2__SCAN_IN, INSTQUEUE_REG_10__1__SCAN_IN, INSTQUEUE_REG_10__0__SCAN_IN, INSTQUEUE_REG_9__7__SCAN_IN, INSTQUEUE_REG_9__6__SCAN_IN, INSTQUEUE_REG_9__5__SCAN_IN, INSTQUEUE_REG_9__4__SCAN_IN, INSTQUEUE_REG_9__3__SCAN_IN, INSTQUEUE_REG_9__2__SCAN_IN, INSTQUEUE_REG_9__1__SCAN_IN, INSTQUEUE_REG_9__0__SCAN_IN, INSTQUEUE_REG_8__7__SCAN_IN, INSTQUEUE_REG_8__6__SCAN_IN, INSTQUEUE_REG_8__5__SCAN_IN, INSTQUEUE_REG_8__4__SCAN_IN, INSTQUEUE_REG_8__3__SCAN_IN, INSTQUEUE_REG_8__2__SCAN_IN, INSTQUEUE_REG_8__1__SCAN_IN, INSTQUEUE_REG_8__0__SCAN_IN, INSTQUEUE_REG_7__7__SCAN_IN, INSTQUEUE_REG_7__6__SCAN_IN, INSTQUEUE_REG_7__5__SCAN_IN, INSTQUEUE_REG_7__4__SCAN_IN, INSTQUEUE_REG_7__3__SCAN_IN, INSTQUEUE_REG_7__2__SCAN_IN, INSTQUEUE_REG_7__1__SCAN_IN, INSTQUEUE_REG_7__0__SCAN_IN, INSTQUEUE_REG_6__7__SCAN_IN, INSTQUEUE_REG_6__6__SCAN_IN, INSTQUEUE_REG_6__5__SCAN_IN, INSTQUEUE_REG_6__4__SCAN_IN, INSTQUEUE_REG_6__3__SCAN_IN, INSTQUEUE_REG_6__2__SCAN_IN, INSTQUEUE_REG_6__1__SCAN_IN, INSTQUEUE_REG_6__0__SCAN_IN, INSTQUEUE_REG_5__7__SCAN_IN, INSTQUEUE_REG_5__6__SCAN_IN, INSTQUEUE_REG_5__5__SCAN_IN, INSTQUEUE_REG_5__4__SCAN_IN, INSTQUEUE_REG_5__3__SCAN_IN, INSTQUEUE_REG_5__2__SCAN_IN, INSTQUEUE_REG_5__1__SCAN_IN, INSTQUEUE_REG_5__0__SCAN_IN, INSTQUEUE_REG_4__7__SCAN_IN, INSTQUEUE_REG_4__6__SCAN_IN, INSTQUEUE_REG_4__5__SCAN_IN, INSTQUEUE_REG_4__4__SCAN_IN, INSTQUEUE_REG_4__3__SCAN_IN, INSTQUEUE_REG_4__2__SCAN_IN, INSTQUEUE_REG_4__1__SCAN_IN, INSTQUEUE_REG_4__0__SCAN_IN, INSTQUEUE_REG_3__7__SCAN_IN, INSTQUEUE_REG_3__6__SCAN_IN, INSTQUEUE_REG_3__5__SCAN_IN, INSTQUEUE_REG_3__4__SCAN_IN, INSTQUEUE_REG_3__3__SCAN_IN, INSTQUEUE_REG_3__2__SCAN_IN, INSTQUEUE_REG_3__1__SCAN_IN, INSTQUEUE_REG_3__0__SCAN_IN, INSTQUEUE_REG_2__7__SCAN_IN, INSTQUEUE_REG_2__6__SCAN_IN, INSTQUEUE_REG_2__5__SCAN_IN, INSTQUEUE_REG_2__4__SCAN_IN, INSTQUEUE_REG_2__3__SCAN_IN, INSTQUEUE_REG_2__2__SCAN_IN, INSTQUEUE_REG_2__1__SCAN_IN, INSTQUEUE_REG_2__0__SCAN_IN, INSTQUEUE_REG_1__7__SCAN_IN, INSTQUEUE_REG_1__6__SCAN_IN, INSTQUEUE_REG_1__5__SCAN_IN, INSTQUEUE_REG_1__4__SCAN_IN, INSTQUEUE_REG_1__3__SCAN_IN, INSTQUEUE_REG_1__2__SCAN_IN, INSTQUEUE_REG_1__1__SCAN_IN, INSTQUEUE_REG_1__0__SCAN_IN, INSTQUEUE_REG_0__7__SCAN_IN, INSTQUEUE_REG_0__6__SCAN_IN, INSTQUEUE_REG_0__5__SCAN_IN, INSTQUEUE_REG_0__4__SCAN_IN, INSTQUEUE_REG_0__3__SCAN_IN, INSTQUEUE_REG_0__2__SCAN_IN, INSTQUEUE_REG_0__1__SCAN_IN, INSTQUEUE_REG_0__0__SCAN_IN, INSTQUEUERD_ADDR_REG_4__SCAN_IN, INSTQUEUERD_ADDR_REG_3__SCAN_IN, INSTQUEUERD_ADDR_REG_2__SCAN_IN, INSTQUEUERD_ADDR_REG_1__SCAN_IN, INSTQUEUERD_ADDR_REG_0__SCAN_IN, INSTQUEUEWR_ADDR_REG_4__SCAN_IN, INSTQUEUEWR_ADDR_REG_3__SCAN_IN, INSTQUEUEWR_ADDR_REG_2__SCAN_IN, INSTQUEUEWR_ADDR_REG_1__SCAN_IN, INSTQUEUEWR_ADDR_REG_0__SCAN_IN, INSTADDRPOINTER_REG_0__SCAN_IN, INSTADDRPOINTER_REG_1__SCAN_IN, INSTADDRPOINTER_REG_2__SCAN_IN, INSTADDRPOINTER_REG_3__SCAN_IN, INSTADDRPOINTER_REG_4__SCAN_IN, INSTADDRPOINTER_REG_5__SCAN_IN, INSTADDRPOINTER_REG_6__SCAN_IN, INSTADDRPOINTER_REG_7__SCAN_IN, INSTADDRPOINTER_REG_8__SCAN_IN, INSTADDRPOINTER_REG_9__SCAN_IN, INSTADDRPOINTER_REG_10__SCAN_IN, INSTADDRPOINTER_REG_11__SCAN_IN, INSTADDRPOINTER_REG_12__SCAN_IN, INSTADDRPOINTER_REG_13__SCAN_IN, INSTADDRPOINTER_REG_14__SCAN_IN, INSTADDRPOINTER_REG_15__SCAN_IN, INSTADDRPOINTER_REG_16__SCAN_IN, INSTADDRPOINTER_REG_17__SCAN_IN, INSTADDRPOINTER_REG_18__SCAN_IN, INSTADDRPOINTER_REG_19__SCAN_IN, INSTADDRPOINTER_REG_20__SCAN_IN, INSTADDRPOINTER_REG_21__SCAN_IN, INSTADDRPOINTER_REG_22__SCAN_IN, INSTADDRPOINTER_REG_23__SCAN_IN, INSTADDRPOINTER_REG_24__SCAN_IN, INSTADDRPOINTER_REG_25__SCAN_IN, INSTADDRPOINTER_REG_26__SCAN_IN, INSTADDRPOINTER_REG_27__SCAN_IN, INSTADDRPOINTER_REG_28__SCAN_IN, INSTADDRPOINTER_REG_29__SCAN_IN, INSTADDRPOINTER_REG_30__SCAN_IN, INSTADDRPOINTER_REG_31__SCAN_IN, PHYADDRPOINTER_REG_0__SCAN_IN, PHYADDRPOINTER_REG_1__SCAN_IN, PHYADDRPOINTER_REG_2__SCAN_IN, PHYADDRPOINTER_REG_3__SCAN_IN, PHYADDRPOINTER_REG_4__SCAN_IN, PHYADDRPOINTER_REG_5__SCAN_IN, PHYADDRPOINTER_REG_6__SCAN_IN, PHYADDRPOINTER_REG_7__SCAN_IN, PHYADDRPOINTER_REG_8__SCAN_IN, PHYADDRPOINTER_REG_9__SCAN_IN, PHYADDRPOINTER_REG_10__SCAN_IN, PHYADDRPOINTER_REG_11__SCAN_IN, PHYADDRPOINTER_REG_12__SCAN_IN, PHYADDRPOINTER_REG_13__SCAN_IN, PHYADDRPOINTER_REG_14__SCAN_IN, PHYADDRPOINTER_REG_15__SCAN_IN, PHYADDRPOINTER_REG_16__SCAN_IN, PHYADDRPOINTER_REG_17__SCAN_IN, PHYADDRPOINTER_REG_18__SCAN_IN, PHYADDRPOINTER_REG_19__SCAN_IN, PHYADDRPOINTER_REG_20__SCAN_IN, PHYADDRPOINTER_REG_21__SCAN_IN, PHYADDRPOINTER_REG_22__SCAN_IN, PHYADDRPOINTER_REG_23__SCAN_IN, PHYADDRPOINTER_REG_24__SCAN_IN, PHYADDRPOINTER_REG_25__SCAN_IN, PHYADDRPOINTER_REG_26__SCAN_IN, PHYADDRPOINTER_REG_27__SCAN_IN, PHYADDRPOINTER_REG_28__SCAN_IN, PHYADDRPOINTER_REG_29__SCAN_IN, PHYADDRPOINTER_REG_30__SCAN_IN, PHYADDRPOINTER_REG_31__SCAN_IN, LWORD_REG_15__SCAN_IN, LWORD_REG_14__SCAN_IN, LWORD_REG_13__SCAN_IN, LWORD_REG_12__SCAN_IN, LWORD_REG_11__SCAN_IN, LWORD_REG_10__SCAN_IN, LWORD_REG_9__SCAN_IN, LWORD_REG_8__SCAN_IN, LWORD_REG_7__SCAN_IN, LWORD_REG_6__SCAN_IN, LWORD_REG_5__SCAN_IN, LWORD_REG_4__SCAN_IN, LWORD_REG_3__SCAN_IN, LWORD_REG_2__SCAN_IN, LWORD_REG_1__SCAN_IN, LWORD_REG_0__SCAN_IN, UWORD_REG_14__SCAN_IN, UWORD_REG_13__SCAN_IN, UWORD_REG_12__SCAN_IN, UWORD_REG_11__SCAN_IN, UWORD_REG_10__SCAN_IN, UWORD_REG_9__SCAN_IN, UWORD_REG_8__SCAN_IN, UWORD_REG_7__SCAN_IN, UWORD_REG_6__SCAN_IN, UWORD_REG_5__SCAN_IN, UWORD_REG_4__SCAN_IN, UWORD_REG_3__SCAN_IN, UWORD_REG_2__SCAN_IN, UWORD_REG_1__SCAN_IN, UWORD_REG_0__SCAN_IN, EAX_REG_0__SCAN_IN, EAX_REG_1__SCAN_IN, EAX_REG_2__SCAN_IN, EAX_REG_3__SCAN_IN, EAX_REG_4__SCAN_IN, EAX_REG_5__SCAN_IN, EAX_REG_6__SCAN_IN, EAX_REG_7__SCAN_IN, EAX_REG_8__SCAN_IN, EAX_REG_9__SCAN_IN, EAX_REG_10__SCAN_IN, EAX_REG_11__SCAN_IN, EAX_REG_12__SCAN_IN, EAX_REG_13__SCAN_IN, EAX_REG_14__SCAN_IN, EAX_REG_15__SCAN_IN, EAX_REG_16__SCAN_IN, EAX_REG_17__SCAN_IN, EAX_REG_18__SCAN_IN, EAX_REG_19__SCAN_IN, EAX_REG_20__SCAN_IN, EAX_REG_21__SCAN_IN, EAX_REG_22__SCAN_IN, EAX_REG_23__SCAN_IN, EAX_REG_24__SCAN_IN, EAX_REG_25__SCAN_IN, EAX_REG_26__SCAN_IN, EAX_REG_27__SCAN_IN, EAX_REG_28__SCAN_IN, EAX_REG_29__SCAN_IN, EAX_REG_30__SCAN_IN, EAX_REG_31__SCAN_IN, EBX_REG_0__SCAN_IN, EBX_REG_1__SCAN_IN, EBX_REG_2__SCAN_IN, EBX_REG_3__SCAN_IN, EBX_REG_4__SCAN_IN, EBX_REG_5__SCAN_IN, EBX_REG_6__SCAN_IN, EBX_REG_7__SCAN_IN, EBX_REG_8__SCAN_IN, EBX_REG_9__SCAN_IN, EBX_REG_10__SCAN_IN, EBX_REG_11__SCAN_IN, EBX_REG_12__SCAN_IN, EBX_REG_13__SCAN_IN, EBX_REG_14__SCAN_IN, EBX_REG_15__SCAN_IN, EBX_REG_16__SCAN_IN, EBX_REG_17__SCAN_IN, EBX_REG_18__SCAN_IN, EBX_REG_19__SCAN_IN, EBX_REG_20__SCAN_IN, EBX_REG_21__SCAN_IN, EBX_REG_22__SCAN_IN, EBX_REG_23__SCAN_IN, EBX_REG_24__SCAN_IN, EBX_REG_25__SCAN_IN, EBX_REG_26__SCAN_IN, EBX_REG_27__SCAN_IN, EBX_REG_28__SCAN_IN, EBX_REG_29__SCAN_IN, EBX_REG_30__SCAN_IN, EBX_REG_31__SCAN_IN, REIP_REG_0__SCAN_IN, REIP_REG_1__SCAN_IN, REIP_REG_2__SCAN_IN, REIP_REG_3__SCAN_IN, REIP_REG_4__SCAN_IN, REIP_REG_5__SCAN_IN, REIP_REG_6__SCAN_IN, REIP_REG_7__SCAN_IN, REIP_REG_8__SCAN_IN, REIP_REG_9__SCAN_IN, REIP_REG_10__SCAN_IN, REIP_REG_11__SCAN_IN, REIP_REG_12__SCAN_IN, REIP_REG_13__SCAN_IN, REIP_REG_14__SCAN_IN, REIP_REG_15__SCAN_IN, perturb_signal, restore_signal, DATAO_REG_25__SCAN_IN_BUFF, DATAO_REG_5__SCAN_IN_BUFF, DATAO_REG_28__SCAN_IN_BUFF, DATAO_REG_21__SCAN_IN_BUFF, BE_N_REG_0__SCAN_IN_BUFF, ADDRESS_REG_23__SCAN_IN_BUFF, ADDRESS_REG_17__SCAN_IN_BUFF, ADDRESS_REG_2__SCAN_IN_BUFF, DATAO_REG_30__SCAN_IN_BUFF, BE_N_REG_1__SCAN_IN_BUFF, ADDRESS_REG_1__SCAN_IN_BUFF, DATAO_REG_8__SCAN_IN_BUFF, DATAO_REG_23__SCAN_IN_BUFF, DATAO_REG_10__SCAN_IN_BUFF, ADDRESS_REG_22__SCAN_IN_BUFF, ADDRESS_REG_11__SCAN_IN_BUFF, ADDRESS_REG_3__SCAN_IN_BUFF, BE_N_REG_3__SCAN_IN_BUFF, DATAO_REG_27__SCAN_IN_BUFF, ADDRESS_REG_10__SCAN_IN_BUFF, ADDRESS_REG_28__SCAN_IN_BUFF, DATAO_REG_12__SCAN_IN_BUFF, BE_N_REG_2__SCAN_IN_BUFF, ADDRESS_REG_13__SCAN_IN_BUFF, DATAO_REG_13__SCAN_IN_BUFF, ADDRESS_REG_20__SCAN_IN_BUFF, DATAO_REG_24__SCAN_IN_BUFF, DATAO_REG_9__SCAN_IN_BUFF, DATAO_REG_7__SCAN_IN_BUFF, DATAO_REG_11__SCAN_IN_BUFF, ADDRESS_REG_19__SCAN_IN_BUFF, ADDRESS_REG_27__SCAN_IN_BUFF, ADDRESS_REG_25__SCAN_IN_BUFF, ADDRESS_REG_29__SCAN_IN_BUFF, ADDRESS_REG_5__SCAN_IN_BUFF, ADDRESS_REG_7__SCAN_IN_BUFF, ADDRESS_REG_8__SCAN_IN_BUFF, ADDRESS_REG_21__SCAN_IN_BUFF, DATAO_REG_20__SCAN_IN_BUFF, DATAO_REG_17__SCAN_IN_BUFF, DATAO_REG_6__SCAN_IN_BUFF, ADDRESS_REG_14__SCAN_IN_BUFF, DATAO_REG_19__SCAN_IN_BUFF, ADS_N_REG_SCAN_IN_BUFF, DATAO_REG_15__SCAN_IN_BUFF, DATAO_REG_26__SCAN_IN_BUFF, DATAO_REG_3__SCAN_IN_BUFF, DATAO_REG_1__SCAN_IN_BUFF, ADDRESS_REG_26__SCAN_IN_BUFF, ADDRESS_REG_18__SCAN_IN_BUFF, M_IO_N_REG_SCAN_IN_BUFF, DATAO_REG_31__SCAN_IN_BUFF, ADDRESS_REG_16__SCAN_IN_BUFF, ADDRESS_REG_9__SCAN_IN_BUFF, ADDRESS_REG_12__SCAN_IN_BUFF, DATAO_REG_29__SCAN_IN_BUFF, DATAO_REG_0__SCAN_IN_BUFF, ADDRESS_REG_4__SCAN_IN_BUFF, D_C_N_REG_SCAN_IN_BUFF, DATAO_REG_4__SCAN_IN_BUFF, ADDRESS_REG_6__SCAN_IN_BUFF, DATAO_REG_2__SCAN_IN_BUFF, ADDRESS_REG_0__SCAN_IN_BUFF, DATAO_REG_18__SCAN_IN_BUFF, DATAO_REG_16__SCAN_IN_BUFF, ADDRESS_REG_24__SCAN_IN_BUFF, DATAO_REG_14__SCAN_IN_BUFF, W_R_N_REG_SCAN_IN_BUFF, ADDRESS_REG_15__SCAN_IN_BUFF, DATAO_REG_22__SCAN_IN_BUFF, U3445, U3446, U3447, U3448, U3213, U3212, U3211, U3210, U3209, U3208, U3207, U3206, U3205, U3204, U3203, U3202, U3201, U3200, U3199, U3198, U3197, U3196, U3195, U3194, U3193, U3192, U3191, U3190, U3189, U3188, U3187, U3186, U3185, U3184, U3183, U3182, U3181, U3451, U3452, U3180, U3179, U3178, U3177, U3176, U3175, U3174, U3173, U3172, U3171, U3170, U3169, U3168, U3167, U3166, U3165, U3164, U3163, U3162, U3161, U3160, U3159, U3158, U3157, U3156, U3155, U3154, U3153, U3152, U3151, U3453, U3150, U3149, U3148, U3147, U3146, U3145, U3144, U3143, U3142, U3141, U3140, U3139, U3138, U3137, U3136, U3135, U3134, U3133, U3132, U3131, U3130, U3129, U3128, U3127, U3126, U3125, U3124, U3123, U3122, U3121, U3120, U3119, U3118, U3117, U3116, U3115, U3114, U3113, U3112, U3111, U3110, U3109, U3108, U3107, U3106, U3105, U3104, U3103, U3102, U3101, U3100, U3099, U3098, U3097, U3096, U3095, U3094, U3093, U3092, U3091, U3090, U3089, U3088, U3087, U3086, U3085, U3084, U3083, U3082, U3081, U3080, U3079, U3078, U3077, U3076, U3075, U3074, U3073, U3072, U3071, U3070, U3069, U3068, U3067, U3066, U3065, U3064, U3063, U3062, U3061, U3060, U3059, U3058, U3057, U3056, U3055, U3054, U3053, U3052, U3051, U3050, U3049, U3048, U3047, U3046, U3045, U3044, U3043, U3042, U3041, U3040, U3039, U3038, U3037, U3036, U3035, U3034, U3033, U3032, U3031, U3030, U3029, U3028, U3027, U3026, U3025, U3024, U3023, U3022, U3021, U3020, U3455, U3456, U3459, U3460, U3461, U3019, U3462, U3463, U3464, U3465, U3018, U3017, U3016, U3015, U3014, U3013, U3012, U3011, U3010, U3009, U3008, U3007, U3006, U3005, U3004, U3003, U3002, U3001, U3000, U2999, U2998, U2997, U2996, U2995, U2994, U2993, U2992, U2991, U2990, U2989, U2988, U2987, U2986, U2985, U2984, U2983, U2982, U2981, U2980, U2979, U2978, U2977, U2976, U2975, U2974, U2973, U2972, U2971, U2970, U2969, U2968, U2967, U2966, U2965, U2964, U2963, U2962, U2961, U2960, U2959, U2958, U2957, U2956, U2955, U2954, U2953, U2952, U2951, U2950, U2949, U2948, U2947, U2946, U2945, U2944, U2943, U2942, U2941, U2940, U2939, U2938, U2937, U2936, U2935, U2934, U2933, U2932, U2931, U2930, U2929, U2928, U2927, U2926, U2925, U2924, U2923, U2922, U2921, U2920, U2919, U2918, U2917, U2916, U2915, U2914, U2913, U2912, U2911, U2910, U2909, U2908, U2907, U2906, U2905, U2904, U2903, U2902, U2901, U2900, U2899, U2898, U2897, U2896, U2895, U2894, U2893, U2892, U2891, U2890, U2889, U2888, U2887, U2886, U2885, U2884, U2883, U2882, U2881, U2880, U2879, U2878, U2877, U2876, U2875, U2874, U2873, U2872, U2871, U2870, U2869, U2868, U2867, U2866, U2865, U2864, U2863, U2862, U2861, U2860, U2859, U2858, U2857, U2856, U2855, U2854, U2853, U2852, U2851, U2850, U2849, U2848, U2847, U2846, U2845, U2844, U2843, U2842, U2841, U2840, U2839, U2838, U2837, U2836, U2835, U2834, U2833, U2832, U2831, U2830, U2829, U2828, U2827, U2826, U2825, U2824, U2823, U2822, U2821, U2820, U2819, U2818, U2817, U2816, U2815, U2814, U2813, U2812, U2811, U2810, U2809, U2808, U2807, U2806, U2805, U2804, U2803, U2802, U2801, U2800, U2799, U2798, U2797, U2796, U2795, U3468, U2794, U3469, U3470, U2793, U3471, U2792, U3472, U2791, U3473, U2790, U2789, U3474, U2788);

  input DATAO_REG_25__SCAN_IN, DATAO_REG_5__SCAN_IN, DATAO_REG_28__SCAN_IN, DATAO_REG_21__SCAN_IN, BE_N_REG_0__SCAN_IN, ADDRESS_REG_23__SCAN_IN, ADDRESS_REG_17__SCAN_IN, ADDRESS_REG_2__SCAN_IN, DATAO_REG_30__SCAN_IN, BE_N_REG_1__SCAN_IN, ADDRESS_REG_1__SCAN_IN, DATAO_REG_8__SCAN_IN, DATAO_REG_23__SCAN_IN, DATAO_REG_10__SCAN_IN, ADDRESS_REG_22__SCAN_IN, ADDRESS_REG_11__SCAN_IN, ADDRESS_REG_3__SCAN_IN, BE_N_REG_3__SCAN_IN, DATAO_REG_27__SCAN_IN, ADDRESS_REG_10__SCAN_IN, ADDRESS_REG_28__SCAN_IN, DATAO_REG_12__SCAN_IN, BE_N_REG_2__SCAN_IN, ADDRESS_REG_13__SCAN_IN, DATAO_REG_13__SCAN_IN, ADDRESS_REG_20__SCAN_IN, DATAO_REG_24__SCAN_IN, DATAO_REG_9__SCAN_IN, DATAO_REG_7__SCAN_IN, DATAO_REG_11__SCAN_IN, ADDRESS_REG_19__SCAN_IN, ADDRESS_REG_27__SCAN_IN, ADDRESS_REG_25__SCAN_IN, ADDRESS_REG_29__SCAN_IN, ADDRESS_REG_5__SCAN_IN, ADDRESS_REG_7__SCAN_IN, ADDRESS_REG_8__SCAN_IN, ADDRESS_REG_21__SCAN_IN, DATAO_REG_20__SCAN_IN, DATAO_REG_17__SCAN_IN, DATAO_REG_6__SCAN_IN, ADDRESS_REG_14__SCAN_IN, DATAO_REG_19__SCAN_IN, ADS_N_REG_SCAN_IN, DATAO_REG_15__SCAN_IN, DATAO_REG_26__SCAN_IN, DATAO_REG_3__SCAN_IN, DATAO_REG_1__SCAN_IN, ADDRESS_REG_26__SCAN_IN, ADDRESS_REG_18__SCAN_IN, M_IO_N_REG_SCAN_IN, DATAO_REG_31__SCAN_IN, ADDRESS_REG_16__SCAN_IN, ADDRESS_REG_9__SCAN_IN, ADDRESS_REG_12__SCAN_IN, DATAO_REG_29__SCAN_IN, DATAO_REG_0__SCAN_IN, ADDRESS_REG_4__SCAN_IN, D_C_N_REG_SCAN_IN, DATAO_REG_4__SCAN_IN, ADDRESS_REG_6__SCAN_IN, DATAO_REG_2__SCAN_IN, ADDRESS_REG_0__SCAN_IN, DATAO_REG_18__SCAN_IN, DATAO_REG_16__SCAN_IN, ADDRESS_REG_24__SCAN_IN, DATAO_REG_14__SCAN_IN, W_R_N_REG_SCAN_IN, ADDRESS_REG_15__SCAN_IN, DATAO_REG_22__SCAN_IN, DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, DATAI_27_, DATAI_26_, DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, DATAI_21_, DATAI_20_, DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, DATAI_15_, DATAI_14_, DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, DATAI_9_, DATAI_8_, DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, DATAI_2_, DATAI_1_, DATAI_0_, MEMORYFETCH_REG_SCAN_IN, NA_N, BS16_N, READY_N, HOLD, READREQUEST_REG_SCAN_IN, CODEFETCH_REG_SCAN_IN, REQUESTPENDING_REG_SCAN_IN, STATEBS16_REG_SCAN_IN, MORE_REG_SCAN_IN, FLUSH_REG_SCAN_IN, BYTEENABLE_REG_0__SCAN_IN, BYTEENABLE_REG_1__SCAN_IN, BYTEENABLE_REG_2__SCAN_IN, BYTEENABLE_REG_3__SCAN_IN, REIP_REG_31__SCAN_IN, REIP_REG_30__SCAN_IN, REIP_REG_29__SCAN_IN, REIP_REG_28__SCAN_IN, REIP_REG_27__SCAN_IN, REIP_REG_26__SCAN_IN, REIP_REG_25__SCAN_IN, REIP_REG_24__SCAN_IN, REIP_REG_23__SCAN_IN, REIP_REG_22__SCAN_IN, REIP_REG_21__SCAN_IN, REIP_REG_20__SCAN_IN, REIP_REG_19__SCAN_IN, REIP_REG_18__SCAN_IN, REIP_REG_17__SCAN_IN, REIP_REG_16__SCAN_IN, STATE_REG_2__SCAN_IN, STATE_REG_1__SCAN_IN, STATE_REG_0__SCAN_IN, DATAWIDTH_REG_0__SCAN_IN, DATAWIDTH_REG_1__SCAN_IN, DATAWIDTH_REG_2__SCAN_IN, DATAWIDTH_REG_3__SCAN_IN, DATAWIDTH_REG_4__SCAN_IN, DATAWIDTH_REG_5__SCAN_IN, DATAWIDTH_REG_6__SCAN_IN, DATAWIDTH_REG_7__SCAN_IN, DATAWIDTH_REG_8__SCAN_IN, DATAWIDTH_REG_9__SCAN_IN, DATAWIDTH_REG_10__SCAN_IN, DATAWIDTH_REG_11__SCAN_IN, DATAWIDTH_REG_12__SCAN_IN, DATAWIDTH_REG_13__SCAN_IN, DATAWIDTH_REG_14__SCAN_IN, DATAWIDTH_REG_15__SCAN_IN, DATAWIDTH_REG_16__SCAN_IN, DATAWIDTH_REG_17__SCAN_IN, DATAWIDTH_REG_18__SCAN_IN, DATAWIDTH_REG_19__SCAN_IN, DATAWIDTH_REG_20__SCAN_IN, DATAWIDTH_REG_21__SCAN_IN, DATAWIDTH_REG_22__SCAN_IN, DATAWIDTH_REG_23__SCAN_IN, DATAWIDTH_REG_24__SCAN_IN, DATAWIDTH_REG_25__SCAN_IN, DATAWIDTH_REG_26__SCAN_IN, DATAWIDTH_REG_27__SCAN_IN, DATAWIDTH_REG_28__SCAN_IN, DATAWIDTH_REG_29__SCAN_IN, DATAWIDTH_REG_30__SCAN_IN, DATAWIDTH_REG_31__SCAN_IN, STATE2_REG_3__SCAN_IN, STATE2_REG_2__SCAN_IN, STATE2_REG_1__SCAN_IN, STATE2_REG_0__SCAN_IN, INSTQUEUE_REG_15__7__SCAN_IN, INSTQUEUE_REG_15__6__SCAN_IN, INSTQUEUE_REG_15__5__SCAN_IN, INSTQUEUE_REG_15__4__SCAN_IN, INSTQUEUE_REG_15__3__SCAN_IN, INSTQUEUE_REG_15__2__SCAN_IN, INSTQUEUE_REG_15__1__SCAN_IN, INSTQUEUE_REG_15__0__SCAN_IN, INSTQUEUE_REG_14__7__SCAN_IN, INSTQUEUE_REG_14__6__SCAN_IN, INSTQUEUE_REG_14__5__SCAN_IN, INSTQUEUE_REG_14__4__SCAN_IN, INSTQUEUE_REG_14__3__SCAN_IN, INSTQUEUE_REG_14__2__SCAN_IN, INSTQUEUE_REG_14__1__SCAN_IN, INSTQUEUE_REG_14__0__SCAN_IN, INSTQUEUE_REG_13__7__SCAN_IN, INSTQUEUE_REG_13__6__SCAN_IN, INSTQUEUE_REG_13__5__SCAN_IN, INSTQUEUE_REG_13__4__SCAN_IN, INSTQUEUE_REG_13__3__SCAN_IN, INSTQUEUE_REG_13__2__SCAN_IN, INSTQUEUE_REG_13__1__SCAN_IN, INSTQUEUE_REG_13__0__SCAN_IN, INSTQUEUE_REG_12__7__SCAN_IN, INSTQUEUE_REG_12__6__SCAN_IN, INSTQUEUE_REG_12__5__SCAN_IN, INSTQUEUE_REG_12__4__SCAN_IN, INSTQUEUE_REG_12__3__SCAN_IN, INSTQUEUE_REG_12__2__SCAN_IN, INSTQUEUE_REG_12__1__SCAN_IN, INSTQUEUE_REG_12__0__SCAN_IN, INSTQUEUE_REG_11__7__SCAN_IN, INSTQUEUE_REG_11__6__SCAN_IN, INSTQUEUE_REG_11__5__SCAN_IN, INSTQUEUE_REG_11__4__SCAN_IN, INSTQUEUE_REG_11__3__SCAN_IN, INSTQUEUE_REG_11__2__SCAN_IN, INSTQUEUE_REG_11__1__SCAN_IN, INSTQUEUE_REG_11__0__SCAN_IN, INSTQUEUE_REG_10__7__SCAN_IN, INSTQUEUE_REG_10__6__SCAN_IN, INSTQUEUE_REG_10__5__SCAN_IN, INSTQUEUE_REG_10__4__SCAN_IN, INSTQUEUE_REG_10__3__SCAN_IN, INSTQUEUE_REG_10__2__SCAN_IN, INSTQUEUE_REG_10__1__SCAN_IN, INSTQUEUE_REG_10__0__SCAN_IN, INSTQUEUE_REG_9__7__SCAN_IN, INSTQUEUE_REG_9__6__SCAN_IN, INSTQUEUE_REG_9__5__SCAN_IN, INSTQUEUE_REG_9__4__SCAN_IN, INSTQUEUE_REG_9__3__SCAN_IN, INSTQUEUE_REG_9__2__SCAN_IN, INSTQUEUE_REG_9__1__SCAN_IN, INSTQUEUE_REG_9__0__SCAN_IN, INSTQUEUE_REG_8__7__SCAN_IN, INSTQUEUE_REG_8__6__SCAN_IN, INSTQUEUE_REG_8__5__SCAN_IN, INSTQUEUE_REG_8__4__SCAN_IN, INSTQUEUE_REG_8__3__SCAN_IN, INSTQUEUE_REG_8__2__SCAN_IN, INSTQUEUE_REG_8__1__SCAN_IN, INSTQUEUE_REG_8__0__SCAN_IN, INSTQUEUE_REG_7__7__SCAN_IN, INSTQUEUE_REG_7__6__SCAN_IN, INSTQUEUE_REG_7__5__SCAN_IN, INSTQUEUE_REG_7__4__SCAN_IN, INSTQUEUE_REG_7__3__SCAN_IN, INSTQUEUE_REG_7__2__SCAN_IN, INSTQUEUE_REG_7__1__SCAN_IN, INSTQUEUE_REG_7__0__SCAN_IN, INSTQUEUE_REG_6__7__SCAN_IN, INSTQUEUE_REG_6__6__SCAN_IN, INSTQUEUE_REG_6__5__SCAN_IN, INSTQUEUE_REG_6__4__SCAN_IN, INSTQUEUE_REG_6__3__SCAN_IN, INSTQUEUE_REG_6__2__SCAN_IN, INSTQUEUE_REG_6__1__SCAN_IN, INSTQUEUE_REG_6__0__SCAN_IN, INSTQUEUE_REG_5__7__SCAN_IN, INSTQUEUE_REG_5__6__SCAN_IN, INSTQUEUE_REG_5__5__SCAN_IN, INSTQUEUE_REG_5__4__SCAN_IN, INSTQUEUE_REG_5__3__SCAN_IN, INSTQUEUE_REG_5__2__SCAN_IN, INSTQUEUE_REG_5__1__SCAN_IN, INSTQUEUE_REG_5__0__SCAN_IN, INSTQUEUE_REG_4__7__SCAN_IN, INSTQUEUE_REG_4__6__SCAN_IN, INSTQUEUE_REG_4__5__SCAN_IN, INSTQUEUE_REG_4__4__SCAN_IN, INSTQUEUE_REG_4__3__SCAN_IN, INSTQUEUE_REG_4__2__SCAN_IN, INSTQUEUE_REG_4__1__SCAN_IN, INSTQUEUE_REG_4__0__SCAN_IN, INSTQUEUE_REG_3__7__SCAN_IN, INSTQUEUE_REG_3__6__SCAN_IN, INSTQUEUE_REG_3__5__SCAN_IN, INSTQUEUE_REG_3__4__SCAN_IN, INSTQUEUE_REG_3__3__SCAN_IN, INSTQUEUE_REG_3__2__SCAN_IN, INSTQUEUE_REG_3__1__SCAN_IN, INSTQUEUE_REG_3__0__SCAN_IN, INSTQUEUE_REG_2__7__SCAN_IN, INSTQUEUE_REG_2__6__SCAN_IN, INSTQUEUE_REG_2__5__SCAN_IN, INSTQUEUE_REG_2__4__SCAN_IN, INSTQUEUE_REG_2__3__SCAN_IN, INSTQUEUE_REG_2__2__SCAN_IN, INSTQUEUE_REG_2__1__SCAN_IN, INSTQUEUE_REG_2__0__SCAN_IN, INSTQUEUE_REG_1__7__SCAN_IN, INSTQUEUE_REG_1__6__SCAN_IN, INSTQUEUE_REG_1__5__SCAN_IN, INSTQUEUE_REG_1__4__SCAN_IN, INSTQUEUE_REG_1__3__SCAN_IN, INSTQUEUE_REG_1__2__SCAN_IN, INSTQUEUE_REG_1__1__SCAN_IN, INSTQUEUE_REG_1__0__SCAN_IN, INSTQUEUE_REG_0__7__SCAN_IN, INSTQUEUE_REG_0__6__SCAN_IN, INSTQUEUE_REG_0__5__SCAN_IN, INSTQUEUE_REG_0__4__SCAN_IN, INSTQUEUE_REG_0__3__SCAN_IN, INSTQUEUE_REG_0__2__SCAN_IN, INSTQUEUE_REG_0__1__SCAN_IN, INSTQUEUE_REG_0__0__SCAN_IN, INSTQUEUERD_ADDR_REG_4__SCAN_IN, INSTQUEUERD_ADDR_REG_3__SCAN_IN, INSTQUEUERD_ADDR_REG_2__SCAN_IN, INSTQUEUERD_ADDR_REG_1__SCAN_IN, INSTQUEUERD_ADDR_REG_0__SCAN_IN, INSTQUEUEWR_ADDR_REG_4__SCAN_IN, INSTQUEUEWR_ADDR_REG_3__SCAN_IN, INSTQUEUEWR_ADDR_REG_2__SCAN_IN, INSTQUEUEWR_ADDR_REG_1__SCAN_IN, INSTQUEUEWR_ADDR_REG_0__SCAN_IN, INSTADDRPOINTER_REG_0__SCAN_IN, INSTADDRPOINTER_REG_1__SCAN_IN, INSTADDRPOINTER_REG_2__SCAN_IN, INSTADDRPOINTER_REG_3__SCAN_IN, INSTADDRPOINTER_REG_4__SCAN_IN, INSTADDRPOINTER_REG_5__SCAN_IN, INSTADDRPOINTER_REG_6__SCAN_IN, INSTADDRPOINTER_REG_7__SCAN_IN, INSTADDRPOINTER_REG_8__SCAN_IN, INSTADDRPOINTER_REG_9__SCAN_IN, INSTADDRPOINTER_REG_10__SCAN_IN, INSTADDRPOINTER_REG_11__SCAN_IN, INSTADDRPOINTER_REG_12__SCAN_IN, INSTADDRPOINTER_REG_13__SCAN_IN, INSTADDRPOINTER_REG_14__SCAN_IN, INSTADDRPOINTER_REG_15__SCAN_IN, INSTADDRPOINTER_REG_16__SCAN_IN, INSTADDRPOINTER_REG_17__SCAN_IN, INSTADDRPOINTER_REG_18__SCAN_IN, INSTADDRPOINTER_REG_19__SCAN_IN, INSTADDRPOINTER_REG_20__SCAN_IN, INSTADDRPOINTER_REG_21__SCAN_IN, INSTADDRPOINTER_REG_22__SCAN_IN, INSTADDRPOINTER_REG_23__SCAN_IN, INSTADDRPOINTER_REG_24__SCAN_IN, INSTADDRPOINTER_REG_25__SCAN_IN, INSTADDRPOINTER_REG_26__SCAN_IN, INSTADDRPOINTER_REG_27__SCAN_IN, INSTADDRPOINTER_REG_28__SCAN_IN, INSTADDRPOINTER_REG_29__SCAN_IN, INSTADDRPOINTER_REG_30__SCAN_IN, INSTADDRPOINTER_REG_31__SCAN_IN, PHYADDRPOINTER_REG_0__SCAN_IN, PHYADDRPOINTER_REG_1__SCAN_IN, PHYADDRPOINTER_REG_2__SCAN_IN, PHYADDRPOINTER_REG_3__SCAN_IN, PHYADDRPOINTER_REG_4__SCAN_IN, PHYADDRPOINTER_REG_5__SCAN_IN, PHYADDRPOINTER_REG_6__SCAN_IN, PHYADDRPOINTER_REG_7__SCAN_IN, PHYADDRPOINTER_REG_8__SCAN_IN, PHYADDRPOINTER_REG_9__SCAN_IN, PHYADDRPOINTER_REG_10__SCAN_IN, PHYADDRPOINTER_REG_11__SCAN_IN, PHYADDRPOINTER_REG_12__SCAN_IN, PHYADDRPOINTER_REG_13__SCAN_IN, PHYADDRPOINTER_REG_14__SCAN_IN, PHYADDRPOINTER_REG_15__SCAN_IN, PHYADDRPOINTER_REG_16__SCAN_IN, PHYADDRPOINTER_REG_17__SCAN_IN, PHYADDRPOINTER_REG_18__SCAN_IN, PHYADDRPOINTER_REG_19__SCAN_IN, PHYADDRPOINTER_REG_20__SCAN_IN, PHYADDRPOINTER_REG_21__SCAN_IN, PHYADDRPOINTER_REG_22__SCAN_IN, PHYADDRPOINTER_REG_23__SCAN_IN, PHYADDRPOINTER_REG_24__SCAN_IN, PHYADDRPOINTER_REG_25__SCAN_IN, PHYADDRPOINTER_REG_26__SCAN_IN, PHYADDRPOINTER_REG_27__SCAN_IN, PHYADDRPOINTER_REG_28__SCAN_IN, PHYADDRPOINTER_REG_29__SCAN_IN, PHYADDRPOINTER_REG_30__SCAN_IN, PHYADDRPOINTER_REG_31__SCAN_IN, LWORD_REG_15__SCAN_IN, LWORD_REG_14__SCAN_IN, LWORD_REG_13__SCAN_IN, LWORD_REG_12__SCAN_IN, LWORD_REG_11__SCAN_IN, LWORD_REG_10__SCAN_IN, LWORD_REG_9__SCAN_IN, LWORD_REG_8__SCAN_IN, LWORD_REG_7__SCAN_IN, LWORD_REG_6__SCAN_IN, LWORD_REG_5__SCAN_IN, LWORD_REG_4__SCAN_IN, LWORD_REG_3__SCAN_IN, LWORD_REG_2__SCAN_IN, LWORD_REG_1__SCAN_IN, LWORD_REG_0__SCAN_IN, UWORD_REG_14__SCAN_IN, UWORD_REG_13__SCAN_IN, UWORD_REG_12__SCAN_IN, UWORD_REG_11__SCAN_IN, UWORD_REG_10__SCAN_IN, UWORD_REG_9__SCAN_IN, UWORD_REG_8__SCAN_IN, UWORD_REG_7__SCAN_IN, UWORD_REG_6__SCAN_IN, UWORD_REG_5__SCAN_IN, UWORD_REG_4__SCAN_IN, UWORD_REG_3__SCAN_IN, UWORD_REG_2__SCAN_IN, UWORD_REG_1__SCAN_IN, UWORD_REG_0__SCAN_IN, EAX_REG_0__SCAN_IN, EAX_REG_1__SCAN_IN, EAX_REG_2__SCAN_IN, EAX_REG_3__SCAN_IN, EAX_REG_4__SCAN_IN, EAX_REG_5__SCAN_IN, EAX_REG_6__SCAN_IN, EAX_REG_7__SCAN_IN, EAX_REG_8__SCAN_IN, EAX_REG_9__SCAN_IN, EAX_REG_10__SCAN_IN, EAX_REG_11__SCAN_IN, EAX_REG_12__SCAN_IN, EAX_REG_13__SCAN_IN, EAX_REG_14__SCAN_IN, EAX_REG_15__SCAN_IN, EAX_REG_16__SCAN_IN, EAX_REG_17__SCAN_IN, EAX_REG_18__SCAN_IN, EAX_REG_19__SCAN_IN, EAX_REG_20__SCAN_IN, EAX_REG_21__SCAN_IN, EAX_REG_22__SCAN_IN, EAX_REG_23__SCAN_IN, EAX_REG_24__SCAN_IN, EAX_REG_25__SCAN_IN, EAX_REG_26__SCAN_IN, EAX_REG_27__SCAN_IN, EAX_REG_28__SCAN_IN, EAX_REG_29__SCAN_IN, EAX_REG_30__SCAN_IN, EAX_REG_31__SCAN_IN, EBX_REG_0__SCAN_IN, EBX_REG_1__SCAN_IN, EBX_REG_2__SCAN_IN, EBX_REG_3__SCAN_IN, EBX_REG_4__SCAN_IN, EBX_REG_5__SCAN_IN, EBX_REG_6__SCAN_IN, EBX_REG_7__SCAN_IN, EBX_REG_8__SCAN_IN, EBX_REG_9__SCAN_IN, EBX_REG_10__SCAN_IN, EBX_REG_11__SCAN_IN, EBX_REG_12__SCAN_IN, EBX_REG_13__SCAN_IN, EBX_REG_14__SCAN_IN, EBX_REG_15__SCAN_IN, EBX_REG_16__SCAN_IN, EBX_REG_17__SCAN_IN, EBX_REG_18__SCAN_IN, EBX_REG_19__SCAN_IN, EBX_REG_20__SCAN_IN, EBX_REG_21__SCAN_IN, EBX_REG_22__SCAN_IN, EBX_REG_23__SCAN_IN, EBX_REG_24__SCAN_IN, EBX_REG_25__SCAN_IN, EBX_REG_26__SCAN_IN, EBX_REG_27__SCAN_IN, EBX_REG_28__SCAN_IN, EBX_REG_29__SCAN_IN, EBX_REG_30__SCAN_IN, EBX_REG_31__SCAN_IN, REIP_REG_0__SCAN_IN, REIP_REG_1__SCAN_IN, REIP_REG_2__SCAN_IN, REIP_REG_3__SCAN_IN, REIP_REG_4__SCAN_IN, REIP_REG_5__SCAN_IN, REIP_REG_6__SCAN_IN, REIP_REG_7__SCAN_IN, REIP_REG_8__SCAN_IN, REIP_REG_9__SCAN_IN, REIP_REG_10__SCAN_IN, REIP_REG_11__SCAN_IN, REIP_REG_12__SCAN_IN, REIP_REG_13__SCAN_IN, REIP_REG_14__SCAN_IN, REIP_REG_15__SCAN_IN, perturb_signal, restore_signal;
  output DATAO_REG_25__SCAN_IN_BUFF, DATAO_REG_5__SCAN_IN_BUFF, DATAO_REG_28__SCAN_IN_BUFF, DATAO_REG_21__SCAN_IN_BUFF, BE_N_REG_0__SCAN_IN_BUFF, ADDRESS_REG_23__SCAN_IN_BUFF, ADDRESS_REG_17__SCAN_IN_BUFF, ADDRESS_REG_2__SCAN_IN_BUFF, DATAO_REG_30__SCAN_IN_BUFF, BE_N_REG_1__SCAN_IN_BUFF, ADDRESS_REG_1__SCAN_IN_BUFF, DATAO_REG_8__SCAN_IN_BUFF, DATAO_REG_23__SCAN_IN_BUFF, DATAO_REG_10__SCAN_IN_BUFF, ADDRESS_REG_22__SCAN_IN_BUFF, ADDRESS_REG_11__SCAN_IN_BUFF, ADDRESS_REG_3__SCAN_IN_BUFF, BE_N_REG_3__SCAN_IN_BUFF, DATAO_REG_27__SCAN_IN_BUFF, ADDRESS_REG_10__SCAN_IN_BUFF, ADDRESS_REG_28__SCAN_IN_BUFF, DATAO_REG_12__SCAN_IN_BUFF, BE_N_REG_2__SCAN_IN_BUFF, ADDRESS_REG_13__SCAN_IN_BUFF, DATAO_REG_13__SCAN_IN_BUFF, ADDRESS_REG_20__SCAN_IN_BUFF, DATAO_REG_24__SCAN_IN_BUFF, DATAO_REG_9__SCAN_IN_BUFF, DATAO_REG_7__SCAN_IN_BUFF, DATAO_REG_11__SCAN_IN_BUFF, ADDRESS_REG_19__SCAN_IN_BUFF, ADDRESS_REG_27__SCAN_IN_BUFF, ADDRESS_REG_25__SCAN_IN_BUFF, ADDRESS_REG_29__SCAN_IN_BUFF, ADDRESS_REG_5__SCAN_IN_BUFF, ADDRESS_REG_7__SCAN_IN_BUFF, ADDRESS_REG_8__SCAN_IN_BUFF, ADDRESS_REG_21__SCAN_IN_BUFF, DATAO_REG_20__SCAN_IN_BUFF, DATAO_REG_17__SCAN_IN_BUFF, DATAO_REG_6__SCAN_IN_BUFF, ADDRESS_REG_14__SCAN_IN_BUFF, DATAO_REG_19__SCAN_IN_BUFF, ADS_N_REG_SCAN_IN_BUFF, DATAO_REG_15__SCAN_IN_BUFF, DATAO_REG_26__SCAN_IN_BUFF, DATAO_REG_3__SCAN_IN_BUFF, DATAO_REG_1__SCAN_IN_BUFF, ADDRESS_REG_26__SCAN_IN_BUFF, ADDRESS_REG_18__SCAN_IN_BUFF, M_IO_N_REG_SCAN_IN_BUFF, DATAO_REG_31__SCAN_IN_BUFF, ADDRESS_REG_16__SCAN_IN_BUFF, ADDRESS_REG_9__SCAN_IN_BUFF, ADDRESS_REG_12__SCAN_IN_BUFF, DATAO_REG_29__SCAN_IN_BUFF, DATAO_REG_0__SCAN_IN_BUFF, ADDRESS_REG_4__SCAN_IN_BUFF, D_C_N_REG_SCAN_IN_BUFF, DATAO_REG_4__SCAN_IN_BUFF, ADDRESS_REG_6__SCAN_IN_BUFF, DATAO_REG_2__SCAN_IN_BUFF, ADDRESS_REG_0__SCAN_IN_BUFF, DATAO_REG_18__SCAN_IN_BUFF, DATAO_REG_16__SCAN_IN_BUFF, ADDRESS_REG_24__SCAN_IN_BUFF, DATAO_REG_14__SCAN_IN_BUFF, W_R_N_REG_SCAN_IN_BUFF, ADDRESS_REG_15__SCAN_IN_BUFF, DATAO_REG_22__SCAN_IN_BUFF, U3445, U3446, U3447, U3448, U3213, U3212, U3211, U3210, U3209, U3208, U3207, U3206, U3205, U3204, U3203, U3202, U3201, U3200, U3199, U3198, U3197, U3196, U3195, U3194, U3193, U3192, U3191, U3190, U3189, U3188, U3187, U3186, U3185, U3184, U3183, U3182, U3181, U3451, U3452, U3180, U3179, U3178, U3177, U3176, U3175, U3174, U3173, U3172, U3171, U3170, U3169, U3168, U3167, U3166, U3165, U3164, U3163, U3162, U3161, U3160, U3159, U3158, U3157, U3156, U3155, U3154, U3153, U3152, U3151, U3453, U3150, U3149, U3148, U3147, U3146, U3145, U3144, U3143, U3142, U3141, U3140, U3139, U3138, U3137, U3136, U3135, U3134, U3133, U3132, U3131, U3130, U3129, U3128, U3127, U3126, U3125, U3124, U3123, U3122, U3121, U3120, U3119, U3118, U3117, U3116, U3115, U3114, U3113, U3112, U3111, U3110, U3109, U3108, U3107, U3106, U3105, U3104, U3103, U3102, U3101, U3100, U3099, U3098, U3097, U3096, U3095, U3094, U3093, U3092, U3091, U3090, U3089, U3088, U3087, U3086, U3085, U3084, U3083, U3082, U3081, U3080, U3079, U3078, U3077, U3076, U3075, U3074, U3073, U3072, U3071, U3070, U3069, U3068, U3067, U3066, U3065, U3064, U3063, U3062, U3061, U3060, U3059, U3058, U3057, U3056, U3055, U3054, U3053, U3052, U3051, U3050, U3049, U3048, U3047, U3046, U3045, U3044, U3043, U3042, U3041, U3040, U3039, U3038, U3037, U3036, U3035, U3034, U3033, U3032, U3031, U3030, U3029, U3028, U3027, U3026, U3025, U3024, U3023, U3022, U3021, U3020, U3455, U3456, U3459, U3460, U3461, U3019, U3462, U3463, U3464, U3465, U3018, U3017, U3016, U3015, U3014, U3013, U3012, U3011, U3010, U3009, U3008, U3007, U3006, U3005, U3004, U3003, U3002, U3001, U3000, U2999, U2998, U2997, U2996, U2995, U2994, U2993, U2992, U2991, U2990, U2989, U2988, U2987, U2986, U2985, U2984, U2983, U2982, U2981, U2980, U2979, U2978, U2977, U2976, U2975, U2974, U2973, U2972, U2971, U2970, U2969, U2968, U2967, U2966, U2965, U2964, U2963, U2962, U2961, U2960, U2959, U2958, U2957, U2956, U2955, U2954, U2953, U2952, U2951, U2950, U2949, U2948, U2947, U2946, U2945, U2944, U2943, U2942, U2941, U2940, U2939, U2938, U2937, U2936, U2935, U2934, U2933, U2932, U2931, U2930, U2929, U2928, U2927, U2926, U2925, U2924, U2923, U2922, U2921, U2920, U2919, U2918, U2917, U2916, U2915, U2914, U2913, U2912, U2911, U2910, U2909, U2908, U2907, U2906, U2905, U2904, U2903, U2902, U2901, U2900, U2899, U2898, U2897, U2896, U2895, U2894, U2893, U2892, U2891, U2890, U2889, U2888, U2887, U2886, U2885, U2884, U2883, U2882, U2881, U2880, U2879, U2878, U2877, U2876, U2875, U2874, U2873, U2872, U2871, U2870, U2869, U2868, U2867, U2866, U2865, U2864, U2863, U2862, U2861, U2860, U2859, U2858, U2857, U2856, U2855, U2854, U2853, U2852, U2851, U2850, U2849, U2848, U2847, U2846, U2845, U2844, U2843, U2842, U2841, U2840, U2839, U2838, U2837, U2836, U2835, U2834, U2833, U2832, U2831, U2830, U2829, U2828, U2827, U2826, U2825, U2824, U2823, U2822, U2821, U2820, U2819, U2818, U2817, U2816, U2815, U2814, U2813, U2812, U2811, U2810, U2809, U2808, U2807, U2806, U2805, U2804, U2803, U2802, U2801, U2800, U2799, U2798, U2797, U2796, U2795, U3468, U2794, U3469, U3470, U2793, U3471, U2792, U3472, U2791, U3473, U2790, U2789, U3474, U2788;
  wire ADD_371_U10, ADD_371_U11, ADD_371_U12, ADD_371_U13, ADD_371_U14, ADD_371_U15, ADD_371_U16, ADD_371_U17, ADD_371_U18, ADD_371_U19, ADD_371_U20, ADD_371_U21, ADD_371_U22, ADD_371_U23, ADD_371_U24, ADD_371_U25, ADD_371_U26, ADD_371_U27, ADD_371_U28, ADD_371_U29, ADD_371_U30, ADD_371_U31, ADD_371_U32, ADD_371_U33, ADD_371_U34, ADD_371_U35, ADD_371_U36, ADD_371_U37, ADD_371_U38, ADD_371_U39, ADD_371_U4, ADD_371_U40, ADD_371_U41, ADD_371_U42, ADD_371_U43, ADD_371_U44, ADD_371_U5, ADD_371_U6, ADD_371_U7, ADD_371_U8, ADD_371_U9, ADD_405_U10, ADD_405_U100, ADD_405_U101, ADD_405_U102, ADD_405_U103, ADD_405_U104, ADD_405_U105, ADD_405_U106, ADD_405_U107, ADD_405_U108, ADD_405_U109, ADD_405_U11, ADD_405_U110, ADD_405_U111, ADD_405_U112, ADD_405_U113, ADD_405_U114, ADD_405_U115, ADD_405_U116, ADD_405_U117, ADD_405_U118, ADD_405_U119, ADD_405_U12, ADD_405_U120, ADD_405_U121, ADD_405_U122, ADD_405_U123, ADD_405_U124, ADD_405_U125, ADD_405_U126, ADD_405_U127, ADD_405_U128, ADD_405_U129, ADD_405_U13, ADD_405_U130, ADD_405_U131, ADD_405_U132, ADD_405_U133, ADD_405_U134, ADD_405_U135, ADD_405_U136, ADD_405_U137, ADD_405_U138, ADD_405_U139, ADD_405_U14, ADD_405_U140, ADD_405_U141, ADD_405_U142, ADD_405_U143, ADD_405_U144, ADD_405_U145, ADD_405_U146, ADD_405_U147, ADD_405_U148, ADD_405_U149, ADD_405_U15, ADD_405_U150, ADD_405_U151, ADD_405_U152, ADD_405_U153, ADD_405_U154, ADD_405_U155, ADD_405_U156, ADD_405_U157, ADD_405_U158, ADD_405_U159, ADD_405_U16, ADD_405_U160, ADD_405_U161, ADD_405_U162, ADD_405_U163, ADD_405_U164, ADD_405_U165, ADD_405_U166, ADD_405_U167, ADD_405_U168, ADD_405_U169, ADD_405_U17, ADD_405_U170, ADD_405_U171, ADD_405_U172, ADD_405_U173, ADD_405_U174, ADD_405_U175, ADD_405_U176, ADD_405_U177, ADD_405_U178, ADD_405_U179, ADD_405_U18, ADD_405_U180, ADD_405_U181, ADD_405_U182, ADD_405_U183, ADD_405_U184, ADD_405_U185, ADD_405_U186, ADD_405_U19, ADD_405_U20, ADD_405_U21, ADD_405_U22, ADD_405_U23, ADD_405_U24, ADD_405_U25, ADD_405_U26, ADD_405_U27, ADD_405_U28, ADD_405_U29, ADD_405_U30, ADD_405_U31, ADD_405_U32, ADD_405_U33, ADD_405_U34, ADD_405_U35, ADD_405_U36, ADD_405_U37, ADD_405_U38, ADD_405_U39, ADD_405_U4, ADD_405_U40, ADD_405_U41, ADD_405_U42, ADD_405_U43, ADD_405_U44, ADD_405_U45, ADD_405_U46, ADD_405_U47, ADD_405_U48, ADD_405_U49, ADD_405_U5, ADD_405_U50, ADD_405_U51, ADD_405_U52, ADD_405_U53, ADD_405_U54, ADD_405_U55, ADD_405_U56, ADD_405_U57, ADD_405_U58, ADD_405_U59, ADD_405_U6, ADD_405_U60, ADD_405_U61, ADD_405_U62, ADD_405_U63, ADD_405_U64, ADD_405_U65, ADD_405_U66, ADD_405_U67, ADD_405_U68, ADD_405_U69, ADD_405_U7, ADD_405_U70, ADD_405_U71, ADD_405_U72, ADD_405_U73, ADD_405_U74, ADD_405_U75, ADD_405_U76, ADD_405_U77, ADD_405_U78, ADD_405_U79, ADD_405_U8, ADD_405_U80, ADD_405_U81, ADD_405_U82, ADD_405_U83, ADD_405_U84, ADD_405_U85, ADD_405_U86, ADD_405_U87, ADD_405_U88, ADD_405_U89, ADD_405_U9, ADD_405_U90, ADD_405_U91, ADD_405_U92, ADD_405_U93, ADD_405_U94, ADD_405_U95, ADD_405_U96, ADD_405_U97, ADD_405_U98, ADD_405_U99, ADD_515_U10, ADD_515_U100, ADD_515_U101, ADD_515_U102, ADD_515_U103, ADD_515_U104, ADD_515_U105, ADD_515_U106, ADD_515_U107, ADD_515_U108, ADD_515_U109, ADD_515_U11, ADD_515_U110, ADD_515_U111, ADD_515_U112, ADD_515_U113, ADD_515_U114, ADD_515_U115, ADD_515_U116, ADD_515_U117, ADD_515_U118, ADD_515_U119, ADD_515_U12, ADD_515_U120, ADD_515_U121, ADD_515_U122, ADD_515_U123, ADD_515_U124, ADD_515_U125, ADD_515_U126, ADD_515_U127, ADD_515_U128, ADD_515_U129, ADD_515_U13, ADD_515_U130, ADD_515_U131, ADD_515_U132, ADD_515_U133, ADD_515_U134, ADD_515_U135, ADD_515_U136, ADD_515_U137, ADD_515_U138, ADD_515_U139, ADD_515_U14, ADD_515_U140, ADD_515_U141, ADD_515_U142, ADD_515_U143, ADD_515_U144, ADD_515_U145, ADD_515_U146, ADD_515_U147, ADD_515_U148, ADD_515_U149, ADD_515_U15, ADD_515_U150, ADD_515_U151, ADD_515_U152, ADD_515_U153, ADD_515_U154, ADD_515_U155, ADD_515_U156, ADD_515_U157, ADD_515_U158, ADD_515_U159, ADD_515_U16, ADD_515_U160, ADD_515_U161, ADD_515_U162, ADD_515_U163, ADD_515_U164, ADD_515_U165, ADD_515_U166, ADD_515_U167, ADD_515_U168, ADD_515_U169, ADD_515_U17, ADD_515_U170, ADD_515_U171, ADD_515_U172, ADD_515_U173, ADD_515_U174, ADD_515_U175, ADD_515_U176, ADD_515_U177, ADD_515_U178, ADD_515_U179, ADD_515_U18, ADD_515_U180, ADD_515_U181, ADD_515_U182, ADD_515_U19, ADD_515_U20, ADD_515_U21, ADD_515_U22, ADD_515_U23, ADD_515_U24, ADD_515_U25, ADD_515_U26, ADD_515_U27, ADD_515_U28, ADD_515_U29, ADD_515_U30, ADD_515_U31, ADD_515_U32, ADD_515_U33, ADD_515_U34, ADD_515_U35, ADD_515_U36, ADD_515_U37, ADD_515_U38, ADD_515_U39, ADD_515_U4, ADD_515_U40, ADD_515_U41, ADD_515_U42, ADD_515_U43, ADD_515_U44, ADD_515_U45, ADD_515_U46, ADD_515_U47, ADD_515_U48, ADD_515_U49, ADD_515_U5, ADD_515_U50, ADD_515_U51, ADD_515_U52, ADD_515_U53, ADD_515_U54, ADD_515_U55, ADD_515_U56, ADD_515_U57, ADD_515_U58, ADD_515_U59, ADD_515_U6, ADD_515_U60, ADD_515_U61, ADD_515_U62, ADD_515_U63, ADD_515_U64, ADD_515_U65, ADD_515_U66, ADD_515_U67, ADD_515_U68, ADD_515_U69, ADD_515_U7, ADD_515_U70, ADD_515_U71, ADD_515_U72, ADD_515_U73, ADD_515_U74, ADD_515_U75, ADD_515_U76, ADD_515_U77, ADD_515_U78, ADD_515_U79, ADD_515_U8, ADD_515_U80, ADD_515_U81, ADD_515_U82, ADD_515_U83, ADD_515_U84, ADD_515_U85, ADD_515_U86, ADD_515_U87, ADD_515_U88, ADD_515_U89, ADD_515_U9, ADD_515_U90, ADD_515_U91, ADD_515_U92, ADD_515_U93, ADD_515_U94, ADD_515_U95, ADD_515_U96, ADD_515_U97, ADD_515_U98, ADD_515_U99, GTE_485_U6, GTE_485_U7, LT_563_1260_U6, LT_563_1260_U7, LT_563_1260_U8, LT_563_1260_U9, LT_563_U10, LT_563_U11, LT_563_U12, LT_563_U13, LT_563_U14, LT_563_U15, LT_563_U16, LT_563_U17, LT_563_U18, LT_563_U19, LT_563_U20, LT_563_U21, LT_563_U22, LT_563_U23, LT_563_U24, LT_563_U25, LT_563_U26, LT_563_U27, LT_563_U28, LT_563_U6, LT_563_U7, LT_563_U8, LT_563_U9, LT_589_U6, LT_589_U7, LT_589_U8, R2027_U10, R2027_U100, R2027_U101, R2027_U102, R2027_U103, R2027_U104, R2027_U105, R2027_U106, R2027_U107, R2027_U108, R2027_U109, R2027_U11, R2027_U110, R2027_U111, R2027_U112, R2027_U113, R2027_U114, R2027_U115, R2027_U116, R2027_U117, R2027_U118, R2027_U119, R2027_U12, R2027_U120, R2027_U121, R2027_U122, R2027_U123, R2027_U124, R2027_U125, R2027_U126, R2027_U127, R2027_U128, R2027_U129, R2027_U13, R2027_U130, R2027_U131, R2027_U132, R2027_U133, R2027_U134, R2027_U135, R2027_U136, R2027_U137, R2027_U138, R2027_U139, R2027_U14, R2027_U140, R2027_U141, R2027_U142, R2027_U143, R2027_U144, R2027_U145, R2027_U146, R2027_U147, R2027_U148, R2027_U149, R2027_U15, R2027_U150, R2027_U151, R2027_U152, R2027_U153, R2027_U154, R2027_U155, R2027_U156, R2027_U157, R2027_U158, R2027_U159, R2027_U16, R2027_U160, R2027_U161, R2027_U162, R2027_U163, R2027_U164, R2027_U165, R2027_U166, R2027_U167, R2027_U168, R2027_U169, R2027_U17, R2027_U170, R2027_U171, R2027_U172, R2027_U173, R2027_U174, R2027_U175, R2027_U176, R2027_U177, R2027_U178, R2027_U179, R2027_U18, R2027_U180, R2027_U181, R2027_U182, R2027_U183, R2027_U184, R2027_U185, R2027_U186, R2027_U187, R2027_U188, R2027_U189, R2027_U19, R2027_U190, R2027_U191, R2027_U192, R2027_U193, R2027_U194, R2027_U195, R2027_U196, R2027_U197, R2027_U198, R2027_U199, R2027_U20, R2027_U200, R2027_U201, R2027_U202, R2027_U21, R2027_U22, R2027_U23, R2027_U24, R2027_U25, R2027_U26, R2027_U27, R2027_U28, R2027_U29, R2027_U30, R2027_U31, R2027_U32, R2027_U33, R2027_U34, R2027_U35, R2027_U36, R2027_U37, R2027_U38, R2027_U39, R2027_U40, R2027_U41, R2027_U42, R2027_U43, R2027_U44, R2027_U45, R2027_U46, R2027_U47, R2027_U48, R2027_U49, R2027_U5, R2027_U50, R2027_U51, R2027_U52, R2027_U53, R2027_U54, R2027_U55, R2027_U56, R2027_U57, R2027_U58, R2027_U59, R2027_U6, R2027_U60, R2027_U61, R2027_U62, R2027_U63, R2027_U64, R2027_U65, R2027_U66, R2027_U67, R2027_U68, R2027_U69, R2027_U7, R2027_U70, R2027_U71, R2027_U72, R2027_U73, R2027_U74, R2027_U75, R2027_U76, R2027_U77, R2027_U78, R2027_U79, R2027_U8, R2027_U80, R2027_U81, R2027_U82, R2027_U83, R2027_U84, R2027_U85, R2027_U86, R2027_U87, R2027_U88, R2027_U89, R2027_U9, R2027_U90, R2027_U91, R2027_U92, R2027_U93, R2027_U94, R2027_U95, R2027_U96, R2027_U97, R2027_U98, R2027_U99, R2096_U10, R2096_U100, R2096_U101, R2096_U102, R2096_U103, R2096_U104, R2096_U105, R2096_U106, R2096_U107, R2096_U108, R2096_U109, R2096_U11, R2096_U110, R2096_U111, R2096_U112, R2096_U113, R2096_U114, R2096_U115, R2096_U116, R2096_U117, R2096_U118, R2096_U119, R2096_U12, R2096_U120, R2096_U121, R2096_U122, R2096_U123, R2096_U124, R2096_U125, R2096_U126, R2096_U127, R2096_U128, R2096_U129, R2096_U13, R2096_U130, R2096_U131, R2096_U132, R2096_U133, R2096_U134, R2096_U135, R2096_U136, R2096_U137, R2096_U138, R2096_U139, R2096_U14, R2096_U140, R2096_U141, R2096_U142, R2096_U143, R2096_U144, R2096_U145, R2096_U146, R2096_U147, R2096_U148, R2096_U149, R2096_U15, R2096_U150, R2096_U151, R2096_U152, R2096_U153, R2096_U154, R2096_U155, R2096_U156, R2096_U157, R2096_U158, R2096_U159, R2096_U16, R2096_U160, R2096_U161, R2096_U162, R2096_U163, R2096_U164, R2096_U165, R2096_U166, R2096_U167, R2096_U168, R2096_U169, R2096_U17, R2096_U170, R2096_U171, R2096_U172, R2096_U173, R2096_U174, R2096_U175, R2096_U176, R2096_U177, R2096_U178, R2096_U179, R2096_U18, R2096_U180, R2096_U181, R2096_U182, R2096_U19, R2096_U20, R2096_U21, R2096_U22, R2096_U23, R2096_U24, R2096_U25, R2096_U26, R2096_U27, R2096_U28, R2096_U29, R2096_U30, R2096_U31, R2096_U32, R2096_U33, R2096_U34, R2096_U35, R2096_U36, R2096_U37, R2096_U38, R2096_U39, R2096_U4, R2096_U40, R2096_U41, R2096_U42, R2096_U43, R2096_U44, R2096_U45, R2096_U46, R2096_U47, R2096_U48, R2096_U49, R2096_U5, R2096_U50, R2096_U51, R2096_U52, R2096_U53, R2096_U54, R2096_U55, R2096_U56, R2096_U57, R2096_U58, R2096_U59, R2096_U6, R2096_U60, R2096_U61, R2096_U62, R2096_U63, R2096_U64, R2096_U65, R2096_U66, R2096_U67, R2096_U68, R2096_U69, R2096_U7, R2096_U70, R2096_U71, R2096_U72, R2096_U73, R2096_U74, R2096_U75, R2096_U76, R2096_U77, R2096_U78, R2096_U79, R2096_U8, R2096_U80, R2096_U81, R2096_U82, R2096_U83, R2096_U84, R2096_U85, R2096_U86, R2096_U87, R2096_U88, R2096_U89, R2096_U9, R2096_U90, R2096_U91, R2096_U92, R2096_U93, R2096_U94, R2096_U95, R2096_U96, R2096_U97, R2096_U98, R2096_U99, R2099_U10, R2099_U100, R2099_U101, R2099_U102, R2099_U103, R2099_U104, R2099_U105, R2099_U106, R2099_U107, R2099_U108, R2099_U109, R2099_U11, R2099_U110, R2099_U111, R2099_U112, R2099_U113, R2099_U114, R2099_U115, R2099_U116, R2099_U117, R2099_U118, R2099_U119, R2099_U12, R2099_U120, R2099_U121, R2099_U122, R2099_U123, R2099_U124, R2099_U125, R2099_U126, R2099_U127, R2099_U128, R2099_U129, R2099_U13, R2099_U130, R2099_U131, R2099_U132, R2099_U133, R2099_U134, R2099_U135, R2099_U136, R2099_U137, R2099_U138, R2099_U139, R2099_U14, R2099_U140, R2099_U141, R2099_U142, R2099_U143, R2099_U144, R2099_U145, R2099_U146, R2099_U147, R2099_U148, R2099_U149, R2099_U15, R2099_U150, R2099_U151, R2099_U152, R2099_U153, R2099_U154, R2099_U155, R2099_U156, R2099_U157, R2099_U158, R2099_U159, R2099_U16, R2099_U160, R2099_U161, R2099_U162, R2099_U163, R2099_U164, R2099_U165, R2099_U166, R2099_U167, R2099_U168, R2099_U169, R2099_U17, R2099_U170, R2099_U171, R2099_U172, R2099_U173, R2099_U174, R2099_U175, R2099_U176, R2099_U177, R2099_U178, R2099_U179, R2099_U18, R2099_U180, R2099_U181, R2099_U182, R2099_U183, R2099_U184, R2099_U185, R2099_U186, R2099_U187, R2099_U188, R2099_U189, R2099_U19, R2099_U190, R2099_U191, R2099_U192, R2099_U193, R2099_U194, R2099_U195, R2099_U196, R2099_U197, R2099_U198, R2099_U199, R2099_U20, R2099_U200, R2099_U201, R2099_U202, R2099_U203, R2099_U204, R2099_U205, R2099_U206, R2099_U207, R2099_U208, R2099_U209, R2099_U21, R2099_U210, R2099_U211, R2099_U212, R2099_U213, R2099_U214, R2099_U215, R2099_U216, R2099_U217, R2099_U218, R2099_U219, R2099_U22, R2099_U220, R2099_U221, R2099_U222, R2099_U223, R2099_U224, R2099_U225, R2099_U226, R2099_U227, R2099_U228, R2099_U229, R2099_U23, R2099_U230, R2099_U231, R2099_U232, R2099_U233, R2099_U234, R2099_U235, R2099_U236, R2099_U237, R2099_U238, R2099_U239, R2099_U24, R2099_U240, R2099_U241, R2099_U242, R2099_U243, R2099_U244, R2099_U245, R2099_U246, R2099_U247, R2099_U248, R2099_U249, R2099_U25, R2099_U250, R2099_U251, R2099_U252, R2099_U253, R2099_U254, R2099_U255, R2099_U256, R2099_U257, R2099_U258, R2099_U259, R2099_U26, R2099_U260, R2099_U261, R2099_U262, R2099_U263, R2099_U264, R2099_U265, R2099_U266, R2099_U267, R2099_U268, R2099_U269, R2099_U27, R2099_U270, R2099_U271, R2099_U272, R2099_U273, R2099_U274, R2099_U275, R2099_U276, R2099_U277, R2099_U278, R2099_U279, R2099_U28, R2099_U280, R2099_U281, R2099_U282, R2099_U283, R2099_U284, R2099_U285, R2099_U286, R2099_U287, R2099_U288, R2099_U289, R2099_U29, R2099_U290, R2099_U291, R2099_U292, R2099_U293, R2099_U294, R2099_U295, R2099_U296, R2099_U297, R2099_U298, R2099_U299, R2099_U30, R2099_U300, R2099_U301, R2099_U302, R2099_U303, R2099_U304, R2099_U305, R2099_U306, R2099_U307, R2099_U308, R2099_U309, R2099_U31, R2099_U310, R2099_U311, R2099_U312, R2099_U313, R2099_U314, R2099_U315, R2099_U316, R2099_U317, R2099_U318, R2099_U319, R2099_U32, R2099_U320, R2099_U321, R2099_U322, R2099_U323, R2099_U324, R2099_U325, R2099_U326, R2099_U327, R2099_U328, R2099_U329, R2099_U33, R2099_U330, R2099_U331, R2099_U332, R2099_U333, R2099_U334, R2099_U335, R2099_U336, R2099_U337, R2099_U338, R2099_U339, R2099_U34, R2099_U340, R2099_U341, R2099_U342, R2099_U343, R2099_U344, R2099_U345, R2099_U346, R2099_U347, R2099_U348, R2099_U349, R2099_U35, R2099_U36, R2099_U37, R2099_U38, R2099_U39, R2099_U4, R2099_U40, R2099_U41, R2099_U42, R2099_U43, R2099_U44, R2099_U45, R2099_U46, R2099_U47, R2099_U48, R2099_U49, R2099_U5, R2099_U50, R2099_U51, R2099_U52, R2099_U53, R2099_U54, R2099_U55, R2099_U56, R2099_U57, R2099_U58, R2099_U59, R2099_U6, R2099_U60, R2099_U61, R2099_U62, R2099_U63, R2099_U64, R2099_U65, R2099_U66, R2099_U67, R2099_U68, R2099_U69, R2099_U7, R2099_U70, R2099_U71, R2099_U72, R2099_U73, R2099_U74, R2099_U75, R2099_U76, R2099_U77, R2099_U78, R2099_U79, R2099_U8, R2099_U80, R2099_U81, R2099_U82, R2099_U83, R2099_U84, R2099_U85, R2099_U86, R2099_U87, R2099_U88, R2099_U89, R2099_U9, R2099_U90, R2099_U91, R2099_U92, R2099_U93, R2099_U94, R2099_U95, R2099_U96, R2099_U97, R2099_U98, R2099_U99, R2144_U10, R2144_U100, R2144_U101, R2144_U102, R2144_U103, R2144_U104, R2144_U105, R2144_U106, R2144_U107, R2144_U108, R2144_U109, R2144_U11, R2144_U110, R2144_U111, R2144_U112, R2144_U113, R2144_U114, R2144_U115, R2144_U116, R2144_U117, R2144_U118, R2144_U119, R2144_U12, R2144_U120, R2144_U121, R2144_U122, R2144_U123, R2144_U124, R2144_U125, R2144_U126, R2144_U127, R2144_U128, R2144_U129, R2144_U13, R2144_U130, R2144_U131, R2144_U132, R2144_U133, R2144_U134, R2144_U135, R2144_U136, R2144_U137, R2144_U138, R2144_U139, R2144_U14, R2144_U140, R2144_U141, R2144_U142, R2144_U143, R2144_U144, R2144_U145, R2144_U146, R2144_U147, R2144_U148, R2144_U149, R2144_U15, R2144_U150, R2144_U151, R2144_U152, R2144_U153, R2144_U154, R2144_U155, R2144_U156, R2144_U157, R2144_U158, R2144_U159, R2144_U16, R2144_U160, R2144_U161, R2144_U162, R2144_U163, R2144_U164, R2144_U165, R2144_U166, R2144_U167, R2144_U168, R2144_U169, R2144_U17, R2144_U170, R2144_U171, R2144_U172, R2144_U173, R2144_U174, R2144_U175, R2144_U176, R2144_U177, R2144_U178, R2144_U179, R2144_U18, R2144_U180, R2144_U181, R2144_U182, R2144_U183, R2144_U184, R2144_U185, R2144_U186, R2144_U187, R2144_U188, R2144_U189, R2144_U19, R2144_U190, R2144_U191, R2144_U192, R2144_U193, R2144_U194, R2144_U195, R2144_U196, R2144_U197, R2144_U198, R2144_U199, R2144_U20, R2144_U200, R2144_U201, R2144_U202, R2144_U203, R2144_U204, R2144_U205, R2144_U206, R2144_U207, R2144_U208, R2144_U209, R2144_U21, R2144_U210, R2144_U211, R2144_U212, R2144_U213, R2144_U214, R2144_U215, R2144_U216, R2144_U217, R2144_U218, R2144_U219, R2144_U22, R2144_U220, R2144_U221, R2144_U222, R2144_U223, R2144_U224, R2144_U225, R2144_U226, R2144_U227, R2144_U228, R2144_U229, R2144_U23, R2144_U230, R2144_U231, R2144_U232, R2144_U233, R2144_U234, R2144_U235, R2144_U236, R2144_U237, R2144_U238, R2144_U239, R2144_U24, R2144_U240, R2144_U241, R2144_U242, R2144_U243, R2144_U244, R2144_U245, R2144_U246, R2144_U247, R2144_U248, R2144_U249, R2144_U25, R2144_U250, R2144_U251, R2144_U252, R2144_U253, R2144_U254, R2144_U255, R2144_U256, R2144_U257, R2144_U258, R2144_U259, R2144_U26, R2144_U260, R2144_U27, R2144_U28, R2144_U29, R2144_U30, R2144_U31, R2144_U32, R2144_U33, R2144_U34, R2144_U35, R2144_U36, R2144_U37, R2144_U38, R2144_U39, R2144_U40, R2144_U41, R2144_U42, R2144_U43, R2144_U44, R2144_U45, R2144_U46, R2144_U47, R2144_U48, R2144_U49, R2144_U5, R2144_U50, R2144_U51, R2144_U52, R2144_U53, R2144_U54, R2144_U55, R2144_U56, R2144_U57, R2144_U58, R2144_U59, R2144_U6, R2144_U60, R2144_U61, R2144_U62, R2144_U63, R2144_U64, R2144_U65, R2144_U66, R2144_U67, R2144_U68, R2144_U69, R2144_U7, R2144_U70, R2144_U71, R2144_U72, R2144_U73, R2144_U74, R2144_U75, R2144_U76, R2144_U77, R2144_U78, R2144_U79, R2144_U8, R2144_U80, R2144_U81, R2144_U82, R2144_U83, R2144_U84, R2144_U85, R2144_U86, R2144_U87, R2144_U88, R2144_U89, R2144_U9, R2144_U90, R2144_U91, R2144_U92, R2144_U93, R2144_U94, R2144_U95, R2144_U96, R2144_U97, R2144_U98, R2144_U99, R2167_U10, R2167_U11, R2167_U12, R2167_U13, R2167_U14, R2167_U15, R2167_U16, R2167_U17, R2167_U18, R2167_U19, R2167_U20, R2167_U21, R2167_U22, R2167_U23, R2167_U24, R2167_U25, R2167_U26, R2167_U27, R2167_U28, R2167_U29, R2167_U30, R2167_U31, R2167_U32, R2167_U33, R2167_U34, R2167_U35, R2167_U36, R2167_U37, R2167_U38, R2167_U39, R2167_U40, R2167_U41, R2167_U42, R2167_U43, R2167_U44, R2167_U45, R2167_U46, R2167_U47, R2167_U48, R2167_U49, R2167_U50, R2167_U6, R2167_U7, R2167_U8, R2167_U9, R2182_U10, R2182_U11, R2182_U12, R2182_U13, R2182_U14, R2182_U15, R2182_U16, R2182_U17, R2182_U18, R2182_U19, R2182_U20, R2182_U21, R2182_U22, R2182_U23, R2182_U24, R2182_U25, R2182_U26, R2182_U27, R2182_U28, R2182_U29, R2182_U30, R2182_U31, R2182_U32, R2182_U33, R2182_U34, R2182_U35, R2182_U36, R2182_U37, R2182_U38, R2182_U39, R2182_U40, R2182_U41, R2182_U42, R2182_U43, R2182_U44, R2182_U45, R2182_U46, R2182_U47, R2182_U48, R2182_U49, R2182_U5, R2182_U50, R2182_U51, R2182_U52, R2182_U53, R2182_U54, R2182_U55, R2182_U56, R2182_U57, R2182_U58, R2182_U59, R2182_U6, R2182_U60, R2182_U61, R2182_U62, R2182_U63, R2182_U64, R2182_U65, R2182_U66, R2182_U67, R2182_U68, R2182_U69, R2182_U7, R2182_U70, R2182_U71, R2182_U72, R2182_U73, R2182_U74, R2182_U75, R2182_U76, R2182_U77, R2182_U78, R2182_U79, R2182_U8, R2182_U80, R2182_U81, R2182_U82, R2182_U83, R2182_U84, R2182_U85, R2182_U86, R2182_U9, R2238_U10, R2238_U11, R2238_U12, R2238_U13, R2238_U14, R2238_U15, R2238_U16, R2238_U17, R2238_U18, R2238_U19, R2238_U20, R2238_U21, R2238_U22, R2238_U23, R2238_U24, R2238_U25, R2238_U26, R2238_U27, R2238_U28, R2238_U29, R2238_U30, R2238_U31, R2238_U32, R2238_U33, R2238_U34, R2238_U35, R2238_U36, R2238_U37, R2238_U38, R2238_U39, R2238_U40, R2238_U41, R2238_U42, R2238_U43, R2238_U44, R2238_U45, R2238_U46, R2238_U47, R2238_U48, R2238_U49, R2238_U50, R2238_U51, R2238_U52, R2238_U53, R2238_U54, R2238_U55, R2238_U56, R2238_U57, R2238_U58, R2238_U59, R2238_U6, R2238_U60, R2238_U61, R2238_U62, R2238_U63, R2238_U64, R2238_U65, R2238_U66, R2238_U7, R2238_U8, R2238_U9, R2278_U10, R2278_U100, R2278_U101, R2278_U102, R2278_U103, R2278_U104, R2278_U105, R2278_U106, R2278_U107, R2278_U108, R2278_U109, R2278_U11, R2278_U110, R2278_U111, R2278_U112, R2278_U113, R2278_U114, R2278_U115, R2278_U116, R2278_U117, R2278_U118, R2278_U119, R2278_U12, R2278_U120, R2278_U121, R2278_U122, R2278_U123, R2278_U124, R2278_U125, R2278_U126, R2278_U127, R2278_U128, R2278_U129, R2278_U13, R2278_U130, R2278_U131, R2278_U132, R2278_U133, R2278_U134, R2278_U135, R2278_U136, R2278_U137, R2278_U138, R2278_U139, R2278_U14, R2278_U140, R2278_U141, R2278_U142, R2278_U143, R2278_U144, R2278_U145, R2278_U146, R2278_U147, R2278_U148, R2278_U149, R2278_U15, R2278_U150, R2278_U151, R2278_U152, R2278_U153, R2278_U154, R2278_U155, R2278_U156, R2278_U157, R2278_U158, R2278_U159, R2278_U16, R2278_U160, R2278_U161, R2278_U162, R2278_U163, R2278_U164, R2278_U165, R2278_U166, R2278_U167, R2278_U168, R2278_U169, R2278_U17, R2278_U170, R2278_U171, R2278_U172, R2278_U173, R2278_U174, R2278_U175, R2278_U176, R2278_U177, R2278_U178, R2278_U179, R2278_U18, R2278_U180, R2278_U181, R2278_U182, R2278_U183, R2278_U184, R2278_U185, R2278_U186, R2278_U187, R2278_U188, R2278_U189, R2278_U19, R2278_U190, R2278_U191, R2278_U192, R2278_U193, R2278_U194, R2278_U195, R2278_U196, R2278_U197, R2278_U198, R2278_U199, R2278_U20, R2278_U200, R2278_U201, R2278_U202, R2278_U203, R2278_U204, R2278_U205, R2278_U206, R2278_U207, R2278_U208, R2278_U209, R2278_U21, R2278_U210, R2278_U211, R2278_U212, R2278_U213, R2278_U214, R2278_U215, R2278_U216, R2278_U217, R2278_U218, R2278_U219, R2278_U22, R2278_U220, R2278_U221, R2278_U222, R2278_U223, R2278_U224, R2278_U225, R2278_U226, R2278_U227, R2278_U228, R2278_U229, R2278_U23, R2278_U230, R2278_U231, R2278_U232, R2278_U233, R2278_U234, R2278_U235, R2278_U236, R2278_U237, R2278_U238, R2278_U239, R2278_U24, R2278_U240, R2278_U241, R2278_U242, R2278_U243, R2278_U244, R2278_U245, R2278_U246, R2278_U247, R2278_U248, R2278_U249, R2278_U25, R2278_U250, R2278_U251, R2278_U252, R2278_U253, R2278_U254, R2278_U255, R2278_U256, R2278_U257, R2278_U258, R2278_U259, R2278_U26, R2278_U260, R2278_U261, R2278_U262, R2278_U263, R2278_U264, R2278_U265, R2278_U266, R2278_U267, R2278_U268, R2278_U269, R2278_U27, R2278_U270, R2278_U271, R2278_U272, R2278_U273, R2278_U274, R2278_U275, R2278_U276, R2278_U277, R2278_U278, R2278_U279, R2278_U28, R2278_U280, R2278_U281, R2278_U282, R2278_U283, R2278_U284, R2278_U285, R2278_U286, R2278_U287, R2278_U288, R2278_U289, R2278_U29, R2278_U290, R2278_U291, R2278_U292, R2278_U293, R2278_U294, R2278_U295, R2278_U296, R2278_U297, R2278_U298, R2278_U299, R2278_U30, R2278_U300, R2278_U301, R2278_U302, R2278_U303, R2278_U304, R2278_U305, R2278_U306, R2278_U307, R2278_U308, R2278_U309, R2278_U31, R2278_U310, R2278_U311, R2278_U312, R2278_U313, R2278_U314, R2278_U315, R2278_U316, R2278_U317, R2278_U318, R2278_U319, R2278_U32, R2278_U320, R2278_U321, R2278_U322, R2278_U323, R2278_U324, R2278_U325, R2278_U326, R2278_U327, R2278_U328, R2278_U329, R2278_U33, R2278_U330, R2278_U331, R2278_U332, R2278_U333, R2278_U334, R2278_U335, R2278_U336, R2278_U337, R2278_U338, R2278_U339, R2278_U34, R2278_U340, R2278_U341, R2278_U342, R2278_U343, R2278_U344, R2278_U345, R2278_U346, R2278_U347, R2278_U348, R2278_U349, R2278_U35, R2278_U350, R2278_U351, R2278_U352, R2278_U353, R2278_U354, R2278_U355, R2278_U356, R2278_U357, R2278_U358, R2278_U359, R2278_U36, R2278_U360, R2278_U361, R2278_U362, R2278_U363, R2278_U364, R2278_U365, R2278_U366, R2278_U367, R2278_U368, R2278_U369, R2278_U37, R2278_U370, R2278_U371, R2278_U372, R2278_U373, R2278_U374, R2278_U375, R2278_U376, R2278_U377, R2278_U378, R2278_U379, R2278_U38, R2278_U380, R2278_U381, R2278_U382, R2278_U383, R2278_U384, R2278_U385, R2278_U386, R2278_U387, R2278_U388, R2278_U389, R2278_U39, R2278_U390, R2278_U391, R2278_U392, R2278_U393, R2278_U394, R2278_U395, R2278_U396, R2278_U397, R2278_U398, R2278_U399, R2278_U40, R2278_U400, R2278_U401, R2278_U402, R2278_U403, R2278_U404, R2278_U405, R2278_U406, R2278_U407, R2278_U408, R2278_U409, R2278_U41, R2278_U410, R2278_U411, R2278_U412, R2278_U413, R2278_U414, R2278_U415, R2278_U416, R2278_U417, R2278_U418, R2278_U419, R2278_U42, R2278_U420, R2278_U421, R2278_U422, R2278_U43, R2278_U44, R2278_U45, R2278_U46, R2278_U47, R2278_U48, R2278_U49, R2278_U5, R2278_U50, R2278_U51, R2278_U52, R2278_U53, R2278_U54, R2278_U55, R2278_U56, R2278_U57, R2278_U58, R2278_U59, R2278_U6, R2278_U60, R2278_U61, R2278_U62, R2278_U63, R2278_U64, R2278_U65, R2278_U66, R2278_U67, R2278_U68, R2278_U69, R2278_U7, R2278_U70, R2278_U71, R2278_U72, R2278_U73, R2278_U74, R2278_U75, R2278_U76, R2278_U77, R2278_U78, R2278_U79, R2278_U8, R2278_U80, R2278_U81, R2278_U82, R2278_U83, R2278_U84, R2278_U85, R2278_U86, R2278_U87, R2278_U88, R2278_U89, R2278_U9, R2278_U90, R2278_U91, R2278_U92, R2278_U93, R2278_U94, R2278_U95, R2278_U96, R2278_U97, R2278_U98, R2278_U99, R2337_U10, R2337_U100, R2337_U101, R2337_U102, R2337_U103, R2337_U104, R2337_U105, R2337_U106, R2337_U107, R2337_U108, R2337_U109, R2337_U11, R2337_U110, R2337_U111, R2337_U112, R2337_U113, R2337_U114, R2337_U115, R2337_U116, R2337_U117, R2337_U118, R2337_U119, R2337_U12, R2337_U120, R2337_U121, R2337_U122, R2337_U123, R2337_U124, R2337_U125, R2337_U126, R2337_U127, R2337_U128, R2337_U129, R2337_U13, R2337_U130, R2337_U131, R2337_U132, R2337_U133, R2337_U134, R2337_U135, R2337_U136, R2337_U137, R2337_U138, R2337_U139, R2337_U14, R2337_U140, R2337_U141, R2337_U142, R2337_U143, R2337_U144, R2337_U145, R2337_U146, R2337_U147, R2337_U148, R2337_U149, R2337_U15, R2337_U150, R2337_U151, R2337_U152, R2337_U153, R2337_U154, R2337_U155, R2337_U156, R2337_U157, R2337_U158, R2337_U159, R2337_U16, R2337_U160, R2337_U161, R2337_U162, R2337_U163, R2337_U164, R2337_U165, R2337_U166, R2337_U167, R2337_U168, R2337_U169, R2337_U17, R2337_U170, R2337_U171, R2337_U172, R2337_U173, R2337_U174, R2337_U175, R2337_U176, R2337_U177, R2337_U178, R2337_U179, R2337_U18, R2337_U180, R2337_U181, R2337_U182, R2337_U183, R2337_U184, R2337_U185, R2337_U186, R2337_U187, R2337_U188, R2337_U189, R2337_U19, R2337_U190, R2337_U191, R2337_U192, R2337_U193, R2337_U20, R2337_U21, R2337_U22, R2337_U23, R2337_U24, R2337_U25, R2337_U26, R2337_U27, R2337_U28, R2337_U29, R2337_U30, R2337_U31, R2337_U32, R2337_U33, R2337_U34, R2337_U35, R2337_U36, R2337_U37, R2337_U38, R2337_U39, R2337_U40, R2337_U41, R2337_U42, R2337_U43, R2337_U44, R2337_U45, R2337_U46, R2337_U47, R2337_U48, R2337_U49, R2337_U5, R2337_U50, R2337_U51, R2337_U52, R2337_U53, R2337_U54, R2337_U55, R2337_U56, R2337_U57, R2337_U58, R2337_U59, R2337_U6, R2337_U60, R2337_U61, R2337_U62, R2337_U63, R2337_U64, R2337_U65, R2337_U66, R2337_U67, R2337_U68, R2337_U69, R2337_U7, R2337_U70, R2337_U71, R2337_U72, R2337_U73, R2337_U74, R2337_U75, R2337_U76, R2337_U77, R2337_U78, R2337_U79, R2337_U8, R2337_U80, R2337_U81, R2337_U82, R2337_U83, R2337_U84, R2337_U85, R2337_U86, R2337_U87, R2337_U88, R2337_U89, R2337_U9, R2337_U90, R2337_U91, R2337_U92, R2337_U93, R2337_U94, R2337_U95, R2337_U96, R2337_U97, R2337_U98, R2337_U99, R2358_U10, R2358_U100, R2358_U101, R2358_U102, R2358_U103, R2358_U104, R2358_U105, R2358_U106, R2358_U107, R2358_U108, R2358_U109, R2358_U11, R2358_U110, R2358_U111, R2358_U112, R2358_U113, R2358_U114, R2358_U115, R2358_U116, R2358_U117, R2358_U118, R2358_U119, R2358_U12, R2358_U120, R2358_U121, R2358_U122, R2358_U123, R2358_U124, R2358_U125, R2358_U126, R2358_U127, R2358_U128, R2358_U129, R2358_U13, R2358_U130, R2358_U131, R2358_U132, R2358_U133, R2358_U134, R2358_U135, R2358_U136, R2358_U137, R2358_U138, R2358_U139, R2358_U14, R2358_U140, R2358_U141, R2358_U142, R2358_U143, R2358_U144, R2358_U145, R2358_U146, R2358_U147, R2358_U148, R2358_U149, R2358_U15, R2358_U150, R2358_U151, R2358_U152, R2358_U153, R2358_U154, R2358_U155, R2358_U156, R2358_U157, R2358_U158, R2358_U159, R2358_U16, R2358_U160, R2358_U161, R2358_U162, R2358_U163, R2358_U164, R2358_U165, R2358_U166, R2358_U167, R2358_U168, R2358_U169, R2358_U17, R2358_U170, R2358_U171, R2358_U172, R2358_U173, R2358_U174, R2358_U175, R2358_U176, R2358_U177, R2358_U178, R2358_U179, R2358_U18, R2358_U180, R2358_U181, R2358_U182, R2358_U183, R2358_U184, R2358_U185, R2358_U186, R2358_U187, R2358_U188, R2358_U189, R2358_U19, R2358_U190, R2358_U191, R2358_U192, R2358_U193, R2358_U194, R2358_U195, R2358_U196, R2358_U197, R2358_U198, R2358_U199, R2358_U20, R2358_U200, R2358_U201, R2358_U202, R2358_U203, R2358_U204, R2358_U205, R2358_U206, R2358_U207, R2358_U208, R2358_U209, R2358_U21, R2358_U210, R2358_U211, R2358_U212, R2358_U213, R2358_U214, R2358_U215, R2358_U216, R2358_U217, R2358_U218, R2358_U219, R2358_U22, R2358_U220, R2358_U221, R2358_U222, R2358_U223, R2358_U224, R2358_U225, R2358_U226, R2358_U227, R2358_U228, R2358_U229, R2358_U23, R2358_U230, R2358_U231, R2358_U232, R2358_U233, R2358_U234, R2358_U235, R2358_U236, R2358_U237, R2358_U238, R2358_U239, R2358_U24, R2358_U240, R2358_U241, R2358_U242, R2358_U243, R2358_U244, R2358_U245, R2358_U246, R2358_U247, R2358_U248, R2358_U249, R2358_U25, R2358_U250, R2358_U251, R2358_U252, R2358_U253, R2358_U254, R2358_U255, R2358_U256, R2358_U257, R2358_U258, R2358_U259, R2358_U26, R2358_U260, R2358_U261, R2358_U262, R2358_U263, R2358_U264, R2358_U265, R2358_U266, R2358_U267, R2358_U268, R2358_U269, R2358_U27, R2358_U270, R2358_U271, R2358_U272, R2358_U273, R2358_U274, R2358_U275, R2358_U276, R2358_U277, R2358_U278, R2358_U279, R2358_U28, R2358_U280, R2358_U281, R2358_U282, R2358_U283, R2358_U284, R2358_U285, R2358_U286, R2358_U287, R2358_U288, R2358_U289, R2358_U29, R2358_U290, R2358_U291, R2358_U292, R2358_U293, R2358_U294, R2358_U295, R2358_U296, R2358_U297, R2358_U298, R2358_U299, R2358_U30, R2358_U300, R2358_U301, R2358_U302, R2358_U303, R2358_U304, R2358_U305, R2358_U306, R2358_U307, R2358_U308, R2358_U309, R2358_U31, R2358_U310, R2358_U311, R2358_U312, R2358_U313, R2358_U314, R2358_U315, R2358_U316, R2358_U317, R2358_U318, R2358_U319, R2358_U32, R2358_U320, R2358_U321, R2358_U322, R2358_U323, R2358_U324, R2358_U325, R2358_U326, R2358_U327, R2358_U328, R2358_U329, R2358_U33, R2358_U330, R2358_U331, R2358_U332, R2358_U333, R2358_U334, R2358_U335, R2358_U336, R2358_U337, R2358_U338, R2358_U339, R2358_U34, R2358_U340, R2358_U341, R2358_U342, R2358_U343, R2358_U344, R2358_U345, R2358_U346, R2358_U347, R2358_U348, R2358_U349, R2358_U35, R2358_U350, R2358_U351, R2358_U352, R2358_U353, R2358_U354, R2358_U355, R2358_U356, R2358_U357, R2358_U358, R2358_U359, R2358_U36, R2358_U360, R2358_U361, R2358_U362, R2358_U363, R2358_U364, R2358_U365, R2358_U366, R2358_U367, R2358_U368, R2358_U369, R2358_U37, R2358_U370, R2358_U371, R2358_U372, R2358_U373, R2358_U374, R2358_U375, R2358_U376, R2358_U377, R2358_U378, R2358_U379, R2358_U38, R2358_U380, R2358_U381, R2358_U382, R2358_U383, R2358_U384, R2358_U385, R2358_U386, R2358_U387, R2358_U388, R2358_U389, R2358_U39, R2358_U390, R2358_U391, R2358_U392, R2358_U393, R2358_U394, R2358_U395, R2358_U396, R2358_U397, R2358_U398, R2358_U399, R2358_U40, R2358_U400, R2358_U401, R2358_U402, R2358_U403, R2358_U404, R2358_U405, R2358_U406, R2358_U407, R2358_U408, R2358_U409, R2358_U41, R2358_U410, R2358_U411, R2358_U412, R2358_U413, R2358_U414, R2358_U415, R2358_U416, R2358_U417, R2358_U418, R2358_U419, R2358_U42, R2358_U420, R2358_U421, R2358_U422, R2358_U423, R2358_U424, R2358_U425, R2358_U426, R2358_U427, R2358_U428, R2358_U429, R2358_U43, R2358_U430, R2358_U431, R2358_U432, R2358_U433, R2358_U434, R2358_U435, R2358_U436, R2358_U437, R2358_U438, R2358_U439, R2358_U44, R2358_U440, R2358_U441, R2358_U442, R2358_U443, R2358_U444, R2358_U445, R2358_U446, R2358_U447, R2358_U448, R2358_U449, R2358_U45, R2358_U450, R2358_U451, R2358_U452, R2358_U453, R2358_U454, R2358_U455, R2358_U456, R2358_U457, R2358_U458, R2358_U459, R2358_U46, R2358_U460, R2358_U461, R2358_U462, R2358_U463, R2358_U464, R2358_U465, R2358_U466, R2358_U467, R2358_U468, R2358_U469, R2358_U47, R2358_U470, R2358_U471, R2358_U472, R2358_U473, R2358_U474, R2358_U475, R2358_U476, R2358_U477, R2358_U478, R2358_U479, R2358_U48, R2358_U480, R2358_U481, R2358_U482, R2358_U483, R2358_U484, R2358_U485, R2358_U486, R2358_U487, R2358_U488, R2358_U489, R2358_U49, R2358_U490, R2358_U491, R2358_U492, R2358_U493, R2358_U494, R2358_U495, R2358_U496, R2358_U497, R2358_U498, R2358_U499, R2358_U5, R2358_U50, R2358_U500, R2358_U501, R2358_U502, R2358_U503, R2358_U504, R2358_U505, R2358_U506, R2358_U507, R2358_U508, R2358_U509, R2358_U51, R2358_U510, R2358_U511, R2358_U512, R2358_U513, R2358_U514, R2358_U515, R2358_U516, R2358_U517, R2358_U518, R2358_U519, R2358_U52, R2358_U520, R2358_U521, R2358_U522, R2358_U523, R2358_U524, R2358_U525, R2358_U526, R2358_U527, R2358_U528, R2358_U529, R2358_U53, R2358_U530, R2358_U531, R2358_U532, R2358_U533, R2358_U534, R2358_U535, R2358_U536, R2358_U537, R2358_U538, R2358_U539, R2358_U54, R2358_U540, R2358_U541, R2358_U542, R2358_U543, R2358_U544, R2358_U545, R2358_U546, R2358_U547, R2358_U548, R2358_U549, R2358_U55, R2358_U550, R2358_U551, R2358_U552, R2358_U553, R2358_U554, R2358_U555, R2358_U556, R2358_U557, R2358_U558, R2358_U559, R2358_U56, R2358_U560, R2358_U561, R2358_U562, R2358_U563, R2358_U564, R2358_U565, R2358_U566, R2358_U567, R2358_U568, R2358_U569, R2358_U57, R2358_U570, R2358_U571, R2358_U572, R2358_U573, R2358_U574, R2358_U575, R2358_U576, R2358_U577, R2358_U578, R2358_U579, R2358_U58, R2358_U580, R2358_U581, R2358_U582, R2358_U583, R2358_U584, R2358_U585, R2358_U586, R2358_U587, R2358_U588, R2358_U589, R2358_U59, R2358_U590, R2358_U591, R2358_U592, R2358_U593, R2358_U594, R2358_U595, R2358_U596, R2358_U597, R2358_U598, R2358_U599, R2358_U6, R2358_U60, R2358_U600, R2358_U601, R2358_U602, R2358_U603, R2358_U604, R2358_U605, R2358_U606, R2358_U607, R2358_U608, R2358_U609, R2358_U61, R2358_U610, R2358_U611, R2358_U612, R2358_U613, R2358_U614, R2358_U615, R2358_U616, R2358_U617, R2358_U618, R2358_U619, R2358_U62, R2358_U620, R2358_U621, R2358_U622, R2358_U623, R2358_U624, R2358_U625, R2358_U626, R2358_U627, R2358_U628, R2358_U629, R2358_U63, R2358_U630, R2358_U631, R2358_U632, R2358_U633, R2358_U634, R2358_U635, R2358_U636, R2358_U637, R2358_U638, R2358_U639, R2358_U64, R2358_U640, R2358_U641, R2358_U642, R2358_U643, R2358_U644, R2358_U645, R2358_U646, R2358_U647, R2358_U648, R2358_U649, R2358_U65, R2358_U650, R2358_U651, R2358_U652, R2358_U653, R2358_U654, R2358_U66, R2358_U67, R2358_U68, R2358_U69, R2358_U7, R2358_U70, R2358_U71, R2358_U72, R2358_U73, R2358_U74, R2358_U75, R2358_U76, R2358_U77, R2358_U78, R2358_U79, R2358_U8, R2358_U80, R2358_U81, R2358_U82, R2358_U83, R2358_U84, R2358_U85, R2358_U86, R2358_U87, R2358_U88, R2358_U89, R2358_U9, R2358_U90, R2358_U91, R2358_U92, R2358_U93, R2358_U94, R2358_U95, R2358_U96, R2358_U97, R2358_U98, R2358_U99, R584_U6, R584_U7, R584_U8, R584_U9, SUB_357_U10, SUB_357_U11, SUB_357_U12, SUB_357_U13, SUB_357_U6, SUB_357_U7, SUB_357_U8, SUB_357_U9, SUB_450_U10, SUB_450_U11, SUB_450_U12, SUB_450_U13, SUB_450_U14, SUB_450_U15, SUB_450_U16, SUB_450_U17, SUB_450_U18, SUB_450_U19, SUB_450_U20, SUB_450_U21, SUB_450_U22, SUB_450_U23, SUB_450_U24, SUB_450_U25, SUB_450_U26, SUB_450_U27, SUB_450_U28, SUB_450_U29, SUB_450_U30, SUB_450_U31, SUB_450_U32, SUB_450_U33, SUB_450_U34, SUB_450_U35, SUB_450_U36, SUB_450_U37, SUB_450_U38, SUB_450_U39, SUB_450_U40, SUB_450_U41, SUB_450_U42, SUB_450_U43, SUB_450_U44, SUB_450_U45, SUB_450_U46, SUB_450_U47, SUB_450_U48, SUB_450_U49, SUB_450_U50, SUB_450_U51, SUB_450_U52, SUB_450_U53, SUB_450_U54, SUB_450_U55, SUB_450_U56, SUB_450_U57, SUB_450_U58, SUB_450_U59, SUB_450_U6, SUB_450_U60, SUB_450_U61, SUB_450_U62, SUB_450_U63, SUB_450_U64, SUB_450_U65, SUB_450_U66, SUB_450_U7, SUB_450_U8, SUB_450_U9, SUB_580_U10, SUB_580_U6, SUB_580_U7, SUB_580_U8, SUB_580_U9, U2352, U2353, U2354, U2355, U2356, U2357, U2358, U2359, U2360, U2361, U2362, U2363, U2364, U2365, U2366, U2367, U2368, U2369, U2370, U2371, U2372, U2373, U2374, U2375, U2376, U2377, U2378, U2379, U2380, U2381, U2382, U2383, U2384, U2385, U2386, U2387, U2388, U2389, U2390, U2391, U2392, U2393, U2394, U2395, U2396, U2397, U2398, U2399, U2400, U2401, U2402, U2403, U2404, U2405, U2406, U2407, U2408, U2409, U2410, U2411, U2412, U2413, U2414, U2415, U2416, U2417, U2418, U2419, U2420, U2421, U2422, U2423, U2424, U2425, U2426, U2427, U2428, U2429, U2430, U2431, U2432, U2433, U2434, U2435, U2436, U2437, U2438, U2439, U2440, U2441, U2442, U2443, U2444, U2445, U2446, U2447, U2448, U2449, U2450, U2451, U2452, U2453, U2454, U2455, U2456, U2457, U2458, U2459, U2460, U2461, U2462, U2463, U2464, U2465, U2466, U2467, U2468, U2469, U2470, U2471, U2472, U2473, U2474, U2475, U2476, U2477, U2478, U2479, U2480, U2481, U2482, U2483, U2484, U2485, U2486, U2487, U2488, U2489, U2490, U2491, U2492, U2493, U2494, U2495, U2496, U2497, U2498, U2499, U2500, U2501, U2502, U2503, U2504, U2505, U2506, U2507, U2508, U2509, U2510, U2511, U2512, U2513, U2514, U2515, U2516, U2517, U2518, U2519, U2520, U2521, U2522, U2523, U2524, U2525, U2526, U2527, U2528, U2529, U2530, U2531, U2532, U2533, U2534, U2535, U2536, U2537, U2538, U2539, U2540, U2541, U2542, U2543, U2544, U2545, U2546, U2547, U2548, U2549, U2550, U2551, U2552, U2553, U2554, U2555, U2556, U2557, U2558, U2559, U2560, U2561, U2562, U2563, U2564, U2565, U2566, U2567, U2568, U2569, U2570, U2571, U2572, U2573, U2574, U2575, U2576, U2577, U2578, U2579, U2580, U2581, U2582, U2583, U2584, U2585, U2586, U2587, U2588, U2589, U2590, U2591, U2592, U2593, U2594, U2595, U2596, U2597, U2598, U2599, U2600, U2601, U2602, U2603, U2604, U2605, U2606, U2607, U2608, U2609, U2610, U2611, U2612, U2613, U2614, U2615, U2616, U2617, U2618, U2620, U2621, U2622, U2623, U2624, U2625, U2626, U2627, U2628, U2629, U2630, U2631, U2632, U2633, U2634, U2635, U2636, U2637, U2638, U2639, U2640, U2641, U2642, U2643, U2644, U2645, U2646, U2647, U2648, U2649, U2650, U2651, U2652, U2653, U2654, U2655, U2656, U2657, U2658, U2659, U2660, U2661, U2662, U2663, U2664, U2665, U2666, U2667, U2668, U2669, U2670, U2671, U2672, U2673, U2674, U2675, U2676, U2677, U2678, U2679, U2680, U2681, U2682, U2683, U2684, U2685, U2686, U2687, U2688, U2689, U2690, U2691, U2692, U2693, U2694, U2695, U2696, U2697, U2698, U2699, U2700, U2701, U2702, U2703, U2704, U2705, U2706, U2707, U2708, U2709, U2710, U2711, U2712, U2713, U2714, U2715, U2716, U2717, U2718, U2719, U2720, U2721, U2722, U2723, U2724, U2725, U2726, U2727, U2728, U2729, U2730, U2731, U2732, U2733, U2734, U2735, U2736, U2737, U2738, U2739, U2740, U2741, U2742, U2743, U2744, U2745, U2746, U2747, U2748, U2749, U2750, U2751, U2752, U2753, U2754, U2755, U2756, U2757, U2758, U2759, U2760, U2761, U2762, U2763, U2764, U2765, U2766, U2767, U2768, U2769, U2770, U2771, U2772, U2773, U2774, U2775, U2776, U2777, U2778, U2779, U2780, U2781, U2782, U2783, U2784, U2785, U2786, U2787, U3214, U3215, U3216, U3217, U3218, U3219, U3220, U3221, U3222, U3223, U3224, U3225, U3226, U3227, U3228, U3229, U3230, U3231, U3232, U3233, U3234, U3235, U3236, U3237, U3238, U3239, U3240, U3241, U3242, U3243, U3244, U3245, U3246, U3247, U3248, U3249, U3250, U3251, U3252, U3253, U3254, U3255, U3256, U3257, U3258, U3259, U3260, U3261, U3262, U3263, U3264, U3265, U3266, U3267, U3268, U3269, U3270, U3271, U3272, U3273, U3274, U3275, U3276, U3277, U3278, U3279, U3280, U3281, U3282, U3283, U3284, U3285, U3286, U3287, U3288, U3289, U3290, U3291, U3292, U3293, U3294, U3295, U3296, U3297, U3298, U3299, U3300, U3301, U3302, U3303, U3304, U3305, U3306, U3307, U3308, U3309, U3310, U3311, U3312, U3313, U3314, U3315, U3316, U3317, U3318, U3319, U3320, U3321, U3322, U3323, U3324, U3325, U3326, U3327, U3328, U3329, U3330, U3331, U3332, U3333, U3334, U3335, U3336, U3337, U3338, U3339, U3340, U3341, U3342, U3343, U3344, U3345, U3346, U3347, U3348, U3349, U3350, U3351, U3352, U3353, U3354, U3355, U3356, U3357, U3358, U3359, U3360, U3361, U3362, U3363, U3364, U3365, U3366, U3367, U3368, U3369, U3370, U3371, U3372, U3373, U3374, U3375, U3376, U3377, U3378, U3379, U3380, U3381, U3382, U3383, U3384, U3385, U3386, U3387, U3388, U3389, U3390, U3391, U3392, U3393, U3394, U3395, U3396, U3397, U3398, U3399, U3400, U3401, U3402, U3403, U3404, U3405, U3406, U3407, U3408, U3409, U3410, U3411, U3412, U3413, U3414, U3415, U3416, U3417, U3418, U3419, U3420, U3421, U3422, U3423, U3424, U3425, U3426, U3427, U3428, U3429, U3430, U3431, U3432, U3433, U3434, U3435, U3436, U3437, U3438, U3439, U3440, U3441, U3442, U3443, U3444, U3449, U3450, U3454, U3457, U3458, U3466, U3467, U3475, U3476, U3477, U3478, U3479, U3480, U3481, U3482, U3483, U3484, U3485, U3486, U3487, U3488, U3489, U3490, U3491, U3492, U3493, U3494, U3495, U3496, U3497, U3498, U3499, U3500, U3501, U3502, U3503, U3504, U3505, U3506, U3507, U3508, U3509, U3510, U3511, U3512, U3513, U3514, U3515, U3516, U3517, U3518, U3519, U3520, U3521, U3522, U3523, U3524, U3525, U3526, U3527, U3528, U3529, U3530, U3531, U3532, U3533, U3534, U3535, U3536, U3537, U3538, U3539, U3540, U3541, U3542, U3543, U3544, U3545, U3546, U3547, U3548, U3549, U3550, U3551, U3552, U3553, U3554, U3555, U3556, U3557, U3558, U3559, U3560, U3561, U3562, U3563, U3564, U3565, U3566, U3567, U3568, U3569, U3570, U3571, U3572, U3573, U3574, U3575, U3576, U3577, U3578, U3579, U3580, U3581, U3582, U3583, U3584, U3585, U3586, U3587, U3588, U3589, U3590, U3591, U3592, U3593, U3594, U3595, U3596, U3597, U3598, U3599, U3600, U3601, U3602, U3603, U3604, U3605, U3606, U3607, U3608, U3609, U3610, U3611, U3612, U3613, U3614, U3615, U3616, U3617, U3618, U3619, U3620, U3621, U3622, U3623, U3624, U3625, U3626, U3627, U3628, U3629, U3630, U3631, U3632, U3633, U3634, U3635, U3636, U3637, U3638, U3639, U3640, U3641, U3642, U3643, U3644, U3645, U3646, U3647, U3648, U3649, U3650, U3651, U3652, U3653, U3654, U3655, U3656, U3657, U3658, U3659, U3660, U3661, U3662, U3663, U3664, U3665, U3666, U3667, U3668, U3669, U3670, U3671, U3672, U3673, U3674, U3675, U3676, U3677, U3678, U3679, U3680, U3681, U3682, U3683, U3684, U3685, U3686, U3687, U3688, U3689, U3690, U3691, U3692, U3693, U3694, U3695, U3696, U3697, U3698, U3699, U3700, U3701, U3702, U3703, U3704, U3705, U3706, U3707, U3708, U3709, U3710, U3711, U3712, U3713, U3714, U3715, U3716, U3717, U3718, U3719, U3720, U3721, U3722, U3723, U3724, U3725, U3726, U3727, U3728, U3729, U3730, U3731, U3732, U3733, U3734, U3735, U3736, U3737, U3738, U3739, U3740, U3741, U3742, U3743, U3744, U3745, U3746, U3747, U3748, U3749, U3750, U3751, U3752, U3753, U3754, U3755, U3756, U3757, U3758, U3759, U3760, U3761, U3762, U3763, U3764, U3765, U3766, U3767, U3768, U3769, U3770, U3771, U3772, U3773, U3774, U3775, U3776, U3777, U3778, U3779, U3780, U3781, U3782, U3783, U3784, U3785, U3786, U3787, U3788, U3789, U3790, U3791, U3792, U3793, U3794, U3795, U3796, U3797, U3798, U3799, U3800, U3801, U3802, U3803, U3804, U3805, U3806, U3807, U3808, U3809, U3810, U3811, U3812, U3813, U3814, U3815, U3816, U3817, U3818, U3819, U3820, U3821, U3822, U3823, U3824, U3825, U3826, U3827, U3828, U3829, U3830, U3831, U3832, U3833, U3834, U3835, U3836, U3837, U3838, U3839, U3840, U3841, U3842, U3843, U3844, U3845, U3846, U3847, U3848, U3849, U3850, U3851, U3852, U3853, U3854, U3855, U3856, U3857, U3858, U3859, U3860, U3861, U3862, U3863, U3864, U3865, U3866, U3867, U3868, U3869, U3870, U3871, U3872, U3873, U3874, U3875, U3876, U3877, U3878, U3879, U3880, U3881, U3882, U3883, U3884, U3885, U3886, U3887, U3888, U3889, U3890, U3891, U3892, U3893, U3894, U3895, U3896, U3897, U3898, U3899, U3900, U3901, U3902, U3903, U3904, U3905, U3906, U3907, U3908, U3909, U3910, U3911, U3912, U3913, U3914, U3915, U3916, U3917, U3918, U3919, U3920, U3921, U3922, U3923, U3924, U3925, U3926, U3927, U3928, U3929, U3930, U3931, U3932, U3933, U3934, U3935, U3936, U3937, U3938, U3939, U3940, U3941, U3942, U3943, U3944, U3945, U3946, U3947, U3948, U3949, U3950, U3951, U3952, U3953, U3954, U3955, U3956, U3957, U3958, U3959, U3960, U3961, U3962, U3963, U3964, U3965, U3966, U3967, U3968, U3969, U3970, U3971, U3972, U3973, U3974, U3975, U3976, U3977, U3978, U3979, U3980, U3981, U3982, U3983, U3984, U3985, U3986, U3987, U3988, U3989, U3990, U3991, U3992, U3993, U3994, U3995, U3996, U3997, U3998, U3999, U4000, U4001, U4002, U4003, U4004, U4005, U4006, U4007, U4008, U4009, U4010, U4011, U4012, U4013, U4014, U4015, U4016, U4017, U4018, U4019, U4020, U4021, U4022, U4023, U4024, U4025, U4026, U4027, U4028, U4029, U4030, U4031, U4032, U4033, U4034, U4035, U4036, U4037, U4038, U4039, U4040, U4041, U4042, U4043, U4044, U4045, U4046, U4047, U4048, U4049, U4050, U4051, U4052, U4053, U4054, U4055, U4056, U4057, U4058, U4059, U4060, U4061, U4062, U4063, U4064, U4065, U4066, U4067, U4068, U4069, U4070, U4071, U4072, U4073, U4074, U4075, U4076, U4077, U4078, U4079, U4080, U4081, U4082, U4083, U4084, U4085, U4086, U4087, U4088, U4089, U4090, U4091, U4092, U4093, U4094, U4095, U4096, U4097, U4098, U4099, U4100, U4101, U4102, U4103, U4104, U4105, U4106, U4107, U4108, U4109, U4110, U4111, U4112, U4113, U4114, U4115, U4116, U4117, U4118, U4119, U4120, U4121, U4122, U4123, U4124, U4125, U4126, U4127, U4128, U4129, U4130, U4131, U4132, U4133, U4134, U4135, U4136, U4137, U4138, U4139, U4140, U4141, U4142, U4143, U4144, U4145, U4146, U4147, U4148, U4149, U4150, U4151, U4152, U4153, U4154, U4155, U4156, U4157, U4158, U4159, U4160, U4161, U4162, U4163, U4164, U4165, U4166, U4167, U4168, U4169, U4170, U4171, U4172, U4173, U4174, U4175, U4176, U4177, U4178, U4179, U4180, U4181, U4182, U4183, U4184, U4185, U4186, U4187, U4188, U4189, U4190, U4191, U4192, U4193, U4194, U4195, U4196, U4197, U4198, U4199, U4200, U4201, U4202, U4203, U4204, U4205, U4206, U4207, U4208, U4209, U4210, U4211, U4212, U4213, U4214, U4215, U4216, U4217, U4218, U4219, U4220, U4221, U4222, U4223, U4224, U4225, U4226, U4227, U4228, U4229, U4230, U4231, U4232, U4233, U4234, U4235, U4236, U4237, U4238, U4239, U4240, U4241, U4242, U4243, U4244, U4245, U4246, U4247, U4248, U4249, U4250, U4251, U4252, U4253, U4254, U4255, U4256, U4257, U4258, U4259, U4260, U4261, U4262, U4263, U4264, U4265, U4266, U4267, U4268, U4269, U4270, U4271, U4272, U4273, U4274, U4275, U4276, U4277, U4278, U4279, U4280, U4281, U4282, U4283, U4284, U4285, U4286, U4287, U4288, U4289, U4290, U4291, U4292, U4293, U4294, U4295, U4296, U4297, U4298, U4299, U4300, U4301, U4302, U4303, U4304, U4305, U4306, U4307, U4308, U4309, U4310, U4311, U4312, U4313, U4314, U4315, U4316, U4317, U4318, U4319, U4320, U4321, U4322, U4323, U4324, U4325, U4326, U4327, U4328, U4329, U4330, U4331, U4332, U4333, U4334, U4335, U4336, U4337, U4338, U4339, U4340, U4341, U4342, U4343, U4344, U4345, U4346, U4347, U4348, U4349, U4350, U4351, U4352, U4353, U4354, U4355, U4356, U4357, U4358, U4359, U4360, U4361, U4362, U4363, U4364, U4365, U4366, U4367, U4368, U4369, U4370, U4371, U4372, U4373, U4374, U4375, U4376, U4377, U4378, U4379, U4380, U4381, U4382, U4383, U4384, U4385, U4386, U4387, U4388, U4389, U4390, U4391, U4392, U4393, U4394, U4395, U4396, U4397, U4398, U4399, U4400, U4401, U4402, U4403, U4404, U4405, U4406, U4407, U4408, U4409, U4410, U4411, U4412, U4413, U4414, U4415, U4416, U4417, U4418, U4419, U4420, U4421, U4422, U4423, U4424, U4425, U4426, U4427, U4428, U4429, U4430, U4431, U4432, U4433, U4434, U4435, U4436, U4437, U4438, U4439, U4440, U4441, U4442, U4443, U4444, U4445, U4446, U4447, U4448, U4449, U4450, U4451, U4452, U4453, U4454, U4455, U4456, U4457, U4458, U4459, U4460, U4461, U4462, U4463, U4464, U4465, U4466, U4467, U4468, U4469, U4470, U4471, U4472, U4473, U4474, U4475, U4476, U4477, U4478, U4479, U4480, U4481, U4482, U4483, U4484, U4485, U4486, U4487, U4488, U4489, U4490, U4491, U4492, U4493, U4494, U4495, U4496, U4497, U4498, U4499, U4500, U4501, U4502, U4503, U4504, U4505, U4506, U4507, U4508, U4509, U4510, U4511, U4512, U4513, U4514, U4515, U4516, U4517, U4518, U4519, U4520, U4521, U4522, U4523, U4524, U4525, U4526, U4527, U4528, U4529, U4530, U4531, U4532, U4533, U4534, U4535, U4536, U4537, U4538, U4539, U4540, U4541, U4542, U4543, U4544, U4545, U4546, U4547, U4548, U4549, U4550, U4551, U4552, U4553, U4554, U4555, U4556, U4557, U4558, U4559, U4560, U4561, U4562, U4563, U4564, U4565, U4566, U4567, U4568, U4569, U4570, U4571, U4572, U4573, U4574, U4575, U4576, U4577, U4578, U4579, U4580, U4581, U4582, U4583, U4584, U4585, U4586, U4587, U4588, U4589, U4590, U4591, U4592, U4593, U4594, U4595, U4596, U4597, U4598, U4599, U4600, U4601, U4602, U4603, U4604, U4605, U4606, U4607, U4608, U4609, U4610, U4611, U4612, U4613, U4614, U4615, U4616, U4617, U4618, U4619, U4620, U4621, U4622, U4623, U4624, U4625, U4626, U4627, U4628, U4629, U4630, U4631, U4632, U4633, U4634, U4635, U4636, U4637, U4638, U4639, U4640, U4641, U4642, U4643, U4644, U4645, U4646, U4647, U4648, U4649, U4650, U4651, U4652, U4653, U4654, U4655, U4656, U4657, U4658, U4659, U4660, U4661, U4662, U4663, U4664, U4665, U4666, U4667, U4668, U4669, U4670, U4671, U4672, U4673, U4674, U4675, U4676, U4677, U4678, U4679, U4680, U4681, U4682, U4683, U4684, U4685, U4686, U4687, U4688, U4689, U4690, U4691, U4692, U4693, U4694, U4695, U4696, U4697, U4698, U4699, U4700, U4701, U4702, U4703, U4704, U4705, U4706, U4707, U4708, U4709, U4710, U4711, U4712, U4713, U4714, U4715, U4716, U4717, U4718, U4719, U4720, U4721, U4722, U4723, U4724, U4725, U4726, U4727, U4728, U4729, U4730, U4731, U4732, U4733, U4734, U4735, U4736, U4737, U4738, U4739, U4740, U4741, U4742, U4743, U4744, U4745, U4746, U4747, U4748, U4749, U4750, U4751, U4752, U4753, U4754, U4755, U4756, U4757, U4758, U4759, U4760, U4761, U4762, U4763, U4764, U4765, U4766, U4767, U4768, U4769, U4770, U4771, U4772, U4773, U4774, U4775, U4776, U4777, U4778, U4779, U4780, U4781, U4782, U4783, U4784, U4785, U4786, U4787, U4788, U4789, U4790, U4791, U4792, U4793, U4794, U4795, U4796, U4797, U4798, U4799, U4800, U4801, U4802, U4803, U4804, U4805, U4806, U4807, U4808, U4809, U4810, U4811, U4812, U4813, U4814, U4815, U4816, U4817, U4818, U4819, U4820, U4821, U4822, U4823, U4824, U4825, U4826, U4827, U4828, U4829, U4830, U4831, U4832, U4833, U4834, U4835, U4836, U4837, U4838, U4839, U4840, U4841, U4842, U4843, U4844, U4845, U4846, U4847, U4848, U4849, U4850, U4851, U4852, U4853, U4854, U4855, U4856, U4857, U4858, U4859, U4860, U4861, U4862, U4863, U4864, U4865, U4866, U4867, U4868, U4869, U4870, U4871, U4872, U4873, U4874, U4875, U4876, U4877, U4878, U4879, U4880, U4881, U4882, U4883, U4884, U4885, U4886, U4887, U4888, U4889, U4890, U4891, U4892, U4893, U4894, U4895, U4896, U4897, U4898, U4899, U4900, U4901, U4902, U4903, U4904, U4905, U4906, U4907, U4908, U4909, U4910, U4911, U4912, U4913, U4914, U4915, U4916, U4917, U4918, U4919, U4920, U4921, U4922, U4923, U4924, U4925, U4926, U4927, U4928, U4929, U4930, U4931, U4932, U4933, U4934, U4935, U4936, U4937, U4938, U4939, U4940, U4941, U4942, U4943, U4944, U4945, U4946, U4947, U4948, U4949, U4950, U4951, U4952, U4953, U4954, U4955, U4956, U4957, U4958, U4959, U4960, U4961, U4962, U4963, U4964, U4965, U4966, U4967, U4968, U4969, U4970, U4971, U4972, U4973, U4974, U4975, U4976, U4977, U4978, U4979, U4980, U4981, U4982, U4983, U4984, U4985, U4986, U4987, U4988, U4989, U4990, U4991, U4992, U4993, U4994, U4995, U4996, U4997, U4998, U4999, U5000, U5001, U5002, U5003, U5004, U5005, U5006, U5007, U5008, U5009, U5010, U5011, U5012, U5013, U5014, U5015, U5016, U5017, U5018, U5019, U5020, U5021, U5022, U5023, U5024, U5025, U5026, U5027, U5028, U5029, U5030, U5031, U5032, U5033, U5034, U5035, U5036, U5037, U5038, U5039, U5040, U5041, U5042, U5043, U5044, U5045, U5046, U5047, U5048, U5049, U5050, U5051, U5052, U5053, U5054, U5055, U5056, U5057, U5058, U5059, U5060, U5061, U5062, U5063, U5064, U5065, U5066, U5067, U5068, U5069, U5070, U5071, U5072, U5073, U5074, U5075, U5076, U5077, U5078, U5079, U5080, U5081, U5082, U5083, U5084, U5085, U5086, U5087, U5088, U5089, U5090, U5091, U5092, U5093, U5094, U5095, U5096, U5097, U5098, U5099, U5100, U5101, U5102, U5103, U5104, U5105, U5106, U5107, U5108, U5109, U5110, U5111, U5112, U5113, U5114, U5115, U5116, U5117, U5118, U5119, U5120, U5121, U5122, U5123, U5124, U5125, U5126, U5127, U5128, U5129, U5130, U5131, U5132, U5133, U5134, U5135, U5136, U5137, U5138, U5139, U5140, U5141, U5142, U5143, U5144, U5145, U5146, U5147, U5148, U5149, U5150, U5151, U5152, U5153, U5154, U5155, U5156, U5157, U5158, U5159, U5160, U5161, U5162, U5163, U5164, U5165, U5166, U5167, U5168, U5169, U5170, U5171, U5172, U5173, U5174, U5175, U5176, U5177, U5178, U5179, U5180, U5181, U5182, U5183, U5184, U5185, U5186, U5187, U5188, U5189, U5190, U5191, U5192, U5193, U5194, U5195, U5196, U5197, U5198, U5199, U5200, U5201, U5202, U5203, U5204, U5205, U5206, U5207, U5208, U5209, U5210, U5211, U5212, U5213, U5214, U5215, U5216, U5217, U5218, U5219, U5220, U5221, U5222, U5223, U5224, U5225, U5226, U5227, U5228, U5229, U5230, U5231, U5232, U5233, U5234, U5235, U5236, U5237, U5238, U5239, U5240, U5241, U5242, U5243, U5244, U5245, U5246, U5247, U5248, U5249, U5250, U5251, U5252, U5253, U5254, U5255, U5256, U5257, U5258, U5259, U5260, U5261, U5262, U5263, U5264, U5265, U5266, U5267, U5268, U5269, U5270, U5271, U5272, U5273, U5274, U5275, U5276, U5277, U5278, U5279, U5280, U5281, U5282, U5283, U5284, U5285, U5286, U5287, U5288, U5289, U5290, U5291, U5292, U5293, U5294, U5295, U5296, U5297, U5298, U5299, U5300, U5301, U5302, U5303, U5304, U5305, U5306, U5307, U5308, U5309, U5310, U5311, U5312, U5313, U5314, U5315, U5316, U5317, U5318, U5319, U5320, U5321, U5322, U5323, U5324, U5325, U5326, U5327, U5328, U5329, U5330, U5331, U5332, U5333, U5334, U5335, U5336, U5337, U5338, U5339, U5340, U5341, U5342, U5343, U5344, U5345, U5346, U5347, U5348, U5349, U5350, U5351, U5352, U5353, U5354, U5355, U5356, U5357, U5358, U5359, U5360, U5361, U5362, U5363, U5364, U5365, U5366, U5367, U5368, U5369, U5370, U5371, U5372, U5373, U5374, U5375, U5376, U5377, U5378, U5379, U5380, U5381, U5382, U5383, U5384, U5385, U5386, U5387, U5388, U5389, U5390, U5391, U5392, U5393, U5394, U5395, U5396, U5397, U5398, U5399, U5400, U5401, U5402, U5403, U5404, U5405, U5406, U5407, U5408, U5409, U5410, U5411, U5412, U5413, U5414, U5415, U5416, U5417, U5418, U5419, U5420, U5421, U5422, U5423, U5424, U5425, U5426, U5427, U5428, U5429, U5430, U5431, U5432, U5433, U5434, U5435, U5436, U5437, U5438, U5439, U5440, U5441, U5442, U5443, U5444, U5445, U5446, U5447, U5448, U5449, U5450, U5451, U5452, U5453, U5454, U5455, U5456, U5457, U5458, U5459, U5460, U5461, U5462, U5463, U5464, U5465, U5466, U5467, U5468, U5469, U5470, U5471, U5472, U5473, U5474, U5475, U5476, U5477, U5478, U5479, U5480, U5481, U5482, U5483, U5484, U5485, U5486, U5487, U5488, U5489, U5490, U5491, U5492, U5493, U5494, U5495, U5496, U5497, U5498, U5499, U5500, U5501, U5502, U5503, U5504, U5505, U5506, U5507, U5508, U5509, U5510, U5511, U5512, U5513, U5514, U5515, U5516, U5517, U5518, U5519, U5520, U5521, U5522, U5523, U5524, U5525, U5526, U5527, U5528, U5529, U5530, U5531, U5532, U5533, U5534, U5535, U5536, U5537, U5538, U5539, U5540, U5541, U5542, U5543, U5544, U5545, U5546, U5547, U5548, U5549, U5550, U5551, U5552, U5553, U5554, U5555, U5556, U5557, U5558, U5559, U5560, U5561, U5562, U5563, U5564, U5565, U5566, U5567, U5568, U5569, U5570, U5571, U5572, U5573, U5574, U5575, U5576, U5577, U5578, U5579, U5580, U5581, U5582, U5583, U5584, U5585, U5586, U5587, U5588, U5589, U5590, U5591, U5592, U5593, U5594, U5595, U5596, U5597, U5598, U5599, U5600, U5601, U5602, U5603, U5604, U5605, U5606, U5607, U5608, U5609, U5610, U5611, U5612, U5613, U5614, U5615, U5616, U5617, U5618, U5619, U5620, U5621, U5622, U5623, U5624, U5625, U5626, U5627, U5628, U5629, U5630, U5631, U5632, U5633, U5634, U5635, U5636, U5637, U5638, U5639, U5640, U5641, U5642, U5643, U5644, U5645, U5646, U5647, U5648, U5649, U5650, U5651, U5652, U5653, U5654, U5655, U5656, U5657, U5658, U5659, U5660, U5661, U5662, U5663, U5664, U5665, U5666, U5667, U5668, U5669, U5670, U5671, U5672, U5673, U5674, U5675, U5676, U5677, U5678, U5679, U5680, U5681, U5682, U5683, U5684, U5685, U5686, U5687, U5688, U5689, U5690, U5691, U5692, U5693, U5694, U5695, U5696, U5697, U5698, U5699, U5700, U5701, U5702, U5703, U5704, U5705, U5706, U5707, U5708, U5709, U5710, U5711, U5712, U5713, U5714, U5715, U5716, U5717, U5718, U5719, U5720, U5721, U5722, U5723, U5724, U5725, U5726, U5727, U5728, U5729, U5730, U5731, U5732, U5733, U5734, U5735, U5736, U5737, U5738, U5739, U5740, U5741, U5742, U5743, U5744, U5745, U5746, U5747, U5748, U5749, U5750, U5751, U5752, U5753, U5754, U5755, U5756, U5757, U5758, U5759, U5760, U5761, U5762, U5763, U5764, U5765, U5766, U5767, U5768, U5769, U5770, U5771, U5772, U5773, U5774, U5775, U5776, U5777, U5778, U5779, U5780, U5781, U5782, U5783, U5784, U5785, U5786, U5787, U5788, U5789, U5790, U5791, U5792, U5793, U5794, U5795, U5796, U5797, U5798, U5799, U5800, U5801, U5802, U5803, U5804, U5805, U5806, U5807, U5808, U5809, U5810, U5811, U5812, U5813, U5814, U5815, U5816, U5817, U5818, U5819, U5820, U5821, U5822, U5823, U5824, U5825, U5826, U5827, U5828, U5829, U5830, U5831, U5832, U5833, U5834, U5835, U5836, U5837, U5838, U5839, U5840, U5841, U5842, U5843, U5844, U5845, U5846, U5847, U5848, U5849, U5850, U5851, U5852, U5853, U5854, U5855, U5856, U5857, U5858, U5859, U5860, U5861, U5862, U5863, U5864, U5865, U5866, U5867, U5868, U5869, U5870, U5871, U5872, U5873, U5874, U5875, U5876, U5877, U5878, U5879, U5880, U5881, U5882, U5883, U5884, U5885, U5886, U5887, U5888, U5889, U5890, U5891, U5892, U5893, U5894, U5895, U5896, U5897, U5898, U5899, U5900, U5901, U5902, U5903, U5904, U5905, U5906, U5907, U5908, U5909, U5910, U5911, U5912, U5913, U5914, U5915, U5916, U5917, U5918, U5919, U5920, U5921, U5922, U5923, U5924, U5925, U5926, U5927, U5928, U5929, U5930, U5931, U5932, U5933, U5934, U5935, U5936, U5937, U5938, U5939, U5940, U5941, U5942, U5943, U5944, U5945, U5946, U5947, U5948, U5949, U5950, U5951, U5952, U5953, U5954, U5955, U5956, U5957, U5958, U5959, U5960, U5961, U5962, U5963, U5964, U5965, U5966, U5967, U5968, U5969, U5970, U5971, U5972, U5973, U5974, U5975, U5976, U5977, U5978, U5979, U5980, U5981, U5982, U5983, U5984, U5985, U5986, U5987, U5988, U5989, U5990, U5991, U5992, U5993, U5994, U5995, U5996, U5997, U5998, U5999, U6000, U6001, U6002, U6003, U6004, U6005, U6006, U6007, U6008, U6009, U6010, U6011, U6012, U6013, U6014, U6015, U6016, U6017, U6018, U6019, U6020, U6021, U6022, U6023, U6024, U6025, U6026, U6027, U6028, U6029, U6030, U6031, U6032, U6033, U6034, U6035, U6036, U6037, U6038, U6039, U6040, U6041, U6042, U6043, U6044, U6045, U6046, U6047, U6048, U6049, U6050, U6051, U6052, U6053, U6054, U6055, U6056, U6057, U6058, U6059, U6060, U6061, U6062, U6063, U6064, U6065, U6066, U6067, U6068, U6069, U6070, U6071, U6072, U6073, U6074, U6075, U6076, U6077, U6078, U6079, U6080, U6081, U6082, U6083, U6084, U6085, U6086, U6087, U6088, U6089, U6090, U6091, U6092, U6093, U6094, U6095, U6096, U6097, U6098, U6099, U6100, U6101, U6102, U6103, U6104, U6105, U6106, U6107, U6108, U6109, U6110, U6111, U6112, U6113, U6114, U6115, U6116, U6117, U6118, U6119, U6120, U6121, U6122, U6123, U6124, U6125, U6126, U6127, U6128, U6129, U6130, U6131, U6132, U6133, U6134, U6135, U6136, U6137, U6138, U6139, U6140, U6141, U6142, U6143, U6144, U6145, U6146, U6147, U6148, U6149, U6150, U6151, U6152, U6153, U6154, U6155, U6156, U6157, U6158, U6159, U6160, U6161, U6162, U6163, U6164, U6165, U6166, U6167, U6168, U6169, U6170, U6171, U6172, U6173, U6174, U6175, U6176, U6177, U6178, U6179, U6180, U6181, U6182, U6183, U6184, U6185, U6186, U6187, U6188, U6189, U6190, U6191, U6192, U6193, U6194, U6195, U6196, U6197, U6198, U6199, U6200, U6201, U6202, U6203, U6204, U6205, U6206, U6207, U6208, U6209, U6210, U6211, U6212, U6213, U6214, U6215, U6216, U6217, U6218, U6219, U6220, U6221, U6222, U6223, U6224, U6225, U6226, U6227, U6228, U6229, U6230, U6231, U6232, U6233, U6234, U6235, U6236, U6237, U6238, U6239, U6240, U6241, U6242, U6243, U6244, U6245, U6246, U6247, U6248, U6249, U6250, U6251, U6252, U6253, U6254, U6255, U6256, U6257, U6258, U6259, U6260, U6261, U6262, U6263, U6264, U6265, U6266, U6267, U6268, U6269, U6270, U6271, U6272, U6273, U6274, U6275, U6276, U6277, U6278, U6279, U6280, U6281, U6282, U6283, U6284, U6285, U6286, U6287, U6288, U6289, U6290, U6291, U6292, U6293, U6294, U6295, U6296, U6297, U6298, U6299, U6300, U6301, U6302, U6303, U6304, U6305, U6306, U6307, U6308, U6309, U6310, U6311, U6312, U6313, U6314, U6315, U6316, U6317, U6318, U6319, U6320, U6321, U6322, U6323, U6324, U6325, U6326, U6327, U6328, U6329, U6330, U6331, U6332, U6333, U6334, U6335, U6336, U6337, U6338, U6339, U6340, U6341, U6342, U6343, U6344, U6345, U6346, U6347, U6348, U6349, U6350, U6351, U6352, U6353, U6354, U6355, U6356, U6357, U6358, U6359, U6360, U6361, U6362, U6363, U6364, U6365, U6366, U6367, U6368, U6369, U6370, U6371, U6372, U6373, U6374, U6375, U6376, U6377, U6378, U6379, U6380, U6381, U6382, U6383, U6384, U6385, U6386, U6387, U6388, U6389, U6390, U6391, U6392, U6393, U6394, U6395, U6396, U6397, U6398, U6399, U6400, U6401, U6402, U6403, U6404, U6405, U6406, U6407, U6408, U6409, U6410, U6411, U6412, U6413, U6414, U6415, U6416, U6417, U6418, U6419, U6420, U6421, U6422, U6423, U6424, U6425, U6426, U6427, U6428, U6429, U6430, U6431, U6432, U6433, U6434, U6435, U6436, U6437, U6438, U6439, U6440, U6441, U6442, U6443, U6444, U6445, U6446, U6447, U6448, U6449, U6450, U6451, U6452, U6453, U6454, U6455, U6456, U6457, U6458, U6459, U6460, U6461, U6462, U6463, U6464, U6465, U6466, U6467, U6468, U6469, U6470, U6471, U6472, U6473, U6474, U6475, U6476, U6477, U6478, U6479, U6480, U6481, U6482, U6483, U6484, U6485, U6486, U6487, U6488, U6489, U6490, U6491, U6492, U6493, U6494, U6495, U6496, U6497, U6498, U6499, U6500, U6501, U6502, U6503, U6504, U6505, U6506, U6507, U6508, U6509, U6510, U6511, U6512, U6513, U6514, U6515, U6516, U6517, U6518, U6519, U6520, U6521, U6522, U6523, U6524, U6525, U6526, U6527, U6528, U6529, U6530, U6531, U6532, U6533, U6534, U6535, U6536, U6537, U6538, U6539, U6540, U6541, U6542, U6543, U6544, U6545, U6546, U6547, U6548, U6549, U6550, U6551, U6552, U6553, U6554, U6555, U6556, U6557, U6558, U6559, U6560, U6561, U6562, U6563, U6564, U6565, U6566, U6567, U6568, U6569, U6570, U6571, U6572, U6573, U6574, U6575, U6576, U6577, U6578, U6579, U6580, U6581, U6582, U6583, U6584, U6585, U6586, U6587, U6588, U6589, U6590, U6591, U6592, U6593, U6594, U6595, U6596, U6597, U6598, U6599, U6600, U6601, U6602, U6603, U6604, U6605, U6606, U6607, U6608, U6609, U6610, U6611, U6612, U6613, U6614, U6615, U6616, U6617, U6618, U6619, U6620, U6621, U6622, U6623, U6624, U6625, U6626, U6627, U6628, U6629, U6630, U6631, U6632, U6633, U6634, U6635, U6636, U6637, U6638, U6639, U6640, U6641, U6642, U6643, U6644, U6645, U6646, U6647, U6648, U6649, U6650, U6651, U6652, U6653, U6654, U6655, U6656, U6657, U6658, U6659, U6660, U6661, U6662, U6663, U6664, U6665, U6666, U6667, U6668, U6669, U6670, U6671, U6672, U6673, U6674, U6675, U6676, U6677, U6678, U6679, U6680, U6681, U6682, U6683, U6684, U6685, U6686, U6687, U6688, U6689, U6690, U6691, U6692, U6693, U6694, U6695, U6696, U6697, U6698, U6699, U6700, U6701, U6702, U6703, U6704, U6705, U6706, U6707, U6708, U6709, U6710, U6711, U6712, U6713, U6714, U6715, U6716, U6717, U6718, U6719, U6720, U6721, U6722, U6723, U6724, U6725, U6726, U6727, U6728, U6729, U6730, U6731, U6732, U6733, U6734, U6735, U6736, U6737, U6738, U6739, U6740, U6741, U6742, U6743, U6744, U6745, U6746, U6747, U6748, U6749, U6750, U6751, U6752, U6753, U6754, U6755, U6756, U6757, U6758, U6759, U6760, U6761, U6762, U6763, U6764, U6765, U6766, U6767, U6768, U6769, U6770, U6771, U6772, U6773, U6774, U6775, U6776, U6777, U6778, U6779, U6780, U6781, U6782, U6783, U6784, U6785, U6786, U6787, U6788, U6789, U6790, U6791, U6792, U6793, U6794, U6795, U6796, U6797, U6798, U6799, U6800, U6801, U6802, U6803, U6804, U6805, U6806, U6807, U6808, U6809, U6810, U6811, U6812, U6813, U6814, U6815, U6816, U6817, U6818, U6819, U6820, U6821, U6822, U6823, U6824, U6825, U6826, U6827, U6828, U6829, U6830, U6831, U6832, U6833, U6834, U6835, U6836, U6837, U6838, U6839, U6840, U6841, U6842, U6843, U6844, U6845, U6846, U6847, U6848, U6849, U6850, U6851, U6852, U6853, U6854, U6855, U6856, U6857, U6858, U6859, U6860, U6861, U6862, U6863, U6864, U6865, U6866, U6867, U6868, U6869, U6870, U6871, U6872, U6873, U6874, U6875, U6876, U6877, U6878, U6879, U6880, U6881, U6882, U6883, U6884, U6885, U6886, U6887, U6888, U6889, U6890, U6891, U6892, U6893, U6894, U6895, U6896, U6897, U6898, U6899, U6900, U6901, U6902, U6903, U6904, U6905, U6906, U6907, U6908, U6909, U6910, U6911, U6912, U6913, U6914, U6915, U6916, U6917, U6918, U6919, U6920, U6921, U6922, U6923, U6924, U6925, U6926, U6927, U6928, U6929, U6930, U6931, U6932, U6933, U6934, U6935, U6936, U6937, U6938, U6939, U6940, U6941, U6942, U6943, U6944, U6945, U6946, U6947, U6948, U6949, U6950, U6951, U6952, U6953, U6954, U6955, U6956, U6957, U6958, U6959, U6960, U6961, U6962, U6963, U6964, U6965, U6966, U6967, U6968, U6969, U6970, U6971, U6972, U6973, U6974, U6975, U6976, U6977, U6978, U6979, U6980, U6981, U6982, U6983, U6984, U6985, U6986, U6987, U6988, U6989, U6990, U6991, U6992, U6993, U6994, U6995, U6996, U6997, U6998, U6999, U7000, U7001, U7002, U7003, U7004, U7005, U7006, U7007, U7008, U7009, U7010, U7011, U7012, U7013, U7014, U7015, U7016, U7017, U7018, U7019, U7020, U7021, U7022, U7023, U7024, U7025, U7026, U7027, U7028, U7029, U7030, U7031, U7032, U7033, U7034, U7035, U7036, U7037, U7038, U7039, U7040, U7041, U7042, U7043, U7044, U7045, U7046, U7047, U7048, U7049, U7050, U7051, U7052, U7053, U7054, U7055, U7056, U7057, U7058, U7059, U7060, U7061, U7062, U7063, U7064, U7065, U7066, U7067, U7068, U7069, U7070, U7071, U7072, U7073, U7074, U7075, U7076, U7077, U7078, U7079, U7080, U7081, U7082, U7083, U7084, U7085, U7086, U7087, U7088, U7089, U7090, U7091, U7092, U7093, U7094, U7095, U7096, U7097, U7098, U7099, U7100, U7101, U7102, U7103, U7104, U7105, U7106, U7107, U7108, U7109, U7110, U7111, U7112, U7113, U7114, U7115, U7116, U7117, U7118, U7119, U7120, U7121, U7122, U7123, U7124, U7125, U7126, U7127, U7128, U7129, U7130, U7131, U7132, U7133, U7134, U7135, U7136, U7137, U7138, U7139, U7140, U7141, U7142, U7143, U7144, U7145, U7146, U7147, U7148, U7149, U7150, U7151, U7152, U7153, U7154, U7155, U7156, U7157, U7158, U7159, U7160, U7161, U7162, U7163, U7164, U7165, U7166, U7167, U7168, U7169, U7170, U7171, U7172, U7173, U7174, U7175, U7176, U7177, U7178, U7179, U7180, U7181, U7182, U7183, U7184, U7185, U7186, U7187, U7188, U7189, U7190, U7191, U7192, U7193, U7194, U7195, U7196, U7197, U7198, U7199, U7200, U7201, U7202, U7203, U7204, U7205, U7206, U7207, U7208, U7209, U7210, U7211, U7212, U7213, U7214, U7215, U7216, U7217, U7218, U7219, U7220, U7221, U7222, U7223, U7224, U7225, U7226, U7227, U7228, U7229, U7230, U7231, U7232, U7233, U7234, U7235, U7236, U7237, U7238, U7239, U7240, U7241, U7242, U7243, U7244, U7245, U7246, U7247, U7248, U7249, U7250, U7251, U7252, U7253, U7254, U7255, U7256, U7257, U7258, U7259, U7260, U7261, U7262, U7263, U7264, U7265, U7266, U7267, U7268, U7269, U7270, U7271, U7272, U7273, U7274, U7275, U7276, U7277, U7278, U7279, U7280, U7281, U7282, U7283, U7284, U7285, U7286, U7287, U7288, U7289, U7290, U7291, U7292, U7293, U7294, U7295, U7296, U7297, U7298, U7299, U7300, U7301, U7302, U7303, U7304, U7305, U7306, U7307, U7308, U7309, U7310, U7311, U7312, U7313, U7314, U7315, U7316, U7317, U7318, U7319, U7320, U7321, U7322, U7323, U7324, U7325, U7326, U7327, U7328, U7329, U7330, U7331, U7332, U7333, U7334, U7335, U7336, U7337, U7338, U7339, U7340, U7341, U7342, U7343, U7344, U7345, U7346, U7347, U7348, U7349, U7350, U7351, U7352, U7353, U7354, U7355, U7356, U7357, U7358, U7359, U7360, U7361, U7362, U7363, U7364, U7365, U7366, U7367, U7368, U7369, U7370, U7371, U7372, U7373, U7374, U7375, U7376, U7377, U7378, U7379, U7380, U7381, U7382, U7383, U7384, U7385, U7386, U7387, U7388, U7389, U7390, U7391, U7392, U7393, U7394, U7395, U7396, U7397, U7398, U7399, U7400, U7401, U7402, U7403, U7404, U7405, U7406, U7407, U7408, U7409, U7410, U7411, U7412, U7413, U7414, U7415, U7416, U7417, U7418, U7419, U7420, U7421, U7422, U7423, U7424, U7425, U7426, U7427, U7428, U7429, U7430, U7431, U7432, U7433, U7434, U7435, U7436, U7437, U7438, U7439, U7440, U7441, U7442, U7443, U7444, U7445, U7446, U7447, U7448, U7449, U7450, U7451, U7452, U7453, U7454, U7455, U7456, U7457, U7458, U7459, U7460, U7461, U7462, U7463, U7464, U7465, U7466, U7467, U7468, U7469, U7470, U7471, U7472, U7473, U7474, U7475, U7476, U7477, U7478, U7479, U7480, U7481, U7482, U7483, U7484, U7485, U7486, U7487, U7488, U7489, U7490, U7491, U7492, U7493, U7494, U7495, U7496, U7497, U7498, U7499, U7500, U7501, U7502, U7503, U7504, U7505, U7506, U7507, U7508, U7509, U7510, U7511, U7512, U7513, U7514, U7515, U7516, U7517, U7518, U7519, U7520, U7521, U7522, U7523, U7524, U7525, U7526, U7527, U7528, U7529, U7530, U7531, U7532, U7533, U7534, U7535, U7536, U7537, U7538, U7539, U7540, U7541, U7542, U7543, U7544, U7545, U7546, U7547, U7548, U7549, U7550, U7551, U7552, U7553, U7554, U7555, U7556, U7557, U7558, U7559, U7560, U7561, U7562, U7563, U7564, U7565, U7566, U7567, U7568, U7569, U7570, U7571, U7572, U7573, U7574, U7575, U7576, U7577, U7578, U7579, U7580, U7581, U7582, U7583, U7584, U7585, U7586, U7587, U7588, U7589, U7590, U7591, U7592, U7593, U7594, U7595, U7596, U7597, U7598, U7599, U7600, U7601, U7602, U7603, U7604, U7605, U7606, U7607, U7608, U7609, U7610, U7611, U7612, U7613, U7614, U7615, U7616, U7617, U7618, U7619, U7620, U7621, U7622, U7623, U7624, U7625, U7626, U7627, U7628, U7629, U7630, U7631, U7632, U7633, U7634, U7635, U7636, U7637, U7638, U7639, U7640, U7641, U7642, U7643, U7644, U7645, U7646, U7647, U7648, U7649, U7650, U7651, U7652, U7653, U7654, U7655, U7656, U7657, U7658, U7659, U7660, U7661, U7662, U7663, U7664, U7665, U7666, U7667, U7668, U7669, U7670, U7671, U7672, U7673, U7674, U7675, U7676, U7677, U7678, U7679, U7680, U7681, U7682, U7683, U7684, U7685, U7686, U7687, U7688, U7689, U7690, U7691, U7692, U7693, U7694, U7695, U7696, U7697, U7698, U7699, U7700, U7701, U7702, U7703, U7704, U7705, U7706, U7707, U7708, U7709, U7710, U7711, U7712, U7713, U7714, U7715, U7716, U7717, U7718, U7719, U7720, U7721, U7722, U7723, U7724, U7725, U7726, U7727, U7728, U7729, U7730, U7731, U7732, U7733, U7734, U7735, U7736, U7737, U7738, U7739, U7740, U7741, U7742, U7743, U7744, U7745, U7746, U7747, U7748, U7749, U7750, U7751, U7752, U7753, U7754, U7755, U7756, U7757, U7758, U7759, U7760, U7761, U7762, U7763, U7764, U7765, U7766, U7767, U7768, U7769, U7770, U7771, U7772, U7773, U7774, U7775, U7776, U7777, U7778, U7779, U7780, U7781, U7782, U2995_in, U2995_pert;

  buf ginst1 (ADDRESS_REG_0__SCAN_IN_BUFF, ADDRESS_REG_0__SCAN_IN);
  buf ginst2 (ADDRESS_REG_10__SCAN_IN_BUFF, ADDRESS_REG_10__SCAN_IN);
  buf ginst3 (ADDRESS_REG_11__SCAN_IN_BUFF, ADDRESS_REG_11__SCAN_IN);
  buf ginst4 (ADDRESS_REG_12__SCAN_IN_BUFF, ADDRESS_REG_12__SCAN_IN);
  buf ginst5 (ADDRESS_REG_13__SCAN_IN_BUFF, ADDRESS_REG_13__SCAN_IN);
  buf ginst6 (ADDRESS_REG_14__SCAN_IN_BUFF, ADDRESS_REG_14__SCAN_IN);
  buf ginst7 (ADDRESS_REG_15__SCAN_IN_BUFF, ADDRESS_REG_15__SCAN_IN);
  buf ginst8 (ADDRESS_REG_16__SCAN_IN_BUFF, ADDRESS_REG_16__SCAN_IN);
  buf ginst9 (ADDRESS_REG_17__SCAN_IN_BUFF, ADDRESS_REG_17__SCAN_IN);
  buf ginst10 (ADDRESS_REG_18__SCAN_IN_BUFF, ADDRESS_REG_18__SCAN_IN);
  buf ginst11 (ADDRESS_REG_19__SCAN_IN_BUFF, ADDRESS_REG_19__SCAN_IN);
  buf ginst12 (ADDRESS_REG_1__SCAN_IN_BUFF, ADDRESS_REG_1__SCAN_IN);
  buf ginst13 (ADDRESS_REG_20__SCAN_IN_BUFF, ADDRESS_REG_20__SCAN_IN);
  buf ginst14 (ADDRESS_REG_21__SCAN_IN_BUFF, ADDRESS_REG_21__SCAN_IN);
  buf ginst15 (ADDRESS_REG_22__SCAN_IN_BUFF, ADDRESS_REG_22__SCAN_IN);
  buf ginst16 (ADDRESS_REG_23__SCAN_IN_BUFF, ADDRESS_REG_23__SCAN_IN);
  buf ginst17 (ADDRESS_REG_24__SCAN_IN_BUFF, ADDRESS_REG_24__SCAN_IN);
  buf ginst18 (ADDRESS_REG_25__SCAN_IN_BUFF, ADDRESS_REG_25__SCAN_IN);
  buf ginst19 (ADDRESS_REG_26__SCAN_IN_BUFF, ADDRESS_REG_26__SCAN_IN);
  buf ginst20 (ADDRESS_REG_27__SCAN_IN_BUFF, ADDRESS_REG_27__SCAN_IN);
  buf ginst21 (ADDRESS_REG_28__SCAN_IN_BUFF, ADDRESS_REG_28__SCAN_IN);
  buf ginst22 (ADDRESS_REG_29__SCAN_IN_BUFF, ADDRESS_REG_29__SCAN_IN);
  buf ginst23 (ADDRESS_REG_2__SCAN_IN_BUFF, ADDRESS_REG_2__SCAN_IN);
  buf ginst24 (ADDRESS_REG_3__SCAN_IN_BUFF, ADDRESS_REG_3__SCAN_IN);
  buf ginst25 (ADDRESS_REG_4__SCAN_IN_BUFF, ADDRESS_REG_4__SCAN_IN);
  buf ginst26 (ADDRESS_REG_5__SCAN_IN_BUFF, ADDRESS_REG_5__SCAN_IN);
  buf ginst27 (ADDRESS_REG_6__SCAN_IN_BUFF, ADDRESS_REG_6__SCAN_IN);
  buf ginst28 (ADDRESS_REG_7__SCAN_IN_BUFF, ADDRESS_REG_7__SCAN_IN);
  buf ginst29 (ADDRESS_REG_8__SCAN_IN_BUFF, ADDRESS_REG_8__SCAN_IN);
  buf ginst30 (ADDRESS_REG_9__SCAN_IN_BUFF, ADDRESS_REG_9__SCAN_IN);
  not ginst31 (ADD_371_U10, U3218);
  nand ginst32 (ADD_371_U11, ADD_371_U28, U3218);
  not ginst33 (ADD_371_U12, U3219);
  nand ginst34 (ADD_371_U13, ADD_371_U29, U3219);
  not ginst35 (ADD_371_U14, U3221);
  not ginst36 (ADD_371_U15, U3220);
  not ginst37 (ADD_371_U16, U3216);
  nand ginst38 (ADD_371_U17, ADD_371_U33, ADD_371_U34);
  nand ginst39 (ADD_371_U18, ADD_371_U35, ADD_371_U36);
  nand ginst40 (ADD_371_U19, ADD_371_U37, ADD_371_U38);
  nand ginst41 (ADD_371_U20, ADD_371_U39, ADD_371_U40);
  nand ginst42 (ADD_371_U21, ADD_371_U43, ADD_371_U44);
  and ginst43 (ADD_371_U22, U3220, U3221);
  nand ginst44 (ADD_371_U23, ADD_371_U30, U3220);
  nand ginst45 (ADD_371_U24, ADD_371_U16, ADD_371_U26);
  and ginst46 (ADD_371_U25, ADD_371_U41, ADD_371_U42);
  nand ginst47 (ADD_371_U26, U3214, U3215);
  not ginst48 (ADD_371_U27, ADD_371_U24);
  not ginst49 (ADD_371_U28, ADD_371_U9);
  not ginst50 (ADD_371_U29, ADD_371_U11);
  not ginst51 (ADD_371_U30, ADD_371_U13);
  not ginst52 (ADD_371_U31, ADD_371_U23);
  nand ginst53 (ADD_371_U32, U3214, U3215, U3216);
  nand ginst54 (ADD_371_U33, ADD_371_U23, U3221);
  nand ginst55 (ADD_371_U34, ADD_371_U14, ADD_371_U31);
  nand ginst56 (ADD_371_U35, ADD_371_U13, U3220);
  nand ginst57 (ADD_371_U36, ADD_371_U15, ADD_371_U30);
  nand ginst58 (ADD_371_U37, ADD_371_U11, U3219);
  nand ginst59 (ADD_371_U38, ADD_371_U12, ADD_371_U29);
  nand ginst60 (ADD_371_U39, ADD_371_U9, U3218);
  not ginst61 (ADD_371_U4, U3214);
  nand ginst62 (ADD_371_U40, ADD_371_U10, ADD_371_U28);
  nand ginst63 (ADD_371_U41, ADD_371_U24, U3217);
  nand ginst64 (ADD_371_U42, ADD_371_U27, ADD_371_U8);
  nand ginst65 (ADD_371_U43, ADD_371_U4, U3215);
  nand ginst66 (ADD_371_U44, ADD_371_U7, U3214);
  nand ginst67 (ADD_371_U5, ADD_371_U24, ADD_371_U32);
  and ginst68 (ADD_371_U6, ADD_371_U22, ADD_371_U30);
  not ginst69 (ADD_371_U7, U3215);
  not ginst70 (ADD_371_U8, U3217);
  nand ginst71 (ADD_371_U9, ADD_371_U24, U3217);
  nand ginst72 (ADD_405_U10, INSTADDRPOINTER_REG_4__SCAN_IN, ADD_405_U98);
  not ginst73 (ADD_405_U100, ADD_405_U12);
  not ginst74 (ADD_405_U101, ADD_405_U14);
  not ginst75 (ADD_405_U102, ADD_405_U16);
  not ginst76 (ADD_405_U103, ADD_405_U19);
  not ginst77 (ADD_405_U104, ADD_405_U20);
  not ginst78 (ADD_405_U105, ADD_405_U22);
  not ginst79 (ADD_405_U106, ADD_405_U24);
  not ginst80 (ADD_405_U107, ADD_405_U26);
  not ginst81 (ADD_405_U108, ADD_405_U28);
  not ginst82 (ADD_405_U109, ADD_405_U30);
  not ginst83 (ADD_405_U11, INSTADDRPOINTER_REG_5__SCAN_IN);
  not ginst84 (ADD_405_U110, ADD_405_U32);
  not ginst85 (ADD_405_U111, ADD_405_U34);
  not ginst86 (ADD_405_U112, ADD_405_U36);
  not ginst87 (ADD_405_U113, ADD_405_U38);
  not ginst88 (ADD_405_U114, ADD_405_U40);
  not ginst89 (ADD_405_U115, ADD_405_U42);
  not ginst90 (ADD_405_U116, ADD_405_U44);
  not ginst91 (ADD_405_U117, ADD_405_U46);
  not ginst92 (ADD_405_U118, ADD_405_U48);
  not ginst93 (ADD_405_U119, ADD_405_U50);
  nand ginst94 (ADD_405_U12, INSTADDRPOINTER_REG_5__SCAN_IN, ADD_405_U99);
  not ginst95 (ADD_405_U120, ADD_405_U52);
  not ginst96 (ADD_405_U121, ADD_405_U54);
  not ginst97 (ADD_405_U122, ADD_405_U56);
  not ginst98 (ADD_405_U123, ADD_405_U58);
  not ginst99 (ADD_405_U124, ADD_405_U60);
  not ginst100 (ADD_405_U125, ADD_405_U95);
  nand ginst101 (ADD_405_U126, INSTADDRPOINTER_REG_0__SCAN_IN, INSTADDRPOINTER_REG_1__SCAN_IN, INSTADDRPOINTER_REG_2__SCAN_IN);
  nand ginst102 (ADD_405_U127, INSTADDRPOINTER_REG_9__SCAN_IN, ADD_405_U19);
  nand ginst103 (ADD_405_U128, ADD_405_U103, ADD_405_U18);
  nand ginst104 (ADD_405_U129, INSTADDRPOINTER_REG_8__SCAN_IN, ADD_405_U16);
  not ginst105 (ADD_405_U13, INSTADDRPOINTER_REG_6__SCAN_IN);
  nand ginst106 (ADD_405_U130, ADD_405_U102, ADD_405_U17);
  nand ginst107 (ADD_405_U131, INSTADDRPOINTER_REG_7__SCAN_IN, ADD_405_U14);
  nand ginst108 (ADD_405_U132, ADD_405_U101, ADD_405_U15);
  nand ginst109 (ADD_405_U133, INSTADDRPOINTER_REG_6__SCAN_IN, ADD_405_U12);
  nand ginst110 (ADD_405_U134, ADD_405_U100, ADD_405_U13);
  nand ginst111 (ADD_405_U135, INSTADDRPOINTER_REG_5__SCAN_IN, ADD_405_U10);
  nand ginst112 (ADD_405_U136, ADD_405_U11, ADD_405_U99);
  nand ginst113 (ADD_405_U137, INSTADDRPOINTER_REG_4__SCAN_IN, ADD_405_U8);
  nand ginst114 (ADD_405_U138, ADD_405_U9, ADD_405_U98);
  nand ginst115 (ADD_405_U139, INSTADDRPOINTER_REG_3__SCAN_IN, ADD_405_U92);
  nand ginst116 (ADD_405_U14, INSTADDRPOINTER_REG_6__SCAN_IN, ADD_405_U100);
  nand ginst117 (ADD_405_U140, ADD_405_U7, ADD_405_U97);
  nand ginst118 (ADD_405_U141, INSTADDRPOINTER_REG_31__SCAN_IN, ADD_405_U95);
  nand ginst119 (ADD_405_U142, ADD_405_U125, ADD_405_U94);
  nand ginst120 (ADD_405_U143, INSTADDRPOINTER_REG_30__SCAN_IN, ADD_405_U60);
  nand ginst121 (ADD_405_U144, ADD_405_U124, ADD_405_U61);
  nand ginst122 (ADD_405_U145, INSTADDRPOINTER_REG_29__SCAN_IN, ADD_405_U58);
  nand ginst123 (ADD_405_U146, ADD_405_U123, ADD_405_U59);
  nand ginst124 (ADD_405_U147, INSTADDRPOINTER_REG_28__SCAN_IN, ADD_405_U56);
  nand ginst125 (ADD_405_U148, ADD_405_U122, ADD_405_U57);
  nand ginst126 (ADD_405_U149, INSTADDRPOINTER_REG_27__SCAN_IN, ADD_405_U54);
  not ginst127 (ADD_405_U15, INSTADDRPOINTER_REG_7__SCAN_IN);
  nand ginst128 (ADD_405_U150, ADD_405_U121, ADD_405_U55);
  nand ginst129 (ADD_405_U151, INSTADDRPOINTER_REG_26__SCAN_IN, ADD_405_U52);
  nand ginst130 (ADD_405_U152, ADD_405_U120, ADD_405_U53);
  nand ginst131 (ADD_405_U153, INSTADDRPOINTER_REG_25__SCAN_IN, ADD_405_U50);
  nand ginst132 (ADD_405_U154, ADD_405_U119, ADD_405_U51);
  nand ginst133 (ADD_405_U155, INSTADDRPOINTER_REG_24__SCAN_IN, ADD_405_U48);
  nand ginst134 (ADD_405_U156, ADD_405_U118, ADD_405_U49);
  nand ginst135 (ADD_405_U157, INSTADDRPOINTER_REG_23__SCAN_IN, ADD_405_U46);
  nand ginst136 (ADD_405_U158, ADD_405_U117, ADD_405_U47);
  nand ginst137 (ADD_405_U159, INSTADDRPOINTER_REG_22__SCAN_IN, ADD_405_U44);
  nand ginst138 (ADD_405_U16, INSTADDRPOINTER_REG_7__SCAN_IN, ADD_405_U101);
  nand ginst139 (ADD_405_U160, ADD_405_U116, ADD_405_U45);
  nand ginst140 (ADD_405_U161, INSTADDRPOINTER_REG_21__SCAN_IN, ADD_405_U42);
  nand ginst141 (ADD_405_U162, ADD_405_U115, ADD_405_U43);
  nand ginst142 (ADD_405_U163, INSTADDRPOINTER_REG_20__SCAN_IN, ADD_405_U40);
  nand ginst143 (ADD_405_U164, ADD_405_U114, ADD_405_U41);
  nand ginst144 (ADD_405_U165, INSTADDRPOINTER_REG_1__SCAN_IN, ADD_405_U4);
  nand ginst145 (ADD_405_U166, INSTADDRPOINTER_REG_0__SCAN_IN, ADD_405_U6);
  nand ginst146 (ADD_405_U167, INSTADDRPOINTER_REG_19__SCAN_IN, ADD_405_U38);
  nand ginst147 (ADD_405_U168, ADD_405_U113, ADD_405_U39);
  nand ginst148 (ADD_405_U169, INSTADDRPOINTER_REG_18__SCAN_IN, ADD_405_U36);
  not ginst149 (ADD_405_U17, INSTADDRPOINTER_REG_8__SCAN_IN);
  nand ginst150 (ADD_405_U170, ADD_405_U112, ADD_405_U37);
  nand ginst151 (ADD_405_U171, INSTADDRPOINTER_REG_17__SCAN_IN, ADD_405_U34);
  nand ginst152 (ADD_405_U172, ADD_405_U111, ADD_405_U35);
  nand ginst153 (ADD_405_U173, INSTADDRPOINTER_REG_16__SCAN_IN, ADD_405_U32);
  nand ginst154 (ADD_405_U174, ADD_405_U110, ADD_405_U33);
  nand ginst155 (ADD_405_U175, INSTADDRPOINTER_REG_15__SCAN_IN, ADD_405_U30);
  nand ginst156 (ADD_405_U176, ADD_405_U109, ADD_405_U31);
  nand ginst157 (ADD_405_U177, INSTADDRPOINTER_REG_14__SCAN_IN, ADD_405_U28);
  nand ginst158 (ADD_405_U178, ADD_405_U108, ADD_405_U29);
  nand ginst159 (ADD_405_U179, INSTADDRPOINTER_REG_13__SCAN_IN, ADD_405_U26);
  not ginst160 (ADD_405_U18, INSTADDRPOINTER_REG_9__SCAN_IN);
  nand ginst161 (ADD_405_U180, ADD_405_U107, ADD_405_U27);
  nand ginst162 (ADD_405_U181, INSTADDRPOINTER_REG_12__SCAN_IN, ADD_405_U24);
  nand ginst163 (ADD_405_U182, ADD_405_U106, ADD_405_U25);
  nand ginst164 (ADD_405_U183, INSTADDRPOINTER_REG_11__SCAN_IN, ADD_405_U22);
  nand ginst165 (ADD_405_U184, ADD_405_U105, ADD_405_U23);
  nand ginst166 (ADD_405_U185, INSTADDRPOINTER_REG_10__SCAN_IN, ADD_405_U20);
  nand ginst167 (ADD_405_U186, ADD_405_U104, ADD_405_U21);
  nand ginst168 (ADD_405_U19, INSTADDRPOINTER_REG_8__SCAN_IN, ADD_405_U102);
  nand ginst169 (ADD_405_U20, INSTADDRPOINTER_REG_9__SCAN_IN, ADD_405_U103);
  not ginst170 (ADD_405_U21, INSTADDRPOINTER_REG_10__SCAN_IN);
  nand ginst171 (ADD_405_U22, INSTADDRPOINTER_REG_10__SCAN_IN, ADD_405_U104);
  not ginst172 (ADD_405_U23, INSTADDRPOINTER_REG_11__SCAN_IN);
  nand ginst173 (ADD_405_U24, INSTADDRPOINTER_REG_11__SCAN_IN, ADD_405_U105);
  not ginst174 (ADD_405_U25, INSTADDRPOINTER_REG_12__SCAN_IN);
  nand ginst175 (ADD_405_U26, INSTADDRPOINTER_REG_12__SCAN_IN, ADD_405_U106);
  not ginst176 (ADD_405_U27, INSTADDRPOINTER_REG_13__SCAN_IN);
  nand ginst177 (ADD_405_U28, INSTADDRPOINTER_REG_13__SCAN_IN, ADD_405_U107);
  not ginst178 (ADD_405_U29, INSTADDRPOINTER_REG_14__SCAN_IN);
  nand ginst179 (ADD_405_U30, INSTADDRPOINTER_REG_14__SCAN_IN, ADD_405_U108);
  not ginst180 (ADD_405_U31, INSTADDRPOINTER_REG_15__SCAN_IN);
  nand ginst181 (ADD_405_U32, INSTADDRPOINTER_REG_15__SCAN_IN, ADD_405_U109);
  not ginst182 (ADD_405_U33, INSTADDRPOINTER_REG_16__SCAN_IN);
  nand ginst183 (ADD_405_U34, INSTADDRPOINTER_REG_16__SCAN_IN, ADD_405_U110);
  not ginst184 (ADD_405_U35, INSTADDRPOINTER_REG_17__SCAN_IN);
  nand ginst185 (ADD_405_U36, INSTADDRPOINTER_REG_17__SCAN_IN, ADD_405_U111);
  not ginst186 (ADD_405_U37, INSTADDRPOINTER_REG_18__SCAN_IN);
  nand ginst187 (ADD_405_U38, INSTADDRPOINTER_REG_18__SCAN_IN, ADD_405_U112);
  not ginst188 (ADD_405_U39, INSTADDRPOINTER_REG_19__SCAN_IN);
  not ginst189 (ADD_405_U4, INSTADDRPOINTER_REG_0__SCAN_IN);
  nand ginst190 (ADD_405_U40, INSTADDRPOINTER_REG_19__SCAN_IN, ADD_405_U113);
  not ginst191 (ADD_405_U41, INSTADDRPOINTER_REG_20__SCAN_IN);
  nand ginst192 (ADD_405_U42, INSTADDRPOINTER_REG_20__SCAN_IN, ADD_405_U114);
  not ginst193 (ADD_405_U43, INSTADDRPOINTER_REG_21__SCAN_IN);
  nand ginst194 (ADD_405_U44, INSTADDRPOINTER_REG_21__SCAN_IN, ADD_405_U115);
  not ginst195 (ADD_405_U45, INSTADDRPOINTER_REG_22__SCAN_IN);
  nand ginst196 (ADD_405_U46, INSTADDRPOINTER_REG_22__SCAN_IN, ADD_405_U116);
  not ginst197 (ADD_405_U47, INSTADDRPOINTER_REG_23__SCAN_IN);
  nand ginst198 (ADD_405_U48, INSTADDRPOINTER_REG_23__SCAN_IN, ADD_405_U117);
  not ginst199 (ADD_405_U49, INSTADDRPOINTER_REG_24__SCAN_IN);
  nand ginst200 (ADD_405_U5, ADD_405_U126, ADD_405_U92);
  nand ginst201 (ADD_405_U50, INSTADDRPOINTER_REG_24__SCAN_IN, ADD_405_U118);
  not ginst202 (ADD_405_U51, INSTADDRPOINTER_REG_25__SCAN_IN);
  nand ginst203 (ADD_405_U52, INSTADDRPOINTER_REG_25__SCAN_IN, ADD_405_U119);
  not ginst204 (ADD_405_U53, INSTADDRPOINTER_REG_26__SCAN_IN);
  nand ginst205 (ADD_405_U54, INSTADDRPOINTER_REG_26__SCAN_IN, ADD_405_U120);
  not ginst206 (ADD_405_U55, INSTADDRPOINTER_REG_27__SCAN_IN);
  nand ginst207 (ADD_405_U56, INSTADDRPOINTER_REG_27__SCAN_IN, ADD_405_U121);
  not ginst208 (ADD_405_U57, INSTADDRPOINTER_REG_28__SCAN_IN);
  nand ginst209 (ADD_405_U58, INSTADDRPOINTER_REG_28__SCAN_IN, ADD_405_U122);
  not ginst210 (ADD_405_U59, INSTADDRPOINTER_REG_29__SCAN_IN);
  not ginst211 (ADD_405_U6, INSTADDRPOINTER_REG_1__SCAN_IN);
  nand ginst212 (ADD_405_U60, INSTADDRPOINTER_REG_29__SCAN_IN, ADD_405_U123);
  not ginst213 (ADD_405_U61, INSTADDRPOINTER_REG_30__SCAN_IN);
  not ginst214 (ADD_405_U62, INSTADDRPOINTER_REG_2__SCAN_IN);
  nand ginst215 (ADD_405_U63, ADD_405_U127, ADD_405_U128);
  nand ginst216 (ADD_405_U64, ADD_405_U129, ADD_405_U130);
  nand ginst217 (ADD_405_U65, ADD_405_U131, ADD_405_U132);
  nand ginst218 (ADD_405_U66, ADD_405_U133, ADD_405_U134);
  nand ginst219 (ADD_405_U67, ADD_405_U135, ADD_405_U136);
  nand ginst220 (ADD_405_U68, ADD_405_U137, ADD_405_U138);
  nand ginst221 (ADD_405_U69, ADD_405_U141, ADD_405_U142);
  not ginst222 (ADD_405_U7, INSTADDRPOINTER_REG_3__SCAN_IN);
  nand ginst223 (ADD_405_U70, ADD_405_U143, ADD_405_U144);
  nand ginst224 (ADD_405_U71, ADD_405_U145, ADD_405_U146);
  nand ginst225 (ADD_405_U72, ADD_405_U147, ADD_405_U148);
  nand ginst226 (ADD_405_U73, ADD_405_U149, ADD_405_U150);
  nand ginst227 (ADD_405_U74, ADD_405_U151, ADD_405_U152);
  nand ginst228 (ADD_405_U75, ADD_405_U153, ADD_405_U154);
  nand ginst229 (ADD_405_U76, ADD_405_U155, ADD_405_U156);
  nand ginst230 (ADD_405_U77, ADD_405_U157, ADD_405_U158);
  nand ginst231 (ADD_405_U78, ADD_405_U159, ADD_405_U160);
  nand ginst232 (ADD_405_U79, ADD_405_U161, ADD_405_U162);
  nand ginst233 (ADD_405_U8, INSTADDRPOINTER_REG_3__SCAN_IN, ADD_405_U92);
  nand ginst234 (ADD_405_U80, ADD_405_U163, ADD_405_U164);
  nand ginst235 (ADD_405_U81, ADD_405_U165, ADD_405_U166);
  nand ginst236 (ADD_405_U82, ADD_405_U167, ADD_405_U168);
  nand ginst237 (ADD_405_U83, ADD_405_U169, ADD_405_U170);
  nand ginst238 (ADD_405_U84, ADD_405_U171, ADD_405_U172);
  nand ginst239 (ADD_405_U85, ADD_405_U173, ADD_405_U174);
  nand ginst240 (ADD_405_U86, ADD_405_U175, ADD_405_U176);
  nand ginst241 (ADD_405_U87, ADD_405_U177, ADD_405_U178);
  nand ginst242 (ADD_405_U88, ADD_405_U179, ADD_405_U180);
  nand ginst243 (ADD_405_U89, ADD_405_U181, ADD_405_U182);
  not ginst244 (ADD_405_U9, INSTADDRPOINTER_REG_4__SCAN_IN);
  nand ginst245 (ADD_405_U90, ADD_405_U183, ADD_405_U184);
  nand ginst246 (ADD_405_U91, ADD_405_U185, ADD_405_U186);
  nand ginst247 (ADD_405_U92, ADD_405_U62, ADD_405_U96);
  and ginst248 (ADD_405_U93, ADD_405_U139, ADD_405_U140);
  not ginst249 (ADD_405_U94, INSTADDRPOINTER_REG_31__SCAN_IN);
  nand ginst250 (ADD_405_U95, INSTADDRPOINTER_REG_30__SCAN_IN, ADD_405_U124);
  nand ginst251 (ADD_405_U96, INSTADDRPOINTER_REG_0__SCAN_IN, INSTADDRPOINTER_REG_1__SCAN_IN);
  not ginst252 (ADD_405_U97, ADD_405_U92);
  not ginst253 (ADD_405_U98, ADD_405_U8);
  not ginst254 (ADD_405_U99, ADD_405_U10);
  nand ginst255 (ADD_515_U10, INSTADDRPOINTER_REG_4__SCAN_IN, ADD_515_U95);
  not ginst256 (ADD_515_U100, ADD_515_U19);
  not ginst257 (ADD_515_U101, ADD_515_U20);
  not ginst258 (ADD_515_U102, ADD_515_U22);
  not ginst259 (ADD_515_U103, ADD_515_U24);
  not ginst260 (ADD_515_U104, ADD_515_U26);
  not ginst261 (ADD_515_U105, ADD_515_U28);
  not ginst262 (ADD_515_U106, ADD_515_U30);
  not ginst263 (ADD_515_U107, ADD_515_U32);
  not ginst264 (ADD_515_U108, ADD_515_U34);
  not ginst265 (ADD_515_U109, ADD_515_U36);
  not ginst266 (ADD_515_U11, INSTADDRPOINTER_REG_5__SCAN_IN);
  not ginst267 (ADD_515_U110, ADD_515_U38);
  not ginst268 (ADD_515_U111, ADD_515_U40);
  not ginst269 (ADD_515_U112, ADD_515_U42);
  not ginst270 (ADD_515_U113, ADD_515_U44);
  not ginst271 (ADD_515_U114, ADD_515_U46);
  not ginst272 (ADD_515_U115, ADD_515_U48);
  not ginst273 (ADD_515_U116, ADD_515_U50);
  not ginst274 (ADD_515_U117, ADD_515_U52);
  not ginst275 (ADD_515_U118, ADD_515_U54);
  not ginst276 (ADD_515_U119, ADD_515_U56);
  nand ginst277 (ADD_515_U12, INSTADDRPOINTER_REG_5__SCAN_IN, ADD_515_U96);
  not ginst278 (ADD_515_U120, ADD_515_U58);
  not ginst279 (ADD_515_U121, ADD_515_U60);
  not ginst280 (ADD_515_U122, ADD_515_U93);
  nand ginst281 (ADD_515_U123, INSTADDRPOINTER_REG_9__SCAN_IN, ADD_515_U19);
  nand ginst282 (ADD_515_U124, ADD_515_U100, ADD_515_U18);
  nand ginst283 (ADD_515_U125, INSTADDRPOINTER_REG_8__SCAN_IN, ADD_515_U16);
  nand ginst284 (ADD_515_U126, ADD_515_U17, ADD_515_U99);
  nand ginst285 (ADD_515_U127, INSTADDRPOINTER_REG_7__SCAN_IN, ADD_515_U14);
  nand ginst286 (ADD_515_U128, ADD_515_U15, ADD_515_U98);
  nand ginst287 (ADD_515_U129, INSTADDRPOINTER_REG_6__SCAN_IN, ADD_515_U12);
  not ginst288 (ADD_515_U13, INSTADDRPOINTER_REG_6__SCAN_IN);
  nand ginst289 (ADD_515_U130, ADD_515_U13, ADD_515_U97);
  nand ginst290 (ADD_515_U131, INSTADDRPOINTER_REG_5__SCAN_IN, ADD_515_U10);
  nand ginst291 (ADD_515_U132, ADD_515_U11, ADD_515_U96);
  nand ginst292 (ADD_515_U133, INSTADDRPOINTER_REG_4__SCAN_IN, ADD_515_U8);
  nand ginst293 (ADD_515_U134, ADD_515_U9, ADD_515_U95);
  nand ginst294 (ADD_515_U135, INSTADDRPOINTER_REG_3__SCAN_IN, ADD_515_U6);
  nand ginst295 (ADD_515_U136, ADD_515_U7, ADD_515_U94);
  nand ginst296 (ADD_515_U137, INSTADDRPOINTER_REG_31__SCAN_IN, ADD_515_U93);
  nand ginst297 (ADD_515_U138, ADD_515_U122, ADD_515_U92);
  nand ginst298 (ADD_515_U139, INSTADDRPOINTER_REG_30__SCAN_IN, ADD_515_U60);
  nand ginst299 (ADD_515_U14, INSTADDRPOINTER_REG_6__SCAN_IN, ADD_515_U97);
  nand ginst300 (ADD_515_U140, ADD_515_U121, ADD_515_U61);
  nand ginst301 (ADD_515_U141, INSTADDRPOINTER_REG_2__SCAN_IN, ADD_515_U4);
  nand ginst302 (ADD_515_U142, INSTADDRPOINTER_REG_1__SCAN_IN, ADD_515_U5);
  nand ginst303 (ADD_515_U143, INSTADDRPOINTER_REG_29__SCAN_IN, ADD_515_U58);
  nand ginst304 (ADD_515_U144, ADD_515_U120, ADD_515_U59);
  nand ginst305 (ADD_515_U145, INSTADDRPOINTER_REG_28__SCAN_IN, ADD_515_U56);
  nand ginst306 (ADD_515_U146, ADD_515_U119, ADD_515_U57);
  nand ginst307 (ADD_515_U147, INSTADDRPOINTER_REG_27__SCAN_IN, ADD_515_U54);
  nand ginst308 (ADD_515_U148, ADD_515_U118, ADD_515_U55);
  nand ginst309 (ADD_515_U149, INSTADDRPOINTER_REG_26__SCAN_IN, ADD_515_U52);
  not ginst310 (ADD_515_U15, INSTADDRPOINTER_REG_7__SCAN_IN);
  nand ginst311 (ADD_515_U150, ADD_515_U117, ADD_515_U53);
  nand ginst312 (ADD_515_U151, INSTADDRPOINTER_REG_25__SCAN_IN, ADD_515_U50);
  nand ginst313 (ADD_515_U152, ADD_515_U116, ADD_515_U51);
  nand ginst314 (ADD_515_U153, INSTADDRPOINTER_REG_24__SCAN_IN, ADD_515_U48);
  nand ginst315 (ADD_515_U154, ADD_515_U115, ADD_515_U49);
  nand ginst316 (ADD_515_U155, INSTADDRPOINTER_REG_23__SCAN_IN, ADD_515_U46);
  nand ginst317 (ADD_515_U156, ADD_515_U114, ADD_515_U47);
  nand ginst318 (ADD_515_U157, INSTADDRPOINTER_REG_22__SCAN_IN, ADD_515_U44);
  nand ginst319 (ADD_515_U158, ADD_515_U113, ADD_515_U45);
  nand ginst320 (ADD_515_U159, INSTADDRPOINTER_REG_21__SCAN_IN, ADD_515_U42);
  nand ginst321 (ADD_515_U16, INSTADDRPOINTER_REG_7__SCAN_IN, ADD_515_U98);
  nand ginst322 (ADD_515_U160, ADD_515_U112, ADD_515_U43);
  nand ginst323 (ADD_515_U161, INSTADDRPOINTER_REG_20__SCAN_IN, ADD_515_U40);
  nand ginst324 (ADD_515_U162, ADD_515_U111, ADD_515_U41);
  nand ginst325 (ADD_515_U163, INSTADDRPOINTER_REG_19__SCAN_IN, ADD_515_U38);
  nand ginst326 (ADD_515_U164, ADD_515_U110, ADD_515_U39);
  nand ginst327 (ADD_515_U165, INSTADDRPOINTER_REG_18__SCAN_IN, ADD_515_U36);
  nand ginst328 (ADD_515_U166, ADD_515_U109, ADD_515_U37);
  nand ginst329 (ADD_515_U167, INSTADDRPOINTER_REG_17__SCAN_IN, ADD_515_U34);
  nand ginst330 (ADD_515_U168, ADD_515_U108, ADD_515_U35);
  nand ginst331 (ADD_515_U169, INSTADDRPOINTER_REG_16__SCAN_IN, ADD_515_U32);
  not ginst332 (ADD_515_U17, INSTADDRPOINTER_REG_8__SCAN_IN);
  nand ginst333 (ADD_515_U170, ADD_515_U107, ADD_515_U33);
  nand ginst334 (ADD_515_U171, INSTADDRPOINTER_REG_15__SCAN_IN, ADD_515_U30);
  nand ginst335 (ADD_515_U172, ADD_515_U106, ADD_515_U31);
  nand ginst336 (ADD_515_U173, INSTADDRPOINTER_REG_14__SCAN_IN, ADD_515_U28);
  nand ginst337 (ADD_515_U174, ADD_515_U105, ADD_515_U29);
  nand ginst338 (ADD_515_U175, INSTADDRPOINTER_REG_13__SCAN_IN, ADD_515_U26);
  nand ginst339 (ADD_515_U176, ADD_515_U104, ADD_515_U27);
  nand ginst340 (ADD_515_U177, INSTADDRPOINTER_REG_12__SCAN_IN, ADD_515_U24);
  nand ginst341 (ADD_515_U178, ADD_515_U103, ADD_515_U25);
  nand ginst342 (ADD_515_U179, INSTADDRPOINTER_REG_11__SCAN_IN, ADD_515_U22);
  not ginst343 (ADD_515_U18, INSTADDRPOINTER_REG_9__SCAN_IN);
  nand ginst344 (ADD_515_U180, ADD_515_U102, ADD_515_U23);
  nand ginst345 (ADD_515_U181, INSTADDRPOINTER_REG_10__SCAN_IN, ADD_515_U20);
  nand ginst346 (ADD_515_U182, ADD_515_U101, ADD_515_U21);
  nand ginst347 (ADD_515_U19, INSTADDRPOINTER_REG_8__SCAN_IN, ADD_515_U99);
  nand ginst348 (ADD_515_U20, INSTADDRPOINTER_REG_9__SCAN_IN, ADD_515_U100);
  not ginst349 (ADD_515_U21, INSTADDRPOINTER_REG_10__SCAN_IN);
  nand ginst350 (ADD_515_U22, INSTADDRPOINTER_REG_10__SCAN_IN, ADD_515_U101);
  not ginst351 (ADD_515_U23, INSTADDRPOINTER_REG_11__SCAN_IN);
  nand ginst352 (ADD_515_U24, INSTADDRPOINTER_REG_11__SCAN_IN, ADD_515_U102);
  not ginst353 (ADD_515_U25, INSTADDRPOINTER_REG_12__SCAN_IN);
  nand ginst354 (ADD_515_U26, INSTADDRPOINTER_REG_12__SCAN_IN, ADD_515_U103);
  not ginst355 (ADD_515_U27, INSTADDRPOINTER_REG_13__SCAN_IN);
  nand ginst356 (ADD_515_U28, INSTADDRPOINTER_REG_13__SCAN_IN, ADD_515_U104);
  not ginst357 (ADD_515_U29, INSTADDRPOINTER_REG_14__SCAN_IN);
  nand ginst358 (ADD_515_U30, INSTADDRPOINTER_REG_14__SCAN_IN, ADD_515_U105);
  not ginst359 (ADD_515_U31, INSTADDRPOINTER_REG_15__SCAN_IN);
  nand ginst360 (ADD_515_U32, INSTADDRPOINTER_REG_15__SCAN_IN, ADD_515_U106);
  not ginst361 (ADD_515_U33, INSTADDRPOINTER_REG_16__SCAN_IN);
  nand ginst362 (ADD_515_U34, INSTADDRPOINTER_REG_16__SCAN_IN, ADD_515_U107);
  not ginst363 (ADD_515_U35, INSTADDRPOINTER_REG_17__SCAN_IN);
  nand ginst364 (ADD_515_U36, INSTADDRPOINTER_REG_17__SCAN_IN, ADD_515_U108);
  not ginst365 (ADD_515_U37, INSTADDRPOINTER_REG_18__SCAN_IN);
  nand ginst366 (ADD_515_U38, INSTADDRPOINTER_REG_18__SCAN_IN, ADD_515_U109);
  not ginst367 (ADD_515_U39, INSTADDRPOINTER_REG_19__SCAN_IN);
  not ginst368 (ADD_515_U4, INSTADDRPOINTER_REG_1__SCAN_IN);
  nand ginst369 (ADD_515_U40, INSTADDRPOINTER_REG_19__SCAN_IN, ADD_515_U110);
  not ginst370 (ADD_515_U41, INSTADDRPOINTER_REG_20__SCAN_IN);
  nand ginst371 (ADD_515_U42, INSTADDRPOINTER_REG_20__SCAN_IN, ADD_515_U111);
  not ginst372 (ADD_515_U43, INSTADDRPOINTER_REG_21__SCAN_IN);
  nand ginst373 (ADD_515_U44, INSTADDRPOINTER_REG_21__SCAN_IN, ADD_515_U112);
  not ginst374 (ADD_515_U45, INSTADDRPOINTER_REG_22__SCAN_IN);
  nand ginst375 (ADD_515_U46, INSTADDRPOINTER_REG_22__SCAN_IN, ADD_515_U113);
  not ginst376 (ADD_515_U47, INSTADDRPOINTER_REG_23__SCAN_IN);
  nand ginst377 (ADD_515_U48, INSTADDRPOINTER_REG_23__SCAN_IN, ADD_515_U114);
  not ginst378 (ADD_515_U49, INSTADDRPOINTER_REG_24__SCAN_IN);
  not ginst379 (ADD_515_U5, INSTADDRPOINTER_REG_2__SCAN_IN);
  nand ginst380 (ADD_515_U50, INSTADDRPOINTER_REG_24__SCAN_IN, ADD_515_U115);
  not ginst381 (ADD_515_U51, INSTADDRPOINTER_REG_25__SCAN_IN);
  nand ginst382 (ADD_515_U52, INSTADDRPOINTER_REG_25__SCAN_IN, ADD_515_U116);
  not ginst383 (ADD_515_U53, INSTADDRPOINTER_REG_26__SCAN_IN);
  nand ginst384 (ADD_515_U54, INSTADDRPOINTER_REG_26__SCAN_IN, ADD_515_U117);
  not ginst385 (ADD_515_U55, INSTADDRPOINTER_REG_27__SCAN_IN);
  nand ginst386 (ADD_515_U56, INSTADDRPOINTER_REG_27__SCAN_IN, ADD_515_U118);
  not ginst387 (ADD_515_U57, INSTADDRPOINTER_REG_28__SCAN_IN);
  nand ginst388 (ADD_515_U58, INSTADDRPOINTER_REG_28__SCAN_IN, ADD_515_U119);
  not ginst389 (ADD_515_U59, INSTADDRPOINTER_REG_29__SCAN_IN);
  nand ginst390 (ADD_515_U6, INSTADDRPOINTER_REG_1__SCAN_IN, INSTADDRPOINTER_REG_2__SCAN_IN);
  nand ginst391 (ADD_515_U60, INSTADDRPOINTER_REG_29__SCAN_IN, ADD_515_U120);
  not ginst392 (ADD_515_U61, INSTADDRPOINTER_REG_30__SCAN_IN);
  nand ginst393 (ADD_515_U62, ADD_515_U123, ADD_515_U124);
  nand ginst394 (ADD_515_U63, ADD_515_U125, ADD_515_U126);
  nand ginst395 (ADD_515_U64, ADD_515_U127, ADD_515_U128);
  nand ginst396 (ADD_515_U65, ADD_515_U129, ADD_515_U130);
  nand ginst397 (ADD_515_U66, ADD_515_U131, ADD_515_U132);
  nand ginst398 (ADD_515_U67, ADD_515_U133, ADD_515_U134);
  nand ginst399 (ADD_515_U68, ADD_515_U135, ADD_515_U136);
  nand ginst400 (ADD_515_U69, ADD_515_U137, ADD_515_U138);
  not ginst401 (ADD_515_U7, INSTADDRPOINTER_REG_3__SCAN_IN);
  nand ginst402 (ADD_515_U70, ADD_515_U139, ADD_515_U140);
  nand ginst403 (ADD_515_U71, ADD_515_U141, ADD_515_U142);
  nand ginst404 (ADD_515_U72, ADD_515_U143, ADD_515_U144);
  nand ginst405 (ADD_515_U73, ADD_515_U145, ADD_515_U146);
  nand ginst406 (ADD_515_U74, ADD_515_U147, ADD_515_U148);
  nand ginst407 (ADD_515_U75, ADD_515_U149, ADD_515_U150);
  nand ginst408 (ADD_515_U76, ADD_515_U151, ADD_515_U152);
  nand ginst409 (ADD_515_U77, ADD_515_U153, ADD_515_U154);
  nand ginst410 (ADD_515_U78, ADD_515_U155, ADD_515_U156);
  nand ginst411 (ADD_515_U79, ADD_515_U157, ADD_515_U158);
  nand ginst412 (ADD_515_U8, INSTADDRPOINTER_REG_3__SCAN_IN, ADD_515_U94);
  nand ginst413 (ADD_515_U80, ADD_515_U159, ADD_515_U160);
  nand ginst414 (ADD_515_U81, ADD_515_U161, ADD_515_U162);
  nand ginst415 (ADD_515_U82, ADD_515_U163, ADD_515_U164);
  nand ginst416 (ADD_515_U83, ADD_515_U165, ADD_515_U166);
  nand ginst417 (ADD_515_U84, ADD_515_U167, ADD_515_U168);
  nand ginst418 (ADD_515_U85, ADD_515_U169, ADD_515_U170);
  nand ginst419 (ADD_515_U86, ADD_515_U171, ADD_515_U172);
  nand ginst420 (ADD_515_U87, ADD_515_U173, ADD_515_U174);
  nand ginst421 (ADD_515_U88, ADD_515_U175, ADD_515_U176);
  nand ginst422 (ADD_515_U89, ADD_515_U177, ADD_515_U178);
  not ginst423 (ADD_515_U9, INSTADDRPOINTER_REG_4__SCAN_IN);
  nand ginst424 (ADD_515_U90, ADD_515_U179, ADD_515_U180);
  nand ginst425 (ADD_515_U91, ADD_515_U181, ADD_515_U182);
  not ginst426 (ADD_515_U92, INSTADDRPOINTER_REG_31__SCAN_IN);
  nand ginst427 (ADD_515_U93, INSTADDRPOINTER_REG_30__SCAN_IN, ADD_515_U121);
  not ginst428 (ADD_515_U94, ADD_515_U6);
  not ginst429 (ADD_515_U95, ADD_515_U8);
  not ginst430 (ADD_515_U96, ADD_515_U10);
  not ginst431 (ADD_515_U97, ADD_515_U12);
  not ginst432 (ADD_515_U98, ADD_515_U14);
  not ginst433 (ADD_515_U99, ADD_515_U16);
  buf ginst434 (ADS_N_REG_SCAN_IN_BUFF, ADS_N_REG_SCAN_IN);
  buf ginst435 (BE_N_REG_0__SCAN_IN_BUFF, BE_N_REG_0__SCAN_IN);
  buf ginst436 (BE_N_REG_1__SCAN_IN_BUFF, BE_N_REG_1__SCAN_IN);
  buf ginst437 (BE_N_REG_2__SCAN_IN_BUFF, BE_N_REG_2__SCAN_IN);
  buf ginst438 (BE_N_REG_3__SCAN_IN_BUFF, BE_N_REG_3__SCAN_IN);
  buf ginst439 (DATAO_REG_0__SCAN_IN_BUFF, DATAO_REG_0__SCAN_IN);
  buf ginst440 (DATAO_REG_10__SCAN_IN_BUFF, DATAO_REG_10__SCAN_IN);
  buf ginst441 (DATAO_REG_11__SCAN_IN_BUFF, DATAO_REG_11__SCAN_IN);
  buf ginst442 (DATAO_REG_12__SCAN_IN_BUFF, DATAO_REG_12__SCAN_IN);
  buf ginst443 (DATAO_REG_13__SCAN_IN_BUFF, DATAO_REG_13__SCAN_IN);
  buf ginst444 (DATAO_REG_14__SCAN_IN_BUFF, DATAO_REG_14__SCAN_IN);
  buf ginst445 (DATAO_REG_15__SCAN_IN_BUFF, DATAO_REG_15__SCAN_IN);
  buf ginst446 (DATAO_REG_16__SCAN_IN_BUFF, DATAO_REG_16__SCAN_IN);
  buf ginst447 (DATAO_REG_17__SCAN_IN_BUFF, DATAO_REG_17__SCAN_IN);
  buf ginst448 (DATAO_REG_18__SCAN_IN_BUFF, DATAO_REG_18__SCAN_IN);
  buf ginst449 (DATAO_REG_19__SCAN_IN_BUFF, DATAO_REG_19__SCAN_IN);
  buf ginst450 (DATAO_REG_1__SCAN_IN_BUFF, DATAO_REG_1__SCAN_IN);
  buf ginst451 (DATAO_REG_20__SCAN_IN_BUFF, DATAO_REG_20__SCAN_IN);
  buf ginst452 (DATAO_REG_21__SCAN_IN_BUFF, DATAO_REG_21__SCAN_IN);
  buf ginst453 (DATAO_REG_22__SCAN_IN_BUFF, DATAO_REG_22__SCAN_IN);
  buf ginst454 (DATAO_REG_23__SCAN_IN_BUFF, DATAO_REG_23__SCAN_IN);
  buf ginst455 (DATAO_REG_24__SCAN_IN_BUFF, DATAO_REG_24__SCAN_IN);
  buf ginst456 (DATAO_REG_25__SCAN_IN_BUFF, DATAO_REG_25__SCAN_IN);
  buf ginst457 (DATAO_REG_26__SCAN_IN_BUFF, DATAO_REG_26__SCAN_IN);
  buf ginst458 (DATAO_REG_27__SCAN_IN_BUFF, DATAO_REG_27__SCAN_IN);
  buf ginst459 (DATAO_REG_28__SCAN_IN_BUFF, DATAO_REG_28__SCAN_IN);
  buf ginst460 (DATAO_REG_29__SCAN_IN_BUFF, DATAO_REG_29__SCAN_IN);
  buf ginst461 (DATAO_REG_2__SCAN_IN_BUFF, DATAO_REG_2__SCAN_IN);
  buf ginst462 (DATAO_REG_30__SCAN_IN_BUFF, DATAO_REG_30__SCAN_IN);
  buf ginst463 (DATAO_REG_31__SCAN_IN_BUFF, DATAO_REG_31__SCAN_IN);
  buf ginst464 (DATAO_REG_3__SCAN_IN_BUFF, DATAO_REG_3__SCAN_IN);
  buf ginst465 (DATAO_REG_4__SCAN_IN_BUFF, DATAO_REG_4__SCAN_IN);
  buf ginst466 (DATAO_REG_5__SCAN_IN_BUFF, DATAO_REG_5__SCAN_IN);
  buf ginst467 (DATAO_REG_6__SCAN_IN_BUFF, DATAO_REG_6__SCAN_IN);
  buf ginst468 (DATAO_REG_7__SCAN_IN_BUFF, DATAO_REG_7__SCAN_IN);
  buf ginst469 (DATAO_REG_8__SCAN_IN_BUFF, DATAO_REG_8__SCAN_IN);
  buf ginst470 (DATAO_REG_9__SCAN_IN_BUFF, DATAO_REG_9__SCAN_IN);
  buf ginst471 (D_C_N_REG_SCAN_IN_BUFF, D_C_N_REG_SCAN_IN);
  nor ginst472 (GTE_485_U6, GTE_485_U7, R2238_U6);
  nor ginst473 (GTE_485_U7, R2238_U19, R2238_U20, R2238_U21, R2238_U22);
  and ginst474 (LT_563_1260_U6, LT_563_1260_U8, LT_563_1260_U9);
  not ginst475 (LT_563_1260_U7, U2673);
  nand ginst476 (LT_563_1260_U8, LT_563_1260_U7, R584_U8);
  nand ginst477 (LT_563_1260_U9, LT_563_1260_U7, R584_U9);
  not ginst478 (LT_563_U10, INSTQUEUEWR_ADDR_REG_3__SCAN_IN);
  not ginst479 (LT_563_U11, INSTQUEUEWR_ADDR_REG_4__SCAN_IN);
  not ginst480 (LT_563_U12, U3476);
  and ginst481 (LT_563_U13, LT_563_U21, LT_563_U22);
  and ginst482 (LT_563_U14, LT_563_U24, LT_563_U25);
  not ginst483 (LT_563_U15, U3479);
  not ginst484 (LT_563_U16, U3480);
  nand ginst485 (LT_563_U17, INSTQUEUEWR_ADDR_REG_0__SCAN_IN, LT_563_U15, LT_563_U16);
  nand ginst486 (LT_563_U18, INSTQUEUEWR_ADDR_REG_1__SCAN_IN, LT_563_U15);
  nand ginst487 (LT_563_U19, INSTQUEUEWR_ADDR_REG_2__SCAN_IN, LT_563_U8);
  nand ginst488 (LT_563_U20, LT_563_U17, LT_563_U18, LT_563_U19, LT_563_U28);
  nand ginst489 (LT_563_U21, LT_563_U7, U3478);
  nand ginst490 (LT_563_U22, LT_563_U10, U3477);
  nand ginst491 (LT_563_U23, LT_563_U13, LT_563_U20);
  nand ginst492 (LT_563_U24, INSTQUEUEWR_ADDR_REG_3__SCAN_IN, LT_563_U9);
  nand ginst493 (LT_563_U25, INSTQUEUEWR_ADDR_REG_4__SCAN_IN, LT_563_U12);
  nand ginst494 (LT_563_U26, LT_563_U14, LT_563_U23);
  nand ginst495 (LT_563_U27, LT_563_U11, U3476);
  nand ginst496 (LT_563_U28, INSTQUEUEWR_ADDR_REG_1__SCAN_IN, INSTQUEUEWR_ADDR_REG_0__SCAN_IN, LT_563_U16);
  and ginst497 (LT_563_U6, LT_563_U26, LT_563_U27);
  not ginst498 (LT_563_U7, INSTQUEUEWR_ADDR_REG_2__SCAN_IN);
  not ginst499 (LT_563_U8, U3478);
  not ginst500 (LT_563_U9, U3477);
  or ginst501 (LT_589_U6, LT_589_U8, U2673);
  and ginst502 (LT_589_U7, R584_U6, R584_U7);
  nor ginst503 (LT_589_U8, LT_589_U7, R584_U8, R584_U9);
  buf ginst504 (M_IO_N_REG_SCAN_IN_BUFF, M_IO_N_REG_SCAN_IN);
  nand ginst505 (R2027_U10, INSTADDRPOINTER_REG_0__SCAN_IN, INSTADDRPOINTER_REG_1__SCAN_IN, INSTADDRPOINTER_REG_2__SCAN_IN);
  nand ginst506 (R2027_U100, INSTADDRPOINTER_REG_0__SCAN_IN, INSTADDRPOINTER_REG_1__SCAN_IN);
  nand ginst507 (R2027_U101, INSTADDRPOINTER_REG_27__SCAN_IN, R2027_U122);
  nand ginst508 (R2027_U102, INSTADDRPOINTER_REG_25__SCAN_IN, R2027_U116);
  nand ginst509 (R2027_U103, INSTADDRPOINTER_REG_23__SCAN_IN, R2027_U115);
  nand ginst510 (R2027_U104, INSTADDRPOINTER_REG_21__SCAN_IN, R2027_U121);
  nand ginst511 (R2027_U105, INSTADDRPOINTER_REG_19__SCAN_IN, R2027_U114);
  nand ginst512 (R2027_U106, INSTADDRPOINTER_REG_17__SCAN_IN, R2027_U117);
  nand ginst513 (R2027_U107, INSTADDRPOINTER_REG_15__SCAN_IN, R2027_U124);
  nand ginst514 (R2027_U108, INSTADDRPOINTER_REG_13__SCAN_IN, R2027_U119);
  nand ginst515 (R2027_U109, INSTADDRPOINTER_REG_11__SCAN_IN, R2027_U113);
  not ginst516 (R2027_U11, INSTADDRPOINTER_REG_6__SCAN_IN);
  nand ginst517 (R2027_U110, INSTADDRPOINTER_REG_9__SCAN_IN, R2027_U120);
  not ginst518 (R2027_U111, R2027_U10);
  not ginst519 (R2027_U112, R2027_U13);
  not ginst520 (R2027_U113, R2027_U22);
  not ginst521 (R2027_U114, R2027_U34);
  not ginst522 (R2027_U115, R2027_U40);
  not ginst523 (R2027_U116, R2027_U43);
  not ginst524 (R2027_U117, R2027_U31);
  not ginst525 (R2027_U118, R2027_U16);
  not ginst526 (R2027_U119, R2027_U25);
  not ginst527 (R2027_U12, INSTADDRPOINTER_REG_5__SCAN_IN);
  not ginst528 (R2027_U120, R2027_U17);
  not ginst529 (R2027_U121, R2027_U36);
  not ginst530 (R2027_U122, R2027_U46);
  not ginst531 (R2027_U123, R2027_U48);
  not ginst532 (R2027_U124, R2027_U27);
  not ginst533 (R2027_U125, R2027_U95);
  not ginst534 (R2027_U126, R2027_U96);
  not ginst535 (R2027_U127, R2027_U97);
  not ginst536 (R2027_U128, R2027_U49);
  not ginst537 (R2027_U129, R2027_U99);
  nand ginst538 (R2027_U13, R2027_U111, R2027_U82);
  not ginst539 (R2027_U130, R2027_U100);
  not ginst540 (R2027_U131, R2027_U101);
  not ginst541 (R2027_U132, R2027_U102);
  not ginst542 (R2027_U133, R2027_U103);
  not ginst543 (R2027_U134, R2027_U104);
  not ginst544 (R2027_U135, R2027_U105);
  not ginst545 (R2027_U136, R2027_U106);
  not ginst546 (R2027_U137, R2027_U107);
  not ginst547 (R2027_U138, R2027_U108);
  not ginst548 (R2027_U139, R2027_U109);
  not ginst549 (R2027_U14, INSTADDRPOINTER_REG_8__SCAN_IN);
  not ginst550 (R2027_U140, R2027_U110);
  nand ginst551 (R2027_U141, R2027_U120, R2027_U18);
  nand ginst552 (R2027_U142, INSTADDRPOINTER_REG_9__SCAN_IN, R2027_U17);
  nand ginst553 (R2027_U143, INSTADDRPOINTER_REG_8__SCAN_IN, R2027_U95);
  nand ginst554 (R2027_U144, R2027_U125, R2027_U14);
  nand ginst555 (R2027_U145, R2027_U118, R2027_U15);
  nand ginst556 (R2027_U146, INSTADDRPOINTER_REG_7__SCAN_IN, R2027_U16);
  nand ginst557 (R2027_U147, INSTADDRPOINTER_REG_6__SCAN_IN, R2027_U96);
  nand ginst558 (R2027_U148, R2027_U11, R2027_U126);
  nand ginst559 (R2027_U149, R2027_U112, R2027_U12);
  not ginst560 (R2027_U15, INSTADDRPOINTER_REG_7__SCAN_IN);
  nand ginst561 (R2027_U150, INSTADDRPOINTER_REG_5__SCAN_IN, R2027_U13);
  nand ginst562 (R2027_U151, INSTADDRPOINTER_REG_4__SCAN_IN, R2027_U97);
  nand ginst563 (R2027_U152, R2027_U127, R2027_U8);
  nand ginst564 (R2027_U153, R2027_U111, R2027_U9);
  nand ginst565 (R2027_U154, INSTADDRPOINTER_REG_3__SCAN_IN, R2027_U10);
  nand ginst566 (R2027_U155, INSTADDRPOINTER_REG_31__SCAN_IN, R2027_U99);
  nand ginst567 (R2027_U156, R2027_U129, R2027_U98);
  nand ginst568 (R2027_U157, INSTADDRPOINTER_REG_30__SCAN_IN, R2027_U49);
  nand ginst569 (R2027_U158, R2027_U128, R2027_U50);
  nand ginst570 (R2027_U159, INSTADDRPOINTER_REG_2__SCAN_IN, R2027_U100);
  nand ginst571 (R2027_U16, R2027_U112, R2027_U83);
  nand ginst572 (R2027_U160, R2027_U130, R2027_U6);
  nand ginst573 (R2027_U161, R2027_U123, R2027_U47);
  nand ginst574 (R2027_U162, INSTADDRPOINTER_REG_29__SCAN_IN, R2027_U48);
  nand ginst575 (R2027_U163, INSTADDRPOINTER_REG_28__SCAN_IN, R2027_U101);
  nand ginst576 (R2027_U164, R2027_U131, R2027_U45);
  nand ginst577 (R2027_U165, R2027_U122, R2027_U44);
  nand ginst578 (R2027_U166, INSTADDRPOINTER_REG_27__SCAN_IN, R2027_U46);
  nand ginst579 (R2027_U167, INSTADDRPOINTER_REG_26__SCAN_IN, R2027_U102);
  nand ginst580 (R2027_U168, R2027_U132, R2027_U41);
  nand ginst581 (R2027_U169, R2027_U116, R2027_U42);
  nand ginst582 (R2027_U17, R2027_U118, R2027_U84);
  nand ginst583 (R2027_U170, INSTADDRPOINTER_REG_25__SCAN_IN, R2027_U43);
  nand ginst584 (R2027_U171, INSTADDRPOINTER_REG_24__SCAN_IN, R2027_U103);
  nand ginst585 (R2027_U172, R2027_U133, R2027_U38);
  nand ginst586 (R2027_U173, R2027_U115, R2027_U39);
  nand ginst587 (R2027_U174, INSTADDRPOINTER_REG_23__SCAN_IN, R2027_U40);
  nand ginst588 (R2027_U175, INSTADDRPOINTER_REG_22__SCAN_IN, R2027_U104);
  nand ginst589 (R2027_U176, R2027_U134, R2027_U37);
  nand ginst590 (R2027_U177, R2027_U121, R2027_U35);
  nand ginst591 (R2027_U178, INSTADDRPOINTER_REG_21__SCAN_IN, R2027_U36);
  nand ginst592 (R2027_U179, INSTADDRPOINTER_REG_20__SCAN_IN, R2027_U105);
  not ginst593 (R2027_U18, INSTADDRPOINTER_REG_9__SCAN_IN);
  nand ginst594 (R2027_U180, R2027_U135, R2027_U32);
  nand ginst595 (R2027_U181, INSTADDRPOINTER_REG_0__SCAN_IN, R2027_U7);
  nand ginst596 (R2027_U182, INSTADDRPOINTER_REG_1__SCAN_IN, R2027_U5);
  nand ginst597 (R2027_U183, R2027_U114, R2027_U33);
  nand ginst598 (R2027_U184, INSTADDRPOINTER_REG_19__SCAN_IN, R2027_U34);
  nand ginst599 (R2027_U185, INSTADDRPOINTER_REG_18__SCAN_IN, R2027_U106);
  nand ginst600 (R2027_U186, R2027_U136, R2027_U29);
  nand ginst601 (R2027_U187, R2027_U117, R2027_U30);
  nand ginst602 (R2027_U188, INSTADDRPOINTER_REG_17__SCAN_IN, R2027_U31);
  nand ginst603 (R2027_U189, INSTADDRPOINTER_REG_16__SCAN_IN, R2027_U107);
  not ginst604 (R2027_U19, INSTADDRPOINTER_REG_10__SCAN_IN);
  nand ginst605 (R2027_U190, R2027_U137, R2027_U28);
  nand ginst606 (R2027_U191, R2027_U124, R2027_U26);
  nand ginst607 (R2027_U192, INSTADDRPOINTER_REG_15__SCAN_IN, R2027_U27);
  nand ginst608 (R2027_U193, INSTADDRPOINTER_REG_14__SCAN_IN, R2027_U108);
  nand ginst609 (R2027_U194, R2027_U138, R2027_U23);
  nand ginst610 (R2027_U195, R2027_U119, R2027_U24);
  nand ginst611 (R2027_U196, INSTADDRPOINTER_REG_13__SCAN_IN, R2027_U25);
  nand ginst612 (R2027_U197, INSTADDRPOINTER_REG_12__SCAN_IN, R2027_U109);
  nand ginst613 (R2027_U198, R2027_U139, R2027_U20);
  nand ginst614 (R2027_U199, R2027_U113, R2027_U21);
  not ginst615 (R2027_U20, INSTADDRPOINTER_REG_12__SCAN_IN);
  nand ginst616 (R2027_U200, INSTADDRPOINTER_REG_11__SCAN_IN, R2027_U22);
  nand ginst617 (R2027_U201, INSTADDRPOINTER_REG_10__SCAN_IN, R2027_U110);
  nand ginst618 (R2027_U202, R2027_U140, R2027_U19);
  not ginst619 (R2027_U21, INSTADDRPOINTER_REG_11__SCAN_IN);
  nand ginst620 (R2027_U22, R2027_U120, R2027_U85);
  not ginst621 (R2027_U23, INSTADDRPOINTER_REG_14__SCAN_IN);
  not ginst622 (R2027_U24, INSTADDRPOINTER_REG_13__SCAN_IN);
  nand ginst623 (R2027_U25, R2027_U113, R2027_U86);
  not ginst624 (R2027_U26, INSTADDRPOINTER_REG_15__SCAN_IN);
  nand ginst625 (R2027_U27, R2027_U119, R2027_U87);
  not ginst626 (R2027_U28, INSTADDRPOINTER_REG_16__SCAN_IN);
  not ginst627 (R2027_U29, INSTADDRPOINTER_REG_18__SCAN_IN);
  not ginst628 (R2027_U30, INSTADDRPOINTER_REG_17__SCAN_IN);
  nand ginst629 (R2027_U31, R2027_U124, R2027_U88);
  not ginst630 (R2027_U32, INSTADDRPOINTER_REG_20__SCAN_IN);
  not ginst631 (R2027_U33, INSTADDRPOINTER_REG_19__SCAN_IN);
  nand ginst632 (R2027_U34, R2027_U117, R2027_U89);
  not ginst633 (R2027_U35, INSTADDRPOINTER_REG_21__SCAN_IN);
  nand ginst634 (R2027_U36, R2027_U114, R2027_U90);
  not ginst635 (R2027_U37, INSTADDRPOINTER_REG_22__SCAN_IN);
  not ginst636 (R2027_U38, INSTADDRPOINTER_REG_24__SCAN_IN);
  not ginst637 (R2027_U39, INSTADDRPOINTER_REG_23__SCAN_IN);
  nand ginst638 (R2027_U40, R2027_U121, R2027_U91);
  not ginst639 (R2027_U41, INSTADDRPOINTER_REG_26__SCAN_IN);
  not ginst640 (R2027_U42, INSTADDRPOINTER_REG_25__SCAN_IN);
  nand ginst641 (R2027_U43, R2027_U115, R2027_U92);
  not ginst642 (R2027_U44, INSTADDRPOINTER_REG_27__SCAN_IN);
  not ginst643 (R2027_U45, INSTADDRPOINTER_REG_28__SCAN_IN);
  nand ginst644 (R2027_U46, R2027_U116, R2027_U93);
  not ginst645 (R2027_U47, INSTADDRPOINTER_REG_29__SCAN_IN);
  nand ginst646 (R2027_U48, R2027_U122, R2027_U94);
  nand ginst647 (R2027_U49, INSTADDRPOINTER_REG_29__SCAN_IN, R2027_U123);
  not ginst648 (R2027_U5, INSTADDRPOINTER_REG_0__SCAN_IN);
  not ginst649 (R2027_U50, INSTADDRPOINTER_REG_30__SCAN_IN);
  nand ginst650 (R2027_U51, R2027_U141, R2027_U142);
  nand ginst651 (R2027_U52, R2027_U143, R2027_U144);
  nand ginst652 (R2027_U53, R2027_U145, R2027_U146);
  nand ginst653 (R2027_U54, R2027_U147, R2027_U148);
  nand ginst654 (R2027_U55, R2027_U149, R2027_U150);
  nand ginst655 (R2027_U56, R2027_U151, R2027_U152);
  nand ginst656 (R2027_U57, R2027_U153, R2027_U154);
  nand ginst657 (R2027_U58, R2027_U155, R2027_U156);
  nand ginst658 (R2027_U59, R2027_U157, R2027_U158);
  not ginst659 (R2027_U6, INSTADDRPOINTER_REG_2__SCAN_IN);
  nand ginst660 (R2027_U60, R2027_U159, R2027_U160);
  nand ginst661 (R2027_U61, R2027_U161, R2027_U162);
  nand ginst662 (R2027_U62, R2027_U163, R2027_U164);
  nand ginst663 (R2027_U63, R2027_U165, R2027_U166);
  nand ginst664 (R2027_U64, R2027_U167, R2027_U168);
  nand ginst665 (R2027_U65, R2027_U169, R2027_U170);
  nand ginst666 (R2027_U66, R2027_U171, R2027_U172);
  nand ginst667 (R2027_U67, R2027_U173, R2027_U174);
  nand ginst668 (R2027_U68, R2027_U175, R2027_U176);
  nand ginst669 (R2027_U69, R2027_U177, R2027_U178);
  not ginst670 (R2027_U7, INSTADDRPOINTER_REG_1__SCAN_IN);
  nand ginst671 (R2027_U70, R2027_U179, R2027_U180);
  nand ginst672 (R2027_U71, R2027_U181, R2027_U182);
  nand ginst673 (R2027_U72, R2027_U183, R2027_U184);
  nand ginst674 (R2027_U73, R2027_U185, R2027_U186);
  nand ginst675 (R2027_U74, R2027_U187, R2027_U188);
  nand ginst676 (R2027_U75, R2027_U189, R2027_U190);
  nand ginst677 (R2027_U76, R2027_U191, R2027_U192);
  nand ginst678 (R2027_U77, R2027_U193, R2027_U194);
  nand ginst679 (R2027_U78, R2027_U195, R2027_U196);
  nand ginst680 (R2027_U79, R2027_U197, R2027_U198);
  not ginst681 (R2027_U8, INSTADDRPOINTER_REG_4__SCAN_IN);
  nand ginst682 (R2027_U80, R2027_U199, R2027_U200);
  nand ginst683 (R2027_U81, R2027_U201, R2027_U202);
  and ginst684 (R2027_U82, INSTADDRPOINTER_REG_3__SCAN_IN, INSTADDRPOINTER_REG_4__SCAN_IN);
  and ginst685 (R2027_U83, INSTADDRPOINTER_REG_5__SCAN_IN, INSTADDRPOINTER_REG_6__SCAN_IN);
  and ginst686 (R2027_U84, INSTADDRPOINTER_REG_7__SCAN_IN, INSTADDRPOINTER_REG_8__SCAN_IN);
  and ginst687 (R2027_U85, INSTADDRPOINTER_REG_9__SCAN_IN, INSTADDRPOINTER_REG_10__SCAN_IN);
  and ginst688 (R2027_U86, INSTADDRPOINTER_REG_11__SCAN_IN, INSTADDRPOINTER_REG_12__SCAN_IN);
  and ginst689 (R2027_U87, INSTADDRPOINTER_REG_13__SCAN_IN, INSTADDRPOINTER_REG_14__SCAN_IN);
  and ginst690 (R2027_U88, INSTADDRPOINTER_REG_15__SCAN_IN, INSTADDRPOINTER_REG_16__SCAN_IN);
  and ginst691 (R2027_U89, INSTADDRPOINTER_REG_17__SCAN_IN, INSTADDRPOINTER_REG_18__SCAN_IN);
  not ginst692 (R2027_U9, INSTADDRPOINTER_REG_3__SCAN_IN);
  and ginst693 (R2027_U90, INSTADDRPOINTER_REG_19__SCAN_IN, INSTADDRPOINTER_REG_20__SCAN_IN);
  and ginst694 (R2027_U91, INSTADDRPOINTER_REG_21__SCAN_IN, INSTADDRPOINTER_REG_22__SCAN_IN);
  and ginst695 (R2027_U92, INSTADDRPOINTER_REG_23__SCAN_IN, INSTADDRPOINTER_REG_24__SCAN_IN);
  and ginst696 (R2027_U93, INSTADDRPOINTER_REG_25__SCAN_IN, INSTADDRPOINTER_REG_26__SCAN_IN);
  and ginst697 (R2027_U94, INSTADDRPOINTER_REG_27__SCAN_IN, INSTADDRPOINTER_REG_28__SCAN_IN);
  nand ginst698 (R2027_U95, INSTADDRPOINTER_REG_7__SCAN_IN, R2027_U118);
  nand ginst699 (R2027_U96, INSTADDRPOINTER_REG_5__SCAN_IN, R2027_U112);
  nand ginst700 (R2027_U97, INSTADDRPOINTER_REG_3__SCAN_IN, R2027_U111);
  not ginst701 (R2027_U98, INSTADDRPOINTER_REG_31__SCAN_IN);
  nand ginst702 (R2027_U99, INSTADDRPOINTER_REG_30__SCAN_IN, R2027_U128);
  nand ginst703 (R2096_U10, REIP_REG_4__SCAN_IN, R2096_U95);
  not ginst704 (R2096_U100, R2096_U19);
  not ginst705 (R2096_U101, R2096_U20);
  not ginst706 (R2096_U102, R2096_U22);
  not ginst707 (R2096_U103, R2096_U24);
  not ginst708 (R2096_U104, R2096_U26);
  not ginst709 (R2096_U105, R2096_U28);
  not ginst710 (R2096_U106, R2096_U30);
  not ginst711 (R2096_U107, R2096_U32);
  not ginst712 (R2096_U108, R2096_U34);
  not ginst713 (R2096_U109, R2096_U36);
  not ginst714 (R2096_U11, REIP_REG_5__SCAN_IN);
  not ginst715 (R2096_U110, R2096_U38);
  not ginst716 (R2096_U111, R2096_U40);
  not ginst717 (R2096_U112, R2096_U42);
  not ginst718 (R2096_U113, R2096_U44);
  not ginst719 (R2096_U114, R2096_U46);
  not ginst720 (R2096_U115, R2096_U48);
  not ginst721 (R2096_U116, R2096_U50);
  not ginst722 (R2096_U117, R2096_U52);
  not ginst723 (R2096_U118, R2096_U54);
  not ginst724 (R2096_U119, R2096_U56);
  nand ginst725 (R2096_U12, REIP_REG_5__SCAN_IN, R2096_U96);
  not ginst726 (R2096_U120, R2096_U58);
  not ginst727 (R2096_U121, R2096_U60);
  not ginst728 (R2096_U122, R2096_U93);
  nand ginst729 (R2096_U123, REIP_REG_9__SCAN_IN, R2096_U19);
  nand ginst730 (R2096_U124, R2096_U100, R2096_U18);
  nand ginst731 (R2096_U125, REIP_REG_8__SCAN_IN, R2096_U16);
  nand ginst732 (R2096_U126, R2096_U17, R2096_U99);
  nand ginst733 (R2096_U127, REIP_REG_7__SCAN_IN, R2096_U14);
  nand ginst734 (R2096_U128, R2096_U15, R2096_U98);
  nand ginst735 (R2096_U129, REIP_REG_6__SCAN_IN, R2096_U12);
  not ginst736 (R2096_U13, REIP_REG_6__SCAN_IN);
  nand ginst737 (R2096_U130, R2096_U13, R2096_U97);
  nand ginst738 (R2096_U131, REIP_REG_5__SCAN_IN, R2096_U10);
  nand ginst739 (R2096_U132, R2096_U11, R2096_U96);
  nand ginst740 (R2096_U133, REIP_REG_4__SCAN_IN, R2096_U8);
  nand ginst741 (R2096_U134, R2096_U9, R2096_U95);
  nand ginst742 (R2096_U135, REIP_REG_3__SCAN_IN, R2096_U6);
  nand ginst743 (R2096_U136, R2096_U7, R2096_U94);
  nand ginst744 (R2096_U137, REIP_REG_31__SCAN_IN, R2096_U93);
  nand ginst745 (R2096_U138, R2096_U122, R2096_U92);
  nand ginst746 (R2096_U139, REIP_REG_30__SCAN_IN, R2096_U60);
  nand ginst747 (R2096_U14, REIP_REG_6__SCAN_IN, R2096_U97);
  nand ginst748 (R2096_U140, R2096_U121, R2096_U61);
  nand ginst749 (R2096_U141, REIP_REG_2__SCAN_IN, R2096_U4);
  nand ginst750 (R2096_U142, REIP_REG_1__SCAN_IN, R2096_U5);
  nand ginst751 (R2096_U143, REIP_REG_29__SCAN_IN, R2096_U58);
  nand ginst752 (R2096_U144, R2096_U120, R2096_U59);
  nand ginst753 (R2096_U145, REIP_REG_28__SCAN_IN, R2096_U56);
  nand ginst754 (R2096_U146, R2096_U119, R2096_U57);
  nand ginst755 (R2096_U147, REIP_REG_27__SCAN_IN, R2096_U54);
  nand ginst756 (R2096_U148, R2096_U118, R2096_U55);
  nand ginst757 (R2096_U149, REIP_REG_26__SCAN_IN, R2096_U52);
  not ginst758 (R2096_U15, REIP_REG_7__SCAN_IN);
  nand ginst759 (R2096_U150, R2096_U117, R2096_U53);
  nand ginst760 (R2096_U151, REIP_REG_25__SCAN_IN, R2096_U50);
  nand ginst761 (R2096_U152, R2096_U116, R2096_U51);
  nand ginst762 (R2096_U153, REIP_REG_24__SCAN_IN, R2096_U48);
  nand ginst763 (R2096_U154, R2096_U115, R2096_U49);
  nand ginst764 (R2096_U155, REIP_REG_23__SCAN_IN, R2096_U46);
  nand ginst765 (R2096_U156, R2096_U114, R2096_U47);
  nand ginst766 (R2096_U157, REIP_REG_22__SCAN_IN, R2096_U44);
  nand ginst767 (R2096_U158, R2096_U113, R2096_U45);
  nand ginst768 (R2096_U159, REIP_REG_21__SCAN_IN, R2096_U42);
  nand ginst769 (R2096_U16, REIP_REG_7__SCAN_IN, R2096_U98);
  nand ginst770 (R2096_U160, R2096_U112, R2096_U43);
  nand ginst771 (R2096_U161, REIP_REG_20__SCAN_IN, R2096_U40);
  nand ginst772 (R2096_U162, R2096_U111, R2096_U41);
  nand ginst773 (R2096_U163, REIP_REG_19__SCAN_IN, R2096_U38);
  nand ginst774 (R2096_U164, R2096_U110, R2096_U39);
  nand ginst775 (R2096_U165, REIP_REG_18__SCAN_IN, R2096_U36);
  nand ginst776 (R2096_U166, R2096_U109, R2096_U37);
  nand ginst777 (R2096_U167, REIP_REG_17__SCAN_IN, R2096_U34);
  nand ginst778 (R2096_U168, R2096_U108, R2096_U35);
  nand ginst779 (R2096_U169, REIP_REG_16__SCAN_IN, R2096_U32);
  not ginst780 (R2096_U17, REIP_REG_8__SCAN_IN);
  nand ginst781 (R2096_U170, R2096_U107, R2096_U33);
  nand ginst782 (R2096_U171, REIP_REG_15__SCAN_IN, R2096_U30);
  nand ginst783 (R2096_U172, R2096_U106, R2096_U31);
  nand ginst784 (R2096_U173, REIP_REG_14__SCAN_IN, R2096_U28);
  nand ginst785 (R2096_U174, R2096_U105, R2096_U29);
  nand ginst786 (R2096_U175, REIP_REG_13__SCAN_IN, R2096_U26);
  nand ginst787 (R2096_U176, R2096_U104, R2096_U27);
  nand ginst788 (R2096_U177, REIP_REG_12__SCAN_IN, R2096_U24);
  nand ginst789 (R2096_U178, R2096_U103, R2096_U25);
  nand ginst790 (R2096_U179, REIP_REG_11__SCAN_IN, R2096_U22);
  not ginst791 (R2096_U18, REIP_REG_9__SCAN_IN);
  nand ginst792 (R2096_U180, R2096_U102, R2096_U23);
  nand ginst793 (R2096_U181, REIP_REG_10__SCAN_IN, R2096_U20);
  nand ginst794 (R2096_U182, R2096_U101, R2096_U21);
  nand ginst795 (R2096_U19, REIP_REG_8__SCAN_IN, R2096_U99);
  nand ginst796 (R2096_U20, REIP_REG_9__SCAN_IN, R2096_U100);
  not ginst797 (R2096_U21, REIP_REG_10__SCAN_IN);
  nand ginst798 (R2096_U22, REIP_REG_10__SCAN_IN, R2096_U101);
  not ginst799 (R2096_U23, REIP_REG_11__SCAN_IN);
  nand ginst800 (R2096_U24, REIP_REG_11__SCAN_IN, R2096_U102);
  not ginst801 (R2096_U25, REIP_REG_12__SCAN_IN);
  nand ginst802 (R2096_U26, REIP_REG_12__SCAN_IN, R2096_U103);
  not ginst803 (R2096_U27, REIP_REG_13__SCAN_IN);
  nand ginst804 (R2096_U28, REIP_REG_13__SCAN_IN, R2096_U104);
  not ginst805 (R2096_U29, REIP_REG_14__SCAN_IN);
  nand ginst806 (R2096_U30, REIP_REG_14__SCAN_IN, R2096_U105);
  not ginst807 (R2096_U31, REIP_REG_15__SCAN_IN);
  nand ginst808 (R2096_U32, REIP_REG_15__SCAN_IN, R2096_U106);
  not ginst809 (R2096_U33, REIP_REG_16__SCAN_IN);
  nand ginst810 (R2096_U34, REIP_REG_16__SCAN_IN, R2096_U107);
  not ginst811 (R2096_U35, REIP_REG_17__SCAN_IN);
  nand ginst812 (R2096_U36, REIP_REG_17__SCAN_IN, R2096_U108);
  not ginst813 (R2096_U37, REIP_REG_18__SCAN_IN);
  nand ginst814 (R2096_U38, REIP_REG_18__SCAN_IN, R2096_U109);
  not ginst815 (R2096_U39, REIP_REG_19__SCAN_IN);
  not ginst816 (R2096_U4, REIP_REG_1__SCAN_IN);
  nand ginst817 (R2096_U40, REIP_REG_19__SCAN_IN, R2096_U110);
  not ginst818 (R2096_U41, REIP_REG_20__SCAN_IN);
  nand ginst819 (R2096_U42, REIP_REG_20__SCAN_IN, R2096_U111);
  not ginst820 (R2096_U43, REIP_REG_21__SCAN_IN);
  nand ginst821 (R2096_U44, REIP_REG_21__SCAN_IN, R2096_U112);
  not ginst822 (R2096_U45, REIP_REG_22__SCAN_IN);
  nand ginst823 (R2096_U46, REIP_REG_22__SCAN_IN, R2096_U113);
  not ginst824 (R2096_U47, REIP_REG_23__SCAN_IN);
  nand ginst825 (R2096_U48, REIP_REG_23__SCAN_IN, R2096_U114);
  not ginst826 (R2096_U49, REIP_REG_24__SCAN_IN);
  not ginst827 (R2096_U5, REIP_REG_2__SCAN_IN);
  nand ginst828 (R2096_U50, REIP_REG_24__SCAN_IN, R2096_U115);
  not ginst829 (R2096_U51, REIP_REG_25__SCAN_IN);
  nand ginst830 (R2096_U52, REIP_REG_25__SCAN_IN, R2096_U116);
  not ginst831 (R2096_U53, REIP_REG_26__SCAN_IN);
  nand ginst832 (R2096_U54, REIP_REG_26__SCAN_IN, R2096_U117);
  not ginst833 (R2096_U55, REIP_REG_27__SCAN_IN);
  nand ginst834 (R2096_U56, REIP_REG_27__SCAN_IN, R2096_U118);
  not ginst835 (R2096_U57, REIP_REG_28__SCAN_IN);
  nand ginst836 (R2096_U58, REIP_REG_28__SCAN_IN, R2096_U119);
  not ginst837 (R2096_U59, REIP_REG_29__SCAN_IN);
  nand ginst838 (R2096_U6, REIP_REG_1__SCAN_IN, REIP_REG_2__SCAN_IN);
  nand ginst839 (R2096_U60, REIP_REG_29__SCAN_IN, R2096_U120);
  not ginst840 (R2096_U61, REIP_REG_30__SCAN_IN);
  nand ginst841 (R2096_U62, R2096_U123, R2096_U124);
  nand ginst842 (R2096_U63, R2096_U125, R2096_U126);
  nand ginst843 (R2096_U64, R2096_U127, R2096_U128);
  nand ginst844 (R2096_U65, R2096_U129, R2096_U130);
  nand ginst845 (R2096_U66, R2096_U131, R2096_U132);
  nand ginst846 (R2096_U67, R2096_U133, R2096_U134);
  nand ginst847 (R2096_U68, R2096_U135, R2096_U136);
  nand ginst848 (R2096_U69, R2096_U137, R2096_U138);
  not ginst849 (R2096_U7, REIP_REG_3__SCAN_IN);
  nand ginst850 (R2096_U70, R2096_U139, R2096_U140);
  nand ginst851 (R2096_U71, R2096_U141, R2096_U142);
  nand ginst852 (R2096_U72, R2096_U143, R2096_U144);
  nand ginst853 (R2096_U73, R2096_U145, R2096_U146);
  nand ginst854 (R2096_U74, R2096_U147, R2096_U148);
  nand ginst855 (R2096_U75, R2096_U149, R2096_U150);
  nand ginst856 (R2096_U76, R2096_U151, R2096_U152);
  nand ginst857 (R2096_U77, R2096_U153, R2096_U154);
  nand ginst858 (R2096_U78, R2096_U155, R2096_U156);
  nand ginst859 (R2096_U79, R2096_U157, R2096_U158);
  nand ginst860 (R2096_U8, REIP_REG_3__SCAN_IN, R2096_U94);
  nand ginst861 (R2096_U80, R2096_U159, R2096_U160);
  nand ginst862 (R2096_U81, R2096_U161, R2096_U162);
  nand ginst863 (R2096_U82, R2096_U163, R2096_U164);
  nand ginst864 (R2096_U83, R2096_U165, R2096_U166);
  nand ginst865 (R2096_U84, R2096_U167, R2096_U168);
  nand ginst866 (R2096_U85, R2096_U169, R2096_U170);
  nand ginst867 (R2096_U86, R2096_U171, R2096_U172);
  nand ginst868 (R2096_U87, R2096_U173, R2096_U174);
  nand ginst869 (R2096_U88, R2096_U175, R2096_U176);
  nand ginst870 (R2096_U89, R2096_U177, R2096_U178);
  not ginst871 (R2096_U9, REIP_REG_4__SCAN_IN);
  nand ginst872 (R2096_U90, R2096_U179, R2096_U180);
  nand ginst873 (R2096_U91, R2096_U181, R2096_U182);
  not ginst874 (R2096_U92, REIP_REG_31__SCAN_IN);
  nand ginst875 (R2096_U93, REIP_REG_30__SCAN_IN, R2096_U121);
  not ginst876 (R2096_U94, R2096_U6);
  not ginst877 (R2096_U95, R2096_U8);
  not ginst878 (R2096_U96, R2096_U10);
  not ginst879 (R2096_U97, R2096_U12);
  not ginst880 (R2096_U98, R2096_U14);
  not ginst881 (R2096_U99, R2096_U16);
  nand ginst882 (R2099_U10, R2099_U159, R2099_U91);
  not ginst883 (R2099_U100, U2710);
  not ginst884 (R2099_U101, U2709);
  not ginst885 (R2099_U102, U2708);
  not ginst886 (R2099_U103, U2707);
  not ginst887 (R2099_U104, U2706);
  not ginst888 (R2099_U105, U2705);
  not ginst889 (R2099_U106, U2704);
  not ginst890 (R2099_U107, U2703);
  not ginst891 (R2099_U108, U2701);
  nand ginst892 (R2099_U109, R2099_U159, R2099_U27);
  nand ginst893 (R2099_U11, R2099_U161, R2099_U92);
  nand ginst894 (R2099_U110, R2099_U157, R2099_U28);
  nand ginst895 (R2099_U111, R2099_U155, R2099_U30);
  nand ginst896 (R2099_U112, R2099_U137, R2099_U35);
  not ginst897 (R2099_U113, U2682);
  not ginst898 (R2099_U114, U2683);
  not ginst899 (R2099_U115, U2684);
  not ginst900 (R2099_U116, U2685);
  not ginst901 (R2099_U117, U2686);
  not ginst902 (R2099_U118, U2687);
  not ginst903 (R2099_U119, U2688);
  nand ginst904 (R2099_U12, R2099_U163, R2099_U93);
  not ginst905 (R2099_U120, U2689);
  not ginst906 (R2099_U121, U2690);
  not ginst907 (R2099_U122, U2691);
  not ginst908 (R2099_U123, U2692);
  not ginst909 (R2099_U124, U2700);
  not ginst910 (R2099_U125, U2699);
  not ginst911 (R2099_U126, U2698);
  not ginst912 (R2099_U127, U2697);
  not ginst913 (R2099_U128, U2696);
  not ginst914 (R2099_U129, U2695);
  nand ginst915 (R2099_U13, R2099_U165, R2099_U94);
  not ginst916 (R2099_U130, U2694);
  not ginst917 (R2099_U131, U2693);
  not ginst918 (R2099_U132, U2680);
  not ginst919 (R2099_U133, U2681);
  not ginst920 (R2099_U134, U2679);
  nand ginst921 (R2099_U135, R2099_U180, R2099_U96);
  nand ginst922 (R2099_U136, R2099_U180, R2099_U44);
  nand ginst923 (R2099_U137, R2099_U151, R2099_U152);
  and ginst924 (R2099_U138, R2099_U296, R2099_U297);
  and ginst925 (R2099_U139, R2099_U318, R2099_U319);
  nand ginst926 (R2099_U14, R2099_U167, R2099_U95);
  nand ginst927 (R2099_U140, R2099_U147, R2099_U148);
  nand ginst928 (R2099_U141, R2099_U167, R2099_U56);
  nand ginst929 (R2099_U142, R2099_U165, R2099_U58);
  nand ginst930 (R2099_U143, R2099_U163, R2099_U60);
  nand ginst931 (R2099_U144, R2099_U161, R2099_U62);
  not ginst932 (R2099_U145, R2099_U135);
  or ginst933 (R2099_U146, U4177, U4178);
  nand ginst934 (R2099_U147, R2099_U146, R2099_U32);
  nand ginst935 (R2099_U148, U4177, U4178);
  not ginst936 (R2099_U149, R2099_U140);
  nand ginst937 (R2099_U15, R2099_U169, R2099_U55);
  nand ginst938 (R2099_U150, R2099_U190, R2099_U6);
  nand ginst939 (R2099_U151, R2099_U140, R2099_U150);
  nand ginst940 (R2099_U152, R2099_U33, U2678);
  not ginst941 (R2099_U153, R2099_U137);
  not ginst942 (R2099_U154, R2099_U112);
  not ginst943 (R2099_U155, R2099_U7);
  not ginst944 (R2099_U156, R2099_U111);
  not ginst945 (R2099_U157, R2099_U8);
  not ginst946 (R2099_U158, R2099_U110);
  not ginst947 (R2099_U159, R2099_U9);
  nand ginst948 (R2099_U16, R2099_U170, R2099_U54);
  not ginst949 (R2099_U160, R2099_U109);
  not ginst950 (R2099_U161, R2099_U10);
  not ginst951 (R2099_U162, R2099_U144);
  not ginst952 (R2099_U163, R2099_U11);
  not ginst953 (R2099_U164, R2099_U143);
  not ginst954 (R2099_U165, R2099_U12);
  not ginst955 (R2099_U166, R2099_U142);
  not ginst956 (R2099_U167, R2099_U13);
  not ginst957 (R2099_U168, R2099_U141);
  not ginst958 (R2099_U169, R2099_U14);
  nand ginst959 (R2099_U17, R2099_U171, R2099_U53);
  not ginst960 (R2099_U170, R2099_U15);
  not ginst961 (R2099_U171, R2099_U16);
  not ginst962 (R2099_U172, R2099_U17);
  not ginst963 (R2099_U173, R2099_U18);
  not ginst964 (R2099_U174, R2099_U19);
  not ginst965 (R2099_U175, R2099_U20);
  not ginst966 (R2099_U176, R2099_U21);
  not ginst967 (R2099_U177, R2099_U22);
  not ginst968 (R2099_U178, R2099_U23);
  not ginst969 (R2099_U179, R2099_U24);
  nand ginst970 (R2099_U18, R2099_U172, R2099_U52);
  not ginst971 (R2099_U180, R2099_U25);
  not ginst972 (R2099_U181, R2099_U136);
  nand ginst973 (R2099_U182, R2099_U99, U4178);
  nand ginst974 (R2099_U183, R2099_U4, U2702);
  not ginst975 (R2099_U184, R2099_U27);
  nand ginst976 (R2099_U185, R2099_U100, U4178);
  nand ginst977 (R2099_U186, R2099_U4, U2710);
  not ginst978 (R2099_U187, R2099_U32);
  nand ginst979 (R2099_U188, R2099_U101, U4178);
  nand ginst980 (R2099_U189, R2099_U4, U2709);
  nand ginst981 (R2099_U19, R2099_U173, R2099_U51);
  not ginst982 (R2099_U190, R2099_U33);
  nand ginst983 (R2099_U191, R2099_U102, U4178);
  nand ginst984 (R2099_U192, R2099_U4, U2708);
  not ginst985 (R2099_U193, R2099_U35);
  nand ginst986 (R2099_U194, R2099_U103, U4178);
  nand ginst987 (R2099_U195, R2099_U4, U2707);
  not ginst988 (R2099_U196, R2099_U34);
  nand ginst989 (R2099_U197, R2099_U104, U4178);
  nand ginst990 (R2099_U198, R2099_U4, U2706);
  not ginst991 (R2099_U199, R2099_U30);
  nand ginst992 (R2099_U20, R2099_U174, R2099_U50);
  nand ginst993 (R2099_U200, R2099_U105, U4178);
  nand ginst994 (R2099_U201, R2099_U4, U2705);
  not ginst995 (R2099_U202, R2099_U31);
  nand ginst996 (R2099_U203, R2099_U106, U4178);
  nand ginst997 (R2099_U204, R2099_U4, U2704);
  not ginst998 (R2099_U205, R2099_U28);
  nand ginst999 (R2099_U206, R2099_U107, U4178);
  nand ginst1000 (R2099_U207, R2099_U4, U2703);
  not ginst1001 (R2099_U208, R2099_U29);
  nand ginst1002 (R2099_U209, R2099_U108, U4178);
  nand ginst1003 (R2099_U21, R2099_U175, R2099_U49);
  nand ginst1004 (R2099_U210, R2099_U4, U2701);
  not ginst1005 (R2099_U211, R2099_U26);
  nand ginst1006 (R2099_U212, R2099_U160, R2099_U211);
  nand ginst1007 (R2099_U213, R2099_U109, R2099_U26);
  nand ginst1008 (R2099_U214, R2099_U159, R2099_U184);
  nand ginst1009 (R2099_U215, R2099_U27, R2099_U9);
  nand ginst1010 (R2099_U216, R2099_U158, R2099_U208);
  nand ginst1011 (R2099_U217, R2099_U110, R2099_U29);
  nand ginst1012 (R2099_U218, R2099_U157, R2099_U205);
  nand ginst1013 (R2099_U219, R2099_U28, R2099_U8);
  nand ginst1014 (R2099_U22, R2099_U176, R2099_U48);
  nand ginst1015 (R2099_U220, R2099_U156, R2099_U202);
  nand ginst1016 (R2099_U221, R2099_U111, R2099_U31);
  nand ginst1017 (R2099_U222, R2099_U155, R2099_U199);
  nand ginst1018 (R2099_U223, R2099_U30, R2099_U7);
  nand ginst1019 (R2099_U224, R2099_U154, R2099_U196);
  nand ginst1020 (R2099_U225, R2099_U112, R2099_U34);
  nand ginst1021 (R2099_U226, R2099_U113, U4178);
  nand ginst1022 (R2099_U227, R2099_U4, U2682);
  not ginst1023 (R2099_U228, R2099_U45);
  nand ginst1024 (R2099_U229, R2099_U114, U4178);
  nand ginst1025 (R2099_U23, R2099_U177, R2099_U47);
  nand ginst1026 (R2099_U230, R2099_U4, U2683);
  not ginst1027 (R2099_U231, R2099_U46);
  nand ginst1028 (R2099_U232, R2099_U115, U4178);
  nand ginst1029 (R2099_U233, R2099_U4, U2684);
  not ginst1030 (R2099_U234, R2099_U47);
  nand ginst1031 (R2099_U235, R2099_U116, U4178);
  nand ginst1032 (R2099_U236, R2099_U4, U2685);
  not ginst1033 (R2099_U237, R2099_U48);
  nand ginst1034 (R2099_U238, R2099_U117, U4178);
  nand ginst1035 (R2099_U239, R2099_U4, U2686);
  nand ginst1036 (R2099_U24, R2099_U178, R2099_U46);
  not ginst1037 (R2099_U240, R2099_U49);
  nand ginst1038 (R2099_U241, R2099_U118, U4178);
  nand ginst1039 (R2099_U242, R2099_U4, U2687);
  not ginst1040 (R2099_U243, R2099_U50);
  nand ginst1041 (R2099_U244, R2099_U119, U4178);
  nand ginst1042 (R2099_U245, R2099_U4, U2688);
  not ginst1043 (R2099_U246, R2099_U51);
  nand ginst1044 (R2099_U247, R2099_U120, U4178);
  nand ginst1045 (R2099_U248, R2099_U4, U2689);
  not ginst1046 (R2099_U249, R2099_U52);
  nand ginst1047 (R2099_U25, R2099_U179, R2099_U45);
  nand ginst1048 (R2099_U250, R2099_U121, U4178);
  nand ginst1049 (R2099_U251, R2099_U4, U2690);
  not ginst1050 (R2099_U252, R2099_U53);
  nand ginst1051 (R2099_U253, R2099_U122, U4178);
  nand ginst1052 (R2099_U254, R2099_U4, U2691);
  not ginst1053 (R2099_U255, R2099_U54);
  nand ginst1054 (R2099_U256, R2099_U123, U4178);
  nand ginst1055 (R2099_U257, R2099_U4, U2692);
  not ginst1056 (R2099_U258, R2099_U55);
  nand ginst1057 (R2099_U259, R2099_U124, U4178);
  nand ginst1058 (R2099_U26, R2099_U209, R2099_U210);
  nand ginst1059 (R2099_U260, R2099_U4, U2700);
  not ginst1060 (R2099_U261, R2099_U62);
  nand ginst1061 (R2099_U262, R2099_U125, U4178);
  nand ginst1062 (R2099_U263, R2099_U4, U2699);
  not ginst1063 (R2099_U264, R2099_U63);
  nand ginst1064 (R2099_U265, R2099_U126, U4178);
  nand ginst1065 (R2099_U266, R2099_U4, U2698);
  not ginst1066 (R2099_U267, R2099_U60);
  nand ginst1067 (R2099_U268, R2099_U127, U4178);
  nand ginst1068 (R2099_U269, R2099_U4, U2697);
  nand ginst1069 (R2099_U27, R2099_U182, R2099_U183);
  not ginst1070 (R2099_U270, R2099_U61);
  nand ginst1071 (R2099_U271, R2099_U128, U4178);
  nand ginst1072 (R2099_U272, R2099_U4, U2696);
  not ginst1073 (R2099_U273, R2099_U58);
  nand ginst1074 (R2099_U274, R2099_U129, U4178);
  nand ginst1075 (R2099_U275, R2099_U4, U2695);
  not ginst1076 (R2099_U276, R2099_U59);
  nand ginst1077 (R2099_U277, R2099_U130, U4178);
  nand ginst1078 (R2099_U278, R2099_U4, U2694);
  not ginst1079 (R2099_U279, R2099_U56);
  nand ginst1080 (R2099_U28, R2099_U203, R2099_U204);
  nand ginst1081 (R2099_U280, R2099_U131, U4178);
  nand ginst1082 (R2099_U281, R2099_U4, U2693);
  not ginst1083 (R2099_U282, R2099_U57);
  nand ginst1084 (R2099_U283, R2099_U132, U4178);
  nand ginst1085 (R2099_U284, R2099_U4, U2680);
  not ginst1086 (R2099_U285, R2099_U43);
  nand ginst1087 (R2099_U286, R2099_U133, U4178);
  nand ginst1088 (R2099_U287, R2099_U4, U2681);
  not ginst1089 (R2099_U288, R2099_U44);
  nand ginst1090 (R2099_U289, R2099_U134, U4178);
  nand ginst1091 (R2099_U29, R2099_U206, R2099_U207);
  nand ginst1092 (R2099_U290, R2099_U4, U2679);
  not ginst1093 (R2099_U291, R2099_U97);
  nand ginst1094 (R2099_U292, R2099_U145, R2099_U291);
  nand ginst1095 (R2099_U293, R2099_U135, R2099_U97);
  nand ginst1096 (R2099_U294, R2099_U181, R2099_U285);
  nand ginst1097 (R2099_U295, R2099_U136, R2099_U43);
  nand ginst1098 (R2099_U296, R2099_U153, R2099_U193);
  nand ginst1099 (R2099_U297, R2099_U137, R2099_U35);
  nand ginst1100 (R2099_U298, R2099_U180, R2099_U288);
  nand ginst1101 (R2099_U299, R2099_U25, R2099_U44);
  nand ginst1102 (R2099_U30, R2099_U197, R2099_U198);
  nand ginst1103 (R2099_U300, R2099_U179, R2099_U228);
  nand ginst1104 (R2099_U301, R2099_U24, R2099_U45);
  nand ginst1105 (R2099_U302, R2099_U178, R2099_U231);
  nand ginst1106 (R2099_U303, R2099_U23, R2099_U46);
  nand ginst1107 (R2099_U304, R2099_U177, R2099_U234);
  nand ginst1108 (R2099_U305, R2099_U22, R2099_U47);
  nand ginst1109 (R2099_U306, R2099_U176, R2099_U237);
  nand ginst1110 (R2099_U307, R2099_U21, R2099_U48);
  nand ginst1111 (R2099_U308, R2099_U175, R2099_U240);
  nand ginst1112 (R2099_U309, R2099_U20, R2099_U49);
  nand ginst1113 (R2099_U31, R2099_U200, R2099_U201);
  nand ginst1114 (R2099_U310, R2099_U174, R2099_U243);
  nand ginst1115 (R2099_U311, R2099_U19, R2099_U50);
  nand ginst1116 (R2099_U312, R2099_U173, R2099_U246);
  nand ginst1117 (R2099_U313, R2099_U18, R2099_U51);
  nand ginst1118 (R2099_U314, R2099_U172, R2099_U249);
  nand ginst1119 (R2099_U315, R2099_U17, R2099_U52);
  nand ginst1120 (R2099_U316, R2099_U171, R2099_U252);
  nand ginst1121 (R2099_U317, R2099_U16, R2099_U53);
  nand ginst1122 (R2099_U318, R2099_U190, U2678);
  nand ginst1123 (R2099_U319, R2099_U33, R2099_U6);
  nand ginst1124 (R2099_U32, R2099_U185, R2099_U186);
  nand ginst1125 (R2099_U320, R2099_U190, U2678);
  nand ginst1126 (R2099_U321, R2099_U33, R2099_U6);
  nand ginst1127 (R2099_U322, R2099_U320, R2099_U321);
  nand ginst1128 (R2099_U323, R2099_U139, R2099_U140);
  nand ginst1129 (R2099_U324, R2099_U149, R2099_U322);
  nand ginst1130 (R2099_U325, R2099_U170, R2099_U255);
  nand ginst1131 (R2099_U326, R2099_U15, R2099_U54);
  nand ginst1132 (R2099_U327, R2099_U169, R2099_U258);
  nand ginst1133 (R2099_U328, R2099_U14, R2099_U55);
  nand ginst1134 (R2099_U329, R2099_U168, R2099_U282);
  nand ginst1135 (R2099_U33, R2099_U188, R2099_U189);
  nand ginst1136 (R2099_U330, R2099_U141, R2099_U57);
  nand ginst1137 (R2099_U331, R2099_U167, R2099_U279);
  nand ginst1138 (R2099_U332, R2099_U13, R2099_U56);
  nand ginst1139 (R2099_U333, R2099_U166, R2099_U276);
  nand ginst1140 (R2099_U334, R2099_U142, R2099_U59);
  nand ginst1141 (R2099_U335, R2099_U165, R2099_U273);
  nand ginst1142 (R2099_U336, R2099_U12, R2099_U58);
  nand ginst1143 (R2099_U337, R2099_U164, R2099_U270);
  nand ginst1144 (R2099_U338, R2099_U143, R2099_U61);
  nand ginst1145 (R2099_U339, R2099_U163, R2099_U267);
  nand ginst1146 (R2099_U34, R2099_U194, R2099_U195);
  nand ginst1147 (R2099_U340, R2099_U11, R2099_U60);
  nand ginst1148 (R2099_U341, R2099_U162, R2099_U264);
  nand ginst1149 (R2099_U342, R2099_U144, R2099_U63);
  nand ginst1150 (R2099_U343, R2099_U161, R2099_U261);
  nand ginst1151 (R2099_U344, R2099_U10, R2099_U62);
  nand ginst1152 (R2099_U345, R2099_U4, U4177);
  nand ginst1153 (R2099_U346, R2099_U5, U4178);
  not ginst1154 (R2099_U347, R2099_U98);
  nand ginst1155 (R2099_U348, R2099_U32, R2099_U347);
  nand ginst1156 (R2099_U349, R2099_U187, R2099_U98);
  nand ginst1157 (R2099_U35, R2099_U191, R2099_U192);
  nand ginst1158 (R2099_U36, R2099_U212, R2099_U213);
  nand ginst1159 (R2099_U37, R2099_U214, R2099_U215);
  nand ginst1160 (R2099_U38, R2099_U216, R2099_U217);
  nand ginst1161 (R2099_U39, R2099_U218, R2099_U219);
  not ginst1162 (R2099_U4, U4178);
  nand ginst1163 (R2099_U40, R2099_U220, R2099_U221);
  nand ginst1164 (R2099_U41, R2099_U222, R2099_U223);
  nand ginst1165 (R2099_U42, R2099_U224, R2099_U225);
  nand ginst1166 (R2099_U43, R2099_U283, R2099_U284);
  nand ginst1167 (R2099_U44, R2099_U286, R2099_U287);
  nand ginst1168 (R2099_U45, R2099_U226, R2099_U227);
  nand ginst1169 (R2099_U46, R2099_U229, R2099_U230);
  nand ginst1170 (R2099_U47, R2099_U232, R2099_U233);
  nand ginst1171 (R2099_U48, R2099_U235, R2099_U236);
  nand ginst1172 (R2099_U49, R2099_U238, R2099_U239);
  not ginst1173 (R2099_U5, U4177);
  nand ginst1174 (R2099_U50, R2099_U241, R2099_U242);
  nand ginst1175 (R2099_U51, R2099_U244, R2099_U245);
  nand ginst1176 (R2099_U52, R2099_U247, R2099_U248);
  nand ginst1177 (R2099_U53, R2099_U250, R2099_U251);
  nand ginst1178 (R2099_U54, R2099_U253, R2099_U254);
  nand ginst1179 (R2099_U55, R2099_U256, R2099_U257);
  nand ginst1180 (R2099_U56, R2099_U277, R2099_U278);
  nand ginst1181 (R2099_U57, R2099_U280, R2099_U281);
  nand ginst1182 (R2099_U58, R2099_U271, R2099_U272);
  nand ginst1183 (R2099_U59, R2099_U274, R2099_U275);
  not ginst1184 (R2099_U6, U2678);
  nand ginst1185 (R2099_U60, R2099_U265, R2099_U266);
  nand ginst1186 (R2099_U61, R2099_U268, R2099_U269);
  nand ginst1187 (R2099_U62, R2099_U259, R2099_U260);
  nand ginst1188 (R2099_U63, R2099_U262, R2099_U263);
  nand ginst1189 (R2099_U64, R2099_U292, R2099_U293);
  nand ginst1190 (R2099_U65, R2099_U294, R2099_U295);
  nand ginst1191 (R2099_U66, R2099_U298, R2099_U299);
  nand ginst1192 (R2099_U67, R2099_U300, R2099_U301);
  nand ginst1193 (R2099_U68, R2099_U302, R2099_U303);
  nand ginst1194 (R2099_U69, R2099_U304, R2099_U305);
  nand ginst1195 (R2099_U7, R2099_U137, R2099_U88);
  nand ginst1196 (R2099_U70, R2099_U306, R2099_U307);
  nand ginst1197 (R2099_U71, R2099_U308, R2099_U309);
  nand ginst1198 (R2099_U72, R2099_U310, R2099_U311);
  nand ginst1199 (R2099_U73, R2099_U312, R2099_U313);
  nand ginst1200 (R2099_U74, R2099_U314, R2099_U315);
  nand ginst1201 (R2099_U75, R2099_U316, R2099_U317);
  nand ginst1202 (R2099_U76, R2099_U325, R2099_U326);
  nand ginst1203 (R2099_U77, R2099_U327, R2099_U328);
  nand ginst1204 (R2099_U78, R2099_U329, R2099_U330);
  nand ginst1205 (R2099_U79, R2099_U331, R2099_U332);
  nand ginst1206 (R2099_U8, R2099_U155, R2099_U89);
  nand ginst1207 (R2099_U80, R2099_U333, R2099_U334);
  nand ginst1208 (R2099_U81, R2099_U335, R2099_U336);
  nand ginst1209 (R2099_U82, R2099_U337, R2099_U338);
  nand ginst1210 (R2099_U83, R2099_U339, R2099_U340);
  nand ginst1211 (R2099_U84, R2099_U341, R2099_U342);
  nand ginst1212 (R2099_U85, R2099_U343, R2099_U344);
  nand ginst1213 (R2099_U86, R2099_U348, R2099_U349);
  nand ginst1214 (R2099_U87, R2099_U323, R2099_U324);
  and ginst1215 (R2099_U88, R2099_U34, R2099_U35);
  and ginst1216 (R2099_U89, R2099_U30, R2099_U31);
  nand ginst1217 (R2099_U9, R2099_U157, R2099_U90);
  and ginst1218 (R2099_U90, R2099_U28, R2099_U29);
  and ginst1219 (R2099_U91, R2099_U26, R2099_U27);
  and ginst1220 (R2099_U92, R2099_U62, R2099_U63);
  and ginst1221 (R2099_U93, R2099_U60, R2099_U61);
  and ginst1222 (R2099_U94, R2099_U58, R2099_U59);
  and ginst1223 (R2099_U95, R2099_U56, R2099_U57);
  and ginst1224 (R2099_U96, R2099_U43, R2099_U44);
  nand ginst1225 (R2099_U97, R2099_U289, R2099_U290);
  nand ginst1226 (R2099_U98, R2099_U345, R2099_U346);
  not ginst1227 (R2099_U99, U2702);
  and ginst1228 (R2144_U10, R2144_U212, R2144_U213, R2144_U82);
  nand ginst1229 (R2144_U100, R2144_U28, U2751);
  not ginst1230 (R2144_U101, R2144_U24);
  not ginst1231 (R2144_U102, R2144_U81);
  nand ginst1232 (R2144_U103, R2144_U181, U2745);
  nand ginst1233 (R2144_U104, R2144_U166, R2144_U167, R2144_U17);
  nand ginst1234 (R2144_U105, R2144_U174, R2144_U175, R2144_U20);
  nand ginst1235 (R2144_U106, R2144_U18, R2144_U200, R2144_U201);
  not ginst1236 (R2144_U107, R2144_U21);
  not ginst1237 (R2144_U108, R2144_U23);
  nand ginst1238 (R2144_U109, R2144_U13, R2144_U193, R2144_U194);
  nand ginst1239 (R2144_U11, R2144_U144, R2144_U146);
  nand ginst1240 (R2144_U110, R2144_U16, R2144_U195, R2144_U196);
  nand ginst1241 (R2144_U111, R2144_U199, U2749);
  nand ginst1242 (R2144_U112, R2144_U15, R2144_U188, R2144_U189);
  nand ginst1243 (R2144_U113, R2144_U192, U2752);
  nand ginst1244 (R2144_U114, R2144_U14, R2144_U187);
  nand ginst1245 (R2144_U115, R2144_U112, U2355);
  nand ginst1246 (R2144_U116, R2144_U184, U2750);
  nand ginst1247 (R2144_U117, R2144_U155, R2144_U157);
  nand ginst1248 (R2144_U118, R2144_U117, R2144_U51);
  not ginst1249 (R2144_U119, R2144_U84);
  not ginst1250 (R2144_U12, U2355);
  not ginst1251 (R2144_U120, R2144_U19);
  not ginst1252 (R2144_U121, R2144_U79);
  not ginst1253 (R2144_U122, R2144_U78);
  not ginst1254 (R2144_U123, R2144_U83);
  nand ginst1255 (R2144_U124, R2144_U105, R2144_U83);
  nand ginst1256 (R2144_U125, R2144_U124, R2144_U21);
  nand ginst1257 (R2144_U126, R2144_U23, R2144_U81);
  nand ginst1258 (R2144_U127, R2144_U124, R2144_U60);
  nand ginst1259 (R2144_U128, R2144_U125, R2144_U61);
  nand ginst1260 (R2144_U129, R2144_U112, U2355);
  not ginst1261 (R2144_U13, U2750);
  not ginst1262 (R2144_U130, R2144_U93);
  nand ginst1263 (R2144_U131, R2144_U14, R2144_U187);
  nand ginst1264 (R2144_U132, R2144_U131, R2144_U93);
  not ginst1265 (R2144_U133, R2144_U91);
  nand ginst1266 (R2144_U134, R2144_U109, R2144_U91);
  nand ginst1267 (R2144_U135, R2144_U116, R2144_U134);
  nand ginst1268 (R2144_U136, R2144_U135, R2144_U62);
  nand ginst1269 (R2144_U137, R2144_U110, R2144_U161);
  nand ginst1270 (R2144_U138, R2144_U116, R2144_U134, R2144_U137);
  not ginst1271 (R2144_U139, R2144_U97);
  not ginst1272 (R2144_U14, U2751);
  not ginst1273 (R2144_U140, R2144_U96);
  not ginst1274 (R2144_U141, R2144_U25);
  not ginst1275 (R2144_U142, R2144_U95);
  not ginst1276 (R2144_U143, R2144_U26);
  nand ginst1277 (R2144_U144, R2144_U24, U2355);
  not ginst1278 (R2144_U145, R2144_U144);
  nand ginst1279 (R2144_U146, R2144_U101, R2144_U12);
  not ginst1280 (R2144_U147, R2144_U94);
  not ginst1281 (R2144_U148, R2144_U98);
  nand ginst1282 (R2144_U149, R2144_U105, R2144_U21);
  not ginst1283 (R2144_U15, U2752);
  nand ginst1284 (R2144_U150, R2144_U106, R2144_U19);
  nand ginst1285 (R2144_U151, R2144_U105, R2144_U120, R2144_U7);
  nand ginst1286 (R2144_U152, R2144_U107, R2144_U7);
  nand ginst1287 (R2144_U153, R2144_U108, R2144_U7);
  nand ginst1288 (R2144_U154, R2144_U100, R2144_U113, R2144_U115);
  nand ginst1289 (R2144_U155, R2144_U114, R2144_U154);
  nand ginst1290 (R2144_U156, R2144_U103, R2144_U104);
  nand ginst1291 (R2144_U157, R2144_U184, U2750);
  nand ginst1292 (R2144_U158, R2144_U110, R2144_U117, R2144_U55);
  nand ginst1293 (R2144_U159, R2144_U106, R2144_U199, U2749);
  not ginst1294 (R2144_U16, U2749);
  nand ginst1295 (R2144_U160, R2144_U158, R2144_U58);
  nand ginst1296 (R2144_U161, R2144_U199, U2749);
  nand ginst1297 (R2144_U162, R2144_U184, U2750);
  nand ginst1298 (R2144_U163, R2144_U109, R2144_U116);
  nand ginst1299 (R2144_U164, R2144_U68, U2355);
  nand ginst1300 (R2144_U165, R2144_U12, U2762);
  nand ginst1301 (R2144_U166, R2144_U69, U2355);
  nand ginst1302 (R2144_U167, R2144_U12, U2761);
  nand ginst1303 (R2144_U168, R2144_U70, U2355);
  nand ginst1304 (R2144_U169, R2144_U12, U2763);
  not ginst1305 (R2144_U17, U2745);
  nand ginst1306 (R2144_U170, R2144_U168, R2144_U169);
  nand ginst1307 (R2144_U171, R2144_U68, U2355);
  nand ginst1308 (R2144_U172, R2144_U12, U2762);
  nand ginst1309 (R2144_U173, R2144_U171, R2144_U172);
  nand ginst1310 (R2144_U174, R2144_U70, U2355);
  nand ginst1311 (R2144_U175, R2144_U12, U2763);
  nand ginst1312 (R2144_U176, R2144_U71, U2355);
  nand ginst1313 (R2144_U177, R2144_U12, U2764);
  nand ginst1314 (R2144_U178, R2144_U176, R2144_U177);
  nand ginst1315 (R2144_U179, R2144_U69, U2355);
  not ginst1316 (R2144_U18, U2748);
  nand ginst1317 (R2144_U180, R2144_U12, U2761);
  nand ginst1318 (R2144_U181, R2144_U179, R2144_U180);
  nand ginst1319 (R2144_U182, R2144_U72, U2355);
  nand ginst1320 (R2144_U183, R2144_U12, U2766);
  nand ginst1321 (R2144_U184, R2144_U182, R2144_U183);
  nand ginst1322 (R2144_U185, R2144_U73, U2355);
  nand ginst1323 (R2144_U186, R2144_U12, U2767);
  not ginst1324 (R2144_U187, R2144_U28);
  nand ginst1325 (R2144_U188, R2144_U74, U2355);
  nand ginst1326 (R2144_U189, R2144_U12, U2768);
  nand ginst1327 (R2144_U19, R2144_U178, U2748);
  nand ginst1328 (R2144_U190, R2144_U74, U2355);
  nand ginst1329 (R2144_U191, R2144_U12, U2768);
  nand ginst1330 (R2144_U192, R2144_U190, R2144_U191);
  nand ginst1331 (R2144_U193, R2144_U72, U2355);
  nand ginst1332 (R2144_U194, R2144_U12, U2766);
  nand ginst1333 (R2144_U195, R2144_U75, U2355);
  nand ginst1334 (R2144_U196, R2144_U12, U2765);
  nand ginst1335 (R2144_U197, R2144_U75, U2355);
  nand ginst1336 (R2144_U198, R2144_U12, U2765);
  nand ginst1337 (R2144_U199, R2144_U197, R2144_U198);
  not ginst1338 (R2144_U20, U2747);
  nand ginst1339 (R2144_U200, R2144_U71, U2355);
  nand ginst1340 (R2144_U201, R2144_U12, U2764);
  nand ginst1341 (R2144_U202, R2144_U76, U2355);
  nand ginst1342 (R2144_U203, R2144_U12, U2760);
  not ginst1343 (R2144_U204, R2144_U29);
  nand ginst1344 (R2144_U205, R2144_U77, U2355);
  nand ginst1345 (R2144_U206, R2144_U12, U2759);
  not ginst1346 (R2144_U207, R2144_U27);
  nand ginst1347 (R2144_U208, R2144_U122, R2144_U207);
  nand ginst1348 (R2144_U209, R2144_U27, R2144_U78);
  nand ginst1349 (R2144_U21, R2144_U170, U2747);
  nand ginst1350 (R2144_U210, R2144_U121, R2144_U204);
  nand ginst1351 (R2144_U211, R2144_U29, R2144_U79);
  nand ginst1352 (R2144_U212, R2144_U124, R2144_U23, R2144_U57);
  nand ginst1353 (R2144_U213, R2144_U108, R2144_U5);
  nand ginst1354 (R2144_U214, R2144_U102, R2144_U156);
  nand ginst1355 (R2144_U215, R2144_U160, R2144_U59, R2144_U81);
  nand ginst1356 (R2144_U216, R2144_U149, R2144_U83);
  nand ginst1357 (R2144_U217, R2144_U123, R2144_U44);
  nand ginst1358 (R2144_U218, R2144_U150, R2144_U84);
  nand ginst1359 (R2144_U219, R2144_U119, R2144_U46);
  not ginst1360 (R2144_U22, U2746);
  nand ginst1361 (R2144_U220, R2144_U85, U2355);
  nand ginst1362 (R2144_U221, R2144_U12, U2754);
  not ginst1363 (R2144_U222, R2144_U32);
  nand ginst1364 (R2144_U223, R2144_U86, U2355);
  nand ginst1365 (R2144_U224, R2144_U12, U2753);
  not ginst1366 (R2144_U225, R2144_U31);
  nand ginst1367 (R2144_U226, R2144_U87, U2355);
  nand ginst1368 (R2144_U227, R2144_U12, U2755);
  not ginst1369 (R2144_U228, R2144_U33);
  nand ginst1370 (R2144_U229, R2144_U88, U2355);
  nand ginst1371 (R2144_U23, R2144_U173, U2746);
  nand ginst1372 (R2144_U230, R2144_U12, U2756);
  not ginst1373 (R2144_U231, R2144_U34);
  nand ginst1374 (R2144_U232, R2144_U89, U2355);
  nand ginst1375 (R2144_U233, R2144_U12, U2757);
  not ginst1376 (R2144_U234, R2144_U35);
  nand ginst1377 (R2144_U235, R2144_U90, U2355);
  nand ginst1378 (R2144_U236, R2144_U12, U2758);
  not ginst1379 (R2144_U237, R2144_U36);
  nand ginst1380 (R2144_U238, R2144_U163, R2144_U91);
  nand ginst1381 (R2144_U239, R2144_U133, R2144_U48);
  nand ginst1382 (R2144_U24, R2144_U63, R2144_U79);
  nand ginst1383 (R2144_U240, R2144_U187, U2751);
  nand ginst1384 (R2144_U241, R2144_U14, R2144_U28);
  nand ginst1385 (R2144_U242, R2144_U187, U2751);
  nand ginst1386 (R2144_U243, R2144_U14, R2144_U28);
  nand ginst1387 (R2144_U244, R2144_U242, R2144_U243);
  nand ginst1388 (R2144_U245, R2144_U92, R2144_U93);
  nand ginst1389 (R2144_U246, R2144_U130, R2144_U244);
  nand ginst1390 (R2144_U247, R2144_U147, R2144_U225);
  nand ginst1391 (R2144_U248, R2144_U31, R2144_U94);
  nand ginst1392 (R2144_U249, R2144_U143, R2144_U222);
  nand ginst1393 (R2144_U25, R2144_U6, R2144_U79);
  nand ginst1394 (R2144_U250, R2144_U26, R2144_U32);
  nand ginst1395 (R2144_U251, R2144_U142, R2144_U228);
  nand ginst1396 (R2144_U252, R2144_U33, R2144_U95);
  nand ginst1397 (R2144_U253, R2144_U141, R2144_U231);
  nand ginst1398 (R2144_U254, R2144_U25, R2144_U34);
  nand ginst1399 (R2144_U255, R2144_U140, R2144_U234);
  nand ginst1400 (R2144_U256, R2144_U35, R2144_U96);
  nand ginst1401 (R2144_U257, R2144_U139, R2144_U237);
  nand ginst1402 (R2144_U258, R2144_U36, R2144_U97);
  nand ginst1403 (R2144_U259, R2144_U98, U2355);
  nand ginst1404 (R2144_U26, R2144_U141, R2144_U65);
  nand ginst1405 (R2144_U260, R2144_U12, R2144_U148);
  nand ginst1406 (R2144_U27, R2144_U205, R2144_U206);
  nand ginst1407 (R2144_U28, R2144_U185, R2144_U186);
  nand ginst1408 (R2144_U29, R2144_U202, R2144_U203);
  nand ginst1409 (R2144_U30, R2144_U208, R2144_U209);
  nand ginst1410 (R2144_U31, R2144_U223, R2144_U224);
  nand ginst1411 (R2144_U32, R2144_U220, R2144_U221);
  nand ginst1412 (R2144_U33, R2144_U226, R2144_U227);
  nand ginst1413 (R2144_U34, R2144_U229, R2144_U230);
  nand ginst1414 (R2144_U35, R2144_U232, R2144_U233);
  nand ginst1415 (R2144_U36, R2144_U235, R2144_U236);
  nand ginst1416 (R2144_U37, R2144_U247, R2144_U248);
  nand ginst1417 (R2144_U38, R2144_U249, R2144_U250);
  nand ginst1418 (R2144_U39, R2144_U251, R2144_U252);
  nand ginst1419 (R2144_U40, R2144_U253, R2144_U254);
  nand ginst1420 (R2144_U41, R2144_U255, R2144_U256);
  nand ginst1421 (R2144_U42, R2144_U257, R2144_U258);
  nand ginst1422 (R2144_U43, R2144_U259, R2144_U260);
  and ginst1423 (R2144_U44, R2144_U105, R2144_U21);
  nand ginst1424 (R2144_U45, R2144_U216, R2144_U217);
  and ginst1425 (R2144_U46, R2144_U106, R2144_U19);
  nand ginst1426 (R2144_U47, R2144_U218, R2144_U219);
  and ginst1427 (R2144_U48, R2144_U109, R2144_U162);
  nand ginst1428 (R2144_U49, R2144_U238, R2144_U239);
  and ginst1429 (R2144_U5, R2144_U103, R2144_U104);
  nand ginst1430 (R2144_U50, R2144_U245, R2144_U246);
  and ginst1431 (R2144_U51, R2144_U109, R2144_U110);
  and ginst1432 (R2144_U52, R2144_U105, R2144_U106);
  and ginst1433 (R2144_U53, R2144_U52, R2144_U7);
  and ginst1434 (R2144_U54, R2144_U103, R2144_U151, R2144_U152, R2144_U153);
  and ginst1435 (R2144_U55, R2144_U106, R2144_U109);
  and ginst1436 (R2144_U56, R2144_U159, R2144_U19);
  and ginst1437 (R2144_U57, R2144_U156, R2144_U21);
  and ginst1438 (R2144_U58, R2144_U159, R2144_U19, R2144_U21);
  and ginst1439 (R2144_U59, R2144_U105, R2144_U5);
  and ginst1440 (R2144_U6, R2144_U27, R2144_U29, R2144_U35, R2144_U36);
  and ginst1441 (R2144_U60, R2144_U126, R2144_U21);
  and ginst1442 (R2144_U61, R2144_U23, R2144_U81);
  and ginst1443 (R2144_U62, R2144_U110, R2144_U111);
  and ginst1444 (R2144_U63, R2144_U6, R2144_U64);
  and ginst1445 (R2144_U64, R2144_U31, R2144_U32, R2144_U33, R2144_U34);
  and ginst1446 (R2144_U65, R2144_U33, R2144_U34);
  and ginst1447 (R2144_U66, R2144_U27, R2144_U29, R2144_U36);
  and ginst1448 (R2144_U67, R2144_U27, R2144_U29);
  not ginst1449 (R2144_U68, U2762);
  not ginst1450 (R2144_U69, U2761);
  and ginst1451 (R2144_U7, R2144_U104, R2144_U81);
  not ginst1452 (R2144_U70, U2763);
  not ginst1453 (R2144_U71, U2764);
  not ginst1454 (R2144_U72, U2766);
  not ginst1455 (R2144_U73, U2767);
  not ginst1456 (R2144_U74, U2768);
  not ginst1457 (R2144_U75, U2765);
  not ginst1458 (R2144_U76, U2760);
  not ginst1459 (R2144_U77, U2759);
  nand ginst1460 (R2144_U78, R2144_U29, R2144_U79);
  nand ginst1461 (R2144_U79, R2144_U54, R2144_U99);
  and ginst1462 (R2144_U8, R2144_U136, R2144_U138);
  and ginst1463 (R2144_U80, R2144_U210, R2144_U211);
  nand ginst1464 (R2144_U81, R2144_U164, R2144_U165, R2144_U22);
  and ginst1465 (R2144_U82, R2144_U214, R2144_U215);
  nand ginst1466 (R2144_U83, R2144_U158, R2144_U56);
  nand ginst1467 (R2144_U84, R2144_U111, R2144_U118);
  not ginst1468 (R2144_U85, U2754);
  not ginst1469 (R2144_U86, U2753);
  not ginst1470 (R2144_U87, U2755);
  not ginst1471 (R2144_U88, U2756);
  not ginst1472 (R2144_U89, U2757);
  and ginst1473 (R2144_U9, R2144_U127, R2144_U128);
  not ginst1474 (R2144_U90, U2758);
  nand ginst1475 (R2144_U91, R2144_U100, R2144_U132);
  and ginst1476 (R2144_U92, R2144_U240, R2144_U241);
  nand ginst1477 (R2144_U93, R2144_U113, R2144_U129);
  nand ginst1478 (R2144_U94, R2144_U143, R2144_U32);
  nand ginst1479 (R2144_U95, R2144_U141, R2144_U34);
  nand ginst1480 (R2144_U96, R2144_U66, R2144_U79);
  nand ginst1481 (R2144_U97, R2144_U67, R2144_U79);
  nand ginst1482 (R2144_U98, R2144_U112, R2144_U113);
  nand ginst1483 (R2144_U99, R2144_U53, R2144_U84);
  not ginst1484 (R2167_U10, U2713);
  not ginst1485 (R2167_U11, U2712);
  not ginst1486 (R2167_U12, U2718);
  not ginst1487 (R2167_U13, U2717);
  not ginst1488 (R2167_U14, U2711);
  not ginst1489 (R2167_U15, U2356);
  not ginst1490 (R2167_U16, STATE2_REG_0__SCAN_IN);
  nand ginst1491 (R2167_U17, R2167_U49, R2167_U50);
  and ginst1492 (R2167_U18, R2167_U29, R2167_U30);
  and ginst1493 (R2167_U19, R2167_U32, R2167_U33);
  and ginst1494 (R2167_U20, R2167_U35, R2167_U36);
  and ginst1495 (R2167_U21, R2167_U38, R2167_U39);
  not ginst1496 (R2167_U22, U2721);
  not ginst1497 (R2167_U23, U2722);
  nand ginst1498 (R2167_U24, R2167_U23, U2715);
  nand ginst1499 (R2167_U25, R2167_U22, U2715);
  or ginst1500 (R2167_U26, U2721, U2722);
  nand ginst1501 (R2167_U27, R2167_U8, U2714);
  nand ginst1502 (R2167_U28, R2167_U24, R2167_U25, R2167_U26, R2167_U27);
  nand ginst1503 (R2167_U29, R2167_U7, U2720);
  nand ginst1504 (R2167_U30, R2167_U10, U2719);
  nand ginst1505 (R2167_U31, R2167_U18, R2167_U28);
  nand ginst1506 (R2167_U32, R2167_U9, U2713);
  nand ginst1507 (R2167_U33, R2167_U12, U2712);
  nand ginst1508 (R2167_U34, R2167_U19, R2167_U31);
  nand ginst1509 (R2167_U35, R2167_U11, U2718);
  nand ginst1510 (R2167_U36, R2167_U14, U2717);
  nand ginst1511 (R2167_U37, R2167_U20, R2167_U34);
  nand ginst1512 (R2167_U38, R2167_U13, U2711);
  nand ginst1513 (R2167_U39, R2167_U6, U2356);
  nand ginst1514 (R2167_U40, R2167_U21, R2167_U37);
  nand ginst1515 (R2167_U41, R2167_U15, U2716);
  nand ginst1516 (R2167_U42, R2167_U40, R2167_U41);
  nand ginst1517 (R2167_U43, R2167_U16, U2716);
  nand ginst1518 (R2167_U44, R2167_U42, R2167_U6);
  nand ginst1519 (R2167_U45, R2167_U43, R2167_U44);
  nand ginst1520 (R2167_U46, STATE2_REG_0__SCAN_IN, R2167_U6);
  nand ginst1521 (R2167_U47, R2167_U42, U2716);
  nand ginst1522 (R2167_U48, R2167_U46, R2167_U47);
  nand ginst1523 (R2167_U49, R2167_U15, R2167_U45);
  nand ginst1524 (R2167_U50, R2167_U48, U2356);
  not ginst1525 (R2167_U6, U2716);
  not ginst1526 (R2167_U7, U2714);
  not ginst1527 (R2167_U8, U2720);
  not ginst1528 (R2167_U9, U2719);
  not ginst1529 (R2182_U10, U2742);
  not ginst1530 (R2182_U11, U2741);
  not ginst1531 (R2182_U12, U2740);
  nand ginst1532 (R2182_U13, R2182_U35, R2182_U41);
  not ginst1533 (R2182_U14, U2737);
  not ginst1534 (R2182_U15, U2738);
  nand ginst1535 (R2182_U16, U2723, U2739);
  not ginst1536 (R2182_U17, U2736);
  not ginst1537 (R2182_U18, U2735);
  nand ginst1538 (R2182_U19, R2182_U36, R2182_U49);
  not ginst1539 (R2182_U20, U2734);
  nand ginst1540 (R2182_U21, R2182_U37, R2182_U46);
  nand ginst1541 (R2182_U22, R2182_U48, U2734);
  not ginst1542 (R2182_U23, U2733);
  nand ginst1543 (R2182_U24, R2182_U63, R2182_U64);
  nand ginst1544 (R2182_U25, R2182_U65, R2182_U66);
  nand ginst1545 (R2182_U26, R2182_U67, R2182_U68);
  nand ginst1546 (R2182_U27, R2182_U71, R2182_U72);
  nand ginst1547 (R2182_U28, R2182_U73, R2182_U74);
  nand ginst1548 (R2182_U29, R2182_U75, R2182_U76);
  nand ginst1549 (R2182_U30, R2182_U77, R2182_U78);
  nand ginst1550 (R2182_U31, R2182_U79, R2182_U80);
  nand ginst1551 (R2182_U32, R2182_U81, R2182_U82);
  nand ginst1552 (R2182_U33, R2182_U83, R2182_U84);
  nand ginst1553 (R2182_U34, R2182_U85, R2182_U86);
  and ginst1554 (R2182_U35, U2741, U2742);
  and ginst1555 (R2182_U36, U2737, U2738);
  and ginst1556 (R2182_U37, U2735, U2736);
  nand ginst1557 (R2182_U38, R2182_U41, U2742);
  not ginst1558 (R2182_U39, U2732);
  nand ginst1559 (R2182_U40, R2182_U56, U2733);
  nand ginst1560 (R2182_U41, R2182_U52, R2182_U53);
  and ginst1561 (R2182_U42, R2182_U69, R2182_U70);
  nand ginst1562 (R2182_U43, R2182_U46, U2736);
  nand ginst1563 (R2182_U44, R2182_U49, U2738);
  nand ginst1564 (R2182_U45, R2182_U51, R2182_U62);
  not ginst1565 (R2182_U46, R2182_U19);
  not ginst1566 (R2182_U47, R2182_U13);
  not ginst1567 (R2182_U48, R2182_U21);
  not ginst1568 (R2182_U49, R2182_U16);
  and ginst1569 (R2182_U5, R2182_U47, U2740);
  not ginst1570 (R2182_U50, R2182_U9);
  or ginst1571 (R2182_U51, U2731, U2743);
  nand ginst1572 (R2182_U52, U2731, U2743);
  nand ginst1573 (R2182_U53, R2182_U50, R2182_U51);
  not ginst1574 (R2182_U54, R2182_U41);
  not ginst1575 (R2182_U55, R2182_U38);
  not ginst1576 (R2182_U56, R2182_U22);
  not ginst1577 (R2182_U57, R2182_U40);
  not ginst1578 (R2182_U58, R2182_U43);
  not ginst1579 (R2182_U59, R2182_U44);
  and ginst1580 (R2182_U6, R2182_U16, R2182_U60);
  or ginst1581 (R2182_U60, U2723, U2739);
  not ginst1582 (R2182_U61, R2182_U45);
  nand ginst1583 (R2182_U62, U2731, U2743);
  nand ginst1584 (R2182_U63, R2182_U12, R2182_U47);
  nand ginst1585 (R2182_U64, R2182_U13, U2740);
  nand ginst1586 (R2182_U65, R2182_U38, U2741);
  nand ginst1587 (R2182_U66, R2182_U11, R2182_U55);
  nand ginst1588 (R2182_U67, R2182_U40, U2732);
  nand ginst1589 (R2182_U68, R2182_U39, R2182_U57);
  nand ginst1590 (R2182_U69, R2182_U41, U2742);
  not ginst1591 (R2182_U7, U2744);
  nand ginst1592 (R2182_U70, R2182_U10, R2182_U54);
  nand ginst1593 (R2182_U71, R2182_U22, U2733);
  nand ginst1594 (R2182_U72, R2182_U23, R2182_U56);
  nand ginst1595 (R2182_U73, R2182_U20, R2182_U48);
  nand ginst1596 (R2182_U74, R2182_U21, U2734);
  nand ginst1597 (R2182_U75, R2182_U43, U2735);
  nand ginst1598 (R2182_U76, R2182_U18, R2182_U58);
  nand ginst1599 (R2182_U77, R2182_U17, R2182_U46);
  nand ginst1600 (R2182_U78, R2182_U19, U2736);
  nand ginst1601 (R2182_U79, R2182_U44, U2737);
  not ginst1602 (R2182_U8, U3233);
  nand ginst1603 (R2182_U80, R2182_U14, R2182_U59);
  nand ginst1604 (R2182_U81, R2182_U15, R2182_U49);
  nand ginst1605 (R2182_U82, R2182_U16, U2738);
  nand ginst1606 (R2182_U83, R2182_U45, R2182_U50);
  nand ginst1607 (R2182_U84, R2182_U61, R2182_U9);
  nand ginst1608 (R2182_U85, R2182_U7, U3233);
  nand ginst1609 (R2182_U86, R2182_U8, U2744);
  nand ginst1610 (R2182_U9, U2744, U3233);
  not ginst1611 (R2238_U10, INSTQUEUEWR_ADDR_REG_1__SCAN_IN);
  not ginst1612 (R2238_U11, INSTQUEUERD_ADDR_REG_2__SCAN_IN);
  not ginst1613 (R2238_U12, INSTQUEUEWR_ADDR_REG_2__SCAN_IN);
  not ginst1614 (R2238_U13, INSTQUEUERD_ADDR_REG_3__SCAN_IN);
  not ginst1615 (R2238_U14, INSTQUEUEWR_ADDR_REG_3__SCAN_IN);
  not ginst1616 (R2238_U15, INSTQUEUEWR_ADDR_REG_4__SCAN_IN);
  nand ginst1617 (R2238_U16, R2238_U40, R2238_U41);
  not ginst1618 (R2238_U17, INSTQUEUERD_ADDR_REG_4__SCAN_IN);
  not ginst1619 (R2238_U18, INSTQUEUEWR_ADDR_REG_0__SCAN_IN);
  nand ginst1620 (R2238_U19, R2238_U50, R2238_U51);
  nand ginst1621 (R2238_U20, R2238_U55, R2238_U56);
  nand ginst1622 (R2238_U21, R2238_U60, R2238_U61);
  nand ginst1623 (R2238_U22, R2238_U65, R2238_U66);
  nand ginst1624 (R2238_U23, R2238_U47, R2238_U48);
  nand ginst1625 (R2238_U24, R2238_U52, R2238_U53);
  nand ginst1626 (R2238_U25, R2238_U57, R2238_U58);
  nand ginst1627 (R2238_U26, R2238_U62, R2238_U63);
  nand ginst1628 (R2238_U27, R2238_U36, R2238_U37);
  nand ginst1629 (R2238_U28, R2238_U32, R2238_U33);
  not ginst1630 (R2238_U29, INSTQUEUERD_ADDR_REG_1__SCAN_IN);
  not ginst1631 (R2238_U30, R2238_U9);
  nand ginst1632 (R2238_U31, R2238_U10, R2238_U30);
  nand ginst1633 (R2238_U32, R2238_U29, R2238_U31);
  nand ginst1634 (R2238_U33, INSTQUEUEWR_ADDR_REG_1__SCAN_IN, R2238_U9);
  not ginst1635 (R2238_U34, R2238_U28);
  nand ginst1636 (R2238_U35, INSTQUEUERD_ADDR_REG_2__SCAN_IN, R2238_U12);
  nand ginst1637 (R2238_U36, R2238_U28, R2238_U35);
  nand ginst1638 (R2238_U37, INSTQUEUEWR_ADDR_REG_2__SCAN_IN, R2238_U11);
  not ginst1639 (R2238_U38, R2238_U27);
  nand ginst1640 (R2238_U39, INSTQUEUERD_ADDR_REG_3__SCAN_IN, R2238_U14);
  nand ginst1641 (R2238_U40, R2238_U27, R2238_U39);
  nand ginst1642 (R2238_U41, INSTQUEUEWR_ADDR_REG_3__SCAN_IN, R2238_U13);
  not ginst1643 (R2238_U42, R2238_U16);
  nand ginst1644 (R2238_U43, INSTQUEUEWR_ADDR_REG_4__SCAN_IN, R2238_U17);
  nand ginst1645 (R2238_U44, R2238_U42, R2238_U43);
  nand ginst1646 (R2238_U45, INSTQUEUERD_ADDR_REG_4__SCAN_IN, R2238_U15);
  nand ginst1647 (R2238_U46, INSTQUEUEWR_ADDR_REG_0__SCAN_IN, R2238_U8);
  nand ginst1648 (R2238_U47, INSTQUEUERD_ADDR_REG_4__SCAN_IN, R2238_U15);
  nand ginst1649 (R2238_U48, INSTQUEUEWR_ADDR_REG_4__SCAN_IN, R2238_U17);
  not ginst1650 (R2238_U49, R2238_U23);
  nand ginst1651 (R2238_U50, R2238_U42, R2238_U49);
  nand ginst1652 (R2238_U51, R2238_U16, R2238_U23);
  nand ginst1653 (R2238_U52, INSTQUEUERD_ADDR_REG_3__SCAN_IN, R2238_U14);
  nand ginst1654 (R2238_U53, INSTQUEUEWR_ADDR_REG_3__SCAN_IN, R2238_U13);
  not ginst1655 (R2238_U54, R2238_U24);
  nand ginst1656 (R2238_U55, R2238_U38, R2238_U54);
  nand ginst1657 (R2238_U56, R2238_U24, R2238_U27);
  nand ginst1658 (R2238_U57, INSTQUEUERD_ADDR_REG_2__SCAN_IN, R2238_U12);
  nand ginst1659 (R2238_U58, INSTQUEUEWR_ADDR_REG_2__SCAN_IN, R2238_U11);
  not ginst1660 (R2238_U59, R2238_U25);
  nand ginst1661 (R2238_U6, R2238_U44, R2238_U45);
  nand ginst1662 (R2238_U60, R2238_U34, R2238_U59);
  nand ginst1663 (R2238_U61, R2238_U25, R2238_U28);
  nand ginst1664 (R2238_U62, INSTQUEUERD_ADDR_REG_1__SCAN_IN, R2238_U10);
  nand ginst1665 (R2238_U63, INSTQUEUEWR_ADDR_REG_1__SCAN_IN, R2238_U29);
  not ginst1666 (R2238_U64, R2238_U26);
  nand ginst1667 (R2238_U65, R2238_U30, R2238_U64);
  nand ginst1668 (R2238_U66, R2238_U26, R2238_U9);
  nand ginst1669 (R2238_U7, R2238_U46, R2238_U9);
  not ginst1670 (R2238_U8, INSTQUEUERD_ADDR_REG_0__SCAN_IN);
  nand ginst1671 (R2238_U9, INSTQUEUERD_ADDR_REG_0__SCAN_IN, R2238_U18);
  and ginst1672 (R2278_U10, R2278_U206, R2278_U9);
  nand ginst1673 (R2278_U100, R2278_U167, R2278_U172);
  and ginst1674 (R2278_U101, R2278_U373, R2278_U374);
  nand ginst1675 (R2278_U102, R2278_U324, R2278_U326);
  and ginst1676 (R2278_U103, R2278_U378, R2278_U379);
  nand ginst1677 (R2278_U104, R2278_U321, R2278_U323);
  and ginst1678 (R2278_U105, R2278_U383, R2278_U384);
  nand ginst1679 (R2278_U106, R2278_U248, R2278_U36);
  nand ginst1680 (R2278_U107, R2278_U250, R2278_U251);
  and ginst1681 (R2278_U108, R2278_U385, R2278_U386);
  nand ginst1682 (R2278_U109, R2278_U246, R2278_U36);
  and ginst1683 (R2278_U11, R2278_U10, R2278_U205);
  nand ginst1684 (R2278_U110, R2278_U347, R2278_U59);
  and ginst1685 (R2278_U111, R2278_U387, R2278_U388);
  nand ginst1686 (R2278_U112, R2278_U316, R2278_U67);
  nand ginst1687 (R2278_U113, R2278_U204, R2278_U245);
  and ginst1688 (R2278_U114, R2278_U389, R2278_U390);
  nand ginst1689 (R2278_U115, R2278_U313, R2278_U68);
  nand ginst1690 (R2278_U116, R2278_U242, R2278_U243);
  and ginst1691 (R2278_U117, R2278_U391, R2278_U392);
  nand ginst1692 (R2278_U118, R2278_U311, R2278_U69);
  nand ginst1693 (R2278_U119, R2278_U205, R2278_U240);
  and ginst1694 (R2278_U12, R2278_U11, R2278_U242);
  and ginst1695 (R2278_U120, R2278_U393, R2278_U394);
  nand ginst1696 (R2278_U121, R2278_U309, R2278_U70);
  nand ginst1697 (R2278_U122, R2278_U206, R2278_U238);
  and ginst1698 (R2278_U123, R2278_U395, R2278_U396);
  nand ginst1699 (R2278_U124, R2278_U232, R2278_U233);
  nand ginst1700 (R2278_U125, R2278_U235, R2278_U236);
  and ginst1701 (R2278_U126, R2278_U397, R2278_U398);
  nand ginst1702 (R2278_U127, R2278_U231, R2278_U232);
  nand ginst1703 (R2278_U128, R2278_U345, R2278_U66);
  and ginst1704 (R2278_U129, R2278_U399, R2278_U400);
  and ginst1705 (R2278_U13, R2278_U12, R2278_U204);
  nand ginst1706 (R2278_U130, R2278_U168, R2278_U169);
  nand ginst1707 (R2278_U131, R2278_U207, R2278_U23);
  nand ginst1708 (R2278_U132, R2278_U307, R2278_U343);
  and ginst1709 (R2278_U133, R2278_U403, R2278_U404);
  nand ginst1710 (R2278_U134, R2278_U208, R2278_U229);
  nand ginst1711 (R2278_U135, R2278_U305, R2278_U341);
  and ginst1712 (R2278_U136, R2278_U405, R2278_U406);
  nand ginst1713 (R2278_U137, R2278_U227, R2278_U228);
  nand ginst1714 (R2278_U138, R2278_U24, R2278_U339);
  and ginst1715 (R2278_U139, R2278_U407, R2278_U408);
  and ginst1716 (R2278_U14, R2278_U246, R2278_U250);
  nand ginst1717 (R2278_U140, R2278_U223, R2278_U56);
  nand ginst1718 (R2278_U141, R2278_U225, R2278_U24);
  and ginst1719 (R2278_U142, R2278_U409, R2278_U410);
  nand ginst1720 (R2278_U143, R2278_U280, R2278_U30);
  nand ginst1721 (R2278_U144, R2278_U209, R2278_U210);
  and ginst1722 (R2278_U145, R2278_U411, R2278_U412);
  nand ginst1723 (R2278_U146, R2278_U278, R2278_U31);
  nand ginst1724 (R2278_U147, R2278_U211, R2278_U30);
  and ginst1725 (R2278_U148, R2278_U413, R2278_U414);
  nand ginst1726 (R2278_U149, R2278_U276, R2278_U29);
  and ginst1727 (R2278_U15, R2278_U14, R2278_U253);
  nand ginst1728 (R2278_U150, R2278_U213, R2278_U31);
  and ginst1729 (R2278_U151, R2278_U415, R2278_U416);
  nand ginst1730 (R2278_U152, R2278_U219, R2278_U71);
  nand ginst1731 (R2278_U153, R2278_U221, R2278_U29);
  and ginst1732 (R2278_U154, R2278_U417, R2278_U418);
  nand ginst1733 (R2278_U155, R2278_U28, R2278_U288);
  nand ginst1734 (R2278_U156, R2278_U215, R2278_U216);
  and ginst1735 (R2278_U157, R2278_U419, R2278_U420);
  nand ginst1736 (R2278_U158, R2278_U27, R2278_U286);
  nand ginst1737 (R2278_U159, R2278_U217, R2278_U28);
  and ginst1738 (R2278_U16, R2278_U15, R2278_U256);
  and ginst1739 (R2278_U160, R2278_U421, R2278_U422);
  not ginst1740 (R2278_U161, R2278_U19);
  or ginst1741 (R2278_U162, INSTADDRPOINTER_REG_7__SCAN_IN, U2780);
  nand ginst1742 (R2278_U163, INSTADDRPOINTER_REG_7__SCAN_IN, U2780);
  or ginst1743 (R2278_U164, INSTADDRPOINTER_REG_6__SCAN_IN, U2781);
  nand ginst1744 (R2278_U165, INSTADDRPOINTER_REG_6__SCAN_IN, U2781);
  or ginst1745 (R2278_U166, INSTADDRPOINTER_REG_3__SCAN_IN, U2784);
  or ginst1746 (R2278_U167, INSTADDRPOINTER_REG_2__SCAN_IN, U2785);
  or ginst1747 (R2278_U168, INSTADDRPOINTER_REG_1__SCAN_IN, U2786);
  nand ginst1748 (R2278_U169, INSTADDRPOINTER_REG_1__SCAN_IN, U2786);
  and ginst1749 (R2278_U17, R2278_U19, R2278_U292);
  nand ginst1750 (R2278_U170, R2278_U161, R2278_U168);
  not ginst1751 (R2278_U171, R2278_U99);
  nand ginst1752 (R2278_U172, INSTADDRPOINTER_REG_2__SCAN_IN, U2785);
  nand ginst1753 (R2278_U173, R2278_U299, R2278_U99);
  not ginst1754 (R2278_U174, R2278_U90);
  nand ginst1755 (R2278_U175, INSTADDRPOINTER_REG_3__SCAN_IN, U2784);
  nand ginst1756 (R2278_U176, R2278_U166, R2278_U300);
  not ginst1757 (R2278_U177, R2278_U87);
  or ginst1758 (R2278_U178, INSTADDRPOINTER_REG_4__SCAN_IN, U2783);
  or ginst1759 (R2278_U179, INSTADDRPOINTER_REG_5__SCAN_IN, U2782);
  nand ginst1760 (R2278_U18, INSTADDRPOINTER_REG_4__SCAN_IN, U2783);
  not ginst1761 (R2278_U180, R2278_U20);
  not ginst1762 (R2278_U181, R2278_U18);
  nand ginst1763 (R2278_U182, R2278_U162, R2278_U164, R2278_U179, R2278_U181);
  nand ginst1764 (R2278_U183, R2278_U43, R2278_U44, R2278_U87);
  not ginst1765 (R2278_U184, R2278_U75);
  or ginst1766 (R2278_U185, INSTADDRPOINTER_REG_8__SCAN_IN, U2779);
  not ginst1767 (R2278_U186, R2278_U26);
  nand ginst1768 (R2278_U187, R2278_U185, R2278_U75);
  not ginst1769 (R2278_U188, R2278_U72);
  or ginst1770 (R2278_U189, INSTADDRPOINTER_REG_9__SCAN_IN, U2778);
  nand ginst1771 (R2278_U19, INSTADDRPOINTER_REG_0__SCAN_IN, U2787);
  not ginst1772 (R2278_U190, R2278_U27);
  not ginst1773 (R2278_U191, R2278_U73);
  not ginst1774 (R2278_U192, R2278_U76);
  nand ginst1775 (R2278_U193, R2278_U178, R2278_U87);
  not ginst1776 (R2278_U194, R2278_U84);
  nand ginst1777 (R2278_U195, R2278_U179, R2278_U84);
  not ginst1778 (R2278_U196, R2278_U81);
  nand ginst1779 (R2278_U197, R2278_U164, R2278_U81);
  not ginst1780 (R2278_U198, R2278_U78);
  not ginst1781 (R2278_U199, R2278_U79);
  nand ginst1782 (R2278_U20, INSTADDRPOINTER_REG_5__SCAN_IN, U2782);
  not ginst1783 (R2278_U200, R2278_U82);
  not ginst1784 (R2278_U201, R2278_U85);
  not ginst1785 (R2278_U202, R2278_U88);
  not ginst1786 (R2278_U203, R2278_U91);
  or ginst1787 (R2278_U204, INSTADDRPOINTER_REG_25__SCAN_IN, U2770);
  or ginst1788 (R2278_U205, INSTADDRPOINTER_REG_23__SCAN_IN, U2770);
  or ginst1789 (R2278_U206, INSTADDRPOINTER_REG_22__SCAN_IN, U2770);
  or ginst1790 (R2278_U207, INSTADDRPOINTER_REG_19__SCAN_IN, U2770);
  or ginst1791 (R2278_U208, INSTADDRPOINTER_REG_18__SCAN_IN, U2770);
  or ginst1792 (R2278_U209, INSTADDRPOINTER_REG_15__SCAN_IN, U2772);
  not ginst1793 (R2278_U21, INSTADDRPOINTER_REG_30__SCAN_IN);
  nand ginst1794 (R2278_U210, INSTADDRPOINTER_REG_15__SCAN_IN, U2772);
  or ginst1795 (R2278_U211, INSTADDRPOINTER_REG_14__SCAN_IN, U2773);
  not ginst1796 (R2278_U212, R2278_U30);
  or ginst1797 (R2278_U213, INSTADDRPOINTER_REG_13__SCAN_IN, U2774);
  not ginst1798 (R2278_U214, R2278_U31);
  or ginst1799 (R2278_U215, INSTADDRPOINTER_REG_11__SCAN_IN, U2776);
  nand ginst1800 (R2278_U216, INSTADDRPOINTER_REG_11__SCAN_IN, U2776);
  or ginst1801 (R2278_U217, INSTADDRPOINTER_REG_10__SCAN_IN, U2777);
  not ginst1802 (R2278_U218, R2278_U28);
  nand ginst1803 (R2278_U219, R2278_U335, R2278_U52);
  not ginst1804 (R2278_U22, U2770);
  not ginst1805 (R2278_U220, R2278_U152);
  or ginst1806 (R2278_U221, INSTADDRPOINTER_REG_12__SCAN_IN, U2775);
  not ginst1807 (R2278_U222, R2278_U29);
  nand ginst1808 (R2278_U223, R2278_U338, R2278_U55);
  not ginst1809 (R2278_U224, R2278_U140);
  or ginst1810 (R2278_U225, INSTADDRPOINTER_REG_16__SCAN_IN, U2771);
  not ginst1811 (R2278_U226, R2278_U24);
  or ginst1812 (R2278_U227, INSTADDRPOINTER_REG_17__SCAN_IN, U2770);
  nand ginst1813 (R2278_U228, INSTADDRPOINTER_REG_17__SCAN_IN, U2770);
  nand ginst1814 (R2278_U229, INSTADDRPOINTER_REG_18__SCAN_IN, U2770);
  nand ginst1815 (R2278_U23, INSTADDRPOINTER_REG_19__SCAN_IN, U2770);
  not ginst1816 (R2278_U230, R2278_U23);
  or ginst1817 (R2278_U231, INSTADDRPOINTER_REG_20__SCAN_IN, U2770);
  nand ginst1818 (R2278_U232, INSTADDRPOINTER_REG_20__SCAN_IN, U2770);
  nand ginst1819 (R2278_U233, R2278_U128, R2278_U231);
  not ginst1820 (R2278_U234, R2278_U124);
  or ginst1821 (R2278_U235, INSTADDRPOINTER_REG_21__SCAN_IN, U2770);
  nand ginst1822 (R2278_U236, INSTADDRPOINTER_REG_21__SCAN_IN, U2770);
  not ginst1823 (R2278_U237, R2278_U121);
  nand ginst1824 (R2278_U238, INSTADDRPOINTER_REG_22__SCAN_IN, U2770);
  not ginst1825 (R2278_U239, R2278_U118);
  nand ginst1826 (R2278_U24, INSTADDRPOINTER_REG_16__SCAN_IN, U2771);
  nand ginst1827 (R2278_U240, INSTADDRPOINTER_REG_23__SCAN_IN, U2770);
  not ginst1828 (R2278_U241, R2278_U115);
  or ginst1829 (R2278_U242, INSTADDRPOINTER_REG_24__SCAN_IN, U2770);
  nand ginst1830 (R2278_U243, INSTADDRPOINTER_REG_24__SCAN_IN, U2770);
  not ginst1831 (R2278_U244, R2278_U112);
  nand ginst1832 (R2278_U245, INSTADDRPOINTER_REG_25__SCAN_IN, U2770);
  or ginst1833 (R2278_U246, INSTADDRPOINTER_REG_26__SCAN_IN, U2770);
  not ginst1834 (R2278_U247, R2278_U36);
  nand ginst1835 (R2278_U248, R2278_U110, R2278_U246);
  not ginst1836 (R2278_U249, R2278_U106);
  nand ginst1837 (R2278_U25, R2278_U207, R2278_U40);
  or ginst1838 (R2278_U250, INSTADDRPOINTER_REG_27__SCAN_IN, U2770);
  nand ginst1839 (R2278_U251, INSTADDRPOINTER_REG_27__SCAN_IN, U2770);
  not ginst1840 (R2278_U252, R2278_U104);
  or ginst1841 (R2278_U253, INSTADDRPOINTER_REG_28__SCAN_IN, U2770);
  nand ginst1842 (R2278_U254, INSTADDRPOINTER_REG_28__SCAN_IN, U2770);
  not ginst1843 (R2278_U255, R2278_U102);
  or ginst1844 (R2278_U256, INSTADDRPOINTER_REG_29__SCAN_IN, U2770);
  nand ginst1845 (R2278_U257, INSTADDRPOINTER_REG_29__SCAN_IN, U2770);
  not ginst1846 (R2278_U258, R2278_U97);
  or ginst1847 (R2278_U259, INSTADDRPOINTER_REG_30__SCAN_IN, U2770);
  nand ginst1848 (R2278_U26, INSTADDRPOINTER_REG_8__SCAN_IN, U2779);
  nand ginst1849 (R2278_U260, INSTADDRPOINTER_REG_30__SCAN_IN, U2770);
  not ginst1850 (R2278_U261, R2278_U95);
  not ginst1851 (R2278_U262, R2278_U100);
  not ginst1852 (R2278_U263, R2278_U107);
  not ginst1853 (R2278_U264, R2278_U109);
  not ginst1854 (R2278_U265, R2278_U113);
  not ginst1855 (R2278_U266, R2278_U116);
  not ginst1856 (R2278_U267, R2278_U119);
  not ginst1857 (R2278_U268, R2278_U122);
  not ginst1858 (R2278_U269, R2278_U125);
  nand ginst1859 (R2278_U27, INSTADDRPOINTER_REG_9__SCAN_IN, U2778);
  not ginst1860 (R2278_U270, R2278_U127);
  not ginst1861 (R2278_U271, R2278_U130);
  not ginst1862 (R2278_U272, R2278_U131);
  not ginst1863 (R2278_U273, R2278_U134);
  not ginst1864 (R2278_U274, R2278_U137);
  not ginst1865 (R2278_U275, R2278_U141);
  nand ginst1866 (R2278_U276, R2278_U152, R2278_U221);
  not ginst1867 (R2278_U277, R2278_U149);
  nand ginst1868 (R2278_U278, R2278_U149, R2278_U213);
  not ginst1869 (R2278_U279, R2278_U146);
  nand ginst1870 (R2278_U28, INSTADDRPOINTER_REG_10__SCAN_IN, U2777);
  nand ginst1871 (R2278_U280, R2278_U146, R2278_U211);
  not ginst1872 (R2278_U281, R2278_U143);
  not ginst1873 (R2278_U282, R2278_U144);
  not ginst1874 (R2278_U283, R2278_U147);
  not ginst1875 (R2278_U284, R2278_U150);
  not ginst1876 (R2278_U285, R2278_U153);
  nand ginst1877 (R2278_U286, R2278_U189, R2278_U72);
  not ginst1878 (R2278_U287, R2278_U158);
  nand ginst1879 (R2278_U288, R2278_U158, R2278_U217);
  not ginst1880 (R2278_U289, R2278_U155);
  nand ginst1881 (R2278_U29, INSTADDRPOINTER_REG_12__SCAN_IN, U2775);
  not ginst1882 (R2278_U290, R2278_U156);
  not ginst1883 (R2278_U291, R2278_U159);
  or ginst1884 (R2278_U292, INSTADDRPOINTER_REG_0__SCAN_IN, U2787);
  nand ginst1885 (R2278_U293, R2278_U5, R2278_U53);
  nand ginst1886 (R2278_U294, R2278_U209, R2278_U211, R2278_U213, R2278_U222);
  nand ginst1887 (R2278_U295, R2278_U190, R2278_U5);
  nand ginst1888 (R2278_U296, R2278_U218, R2278_U5);
  nand ginst1889 (R2278_U297, R2278_U209, R2278_U212);
  nand ginst1890 (R2278_U298, R2278_U209, R2278_U211, R2278_U214);
  or ginst1891 (R2278_U299, INSTADDRPOINTER_REG_2__SCAN_IN, U2785);
  nand ginst1892 (R2278_U30, INSTADDRPOINTER_REG_14__SCAN_IN, U2773);
  nand ginst1893 (R2278_U300, R2278_U172, R2278_U173);
  nand ginst1894 (R2278_U301, INSTADDRPOINTER_REG_6__SCAN_IN, R2278_U162, U2781);
  nand ginst1895 (R2278_U302, R2278_U162, R2278_U164, R2278_U180);
  or ginst1896 (R2278_U303, INSTADDRPOINTER_REG_6__SCAN_IN, U2781);
  nand ginst1897 (R2278_U304, R2278_U226, R2278_U227);
  not ginst1898 (R2278_U305, R2278_U41);
  nand ginst1899 (R2278_U306, R2278_U208, R2278_U41);
  not ginst1900 (R2278_U307, R2278_U40);
  not ginst1901 (R2278_U308, R2278_U25);
  nand ginst1902 (R2278_U309, R2278_U128, R2278_U9);
  nand ginst1903 (R2278_U31, INSTADDRPOINTER_REG_13__SCAN_IN, U2774);
  nand ginst1904 (R2278_U310, R2278_U235, R2278_U47);
  nand ginst1905 (R2278_U311, R2278_U10, R2278_U128);
  nand ginst1906 (R2278_U312, R2278_U206, R2278_U334);
  nand ginst1907 (R2278_U313, R2278_U11, R2278_U128);
  nand ginst1908 (R2278_U314, R2278_U238, R2278_U312);
  nand ginst1909 (R2278_U315, R2278_U205, R2278_U314);
  nand ginst1910 (R2278_U316, R2278_U12, R2278_U128);
  nand ginst1911 (R2278_U317, R2278_U240, R2278_U315);
  nand ginst1912 (R2278_U318, R2278_U242, R2278_U317);
  nand ginst1913 (R2278_U319, R2278_U243, R2278_U318);
  not ginst1914 (R2278_U32, INSTADDRPOINTER_REG_29__SCAN_IN);
  nand ginst1915 (R2278_U320, R2278_U204, R2278_U319);
  nand ginst1916 (R2278_U321, R2278_U110, R2278_U14);
  nand ginst1917 (R2278_U322, R2278_U247, R2278_U250);
  not ginst1918 (R2278_U323, R2278_U39);
  nand ginst1919 (R2278_U324, R2278_U110, R2278_U15);
  nand ginst1920 (R2278_U325, R2278_U253, R2278_U39);
  not ginst1921 (R2278_U326, R2278_U38);
  nand ginst1922 (R2278_U327, R2278_U110, R2278_U16);
  nand ginst1923 (R2278_U328, R2278_U256, R2278_U38);
  not ginst1924 (R2278_U329, R2278_U37);
  not ginst1925 (R2278_U33, U2770);
  nand ginst1926 (R2278_U330, R2278_U110, R2278_U60);
  nand ginst1927 (R2278_U331, R2278_U259, R2278_U37);
  nand ginst1928 (R2278_U332, R2278_U13, R2278_U230);
  nand ginst1929 (R2278_U333, R2278_U13, R2278_U308);
  nand ginst1930 (R2278_U334, R2278_U236, R2278_U310);
  nand ginst1931 (R2278_U335, R2278_U302, R2278_U336, R2278_U50);
  nand ginst1932 (R2278_U336, R2278_U48, R2278_U49, R2278_U87);
  or ginst1933 (R2278_U337, INSTADDRPOINTER_REG_6__SCAN_IN, U2781);
  nand ginst1934 (R2278_U338, R2278_U219, R2278_U54);
  nand ginst1935 (R2278_U339, R2278_U140, R2278_U225);
  not ginst1936 (R2278_U34, INSTADDRPOINTER_REG_28__SCAN_IN);
  not ginst1937 (R2278_U340, R2278_U138);
  nand ginst1938 (R2278_U341, R2278_U140, R2278_U6);
  not ginst1939 (R2278_U342, R2278_U135);
  nand ginst1940 (R2278_U343, R2278_U140, R2278_U7);
  not ginst1941 (R2278_U344, R2278_U132);
  nand ginst1942 (R2278_U345, R2278_U140, R2278_U8);
  not ginst1943 (R2278_U346, R2278_U128);
  nand ginst1944 (R2278_U347, R2278_U140, R2278_U57);
  not ginst1945 (R2278_U348, R2278_U110);
  nand ginst1946 (R2278_U349, R2278_U188, R2278_U73);
  not ginst1947 (R2278_U35, U2770);
  nand ginst1948 (R2278_U350, R2278_U191, R2278_U72);
  nand ginst1949 (R2278_U351, R2278_U184, R2278_U76);
  nand ginst1950 (R2278_U352, R2278_U192, R2278_U75);
  nand ginst1951 (R2278_U353, R2278_U198, R2278_U79);
  nand ginst1952 (R2278_U354, R2278_U199, R2278_U78);
  nand ginst1953 (R2278_U355, R2278_U196, R2278_U82);
  nand ginst1954 (R2278_U356, R2278_U200, R2278_U81);
  nand ginst1955 (R2278_U357, R2278_U194, R2278_U85);
  nand ginst1956 (R2278_U358, R2278_U201, R2278_U84);
  nand ginst1957 (R2278_U359, R2278_U177, R2278_U88);
  nand ginst1958 (R2278_U36, INSTADDRPOINTER_REG_26__SCAN_IN, U2770);
  nand ginst1959 (R2278_U360, R2278_U202, R2278_U87);
  nand ginst1960 (R2278_U361, R2278_U174, R2278_U91);
  nand ginst1961 (R2278_U362, R2278_U203, R2278_U90);
  nand ginst1962 (R2278_U363, R2278_U94, U2769);
  nand ginst1963 (R2278_U364, INSTADDRPOINTER_REG_31__SCAN_IN, R2278_U93);
  not ginst1964 (R2278_U365, R2278_U62);
  nand ginst1965 (R2278_U366, R2278_U261, R2278_U365);
  nand ginst1966 (R2278_U367, R2278_U62, R2278_U95);
  nand ginst1967 (R2278_U368, R2278_U21, U2770);
  nand ginst1968 (R2278_U369, INSTADDRPOINTER_REG_30__SCAN_IN, R2278_U22);
  nand ginst1969 (R2278_U37, R2278_U257, R2278_U328);
  not ginst1970 (R2278_U370, R2278_U63);
  nand ginst1971 (R2278_U371, R2278_U258, R2278_U370);
  nand ginst1972 (R2278_U372, R2278_U63, R2278_U97);
  nand ginst1973 (R2278_U373, R2278_U100, R2278_U171);
  nand ginst1974 (R2278_U374, R2278_U262, R2278_U99);
  nand ginst1975 (R2278_U375, R2278_U32, U2770);
  nand ginst1976 (R2278_U376, INSTADDRPOINTER_REG_29__SCAN_IN, R2278_U33);
  not ginst1977 (R2278_U377, R2278_U64);
  nand ginst1978 (R2278_U378, R2278_U255, R2278_U377);
  nand ginst1979 (R2278_U379, R2278_U102, R2278_U64);
  nand ginst1980 (R2278_U38, R2278_U254, R2278_U325);
  nand ginst1981 (R2278_U380, R2278_U34, U2770);
  nand ginst1982 (R2278_U381, INSTADDRPOINTER_REG_28__SCAN_IN, R2278_U35);
  not ginst1983 (R2278_U382, R2278_U65);
  nand ginst1984 (R2278_U383, R2278_U252, R2278_U382);
  nand ginst1985 (R2278_U384, R2278_U104, R2278_U65);
  nand ginst1986 (R2278_U385, R2278_U107, R2278_U249);
  nand ginst1987 (R2278_U386, R2278_U106, R2278_U263);
  nand ginst1988 (R2278_U387, R2278_U110, R2278_U264);
  nand ginst1989 (R2278_U388, R2278_U109, R2278_U348);
  nand ginst1990 (R2278_U389, R2278_U113, R2278_U244);
  nand ginst1991 (R2278_U39, R2278_U251, R2278_U322);
  nand ginst1992 (R2278_U390, R2278_U112, R2278_U265);
  nand ginst1993 (R2278_U391, R2278_U116, R2278_U241);
  nand ginst1994 (R2278_U392, R2278_U115, R2278_U266);
  nand ginst1995 (R2278_U393, R2278_U119, R2278_U239);
  nand ginst1996 (R2278_U394, R2278_U118, R2278_U267);
  nand ginst1997 (R2278_U395, R2278_U122, R2278_U237);
  nand ginst1998 (R2278_U396, R2278_U121, R2278_U268);
  nand ginst1999 (R2278_U397, R2278_U125, R2278_U234);
  nand ginst2000 (R2278_U398, R2278_U124, R2278_U269);
  nand ginst2001 (R2278_U399, R2278_U128, R2278_U270);
  nand ginst2002 (R2278_U40, R2278_U229, R2278_U306);
  nand ginst2003 (R2278_U400, R2278_U127, R2278_U346);
  nand ginst2004 (R2278_U401, R2278_U130, R2278_U161);
  nand ginst2005 (R2278_U402, R2278_U19, R2278_U271);
  nand ginst2006 (R2278_U403, R2278_U132, R2278_U272);
  nand ginst2007 (R2278_U404, R2278_U131, R2278_U344);
  nand ginst2008 (R2278_U405, R2278_U135, R2278_U273);
  nand ginst2009 (R2278_U406, R2278_U134, R2278_U342);
  nand ginst2010 (R2278_U407, R2278_U138, R2278_U274);
  nand ginst2011 (R2278_U408, R2278_U137, R2278_U340);
  nand ginst2012 (R2278_U409, R2278_U141, R2278_U224);
  nand ginst2013 (R2278_U41, R2278_U228, R2278_U304);
  nand ginst2014 (R2278_U410, R2278_U140, R2278_U275);
  nand ginst2015 (R2278_U411, R2278_U144, R2278_U281);
  nand ginst2016 (R2278_U412, R2278_U143, R2278_U282);
  nand ginst2017 (R2278_U413, R2278_U147, R2278_U279);
  nand ginst2018 (R2278_U414, R2278_U146, R2278_U283);
  nand ginst2019 (R2278_U415, R2278_U150, R2278_U277);
  nand ginst2020 (R2278_U416, R2278_U149, R2278_U284);
  nand ginst2021 (R2278_U417, R2278_U153, R2278_U220);
  nand ginst2022 (R2278_U418, R2278_U152, R2278_U285);
  nand ginst2023 (R2278_U419, R2278_U156, R2278_U289);
  nand ginst2024 (R2278_U42, R2278_U401, R2278_U402);
  nand ginst2025 (R2278_U420, R2278_U155, R2278_U290);
  nand ginst2026 (R2278_U421, R2278_U159, R2278_U287);
  nand ginst2027 (R2278_U422, R2278_U158, R2278_U291);
  and ginst2028 (R2278_U43, R2278_U162, R2278_U178);
  and ginst2029 (R2278_U44, R2278_U179, R2278_U303);
  and ginst2030 (R2278_U45, R2278_U163, R2278_U182);
  and ginst2031 (R2278_U46, R2278_U301, R2278_U302);
  and ginst2032 (R2278_U47, INSTADDRPOINTER_REG_20__SCAN_IN, U2770);
  and ginst2033 (R2278_U48, R2278_U162, R2278_U178);
  and ginst2034 (R2278_U49, R2278_U179, R2278_U337);
  and ginst2035 (R2278_U5, R2278_U215, R2278_U217);
  and ginst2036 (R2278_U50, R2278_U163, R2278_U182, R2278_U301);
  and ginst2037 (R2278_U51, R2278_U185, R2278_U189);
  and ginst2038 (R2278_U52, R2278_U5, R2278_U51);
  and ginst2039 (R2278_U53, R2278_U186, R2278_U189);
  and ginst2040 (R2278_U54, R2278_U216, R2278_U293, R2278_U295, R2278_U296);
  and ginst2041 (R2278_U55, R2278_U209, R2278_U211, R2278_U213, R2278_U221);
  and ginst2042 (R2278_U56, R2278_U210, R2278_U294, R2278_U297, R2278_U298);
  and ginst2043 (R2278_U57, R2278_U13, R2278_U8);
  and ginst2044 (R2278_U58, R2278_U245, R2278_U332);
  and ginst2045 (R2278_U59, R2278_U320, R2278_U333, R2278_U58);
  and ginst2046 (R2278_U6, R2278_U225, R2278_U227);
  and ginst2047 (R2278_U60, R2278_U16, R2278_U259);
  and ginst2048 (R2278_U61, R2278_U260, R2278_U331);
  nand ginst2049 (R2278_U62, R2278_U363, R2278_U364);
  nand ginst2050 (R2278_U63, R2278_U368, R2278_U369);
  nand ginst2051 (R2278_U64, R2278_U375, R2278_U376);
  nand ginst2052 (R2278_U65, R2278_U380, R2278_U381);
  and ginst2053 (R2278_U66, R2278_U23, R2278_U25);
  and ginst2054 (R2278_U67, R2278_U243, R2278_U318);
  and ginst2055 (R2278_U68, R2278_U240, R2278_U315);
  and ginst2056 (R2278_U69, R2278_U238, R2278_U312);
  and ginst2057 (R2278_U7, R2278_U208, R2278_U6);
  and ginst2058 (R2278_U70, R2278_U236, R2278_U310);
  and ginst2059 (R2278_U71, R2278_U216, R2278_U293, R2278_U295, R2278_U296);
  nand ginst2060 (R2278_U72, R2278_U187, R2278_U26);
  nand ginst2061 (R2278_U73, R2278_U189, R2278_U27);
  and ginst2062 (R2278_U74, R2278_U349, R2278_U350);
  nand ginst2063 (R2278_U75, R2278_U183, R2278_U45, R2278_U46);
  nand ginst2064 (R2278_U76, R2278_U185, R2278_U26);
  and ginst2065 (R2278_U77, R2278_U351, R2278_U352);
  nand ginst2066 (R2278_U78, R2278_U165, R2278_U197);
  nand ginst2067 (R2278_U79, R2278_U162, R2278_U163);
  and ginst2068 (R2278_U8, R2278_U207, R2278_U7);
  and ginst2069 (R2278_U80, R2278_U353, R2278_U354);
  nand ginst2070 (R2278_U81, R2278_U195, R2278_U20);
  nand ginst2071 (R2278_U82, R2278_U164, R2278_U165);
  and ginst2072 (R2278_U83, R2278_U355, R2278_U356);
  nand ginst2073 (R2278_U84, R2278_U18, R2278_U193);
  nand ginst2074 (R2278_U85, R2278_U179, R2278_U20);
  and ginst2075 (R2278_U86, R2278_U357, R2278_U358);
  nand ginst2076 (R2278_U87, R2278_U175, R2278_U176);
  nand ginst2077 (R2278_U88, R2278_U178, R2278_U18);
  and ginst2078 (R2278_U89, R2278_U359, R2278_U360);
  and ginst2079 (R2278_U9, R2278_U231, R2278_U235);
  nand ginst2080 (R2278_U90, R2278_U172, R2278_U173);
  nand ginst2081 (R2278_U91, R2278_U166, R2278_U175);
  and ginst2082 (R2278_U92, R2278_U361, R2278_U362);
  not ginst2083 (R2278_U93, U2769);
  not ginst2084 (R2278_U94, INSTADDRPOINTER_REG_31__SCAN_IN);
  nand ginst2085 (R2278_U95, R2278_U330, R2278_U61);
  and ginst2086 (R2278_U96, R2278_U366, R2278_U367);
  nand ginst2087 (R2278_U97, R2278_U327, R2278_U329);
  and ginst2088 (R2278_U98, R2278_U371, R2278_U372);
  nand ginst2089 (R2278_U99, R2278_U169, R2278_U170);
  nand ginst2090 (R2337_U10, PHYADDRPOINTER_REG_1__SCAN_IN, PHYADDRPOINTER_REG_2__SCAN_IN, PHYADDRPOINTER_REG_3__SCAN_IN, PHYADDRPOINTER_REG_4__SCAN_IN, PHYADDRPOINTER_REG_5__SCAN_IN);
  nand ginst2091 (R2337_U100, PHYADDRPOINTER_REG_18__SCAN_IN, R2337_U120);
  nand ginst2092 (R2337_U101, PHYADDRPOINTER_REG_16__SCAN_IN, R2337_U118);
  nand ginst2093 (R2337_U102, PHYADDRPOINTER_REG_14__SCAN_IN, R2337_U116);
  nand ginst2094 (R2337_U103, PHYADDRPOINTER_REG_12__SCAN_IN, R2337_U114);
  nand ginst2095 (R2337_U104, PHYADDRPOINTER_REG_10__SCAN_IN, R2337_U112);
  not ginst2096 (R2337_U105, R2337_U94);
  not ginst2097 (R2337_U106, R2337_U16);
  not ginst2098 (R2337_U107, R2337_U93);
  not ginst2099 (R2337_U108, R2337_U10);
  not ginst2100 (R2337_U109, R2337_U92);
  not ginst2101 (R2337_U11, PHYADDRPOINTER_REG_7__SCAN_IN);
  not ginst2102 (R2337_U110, R2337_U13);
  not ginst2103 (R2337_U111, R2337_U91);
  not ginst2104 (R2337_U112, R2337_U17);
  not ginst2105 (R2337_U113, R2337_U104);
  not ginst2106 (R2337_U114, R2337_U20);
  not ginst2107 (R2337_U115, R2337_U103);
  not ginst2108 (R2337_U116, R2337_U23);
  not ginst2109 (R2337_U117, R2337_U102);
  not ginst2110 (R2337_U118, R2337_U26);
  not ginst2111 (R2337_U119, R2337_U101);
  not ginst2112 (R2337_U12, PHYADDRPOINTER_REG_6__SCAN_IN);
  not ginst2113 (R2337_U120, R2337_U29);
  not ginst2114 (R2337_U121, R2337_U100);
  not ginst2115 (R2337_U122, R2337_U32);
  not ginst2116 (R2337_U123, R2337_U99);
  not ginst2117 (R2337_U124, R2337_U35);
  not ginst2118 (R2337_U125, R2337_U98);
  not ginst2119 (R2337_U126, R2337_U38);
  not ginst2120 (R2337_U127, R2337_U97);
  not ginst2121 (R2337_U128, R2337_U41);
  not ginst2122 (R2337_U129, R2337_U43);
  nand ginst2123 (R2337_U13, R2337_U108, R2337_U81);
  not ginst2124 (R2337_U130, R2337_U45);
  not ginst2125 (R2337_U131, R2337_U47);
  not ginst2126 (R2337_U132, R2337_U49);
  not ginst2127 (R2337_U133, R2337_U96);
  nand ginst2128 (R2337_U134, PHYADDRPOINTER_REG_9__SCAN_IN, R2337_U91);
  nand ginst2129 (R2337_U135, R2337_U111, R2337_U15);
  nand ginst2130 (R2337_U136, PHYADDRPOINTER_REG_8__SCAN_IN, R2337_U13);
  nand ginst2131 (R2337_U137, R2337_U110, R2337_U14);
  nand ginst2132 (R2337_U138, PHYADDRPOINTER_REG_7__SCAN_IN, R2337_U92);
  nand ginst2133 (R2337_U139, R2337_U109, R2337_U11);
  not ginst2134 (R2337_U14, PHYADDRPOINTER_REG_8__SCAN_IN);
  nand ginst2135 (R2337_U140, PHYADDRPOINTER_REG_6__SCAN_IN, R2337_U10);
  nand ginst2136 (R2337_U141, R2337_U108, R2337_U12);
  nand ginst2137 (R2337_U142, PHYADDRPOINTER_REG_5__SCAN_IN, R2337_U93);
  nand ginst2138 (R2337_U143, R2337_U107, R2337_U6);
  nand ginst2139 (R2337_U144, PHYADDRPOINTER_REG_4__SCAN_IN, R2337_U16);
  nand ginst2140 (R2337_U145, R2337_U106, R2337_U7);
  nand ginst2141 (R2337_U146, PHYADDRPOINTER_REG_3__SCAN_IN, R2337_U94);
  nand ginst2142 (R2337_U147, R2337_U105, R2337_U8);
  nand ginst2143 (R2337_U148, PHYADDRPOINTER_REG_31__SCAN_IN, R2337_U96);
  nand ginst2144 (R2337_U149, R2337_U133, R2337_U95);
  not ginst2145 (R2337_U15, PHYADDRPOINTER_REG_9__SCAN_IN);
  nand ginst2146 (R2337_U150, PHYADDRPOINTER_REG_30__SCAN_IN, R2337_U49);
  nand ginst2147 (R2337_U151, R2337_U132, R2337_U50);
  nand ginst2148 (R2337_U152, PHYADDRPOINTER_REG_1__SCAN_IN, R2337_U9);
  nand ginst2149 (R2337_U153, PHYADDRPOINTER_REG_2__SCAN_IN, R2337_U5);
  nand ginst2150 (R2337_U154, PHYADDRPOINTER_REG_29__SCAN_IN, R2337_U47);
  nand ginst2151 (R2337_U155, R2337_U131, R2337_U48);
  nand ginst2152 (R2337_U156, PHYADDRPOINTER_REG_28__SCAN_IN, R2337_U45);
  nand ginst2153 (R2337_U157, R2337_U130, R2337_U46);
  nand ginst2154 (R2337_U158, PHYADDRPOINTER_REG_27__SCAN_IN, R2337_U43);
  nand ginst2155 (R2337_U159, R2337_U129, R2337_U44);
  nand ginst2156 (R2337_U16, PHYADDRPOINTER_REG_1__SCAN_IN, PHYADDRPOINTER_REG_2__SCAN_IN, PHYADDRPOINTER_REG_3__SCAN_IN);
  nand ginst2157 (R2337_U160, PHYADDRPOINTER_REG_26__SCAN_IN, R2337_U41);
  nand ginst2158 (R2337_U161, R2337_U128, R2337_U42);
  nand ginst2159 (R2337_U162, PHYADDRPOINTER_REG_25__SCAN_IN, R2337_U97);
  nand ginst2160 (R2337_U163, R2337_U127, R2337_U39);
  nand ginst2161 (R2337_U164, PHYADDRPOINTER_REG_24__SCAN_IN, R2337_U38);
  nand ginst2162 (R2337_U165, R2337_U126, R2337_U40);
  nand ginst2163 (R2337_U166, PHYADDRPOINTER_REG_23__SCAN_IN, R2337_U98);
  nand ginst2164 (R2337_U167, R2337_U125, R2337_U36);
  nand ginst2165 (R2337_U168, PHYADDRPOINTER_REG_22__SCAN_IN, R2337_U35);
  nand ginst2166 (R2337_U169, R2337_U124, R2337_U37);
  nand ginst2167 (R2337_U17, R2337_U110, R2337_U82);
  nand ginst2168 (R2337_U170, PHYADDRPOINTER_REG_21__SCAN_IN, R2337_U99);
  nand ginst2169 (R2337_U171, R2337_U123, R2337_U33);
  nand ginst2170 (R2337_U172, PHYADDRPOINTER_REG_20__SCAN_IN, R2337_U32);
  nand ginst2171 (R2337_U173, R2337_U122, R2337_U34);
  nand ginst2172 (R2337_U174, PHYADDRPOINTER_REG_19__SCAN_IN, R2337_U100);
  nand ginst2173 (R2337_U175, R2337_U121, R2337_U30);
  nand ginst2174 (R2337_U176, PHYADDRPOINTER_REG_18__SCAN_IN, R2337_U29);
  nand ginst2175 (R2337_U177, R2337_U120, R2337_U31);
  nand ginst2176 (R2337_U178, PHYADDRPOINTER_REG_17__SCAN_IN, R2337_U101);
  nand ginst2177 (R2337_U179, R2337_U119, R2337_U27);
  not ginst2178 (R2337_U18, PHYADDRPOINTER_REG_11__SCAN_IN);
  nand ginst2179 (R2337_U180, PHYADDRPOINTER_REG_16__SCAN_IN, R2337_U26);
  nand ginst2180 (R2337_U181, R2337_U118, R2337_U28);
  nand ginst2181 (R2337_U182, PHYADDRPOINTER_REG_15__SCAN_IN, R2337_U102);
  nand ginst2182 (R2337_U183, R2337_U117, R2337_U24);
  nand ginst2183 (R2337_U184, PHYADDRPOINTER_REG_14__SCAN_IN, R2337_U23);
  nand ginst2184 (R2337_U185, R2337_U116, R2337_U25);
  nand ginst2185 (R2337_U186, PHYADDRPOINTER_REG_13__SCAN_IN, R2337_U103);
  nand ginst2186 (R2337_U187, R2337_U115, R2337_U21);
  nand ginst2187 (R2337_U188, PHYADDRPOINTER_REG_12__SCAN_IN, R2337_U20);
  nand ginst2188 (R2337_U189, R2337_U114, R2337_U22);
  not ginst2189 (R2337_U19, PHYADDRPOINTER_REG_10__SCAN_IN);
  nand ginst2190 (R2337_U190, PHYADDRPOINTER_REG_11__SCAN_IN, R2337_U104);
  nand ginst2191 (R2337_U191, R2337_U113, R2337_U18);
  nand ginst2192 (R2337_U192, PHYADDRPOINTER_REG_10__SCAN_IN, R2337_U17);
  nand ginst2193 (R2337_U193, R2337_U112, R2337_U19);
  nand ginst2194 (R2337_U20, R2337_U112, R2337_U83);
  not ginst2195 (R2337_U21, PHYADDRPOINTER_REG_13__SCAN_IN);
  not ginst2196 (R2337_U22, PHYADDRPOINTER_REG_12__SCAN_IN);
  nand ginst2197 (R2337_U23, R2337_U114, R2337_U84);
  not ginst2198 (R2337_U24, PHYADDRPOINTER_REG_15__SCAN_IN);
  not ginst2199 (R2337_U25, PHYADDRPOINTER_REG_14__SCAN_IN);
  nand ginst2200 (R2337_U26, R2337_U116, R2337_U85);
  not ginst2201 (R2337_U27, PHYADDRPOINTER_REG_17__SCAN_IN);
  not ginst2202 (R2337_U28, PHYADDRPOINTER_REG_16__SCAN_IN);
  nand ginst2203 (R2337_U29, R2337_U118, R2337_U86);
  not ginst2204 (R2337_U30, PHYADDRPOINTER_REG_19__SCAN_IN);
  not ginst2205 (R2337_U31, PHYADDRPOINTER_REG_18__SCAN_IN);
  nand ginst2206 (R2337_U32, R2337_U120, R2337_U87);
  not ginst2207 (R2337_U33, PHYADDRPOINTER_REG_21__SCAN_IN);
  not ginst2208 (R2337_U34, PHYADDRPOINTER_REG_20__SCAN_IN);
  nand ginst2209 (R2337_U35, R2337_U122, R2337_U88);
  not ginst2210 (R2337_U36, PHYADDRPOINTER_REG_23__SCAN_IN);
  not ginst2211 (R2337_U37, PHYADDRPOINTER_REG_22__SCAN_IN);
  nand ginst2212 (R2337_U38, R2337_U124, R2337_U89);
  not ginst2213 (R2337_U39, PHYADDRPOINTER_REG_25__SCAN_IN);
  not ginst2214 (R2337_U40, PHYADDRPOINTER_REG_24__SCAN_IN);
  nand ginst2215 (R2337_U41, R2337_U126, R2337_U90);
  not ginst2216 (R2337_U42, PHYADDRPOINTER_REG_26__SCAN_IN);
  nand ginst2217 (R2337_U43, PHYADDRPOINTER_REG_26__SCAN_IN, R2337_U128);
  not ginst2218 (R2337_U44, PHYADDRPOINTER_REG_27__SCAN_IN);
  nand ginst2219 (R2337_U45, PHYADDRPOINTER_REG_27__SCAN_IN, R2337_U129);
  not ginst2220 (R2337_U46, PHYADDRPOINTER_REG_28__SCAN_IN);
  nand ginst2221 (R2337_U47, PHYADDRPOINTER_REG_28__SCAN_IN, R2337_U130);
  not ginst2222 (R2337_U48, PHYADDRPOINTER_REG_29__SCAN_IN);
  nand ginst2223 (R2337_U49, PHYADDRPOINTER_REG_29__SCAN_IN, R2337_U131);
  not ginst2224 (R2337_U5, PHYADDRPOINTER_REG_1__SCAN_IN);
  not ginst2225 (R2337_U50, PHYADDRPOINTER_REG_30__SCAN_IN);
  nand ginst2226 (R2337_U51, R2337_U134, R2337_U135);
  nand ginst2227 (R2337_U52, R2337_U136, R2337_U137);
  nand ginst2228 (R2337_U53, R2337_U138, R2337_U139);
  nand ginst2229 (R2337_U54, R2337_U140, R2337_U141);
  nand ginst2230 (R2337_U55, R2337_U142, R2337_U143);
  nand ginst2231 (R2337_U56, R2337_U144, R2337_U145);
  nand ginst2232 (R2337_U57, R2337_U146, R2337_U147);
  nand ginst2233 (R2337_U58, R2337_U148, R2337_U149);
  nand ginst2234 (R2337_U59, R2337_U150, R2337_U151);
  not ginst2235 (R2337_U6, PHYADDRPOINTER_REG_5__SCAN_IN);
  nand ginst2236 (R2337_U60, R2337_U152, R2337_U153);
  nand ginst2237 (R2337_U61, R2337_U154, R2337_U155);
  nand ginst2238 (R2337_U62, R2337_U156, R2337_U157);
  nand ginst2239 (R2337_U63, R2337_U158, R2337_U159);
  nand ginst2240 (R2337_U64, R2337_U160, R2337_U161);
  nand ginst2241 (R2337_U65, R2337_U162, R2337_U163);
  nand ginst2242 (R2337_U66, R2337_U164, R2337_U165);
  nand ginst2243 (R2337_U67, R2337_U166, R2337_U167);
  nand ginst2244 (R2337_U68, R2337_U168, R2337_U169);
  nand ginst2245 (R2337_U69, R2337_U170, R2337_U171);
  not ginst2246 (R2337_U7, PHYADDRPOINTER_REG_4__SCAN_IN);
  nand ginst2247 (R2337_U70, R2337_U172, R2337_U173);
  nand ginst2248 (R2337_U71, R2337_U174, R2337_U175);
  nand ginst2249 (R2337_U72, R2337_U176, R2337_U177);
  nand ginst2250 (R2337_U73, R2337_U178, R2337_U179);
  nand ginst2251 (R2337_U74, R2337_U180, R2337_U181);
  nand ginst2252 (R2337_U75, R2337_U182, R2337_U183);
  nand ginst2253 (R2337_U76, R2337_U184, R2337_U185);
  nand ginst2254 (R2337_U77, R2337_U186, R2337_U187);
  nand ginst2255 (R2337_U78, R2337_U188, R2337_U189);
  nand ginst2256 (R2337_U79, R2337_U190, R2337_U191);
  not ginst2257 (R2337_U8, PHYADDRPOINTER_REG_3__SCAN_IN);
  nand ginst2258 (R2337_U80, R2337_U192, R2337_U193);
  and ginst2259 (R2337_U81, PHYADDRPOINTER_REG_6__SCAN_IN, PHYADDRPOINTER_REG_7__SCAN_IN);
  and ginst2260 (R2337_U82, PHYADDRPOINTER_REG_8__SCAN_IN, PHYADDRPOINTER_REG_9__SCAN_IN);
  and ginst2261 (R2337_U83, PHYADDRPOINTER_REG_10__SCAN_IN, PHYADDRPOINTER_REG_11__SCAN_IN);
  and ginst2262 (R2337_U84, PHYADDRPOINTER_REG_12__SCAN_IN, PHYADDRPOINTER_REG_13__SCAN_IN);
  and ginst2263 (R2337_U85, PHYADDRPOINTER_REG_14__SCAN_IN, PHYADDRPOINTER_REG_15__SCAN_IN);
  and ginst2264 (R2337_U86, PHYADDRPOINTER_REG_16__SCAN_IN, PHYADDRPOINTER_REG_17__SCAN_IN);
  and ginst2265 (R2337_U87, PHYADDRPOINTER_REG_18__SCAN_IN, PHYADDRPOINTER_REG_19__SCAN_IN);
  and ginst2266 (R2337_U88, PHYADDRPOINTER_REG_20__SCAN_IN, PHYADDRPOINTER_REG_21__SCAN_IN);
  and ginst2267 (R2337_U89, PHYADDRPOINTER_REG_22__SCAN_IN, PHYADDRPOINTER_REG_23__SCAN_IN);
  not ginst2268 (R2337_U9, PHYADDRPOINTER_REG_2__SCAN_IN);
  and ginst2269 (R2337_U90, PHYADDRPOINTER_REG_24__SCAN_IN, PHYADDRPOINTER_REG_25__SCAN_IN);
  nand ginst2270 (R2337_U91, PHYADDRPOINTER_REG_8__SCAN_IN, R2337_U110);
  nand ginst2271 (R2337_U92, PHYADDRPOINTER_REG_6__SCAN_IN, R2337_U108);
  nand ginst2272 (R2337_U93, PHYADDRPOINTER_REG_4__SCAN_IN, R2337_U106);
  nand ginst2273 (R2337_U94, PHYADDRPOINTER_REG_1__SCAN_IN, PHYADDRPOINTER_REG_2__SCAN_IN);
  not ginst2274 (R2337_U95, PHYADDRPOINTER_REG_31__SCAN_IN);
  nand ginst2275 (R2337_U96, PHYADDRPOINTER_REG_30__SCAN_IN, R2337_U132);
  nand ginst2276 (R2337_U97, PHYADDRPOINTER_REG_24__SCAN_IN, R2337_U126);
  nand ginst2277 (R2337_U98, PHYADDRPOINTER_REG_22__SCAN_IN, R2337_U124);
  nand ginst2278 (R2337_U99, PHYADDRPOINTER_REG_20__SCAN_IN, R2337_U122);
  and ginst2279 (R2358_U10, R2358_U253, R2358_U304);
  and ginst2280 (R2358_U100, R2358_U284, R2358_U285);
  nand ginst2281 (R2358_U101, R2358_U618, R2358_U619);
  and ginst2282 (R2358_U102, R2358_U283, R2358_U293);
  nand ginst2283 (R2358_U103, R2358_U620, R2358_U621);
  and ginst2284 (R2358_U104, R2358_U319, R2358_U320);
  nand ginst2285 (R2358_U105, R2358_U622, R2358_U623);
  and ginst2286 (R2358_U106, R2358_U321, R2358_U322);
  nand ginst2287 (R2358_U107, R2358_U624, R2358_U625);
  and ginst2288 (R2358_U108, R2358_U323, R2358_U324);
  nand ginst2289 (R2358_U109, R2358_U626, R2358_U627);
  and ginst2290 (R2358_U11, R2358_U301, R2358_U303);
  nand ginst2291 (R2358_U110, R2358_U631, R2358_U632);
  and ginst2292 (R2358_U111, R2358_U232, R2358_U233);
  nand ginst2293 (R2358_U112, R2358_U633, R2358_U634);
  and ginst2294 (R2358_U113, R2358_U316, R2358_U317);
  nand ginst2295 (R2358_U114, R2358_U635, R2358_U636);
  and ginst2296 (R2358_U115, R2358_U294, R2358_U295);
  nand ginst2297 (R2358_U116, R2358_U637, R2358_U638);
  and ginst2298 (R2358_U117, R2358_U296, R2358_U59);
  nand ginst2299 (R2358_U118, R2358_U639, R2358_U640);
  nand ginst2300 (R2358_U119, R2358_U644, R2358_U645);
  and ginst2301 (R2358_U12, R2358_U7, R2358_U8);
  nand ginst2302 (R2358_U120, R2358_U649, R2358_U650);
  and ginst2303 (R2358_U121, R2358_U310, R2358_U53);
  nand ginst2304 (R2358_U122, R2358_U651, R2358_U652);
  and ginst2305 (R2358_U123, R2358_U232, R2358_U235);
  and ginst2306 (R2358_U124, R2358_U229, R2358_U231);
  and ginst2307 (R2358_U125, R2358_U243, R2358_U244);
  and ginst2308 (R2358_U126, R2358_U245, R2358_U249);
  and ginst2309 (R2358_U127, R2358_U222, R2358_U245);
  and ginst2310 (R2358_U128, R2358_U265, R2358_U31);
  and ginst2311 (R2358_U129, R2358_U230, R2358_U231);
  and ginst2312 (R2358_U13, R2358_U527, R2358_U528);
  and ginst2313 (R2358_U130, R2358_U282, R2358_U285);
  and ginst2314 (R2358_U131, R2358_U288, R2358_U289);
  and ginst2315 (R2358_U132, R2358_U279, R2358_U281);
  and ginst2316 (R2358_U133, R2358_U323, R2358_U326);
  and ginst2317 (R2358_U134, R2358_U319, R2358_U322);
  and ginst2318 (R2358_U135, R2358_U277, R2358_U279);
  and ginst2319 (R2358_U136, R2358_U10, R2358_U11);
  and ginst2320 (R2358_U137, R2358_U425, R2358_U432);
  and ginst2321 (R2358_U138, R2358_U224, R2358_U310);
  and ginst2322 (R2358_U139, R2358_U311, R2358_U415);
  and ginst2323 (R2358_U14, R2358_U378, R2358_U379);
  and ginst2324 (R2358_U140, R2358_U411, R2358_U420);
  and ginst2325 (R2358_U141, R2358_U319, R2358_U322);
  and ginst2326 (R2358_U142, R2358_U313, R2358_U317);
  and ginst2327 (R2358_U143, R2358_U12, R2358_U426);
  and ginst2328 (R2358_U144, R2358_U278, R2358_U402);
  and ginst2329 (R2358_U145, R2358_U144, R2358_U406, R2358_U430);
  and ginst2330 (R2358_U146, R2358_U411, R2358_U420);
  and ginst2331 (R2358_U147, R2358_U313, R2358_U317);
  and ginst2332 (R2358_U148, R2358_U149, R2358_U7);
  and ginst2333 (R2358_U149, R2358_U147, R2358_U9);
  and ginst2334 (R2358_U15, R2358_U374, R2358_U376);
  and ginst2335 (R2358_U150, R2358_U422, R2358_U439);
  and ginst2336 (R2358_U151, R2358_U279, R2358_U5);
  and ginst2337 (R2358_U152, R2358_U282, R2358_U285, R2358_U293);
  and ginst2338 (R2358_U153, R2358_U287, R2358_U289);
  and ginst2339 (R2358_U154, R2358_U283, R2358_U284);
  and ginst2340 (R2358_U155, R2358_U156, R2358_U434);
  and ginst2341 (R2358_U156, R2358_U324, R2358_U6);
  and ginst2342 (R2358_U157, R2358_U418, R2358_U46);
  and ginst2343 (R2358_U158, R2358_U326, R2358_U6);
  and ginst2344 (R2358_U159, R2358_U313, R2358_U9);
  and ginst2345 (R2358_U16, R2358_U367, R2358_U370);
  and ginst2346 (R2358_U160, R2358_U224, R2358_U299, R2358_U300);
  and ginst2347 (R2358_U161, R2358_U227, R2358_U369);
  and ginst2348 (R2358_U162, R2358_U302, R2358_U303);
  and ginst2349 (R2358_U163, R2358_U307, R2358_U375);
  not ginst2350 (R2358_U164, U2612);
  and ginst2351 (R2358_U165, R2358_U443, R2358_U444);
  not ginst2352 (R2358_U166, U2610);
  not ginst2353 (R2358_U167, U2609);
  not ginst2354 (R2358_U168, U2667);
  not ginst2355 (R2358_U169, U2668);
  and ginst2356 (R2358_U17, R2358_U359, R2358_U360);
  not ginst2357 (R2358_U170, U2670);
  not ginst2358 (R2358_U171, U2671);
  not ginst2359 (R2358_U172, U2672);
  not ginst2360 (R2358_U173, U2669);
  not ginst2361 (R2358_U174, U2611);
  nand ginst2362 (R2358_U175, R2358_U255, R2358_U49);
  nand ginst2363 (R2358_U176, R2358_U126, R2358_U250, R2358_U251);
  nand ginst2364 (R2358_U177, R2358_U247, R2358_U257);
  nand ginst2365 (R2358_U178, R2358_U230, R2358_U240);
  not ginst2366 (R2358_U179, U2651);
  and ginst2367 (R2358_U18, R2358_U352, R2358_U354);
  and ginst2368 (R2358_U180, R2358_U504, R2358_U505);
  not ginst2369 (R2358_U181, U2613);
  not ginst2370 (R2358_U182, U2614);
  not ginst2371 (R2358_U183, U2617);
  not ginst2372 (R2358_U184, U2615);
  not ginst2373 (R2358_U185, U2616);
  not ginst2374 (R2358_U186, U2618);
  not ginst2375 (R2358_U187, U2664);
  not ginst2376 (R2358_U188, U2665);
  not ginst2377 (R2358_U189, U2666);
  and ginst2378 (R2358_U19, R2358_U335, R2358_U336);
  not ginst2379 (R2358_U190, U2663);
  not ginst2380 (R2358_U191, U2658);
  not ginst2381 (R2358_U192, U2659);
  not ginst2382 (R2358_U193, U2660);
  not ginst2383 (R2358_U194, U2661);
  not ginst2384 (R2358_U195, U2662);
  not ginst2385 (R2358_U196, U2654);
  not ginst2386 (R2358_U197, U2655);
  not ginst2387 (R2358_U198, U2656);
  not ginst2388 (R2358_U199, U2657);
  and ginst2389 (R2358_U20, R2358_U274, R2358_U276);
  not ginst2390 (R2358_U200, U2652);
  not ginst2391 (R2358_U201, U2653);
  nand ginst2392 (R2358_U202, R2358_U145, R2358_U429);
  nand ginst2393 (R2358_U203, R2358_U292, R2358_U332);
  nand ginst2394 (R2358_U204, R2358_U337, R2358_U338);
  nand ginst2395 (R2358_U205, R2358_U153, R2358_U340);
  nand ginst2396 (R2358_U206, R2358_U285, R2358_U344);
  nand ginst2397 (R2358_U207, R2358_U283, R2358_U342);
  nand ginst2398 (R2358_U208, R2358_U150, R2358_U421);
  nand ginst2399 (R2358_U209, R2358_U321, R2358_U347);
  and ginst2400 (R2358_U21, R2358_U262, R2358_U266);
  nand ginst2401 (R2358_U210, R2358_U345, R2358_U437);
  nand ginst2402 (R2358_U211, R2358_U325, R2358_U350);
  nand ginst2403 (R2358_U212, R2358_U236, R2358_U268);
  nand ginst2404 (R2358_U213, R2358_U409, R2358_U412);
  nand ginst2405 (R2358_U214, R2358_U356, R2358_U59);
  nand ginst2406 (R2358_U215, R2358_U61, R2358_U70);
  nand ginst2407 (R2358_U216, R2358_U361, R2358_U53);
  nand ginst2408 (R2358_U217, R2358_U137, R2358_U431);
  nand ginst2409 (R2358_U218, R2358_U235, R2358_U236);
  nand ginst2410 (R2358_U219, R2358_U138, R2358_U139, R2358_U217);
  not ginst2411 (R2358_U22, U2352);
  not ginst2412 (R2358_U220, R2358_U211);
  not ginst2413 (R2358_U221, R2358_U206);
  nand ginst2414 (R2358_U222, R2358_U403, R2358_U404);
  not ginst2415 (R2358_U223, R2358_U51);
  nand ginst2416 (R2358_U224, R2358_U521, R2358_U54);
  not ginst2417 (R2358_U225, R2358_U46);
  nand ginst2418 (R2358_U226, R2358_U329, R2358_U349);
  nand ginst2419 (R2358_U227, R2358_U79, U2636);
  not ginst2420 (R2358_U228, R2358_U31);
  nand ginst2421 (R2358_U229, R2358_U28, R2358_U479, R2358_U480);
  not ginst2422 (R2358_U23, U2643);
  nand ginst2423 (R2358_U230, R2358_U485, U2647);
  nand ginst2424 (R2358_U231, R2358_U30, R2358_U481, R2358_U482);
  nand ginst2425 (R2358_U232, R2358_U27, R2358_U475, R2358_U476);
  nand ginst2426 (R2358_U233, R2358_U471, U2649);
  nand ginst2427 (R2358_U234, R2358_U468, U2648);
  nand ginst2428 (R2358_U235, R2358_U29, R2358_U477, R2358_U478);
  nand ginst2429 (R2358_U236, R2358_U474, U2650);
  nand ginst2430 (R2358_U237, R2358_U22, R2358_U236);
  nand ginst2431 (R2358_U238, R2358_U123, R2358_U237);
  nand ginst2432 (R2358_U239, R2358_U233, R2358_U234, R2358_U238);
  not ginst2433 (R2358_U24, U2644);
  nand ginst2434 (R2358_U240, R2358_U124, R2358_U239);
  not ginst2435 (R2358_U241, R2358_U178);
  nand ginst2436 (R2358_U242, R2358_U23, R2358_U451, R2358_U452);
  nand ginst2437 (R2358_U243, R2358_U25, R2358_U462, R2358_U463);
  nand ginst2438 (R2358_U244, R2358_U26, R2358_U464, R2358_U465);
  nand ginst2439 (R2358_U245, R2358_U450, U2643);
  nand ginst2440 (R2358_U246, R2358_U458, U2645);
  nand ginst2441 (R2358_U247, R2358_U461, U2646);
  nand ginst2442 (R2358_U248, R2358_U246, R2358_U247);
  nand ginst2443 (R2358_U249, R2358_U222, R2358_U243, R2358_U248);
  not ginst2444 (R2358_U25, U2645);
  nand ginst2445 (R2358_U250, R2358_U125, R2358_U178, R2358_U222);
  nand ginst2446 (R2358_U251, R2358_U228, R2358_U242);
  not ginst2447 (R2358_U252, R2358_U176);
  nand ginst2448 (R2358_U253, R2358_U32, R2358_U486, R2358_U487);
  not ginst2449 (R2358_U254, R2358_U49);
  nand ginst2450 (R2358_U255, R2358_U176, R2358_U253);
  not ginst2451 (R2358_U256, R2358_U175);
  nand ginst2452 (R2358_U257, R2358_U178, R2358_U244);
  not ginst2453 (R2358_U258, R2358_U177);
  nand ginst2454 (R2358_U259, R2358_U177, R2358_U243);
  not ginst2455 (R2358_U26, U2646);
  not ginst2456 (R2358_U260, R2358_U34);
  nand ginst2457 (R2358_U261, R2358_U260, R2358_U31);
  nand ginst2458 (R2358_U262, R2358_U127, R2358_U261);
  nand ginst2459 (R2358_U263, R2358_U24, R2358_U455);
  nand ginst2460 (R2358_U264, R2358_U263, R2358_U34);
  nand ginst2461 (R2358_U265, R2358_U242, R2358_U245);
  nand ginst2462 (R2358_U266, R2358_U128, R2358_U264);
  nand ginst2463 (R2358_U267, R2358_U24, R2358_U455);
  nand ginst2464 (R2358_U268, R2358_U235, U2352);
  not ginst2465 (R2358_U269, R2358_U212);
  not ginst2466 (R2358_U27, U2649);
  nand ginst2467 (R2358_U270, R2358_U212, R2358_U232);
  not ginst2468 (R2358_U271, R2358_U64);
  not ginst2469 (R2358_U272, R2358_U65);
  nand ginst2470 (R2358_U273, R2358_U234, R2358_U65);
  nand ginst2471 (R2358_U274, R2358_U129, R2358_U273);
  nand ginst2472 (R2358_U275, R2358_U230, R2358_U231);
  nand ginst2473 (R2358_U276, R2358_U234, R2358_U275, R2358_U65);
  nand ginst2474 (R2358_U277, R2358_U35, R2358_U562, R2358_U563);
  nand ginst2475 (R2358_U278, R2358_U580, U2620);
  nand ginst2476 (R2358_U279, R2358_U40, R2358_U564, R2358_U565);
  not ginst2477 (R2358_U28, U2648);
  nand ginst2478 (R2358_U280, R2358_U595, U2621);
  nand ginst2479 (R2358_U281, R2358_U38, R2358_U554, R2358_U555);
  nand ginst2480 (R2358_U282, R2358_U39, R2358_U556, R2358_U557);
  nand ginst2481 (R2358_U283, R2358_U583, U2625);
  nand ginst2482 (R2358_U284, R2358_U586, U2624);
  nand ginst2483 (R2358_U285, R2358_U37, R2358_U558, R2358_U559);
  nand ginst2484 (R2358_U286, R2358_U283, R2358_U284);
  nand ginst2485 (R2358_U287, R2358_U130, R2358_U286);
  nand ginst2486 (R2358_U288, R2358_U592, U2622);
  nand ginst2487 (R2358_U289, R2358_U589, U2623);
  not ginst2488 (R2358_U29, U2650);
  nand ginst2489 (R2358_U290, R2358_U131, R2358_U287);
  nand ginst2490 (R2358_U291, R2358_U132, R2358_U290);
  not ginst2491 (R2358_U292, R2358_U63);
  nand ginst2492 (R2358_U293, R2358_U36, R2358_U560, R2358_U561);
  nand ginst2493 (R2358_U294, R2358_U535, R2358_U536, R2358_U57);
  nand ginst2494 (R2358_U295, R2358_U604, U2632);
  nand ginst2495 (R2358_U296, R2358_U537, R2358_U538, R2358_U58);
  not ginst2496 (R2358_U297, R2358_U59);
  not ginst2497 (R2358_U298, R2358_U61);
  nand ginst2498 (R2358_U299, R2358_U13, R2358_U71);
  not ginst2499 (R2358_U30, U2647);
  nand ginst2500 (R2358_U300, R2358_U81, U2635);
  nand ginst2501 (R2358_U301, R2358_U48, R2358_U509, R2358_U510);
  nand ginst2502 (R2358_U302, R2358_U515, U2639);
  nand ginst2503 (R2358_U303, R2358_U47, R2358_U511, R2358_U512);
  nand ginst2504 (R2358_U304, R2358_U33, R2358_U442);
  nand ginst2505 (R2358_U305, R2358_U76, U2641);
  not ginst2506 (R2358_U306, R2358_U74);
  nand ginst2507 (R2358_U307, R2358_U518, U2640);
  not ginst2508 (R2358_U308, R2358_U217);
  not ginst2509 (R2358_U309, R2358_U53);
  nand ginst2510 (R2358_U31, R2358_U77, U2644);
  nand ginst2511 (R2358_U310, R2358_U52, R2358_U522, R2358_U523);
  nand ginst2512 (R2358_U311, R2358_U50, R2358_U526);
  not ginst2513 (R2358_U312, R2358_U67);
  nand ginst2514 (R2358_U313, R2358_U539, R2358_U540, R2358_U60);
  not ginst2515 (R2358_U314, R2358_U70);
  not ginst2516 (R2358_U315, R2358_U213);
  nand ginst2517 (R2358_U316, R2358_U598, U2631);
  nand ginst2518 (R2358_U317, R2358_U541, R2358_U542, R2358_U56);
  not ginst2519 (R2358_U318, R2358_U68);
  nand ginst2520 (R2358_U319, R2358_U41, R2358_U543, R2358_U544);
  not ginst2521 (R2358_U32, U2642);
  nand ginst2522 (R2358_U320, R2358_U568, U2626);
  nand ginst2523 (R2358_U321, R2358_U571, U2627);
  nand ginst2524 (R2358_U322, R2358_U42, R2358_U545, R2358_U546);
  nand ginst2525 (R2358_U323, R2358_U574, U2628);
  nand ginst2526 (R2358_U324, R2358_U43, R2358_U547, R2358_U548);
  nand ginst2527 (R2358_U325, R2358_U44, R2358_U549, R2358_U550);
  nand ginst2528 (R2358_U326, R2358_U577, U2629);
  nand ginst2529 (R2358_U327, R2358_U225, R2358_U325);
  nand ginst2530 (R2358_U328, R2358_U321, R2358_U437);
  nand ginst2531 (R2358_U329, R2358_U45, R2358_U553);
  not ginst2532 (R2358_U33, U2641);
  not ginst2533 (R2358_U330, R2358_U202);
  not ginst2534 (R2358_U331, R2358_U208);
  nand ginst2535 (R2358_U332, R2358_U151, R2358_U208);
  not ginst2536 (R2358_U333, R2358_U203);
  nand ginst2537 (R2358_U334, R2358_U229, R2358_U234);
  nand ginst2538 (R2358_U335, R2358_U271, R2358_U334);
  nand ginst2539 (R2358_U336, R2358_U234, R2358_U272);
  nand ginst2540 (R2358_U337, R2358_U281, R2358_U290);
  nand ginst2541 (R2358_U338, R2358_U208, R2358_U5);
  not ginst2542 (R2358_U339, R2358_U204);
  nand ginst2543 (R2358_U34, R2358_U246, R2358_U259);
  nand ginst2544 (R2358_U340, R2358_U152, R2358_U208);
  not ginst2545 (R2358_U341, R2358_U205);
  nand ginst2546 (R2358_U342, R2358_U208, R2358_U293);
  not ginst2547 (R2358_U343, R2358_U207);
  nand ginst2548 (R2358_U344, R2358_U154, R2358_U342);
  nand ginst2549 (R2358_U345, R2358_U155, R2358_U433);
  not ginst2550 (R2358_U346, R2358_U210);
  nand ginst2551 (R2358_U347, R2358_U210, R2358_U322);
  not ginst2552 (R2358_U348, R2358_U209);
  nand ginst2553 (R2358_U349, R2358_U157, R2358_U416);
  not ginst2554 (R2358_U35, U2620);
  nand ginst2555 (R2358_U350, R2358_U226, R2358_U326);
  nand ginst2556 (R2358_U351, R2358_U318, R2358_U46);
  nand ginst2557 (R2358_U352, R2358_U158, R2358_U351);
  nand ginst2558 (R2358_U353, R2358_U325, R2358_U326);
  nand ginst2559 (R2358_U354, R2358_U226, R2358_U353);
  not ginst2560 (R2358_U355, R2358_U215);
  nand ginst2561 (R2358_U356, R2358_U215, R2358_U296);
  not ginst2562 (R2358_U357, R2358_U214);
  nand ginst2563 (R2358_U358, R2358_U313, R2358_U61);
  nand ginst2564 (R2358_U359, R2358_U312, R2358_U358);
  not ginst2565 (R2358_U36, U2625);
  nand ginst2566 (R2358_U360, R2358_U314, R2358_U61);
  nand ginst2567 (R2358_U361, R2358_U217, R2358_U310);
  not ginst2568 (R2358_U362, R2358_U216);
  nand ginst2569 (R2358_U363, R2358_U50, R2358_U526);
  nand ginst2570 (R2358_U364, R2358_U216, R2358_U363);
  not ginst2571 (R2358_U365, R2358_U72);
  nand ginst2572 (R2358_U366, R2358_U227, R2358_U365);
  nand ginst2573 (R2358_U367, R2358_U160, R2358_U366);
  nand ginst2574 (R2358_U368, R2358_U224, R2358_U72);
  nand ginst2575 (R2358_U369, R2358_U299, R2358_U300);
  not ginst2576 (R2358_U37, U2624);
  nand ginst2577 (R2358_U370, R2358_U161, R2358_U368);
  nand ginst2578 (R2358_U371, R2358_U50, R2358_U526);
  not ginst2579 (R2358_U372, R2358_U75);
  nand ginst2580 (R2358_U373, R2358_U307, R2358_U75);
  nand ginst2581 (R2358_U374, R2358_U162, R2358_U373);
  nand ginst2582 (R2358_U375, R2358_U302, R2358_U303);
  nand ginst2583 (R2358_U376, R2358_U163, R2358_U75);
  nand ginst2584 (R2358_U377, R2358_U301, R2358_U307);
  nand ginst2585 (R2358_U378, R2358_U306, R2358_U377);
  nand ginst2586 (R2358_U379, R2358_U307, R2358_U372);
  not ginst2587 (R2358_U38, U2622);
  not ginst2588 (R2358_U380, R2358_U218);
  nand ginst2589 (R2358_U381, R2358_U253, R2358_U49);
  nand ginst2590 (R2358_U382, R2358_U267, R2358_U31);
  nand ginst2591 (R2358_U383, R2358_U243, R2358_U246);
  nand ginst2592 (R2358_U384, R2358_U244, R2358_U247);
  nand ginst2593 (R2358_U385, R2358_U277, R2358_U278);
  nand ginst2594 (R2358_U386, R2358_U279, R2358_U280);
  nand ginst2595 (R2358_U387, R2358_U281, R2358_U288);
  nand ginst2596 (R2358_U388, R2358_U282, R2358_U289);
  nand ginst2597 (R2358_U389, R2358_U284, R2358_U285);
  not ginst2598 (R2358_U39, U2623);
  nand ginst2599 (R2358_U390, R2358_U283, R2358_U293);
  nand ginst2600 (R2358_U391, R2358_U319, R2358_U320);
  nand ginst2601 (R2358_U392, R2358_U321, R2358_U322);
  nand ginst2602 (R2358_U393, R2358_U323, R2358_U324);
  nand ginst2603 (R2358_U394, R2358_U329, R2358_U46);
  nand ginst2604 (R2358_U395, R2358_U232, R2358_U233);
  nand ginst2605 (R2358_U396, R2358_U316, R2358_U317);
  nand ginst2606 (R2358_U397, R2358_U294, R2358_U295);
  nand ginst2607 (R2358_U398, R2358_U296, R2358_U59);
  nand ginst2608 (R2358_U399, R2358_U224, R2358_U227);
  not ginst2609 (R2358_U40, U2621);
  nand ginst2610 (R2358_U400, R2358_U371, R2358_U51);
  nand ginst2611 (R2358_U401, R2358_U310, R2358_U53);
  nand ginst2612 (R2358_U402, R2358_U277, R2358_U63);
  nand ginst2613 (R2358_U403, R2358_U242, R2358_U77);
  nand ginst2614 (R2358_U404, R2358_U242, U2644);
  nand ginst2615 (R2358_U405, R2358_U518, U2640);
  nand ginst2616 (R2358_U406, R2358_U62, R2358_U8);
  nand ginst2617 (R2358_U407, R2358_U297, R2358_U9);
  nand ginst2618 (R2358_U408, R2358_U298, R2358_U9);
  nand ginst2619 (R2358_U409, R2358_U159, R2358_U67);
  not ginst2620 (R2358_U41, U2626);
  nand ginst2621 (R2358_U410, R2358_U223, R2358_U224, R2358_U299);
  nand ginst2622 (R2358_U411, R2358_U224, R2358_U299, R2358_U309, R2358_U311);
  not ginst2623 (R2358_U412, R2358_U69);
  nand ginst2624 (R2358_U413, R2358_U10, R2358_U176);
  nand ginst2625 (R2358_U414, R2358_U254, R2358_U304);
  nand ginst2626 (R2358_U415, R2358_U13, R2358_U71);
  nand ginst2627 (R2358_U416, R2358_U426, R2358_U67);
  nand ginst2628 (R2358_U417, R2358_U317, R2358_U69);
  not ginst2629 (R2358_U418, R2358_U66);
  nand ginst2630 (R2358_U419, R2358_U13, R2358_U71);
  not ginst2631 (R2358_U42, U2627);
  nand ginst2632 (R2358_U420, R2358_U419, R2358_U427, R2358_U428);
  nand ginst2633 (R2358_U421, R2358_U148, R2358_U67);
  nand ginst2634 (R2358_U422, R2358_U66, R2358_U7);
  not ginst2635 (R2358_U423, R2358_U73);
  nand ginst2636 (R2358_U424, R2358_U302, R2358_U405);
  nand ginst2637 (R2358_U425, R2358_U303, R2358_U424);
  not ginst2638 (R2358_U426, R2358_U55);
  nand ginst2639 (R2358_U427, R2358_U227, R2358_U71);
  nand ginst2640 (R2358_U428, R2358_U227, R2358_U534);
  nand ginst2641 (R2358_U429, R2358_U143, R2358_U435);
  not ginst2642 (R2358_U43, U2628);
  nand ginst2643 (R2358_U430, R2358_U12, R2358_U66);
  nand ginst2644 (R2358_U431, R2358_U136, R2358_U176);
  nand ginst2645 (R2358_U432, R2358_U11, R2358_U73);
  nand ginst2646 (R2358_U433, R2358_U312, R2358_U418);
  nand ginst2647 (R2358_U434, R2358_U418, R2358_U55);
  nand ginst2648 (R2358_U435, R2358_U140, R2358_U219, R2358_U410);
  nand ginst2649 (R2358_U436, R2358_U133, R2358_U327);
  nand ginst2650 (R2358_U437, R2358_U324, R2358_U436);
  nand ginst2651 (R2358_U438, R2358_U134, R2358_U328);
  not ginst2652 (R2358_U439, R2358_U62);
  not ginst2653 (R2358_U44, U2629);
  nand ginst2654 (R2358_U440, R2358_U164, U2352);
  nand ginst2655 (R2358_U441, R2358_U22, U2612);
  not ginst2656 (R2358_U442, R2358_U76);
  nand ginst2657 (R2358_U443, R2358_U442, U2641);
  nand ginst2658 (R2358_U444, R2358_U33, R2358_U76);
  nand ginst2659 (R2358_U445, R2358_U442, U2641);
  nand ginst2660 (R2358_U446, R2358_U33, R2358_U76);
  nand ginst2661 (R2358_U447, R2358_U445, R2358_U446);
  nand ginst2662 (R2358_U448, R2358_U166, U2352);
  nand ginst2663 (R2358_U449, R2358_U22, U2610);
  not ginst2664 (R2358_U45, U2630);
  nand ginst2665 (R2358_U450, R2358_U448, R2358_U449);
  nand ginst2666 (R2358_U451, R2358_U166, U2352);
  nand ginst2667 (R2358_U452, R2358_U22, U2610);
  nand ginst2668 (R2358_U453, R2358_U167, U2352);
  nand ginst2669 (R2358_U454, R2358_U22, U2609);
  not ginst2670 (R2358_U455, R2358_U77);
  nand ginst2671 (R2358_U456, R2358_U168, U2352);
  nand ginst2672 (R2358_U457, R2358_U22, U2667);
  nand ginst2673 (R2358_U458, R2358_U456, R2358_U457);
  nand ginst2674 (R2358_U459, R2358_U169, U2352);
  nand ginst2675 (R2358_U46, R2358_U78, U2630);
  nand ginst2676 (R2358_U460, R2358_U22, U2668);
  nand ginst2677 (R2358_U461, R2358_U459, R2358_U460);
  nand ginst2678 (R2358_U462, R2358_U168, U2352);
  nand ginst2679 (R2358_U463, R2358_U22, U2667);
  nand ginst2680 (R2358_U464, R2358_U169, U2352);
  nand ginst2681 (R2358_U465, R2358_U22, U2668);
  nand ginst2682 (R2358_U466, R2358_U170, U2352);
  nand ginst2683 (R2358_U467, R2358_U22, U2670);
  nand ginst2684 (R2358_U468, R2358_U466, R2358_U467);
  nand ginst2685 (R2358_U469, R2358_U171, U2352);
  not ginst2686 (R2358_U47, U2639);
  nand ginst2687 (R2358_U470, R2358_U22, U2671);
  nand ginst2688 (R2358_U471, R2358_U469, R2358_U470);
  nand ginst2689 (R2358_U472, R2358_U172, U2352);
  nand ginst2690 (R2358_U473, R2358_U22, U2672);
  nand ginst2691 (R2358_U474, R2358_U472, R2358_U473);
  nand ginst2692 (R2358_U475, R2358_U171, U2352);
  nand ginst2693 (R2358_U476, R2358_U22, U2671);
  nand ginst2694 (R2358_U477, R2358_U172, U2352);
  nand ginst2695 (R2358_U478, R2358_U22, U2672);
  nand ginst2696 (R2358_U479, R2358_U170, U2352);
  not ginst2697 (R2358_U48, U2640);
  nand ginst2698 (R2358_U480, R2358_U22, U2670);
  nand ginst2699 (R2358_U481, R2358_U173, U2352);
  nand ginst2700 (R2358_U482, R2358_U22, U2669);
  nand ginst2701 (R2358_U483, R2358_U173, U2352);
  nand ginst2702 (R2358_U484, R2358_U22, U2669);
  nand ginst2703 (R2358_U485, R2358_U483, R2358_U484);
  nand ginst2704 (R2358_U486, R2358_U174, U2352);
  nand ginst2705 (R2358_U487, R2358_U22, U2611);
  nand ginst2706 (R2358_U488, R2358_U174, U2352);
  nand ginst2707 (R2358_U489, R2358_U22, U2611);
  nand ginst2708 (R2358_U49, R2358_U490, U2642);
  nand ginst2709 (R2358_U490, R2358_U488, R2358_U489);
  nand ginst2710 (R2358_U491, R2358_U165, R2358_U175);
  nand ginst2711 (R2358_U492, R2358_U256, R2358_U447);
  nand ginst2712 (R2358_U493, R2358_U176, R2358_U381);
  nand ginst2713 (R2358_U494, R2358_U252, R2358_U84);
  nand ginst2714 (R2358_U495, R2358_U455, U2644);
  nand ginst2715 (R2358_U496, R2358_U24, R2358_U77);
  nand ginst2716 (R2358_U497, R2358_U495, R2358_U496);
  nand ginst2717 (R2358_U498, R2358_U34, R2358_U382);
  nand ginst2718 (R2358_U499, R2358_U260, R2358_U497);
  and ginst2719 (R2358_U5, R2358_U281, R2358_U282, R2358_U285, R2358_U293);
  not ginst2720 (R2358_U50, U2637);
  nand ginst2721 (R2358_U500, R2358_U177, R2358_U383);
  nand ginst2722 (R2358_U501, R2358_U258, R2358_U87);
  nand ginst2723 (R2358_U502, R2358_U178, R2358_U384);
  nand ginst2724 (R2358_U503, R2358_U241, R2358_U89);
  nand ginst2725 (R2358_U504, R2358_U179, U2352);
  nand ginst2726 (R2358_U505, R2358_U22, U2651);
  nand ginst2727 (R2358_U506, R2358_U179, U2352);
  nand ginst2728 (R2358_U507, R2358_U22, U2651);
  nand ginst2729 (R2358_U508, R2358_U506, R2358_U507);
  nand ginst2730 (R2358_U509, R2358_U181, U2352);
  nand ginst2731 (R2358_U51, R2358_U80, U2637);
  nand ginst2732 (R2358_U510, R2358_U22, U2613);
  nand ginst2733 (R2358_U511, R2358_U182, U2352);
  nand ginst2734 (R2358_U512, R2358_U22, U2614);
  nand ginst2735 (R2358_U513, R2358_U182, U2352);
  nand ginst2736 (R2358_U514, R2358_U22, U2614);
  nand ginst2737 (R2358_U515, R2358_U513, R2358_U514);
  nand ginst2738 (R2358_U516, R2358_U181, U2352);
  nand ginst2739 (R2358_U517, R2358_U22, U2613);
  nand ginst2740 (R2358_U518, R2358_U516, R2358_U517);
  nand ginst2741 (R2358_U519, R2358_U183, U2352);
  not ginst2742 (R2358_U52, U2638);
  nand ginst2743 (R2358_U520, R2358_U22, U2617);
  not ginst2744 (R2358_U521, R2358_U79);
  nand ginst2745 (R2358_U522, R2358_U184, U2352);
  nand ginst2746 (R2358_U523, R2358_U22, U2615);
  nand ginst2747 (R2358_U524, R2358_U185, U2352);
  nand ginst2748 (R2358_U525, R2358_U22, U2616);
  not ginst2749 (R2358_U526, R2358_U80);
  nand ginst2750 (R2358_U527, R2358_U186, U2352);
  nand ginst2751 (R2358_U528, R2358_U22, U2618);
  nand ginst2752 (R2358_U529, R2358_U184, U2352);
  nand ginst2753 (R2358_U53, R2358_U531, U2638);
  nand ginst2754 (R2358_U530, R2358_U22, U2615);
  nand ginst2755 (R2358_U531, R2358_U529, R2358_U530);
  nand ginst2756 (R2358_U532, R2358_U186, U2352);
  nand ginst2757 (R2358_U533, R2358_U22, U2618);
  not ginst2758 (R2358_U534, R2358_U81);
  nand ginst2759 (R2358_U535, R2358_U187, U2352);
  nand ginst2760 (R2358_U536, R2358_U22, U2664);
  nand ginst2761 (R2358_U537, R2358_U188, U2352);
  nand ginst2762 (R2358_U538, R2358_U22, U2665);
  nand ginst2763 (R2358_U539, R2358_U189, U2352);
  not ginst2764 (R2358_U54, U2636);
  nand ginst2765 (R2358_U540, R2358_U22, U2666);
  nand ginst2766 (R2358_U541, R2358_U190, U2352);
  nand ginst2767 (R2358_U542, R2358_U22, U2663);
  nand ginst2768 (R2358_U543, R2358_U191, U2352);
  nand ginst2769 (R2358_U544, R2358_U22, U2658);
  nand ginst2770 (R2358_U545, R2358_U192, U2352);
  nand ginst2771 (R2358_U546, R2358_U22, U2659);
  nand ginst2772 (R2358_U547, R2358_U193, U2352);
  nand ginst2773 (R2358_U548, R2358_U22, U2660);
  nand ginst2774 (R2358_U549, R2358_U194, U2352);
  nand ginst2775 (R2358_U55, R2358_U142, R2358_U9);
  nand ginst2776 (R2358_U550, R2358_U22, U2661);
  nand ginst2777 (R2358_U551, R2358_U195, U2352);
  nand ginst2778 (R2358_U552, R2358_U22, U2662);
  not ginst2779 (R2358_U553, R2358_U78);
  nand ginst2780 (R2358_U554, R2358_U196, U2352);
  nand ginst2781 (R2358_U555, R2358_U22, U2654);
  nand ginst2782 (R2358_U556, R2358_U197, U2352);
  nand ginst2783 (R2358_U557, R2358_U22, U2655);
  nand ginst2784 (R2358_U558, R2358_U198, U2352);
  nand ginst2785 (R2358_U559, R2358_U22, U2656);
  not ginst2786 (R2358_U56, U2631);
  nand ginst2787 (R2358_U560, R2358_U199, U2352);
  nand ginst2788 (R2358_U561, R2358_U22, U2657);
  nand ginst2789 (R2358_U562, R2358_U200, U2352);
  nand ginst2790 (R2358_U563, R2358_U22, U2652);
  nand ginst2791 (R2358_U564, R2358_U201, U2352);
  nand ginst2792 (R2358_U565, R2358_U22, U2653);
  nand ginst2793 (R2358_U566, R2358_U191, U2352);
  nand ginst2794 (R2358_U567, R2358_U22, U2658);
  nand ginst2795 (R2358_U568, R2358_U566, R2358_U567);
  nand ginst2796 (R2358_U569, R2358_U192, U2352);
  not ginst2797 (R2358_U57, U2632);
  nand ginst2798 (R2358_U570, R2358_U22, U2659);
  nand ginst2799 (R2358_U571, R2358_U569, R2358_U570);
  nand ginst2800 (R2358_U572, R2358_U193, U2352);
  nand ginst2801 (R2358_U573, R2358_U22, U2660);
  nand ginst2802 (R2358_U574, R2358_U572, R2358_U573);
  nand ginst2803 (R2358_U575, R2358_U194, U2352);
  nand ginst2804 (R2358_U576, R2358_U22, U2661);
  nand ginst2805 (R2358_U577, R2358_U575, R2358_U576);
  nand ginst2806 (R2358_U578, R2358_U200, U2352);
  nand ginst2807 (R2358_U579, R2358_U22, U2652);
  not ginst2808 (R2358_U58, U2633);
  nand ginst2809 (R2358_U580, R2358_U578, R2358_U579);
  nand ginst2810 (R2358_U581, R2358_U199, U2352);
  nand ginst2811 (R2358_U582, R2358_U22, U2657);
  nand ginst2812 (R2358_U583, R2358_U581, R2358_U582);
  nand ginst2813 (R2358_U584, R2358_U198, U2352);
  nand ginst2814 (R2358_U585, R2358_U22, U2656);
  nand ginst2815 (R2358_U586, R2358_U584, R2358_U585);
  nand ginst2816 (R2358_U587, R2358_U197, U2352);
  nand ginst2817 (R2358_U588, R2358_U22, U2655);
  nand ginst2818 (R2358_U589, R2358_U587, R2358_U588);
  nand ginst2819 (R2358_U59, R2358_U607, U2633);
  nand ginst2820 (R2358_U590, R2358_U196, U2352);
  nand ginst2821 (R2358_U591, R2358_U22, U2654);
  nand ginst2822 (R2358_U592, R2358_U590, R2358_U591);
  nand ginst2823 (R2358_U593, R2358_U201, U2352);
  nand ginst2824 (R2358_U594, R2358_U22, U2653);
  nand ginst2825 (R2358_U595, R2358_U593, R2358_U594);
  nand ginst2826 (R2358_U596, R2358_U190, U2352);
  nand ginst2827 (R2358_U597, R2358_U22, U2663);
  nand ginst2828 (R2358_U598, R2358_U596, R2358_U597);
  nand ginst2829 (R2358_U599, R2358_U189, U2352);
  and ginst2830 (R2358_U6, R2358_U325, R2358_U329);
  not ginst2831 (R2358_U60, U2634);
  nand ginst2832 (R2358_U600, R2358_U22, U2666);
  nand ginst2833 (R2358_U601, R2358_U599, R2358_U600);
  nand ginst2834 (R2358_U602, R2358_U187, U2352);
  nand ginst2835 (R2358_U603, R2358_U22, U2664);
  nand ginst2836 (R2358_U604, R2358_U602, R2358_U603);
  nand ginst2837 (R2358_U605, R2358_U188, U2352);
  nand ginst2838 (R2358_U606, R2358_U22, U2665);
  nand ginst2839 (R2358_U607, R2358_U605, R2358_U606);
  nand ginst2840 (R2358_U608, R2358_U180, R2358_U202);
  nand ginst2841 (R2358_U609, R2358_U330, R2358_U508);
  nand ginst2842 (R2358_U61, R2358_U601, U2634);
  nand ginst2843 (R2358_U610, R2358_U203, R2358_U385);
  nand ginst2844 (R2358_U611, R2358_U333, R2358_U92);
  nand ginst2845 (R2358_U612, R2358_U204, R2358_U386);
  nand ginst2846 (R2358_U613, R2358_U339, R2358_U94);
  nand ginst2847 (R2358_U614, R2358_U205, R2358_U387);
  nand ginst2848 (R2358_U615, R2358_U341, R2358_U96);
  nand ginst2849 (R2358_U616, R2358_U221, R2358_U388);
  nand ginst2850 (R2358_U617, R2358_U206, R2358_U98);
  nand ginst2851 (R2358_U618, R2358_U207, R2358_U389);
  nand ginst2852 (R2358_U619, R2358_U100, R2358_U343);
  nand ginst2853 (R2358_U62, R2358_U320, R2358_U438);
  nand ginst2854 (R2358_U620, R2358_U208, R2358_U390);
  nand ginst2855 (R2358_U621, R2358_U102, R2358_U331);
  nand ginst2856 (R2358_U622, R2358_U209, R2358_U391);
  nand ginst2857 (R2358_U623, R2358_U104, R2358_U348);
  nand ginst2858 (R2358_U624, R2358_U210, R2358_U392);
  nand ginst2859 (R2358_U625, R2358_U106, R2358_U346);
  nand ginst2860 (R2358_U626, R2358_U220, R2358_U393);
  nand ginst2861 (R2358_U627, R2358_U108, R2358_U211);
  nand ginst2862 (R2358_U628, R2358_U553, U2630);
  nand ginst2863 (R2358_U629, R2358_U45, R2358_U78);
  nand ginst2864 (R2358_U63, R2358_U280, R2358_U291);
  nand ginst2865 (R2358_U630, R2358_U628, R2358_U629);
  nand ginst2866 (R2358_U631, R2358_U394, R2358_U68);
  nand ginst2867 (R2358_U632, R2358_U318, R2358_U630);
  nand ginst2868 (R2358_U633, R2358_U212, R2358_U395);
  nand ginst2869 (R2358_U634, R2358_U111, R2358_U269);
  nand ginst2870 (R2358_U635, R2358_U213, R2358_U396);
  nand ginst2871 (R2358_U636, R2358_U113, R2358_U315);
  nand ginst2872 (R2358_U637, R2358_U214, R2358_U397);
  nand ginst2873 (R2358_U638, R2358_U115, R2358_U357);
  nand ginst2874 (R2358_U639, R2358_U215, R2358_U398);
  nand ginst2875 (R2358_U64, R2358_U233, R2358_U270);
  nand ginst2876 (R2358_U640, R2358_U117, R2358_U355);
  nand ginst2877 (R2358_U641, R2358_U521, U2636);
  nand ginst2878 (R2358_U642, R2358_U54, R2358_U79);
  nand ginst2879 (R2358_U643, R2358_U641, R2358_U642);
  nand ginst2880 (R2358_U644, R2358_U399, R2358_U72);
  nand ginst2881 (R2358_U645, R2358_U365, R2358_U643);
  nand ginst2882 (R2358_U646, R2358_U526, U2637);
  nand ginst2883 (R2358_U647, R2358_U50, R2358_U80);
  nand ginst2884 (R2358_U648, R2358_U646, R2358_U647);
  nand ginst2885 (R2358_U649, R2358_U216, R2358_U400);
  nand ginst2886 (R2358_U65, R2358_U229, R2358_U64);
  nand ginst2887 (R2358_U650, R2358_U362, R2358_U648);
  nand ginst2888 (R2358_U651, R2358_U217, R2358_U401);
  nand ginst2889 (R2358_U652, R2358_U121, R2358_U308);
  nand ginst2890 (R2358_U653, R2358_U218, U2352);
  nand ginst2891 (R2358_U654, R2358_U22, R2358_U380);
  nand ginst2892 (R2358_U66, R2358_U316, R2358_U417);
  nand ginst2893 (R2358_U67, R2358_U146, R2358_U219, R2358_U410);
  nand ginst2894 (R2358_U68, R2358_U416, R2358_U418);
  nand ginst2895 (R2358_U69, R2358_U295, R2358_U407, R2358_U408);
  and ginst2896 (R2358_U7, R2358_U141, R2358_U324, R2358_U6);
  nand ginst2897 (R2358_U70, R2358_U313, R2358_U67);
  not ginst2898 (R2358_U71, U2635);
  nand ginst2899 (R2358_U72, R2358_U364, R2358_U51);
  nand ginst2900 (R2358_U73, R2358_U305, R2358_U414);
  nand ginst2901 (R2358_U74, R2358_U413, R2358_U423);
  nand ginst2902 (R2358_U75, R2358_U301, R2358_U74);
  nand ginst2903 (R2358_U76, R2358_U440, R2358_U441);
  nand ginst2904 (R2358_U77, R2358_U453, R2358_U454);
  nand ginst2905 (R2358_U78, R2358_U551, R2358_U552);
  nand ginst2906 (R2358_U79, R2358_U519, R2358_U520);
  and ginst2907 (R2358_U8, R2358_U135, R2358_U5);
  nand ginst2908 (R2358_U80, R2358_U524, R2358_U525);
  nand ginst2909 (R2358_U81, R2358_U532, R2358_U533);
  nand ginst2910 (R2358_U82, R2358_U653, R2358_U654);
  nand ginst2911 (R2358_U83, R2358_U491, R2358_U492);
  and ginst2912 (R2358_U84, R2358_U253, R2358_U49);
  nand ginst2913 (R2358_U85, R2358_U493, R2358_U494);
  nand ginst2914 (R2358_U86, R2358_U498, R2358_U499);
  and ginst2915 (R2358_U87, R2358_U243, R2358_U246);
  nand ginst2916 (R2358_U88, R2358_U500, R2358_U501);
  and ginst2917 (R2358_U89, R2358_U244, R2358_U247);
  and ginst2918 (R2358_U9, R2358_U294, R2358_U296);
  nand ginst2919 (R2358_U90, R2358_U502, R2358_U503);
  nand ginst2920 (R2358_U91, R2358_U608, R2358_U609);
  and ginst2921 (R2358_U92, R2358_U277, R2358_U278);
  nand ginst2922 (R2358_U93, R2358_U610, R2358_U611);
  and ginst2923 (R2358_U94, R2358_U279, R2358_U280);
  nand ginst2924 (R2358_U95, R2358_U612, R2358_U613);
  and ginst2925 (R2358_U96, R2358_U281, R2358_U288);
  nand ginst2926 (R2358_U97, R2358_U614, R2358_U615);
  and ginst2927 (R2358_U98, R2358_U282, R2358_U289);
  nand ginst2928 (R2358_U99, R2358_U616, R2358_U617);
  not ginst2929 (R584_U6, U2676);
  not ginst2930 (R584_U7, U2677);
  not ginst2931 (R584_U8, U2674);
  not ginst2932 (R584_U9, U2675);
  not ginst2933 (SUB_357_U10, U3214);
  not ginst2934 (SUB_357_U11, U3217);
  not ginst2935 (SUB_357_U12, U3216);
  not ginst2936 (SUB_357_U13, U3218);
  not ginst2937 (SUB_357_U6, U3220);
  not ginst2938 (SUB_357_U7, U3215);
  not ginst2939 (SUB_357_U8, U3221);
  not ginst2940 (SUB_357_U9, U3219);
  not ginst2941 (SUB_450_U10, INSTQUEUEWR_ADDR_REG_1__SCAN_IN);
  not ginst2942 (SUB_450_U11, INSTQUEUERD_ADDR_REG_2__SCAN_IN);
  not ginst2943 (SUB_450_U12, INSTQUEUEWR_ADDR_REG_2__SCAN_IN);
  not ginst2944 (SUB_450_U13, INSTQUEUERD_ADDR_REG_3__SCAN_IN);
  not ginst2945 (SUB_450_U14, INSTQUEUEWR_ADDR_REG_3__SCAN_IN);
  not ginst2946 (SUB_450_U15, INSTQUEUEWR_ADDR_REG_4__SCAN_IN);
  nand ginst2947 (SUB_450_U16, SUB_450_U40, SUB_450_U41);
  not ginst2948 (SUB_450_U17, INSTQUEUERD_ADDR_REG_4__SCAN_IN);
  not ginst2949 (SUB_450_U18, INSTQUEUEWR_ADDR_REG_0__SCAN_IN);
  nand ginst2950 (SUB_450_U19, SUB_450_U50, SUB_450_U51);
  nand ginst2951 (SUB_450_U20, SUB_450_U55, SUB_450_U56);
  nand ginst2952 (SUB_450_U21, SUB_450_U60, SUB_450_U61);
  nand ginst2953 (SUB_450_U22, SUB_450_U65, SUB_450_U66);
  nand ginst2954 (SUB_450_U23, SUB_450_U47, SUB_450_U48);
  nand ginst2955 (SUB_450_U24, SUB_450_U52, SUB_450_U53);
  nand ginst2956 (SUB_450_U25, SUB_450_U57, SUB_450_U58);
  nand ginst2957 (SUB_450_U26, SUB_450_U62, SUB_450_U63);
  nand ginst2958 (SUB_450_U27, SUB_450_U36, SUB_450_U37);
  nand ginst2959 (SUB_450_U28, SUB_450_U32, SUB_450_U33);
  not ginst2960 (SUB_450_U29, INSTQUEUERD_ADDR_REG_1__SCAN_IN);
  not ginst2961 (SUB_450_U30, SUB_450_U9);
  nand ginst2962 (SUB_450_U31, SUB_450_U10, SUB_450_U30);
  nand ginst2963 (SUB_450_U32, SUB_450_U29, SUB_450_U31);
  nand ginst2964 (SUB_450_U33, INSTQUEUEWR_ADDR_REG_1__SCAN_IN, SUB_450_U9);
  not ginst2965 (SUB_450_U34, SUB_450_U28);
  nand ginst2966 (SUB_450_U35, INSTQUEUERD_ADDR_REG_2__SCAN_IN, SUB_450_U12);
  nand ginst2967 (SUB_450_U36, SUB_450_U28, SUB_450_U35);
  nand ginst2968 (SUB_450_U37, INSTQUEUEWR_ADDR_REG_2__SCAN_IN, SUB_450_U11);
  not ginst2969 (SUB_450_U38, SUB_450_U27);
  nand ginst2970 (SUB_450_U39, INSTQUEUERD_ADDR_REG_3__SCAN_IN, SUB_450_U14);
  nand ginst2971 (SUB_450_U40, SUB_450_U27, SUB_450_U39);
  nand ginst2972 (SUB_450_U41, INSTQUEUEWR_ADDR_REG_3__SCAN_IN, SUB_450_U13);
  not ginst2973 (SUB_450_U42, SUB_450_U16);
  nand ginst2974 (SUB_450_U43, INSTQUEUEWR_ADDR_REG_4__SCAN_IN, SUB_450_U17);
  nand ginst2975 (SUB_450_U44, SUB_450_U42, SUB_450_U43);
  nand ginst2976 (SUB_450_U45, INSTQUEUERD_ADDR_REG_4__SCAN_IN, SUB_450_U15);
  nand ginst2977 (SUB_450_U46, INSTQUEUEWR_ADDR_REG_0__SCAN_IN, SUB_450_U8);
  nand ginst2978 (SUB_450_U47, INSTQUEUERD_ADDR_REG_4__SCAN_IN, SUB_450_U15);
  nand ginst2979 (SUB_450_U48, INSTQUEUEWR_ADDR_REG_4__SCAN_IN, SUB_450_U17);
  not ginst2980 (SUB_450_U49, SUB_450_U23);
  nand ginst2981 (SUB_450_U50, SUB_450_U42, SUB_450_U49);
  nand ginst2982 (SUB_450_U51, SUB_450_U16, SUB_450_U23);
  nand ginst2983 (SUB_450_U52, INSTQUEUERD_ADDR_REG_3__SCAN_IN, SUB_450_U14);
  nand ginst2984 (SUB_450_U53, INSTQUEUEWR_ADDR_REG_3__SCAN_IN, SUB_450_U13);
  not ginst2985 (SUB_450_U54, SUB_450_U24);
  nand ginst2986 (SUB_450_U55, SUB_450_U38, SUB_450_U54);
  nand ginst2987 (SUB_450_U56, SUB_450_U24, SUB_450_U27);
  nand ginst2988 (SUB_450_U57, INSTQUEUERD_ADDR_REG_2__SCAN_IN, SUB_450_U12);
  nand ginst2989 (SUB_450_U58, INSTQUEUEWR_ADDR_REG_2__SCAN_IN, SUB_450_U11);
  not ginst2990 (SUB_450_U59, SUB_450_U25);
  nand ginst2991 (SUB_450_U6, SUB_450_U44, SUB_450_U45);
  nand ginst2992 (SUB_450_U60, SUB_450_U34, SUB_450_U59);
  nand ginst2993 (SUB_450_U61, SUB_450_U25, SUB_450_U28);
  nand ginst2994 (SUB_450_U62, INSTQUEUERD_ADDR_REG_1__SCAN_IN, SUB_450_U10);
  nand ginst2995 (SUB_450_U63, INSTQUEUEWR_ADDR_REG_1__SCAN_IN, SUB_450_U29);
  not ginst2996 (SUB_450_U64, SUB_450_U26);
  nand ginst2997 (SUB_450_U65, SUB_450_U30, SUB_450_U64);
  nand ginst2998 (SUB_450_U66, SUB_450_U26, SUB_450_U9);
  nand ginst2999 (SUB_450_U7, SUB_450_U46, SUB_450_U9);
  not ginst3000 (SUB_450_U8, INSTQUEUERD_ADDR_REG_0__SCAN_IN);
  nand ginst3001 (SUB_450_U9, INSTQUEUERD_ADDR_REG_0__SCAN_IN, SUB_450_U18);
  nand ginst3002 (SUB_580_U10, INSTADDRPOINTER_REG_0__SCAN_IN, SUB_580_U7);
  nand ginst3003 (SUB_580_U6, SUB_580_U10, SUB_580_U9);
  not ginst3004 (SUB_580_U7, INSTADDRPOINTER_REG_1__SCAN_IN);
  not ginst3005 (SUB_580_U8, INSTADDRPOINTER_REG_0__SCAN_IN);
  nand ginst3006 (SUB_580_U9, INSTADDRPOINTER_REG_1__SCAN_IN, SUB_580_U8);
  nor ginst3007 (U2352, STATEBS16_REG_SCAN_IN, STATE2_REG_2__SCAN_IN);
  and ginst3008 (U2353, STATE2_REG_2__SCAN_IN, U4219);
  and ginst3009 (U2354, U4253, U4465);
  and ginst3010 (U2355, U2450, U3221);
  and ginst3011 (U2356, R2238_U6, U4180);
  and ginst3012 (U2357, R2167_U17, U3853, U5947);
  and ginst3013 (U2358, U2388, U4212);
  and ginst3014 (U2359, STATE2_REG_2__SCAN_IN, U3418);
  and ginst3015 (U2360, STATE2_REG_2__SCAN_IN, U3401);
  and ginst3016 (U2361, STATE2_REG_3__SCAN_IN, U4212);
  and ginst3017 (U2362, U2359, U4196);
  and ginst3018 (U2363, U2359, U4198);
  and ginst3019 (U2364, U3403, U3852);
  and ginst3020 (U2365, U3403, U4249);
  and ginst3021 (U2366, STATE2_REG_1__SCAN_IN, U3417, U3418);
  and ginst3022 (U2367, STATE2_REG_1__SCAN_IN, R2337_U58, U3418);
  and ginst3023 (U2368, STATE2_REG_0__SCAN_IN, U4223);
  and ginst3024 (U2369, U2362, U4485);
  and ginst3025 (U2370, U3250, U3401);
  and ginst3026 (U2371, U4210, U4437);
  and ginst3027 (U2372, STATE2_REG_0__SCAN_IN, U3403);
  and ginst3028 (U2373, STATE2_REG_3__SCAN_IN, U3418);
  and ginst3029 (U2374, U2360, U4202);
  and ginst3030 (U2375, U2360, U4204);
  and ginst3031 (U2376, U3403, U5786);
  and ginst3032 (U2377, U3401, U3750);
  and ginst3033 (U2378, U2360, U5557);
  and ginst3034 (U2379, U2363, U3267);
  and ginst3035 (U2380, U2360, U7596);
  and ginst3036 (U2381, U2357, U3258);
  and ginst3037 (U2382, U2357, U4465);
  and ginst3038 (U2383, U3378, U4210);
  and ginst3039 (U2384, STATE2_REG_0__SCAN_IN, U3404);
  and ginst3040 (U2385, U3281, U3404);
  and ginst3041 (U2386, U3410, U4211);
  and ginst3042 (U2387, U3872, U4211);
  and ginst3043 (U2388, STATEBS16_REG_SCAN_IN, U4197);
  and ginst3044 (U2389, U2452, U7482);
  and ginst3045 (U2390, DATAI_0_, U4212);
  and ginst3046 (U2391, DATAI_1_, U4212);
  and ginst3047 (U2392, DATAI_2_, U4212);
  and ginst3048 (U2393, DATAI_3_, U4212);
  and ginst3049 (U2394, DATAI_4_, U4212);
  and ginst3050 (U2395, DATAI_5_, U4212);
  and ginst3051 (U2396, DATAI_6_, U4212);
  and ginst3052 (U2397, DATAI_7_, U4212);
  and ginst3053 (U2398, DATAI_24_, U2358);
  and ginst3054 (U2399, DATAI_16_, U2358);
  and ginst3055 (U2400, DATAI_25_, U2358);
  and ginst3056 (U2401, DATAI_17_, U2358);
  and ginst3057 (U2402, DATAI_26_, U2358);
  and ginst3058 (U2403, DATAI_18_, U2358);
  and ginst3059 (U2404, DATAI_27_, U2358);
  and ginst3060 (U2405, DATAI_19_, U2358);
  and ginst3061 (U2406, DATAI_28_, U2358);
  and ginst3062 (U2407, DATAI_20_, U2358);
  and ginst3063 (U2408, DATAI_29_, U2358);
  and ginst3064 (U2409, DATAI_21_, U2358);
  and ginst3065 (U2410, DATAI_30_, U2358);
  and ginst3066 (U2411, DATAI_22_, U2358);
  and ginst3067 (U2412, DATAI_31_, U2358);
  and ginst3068 (U2413, DATAI_23_, U2358);
  and ginst3069 (U2414, U2361, U3258);
  and ginst3070 (U2415, U2361, U3378);
  and ginst3071 (U2416, U2361, U3264);
  and ginst3072 (U2417, U2361, U3271);
  and ginst3073 (U2418, U2361, U3270);
  and ginst3074 (U2419, U2361, U3265);
  and ginst3075 (U2420, U2361, U4161);
  and ginst3076 (U2421, U2361, U4159);
  and ginst3077 (U2422, U4211, U5449);
  and ginst3078 (U2423, U4211, U4219);
  and ginst3079 (U2424, U2384, U3271);
  and ginst3080 (U2425, U2368, U2448);
  and ginst3081 (U2426, U3418, U3877);
  nor ginst3082 (U2427, STATE2_REG_3__SCAN_IN, STATE2_REG_1__SCAN_IN);
  and ginst3083 (U2428, STATE2_REG_2__SCAN_IN, STATE2_REG_1__SCAN_IN);
  and ginst3084 (U2429, U3418, U6354);
  and ginst3085 (U2430, STATE2_REG_1__SCAN_IN, U3374);
  and ginst3086 (U2431, U4187, U7482);
  and ginst3087 (U2432, U3347, U3442);
  and ginst3088 (U2433, U3442, U4528);
  and ginst3089 (U2434, U3347, U7684);
  and ginst3090 (U2435, U4528, U7684);
  and ginst3091 (U2436, U3222, U3288);
  and ginst3092 (U2437, U3288, U4531);
  and ginst3093 (U2438, R2182_U25, R2182_U42);
  and ginst3094 (U2439, R2182_U42, U3303);
  and ginst3095 (U2440, R2182_U25, U3304);
  nor ginst3096 (U2441, R2182_U25, R2182_U42);
  and ginst3097 (U2442, R2182_U33, R2182_U34);
  and ginst3098 (U2443, R2182_U33, U3305);
  and ginst3099 (U2444, R2182_U34, U3306);
  nor ginst3100 (U2445, R2182_U33, R2182_U34);
  and ginst3101 (U2446, STATE2_REG_1__SCAN_IN, U3458);
  and ginst3102 (U2447, U2452, U3565);
  and ginst3103 (U2448, R2167_U17, U3271);
  and ginst3104 (U2449, U3258, U4482);
  and ginst3105 (U2450, STATE2_REG_0__SCAN_IN, U4388);
  and ginst3106 (U2451, STATE2_REG_0__SCAN_IN, U4239);
  and ginst3107 (U2452, U3264, U3378, U4161, U4388);
  and ginst3108 (U2453, INSTQUEUERD_ADDR_REG_3__SCAN_IN, INSTQUEUERD_ADDR_REG_2__SCAN_IN, INSTQUEUERD_ADDR_REG_1__SCAN_IN, INSTQUEUERD_ADDR_REG_0__SCAN_IN);
  and ginst3109 (U2454, INSTQUEUERD_ADDR_REG_1__SCAN_IN, U3253);
  and ginst3110 (U2455, INSTQUEUERD_ADDR_REG_3__SCAN_IN, INSTQUEUERD_ADDR_REG_2__SCAN_IN, INSTQUEUERD_ADDR_REG_1__SCAN_IN, U3253);
  and ginst3111 (U2456, INSTQUEUERD_ADDR_REG_0__SCAN_IN, U3252);
  and ginst3112 (U2457, INSTQUEUERD_ADDR_REG_3__SCAN_IN, INSTQUEUERD_ADDR_REG_2__SCAN_IN, INSTQUEUERD_ADDR_REG_0__SCAN_IN, U3252);
  and ginst3113 (U2458, U3495, U4366);
  and ginst3114 (U2459, INSTQUEUERD_ADDR_REG_3__SCAN_IN, INSTQUEUERD_ADDR_REG_1__SCAN_IN, INSTQUEUERD_ADDR_REG_0__SCAN_IN, U3251);
  and ginst3115 (U2460, INSTQUEUERD_ADDR_REG_1__SCAN_IN, U3251, U3253);
  and ginst3116 (U2461, U3493, U3494);
  and ginst3117 (U2462, INSTQUEUERD_ADDR_REG_0__SCAN_IN, U3251, U3252);
  and ginst3118 (U2463, U3491, U3492);
  and ginst3119 (U2464, INSTQUEUERD_ADDR_REG_3__SCAN_IN, U4368);
  and ginst3120 (U2465, U3489, U3490);
  and ginst3121 (U2466, U3487, U3488);
  and ginst3122 (U2467, INSTQUEUERD_ADDR_REG_2__SCAN_IN, U3257, U4366);
  and ginst3123 (U2468, U3485, U3486);
  nor ginst3124 (U2469, INSTQUEUERD_ADDR_REG_3__SCAN_IN, INSTQUEUERD_ADDR_REG_2__SCAN_IN);
  and ginst3125 (U2470, INSTQUEUERD_ADDR_REG_1__SCAN_IN, U2469, U3253);
  and ginst3126 (U2471, INSTQUEUERD_ADDR_REG_0__SCAN_IN, U2469, U3252);
  and ginst3127 (U2472, U3257, U4368);
  and ginst3128 (U2473, U3393, U7667, U7668);
  and ginst3129 (U2474, R2144_U49, U3299);
  and ginst3130 (U2475, U3345, U3441);
  and ginst3131 (U2476, R2144_U49, R2144_U8);
  and ginst3132 (U2477, U2476, U4516);
  and ginst3133 (U2478, INSTQUEUEWR_ADDR_REG_3__SCAN_IN, INSTQUEUEWR_ADDR_REG_2__SCAN_IN);
  and ginst3134 (U2479, INSTQUEUEWR_ADDR_REG_2__SCAN_IN, U3290);
  and ginst3135 (U2480, U3302, U4536);
  and ginst3136 (U2481, U2476, U4512);
  and ginst3137 (U2482, U3314, U4594);
  and ginst3138 (U2483, U2476, U4513);
  and ginst3139 (U2484, U3321, U4653);
  and ginst3140 (U2485, R2144_U43, U4514);
  nor ginst3141 (U2486, R2144_U43, R2144_U50);
  and ginst3142 (U2487, U2476, U2486);
  nor ginst3143 (U2488, INSTQUEUEWR_ADDR_REG_1__SCAN_IN, INSTQUEUEWR_ADDR_REG_0__SCAN_IN);
  and ginst3144 (U2489, U3325, U4710);
  and ginst3145 (U2490, U3345, U7681);
  and ginst3146 (U2491, U4516, U4517);
  and ginst3147 (U2492, U3330, U4768);
  and ginst3148 (U2493, U4512, U4517);
  and ginst3149 (U2494, U3334, U4825);
  and ginst3150 (U2495, U4513, U4517);
  and ginst3151 (U2496, U3337, U4883);
  and ginst3152 (U2497, U2486, U4517);
  and ginst3153 (U2498, U3341, U4940);
  and ginst3154 (U2499, U3441, U4519);
  and ginst3155 (U2500, U3344, U3346);
  and ginst3156 (U2501, U2474, U4512);
  and ginst3157 (U2502, U3351, U5053);
  and ginst3158 (U2503, U2474, U4513);
  and ginst3159 (U2504, U3354, U5111);
  and ginst3160 (U2505, U2474, U2486);
  and ginst3161 (U2506, U3358, U5168);
  and ginst3162 (U2507, U4519, U7681);
  nor ginst3163 (U2508, R2144_U49, R2144_U8);
  and ginst3164 (U2509, U2508, U4516);
  nor ginst3165 (U2510, INSTQUEUEWR_ADDR_REG_3__SCAN_IN, INSTQUEUEWR_ADDR_REG_2__SCAN_IN);
  and ginst3166 (U2511, U3361, U5226);
  and ginst3167 (U2512, U2508, U4512);
  and ginst3168 (U2513, U3365, U5283);
  and ginst3169 (U2514, U2508, U4513);
  and ginst3170 (U2515, U3368, U5341);
  and ginst3171 (U2516, U2486, U2508);
  and ginst3172 (U2517, U3372, U5398);
  and ginst3173 (U2518, U5456, U7687, U7688);
  and ginst3174 (U2519, U3732, U5487);
  and ginst3175 (U2520, U3433, U4207);
  and ginst3176 (U2521, INSTQUEUERD_ADDR_REG_0__SCAN_IN, U3389);
  and ginst3177 (U2522, U5471, U5499);
  and ginst3178 (U2523, U2521, U2522);
  and ginst3179 (U2524, U3253, U3389);
  and ginst3180 (U2525, U2522, U2524);
  and ginst3181 (U2526, INSTQUEUERD_ADDR_REG_0__SCAN_IN, U5507);
  and ginst3182 (U2527, U2522, U2526);
  and ginst3183 (U2528, U3253, U5507);
  and ginst3184 (U2529, U2522, U2528);
  and ginst3185 (U2530, U3388, U5471);
  and ginst3186 (U2531, U2521, U2530);
  and ginst3187 (U2532, U2524, U2530);
  and ginst3188 (U2533, U2526, U2530);
  and ginst3189 (U2534, U2528, U2530);
  and ginst3190 (U2535, U3425, U5499);
  and ginst3191 (U2536, U2521, U2535);
  and ginst3192 (U2537, U2524, U2535);
  and ginst3193 (U2538, U2526, U2535);
  and ginst3194 (U2539, U2528, U2535);
  and ginst3195 (U2540, U3388, U3425);
  and ginst3196 (U2541, U2521, U2540);
  and ginst3197 (U2542, U2524, U2540);
  and ginst3198 (U2543, U2526, U2540);
  and ginst3199 (U2544, U2528, U2540);
  and ginst3200 (U2545, U5468, U7708);
  and ginst3201 (U2546, U2454, U2545);
  and ginst3202 (U2547, U2545, U3486);
  and ginst3203 (U2548, U2545, U4366);
  and ginst3204 (U2549, U2456, U2545);
  and ginst3205 (U2550, U3443, U5468);
  and ginst3206 (U2551, U2454, U2550);
  and ginst3207 (U2552, U2550, U3486);
  and ginst3208 (U2553, U2550, U4366);
  and ginst3209 (U2554, U2456, U2550);
  and ginst3210 (U2555, U3429, U7708);
  and ginst3211 (U2556, U2454, U2555);
  and ginst3212 (U2557, U2555, U3486);
  and ginst3213 (U2558, U2555, U4366);
  and ginst3214 (U2559, U2456, U2555);
  and ginst3215 (U2560, U3429, U3443);
  and ginst3216 (U2561, U2454, U2560);
  and ginst3217 (U2562, U2560, U3486);
  and ginst3218 (U2563, U2560, U4366);
  and ginst3219 (U2564, U2456, U2560);
  and ginst3220 (U2565, U4367, U7053);
  and ginst3221 (U2566, U2460, U7053);
  and ginst3222 (U2567, U2462, U7053);
  and ginst3223 (U2568, U4368, U7053);
  and ginst3224 (U2569, INSTQUEUERD_ADDR_REG_2__SCAN_IN, U7053);
  and ginst3225 (U2570, U2569, U3486);
  and ginst3226 (U2571, U2454, U2569);
  and ginst3227 (U2572, U2456, U2569);
  and ginst3228 (U2573, U2569, U4366);
  and ginst3229 (U2574, U3432, U4367);
  and ginst3230 (U2575, U2460, U3432);
  and ginst3231 (U2576, U2462, U3432);
  and ginst3232 (U2577, U3432, U4368);
  and ginst3233 (U2578, INSTQUEUERD_ADDR_REG_2__SCAN_IN, U3432);
  and ginst3234 (U2579, U2578, U3486);
  and ginst3235 (U2580, U2454, U2578);
  and ginst3236 (U2581, U2456, U2578);
  and ginst3237 (U2582, U2578, U4366);
  and ginst3238 (U2583, U4172, U7778);
  and ginst3239 (U2584, U2524, U2583);
  and ginst3240 (U2585, U2521, U2583);
  and ginst3241 (U2586, U2528, U2583);
  and ginst3242 (U2587, U2526, U2583);
  and ginst3243 (U2588, U3439, U7778);
  and ginst3244 (U2589, U2524, U2588);
  and ginst3245 (U2590, U2521, U2588);
  and ginst3246 (U2591, U2528, U2588);
  and ginst3247 (U2592, U2526, U2588);
  and ginst3248 (U2593, U3444, U4172);
  and ginst3249 (U2594, U2524, U2593);
  and ginst3250 (U2595, U2521, U2593);
  and ginst3251 (U2596, U2528, U2593);
  and ginst3252 (U2597, U2526, U2593);
  and ginst3253 (U2598, U3439, U3444);
  and ginst3254 (U2599, U2524, U2598);
  and ginst3255 (U2600, U2521, U2598);
  and ginst3256 (U2601, U2528, U2598);
  and ginst3257 (U2602, U2526, U2598);
  and ginst3258 (U2603, STATE2_REG_0__SCAN_IN, U3376);
  and ginst3259 (U2604, EBX_REG_31__SCAN_IN, U2379);
  and ginst3260 (U2605, U2607, U3518, U3519, U3520, U3521);
  and ginst3261 (U2606, U3414, U7492);
  and ginst3262 (U2607, U7659, U7660);
  and ginst3263 (U2608, U7774, U7775);
  nand ginst3264 (U2609, U3993, U6744);
  nand ginst3265 (U2610, U3992, U6741);
  nand ginst3266 (U2611, U3991, U6738);
  nand ginst3267 (U2612, U3990, U6735);
  nand ginst3268 (U2613, U4014, U6844);
  nand ginst3269 (U2614, U6841, U6842, U6843);
  nand ginst3270 (U2615, U6838, U6839, U6840);
  nand ginst3271 (U2616, U6835, U6836, U6837);
  nand ginst3272 (U2617, U6832, U6833, U6834);
  nand ginst3273 (U2618, U6829, U6830, U6831);
  and ginst3274 (U2620, R2144_U145, U6734);
  and ginst3275 (U2621, R2144_U145, U6734);
  and ginst3276 (U2622, R2144_U145, U6734);
  and ginst3277 (U2623, R2144_U145, U6734);
  and ginst3278 (U2624, R2144_U145, U6734);
  and ginst3279 (U2625, R2144_U145, U6734);
  and ginst3280 (U2626, R2144_U145, U6734);
  and ginst3281 (U2627, R2144_U145, U6734);
  and ginst3282 (U2628, R2144_U145, U6734);
  and ginst3283 (U2629, R2144_U145, U6734);
  and ginst3284 (U2630, R2144_U145, U6734);
  and ginst3285 (U2631, R2144_U145, U6734);
  and ginst3286 (U2632, R2144_U145, U6734);
  and ginst3287 (U2633, R2144_U145, U6734);
  and ginst3288 (U2634, R2144_U11, U6734);
  and ginst3289 (U2635, R2144_U37, U6734);
  and ginst3290 (U2636, R2144_U38, U6734);
  and ginst3291 (U2637, R2144_U39, U6734);
  and ginst3292 (U2638, R2144_U40, U6734);
  and ginst3293 (U2639, R2144_U41, U6734);
  and ginst3294 (U2640, R2144_U42, U6734);
  and ginst3295 (U2641, R2144_U30, U6734);
  and ginst3296 (U2642, R2144_U80, U6734);
  and ginst3297 (U2643, R2144_U10, U6734);
  and ginst3298 (U2644, R2144_U9, U6734);
  and ginst3299 (U2645, R2144_U45, U6734);
  and ginst3300 (U2646, R2144_U47, U6734);
  and ginst3301 (U2647, R2144_U8, U6734);
  nand ginst3302 (U2648, U3427, U6857);
  and ginst3303 (U2649, R2144_U50, U6734);
  and ginst3304 (U2650, STATE2_REG_2__SCAN_IN, U6858);
  nand ginst3305 (U2651, U6756, U6757, U6758);
  nand ginst3306 (U2652, U3997, U6759);
  nand ginst3307 (U2653, U3999, U6768);
  nand ginst3308 (U2654, U4000, U6772);
  nand ginst3309 (U2655, U4001, U6776);
  nand ginst3310 (U2656, U4002, U6780);
  nand ginst3311 (U2657, U4003, U6784);
  nand ginst3312 (U2658, U4004, U6788);
  nand ginst3313 (U2659, U4005, U6792);
  nand ginst3314 (U2660, U4006, U6796);
  nand ginst3315 (U2661, U4007, U6800);
  nand ginst3316 (U2662, U4008, U6804);
  nand ginst3317 (U2663, U4010, U6813);
  nand ginst3318 (U2664, U4011, U6817);
  nand ginst3319 (U2665, U4012, U6821);
  nand ginst3320 (U2666, U4013, U6825);
  nand ginst3321 (U2667, U3994, U6747);
  nand ginst3322 (U2668, U3996, U6751, U6754, U6755);
  nand ginst3323 (U2669, U3998, U6763, U6766, U6767);
  nand ginst3324 (U2670, U4009, U6808, U6811, U6812);
  nand ginst3325 (U2671, U4015, U6847, U6850, U6851);
  nand ginst3326 (U2672, U6852, U6853, U6854, U6855, U6856);
  nand ginst3327 (U2673, U7445, U7446);
  nand ginst3328 (U2674, U7447, U7448);
  nand ginst3329 (U2675, U4156, U7451);
  nand ginst3330 (U2676, U4157, U7454);
  nand ginst3331 (U2677, U7455, U7781, U7782);
  nand ginst3332 (U2678, U3271, U7444);
  nand ginst3333 (U2679, U7392, U7393);
  nand ginst3334 (U2680, U7394, U7395);
  nand ginst3335 (U2681, U7398, U7399);
  nand ginst3336 (U2682, U7400, U7401);
  nand ginst3337 (U2683, U7402, U7403);
  nand ginst3338 (U2684, U7404, U7405);
  nand ginst3339 (U2685, U7406, U7407);
  nand ginst3340 (U2686, U7408, U7409);
  nand ginst3341 (U2687, U7410, U7411);
  nand ginst3342 (U2688, U7412, U7413);
  nand ginst3343 (U2689, U7414, U7415);
  nand ginst3344 (U2690, U7416, U7417);
  nand ginst3345 (U2691, U7420, U7421);
  nand ginst3346 (U2692, U7422, U7423);
  nand ginst3347 (U2693, U7424, U7425);
  nand ginst3348 (U2694, U7426, U7427);
  nand ginst3349 (U2695, U7428, U7429);
  nand ginst3350 (U2696, U7430, U7431);
  nand ginst3351 (U2697, U7432, U7433);
  nand ginst3352 (U2698, U7434, U7435);
  nand ginst3353 (U2699, U7436, U7437);
  nand ginst3354 (U2700, U7438, U7439);
  nand ginst3355 (U2701, U7380, U7381);
  nand ginst3356 (U2702, U7382, U7383);
  nand ginst3357 (U2703, U7384, U7385);
  nand ginst3358 (U2704, U7386, U7387);
  nand ginst3359 (U2705, U7388, U7389);
  nand ginst3360 (U2706, U7390, U7391);
  nand ginst3361 (U2707, U7396, U7397);
  nand ginst3362 (U2708, U7418, U7419);
  nand ginst3363 (U2709, U7440, U7441);
  nand ginst3364 (U2710, U7442, U7443);
  nand ginst3365 (U2711, U7364, U7365);
  nand ginst3366 (U2712, U7366, U7367);
  nand ginst3367 (U2713, U4153, U4227);
  nand ginst3368 (U2714, U3421, U4154, U7373, U7374);
  nand ginst3369 (U2715, U4155, U4227);
  nand ginst3370 (U2716, U7352, U7353);
  nand ginst3371 (U2717, U7354, U7355);
  nand ginst3372 (U2718, U4149, U7356);
  nand ginst3373 (U2719, U4150, U7358);
  nand ginst3374 (U2720, U4151, U7360);
  nand ginst3375 (U2721, U4152, U7362);
  nand ginst3376 (U2722, U4147, U4180);
  and ginst3377 (U2723, U7071, U7224);
  and ginst3378 (U2724, U7071, U7241);
  and ginst3379 (U2725, U7071, U7258);
  and ginst3380 (U2726, U7071, U7608);
  and ginst3381 (U2727, U7071, U7290);
  and ginst3382 (U2728, U7071, U7307);
  and ginst3383 (U2729, U7071, U7324);
  and ginst3384 (U2730, U7071, U7341);
  nand ginst3385 (U2731, U2606, U7342);
  and ginst3386 (U2732, U7070, U7071);
  and ginst3387 (U2733, U7071, U7102);
  and ginst3388 (U2734, U7071, U7119);
  and ginst3389 (U2735, U7071, U7606);
  and ginst3390 (U2736, U7071, U7151);
  and ginst3391 (U2737, U7071, U7168);
  and ginst3392 (U2738, U7071, U7185);
  and ginst3393 (U2739, U7071, U7202);
  and ginst3394 (U2740, INSTQUEUERD_ADDR_REG_4__SCAN_IN, U7051);
  nand ginst3395 (U2741, U4066, U7084);
  and ginst3396 (U2742, U7479, U7480);
  and ginst3397 (U2743, U7458, U7494);
  and ginst3398 (U2744, U7466, U7467);
  nand ginst3399 (U2745, U7035, U7036);
  nand ginst3400 (U2746, U7037, U7038);
  nand ginst3401 (U2747, U7039, U7040);
  nand ginst3402 (U2748, U7041, U7604);
  nand ginst3403 (U2749, U7042, U7043);
  nand ginst3404 (U2750, U7044, U7045);
  nand ginst3405 (U2751, U4049, U7046);
  nand ginst3406 (U2752, U4050, U7048, U7049);
  and ginst3407 (U2753, U6897, U6945);
  and ginst3408 (U2754, U6897, U6962);
  and ginst3409 (U2755, U6897, U6979);
  and ginst3410 (U2756, U6897, U7603);
  and ginst3411 (U2757, U6897, U7011);
  and ginst3412 (U2758, U6897, U7028);
  and ginst3413 (U2759, U6896, U6897);
  and ginst3414 (U2760, U6897, U6914);
  nand ginst3415 (U2761, U6915, U6916);
  nand ginst3416 (U2762, U6917, U6918);
  nand ginst3417 (U2763, U6919, U6920);
  nand ginst3418 (U2764, U6921, U6922);
  nand ginst3419 (U2765, U6923, U6924, U6925);
  nand ginst3420 (U2766, U6926, U6927, U6928);
  nand ginst3421 (U2767, U7029, U7030, U7031);
  nand ginst3422 (U2768, U7032, U7033, U7034);
  and ginst3423 (U2769, R2144_U145, U4147);
  and ginst3424 (U2770, R2144_U145, U4147);
  and ginst3425 (U2771, R2144_U11, U4147);
  and ginst3426 (U2772, R2144_U37, U4147);
  and ginst3427 (U2773, R2144_U38, U4147);
  and ginst3428 (U2774, R2144_U39, U4147);
  and ginst3429 (U2775, R2144_U40, U4147);
  and ginst3430 (U2776, R2144_U41, U4147);
  and ginst3431 (U2777, R2144_U42, U4147);
  and ginst3432 (U2778, R2144_U30, U4147);
  nand ginst3433 (U2779, U6859, U6860);
  nand ginst3434 (U2780, U6861, U6862);
  nand ginst3435 (U2781, U6863, U6864);
  nand ginst3436 (U2782, U6865, U6866);
  nand ginst3437 (U2783, U6867, U6868);
  nand ginst3438 (U2784, U6869, U6870);
  nand ginst3439 (U2785, U6871, U6872, U6873);
  nand ginst3440 (U2786, U4016, U6874, U6875);
  nand ginst3441 (U2787, U6877, U6878, U6879);
  nand ginst3442 (U2788, U3419, U6605, U7486);
  nand ginst3443 (U2789, U6601, U7638);
  nand ginst3444 (U2790, U6599, U6600);
  nand ginst3445 (U2791, U4231, U7756, U7757);
  nand ginst3446 (U2792, U4231, U7752, U7753);
  nand ginst3447 (U2793, U4236, U6589);
  nand ginst3448 (U2794, U4228, U7744, U7745);
  nand ginst3449 (U2795, U4228, U7734, U7735);
  nand ginst3450 (U2796, U3936, U3937, U6579, U6581, U6583);
  nand ginst3451 (U2797, U3934, U3935, U6572, U6574, U6576);
  nand ginst3452 (U2798, U3932, U3933, U6565, U6567, U6569);
  nand ginst3453 (U2799, U3930, U3931, U6558, U6560, U6562);
  nand ginst3454 (U2800, U3928, U3929, U6551, U6553, U6555);
  nand ginst3455 (U2801, U3926, U3927, U6544, U6546, U6548);
  nand ginst3456 (U2802, U3924, U3925, U6537, U6539, U6541);
  nand ginst3457 (U2803, U3922, U3923, U6530, U6532, U6534);
  nand ginst3458 (U2804, U3920, U3921, U6523, U6525, U6527);
  nand ginst3459 (U2805, U3918, U3919, U6516, U6518, U6520);
  nand ginst3460 (U2806, U3916, U3917, U6509, U6511, U6513);
  nand ginst3461 (U2807, U3914, U3915, U6502, U6504, U6506);
  nand ginst3462 (U2808, U3912, U3913, U6495, U6497, U6499);
  nand ginst3463 (U2809, U3910, U3911, U6488, U6490, U6492);
  nand ginst3464 (U2810, U3908, U3909, U6481, U6483, U6485);
  nand ginst3465 (U2811, U3906, U3907, U6475, U6476, U6478);
  nand ginst3466 (U2812, U3904, U3905, U6468, U6469, U6471);
  nand ginst3467 (U2813, U3902, U3903, U6461, U6462, U6464);
  nand ginst3468 (U2814, U3900, U3901, U6454, U6455, U6457);
  nand ginst3469 (U2815, U3898, U3899, U6447, U6448, U6450);
  nand ginst3470 (U2816, U3896, U3897, U6440, U6441, U6443);
  nand ginst3471 (U2817, U3894, U3895, U6433, U6434, U6436);
  nand ginst3472 (U2818, U3892, U3893, U6426, U6427, U6429);
  nand ginst3473 (U2819, U3890, U3891, U6419, U6420, U6422);
  nand ginst3474 (U2820, U3888, U3889, U6412, U6413, U6415);
  nand ginst3475 (U2821, U3886, U3887, U6405, U6406, U6408);
  nand ginst3476 (U2822, U3884, U3885, U6397, U6398);
  nand ginst3477 (U2823, U3882, U3883, U6389, U6390, U6391);
  nand ginst3478 (U2824, U3881, U6380, U6381, U6382);
  nand ginst3479 (U2825, U3880, U6372, U6373, U6374);
  nand ginst3480 (U2826, U3879, U6364, U6365, U6366);
  nand ginst3481 (U2827, U3878, U6356, U6357, U6358);
  nand ginst3482 (U2828, U6346, U6347);
  nand ginst3483 (U2829, U6343, U6344, U6345);
  nand ginst3484 (U2830, U6340, U6341, U6342);
  nand ginst3485 (U2831, U6337, U6338, U6339);
  nand ginst3486 (U2832, U6334, U6335, U6336);
  nand ginst3487 (U2833, U6331, U6332, U6333);
  nand ginst3488 (U2834, U6328, U6329, U6330);
  nand ginst3489 (U2835, U6325, U6326, U6327);
  nand ginst3490 (U2836, U6322, U6323, U6324);
  nand ginst3491 (U2837, U6319, U6320, U6321);
  nand ginst3492 (U2838, U6316, U6317, U6318);
  nand ginst3493 (U2839, U6313, U6314, U6315);
  nand ginst3494 (U2840, U6310, U6311, U6312);
  nand ginst3495 (U2841, U6307, U6308, U6309);
  nand ginst3496 (U2842, U6304, U6305, U6306);
  nand ginst3497 (U2843, U6301, U6302, U6303);
  nand ginst3498 (U2844, U6298, U6299, U6300);
  nand ginst3499 (U2845, U6295, U6296, U6297);
  nand ginst3500 (U2846, U6292, U6293, U6294);
  nand ginst3501 (U2847, U6289, U6290, U6291);
  nand ginst3502 (U2848, U6286, U6287, U6288);
  nand ginst3503 (U2849, U6283, U6284, U6285);
  nand ginst3504 (U2850, U6280, U6281, U6282);
  nand ginst3505 (U2851, U6277, U6278, U6279);
  nand ginst3506 (U2852, U6274, U6275, U6276);
  nand ginst3507 (U2853, U6271, U6272, U6273);
  nand ginst3508 (U2854, U6268, U6269, U6270);
  nand ginst3509 (U2855, U6265, U6266, U6267);
  nand ginst3510 (U2856, U6262, U6263, U6264);
  nand ginst3511 (U2857, U6259, U6260, U6261);
  nand ginst3512 (U2858, U6256, U6257, U6258);
  nand ginst3513 (U2859, U6253, U6254, U6255);
  nand ginst3514 (U2860, U4164, U6250);
  nand ginst3515 (U2861, U6246, U6247, U6248, U6249);
  nand ginst3516 (U2862, U6242, U6243, U6244, U6245);
  nand ginst3517 (U2863, U6238, U6239, U6240, U6241);
  nand ginst3518 (U2864, U6234, U6235, U6236, U6237);
  nand ginst3519 (U2865, U6230, U6231, U6232, U6233);
  nand ginst3520 (U2866, U6226, U6227, U6228, U6229);
  nand ginst3521 (U2867, U6222, U6223, U6224, U6225);
  nand ginst3522 (U2868, U6218, U6219, U6220, U6221);
  nand ginst3523 (U2869, U6214, U6215, U6216, U6217);
  nand ginst3524 (U2870, U6210, U6211, U6212, U6213);
  nand ginst3525 (U2871, U6206, U6207, U6208, U6209);
  nand ginst3526 (U2872, U6202, U6203, U6204, U6205);
  nand ginst3527 (U2873, U6198, U6199, U6200, U6201);
  nand ginst3528 (U2874, U6194, U6195, U6196, U6197);
  nand ginst3529 (U2875, U6190, U6191, U6192, U6193);
  nand ginst3530 (U2876, U6187, U6188, U6189);
  nand ginst3531 (U2877, U6184, U6185, U6186);
  nand ginst3532 (U2878, U6181, U6182, U6183);
  nand ginst3533 (U2879, U6178, U6179, U6180);
  nand ginst3534 (U2880, U6175, U6176, U6177);
  nand ginst3535 (U2881, U6172, U6173, U6174);
  nand ginst3536 (U2882, U6169, U6170, U6171);
  nand ginst3537 (U2883, U6166, U6167, U6168);
  nand ginst3538 (U2884, U6163, U6164, U6165);
  nand ginst3539 (U2885, U6160, U6161, U6162);
  nand ginst3540 (U2886, U6157, U6158, U6159);
  nand ginst3541 (U2887, U6154, U6155, U6156);
  nand ginst3542 (U2888, U6151, U6152, U6153);
  nand ginst3543 (U2889, U6148, U6149, U6150);
  nand ginst3544 (U2890, U6145, U6146, U6147);
  nand ginst3545 (U2891, U6142, U6143, U6144);
  and ginst3546 (U2892, DATAO_REG_31__SCAN_IN, U6043);
  nand ginst3547 (U2893, U3870, U6134);
  nand ginst3548 (U2894, U3869, U6131);
  nand ginst3549 (U2895, U3868, U6128);
  nand ginst3550 (U2896, U3867, U6125);
  nand ginst3551 (U2897, U3866, U6122);
  nand ginst3552 (U2898, U3865, U6119);
  nand ginst3553 (U2899, U3864, U6116);
  nand ginst3554 (U2900, U3863, U6113);
  nand ginst3555 (U2901, U3862, U6110);
  nand ginst3556 (U2902, U3861, U6107);
  nand ginst3557 (U2903, U3860, U6104);
  nand ginst3558 (U2904, U3859, U6101);
  nand ginst3559 (U2905, U3858, U6098);
  nand ginst3560 (U2906, U3857, U6095);
  nand ginst3561 (U2907, U3856, U6092);
  nand ginst3562 (U2908, U6089, U6090, U6091);
  nand ginst3563 (U2909, U6086, U6087, U6088);
  nand ginst3564 (U2910, U6083, U6084, U6085);
  nand ginst3565 (U2911, U6080, U6081, U6082);
  nand ginst3566 (U2912, U6077, U6078, U6079);
  nand ginst3567 (U2913, U6074, U6075, U6076);
  nand ginst3568 (U2914, U6071, U6072, U6073);
  nand ginst3569 (U2915, U6068, U6069, U6070);
  nand ginst3570 (U2916, U6065, U6066, U6067);
  nand ginst3571 (U2917, U6062, U6063, U6064);
  nand ginst3572 (U2918, U6059, U6060, U6061);
  nand ginst3573 (U2919, U6056, U6057, U6058);
  nand ginst3574 (U2920, U6053, U6054, U6055);
  nand ginst3575 (U2921, U6050, U6051, U6052);
  nand ginst3576 (U2922, U6047, U6048, U6049);
  nand ginst3577 (U2923, U6044, U6045, U6046);
  nand ginst3578 (U2924, U7528, U7530);
  nand ginst3579 (U2925, U7527, U7532);
  nand ginst3580 (U2926, U7526, U7534);
  nand ginst3581 (U2927, U7525, U7536);
  nand ginst3582 (U2928, U7524, U7538);
  nand ginst3583 (U2929, U7523, U7540);
  nand ginst3584 (U2930, U7522, U7542);
  nand ginst3585 (U2931, U7521, U7544);
  nand ginst3586 (U2932, U7520, U7546);
  nand ginst3587 (U2933, U7519, U7548);
  nand ginst3588 (U2934, U7518, U7550);
  nand ginst3589 (U2935, U7517, U7552);
  nand ginst3590 (U2936, U7516, U7554);
  nand ginst3591 (U2937, U7515, U7556);
  nand ginst3592 (U2938, U7514, U7558);
  nand ginst3593 (U2939, U7513, U7560);
  nand ginst3594 (U2940, U7512, U7562);
  nand ginst3595 (U2941, U7511, U7564);
  nand ginst3596 (U2942, U7510, U7566);
  nand ginst3597 (U2943, U7509, U7568);
  nand ginst3598 (U2944, U7508, U7570);
  nand ginst3599 (U2945, U7507, U7572);
  nand ginst3600 (U2946, U7506, U7574);
  nand ginst3601 (U2947, U7505, U7576);
  nand ginst3602 (U2948, U7504, U7578);
  nand ginst3603 (U2949, U7503, U7580);
  nand ginst3604 (U2950, U7502, U7582);
  nand ginst3605 (U2951, U7501, U7584);
  nand ginst3606 (U2952, U7500, U7586);
  nand ginst3607 (U2953, U7499, U7588);
  nand ginst3608 (U2954, U7498, U7590);
  nand ginst3609 (U2955, U5942, U5943, U5944, U5945, U5946);
  nand ginst3610 (U2956, U5937, U5938, U5939, U5940, U5941);
  nand ginst3611 (U2957, U5932, U5933, U5934, U5935, U5936);
  nand ginst3612 (U2958, U5927, U5928, U5929, U5930, U5931);
  nand ginst3613 (U2959, U5922, U5923, U5924, U5925, U5926);
  nand ginst3614 (U2960, U5917, U5918, U5919, U5920, U5921);
  nand ginst3615 (U2961, U5912, U5913, U5914, U5915, U5916);
  nand ginst3616 (U2962, U5907, U5908, U5909, U5910, U5911);
  nand ginst3617 (U2963, U5902, U5903, U5904, U5905, U5906);
  nand ginst3618 (U2964, U5897, U5898, U5899, U5900, U5901);
  nand ginst3619 (U2965, U5892, U5893, U5894, U5895, U5896);
  nand ginst3620 (U2966, U5887, U5888, U5889, U5890, U5891);
  nand ginst3621 (U2967, U5882, U5883, U5884, U5885, U5886);
  nand ginst3622 (U2968, U5877, U5878, U5879, U5880, U5881);
  nand ginst3623 (U2969, U5872, U5873, U5874, U5875, U5876);
  nand ginst3624 (U2970, U5867, U5868, U5869, U5870, U5871);
  nand ginst3625 (U2971, U5862, U5863, U5864, U5865, U5866);
  nand ginst3626 (U2972, U5857, U5858, U5859, U5860, U5861);
  nand ginst3627 (U2973, U5852, U5853, U5854, U5855, U5856);
  nand ginst3628 (U2974, U5847, U5848, U5849, U5850, U5851);
  nand ginst3629 (U2975, U5842, U5843, U5844, U5845, U5846);
  nand ginst3630 (U2976, U5837, U5838, U5839, U5840, U5841);
  nand ginst3631 (U2977, U5832, U5833, U5834, U5835, U5836);
  nand ginst3632 (U2978, U5827, U5828, U5829, U5830, U5831);
  nand ginst3633 (U2979, U5822, U5823, U5824, U5825, U5826);
  nand ginst3634 (U2980, U5817, U5818, U5819, U5820, U5821);
  nand ginst3635 (U2981, U5812, U5813, U5814, U5815, U5816);
  nand ginst3636 (U2982, U5807, U5808, U5809, U5810, U5811);
  nand ginst3637 (U2983, U5802, U5803, U5804, U5805, U5806);
  nand ginst3638 (U2984, U5797, U5798, U5799, U5800, U5801);
  nand ginst3639 (U2985, U5792, U5793, U5794, U5795, U5796);
  nand ginst3640 (U2986, U5787, U5788, U5789, U5790, U5791);
  nand ginst3641 (U2987, U3847, U3849, U5775, U5777);
  nand ginst3642 (U2988, U3844, U3846, U5768, U5770);
  nand ginst3643 (U2989, U3841, U3843, U5761, U5763);
  nand ginst3644 (U2990, U3838, U3840, U5754, U5756);
  nand ginst3645 (U2991, U3835, U3837, U5747, U5749);
  nand ginst3646 (U2992, U3832, U3834, U5740, U5742);
  nand ginst3647 (U2993, U3829, U3831, U5733, U5735);
  nand ginst3648 (U2994, U3826, U3828, U5726, U5728);
  xor ginst3649 (U2995, restore_signal, U2995_pert);
  nand ginst3650 (U2995_in, U3823, U3825, U5719, U5721);
  xor ginst3651 (U2995_pert, U2995_in, perturb_signal);
  nand ginst3652 (U2996, U3820, U3822, U5712, U5714);
  nand ginst3653 (U2997, U3817, U3819, U5705, U5707);
  nand ginst3654 (U2998, U3814, U3816, U5698, U5700);
  nand ginst3655 (U2999, U3811, U3813, U5691, U5693);
  nand ginst3656 (U3000, U3808, U3810, U5684, U5686);
  nand ginst3657 (U3001, U3805, U3807, U5677, U5679);
  nand ginst3658 (U3002, U3802, U3804, U5670, U5672);
  nand ginst3659 (U3003, U3799, U3801, U5663, U5665);
  nand ginst3660 (U3004, U3796, U3798, U5656, U5658);
  nand ginst3661 (U3005, U3793, U3795, U5649, U5651);
  nand ginst3662 (U3006, U3790, U3792, U5644);
  nand ginst3663 (U3007, U3787, U3789, U5637);
  nand ginst3664 (U3008, U3784, U3786, U5630);
  nand ginst3665 (U3009, U3781, U3783, U5623);
  nand ginst3666 (U3010, U3778, U3780, U5616);
  nand ginst3667 (U3011, U3775, U3777, U5609);
  nand ginst3668 (U3012, U3772, U3774, U5602);
  nand ginst3669 (U3013, U3769, U3771, U5595);
  nand ginst3670 (U3014, U3766, U3768, U5588);
  nand ginst3671 (U3015, U3763, U3764);
  nand ginst3672 (U3016, U3759, U3760, U3762);
  nand ginst3673 (U3017, U3755, U3756, U3758);
  nand ginst3674 (U3018, U3751, U3752, U3754);
  and ginst3675 (U3019, INSTQUEUEWR_ADDR_REG_4__SCAN_IN, U5525);
  nand ginst3676 (U3020, U3718, U5447, U5448);
  nand ginst3677 (U3021, U3717, U5442, U5443);
  nand ginst3678 (U3022, U3716, U5437, U5438);
  nand ginst3679 (U3023, U3715, U5432, U5433);
  nand ginst3680 (U3024, U3714, U5428, U7600);
  nand ginst3681 (U3025, U3713, U5423, U5424);
  nand ginst3682 (U3026, U3712, U5418, U5419);
  nand ginst3683 (U3027, U3711, U5413, U5414);
  nand ginst3684 (U3028, U3709, U5391, U5392);
  nand ginst3685 (U3029, U3708, U5386, U5387);
  nand ginst3686 (U3030, U3707, U5381, U5382);
  nand ginst3687 (U3031, U3706, U5376, U5377);
  nand ginst3688 (U3032, U3705, U5371, U5372);
  nand ginst3689 (U3033, U3704, U5366, U5367);
  nand ginst3690 (U3034, U3703, U5361, U5362);
  nand ginst3691 (U3035, U3702, U5356, U5357);
  nand ginst3692 (U3036, U3700, U5333, U5334);
  nand ginst3693 (U3037, U3699, U5328, U5329);
  nand ginst3694 (U3038, U3698, U5323, U5324);
  nand ginst3695 (U3039, U3697, U5318, U5319);
  nand ginst3696 (U3040, U3696, U5313, U5314);
  nand ginst3697 (U3041, U3695, U5308, U5309);
  nand ginst3698 (U3042, U3694, U5303, U5304);
  nand ginst3699 (U3043, U3693, U5298, U5299);
  nand ginst3700 (U3044, U3691, U5276, U5277);
  nand ginst3701 (U3045, U3690, U5271, U5272);
  nand ginst3702 (U3046, U3689, U5266, U5267);
  nand ginst3703 (U3047, U3688, U5261, U5262);
  nand ginst3704 (U3048, U3687, U5256, U5257);
  nand ginst3705 (U3049, U3686, U5251, U5252);
  nand ginst3706 (U3050, U3685, U5246, U5247);
  nand ginst3707 (U3051, U3684, U5241, U5242);
  nand ginst3708 (U3052, U3682, U5218, U5219);
  nand ginst3709 (U3053, U3681, U5213, U5214);
  nand ginst3710 (U3054, U3680, U5208, U5209);
  nand ginst3711 (U3055, U3679, U5203, U5204);
  nand ginst3712 (U3056, U3678, U5198, U5199);
  nand ginst3713 (U3057, U3677, U5193, U5194);
  nand ginst3714 (U3058, U3676, U5188, U5189);
  nand ginst3715 (U3059, U3675, U5183, U5184);
  nand ginst3716 (U3060, U3673, U5161, U5162);
  nand ginst3717 (U3061, U3672, U5156, U5157);
  nand ginst3718 (U3062, U3671, U5151, U5152);
  nand ginst3719 (U3063, U3670, U5146, U5147);
  nand ginst3720 (U3064, U3669, U5141, U5142);
  nand ginst3721 (U3065, U3668, U5136, U5137);
  nand ginst3722 (U3066, U3667, U5131, U5132);
  nand ginst3723 (U3067, U3666, U5126, U5127);
  nand ginst3724 (U3068, U3664, U5103, U5104);
  nand ginst3725 (U3069, U3663, U5098, U5099);
  nand ginst3726 (U3070, U3662, U5093, U5094);
  nand ginst3727 (U3071, U3661, U5088, U5089);
  nand ginst3728 (U3072, U3660, U5083, U5084);
  nand ginst3729 (U3073, U3659, U5078, U5079);
  nand ginst3730 (U3074, U3658, U5073, U5074);
  nand ginst3731 (U3075, U3657, U5068, U5069);
  nand ginst3732 (U3076, U3655, U5046, U5047);
  nand ginst3733 (U3077, U3654, U5041, U5042);
  nand ginst3734 (U3078, U3653, U5036, U5037);
  nand ginst3735 (U3079, U3652, U5031, U5032);
  nand ginst3736 (U3080, U3651, U5026, U5027);
  nand ginst3737 (U3081, U3650, U5021, U5022);
  nand ginst3738 (U3082, U3649, U5016, U5017);
  nand ginst3739 (U3083, U3648, U5011, U5012);
  nand ginst3740 (U3084, U3646, U4990, U4991);
  nand ginst3741 (U3085, U3645, U4985, U4986);
  nand ginst3742 (U3086, U3644, U4980, U4981);
  nand ginst3743 (U3087, U3643, U4975, U4976);
  nand ginst3744 (U3088, U3642, U4970, U4971);
  nand ginst3745 (U3089, U3641, U4965, U4966);
  nand ginst3746 (U3090, U3640, U4960, U4961);
  nand ginst3747 (U3091, U3639, U4955, U4956);
  nand ginst3748 (U3092, U3637, U4933, U4934);
  nand ginst3749 (U3093, U3636, U4928, U4929);
  nand ginst3750 (U3094, U3635, U4923, U4924);
  nand ginst3751 (U3095, U3634, U4918, U4919);
  nand ginst3752 (U3096, U3633, U4913, U4914);
  nand ginst3753 (U3097, U3632, U4908, U4909);
  nand ginst3754 (U3098, U3631, U4903, U4904);
  nand ginst3755 (U3099, U3630, U4898, U4899);
  nand ginst3756 (U3100, U3628, U4875, U4876);
  nand ginst3757 (U3101, U3627, U4870, U4871);
  nand ginst3758 (U3102, U3626, U4865, U4866);
  nand ginst3759 (U3103, U3625, U4860, U4861);
  nand ginst3760 (U3104, U3624, U4855, U4856);
  nand ginst3761 (U3105, U3623, U4850, U4851);
  nand ginst3762 (U3106, U3622, U4845, U4846);
  nand ginst3763 (U3107, U3621, U4840, U4841);
  nand ginst3764 (U3108, U3619, U4818, U4819);
  nand ginst3765 (U3109, U3618, U4813, U4814);
  nand ginst3766 (U3110, U3617, U4808, U4809);
  nand ginst3767 (U3111, U3616, U4803, U4804);
  nand ginst3768 (U3112, U3615, U4798, U4799);
  nand ginst3769 (U3113, U3614, U4793, U4794);
  nand ginst3770 (U3114, U3613, U4788, U4789);
  nand ginst3771 (U3115, U3612, U4783, U4784);
  nand ginst3772 (U3116, U3610, U4760, U4761);
  nand ginst3773 (U3117, U3609, U4755, U4756);
  nand ginst3774 (U3118, U3608, U4750, U4751);
  nand ginst3775 (U3119, U3607, U4745, U4746);
  nand ginst3776 (U3120, U3606, U4740, U4741);
  nand ginst3777 (U3121, U3605, U4735, U4736);
  nand ginst3778 (U3122, U3604, U4730, U4731);
  nand ginst3779 (U3123, U3603, U4725, U4726);
  nand ginst3780 (U3124, U3601, U4703, U4704);
  nand ginst3781 (U3125, U3600, U4698, U4699);
  nand ginst3782 (U3126, U3599, U4693, U4694);
  nand ginst3783 (U3127, U3598, U4688, U4689);
  nand ginst3784 (U3128, U3597, U4683, U4684);
  nand ginst3785 (U3129, U3596, U4678, U4679);
  nand ginst3786 (U3130, U3595, U4673, U4674);
  nand ginst3787 (U3131, U3594, U4668, U4669);
  nand ginst3788 (U3132, U3592, U4644, U4645);
  nand ginst3789 (U3133, U3591, U4639, U4640);
  nand ginst3790 (U3134, U3590, U4634, U4635);
  nand ginst3791 (U3135, U3589, U4629, U4630);
  nand ginst3792 (U3136, U3588, U4624, U4625);
  nand ginst3793 (U3137, U3587, U4619, U4620);
  nand ginst3794 (U3138, U3586, U4614, U4615);
  nand ginst3795 (U3139, U3585, U4609, U4610);
  nand ginst3796 (U3140, U3583, U4586, U4587);
  nand ginst3797 (U3141, U3582, U4581, U4582);
  nand ginst3798 (U3142, U3581, U4576, U4577);
  nand ginst3799 (U3143, U3580, U4571, U4572);
  nand ginst3800 (U3144, U3579, U4566, U4567);
  nand ginst3801 (U3145, U3578, U4561, U4562);
  nand ginst3802 (U3146, U3577, U4556, U4557);
  nand ginst3803 (U3147, U3576, U4551, U4552);
  nand ginst3804 (U3148, U3574, U7677, U7678);
  nand ginst3805 (U3149, U4232, U4506, U4507, U4508);
  nand ginst3806 (U3150, U3570, U4504);
  and ginst3807 (U3151, DATAWIDTH_REG_31__SCAN_IN, U7638);
  and ginst3808 (U3152, DATAWIDTH_REG_30__SCAN_IN, U7638);
  and ginst3809 (U3153, DATAWIDTH_REG_29__SCAN_IN, U7638);
  and ginst3810 (U3154, DATAWIDTH_REG_28__SCAN_IN, U7638);
  and ginst3811 (U3155, DATAWIDTH_REG_27__SCAN_IN, U7638);
  and ginst3812 (U3156, DATAWIDTH_REG_26__SCAN_IN, U7638);
  and ginst3813 (U3157, DATAWIDTH_REG_25__SCAN_IN, U7638);
  and ginst3814 (U3158, DATAWIDTH_REG_24__SCAN_IN, U7638);
  and ginst3815 (U3159, DATAWIDTH_REG_23__SCAN_IN, U7638);
  and ginst3816 (U3160, DATAWIDTH_REG_22__SCAN_IN, U7638);
  and ginst3817 (U3161, DATAWIDTH_REG_21__SCAN_IN, U7638);
  and ginst3818 (U3162, DATAWIDTH_REG_20__SCAN_IN, U7638);
  and ginst3819 (U3163, DATAWIDTH_REG_19__SCAN_IN, U7638);
  and ginst3820 (U3164, DATAWIDTH_REG_18__SCAN_IN, U7638);
  and ginst3821 (U3165, DATAWIDTH_REG_17__SCAN_IN, U7638);
  and ginst3822 (U3166, DATAWIDTH_REG_16__SCAN_IN, U7638);
  and ginst3823 (U3167, DATAWIDTH_REG_15__SCAN_IN, U7638);
  and ginst3824 (U3168, DATAWIDTH_REG_14__SCAN_IN, U7638);
  and ginst3825 (U3169, DATAWIDTH_REG_13__SCAN_IN, U7638);
  and ginst3826 (U3170, DATAWIDTH_REG_12__SCAN_IN, U7638);
  and ginst3827 (U3171, DATAWIDTH_REG_11__SCAN_IN, U7638);
  and ginst3828 (U3172, DATAWIDTH_REG_10__SCAN_IN, U7638);
  and ginst3829 (U3173, DATAWIDTH_REG_9__SCAN_IN, U7638);
  and ginst3830 (U3174, DATAWIDTH_REG_8__SCAN_IN, U7638);
  and ginst3831 (U3175, DATAWIDTH_REG_7__SCAN_IN, U7638);
  and ginst3832 (U3176, DATAWIDTH_REG_6__SCAN_IN, U7638);
  and ginst3833 (U3177, DATAWIDTH_REG_5__SCAN_IN, U7638);
  and ginst3834 (U3178, DATAWIDTH_REG_4__SCAN_IN, U7638);
  and ginst3835 (U3179, DATAWIDTH_REG_3__SCAN_IN, U7638);
  and ginst3836 (U3180, DATAWIDTH_REG_2__SCAN_IN, U7638);
  nand ginst3837 (U3181, U4363, U7634, U7635);
  nand ginst3838 (U3182, U3483, U7632, U7633);
  nand ginst3839 (U3183, U3482, U4357);
  nand ginst3840 (U3184, U4342, U4343, U4344);
  nand ginst3841 (U3185, U4339, U4340, U4341);
  nand ginst3842 (U3186, U4336, U4337, U4338);
  nand ginst3843 (U3187, U4333, U4334, U4335);
  nand ginst3844 (U3188, U4330, U4331, U4332);
  nand ginst3845 (U3189, U4327, U4328, U4329);
  nand ginst3846 (U3190, U4324, U4325, U4326);
  nand ginst3847 (U3191, U4321, U4322, U4323);
  nand ginst3848 (U3192, U4318, U4319, U4320);
  nand ginst3849 (U3193, U4315, U4316, U4317);
  nand ginst3850 (U3194, U4312, U4313, U4314);
  nand ginst3851 (U3195, U4309, U4310, U4311);
  nand ginst3852 (U3196, U4306, U4307, U4308);
  nand ginst3853 (U3197, U4303, U4304, U4305);
  nand ginst3854 (U3198, U4300, U4301, U4302);
  nand ginst3855 (U3199, U4297, U4298, U4299);
  nand ginst3856 (U3200, U4294, U4295, U4296);
  nand ginst3857 (U3201, U4291, U4292, U4293);
  nand ginst3858 (U3202, U4288, U4289, U4290);
  nand ginst3859 (U3203, U4285, U4286, U4287);
  nand ginst3860 (U3204, U4282, U4283, U4284);
  nand ginst3861 (U3205, U4279, U4280, U4281);
  nand ginst3862 (U3206, U4276, U4277, U4278);
  nand ginst3863 (U3207, U4273, U4274, U4275);
  nand ginst3864 (U3208, U4270, U4271, U4272);
  nand ginst3865 (U3209, U4267, U4268, U4269);
  nand ginst3866 (U3210, U4264, U4265, U4266);
  nand ginst3867 (U3211, U4261, U4262, U4263);
  nand ginst3868 (U3212, U4258, U4259, U4260);
  nand ginst3869 (U3213, U4255, U4256, U4257);
  nand ginst3870 (U3214, U3986, U3987, U3988, U3989);
  nand ginst3871 (U3215, U3982, U3983, U3984, U3985);
  nand ginst3872 (U3216, U3978, U3979, U3980, U3981);
  nand ginst3873 (U3217, U3974, U3975, U3976, U3977);
  nand ginst3874 (U3218, U3970, U3971, U3972, U3973);
  nand ginst3875 (U3219, U3966, U3967, U3968, U3969);
  nand ginst3876 (U3220, U3962, U3963, U3964, U3965);
  nand ginst3877 (U3221, U3958, U3959, U3960, U3961);
  nand ginst3878 (U3222, U3310, U3316);
  nand ginst3879 (U3223, U2432, U3222);
  nand ginst3880 (U3224, U2432, U4531);
  nand ginst3881 (U3225, U2434, U3222);
  nand ginst3882 (U3226, U2434, U4531);
  nand ginst3883 (U3227, U2433, U3222);
  nand ginst3884 (U3228, U2433, U4531);
  nand ginst3885 (U3229, U2435, U3222);
  nand ginst3886 (U3230, U2435, U4531);
  nand ginst3887 (U3231, U3378, U3381, U5451);
  nand ginst3888 (U3232, U5452, U7074);
  nand ginst3889 (U3233, U4144, U4146, U7779, U7780);
  not ginst3890 (U3234, REQUESTPENDING_REG_SCAN_IN);
  not ginst3891 (U3235, STATE_REG_1__SCAN_IN);
  nand ginst3892 (U3236, STATE_REG_1__SCAN_IN, U3245);
  nand ginst3893 (U3237, U3238, U4209);
  not ginst3894 (U3238, STATE_REG_2__SCAN_IN);
  nand ginst3895 (U3239, STATE_REG_2__SCAN_IN, U4209);
  not ginst3896 (U3240, REIP_REG_1__SCAN_IN);
  nand ginst3897 (U3241, STATE_REG_1__SCAN_IN, U3238);
  or ginst3898 (U3242, STATE_REG_2__SCAN_IN, STATE_REG_1__SCAN_IN);
  not ginst3899 (U3243, HOLD);
  not ginst3900 (U3244, READY_N);
  not ginst3901 (U3245, STATE_REG_0__SCAN_IN);
  nand ginst3902 (U3246, STATE_REG_0__SCAN_IN, U3247);
  nand ginst3903 (U3247, REQUESTPENDING_REG_SCAN_IN, U3243);
  or ginst3904 (U3248, HOLD, REQUESTPENDING_REG_SCAN_IN);
  not ginst3905 (U3249, STATE2_REG_1__SCAN_IN);
  not ginst3906 (U3250, STATE2_REG_2__SCAN_IN);
  not ginst3907 (U3251, INSTQUEUERD_ADDR_REG_2__SCAN_IN);
  not ginst3908 (U3252, INSTQUEUERD_ADDR_REG_1__SCAN_IN);
  not ginst3909 (U3253, INSTQUEUERD_ADDR_REG_0__SCAN_IN);
  nand ginst3910 (U3254, INSTQUEUERD_ADDR_REG_2__SCAN_IN, INSTQUEUERD_ADDR_REG_1__SCAN_IN, INSTQUEUERD_ADDR_REG_0__SCAN_IN, U3257);
  or ginst3911 (U3255, INSTQUEUERD_ADDR_REG_2__SCAN_IN, INSTQUEUERD_ADDR_REG_1__SCAN_IN, INSTQUEUERD_ADDR_REG_0__SCAN_IN);
  or ginst3912 (U3256, INSTQUEUERD_ADDR_REG_1__SCAN_IN, INSTQUEUERD_ADDR_REG_0__SCAN_IN);
  not ginst3913 (U3257, INSTQUEUERD_ADDR_REG_3__SCAN_IN);
  nand ginst3914 (U3258, U3552, U3553, U3554, U3555);
  nand ginst3915 (U3259, U3245, U4484);
  not ginst3916 (U3260, R2167_U17);
  nand ginst3917 (U3261, INSTQUEUERD_ADDR_REG_2__SCAN_IN, U3257);
  nand ginst3918 (U3262, INSTQUEUERD_ADDR_REG_1__SCAN_IN, INSTQUEUERD_ADDR_REG_0__SCAN_IN);
  nand ginst3919 (U3263, U3504, U3505, U3506, U3507);
  nand ginst3920 (U3264, U3524, U3525, U3526, U3527, U4158);
  nand ginst3921 (U3265, U3542, U3543, U3544, U3545);
  nand ginst3922 (U3266, U3546, U3547);
  or ginst3923 (U3267, READY_N, STATEBS16_REG_SCAN_IN);
  nand ginst3924 (U3268, R2167_U17, U4485);
  nand ginst3925 (U3269, U3271, U4465);
  nand ginst3926 (U3270, U3496, U3497, U3498, U3499);
  nand ginst3927 (U3271, U3548, U3549, U3550, U3551);
  nand ginst3928 (U3272, U2473, U4489);
  nand ginst3929 (U3273, U2389, U3270);
  nand ginst3930 (U3274, U4465, U4482);
  nand ginst3931 (U3275, U2447, U4237);
  nand ginst3932 (U3276, U3265, U3378, U4161, U4448);
  nand ginst3933 (U3277, U3258, U3270);
  nand ginst3934 (U3278, U3271, U4178);
  nand ginst3935 (U3279, U2431, U4244);
  nand ginst3936 (U3280, LT_563_U6, U4166, U4213, U4497, U7614);
  not ginst3937 (U3281, STATE2_REG_0__SCAN_IN);
  nand ginst3938 (U3282, STATE2_REG_0__SCAN_IN, U7592);
  not ginst3939 (U3283, STATE2_REG_3__SCAN_IN);
  nand ginst3940 (U3284, STATE2_REG_2__SCAN_IN, U3249);
  or ginst3941 (U3285, STATE2_REG_2__SCAN_IN, STATE2_REG_1__SCAN_IN);
  nand ginst3942 (U3286, STATE2_REG_3__SCAN_IN, R2167_U17);
  nand ginst3943 (U3287, U3281, U4535);
  not ginst3944 (U3288, INSTQUEUEWR_ADDR_REG_0__SCAN_IN);
  not ginst3945 (U3289, INSTQUEUEWR_ADDR_REG_1__SCAN_IN);
  not ginst3946 (U3290, INSTQUEUEWR_ADDR_REG_3__SCAN_IN);
  not ginst3947 (U3291, INSTQUEUEWR_ADDR_REG_2__SCAN_IN);
  nand ginst3948 (U3292, INSTQUEUEWR_ADDR_REG_1__SCAN_IN, INSTQUEUEWR_ADDR_REG_0__SCAN_IN);
  nand ginst3949 (U3293, U2478, U4521);
  or ginst3950 (U3294, STATE2_REG_3__SCAN_IN, STATE2_REG_2__SCAN_IN);
  not ginst3951 (U3295, STATEBS16_REG_SCAN_IN);
  not ginst3952 (U3296, R2144_U43);
  not ginst3953 (U3297, R2144_U50);
  not ginst3954 (U3298, R2144_U49);
  not ginst3955 (U3299, R2144_U8);
  nand ginst3956 (U3300, R2144_U43, R2144_U50);
  nand ginst3957 (U3301, U3296, U3319);
  nand ginst3958 (U3302, U2475, U4515);
  not ginst3959 (U3303, R2182_U25);
  not ginst3960 (U3304, R2182_U42);
  not ginst3961 (U3305, R2182_U34);
  not ginst3962 (U3306, R2182_U33);
  nand ginst3963 (U3307, U3295, U4197);
  nand ginst3964 (U3308, U3293, U4523);
  nand ginst3965 (U3309, U3293, U4532);
  nand ginst3966 (U3310, INSTQUEUEWR_ADDR_REG_1__SCAN_IN, U3288);
  nand ginst3967 (U3311, U2478, U4530);
  nand ginst3968 (U3312, R2144_U50, U3296);
  nand ginst3969 (U3313, R2144_U43, U3319);
  nand ginst3970 (U3314, U2475, U4588);
  nand ginst3971 (U3315, U3311, U4591);
  nand ginst3972 (U3316, INSTQUEUEWR_ADDR_REG_0__SCAN_IN, U3289);
  nand ginst3973 (U3317, U2478, U4529);
  nand ginst3974 (U3318, R2144_U43, U3297);
  nand ginst3975 (U3319, U3312, U3318);
  nand ginst3976 (U3320, U3296, U4514);
  nand ginst3977 (U3321, U2475, U4646);
  nand ginst3978 (U3322, U3317, U4649);
  nand ginst3979 (U3323, U3317, U4651);
  nand ginst3980 (U3324, U2478, U2488);
  nand ginst3981 (U3325, U2475, U2485);
  nand ginst3982 (U3326, U3324, U4707);
  nand ginst3983 (U3327, INSTQUEUEWR_ADDR_REG_3__SCAN_IN, U3291);
  nand ginst3984 (U3328, U4521, U4526);
  nand ginst3985 (U3329, R2144_U8, U3298);
  nand ginst3986 (U3330, U2490, U4515);
  nand ginst3987 (U3331, U3328, U4764);
  nand ginst3988 (U3332, U3328, U4766);
  nand ginst3989 (U3333, U4526, U4530);
  nand ginst3990 (U3334, U2490, U4588);
  nand ginst3991 (U3335, U3333, U4822);
  nand ginst3992 (U3336, U4526, U4529);
  nand ginst3993 (U3337, U2490, U4646);
  nand ginst3994 (U3338, U3336, U4879);
  nand ginst3995 (U3339, U3336, U4881);
  nand ginst3996 (U3340, U2488, U4526);
  nand ginst3997 (U3341, U2485, U2490);
  nand ginst3998 (U3342, U3340, U4937);
  nand ginst3999 (U3343, U2479, U4521);
  nand ginst4000 (U3344, U2474, U4516);
  nand ginst4001 (U3345, U3329, U3344, U4518);
  nand ginst4002 (U3346, U2499, U4515);
  nand ginst4003 (U3347, U3327, U3343, U4527);
  nand ginst4004 (U3348, U3343, U4993);
  nand ginst4005 (U3349, U3343, U4995);
  nand ginst4006 (U3350, U2479, U4530);
  nand ginst4007 (U3351, U2499, U4588);
  nand ginst4008 (U3352, U3350, U5050);
  nand ginst4009 (U3353, U2479, U4529);
  nand ginst4010 (U3354, U2499, U4646);
  nand ginst4011 (U3355, U3353, U5107);
  nand ginst4012 (U3356, U3353, U5109);
  nand ginst4013 (U3357, U2479, U2488);
  nand ginst4014 (U3358, U2485, U2499);
  nand ginst4015 (U3359, U3357, U5165);
  nand ginst4016 (U3360, U2510, U4521);
  nand ginst4017 (U3361, U2507, U4515);
  nand ginst4018 (U3362, U3360, U5222);
  nand ginst4019 (U3363, U3360, U5224);
  nand ginst4020 (U3364, U2510, U4530);
  nand ginst4021 (U3365, U2507, U4588);
  nand ginst4022 (U3366, U3364, U5280);
  nand ginst4023 (U3367, U2510, U4529);
  nand ginst4024 (U3368, U2507, U4646);
  nand ginst4025 (U3369, U3367, U5337);
  nand ginst4026 (U3370, U3367, U5339);
  nand ginst4027 (U3371, U2488, U2510);
  nand ginst4028 (U3372, U2485, U2507);
  nand ginst4029 (U3373, U3371, U5395);
  not ginst4030 (U3374, FLUSH_REG_SCAN_IN);
  not ginst4031 (U3375, GTE_485_U6);
  nand ginst4032 (U3376, U3265, U3271);
  nand ginst4033 (U3377, U3258, U3271);
  nand ginst4034 (U3378, U3500, U3501, U3502, U3503);
  nand ginst4035 (U3379, U5477, U5478, U7616);
  nand ginst4036 (U3380, U3271, U4387);
  nand ginst4037 (U3381, U2605, U3264);
  nand ginst4038 (U3382, U4387, U4482, U7482);
  nand ginst4039 (U3383, U3729, U4235);
  nand ginst4040 (U3384, U2605, U4387, U4465, U4482, U7482);
  nand ginst4041 (U3385, U2605, U4159, U4388, U4437, U4448);
  nand ginst4042 (U3386, U4187, U4222, U4465);
  nand ginst4043 (U3387, U2447, U2449);
  nand ginst4044 (U3388, U3431, U5498);
  nand ginst4045 (U3389, U3256, U3262);
  not ginst4046 (U3390, LT_589_U6);
  nand ginst4047 (U3391, U3287, U4230, U5524);
  nand ginst4048 (U3392, STATE2_REG_0__SCAN_IN, U3265, U3271);
  nand ginst4049 (U3393, U3258, U3260);
  nand ginst4050 (U3394, U3264, U3378);
  nand ginst4051 (U3395, U2427, U3281);
  nand ginst4052 (U3396, U3378, U4448);
  nand ginst4053 (U3397, U3265, U4241);
  nand ginst4054 (U3398, U2452, U4178);
  nand ginst4055 (U3399, STATE2_REG_2__SCAN_IN, U3258);
  not ginst4056 (U3400, REIP_REG_0__SCAN_IN);
  nand ginst4057 (U3401, U3744, U5550);
  nand ginst4058 (U3402, U4161, U4388);
  nand ginst4059 (U3403, U3851, U4236);
  nand ginst4060 (U3404, U6041, U6042);
  nand ginst4061 (U3405, STATE2_REG_0__SCAN_IN, U4482);
  nand ginst4062 (U3406, U4387, U7482);
  nand ginst4063 (U3407, U4194, U4465);
  nand ginst4064 (U3408, U2431, U4182);
  nand ginst4065 (U3409, STATE2_REG_0__SCAN_IN, U4198);
  nand ginst4066 (U3410, U3378, U4491);
  nand ginst4067 (U3411, U4223, U6141);
  nand ginst4068 (U3412, STATE2_REG_0__SCAN_IN, U4204);
  nand ginst4069 (U3413, U4223, U6252);
  nand ginst4070 (U3414, STATE2_REG_0__SCAN_IN, U2452, U3874, U4237);
  nand ginst4071 (U3415, U2447, U3854);
  not ginst4072 (U3416, EBX_REG_31__SCAN_IN);
  not ginst4073 (U3417, R2337_U58);
  nand ginst4074 (U3418, U3875, U4216);
  nand ginst4075 (U3419, U3249, U4197);
  nand ginst4076 (U3420, U3940, U3943, U3946, U3950);
  nand ginst4077 (U3421, U3258, U4194);
  not ginst4078 (U3422, CODEFETCH_REG_SCAN_IN);
  not ginst4079 (U3423, READREQUEST_REG_SCAN_IN);
  nand ginst4080 (U3424, U2447, U4486);
  nand ginst4081 (U3425, U3254, U5470);
  nand ginst4082 (U3426, STATE2_REG_2__SCAN_IN, U4437);
  nand ginst4083 (U3427, STATEBS16_REG_SCAN_IN, U3250);
  not ginst4084 (U3428, U3221);
  nand ginst4085 (U3429, U5466, U5467);
  nand ginst4086 (U3430, U2450, U3428);
  nand ginst4087 (U3431, INSTQUEUERD_ADDR_REG_1__SCAN_IN, INSTQUEUERD_ADDR_REG_0__SCAN_IN, U3251);
  nand ginst4088 (U3432, U3261, U7052);
  nand ginst4089 (U3433, U4185, U4222);
  nand ginst4090 (U3434, U4219, U4238, U4388);
  nand ginst4091 (U3435, U3265, U4219, U4238);
  nand ginst4092 (U3436, U4465, U4484);
  nand ginst4093 (U3437, U4062, U4063, U4065, U7081);
  nand ginst4094 (U3438, U4242, U4254);
  nand ginst4095 (U3439, U3255, U4171);
  nand ginst4096 (U3440, STATE2_REG_0__SCAN_IN, U2605);
  nand ginst4097 (U3441, U7679, U7680);
  nand ginst4098 (U3442, U7682, U7683);
  nand ginst4099 (U3443, U7706, U7707);
  nand ginst4100 (U3444, U7776, U7777);
  nand ginst4101 (U3445, U7621, U7622);
  nand ginst4102 (U3446, U7623, U7624);
  nand ginst4103 (U3447, U7625, U7626);
  nand ginst4104 (U3448, U7627, U7628);
  nand ginst4105 (U3449, U7636, U7637);
  and ginst4106 (U3450, U3242, U4167);
  nand ginst4107 (U3451, U7639, U7640);
  nand ginst4108 (U3452, U7641, U7642);
  nand ginst4109 (U3453, U7673, U7674);
  and ginst4110 (U3454, R2182_U24, U2427, U4203);
  nand ginst4111 (U3455, U7689, U7690);
  nand ginst4112 (U3456, U7696, U7697);
  nand ginst4113 (U3457, U7698, U7699);
  nand ginst4114 (U3458, U7701, U7702);
  nand ginst4115 (U3459, U7709, U7710);
  nand ginst4116 (U3460, U7711, U7712);
  nand ginst4117 (U3461, U7715, U7716);
  nand ginst4118 (U3462, U7717, U7718);
  nand ginst4119 (U3463, U7722, U7723);
  nand ginst4120 (U3464, U7724, U7725);
  nand ginst4121 (U3465, U7726, U7727);
  and ginst4122 (U3466, R2358_U91, U4437);
  nor ginst4123 (U3467, DATAWIDTH_REG_1__SCAN_IN, REIP_REG_1__SCAN_IN);
  nand ginst4124 (U3468, U7742, U7743);
  nand ginst4125 (U3469, U7746, U7747);
  nand ginst4126 (U3470, U7748, U7749);
  nand ginst4127 (U3471, U7750, U7751);
  nand ginst4128 (U3472, U7754, U7755);
  nand ginst4129 (U3473, U7758, U7759);
  nand ginst4130 (U3474, U7760, U7761);
  and ginst4131 (U3475, R2182_U24, U4203);
  nand ginst4132 (U3476, U7762, U7763);
  nand ginst4133 (U3477, U7764, U7765);
  nand ginst4134 (U3478, U7766, U7767);
  nand ginst4135 (U3479, U7768, U7769);
  nand ginst4136 (U3480, U7770, U7771);
  and ginst4137 (U3481, READY_N, STATE_REG_1__SCAN_IN);
  and ginst4138 (U3482, U3239, U4356);
  and ginst4139 (U3483, U3237, U4358);
  and ginst4140 (U3484, REQUESTPENDING_REG_SCAN_IN, STATE_REG_0__SCAN_IN);
  nor ginst4141 (U3485, INSTQUEUERD_ADDR_REG_3__SCAN_IN, INSTQUEUERD_ADDR_REG_2__SCAN_IN);
  and ginst4142 (U3486, INSTQUEUERD_ADDR_REG_1__SCAN_IN, INSTQUEUERD_ADDR_REG_0__SCAN_IN);
  nor ginst4143 (U3487, INSTQUEUERD_ADDR_REG_3__SCAN_IN, INSTQUEUERD_ADDR_REG_1__SCAN_IN);
  and ginst4144 (U3488, INSTQUEUERD_ADDR_REG_2__SCAN_IN, INSTQUEUERD_ADDR_REG_0__SCAN_IN);
  nor ginst4145 (U3489, INSTQUEUERD_ADDR_REG_3__SCAN_IN, INSTQUEUERD_ADDR_REG_0__SCAN_IN);
  and ginst4146 (U3490, INSTQUEUERD_ADDR_REG_2__SCAN_IN, INSTQUEUERD_ADDR_REG_1__SCAN_IN);
  nor ginst4147 (U3491, INSTQUEUERD_ADDR_REG_2__SCAN_IN, INSTQUEUERD_ADDR_REG_1__SCAN_IN);
  and ginst4148 (U3492, INSTQUEUERD_ADDR_REG_3__SCAN_IN, INSTQUEUERD_ADDR_REG_0__SCAN_IN);
  nor ginst4149 (U3493, INSTQUEUERD_ADDR_REG_2__SCAN_IN, INSTQUEUERD_ADDR_REG_0__SCAN_IN);
  and ginst4150 (U3494, INSTQUEUERD_ADDR_REG_3__SCAN_IN, INSTQUEUERD_ADDR_REG_1__SCAN_IN);
  and ginst4151 (U3495, INSTQUEUERD_ADDR_REG_3__SCAN_IN, INSTQUEUERD_ADDR_REG_2__SCAN_IN);
  and ginst4152 (U3496, U4371, U4372, U4373, U4374);
  and ginst4153 (U3497, U4375, U4376, U4377, U4378);
  and ginst4154 (U3498, U4379, U4380, U4381, U4382);
  and ginst4155 (U3499, U4383, U4384, U4385, U4386);
  and ginst4156 (U3500, U4421, U4422, U4423, U4424);
  and ginst4157 (U3501, U4425, U4426, U4427, U4428);
  and ginst4158 (U3502, U4429, U4430, U4431, U4432);
  and ginst4159 (U3503, U4433, U4434, U4435, U4436);
  and ginst4160 (U3504, U4404, U4405, U4406, U4407);
  and ginst4161 (U3505, U4408, U4409, U4410, U4411);
  and ginst4162 (U3506, U4412, U4413, U4414, U4415);
  and ginst4163 (U3507, U4416, U4417, U4418, U4419);
  nor ginst4164 (U3508, INSTQUEUERD_ADDR_REG_3__SCAN_IN, INSTQUEUERD_ADDR_REG_1__SCAN_IN);
  and ginst4165 (U3509, INSTQUEUE_REG_5__5__SCAN_IN, INSTQUEUERD_ADDR_REG_0__SCAN_IN);
  nor ginst4166 (U3510, INSTQUEUERD_ADDR_REG_3__SCAN_IN, INSTQUEUERD_ADDR_REG_0__SCAN_IN);
  and ginst4167 (U3511, INSTQUEUE_REG_6__5__SCAN_IN, INSTQUEUERD_ADDR_REG_1__SCAN_IN);
  and ginst4168 (U3512, INSTQUEUE_REG_8__5__SCAN_IN, INSTQUEUERD_ADDR_REG_3__SCAN_IN);
  nor ginst4169 (U3513, INSTQUEUERD_ADDR_REG_2__SCAN_IN, INSTQUEUERD_ADDR_REG_0__SCAN_IN);
  and ginst4170 (U3514, INSTQUEUE_REG_10__5__SCAN_IN, INSTQUEUERD_ADDR_REG_3__SCAN_IN);
  and ginst4171 (U3515, INSTQUEUE_REG_12__5__SCAN_IN, INSTQUEUERD_ADDR_REG_3__SCAN_IN);
  nor ginst4172 (U3516, INSTQUEUERD_ADDR_REG_2__SCAN_IN, INSTQUEUERD_ADDR_REG_1__SCAN_IN);
  and ginst4173 (U3517, INSTQUEUE_REG_9__5__SCAN_IN, INSTQUEUERD_ADDR_REG_0__SCAN_IN);
  and ginst4174 (U3518, U4389, U4390, U4391, U4392);
  and ginst4175 (U3519, U4393, U4394, U4395, U4396);
  and ginst4176 (U3520, U4397, U4398, U4399, U4400);
  and ginst4177 (U3521, U4401, U4402);
  nor ginst4178 (U3522, INSTQUEUERD_ADDR_REG_3__SCAN_IN, INSTQUEUERD_ADDR_REG_2__SCAN_IN);
  and ginst4179 (U3523, INSTQUEUE_REG_3__6__SCAN_IN, INSTQUEUERD_ADDR_REG_0__SCAN_IN);
  and ginst4180 (U3524, U4438, U4439, U4440, U4441);
  and ginst4181 (U3525, U4442, U4443, U4444);
  and ginst4182 (U3526, U4445, U4446, U4447);
  and ginst4183 (U3527, U7663, U7664, U7665, U7666);
  nor ginst4184 (U3528, INSTQUEUERD_ADDR_REG_3__SCAN_IN, INSTQUEUERD_ADDR_REG_2__SCAN_IN);
  and ginst4185 (U3529, INSTQUEUE_REG_1__4__SCAN_IN, INSTQUEUERD_ADDR_REG_0__SCAN_IN);
  nor ginst4186 (U3530, INSTQUEUERD_ADDR_REG_1__SCAN_IN, INSTQUEUERD_ADDR_REG_0__SCAN_IN);
  and ginst4187 (U3531, INSTQUEUE_REG_4__4__SCAN_IN, INSTQUEUERD_ADDR_REG_2__SCAN_IN);
  nor ginst4188 (U3532, INSTQUEUERD_ADDR_REG_1__SCAN_IN, INSTQUEUERD_ADDR_REG_0__SCAN_IN);
  and ginst4189 (U3533, INSTQUEUE_REG_12__4__SCAN_IN, INSTQUEUERD_ADDR_REG_2__SCAN_IN);
  and ginst4190 (U3534, INSTQUEUERD_ADDR_REG_2__SCAN_IN, INSTQUEUERD_ADDR_REG_0__SCAN_IN);
  and ginst4191 (U3535, INSTQUEUE_REG_13__4__SCAN_IN, INSTQUEUERD_ADDR_REG_3__SCAN_IN);
  nor ginst4192 (U3536, INSTQUEUERD_ADDR_REG_3__SCAN_IN, INSTQUEUERD_ADDR_REG_0__SCAN_IN);
  and ginst4193 (U3537, INSTQUEUE_REG_6__4__SCAN_IN, INSTQUEUERD_ADDR_REG_2__SCAN_IN);
  and ginst4194 (U3538, INSTQUEUERD_ADDR_REG_2__SCAN_IN, INSTQUEUERD_ADDR_REG_1__SCAN_IN);
  and ginst4195 (U3539, INSTQUEUE_REG_14__4__SCAN_IN, INSTQUEUERD_ADDR_REG_3__SCAN_IN);
  nor ginst4196 (U3540, INSTQUEUERD_ADDR_REG_2__SCAN_IN, INSTQUEUERD_ADDR_REG_1__SCAN_IN);
  and ginst4197 (U3541, INSTQUEUE_REG_9__4__SCAN_IN, INSTQUEUERD_ADDR_REG_3__SCAN_IN);
  and ginst4198 (U3542, U7643, U7644, U7645, U7646);
  and ginst4199 (U3543, U7647, U7648, U7649, U7650);
  and ginst4200 (U3544, U7651, U7652, U7653, U7654);
  and ginst4201 (U3545, U7655, U7656, U7657, U7658);
  and ginst4202 (U3546, U3270, U3378, U7482);
  and ginst4203 (U3547, U2605, U4388, U4448);
  and ginst4204 (U3548, U4466, U4467, U4468, U4469);
  and ginst4205 (U3549, U4470, U4471, U4472, U4473);
  and ginst4206 (U3550, U4474, U4475, U4476, U4477);
  and ginst4207 (U3551, U4478, U4479, U4480, U4481);
  and ginst4208 (U3552, U4449, U4450, U4451, U4452);
  and ginst4209 (U3553, U4453, U4454, U4455, U4456);
  and ginst4210 (U3554, U4457, U4458, U4459, U4460);
  and ginst4211 (U3555, U4461, U4462, U4463, U4464);
  and ginst4212 (U3556, U4196, U4365);
  and ginst4213 (U3557, U4404, U4405, U4406, U4407);
  and ginst4214 (U3558, U4408, U4409, U4410, U4411);
  and ginst4215 (U3559, U4412, U4413, U4414, U4415);
  and ginst4216 (U3560, U4416, U4417, U4418, U4419);
  and ginst4217 (U3561, U4389, U4390, U4391, U4392);
  and ginst4218 (U3562, U4393, U4394, U4395, U4396);
  and ginst4219 (U3563, U4397, U4398, U4399, U4400);
  and ginst4220 (U3564, U4401, U4402);
  and ginst4221 (U3565, U4159, U4387);
  and ginst4222 (U3566, U3270, U4237);
  and ginst4223 (U3567, U3270, U3271, U4388, U7482);
  and ginst4224 (U3568, U3387, U4205);
  and ginst4225 (U3569, STATE2_REG_2__SCAN_IN, U7591);
  and ginst4226 (U3570, U3284, U4503);
  and ginst4227 (U3571, U2427, U3244);
  and ginst4228 (U3572, STATE2_REG_3__SCAN_IN, STATE2_REG_0__SCAN_IN);
  and ginst4229 (U3573, U4229, U4234);
  and ginst4230 (U3574, U3573, U4511);
  and ginst4231 (U3575, U4212, U4540, U4541);
  and ginst4232 (U3576, U4548, U4549, U4550);
  and ginst4233 (U3577, U4553, U4554, U4555);
  and ginst4234 (U3578, U4558, U4559, U4560);
  and ginst4235 (U3579, U4563, U4564, U4565);
  and ginst4236 (U3580, U4568, U4569, U4570);
  and ginst4237 (U3581, U4573, U4574, U4575);
  and ginst4238 (U3582, U4578, U4579, U4580);
  and ginst4239 (U3583, U4583, U4584, U4585);
  and ginst4240 (U3584, U4212, U4598, U4599);
  and ginst4241 (U3585, U4606, U4607, U4608);
  and ginst4242 (U3586, U4611, U4612, U4613);
  and ginst4243 (U3587, U4616, U4617, U4618);
  and ginst4244 (U3588, U4621, U4622, U4623);
  and ginst4245 (U3589, U4626, U4627, U4628);
  and ginst4246 (U3590, U4631, U4632, U4633);
  and ginst4247 (U3591, U4636, U4637, U4638);
  and ginst4248 (U3592, U4641, U4642, U4643);
  and ginst4249 (U3593, U4212, U4657, U4658);
  and ginst4250 (U3594, U4665, U4666, U4667);
  and ginst4251 (U3595, U4670, U4671, U4672);
  and ginst4252 (U3596, U4675, U4676, U4677);
  and ginst4253 (U3597, U4680, U4681, U4682);
  and ginst4254 (U3598, U4685, U4686, U4687);
  and ginst4255 (U3599, U4690, U4691, U4692);
  and ginst4256 (U3600, U4695, U4696, U4697);
  and ginst4257 (U3601, U4700, U4701, U4702);
  and ginst4258 (U3602, U4212, U4714, U4715);
  and ginst4259 (U3603, U4722, U4723, U4724);
  and ginst4260 (U3604, U4727, U4728, U4729);
  and ginst4261 (U3605, U4732, U4733, U4734);
  and ginst4262 (U3606, U4737, U4738, U4739);
  and ginst4263 (U3607, U4742, U4743, U4744);
  and ginst4264 (U3608, U4747, U4748, U4749);
  and ginst4265 (U3609, U4752, U4753, U4754);
  and ginst4266 (U3610, U4757, U4758, U4759);
  and ginst4267 (U3611, U4212, U4772, U4773);
  and ginst4268 (U3612, U4780, U4781, U4782);
  and ginst4269 (U3613, U4785, U4786, U4787);
  and ginst4270 (U3614, U4790, U4791, U4792);
  and ginst4271 (U3615, U4795, U4796, U4797);
  and ginst4272 (U3616, U4800, U4801, U4802);
  and ginst4273 (U3617, U4805, U4806, U4807);
  and ginst4274 (U3618, U4810, U4811, U4812);
  and ginst4275 (U3619, U4815, U4816, U4817);
  and ginst4276 (U3620, U4212, U4829, U4830);
  and ginst4277 (U3621, U4837, U4838, U4839);
  and ginst4278 (U3622, U4842, U4843, U4844);
  and ginst4279 (U3623, U4847, U4848, U4849);
  and ginst4280 (U3624, U4852, U4853, U4854);
  and ginst4281 (U3625, U4857, U4858, U4859);
  and ginst4282 (U3626, U4862, U4863, U4864);
  and ginst4283 (U3627, U4867, U4868, U4869);
  and ginst4284 (U3628, U4872, U4873, U4874);
  and ginst4285 (U3629, U4212, U4887, U4888);
  and ginst4286 (U3630, U4895, U4896, U4897);
  and ginst4287 (U3631, U4900, U4901, U4902);
  and ginst4288 (U3632, U4905, U4906, U4907);
  and ginst4289 (U3633, U4910, U4911, U4912);
  and ginst4290 (U3634, U4915, U4916, U4917);
  and ginst4291 (U3635, U4920, U4921, U4922);
  and ginst4292 (U3636, U4925, U4926, U4927);
  and ginst4293 (U3637, U4930, U4931, U4932);
  and ginst4294 (U3638, U4212, U4944, U4945);
  and ginst4295 (U3639, U4952, U4953, U4954);
  and ginst4296 (U3640, U4957, U4958, U4959);
  and ginst4297 (U3641, U4962, U4963, U4964);
  and ginst4298 (U3642, U4967, U4968, U4969);
  and ginst4299 (U3643, U4972, U4973, U4974);
  and ginst4300 (U3644, U4977, U4978, U4979);
  and ginst4301 (U3645, U4982, U4983, U4984);
  and ginst4302 (U3646, U4987, U4988, U4989);
  and ginst4303 (U3647, U4212, U5000, U5001);
  and ginst4304 (U3648, U5008, U5009, U5010);
  and ginst4305 (U3649, U5013, U5014, U5015);
  and ginst4306 (U3650, U5018, U5019, U5020);
  and ginst4307 (U3651, U5023, U5024, U5025);
  and ginst4308 (U3652, U5028, U5029, U5030);
  and ginst4309 (U3653, U5033, U5034, U5035);
  and ginst4310 (U3654, U5038, U5039, U5040);
  and ginst4311 (U3655, U5043, U5044, U5045);
  and ginst4312 (U3656, U4212, U5057, U5058);
  and ginst4313 (U3657, U5065, U5066, U5067);
  and ginst4314 (U3658, U5070, U5071, U5072);
  and ginst4315 (U3659, U5075, U5076, U5077);
  and ginst4316 (U3660, U5080, U5081, U5082);
  and ginst4317 (U3661, U5085, U5086, U5087);
  and ginst4318 (U3662, U5090, U5091, U5092);
  and ginst4319 (U3663, U5095, U5096, U5097);
  and ginst4320 (U3664, U5100, U5101, U5102);
  and ginst4321 (U3665, U4212, U5115, U5116);
  and ginst4322 (U3666, U5123, U5124, U5125);
  and ginst4323 (U3667, U5128, U5129, U5130);
  and ginst4324 (U3668, U5133, U5134, U5135);
  and ginst4325 (U3669, U5138, U5139, U5140);
  and ginst4326 (U3670, U5143, U5144, U5145);
  and ginst4327 (U3671, U5148, U5149, U5150);
  and ginst4328 (U3672, U5153, U5154, U5155);
  and ginst4329 (U3673, U5158, U5159, U5160);
  and ginst4330 (U3674, U4212, U5172, U5173);
  and ginst4331 (U3675, U5180, U5181, U5182);
  and ginst4332 (U3676, U5185, U5186, U5187);
  and ginst4333 (U3677, U5190, U5191, U5192);
  and ginst4334 (U3678, U5195, U5196, U5197);
  and ginst4335 (U3679, U5200, U5201, U5202);
  and ginst4336 (U3680, U5205, U5206, U5207);
  and ginst4337 (U3681, U5210, U5211, U5212);
  and ginst4338 (U3682, U5215, U5216, U5217);
  and ginst4339 (U3683, U4212, U5230, U5231);
  and ginst4340 (U3684, U5238, U5239, U5240);
  and ginst4341 (U3685, U5243, U5244, U5245);
  and ginst4342 (U3686, U5248, U5249, U5250);
  and ginst4343 (U3687, U5253, U5254, U5255);
  and ginst4344 (U3688, U5258, U5259, U5260);
  and ginst4345 (U3689, U5263, U5264, U5265);
  and ginst4346 (U3690, U5268, U5269, U5270);
  and ginst4347 (U3691, U5273, U5274, U5275);
  and ginst4348 (U3692, U4212, U5287, U5288);
  and ginst4349 (U3693, U5295, U5296, U5297);
  and ginst4350 (U3694, U5300, U5301, U5302);
  and ginst4351 (U3695, U5305, U5306, U5307);
  and ginst4352 (U3696, U5310, U5311, U5312);
  and ginst4353 (U3697, U5315, U5316, U5317);
  and ginst4354 (U3698, U5320, U5321, U5322);
  and ginst4355 (U3699, U5325, U5326, U5327);
  and ginst4356 (U3700, U5330, U5331, U5332);
  and ginst4357 (U3701, U4212, U5345, U5346);
  and ginst4358 (U3702, U5353, U5354, U5355);
  and ginst4359 (U3703, U5358, U5359, U5360);
  and ginst4360 (U3704, U5363, U5364, U5365);
  and ginst4361 (U3705, U5368, U5369, U5370);
  and ginst4362 (U3706, U5373, U5374, U5375);
  and ginst4363 (U3707, U5378, U5379, U5380);
  and ginst4364 (U3708, U5383, U5384, U5385);
  and ginst4365 (U3709, U5388, U5389, U5390);
  and ginst4366 (U3710, U4212, U5402, U5403);
  and ginst4367 (U3711, U5410, U5411, U5412);
  and ginst4368 (U3712, U5415, U5416, U5417);
  and ginst4369 (U3713, U5420, U5421, U5422);
  and ginst4370 (U3714, U5425, U5426, U5427);
  and ginst4371 (U3715, U5429, U5430, U5431);
  and ginst4372 (U3716, U5434, U5435, U5436);
  and ginst4373 (U3717, U5439, U5440, U5441);
  and ginst4374 (U3718, U5444, U5445, U5446);
  and ginst4375 (U3719, FLUSH_REG_SCAN_IN, STATE2_REG_0__SCAN_IN);
  and ginst4376 (U3720, U4387, U4482);
  and ginst4377 (U3721, U3244, U4485);
  and ginst4378 (U3722, U3244, U4198);
  and ginst4379 (U3723, U4205, U7484);
  and ginst4380 (U3724, U5459, U5460);
  and ginst4381 (U3725, U3724, U5458);
  and ginst4382 (U3726, U2518, U3725);
  and ginst4383 (U3727, U4230, U5463);
  and ginst4384 (U3728, U5473, U5474);
  and ginst4385 (U3729, U4388, U4437);
  and ginst4386 (U3730, U3380, U5484);
  and ginst4387 (U3731, U5485, U5486);
  and ginst4388 (U3732, U3730, U3731, U5488, U7615);
  and ginst4389 (U3733, U3384, U4251);
  and ginst4390 (U3734, U2520, U3266, U3275, U3398, U3733);
  and ginst4391 (U3735, U3736, U5490);
  and ginst4392 (U3736, U5492, U5493);
  and ginst4393 (U3737, U5501, U7704, U7705);
  and ginst4394 (U3738, U5510, U5512);
  and ginst4395 (U3739, U5531, U5532);
  and ginst4396 (U3740, U5535, U5536);
  and ginst4397 (U3741, U5540, U5541);
  and ginst4398 (U3742, U3244, U5546);
  and ginst4399 (U3743, U3271, U3394);
  and ginst4400 (U3744, U5549, U5551);
  and ginst4401 (U3745, U3385, U3386, U5555);
  and ginst4402 (U3746, U2520, U3745, U5556);
  and ginst4403 (U3747, U3271, U4174);
  and ginst4404 (U3748, U3275, U3435, U4205);
  and ginst4405 (U3749, U5554, U7495);
  and ginst4406 (U3750, STATE2_REG_2__SCAN_IN, U7496);
  and ginst4407 (U3751, U5558, U5559);
  and ginst4408 (U3752, U5560, U5561);
  and ginst4409 (U3753, U5563, U5564);
  and ginst4410 (U3754, U3753, U5562);
  and ginst4411 (U3755, U5565, U5566);
  and ginst4412 (U3756, U5567, U5568);
  and ginst4413 (U3757, U5570, U5571);
  and ginst4414 (U3758, U3757, U5569);
  and ginst4415 (U3759, U5572, U5573);
  and ginst4416 (U3760, U5574, U5575);
  and ginst4417 (U3761, U5577, U5578);
  and ginst4418 (U3762, U3761, U5576);
  and ginst4419 (U3763, U5579, U5580, U5582);
  and ginst4420 (U3764, U3765, U5581, U5583);
  and ginst4421 (U3765, U5584, U5585);
  and ginst4422 (U3766, U5586, U5587, U5589);
  and ginst4423 (U3767, U5591, U5592);
  and ginst4424 (U3768, U3767, U5590);
  and ginst4425 (U3769, U5593, U5594, U5596);
  and ginst4426 (U3770, U5598, U5599);
  and ginst4427 (U3771, U3770, U5597);
  and ginst4428 (U3772, U5600, U5601, U5603);
  and ginst4429 (U3773, U5605, U5606);
  and ginst4430 (U3774, U3773, U5604);
  and ginst4431 (U3775, U5607, U5608, U5610);
  and ginst4432 (U3776, U5612, U5613);
  and ginst4433 (U3777, U3776, U5611);
  and ginst4434 (U3778, U5614, U5615, U5617);
  and ginst4435 (U3779, U5619, U5620);
  and ginst4436 (U3780, U3779, U5618);
  and ginst4437 (U3781, U5621, U5622, U5624);
  and ginst4438 (U3782, U5626, U5627);
  and ginst4439 (U3783, U3782, U5625);
  and ginst4440 (U3784, U5628, U5629, U5631);
  and ginst4441 (U3785, U5633, U5634);
  and ginst4442 (U3786, U3785, U5632);
  and ginst4443 (U3787, U5635, U5636, U5638);
  and ginst4444 (U3788, U5640, U5641);
  and ginst4445 (U3789, U3788, U5639);
  and ginst4446 (U3790, U5642, U5643, U5645);
  and ginst4447 (U3791, U5647, U5648);
  and ginst4448 (U3792, U3791, U5646);
  and ginst4449 (U3793, U5650, U5652);
  and ginst4450 (U3794, U5654, U5655);
  and ginst4451 (U3795, U3794, U5653);
  and ginst4452 (U3796, U5657, U5659);
  and ginst4453 (U3797, U5661, U5662);
  and ginst4454 (U3798, U3797, U5660);
  and ginst4455 (U3799, U5664, U5666);
  and ginst4456 (U3800, U5668, U5669);
  and ginst4457 (U3801, U3800, U5667);
  and ginst4458 (U3802, U5671, U5673);
  and ginst4459 (U3803, U5675, U5676);
  and ginst4460 (U3804, U3803, U5674);
  and ginst4461 (U3805, U5678, U5680);
  and ginst4462 (U3806, U5682, U5683);
  and ginst4463 (U3807, U3806, U5681);
  and ginst4464 (U3808, U5685, U5687);
  and ginst4465 (U3809, U5689, U5690);
  and ginst4466 (U3810, U3809, U5688);
  and ginst4467 (U3811, U5692, U5694);
  and ginst4468 (U3812, U5696, U5697);
  and ginst4469 (U3813, U3812, U5695);
  and ginst4470 (U3814, U5699, U5701);
  and ginst4471 (U3815, U5703, U5704);
  and ginst4472 (U3816, U3815, U5702);
  and ginst4473 (U3817, U5706, U5708);
  and ginst4474 (U3818, U5710, U5711);
  and ginst4475 (U3819, U3818, U5709);
  and ginst4476 (U3820, U5713, U5715);
  and ginst4477 (U3821, U5717, U5718);
  and ginst4478 (U3822, U3821, U5716);
  and ginst4479 (U3823, U5720, U5722);
  and ginst4480 (U3824, U5724, U5725);
  and ginst4481 (U3825, U3824, U5723);
  and ginst4482 (U3826, U5727, U5729);
  and ginst4483 (U3827, U5731, U5732);
  and ginst4484 (U3828, U3827, U5730);
  and ginst4485 (U3829, U5734, U5736);
  and ginst4486 (U3830, U5738, U5739);
  and ginst4487 (U3831, U3830, U5737);
  and ginst4488 (U3832, U5741, U5743);
  and ginst4489 (U3833, U5745, U5746);
  and ginst4490 (U3834, U3833, U5744);
  and ginst4491 (U3835, U5748, U5750);
  and ginst4492 (U3836, U5752, U5753);
  and ginst4493 (U3837, U3836, U5751);
  and ginst4494 (U3838, U5755, U5757);
  and ginst4495 (U3839, U5759, U5760);
  and ginst4496 (U3840, U3839, U5758);
  and ginst4497 (U3841, U5762, U5764);
  and ginst4498 (U3842, U5766, U5767);
  and ginst4499 (U3843, U3842, U5765);
  and ginst4500 (U3844, U5769, U5771);
  and ginst4501 (U3845, U5773, U5774);
  and ginst4502 (U3846, U3845, U5772);
  and ginst4503 (U3847, U5776, U5778);
  and ginst4504 (U3848, U5780, U5781);
  and ginst4505 (U3849, U3848, U5779);
  and ginst4506 (U3850, U3249, U3270, U7482);
  and ginst4507 (U3851, U3395, U5782);
  and ginst4508 (U3852, STATEBS16_REG_SCAN_IN, STATE2_REG_1__SCAN_IN);
  and ginst4509 (U3853, U2368, U3271);
  and ginst4510 (U3854, STATE2_REG_0__SCAN_IN, U2449);
  and ginst4511 (U3855, U2368, U4196);
  and ginst4512 (U3856, U6093, U6094);
  and ginst4513 (U3857, U6096, U6097);
  and ginst4514 (U3858, U6099, U6100);
  and ginst4515 (U3859, U6102, U6103);
  and ginst4516 (U3860, U6105, U6106);
  and ginst4517 (U3861, U6108, U6109);
  and ginst4518 (U3862, U6111, U6112);
  and ginst4519 (U3863, U6114, U6115);
  and ginst4520 (U3864, U6117, U6118);
  and ginst4521 (U3865, U6120, U6121);
  and ginst4522 (U3866, U6123, U6124);
  and ginst4523 (U3867, U6126, U6127);
  and ginst4524 (U3868, U6129, U6130);
  and ginst4525 (U3869, U6132, U6133);
  and ginst4526 (U3870, U6135, U6136);
  and ginst4527 (U3871, U6138, U6139);
  and ginst4528 (U3872, U2605, U3378);
  and ginst4529 (U3873, STATE2_REG_0__SCAN_IN, U3258, U7482);
  and ginst4530 (U3874, U4159, U4387);
  and ginst4531 (U3875, U4229, U4232, U6350);
  nor ginst4532 (U3876, READY_N, STATEBS16_REG_SCAN_IN);
  and ginst4533 (U3877, U4174, U4482);
  and ginst4534 (U3878, U6359, U6360, U6361, U6362, U6363);
  and ginst4535 (U3879, U6367, U6368, U6369, U6370, U6371);
  and ginst4536 (U3880, U6375, U6376, U6377, U6378, U6379);
  and ginst4537 (U3881, U6383, U6384, U6385, U6386, U6387);
  and ginst4538 (U3882, U4215, U6388);
  and ginst4539 (U3883, U6392, U6393, U6394, U6395);
  and ginst4540 (U3884, U4215, U6396);
  and ginst4541 (U3885, U6399, U6400, U6401, U6402, U6403);
  and ginst4542 (U3886, U4215, U6404);
  and ginst4543 (U3887, U6407, U6409, U6410);
  and ginst4544 (U3888, U4215, U6411);
  and ginst4545 (U3889, U6414, U6416, U6417);
  and ginst4546 (U3890, U4215, U6418);
  and ginst4547 (U3891, U6421, U6423, U6424);
  and ginst4548 (U3892, U4215, U6425);
  and ginst4549 (U3893, U6428, U6430, U6431);
  and ginst4550 (U3894, U4215, U6432);
  and ginst4551 (U3895, U6435, U6437, U6438);
  and ginst4552 (U3896, U4215, U6439);
  and ginst4553 (U3897, U6442, U6444, U6445);
  and ginst4554 (U3898, U4215, U6446);
  and ginst4555 (U3899, U6449, U6451, U6452);
  and ginst4556 (U3900, U4215, U6453);
  and ginst4557 (U3901, U6456, U6458, U6459);
  and ginst4558 (U3902, U4215, U6460);
  and ginst4559 (U3903, U6463, U6465, U6466);
  and ginst4560 (U3904, U4215, U6467);
  and ginst4561 (U3905, U6470, U6472, U6473);
  and ginst4562 (U3906, U4215, U6474);
  and ginst4563 (U3907, U6477, U6479, U6480);
  and ginst4564 (U3908, U4215, U6482);
  and ginst4565 (U3909, U6484, U6486, U6487);
  and ginst4566 (U3910, U4215, U6489);
  and ginst4567 (U3911, U6491, U6493, U6494);
  and ginst4568 (U3912, U4215, U6496);
  and ginst4569 (U3913, U6498, U6500, U6501);
  and ginst4570 (U3914, U6503, U6505);
  and ginst4571 (U3915, U6507, U6508);
  and ginst4572 (U3916, U6510, U6512);
  and ginst4573 (U3917, U6514, U6515);
  and ginst4574 (U3918, U6517, U6519);
  and ginst4575 (U3919, U6521, U6522);
  and ginst4576 (U3920, U6524, U6526);
  and ginst4577 (U3921, U6528, U6529);
  and ginst4578 (U3922, U6531, U6533);
  and ginst4579 (U3923, U6535, U6536);
  and ginst4580 (U3924, U6538, U6540);
  and ginst4581 (U3925, U6542, U6543);
  and ginst4582 (U3926, U6545, U6547);
  and ginst4583 (U3927, U6549, U6550);
  and ginst4584 (U3928, U6552, U6554);
  and ginst4585 (U3929, U6556, U6557);
  and ginst4586 (U3930, U6559, U6561);
  and ginst4587 (U3931, U6563, U6564);
  and ginst4588 (U3932, U6566, U6568);
  and ginst4589 (U3933, U6570, U6571);
  and ginst4590 (U3934, U6573, U6575);
  and ginst4591 (U3935, U6577, U6578);
  and ginst4592 (U3936, U6580, U6582);
  and ginst4593 (U3937, U6584, U6585);
  nor ginst4594 (U3938, DATAWIDTH_REG_2__SCAN_IN, DATAWIDTH_REG_3__SCAN_IN, DATAWIDTH_REG_4__SCAN_IN, DATAWIDTH_REG_5__SCAN_IN);
  nor ginst4595 (U3939, DATAWIDTH_REG_6__SCAN_IN, DATAWIDTH_REG_7__SCAN_IN, DATAWIDTH_REG_8__SCAN_IN, DATAWIDTH_REG_9__SCAN_IN);
  and ginst4596 (U3940, U3938, U3939);
  nor ginst4597 (U3941, DATAWIDTH_REG_10__SCAN_IN, DATAWIDTH_REG_11__SCAN_IN, DATAWIDTH_REG_12__SCAN_IN, DATAWIDTH_REG_13__SCAN_IN);
  nor ginst4598 (U3942, DATAWIDTH_REG_14__SCAN_IN, DATAWIDTH_REG_15__SCAN_IN, DATAWIDTH_REG_16__SCAN_IN, DATAWIDTH_REG_17__SCAN_IN);
  and ginst4599 (U3943, U3941, U3942);
  nor ginst4600 (U3944, DATAWIDTH_REG_18__SCAN_IN, DATAWIDTH_REG_19__SCAN_IN, DATAWIDTH_REG_20__SCAN_IN, DATAWIDTH_REG_21__SCAN_IN);
  nor ginst4601 (U3945, DATAWIDTH_REG_22__SCAN_IN, DATAWIDTH_REG_23__SCAN_IN, DATAWIDTH_REG_24__SCAN_IN, DATAWIDTH_REG_25__SCAN_IN);
  and ginst4602 (U3946, U3944, U3945);
  nor ginst4603 (U3947, DATAWIDTH_REG_26__SCAN_IN, DATAWIDTH_REG_27__SCAN_IN);
  nor ginst4604 (U3948, DATAWIDTH_REG_28__SCAN_IN, DATAWIDTH_REG_29__SCAN_IN);
  nor ginst4605 (U3949, DATAWIDTH_REG_30__SCAN_IN, DATAWIDTH_REG_31__SCAN_IN);
  and ginst4606 (U3950, U3947, U3948, U3949, U6586);
  nor ginst4607 (U3951, DATAWIDTH_REG_0__SCAN_IN, DATAWIDTH_REG_1__SCAN_IN, REIP_REG_0__SCAN_IN);
  and ginst4608 (U3952, STATE2_REG_2__SCAN_IN, U3244);
  and ginst4609 (U3953, U3285, U6596);
  nor ginst4610 (U3954, READY_N, STATE2_REG_0__SCAN_IN);
  and ginst4611 (U3955, U3294, U3395, U6590);
  and ginst4612 (U3956, STATE2_REG_2__SCAN_IN, U3274);
  and ginst4613 (U3957, U4194, U4223);
  and ginst4614 (U3958, U6606, U6607, U6608, U6609);
  and ginst4615 (U3959, U6610, U6611, U6612, U6613);
  and ginst4616 (U3960, U6614, U6615, U6616, U6617);
  and ginst4617 (U3961, U6618, U6619, U6620, U6621);
  and ginst4618 (U3962, U6622, U6623, U6624, U6625);
  and ginst4619 (U3963, U6626, U6627, U6628, U6629);
  and ginst4620 (U3964, U6630, U6631, U6632, U6633);
  and ginst4621 (U3965, U6634, U6635, U6636, U6637);
  and ginst4622 (U3966, U6638, U6639, U6640, U6641);
  and ginst4623 (U3967, U6642, U6643, U6644, U6645);
  and ginst4624 (U3968, U6646, U6647, U6648, U6649);
  and ginst4625 (U3969, U6650, U6651, U6652, U6653);
  and ginst4626 (U3970, U6654, U6655, U6656, U6657);
  and ginst4627 (U3971, U6658, U6659, U6660, U6661);
  and ginst4628 (U3972, U6662, U6663, U6664, U6665);
  and ginst4629 (U3973, U6666, U6667, U6668, U7601);
  and ginst4630 (U3974, U6669, U6670, U6671, U6672);
  and ginst4631 (U3975, U6673, U6674, U6675, U6676);
  and ginst4632 (U3976, U6677, U6678, U6679, U6680);
  and ginst4633 (U3977, U6681, U6682, U6683, U6684);
  and ginst4634 (U3978, U6685, U6686, U6687, U6688);
  and ginst4635 (U3979, U6689, U6690, U6691, U6692);
  and ginst4636 (U3980, U6693, U6694, U6695, U6696);
  and ginst4637 (U3981, U6697, U6698, U6699, U6700);
  and ginst4638 (U3982, U6701, U6702, U6703, U6704);
  and ginst4639 (U3983, U6705, U6706, U6707, U6708);
  and ginst4640 (U3984, U6709, U6710, U6711, U6712);
  and ginst4641 (U3985, U6713, U6714, U6715, U6716);
  and ginst4642 (U3986, U6717, U6718, U6719, U6720);
  and ginst4643 (U3987, U6721, U6722, U6723, U6724);
  and ginst4644 (U3988, U6725, U6726, U6727, U6728);
  and ginst4645 (U3989, U6729, U6730, U6731, U6732);
  and ginst4646 (U3990, U6736, U6737);
  and ginst4647 (U3991, U6739, U6740);
  and ginst4648 (U3992, U6742, U6743);
  and ginst4649 (U3993, U6745, U6746);
  and ginst4650 (U3994, U3995, U6748);
  and ginst4651 (U3995, U6749, U6750);
  and ginst4652 (U3996, U6752, U6753);
  and ginst4653 (U3997, U6760, U6761, U6762);
  and ginst4654 (U3998, U6764, U6765);
  and ginst4655 (U3999, U6769, U6770, U6771);
  and ginst4656 (U4000, U6773, U6774, U6775);
  and ginst4657 (U4001, U6777, U6778, U6779);
  and ginst4658 (U4002, U6781, U6782, U6783);
  and ginst4659 (U4003, U6785, U6786, U6787);
  and ginst4660 (U4004, U6789, U6790, U6791);
  and ginst4661 (U4005, U6793, U6794, U6795);
  and ginst4662 (U4006, U6797, U6798, U6799);
  and ginst4663 (U4007, U6801, U6802, U6803);
  and ginst4664 (U4008, U6805, U6806, U6807);
  and ginst4665 (U4009, U6809, U6810);
  and ginst4666 (U4010, U6814, U6815, U6816);
  and ginst4667 (U4011, U6818, U6819, U6820);
  and ginst4668 (U4012, U6822, U6823, U6824);
  and ginst4669 (U4013, U6826, U6827, U6828);
  and ginst4670 (U4014, U6845, U6846);
  and ginst4671 (U4015, U6848, U6849);
  and ginst4672 (U4016, U3270, U6876, U7482);
  and ginst4673 (U4017, U6880, U6881, U6882, U6883);
  and ginst4674 (U4018, U6884, U6885, U6886, U6887);
  and ginst4675 (U4019, U6888, U6889, U6890, U6891);
  and ginst4676 (U4020, U6892, U6893, U6894, U6895);
  and ginst4677 (U4021, U6898, U6899, U6900, U6901);
  and ginst4678 (U4022, U6902, U6903, U6904, U6905);
  and ginst4679 (U4023, U6906, U6907, U6908, U6909);
  and ginst4680 (U4024, U6910, U6911, U6912, U6913);
  and ginst4681 (U4025, U6929, U6930, U6931, U6932);
  and ginst4682 (U4026, U6933, U6934, U6935, U6936);
  and ginst4683 (U4027, U6937, U6938, U6939, U6940);
  and ginst4684 (U4028, U6941, U6942, U6943, U6944);
  and ginst4685 (U4029, U6946, U6947, U6948, U6949);
  and ginst4686 (U4030, U6950, U6951, U6952, U6953);
  and ginst4687 (U4031, U6954, U6955, U6956, U6957);
  and ginst4688 (U4032, U6958, U6959, U6960, U6961);
  and ginst4689 (U4033, U6963, U6964, U6965, U6966);
  and ginst4690 (U4034, U6967, U6968, U6969, U6970);
  and ginst4691 (U4035, U6971, U6972, U6973, U6974);
  and ginst4692 (U4036, U6975, U6976, U6977, U6978);
  and ginst4693 (U4037, U6980, U6981, U6982, U6983);
  and ginst4694 (U4038, U6984, U6985, U6986, U6987);
  and ginst4695 (U4039, U6988, U6989, U6990, U6991);
  and ginst4696 (U4040, U6992, U6993, U6994, U7602);
  and ginst4697 (U4041, U6995, U6996, U6997, U6998);
  and ginst4698 (U4042, U6999, U7000, U7001, U7002);
  and ginst4699 (U4043, U7003, U7004, U7005, U7006);
  and ginst4700 (U4044, U7007, U7008, U7009, U7010);
  and ginst4701 (U4045, U7012, U7013, U7014, U7015);
  and ginst4702 (U4046, U7016, U7017, U7018, U7019);
  and ginst4703 (U4047, U7020, U7021, U7022, U7023);
  and ginst4704 (U4048, U7024, U7025, U7026, U7027);
  and ginst4705 (U4049, U3430, U7047);
  and ginst4706 (U4050, STATE2_REG_0__SCAN_IN, U7050);
  and ginst4707 (U4051, U7054, U7055, U7056, U7057);
  and ginst4708 (U4052, U7058, U7059, U7060, U7061);
  and ginst4709 (U4053, U7062, U7063, U7064, U7065);
  and ginst4710 (U4054, U7066, U7067, U7068, U7069);
  and ginst4711 (U4055, STATE2_REG_0__SCAN_IN, U4244);
  and ginst4712 (U4056, U4389, U4391, U4392, U4393);
  and ginst4713 (U4057, U4394, U4395, U4396);
  and ginst4714 (U4058, U4397, U4398, U4399, U4400);
  and ginst4715 (U4059, U4401, U4402);
  and ginst4716 (U4060, U3378, U4388);
  and ginst4717 (U4061, STATE2_REG_0__SCAN_IN, U3271);
  and ginst4718 (U4062, U7077, U7078);
  and ginst4719 (U4063, U3421, U7460, U7461);
  and ginst4720 (U4064, U7462, U7463, U7464);
  and ginst4721 (U4065, U2606, U4064, U7465);
  and ginst4722 (U4066, U7083, U7085);
  and ginst4723 (U4067, U7086, U7087, U7088, U7089);
  and ginst4724 (U4068, U7090, U7091, U7092, U7093);
  and ginst4725 (U4069, U7094, U7095, U7096, U7097);
  and ginst4726 (U4070, U7098, U7099, U7100, U7101);
  and ginst4727 (U4071, U7103, U7104, U7105, U7106);
  and ginst4728 (U4072, U7107, U7108, U7109, U7110);
  and ginst4729 (U4073, U7111, U7112, U7113, U7114);
  and ginst4730 (U4074, U7115, U7116, U7117, U7118);
  and ginst4731 (U4075, U7120, U7121, U7122, U7123);
  and ginst4732 (U4076, U7124, U7125, U7126, U7127);
  and ginst4733 (U4077, U7128, U7129, U7130, U7131);
  and ginst4734 (U4078, U7132, U7133);
  and ginst4735 (U4079, U4078, U7134, U7605);
  and ginst4736 (U4080, U7135, U7136, U7137, U7138);
  and ginst4737 (U4081, U7139, U7140, U7141, U7142);
  and ginst4738 (U4082, U7143, U7144, U7145, U7146);
  and ginst4739 (U4083, U7147, U7148, U7149, U7150);
  and ginst4740 (U4084, U7152, U7153, U7154, U7155);
  and ginst4741 (U4085, U7156, U7157, U7158, U7159);
  and ginst4742 (U4086, U7160, U7161, U7162, U7163);
  and ginst4743 (U4087, U7164, U7165, U7166, U7167);
  and ginst4744 (U4088, U7169, U7170, U7171, U7172);
  and ginst4745 (U4089, U7173, U7174, U7175, U7176);
  and ginst4746 (U4090, U7177, U7178, U7179, U7180);
  and ginst4747 (U4091, U7181, U7182, U7183, U7184);
  and ginst4748 (U4092, U7186, U7187, U7188, U7189);
  and ginst4749 (U4093, U7190, U7191, U7192, U7193);
  and ginst4750 (U4094, U7194, U7195, U7196, U7197);
  and ginst4751 (U4095, U7198, U7199, U7200, U7201);
  and ginst4752 (U4096, U3251, U7203);
  and ginst4753 (U4097, U7203, U7204);
  and ginst4754 (U4098, U3252, U7205);
  and ginst4755 (U4099, U3414, U7077);
  and ginst4756 (U4100, U7205, U7206);
  and ginst4757 (U4101, U4100, U7460, U7461);
  and ginst4758 (U4102, U3421, U4099, U4101, U7078);
  and ginst4759 (U4103, U7462, U7464, U7468, U7474);
  and ginst4760 (U4104, U7475, U7476, U7477, U7493);
  and ginst4761 (U4105, U7077, U7078);
  and ginst4762 (U4106, U3421, U7460, U7461);
  and ginst4763 (U4107, U7462, U7463, U7464);
  and ginst4764 (U4108, U2606, U2608, U4107, U7465);
  and ginst4765 (U4109, U7208, U7209, U7210, U7211);
  and ginst4766 (U4110, U7212, U7213, U7214, U7215);
  and ginst4767 (U4111, U7216, U7217, U7218, U7219);
  and ginst4768 (U4112, U7220, U7221, U7222, U7223);
  and ginst4769 (U4113, U7225, U7226, U7227, U7228);
  and ginst4770 (U4114, U7229, U7230, U7231, U7232);
  and ginst4771 (U4115, U7233, U7234, U7235, U7236);
  and ginst4772 (U4116, U7237, U7238, U7239, U7240);
  and ginst4773 (U4117, U7242, U7243, U7244, U7245);
  and ginst4774 (U4118, U7246, U7247, U7248, U7249);
  and ginst4775 (U4119, U7250, U7251, U7252, U7253);
  and ginst4776 (U4120, U7254, U7255, U7256, U7257);
  and ginst4777 (U4121, U7259, U7260, U7261, U7262);
  and ginst4778 (U4122, U7263, U7264, U7265, U7266);
  and ginst4779 (U4123, U7267, U7268, U7269, U7270);
  and ginst4780 (U4124, U7271, U7272, U7273, U7607);
  and ginst4781 (U4125, U7274, U7275, U7276, U7277);
  and ginst4782 (U4126, U7278, U7279, U7280, U7281);
  and ginst4783 (U4127, U7282, U7283, U7284, U7285);
  and ginst4784 (U4128, U7286, U7287, U7288, U7289);
  and ginst4785 (U4129, U7291, U7292, U7293, U7294);
  and ginst4786 (U4130, U7295, U7296, U7297, U7298);
  and ginst4787 (U4131, U7299, U7300, U7301, U7302);
  and ginst4788 (U4132, U7303, U7304, U7305, U7306);
  and ginst4789 (U4133, U7308, U7309, U7310, U7311);
  and ginst4790 (U4134, U7312, U7313, U7314, U7315);
  and ginst4791 (U4135, U7316, U7317, U7318, U7319);
  and ginst4792 (U4136, U7320, U7321, U7322, U7323);
  and ginst4793 (U4137, U7325, U7326, U7327, U7328);
  and ginst4794 (U4138, U7329, U7330, U7331, U7332);
  and ginst4795 (U4139, U7333, U7334, U7335, U7336);
  and ginst4796 (U4140, U7337, U7338, U7339, U7340);
  and ginst4797 (U4141, U3271, U3406);
  and ginst4798 (U4142, U3270, U3378);
  and ginst4799 (U4143, U4251, U7345, U7346);
  and ginst4800 (U4144, U4143, U7347);
  and ginst4801 (U4145, STATE2_REG_0__SCAN_IN, U2427);
  and ginst4802 (U4146, U4145, U7348);
  and ginst4803 (U4147, U3258, U4161);
  and ginst4804 (U4148, STATE2_REG_0__SCAN_IN, U4161);
  and ginst4805 (U4149, STATE2_REG_0__SCAN_IN, U7357);
  and ginst4806 (U4150, U2603, U7359);
  and ginst4807 (U4151, STATE2_REG_0__SCAN_IN, U7361);
  and ginst4808 (U4152, U2603, U7363);
  and ginst4809 (U4153, U7370, U7371);
  and ginst4810 (U4154, U3440, U7372);
  and ginst4811 (U4155, U7375, U7376, U7377);
  and ginst4812 (U4156, U7449, U7450);
  and ginst4813 (U4157, U7452, U7453);
  and ginst4814 (U4158, U7661, U7662);
  nand ginst4815 (U4159, U3557, U3558, U3559, U3560);
  nand ginst4816 (U4160, U3727, U5462);
  nand ginst4817 (U4161, U2607, U3561, U3562, U3563, U3564);
  not ginst4818 (U4162, INSTADDRPOINTER_REG_31__SCAN_IN);
  and ginst4819 (U4163, U7713, U7714);
  and ginst4820 (U4164, U7732, U7733);
  nand ginst4821 (U4165, U2368, U3272);
  nand ginst4822 (U4166, U3378, U4496);
  not ginst4823 (U4167, BS16_N);
  nand ginst4824 (U4168, U3955, U4216);
  nand ginst4825 (U4169, U3419, U4216);
  nand ginst4826 (U4170, U3726, U7685, U7686);
  nand ginst4827 (U4171, INSTQUEUERD_ADDR_REG_2__SCAN_IN, U3256);
  not ginst4828 (U4172, U3439);
  nand ginst4829 (U4173, HOLD, U3244);
  not ginst4830 (U4174, U3399);
  not ginst4831 (U4175, U3427);
  not ginst4832 (U4176, U3426);
  not ginst4833 (U4177, U3380);
  not ginst4834 (U4178, U3277);
  not ginst4835 (U4179, U3436);
  not ginst4836 (U4180, U3392);
  not ginst4837 (U4181, U3421);
  not ginst4838 (U4182, U3407);
  nand ginst4839 (U4183, U3258, U4253);
  nand ginst4840 (U4184, U2605, U4448);
  not ginst4841 (U4185, U3383);
  not ginst4842 (U4186, U3412);
  not ginst4843 (U4187, U3276);
  not ginst4844 (U4188, U3408);
  not ginst4845 (U4189, U3409);
  not ginst4846 (U4190, U3415);
  not ginst4847 (U4191, U3395);
  not ginst4848 (U4192, U3414);
  nand ginst4849 (U4193, U3873, U4177, U4185);
  not ginst4850 (U4194, U3405);
  not ginst4851 (U4195, U3430);
  not ginst4852 (U4196, U3269);
  not ginst4853 (U4197, U3294);
  not ginst4854 (U4198, U3377);
  not ginst4855 (U4199, U3433);
  not ginst4856 (U4200, U3434);
  not ginst4857 (U4201, U3435);
  not ginst4858 (U4202, U3387);
  not ginst4859 (U4203, U3275);
  not ginst4860 (U4204, U3279);
  nand ginst4861 (U4205, U2431, U3566);
  not ginst4862 (U4206, U3386);
  nand ginst4863 (U4207, U3258, U4437);
  not ginst4864 (U4208, U3420);
  not ginst4865 (U4209, U3236);
  not ginst4866 (U4210, U3413);
  not ginst4867 (U4211, U3411);
  not ginst4868 (U4212, U3287);
  not ginst4869 (U4213, LT_563_1260_U6);
  not ginst4870 (U4214, U3307);
  nand ginst4871 (U4215, U3418, U4243);
  nand ginst4872 (U4216, U4223, U7488);
  nand ginst4873 (U4217, U2362, U3259);
  nand ginst4874 (U4218, U2363, U4365);
  not ginst4875 (U4219, U3394);
  not ginst4876 (U4220, U3239);
  not ginst4877 (U4221, U3237);
  not ginst4878 (U4222, U3382);
  not ginst4879 (U4223, U3284);
  not ginst4880 (U4224, U3385);
  not ginst4881 (U4225, U4166);
  not ginst4882 (U4226, U3344);
  nand ginst4883 (U4227, U4465, U7369);
  nand ginst4884 (U4228, U3951, U4208);
  nand ginst4885 (U4229, U3572, U4249);
  nand ginst4886 (U4230, U2428, U3719);
  nand ginst4887 (U4231, U3245, U4352);
  nand ginst4888 (U4232, STATE2_REG_1__SCAN_IN, U2352, U3281);
  nand ginst4889 (U4233, U2428, U3390);
  nand ginst4890 (U4234, READY_N, STATE2_REG_0__SCAN_IN, U3250);
  not ginst4891 (U4235, U3381);
  nand ginst4892 (U4236, U2353, U2448, U2451, U3850);
  not ginst4893 (U4237, U3274);
  not ginst4894 (U4238, U3384);
  not ginst4895 (U4239, U3402);
  not ginst4896 (U4240, U3286);
  not ginst4897 (U4241, U3396);
  not ginst4898 (U4242, U3406);
  not ginst4899 (U4243, U3419);
  not ginst4900 (U4244, U3278);
  not ginst4901 (U4245, U3376);
  not ginst4902 (U4246, U3241);
  not ginst4903 (U4247, U3268);
  not ginst4904 (U4248, U3393);
  not ginst4905 (U4249, U3285);
  not ginst4906 (U4250, U3273);
  nand ginst4907 (U4251, U4224, U4387);
  not ginst4908 (U4252, U3398);
  not ginst4909 (U4253, U3440);
  not ginst4910 (U4254, U3397);
  nand ginst4911 (U4255, REIP_REG_31__SCAN_IN, U4221);
  nand ginst4912 (U4256, REIP_REG_30__SCAN_IN, U4220);
  nand ginst4913 (U4257, ADDRESS_REG_29__SCAN_IN, U3236);
  nand ginst4914 (U4258, REIP_REG_30__SCAN_IN, U4221);
  nand ginst4915 (U4259, REIP_REG_29__SCAN_IN, U4220);
  nand ginst4916 (U4260, ADDRESS_REG_28__SCAN_IN, U3236);
  nand ginst4917 (U4261, REIP_REG_29__SCAN_IN, U4221);
  nand ginst4918 (U4262, REIP_REG_28__SCAN_IN, U4220);
  nand ginst4919 (U4263, ADDRESS_REG_27__SCAN_IN, U3236);
  nand ginst4920 (U4264, REIP_REG_28__SCAN_IN, U4221);
  nand ginst4921 (U4265, REIP_REG_27__SCAN_IN, U4220);
  nand ginst4922 (U4266, ADDRESS_REG_26__SCAN_IN, U3236);
  nand ginst4923 (U4267, REIP_REG_27__SCAN_IN, U4221);
  nand ginst4924 (U4268, REIP_REG_26__SCAN_IN, U4220);
  nand ginst4925 (U4269, ADDRESS_REG_25__SCAN_IN, U3236);
  nand ginst4926 (U4270, REIP_REG_26__SCAN_IN, U4221);
  nand ginst4927 (U4271, REIP_REG_25__SCAN_IN, U4220);
  nand ginst4928 (U4272, ADDRESS_REG_24__SCAN_IN, U3236);
  nand ginst4929 (U4273, REIP_REG_25__SCAN_IN, U4221);
  nand ginst4930 (U4274, REIP_REG_24__SCAN_IN, U4220);
  nand ginst4931 (U4275, ADDRESS_REG_23__SCAN_IN, U3236);
  nand ginst4932 (U4276, REIP_REG_24__SCAN_IN, U4221);
  nand ginst4933 (U4277, REIP_REG_23__SCAN_IN, U4220);
  nand ginst4934 (U4278, ADDRESS_REG_22__SCAN_IN, U3236);
  nand ginst4935 (U4279, REIP_REG_23__SCAN_IN, U4221);
  nand ginst4936 (U4280, REIP_REG_22__SCAN_IN, U4220);
  nand ginst4937 (U4281, ADDRESS_REG_21__SCAN_IN, U3236);
  nand ginst4938 (U4282, REIP_REG_22__SCAN_IN, U4221);
  nand ginst4939 (U4283, REIP_REG_21__SCAN_IN, U4220);
  nand ginst4940 (U4284, ADDRESS_REG_20__SCAN_IN, U3236);
  nand ginst4941 (U4285, REIP_REG_21__SCAN_IN, U4221);
  nand ginst4942 (U4286, REIP_REG_20__SCAN_IN, U4220);
  nand ginst4943 (U4287, ADDRESS_REG_19__SCAN_IN, U3236);
  nand ginst4944 (U4288, REIP_REG_20__SCAN_IN, U4221);
  nand ginst4945 (U4289, REIP_REG_19__SCAN_IN, U4220);
  nand ginst4946 (U4290, ADDRESS_REG_18__SCAN_IN, U3236);
  nand ginst4947 (U4291, REIP_REG_19__SCAN_IN, U4221);
  nand ginst4948 (U4292, REIP_REG_18__SCAN_IN, U4220);
  nand ginst4949 (U4293, ADDRESS_REG_17__SCAN_IN, U3236);
  nand ginst4950 (U4294, REIP_REG_18__SCAN_IN, U4221);
  nand ginst4951 (U4295, REIP_REG_17__SCAN_IN, U4220);
  nand ginst4952 (U4296, ADDRESS_REG_16__SCAN_IN, U3236);
  nand ginst4953 (U4297, REIP_REG_17__SCAN_IN, U4221);
  nand ginst4954 (U4298, REIP_REG_16__SCAN_IN, U4220);
  nand ginst4955 (U4299, ADDRESS_REG_15__SCAN_IN, U3236);
  nand ginst4956 (U4300, REIP_REG_16__SCAN_IN, U4221);
  nand ginst4957 (U4301, REIP_REG_15__SCAN_IN, U4220);
  nand ginst4958 (U4302, ADDRESS_REG_14__SCAN_IN, U3236);
  nand ginst4959 (U4303, REIP_REG_15__SCAN_IN, U4221);
  nand ginst4960 (U4304, REIP_REG_14__SCAN_IN, U4220);
  nand ginst4961 (U4305, ADDRESS_REG_13__SCAN_IN, U3236);
  nand ginst4962 (U4306, REIP_REG_14__SCAN_IN, U4221);
  nand ginst4963 (U4307, REIP_REG_13__SCAN_IN, U4220);
  nand ginst4964 (U4308, ADDRESS_REG_12__SCAN_IN, U3236);
  nand ginst4965 (U4309, REIP_REG_13__SCAN_IN, U4221);
  nand ginst4966 (U4310, REIP_REG_12__SCAN_IN, U4220);
  nand ginst4967 (U4311, ADDRESS_REG_11__SCAN_IN, U3236);
  nand ginst4968 (U4312, REIP_REG_12__SCAN_IN, U4221);
  nand ginst4969 (U4313, REIP_REG_11__SCAN_IN, U4220);
  nand ginst4970 (U4314, ADDRESS_REG_10__SCAN_IN, U3236);
  nand ginst4971 (U4315, REIP_REG_11__SCAN_IN, U4221);
  nand ginst4972 (U4316, REIP_REG_10__SCAN_IN, U4220);
  nand ginst4973 (U4317, ADDRESS_REG_9__SCAN_IN, U3236);
  nand ginst4974 (U4318, REIP_REG_10__SCAN_IN, U4221);
  nand ginst4975 (U4319, REIP_REG_9__SCAN_IN, U4220);
  nand ginst4976 (U4320, ADDRESS_REG_8__SCAN_IN, U3236);
  nand ginst4977 (U4321, REIP_REG_9__SCAN_IN, U4221);
  nand ginst4978 (U4322, REIP_REG_8__SCAN_IN, U4220);
  nand ginst4979 (U4323, ADDRESS_REG_7__SCAN_IN, U3236);
  nand ginst4980 (U4324, REIP_REG_8__SCAN_IN, U4221);
  nand ginst4981 (U4325, REIP_REG_7__SCAN_IN, U4220);
  nand ginst4982 (U4326, ADDRESS_REG_6__SCAN_IN, U3236);
  nand ginst4983 (U4327, REIP_REG_7__SCAN_IN, U4221);
  nand ginst4984 (U4328, REIP_REG_6__SCAN_IN, U4220);
  nand ginst4985 (U4329, ADDRESS_REG_5__SCAN_IN, U3236);
  nand ginst4986 (U4330, REIP_REG_6__SCAN_IN, U4221);
  nand ginst4987 (U4331, REIP_REG_5__SCAN_IN, U4220);
  nand ginst4988 (U4332, ADDRESS_REG_4__SCAN_IN, U3236);
  nand ginst4989 (U4333, REIP_REG_5__SCAN_IN, U4221);
  nand ginst4990 (U4334, REIP_REG_4__SCAN_IN, U4220);
  nand ginst4991 (U4335, ADDRESS_REG_3__SCAN_IN, U3236);
  nand ginst4992 (U4336, REIP_REG_4__SCAN_IN, U4221);
  nand ginst4993 (U4337, REIP_REG_3__SCAN_IN, U4220);
  nand ginst4994 (U4338, ADDRESS_REG_2__SCAN_IN, U3236);
  nand ginst4995 (U4339, REIP_REG_3__SCAN_IN, U4221);
  nand ginst4996 (U4340, REIP_REG_2__SCAN_IN, U4220);
  nand ginst4997 (U4341, ADDRESS_REG_1__SCAN_IN, U3236);
  nand ginst4998 (U4342, REIP_REG_2__SCAN_IN, U4221);
  nand ginst4999 (U4343, REIP_REG_1__SCAN_IN, U4220);
  nand ginst5000 (U4344, ADDRESS_REG_0__SCAN_IN, U3236);
  not ginst5001 (U4345, U3247);
  nand ginst5002 (U4346, U3244, U4345);
  nand ginst5003 (U4347, NA_N, U4246);
  not ginst5004 (U4348, U3248);
  nand ginst5005 (U4349, U3244, U4348);
  or ginst5006 (U4350, NA_N, STATE_REG_0__SCAN_IN);
  nand ginst5007 (U4351, U4350, U7610, U7611);
  not ginst5008 (U4352, U3242);
  nand ginst5009 (U4353, HOLD, U3234, U4352);
  nand ginst5010 (U4354, U3248, U3481);
  nand ginst5011 (U4355, U4353, U4354);
  nand ginst5012 (U4356, STATE_REG_0__SCAN_IN, U4347, U4355);
  nand ginst5013 (U4357, STATE_REG_2__SCAN_IN, U4351);
  nand ginst5014 (U4358, READY_N, U4209);
  nand ginst5015 (U4359, U3484, U7613);
  nand ginst5016 (U4360, STATE_REG_2__SCAN_IN, U3247);
  nand ginst5017 (U4361, NA_N, U3245);
  nand ginst5018 (U4362, U4360, U4361);
  nand ginst5019 (U4363, U3235, U4362);
  nand ginst5020 (U4364, U3242, U4167);
  not ginst5021 (U4365, U3267);
  not ginst5022 (U4366, U3256);
  not ginst5023 (U4367, U3431);
  not ginst5024 (U4368, U3255);
  not ginst5025 (U4369, U3261);
  not ginst5026 (U4370, U3254);
  nand ginst5027 (U4371, INSTQUEUE_REG_7__3__SCAN_IN, U4370);
  nand ginst5028 (U4372, INSTQUEUE_REG_0__3__SCAN_IN, U2472);
  nand ginst5029 (U4373, INSTQUEUE_REG_1__3__SCAN_IN, U2471);
  nand ginst5030 (U4374, INSTQUEUE_REG_2__3__SCAN_IN, U2470);
  nand ginst5031 (U4375, INSTQUEUE_REG_3__3__SCAN_IN, U2468);
  nand ginst5032 (U4376, INSTQUEUE_REG_4__3__SCAN_IN, U2467);
  nand ginst5033 (U4377, INSTQUEUE_REG_5__3__SCAN_IN, U2466);
  nand ginst5034 (U4378, INSTQUEUE_REG_6__3__SCAN_IN, U2465);
  nand ginst5035 (U4379, INSTQUEUE_REG_8__3__SCAN_IN, U2464);
  nand ginst5036 (U4380, INSTQUEUE_REG_9__3__SCAN_IN, U2463);
  nand ginst5037 (U4381, INSTQUEUE_REG_10__3__SCAN_IN, U2461);
  nand ginst5038 (U4382, INSTQUEUE_REG_11__3__SCAN_IN, U2459);
  nand ginst5039 (U4383, INSTQUEUE_REG_12__3__SCAN_IN, U2458);
  nand ginst5040 (U4384, INSTQUEUE_REG_13__3__SCAN_IN, U2457);
  nand ginst5041 (U4385, INSTQUEUE_REG_14__3__SCAN_IN, U2455);
  nand ginst5042 (U4386, INSTQUEUE_REG_15__3__SCAN_IN, U2453);
  not ginst5043 (U4387, U3270);
  not ginst5044 (U4388, U3265);
  nand ginst5045 (U4389, INSTQUEUE_REG_7__5__SCAN_IN, INSTQUEUERD_ADDR_REG_2__SCAN_IN, INSTQUEUERD_ADDR_REG_1__SCAN_IN, INSTQUEUERD_ADDR_REG_0__SCAN_IN, U3257);
  nand ginst5046 (U4390, INSTQUEUE_REG_0__5__SCAN_IN, U3257, U4368);
  nand ginst5047 (U4391, INSTQUEUE_REG_1__5__SCAN_IN, INSTQUEUERD_ADDR_REG_0__SCAN_IN, U2469, U3252);
  nand ginst5048 (U4392, INSTQUEUE_REG_2__5__SCAN_IN, INSTQUEUERD_ADDR_REG_1__SCAN_IN, U2469, U3253);
  nand ginst5049 (U4393, INSTQUEUE_REG_4__5__SCAN_IN, INSTQUEUERD_ADDR_REG_2__SCAN_IN, U3257, U4366);
  nand ginst5050 (U4394, INSTQUEUERD_ADDR_REG_2__SCAN_IN, U3508, U3509);
  nand ginst5051 (U4395, INSTQUEUERD_ADDR_REG_2__SCAN_IN, U3510, U3511);
  nand ginst5052 (U4396, U3512, U4368);
  nand ginst5053 (U4397, INSTQUEUERD_ADDR_REG_1__SCAN_IN, U3513, U3514);
  nand ginst5054 (U4398, INSTQUEUE_REG_11__5__SCAN_IN, INSTQUEUERD_ADDR_REG_3__SCAN_IN, INSTQUEUERD_ADDR_REG_1__SCAN_IN, INSTQUEUERD_ADDR_REG_0__SCAN_IN, U3251);
  nand ginst5055 (U4399, INSTQUEUERD_ADDR_REG_2__SCAN_IN, U3515, U4366);
  nand ginst5056 (U4400, INSTQUEUE_REG_13__5__SCAN_IN, INSTQUEUERD_ADDR_REG_3__SCAN_IN, INSTQUEUERD_ADDR_REG_2__SCAN_IN, INSTQUEUERD_ADDR_REG_0__SCAN_IN, U3252);
  nand ginst5057 (U4401, INSTQUEUE_REG_14__5__SCAN_IN, INSTQUEUERD_ADDR_REG_3__SCAN_IN, INSTQUEUERD_ADDR_REG_2__SCAN_IN, INSTQUEUERD_ADDR_REG_1__SCAN_IN, U3253);
  nand ginst5058 (U4402, INSTQUEUE_REG_15__5__SCAN_IN, INSTQUEUERD_ADDR_REG_3__SCAN_IN, INSTQUEUERD_ADDR_REG_2__SCAN_IN, INSTQUEUERD_ADDR_REG_1__SCAN_IN, INSTQUEUERD_ADDR_REG_0__SCAN_IN);
  not ginst5059 (U4403, U4161);
  nand ginst5060 (U4404, INSTQUEUE_REG_7__2__SCAN_IN, U4370);
  nand ginst5061 (U4405, INSTQUEUE_REG_0__2__SCAN_IN, U2472);
  nand ginst5062 (U4406, INSTQUEUE_REG_1__2__SCAN_IN, U2471);
  nand ginst5063 (U4407, INSTQUEUE_REG_2__2__SCAN_IN, U2470);
  nand ginst5064 (U4408, INSTQUEUE_REG_3__2__SCAN_IN, U2468);
  nand ginst5065 (U4409, INSTQUEUE_REG_4__2__SCAN_IN, U2467);
  nand ginst5066 (U4410, INSTQUEUE_REG_5__2__SCAN_IN, U2466);
  nand ginst5067 (U4411, INSTQUEUE_REG_6__2__SCAN_IN, U2465);
  nand ginst5068 (U4412, INSTQUEUE_REG_8__2__SCAN_IN, U2464);
  nand ginst5069 (U4413, INSTQUEUE_REG_9__2__SCAN_IN, U2463);
  nand ginst5070 (U4414, INSTQUEUE_REG_10__2__SCAN_IN, U2461);
  nand ginst5071 (U4415, INSTQUEUE_REG_11__2__SCAN_IN, U2459);
  nand ginst5072 (U4416, INSTQUEUE_REG_12__2__SCAN_IN, U2458);
  nand ginst5073 (U4417, INSTQUEUE_REG_13__2__SCAN_IN, U2457);
  nand ginst5074 (U4418, INSTQUEUE_REG_14__2__SCAN_IN, U2455);
  nand ginst5075 (U4419, INSTQUEUE_REG_15__2__SCAN_IN, U2453);
  not ginst5076 (U4420, U4159);
  nand ginst5077 (U4421, INSTQUEUE_REG_7__7__SCAN_IN, U4370);
  nand ginst5078 (U4422, INSTQUEUE_REG_0__7__SCAN_IN, U2472);
  nand ginst5079 (U4423, INSTQUEUE_REG_1__7__SCAN_IN, U2471);
  nand ginst5080 (U4424, INSTQUEUE_REG_2__7__SCAN_IN, U2470);
  nand ginst5081 (U4425, INSTQUEUE_REG_3__7__SCAN_IN, U2468);
  nand ginst5082 (U4426, INSTQUEUE_REG_4__7__SCAN_IN, U2467);
  nand ginst5083 (U4427, INSTQUEUE_REG_5__7__SCAN_IN, U2466);
  nand ginst5084 (U4428, INSTQUEUE_REG_6__7__SCAN_IN, U2465);
  nand ginst5085 (U4429, INSTQUEUE_REG_8__7__SCAN_IN, U2464);
  nand ginst5086 (U4430, INSTQUEUE_REG_9__7__SCAN_IN, U2463);
  nand ginst5087 (U4431, INSTQUEUE_REG_10__7__SCAN_IN, U2461);
  nand ginst5088 (U4432, INSTQUEUE_REG_11__7__SCAN_IN, U2459);
  nand ginst5089 (U4433, INSTQUEUE_REG_12__7__SCAN_IN, U2458);
  nand ginst5090 (U4434, INSTQUEUE_REG_13__7__SCAN_IN, U2457);
  nand ginst5091 (U4435, INSTQUEUE_REG_14__7__SCAN_IN, U2455);
  nand ginst5092 (U4436, INSTQUEUE_REG_15__7__SCAN_IN, U2453);
  not ginst5093 (U4437, U3378);
  nand ginst5094 (U4438, INSTQUEUE_REG_7__6__SCAN_IN, U3486, U4369);
  nand ginst5095 (U4439, INSTQUEUE_REG_1__6__SCAN_IN, U2456, U2469);
  nand ginst5096 (U4440, INSTQUEUE_REG_2__6__SCAN_IN, U2454, U2469);
  nand ginst5097 (U4441, INSTQUEUE_REG_4__6__SCAN_IN, U4366, U4369);
  nand ginst5098 (U4442, INSTQUEUE_REG_5__6__SCAN_IN, U2456, U4369);
  nand ginst5099 (U4443, INSTQUEUE_REG_6__6__SCAN_IN, U2454, U4369);
  nand ginst5100 (U4444, INSTQUEUE_REG_12__6__SCAN_IN, U3495, U4366);
  nand ginst5101 (U4445, INSTQUEUE_REG_13__6__SCAN_IN, U2456, U3495);
  nand ginst5102 (U4446, INSTQUEUE_REG_14__6__SCAN_IN, U2454, U3495);
  nand ginst5103 (U4447, INSTQUEUE_REG_15__6__SCAN_IN, U3486, U3495);
  not ginst5104 (U4448, U3264);
  nand ginst5105 (U4449, INSTQUEUE_REG_7__1__SCAN_IN, U4370);
  nand ginst5106 (U4450, INSTQUEUE_REG_0__1__SCAN_IN, U2472);
  nand ginst5107 (U4451, INSTQUEUE_REG_1__1__SCAN_IN, U2471);
  nand ginst5108 (U4452, INSTQUEUE_REG_2__1__SCAN_IN, U2470);
  nand ginst5109 (U4453, INSTQUEUE_REG_3__1__SCAN_IN, U2468);
  nand ginst5110 (U4454, INSTQUEUE_REG_4__1__SCAN_IN, U2467);
  nand ginst5111 (U4455, INSTQUEUE_REG_5__1__SCAN_IN, U2466);
  nand ginst5112 (U4456, INSTQUEUE_REG_6__1__SCAN_IN, U2465);
  nand ginst5113 (U4457, INSTQUEUE_REG_8__1__SCAN_IN, U2464);
  nand ginst5114 (U4458, INSTQUEUE_REG_9__1__SCAN_IN, U2463);
  nand ginst5115 (U4459, INSTQUEUE_REG_10__1__SCAN_IN, U2461);
  nand ginst5116 (U4460, INSTQUEUE_REG_11__1__SCAN_IN, U2459);
  nand ginst5117 (U4461, INSTQUEUE_REG_12__1__SCAN_IN, U2458);
  nand ginst5118 (U4462, INSTQUEUE_REG_13__1__SCAN_IN, U2457);
  nand ginst5119 (U4463, INSTQUEUE_REG_14__1__SCAN_IN, U2455);
  nand ginst5120 (U4464, INSTQUEUE_REG_15__1__SCAN_IN, U2453);
  not ginst5121 (U4465, U3258);
  nand ginst5122 (U4466, INSTQUEUE_REG_7__0__SCAN_IN, U4370);
  nand ginst5123 (U4467, INSTQUEUE_REG_0__0__SCAN_IN, U2472);
  nand ginst5124 (U4468, INSTQUEUE_REG_1__0__SCAN_IN, U2471);
  nand ginst5125 (U4469, INSTQUEUE_REG_2__0__SCAN_IN, U2470);
  nand ginst5126 (U4470, INSTQUEUE_REG_3__0__SCAN_IN, U2468);
  nand ginst5127 (U4471, INSTQUEUE_REG_4__0__SCAN_IN, U2467);
  nand ginst5128 (U4472, INSTQUEUE_REG_5__0__SCAN_IN, U2466);
  nand ginst5129 (U4473, INSTQUEUE_REG_6__0__SCAN_IN, U2465);
  nand ginst5130 (U4474, INSTQUEUE_REG_8__0__SCAN_IN, U2464);
  nand ginst5131 (U4475, INSTQUEUE_REG_9__0__SCAN_IN, U2463);
  nand ginst5132 (U4476, INSTQUEUE_REG_10__0__SCAN_IN, U2461);
  nand ginst5133 (U4477, INSTQUEUE_REG_11__0__SCAN_IN, U2459);
  nand ginst5134 (U4478, INSTQUEUE_REG_12__0__SCAN_IN, U2458);
  nand ginst5135 (U4479, INSTQUEUE_REG_13__0__SCAN_IN, U2457);
  nand ginst5136 (U4480, INSTQUEUE_REG_14__0__SCAN_IN, U2455);
  nand ginst5137 (U4481, INSTQUEUE_REG_15__0__SCAN_IN, U2453);
  not ginst5138 (U4482, U3271);
  nand ginst5139 (U4483, STATE_REG_2__SCAN_IN, U3235);
  nand ginst5140 (U4484, U3241, U4483);
  not ginst5141 (U4485, U3259);
  nand ginst5142 (U4486, U3375, U4465);
  not ginst5143 (U4487, U3424);
  nand ginst5144 (U4488, U3259, U3274, U3377);
  nand ginst5145 (U4489, U3244, U4488);
  not ginst5146 (U4490, U3272);
  nand ginst5147 (U4491, U4161, U4448);
  nand ginst5148 (U4492, U3273, U4184);
  nand ginst5149 (U4493, U3567, U4492);
  nand ginst5150 (U4494, U3568, U4493);
  nand ginst5151 (U4495, U3375, U4203);
  nand ginst5152 (U4496, U4495, U7669, U7670);
  nand ginst5153 (U4497, U2448, U4250);
  or ginst5154 (U4498, MORE_REG_SCAN_IN, FLUSH_REG_SCAN_IN);
  not ginst5155 (U4499, U3280);
  nand ginst5156 (U4500, U3249, U4499);
  nand ginst5157 (U4501, READY_N, STATE2_REG_1__SCAN_IN);
  not ginst5158 (U4502, U3282);
  nand ginst5159 (U4503, STATE2_REG_1__SCAN_IN, U7675, U7676);
  nand ginst5160 (U4504, STATE2_REG_2__SCAN_IN, U3282);
  nand ginst5161 (U4505, U4234, U7592);
  nand ginst5162 (U4506, U3571, U4502);
  nand ginst5163 (U4507, STATE2_REG_1__SCAN_IN, U4505);
  nand ginst5164 (U4508, U2368, U7592);
  nand ginst5165 (U4509, U4240, U4249);
  nand ginst5166 (U4510, U4233, U7592);
  nand ginst5167 (U4511, U2368, U3280);
  not ginst5168 (U4512, U3312);
  not ginst5169 (U4513, U3318);
  not ginst5170 (U4514, U3319);
  not ginst5171 (U4515, U3301);
  not ginst5172 (U4516, U3300);
  not ginst5173 (U4517, U3329);
  nand ginst5174 (U4518, R2144_U8, U3300);
  not ginst5175 (U4519, U3345);
  not ginst5176 (U4520, U3302);
  not ginst5177 (U4521, U3292);
  not ginst5178 (U4522, U3293);
  nand ginst5179 (U4523, U2438, U2442);
  not ginst5180 (U4524, U3308);
  not ginst5181 (U4525, U3343);
  not ginst5182 (U4526, U3327);
  nand ginst5183 (U4527, INSTQUEUEWR_ADDR_REG_3__SCAN_IN, U3292);
  not ginst5184 (U4528, U3347);
  not ginst5185 (U4529, U3316);
  not ginst5186 (U4530, U3310);
  not ginst5187 (U4531, U3222);
  nand ginst5188 (U4532, U2432, U2436);
  not ginst5189 (U4533, U3309);
  nand ginst5190 (U4534, STATE2_REG_1__SCAN_IN, U3250);
  nand ginst5191 (U4535, U3284, U3286, U4534);
  nand ginst5192 (U4536, U2476, U4516);
  nand ginst5193 (U4537, U2358, U2480);
  nand ginst5194 (U4538, U3307, U4537);
  nand ginst5195 (U4539, U4524, U4538);
  nand ginst5196 (U4540, STATE2_REG_3__SCAN_IN, U3293);
  nand ginst5197 (U4541, STATE2_REG_2__SCAN_IN, U4533);
  nand ginst5198 (U4542, U3575, U4539);
  nand ginst5199 (U4543, U2388, U2480);
  nand ginst5200 (U4544, U3307, U4543);
  nand ginst5201 (U4545, U3308, U4544);
  nand ginst5202 (U4546, STATE2_REG_2__SCAN_IN, U3309);
  nand ginst5203 (U4547, U4545, U4546);
  nand ginst5204 (U4548, U2415, U4522);
  nand ginst5205 (U4549, U2413, U2477);
  nand ginst5206 (U4550, U2412, U4520);
  nand ginst5207 (U4551, U2397, U4547);
  nand ginst5208 (U4552, INSTQUEUE_REG_15__7__SCAN_IN, U4542);
  nand ginst5209 (U4553, U2416, U4522);
  nand ginst5210 (U4554, U2411, U2477);
  nand ginst5211 (U4555, U2410, U4520);
  nand ginst5212 (U4556, U2396, U4547);
  nand ginst5213 (U4557, INSTQUEUE_REG_15__6__SCAN_IN, U4542);
  nand ginst5214 (U4558, U2420, U4522);
  nand ginst5215 (U4559, U2409, U2477);
  nand ginst5216 (U4560, U2408, U4520);
  nand ginst5217 (U4561, U2395, U4547);
  nand ginst5218 (U4562, INSTQUEUE_REG_15__5__SCAN_IN, U4542);
  nand ginst5219 (U4563, U2419, U4522);
  nand ginst5220 (U4564, U2407, U2477);
  nand ginst5221 (U4565, U2406, U4520);
  nand ginst5222 (U4566, U2394, U4547);
  nand ginst5223 (U4567, INSTQUEUE_REG_15__4__SCAN_IN, U4542);
  nand ginst5224 (U4568, U2418, U4522);
  nand ginst5225 (U4569, U2405, U2477);
  nand ginst5226 (U4570, U2404, U4520);
  nand ginst5227 (U4571, U2393, U4547);
  nand ginst5228 (U4572, INSTQUEUE_REG_15__3__SCAN_IN, U4542);
  nand ginst5229 (U4573, U2421, U4522);
  nand ginst5230 (U4574, U2403, U2477);
  nand ginst5231 (U4575, U2402, U4520);
  nand ginst5232 (U4576, U2392, U4547);
  nand ginst5233 (U4577, INSTQUEUE_REG_15__2__SCAN_IN, U4542);
  nand ginst5234 (U4578, U2414, U4522);
  nand ginst5235 (U4579, U2401, U2477);
  nand ginst5236 (U4580, U2400, U4520);
  nand ginst5237 (U4581, U2391, U4547);
  nand ginst5238 (U4582, INSTQUEUE_REG_15__1__SCAN_IN, U4542);
  nand ginst5239 (U4583, U2417, U4522);
  nand ginst5240 (U4584, U2399, U2477);
  nand ginst5241 (U4585, U2398, U4520);
  nand ginst5242 (U4586, U2390, U4547);
  nand ginst5243 (U4587, INSTQUEUE_REG_15__0__SCAN_IN, U4542);
  not ginst5244 (U4588, U3313);
  not ginst5245 (U4589, U3314);
  not ginst5246 (U4590, U3311);
  nand ginst5247 (U4591, U2438, U2443);
  not ginst5248 (U4592, U3315);
  not ginst5249 (U4593, U3223);
  nand ginst5250 (U4594, U2476, U4512);
  nand ginst5251 (U4595, U2358, U2482);
  nand ginst5252 (U4596, U3307, U4595);
  nand ginst5253 (U4597, U4592, U4596);
  nand ginst5254 (U4598, STATE2_REG_3__SCAN_IN, U3311);
  nand ginst5255 (U4599, STATE2_REG_2__SCAN_IN, U3223);
  nand ginst5256 (U4600, U3584, U4597);
  nand ginst5257 (U4601, U2388, U2482);
  nand ginst5258 (U4602, U3307, U4601);
  nand ginst5259 (U4603, U3315, U4602);
  nand ginst5260 (U4604, STATE2_REG_2__SCAN_IN, U4593);
  nand ginst5261 (U4605, U4603, U4604);
  nand ginst5262 (U4606, U2415, U4590);
  nand ginst5263 (U4607, U2413, U2481);
  nand ginst5264 (U4608, U2412, U4589);
  nand ginst5265 (U4609, U2397, U4605);
  nand ginst5266 (U4610, INSTQUEUE_REG_14__7__SCAN_IN, U4600);
  nand ginst5267 (U4611, U2416, U4590);
  nand ginst5268 (U4612, U2411, U2481);
  nand ginst5269 (U4613, U2410, U4589);
  nand ginst5270 (U4614, U2396, U4605);
  nand ginst5271 (U4615, INSTQUEUE_REG_14__6__SCAN_IN, U4600);
  nand ginst5272 (U4616, U2420, U4590);
  nand ginst5273 (U4617, U2409, U2481);
  nand ginst5274 (U4618, U2408, U4589);
  nand ginst5275 (U4619, U2395, U4605);
  nand ginst5276 (U4620, INSTQUEUE_REG_14__5__SCAN_IN, U4600);
  nand ginst5277 (U4621, U2419, U4590);
  nand ginst5278 (U4622, U2407, U2481);
  nand ginst5279 (U4623, U2406, U4589);
  nand ginst5280 (U4624, U2394, U4605);
  nand ginst5281 (U4625, INSTQUEUE_REG_14__4__SCAN_IN, U4600);
  nand ginst5282 (U4626, U2418, U4590);
  nand ginst5283 (U4627, U2405, U2481);
  nand ginst5284 (U4628, U2404, U4589);
  nand ginst5285 (U4629, U2393, U4605);
  nand ginst5286 (U4630, INSTQUEUE_REG_14__3__SCAN_IN, U4600);
  nand ginst5287 (U4631, U2421, U4590);
  nand ginst5288 (U4632, U2403, U2481);
  nand ginst5289 (U4633, U2402, U4589);
  nand ginst5290 (U4634, U2392, U4605);
  nand ginst5291 (U4635, INSTQUEUE_REG_14__2__SCAN_IN, U4600);
  nand ginst5292 (U4636, U2414, U4590);
  nand ginst5293 (U4637, U2401, U2481);
  nand ginst5294 (U4638, U2400, U4589);
  nand ginst5295 (U4639, U2391, U4605);
  nand ginst5296 (U4640, INSTQUEUE_REG_14__1__SCAN_IN, U4600);
  nand ginst5297 (U4641, U2417, U4590);
  nand ginst5298 (U4642, U2399, U2481);
  nand ginst5299 (U4643, U2398, U4589);
  nand ginst5300 (U4644, U2390, U4605);
  nand ginst5301 (U4645, INSTQUEUE_REG_14__0__SCAN_IN, U4600);
  not ginst5302 (U4646, U3320);
  not ginst5303 (U4647, U3321);
  not ginst5304 (U4648, U3317);
  nand ginst5305 (U4649, U2438, U2444);
  not ginst5306 (U4650, U3322);
  nand ginst5307 (U4651, U2432, U2437);
  not ginst5308 (U4652, U3323);
  nand ginst5309 (U4653, U2476, U4513);
  nand ginst5310 (U4654, U2358, U2484);
  nand ginst5311 (U4655, U3307, U4654);
  nand ginst5312 (U4656, U4650, U4655);
  nand ginst5313 (U4657, STATE2_REG_3__SCAN_IN, U3317);
  nand ginst5314 (U4658, STATE2_REG_2__SCAN_IN, U4652);
  nand ginst5315 (U4659, U3593, U4656);
  nand ginst5316 (U4660, U2388, U2484);
  nand ginst5317 (U4661, U3307, U4660);
  nand ginst5318 (U4662, U3322, U4661);
  nand ginst5319 (U4663, STATE2_REG_2__SCAN_IN, U3323);
  nand ginst5320 (U4664, U4662, U4663);
  nand ginst5321 (U4665, U2415, U4648);
  nand ginst5322 (U4666, U2413, U2483);
  nand ginst5323 (U4667, U2412, U4647);
  nand ginst5324 (U4668, U2397, U4664);
  nand ginst5325 (U4669, INSTQUEUE_REG_13__7__SCAN_IN, U4659);
  nand ginst5326 (U4670, U2416, U4648);
  nand ginst5327 (U4671, U2411, U2483);
  nand ginst5328 (U4672, U2410, U4647);
  nand ginst5329 (U4673, U2396, U4664);
  nand ginst5330 (U4674, INSTQUEUE_REG_13__6__SCAN_IN, U4659);
  nand ginst5331 (U4675, U2420, U4648);
  nand ginst5332 (U4676, U2409, U2483);
  nand ginst5333 (U4677, U2408, U4647);
  nand ginst5334 (U4678, U2395, U4664);
  nand ginst5335 (U4679, INSTQUEUE_REG_13__5__SCAN_IN, U4659);
  nand ginst5336 (U4680, U2419, U4648);
  nand ginst5337 (U4681, U2407, U2483);
  nand ginst5338 (U4682, U2406, U4647);
  nand ginst5339 (U4683, U2394, U4664);
  nand ginst5340 (U4684, INSTQUEUE_REG_13__4__SCAN_IN, U4659);
  nand ginst5341 (U4685, U2418, U4648);
  nand ginst5342 (U4686, U2405, U2483);
  nand ginst5343 (U4687, U2404, U4647);
  nand ginst5344 (U4688, U2393, U4664);
  nand ginst5345 (U4689, INSTQUEUE_REG_13__3__SCAN_IN, U4659);
  nand ginst5346 (U4690, U2421, U4648);
  nand ginst5347 (U4691, U2403, U2483);
  nand ginst5348 (U4692, U2402, U4647);
  nand ginst5349 (U4693, U2392, U4664);
  nand ginst5350 (U4694, INSTQUEUE_REG_13__2__SCAN_IN, U4659);
  nand ginst5351 (U4695, U2414, U4648);
  nand ginst5352 (U4696, U2401, U2483);
  nand ginst5353 (U4697, U2400, U4647);
  nand ginst5354 (U4698, U2391, U4664);
  nand ginst5355 (U4699, INSTQUEUE_REG_13__1__SCAN_IN, U4659);
  nand ginst5356 (U4700, U2417, U4648);
  nand ginst5357 (U4701, U2399, U2483);
  nand ginst5358 (U4702, U2398, U4647);
  nand ginst5359 (U4703, U2390, U4664);
  nand ginst5360 (U4704, INSTQUEUE_REG_13__0__SCAN_IN, U4659);
  not ginst5361 (U4705, U3325);
  not ginst5362 (U4706, U3324);
  nand ginst5363 (U4707, U2438, U2445);
  not ginst5364 (U4708, U3326);
  not ginst5365 (U4709, U3224);
  nand ginst5366 (U4710, U2476, U2486);
  nand ginst5367 (U4711, U2358, U2489);
  nand ginst5368 (U4712, U3307, U4711);
  nand ginst5369 (U4713, U4708, U4712);
  nand ginst5370 (U4714, STATE2_REG_3__SCAN_IN, U3324);
  nand ginst5371 (U4715, STATE2_REG_2__SCAN_IN, U3224);
  nand ginst5372 (U4716, U3602, U4713);
  nand ginst5373 (U4717, U2388, U2489);
  nand ginst5374 (U4718, U3307, U4717);
  nand ginst5375 (U4719, U3326, U4718);
  nand ginst5376 (U4720, STATE2_REG_2__SCAN_IN, U4709);
  nand ginst5377 (U4721, U4719, U4720);
  nand ginst5378 (U4722, U2415, U4706);
  nand ginst5379 (U4723, U2413, U2487);
  nand ginst5380 (U4724, U2412, U4705);
  nand ginst5381 (U4725, U2397, U4721);
  nand ginst5382 (U4726, INSTQUEUE_REG_12__7__SCAN_IN, U4716);
  nand ginst5383 (U4727, U2416, U4706);
  nand ginst5384 (U4728, U2411, U2487);
  nand ginst5385 (U4729, U2410, U4705);
  nand ginst5386 (U4730, U2396, U4721);
  nand ginst5387 (U4731, INSTQUEUE_REG_12__6__SCAN_IN, U4716);
  nand ginst5388 (U4732, U2420, U4706);
  nand ginst5389 (U4733, U2409, U2487);
  nand ginst5390 (U4734, U2408, U4705);
  nand ginst5391 (U4735, U2395, U4721);
  nand ginst5392 (U4736, INSTQUEUE_REG_12__5__SCAN_IN, U4716);
  nand ginst5393 (U4737, U2419, U4706);
  nand ginst5394 (U4738, U2407, U2487);
  nand ginst5395 (U4739, U2406, U4705);
  nand ginst5396 (U4740, U2394, U4721);
  nand ginst5397 (U4741, INSTQUEUE_REG_12__4__SCAN_IN, U4716);
  nand ginst5398 (U4742, U2418, U4706);
  nand ginst5399 (U4743, U2405, U2487);
  nand ginst5400 (U4744, U2404, U4705);
  nand ginst5401 (U4745, U2393, U4721);
  nand ginst5402 (U4746, INSTQUEUE_REG_12__3__SCAN_IN, U4716);
  nand ginst5403 (U4747, U2421, U4706);
  nand ginst5404 (U4748, U2403, U2487);
  nand ginst5405 (U4749, U2402, U4705);
  nand ginst5406 (U4750, U2392, U4721);
  nand ginst5407 (U4751, INSTQUEUE_REG_12__2__SCAN_IN, U4716);
  nand ginst5408 (U4752, U2414, U4706);
  nand ginst5409 (U4753, U2401, U2487);
  nand ginst5410 (U4754, U2400, U4705);
  nand ginst5411 (U4755, U2391, U4721);
  nand ginst5412 (U4756, INSTQUEUE_REG_12__1__SCAN_IN, U4716);
  nand ginst5413 (U4757, U2417, U4706);
  nand ginst5414 (U4758, U2399, U2487);
  nand ginst5415 (U4759, U2398, U4705);
  nand ginst5416 (U4760, U2390, U4721);
  nand ginst5417 (U4761, INSTQUEUE_REG_12__0__SCAN_IN, U4716);
  not ginst5418 (U4762, U3330);
  not ginst5419 (U4763, U3328);
  nand ginst5420 (U4764, U2440, U2442);
  not ginst5421 (U4765, U3331);
  nand ginst5422 (U4766, U2434, U2436);
  not ginst5423 (U4767, U3332);
  nand ginst5424 (U4768, U4516, U4517);
  nand ginst5425 (U4769, U2358, U2492);
  nand ginst5426 (U4770, U3307, U4769);
  nand ginst5427 (U4771, U4765, U4770);
  nand ginst5428 (U4772, STATE2_REG_3__SCAN_IN, U3328);
  nand ginst5429 (U4773, STATE2_REG_2__SCAN_IN, U4767);
  nand ginst5430 (U4774, U3611, U4771);
  nand ginst5431 (U4775, U2388, U2492);
  nand ginst5432 (U4776, U3307, U4775);
  nand ginst5433 (U4777, U3331, U4776);
  nand ginst5434 (U4778, STATE2_REG_2__SCAN_IN, U3332);
  nand ginst5435 (U4779, U4777, U4778);
  nand ginst5436 (U4780, U2415, U4763);
  nand ginst5437 (U4781, U2413, U2491);
  nand ginst5438 (U4782, U2412, U4762);
  nand ginst5439 (U4783, U2397, U4779);
  nand ginst5440 (U4784, INSTQUEUE_REG_11__7__SCAN_IN, U4774);
  nand ginst5441 (U4785, U2416, U4763);
  nand ginst5442 (U4786, U2411, U2491);
  nand ginst5443 (U4787, U2410, U4762);
  nand ginst5444 (U4788, U2396, U4779);
  nand ginst5445 (U4789, INSTQUEUE_REG_11__6__SCAN_IN, U4774);
  nand ginst5446 (U4790, U2420, U4763);
  nand ginst5447 (U4791, U2409, U2491);
  nand ginst5448 (U4792, U2408, U4762);
  nand ginst5449 (U4793, U2395, U4779);
  nand ginst5450 (U4794, INSTQUEUE_REG_11__5__SCAN_IN, U4774);
  nand ginst5451 (U4795, U2419, U4763);
  nand ginst5452 (U4796, U2407, U2491);
  nand ginst5453 (U4797, U2406, U4762);
  nand ginst5454 (U4798, U2394, U4779);
  nand ginst5455 (U4799, INSTQUEUE_REG_11__4__SCAN_IN, U4774);
  nand ginst5456 (U4800, U2418, U4763);
  nand ginst5457 (U4801, U2405, U2491);
  nand ginst5458 (U4802, U2404, U4762);
  nand ginst5459 (U4803, U2393, U4779);
  nand ginst5460 (U4804, INSTQUEUE_REG_11__3__SCAN_IN, U4774);
  nand ginst5461 (U4805, U2421, U4763);
  nand ginst5462 (U4806, U2403, U2491);
  nand ginst5463 (U4807, U2402, U4762);
  nand ginst5464 (U4808, U2392, U4779);
  nand ginst5465 (U4809, INSTQUEUE_REG_11__2__SCAN_IN, U4774);
  nand ginst5466 (U4810, U2414, U4763);
  nand ginst5467 (U4811, U2401, U2491);
  nand ginst5468 (U4812, U2400, U4762);
  nand ginst5469 (U4813, U2391, U4779);
  nand ginst5470 (U4814, INSTQUEUE_REG_11__1__SCAN_IN, U4774);
  nand ginst5471 (U4815, U2417, U4763);
  nand ginst5472 (U4816, U2399, U2491);
  nand ginst5473 (U4817, U2398, U4762);
  nand ginst5474 (U4818, U2390, U4779);
  nand ginst5475 (U4819, INSTQUEUE_REG_11__0__SCAN_IN, U4774);
  not ginst5476 (U4820, U3334);
  not ginst5477 (U4821, U3333);
  nand ginst5478 (U4822, U2440, U2443);
  not ginst5479 (U4823, U3335);
  not ginst5480 (U4824, U3225);
  nand ginst5481 (U4825, U4512, U4517);
  nand ginst5482 (U4826, U2358, U2494);
  nand ginst5483 (U4827, U3307, U4826);
  nand ginst5484 (U4828, U4823, U4827);
  nand ginst5485 (U4829, STATE2_REG_3__SCAN_IN, U3333);
  nand ginst5486 (U4830, STATE2_REG_2__SCAN_IN, U3225);
  nand ginst5487 (U4831, U3620, U4828);
  nand ginst5488 (U4832, U2388, U2494);
  nand ginst5489 (U4833, U3307, U4832);
  nand ginst5490 (U4834, U3335, U4833);
  nand ginst5491 (U4835, STATE2_REG_2__SCAN_IN, U4824);
  nand ginst5492 (U4836, U4834, U4835);
  nand ginst5493 (U4837, U2415, U4821);
  nand ginst5494 (U4838, U2413, U2493);
  nand ginst5495 (U4839, U2412, U4820);
  nand ginst5496 (U4840, U2397, U4836);
  nand ginst5497 (U4841, INSTQUEUE_REG_10__7__SCAN_IN, U4831);
  nand ginst5498 (U4842, U2416, U4821);
  nand ginst5499 (U4843, U2411, U2493);
  nand ginst5500 (U4844, U2410, U4820);
  nand ginst5501 (U4845, U2396, U4836);
  nand ginst5502 (U4846, INSTQUEUE_REG_10__6__SCAN_IN, U4831);
  nand ginst5503 (U4847, U2420, U4821);
  nand ginst5504 (U4848, U2409, U2493);
  nand ginst5505 (U4849, U2408, U4820);
  nand ginst5506 (U4850, U2395, U4836);
  nand ginst5507 (U4851, INSTQUEUE_REG_10__5__SCAN_IN, U4831);
  nand ginst5508 (U4852, U2419, U4821);
  nand ginst5509 (U4853, U2407, U2493);
  nand ginst5510 (U4854, U2406, U4820);
  nand ginst5511 (U4855, U2394, U4836);
  nand ginst5512 (U4856, INSTQUEUE_REG_10__4__SCAN_IN, U4831);
  nand ginst5513 (U4857, U2418, U4821);
  nand ginst5514 (U4858, U2405, U2493);
  nand ginst5515 (U4859, U2404, U4820);
  nand ginst5516 (U4860, U2393, U4836);
  nand ginst5517 (U4861, INSTQUEUE_REG_10__3__SCAN_IN, U4831);
  nand ginst5518 (U4862, U2421, U4821);
  nand ginst5519 (U4863, U2403, U2493);
  nand ginst5520 (U4864, U2402, U4820);
  nand ginst5521 (U4865, U2392, U4836);
  nand ginst5522 (U4866, INSTQUEUE_REG_10__2__SCAN_IN, U4831);
  nand ginst5523 (U4867, U2414, U4821);
  nand ginst5524 (U4868, U2401, U2493);
  nand ginst5525 (U4869, U2400, U4820);
  nand ginst5526 (U4870, U2391, U4836);
  nand ginst5527 (U4871, INSTQUEUE_REG_10__1__SCAN_IN, U4831);
  nand ginst5528 (U4872, U2417, U4821);
  nand ginst5529 (U4873, U2399, U2493);
  nand ginst5530 (U4874, U2398, U4820);
  nand ginst5531 (U4875, U2390, U4836);
  nand ginst5532 (U4876, INSTQUEUE_REG_10__0__SCAN_IN, U4831);
  not ginst5533 (U4877, U3337);
  not ginst5534 (U4878, U3336);
  nand ginst5535 (U4879, U2440, U2444);
  not ginst5536 (U4880, U3338);
  nand ginst5537 (U4881, U2434, U2437);
  not ginst5538 (U4882, U3339);
  nand ginst5539 (U4883, U4513, U4517);
  nand ginst5540 (U4884, U2358, U2496);
  nand ginst5541 (U4885, U3307, U4884);
  nand ginst5542 (U4886, U4880, U4885);
  nand ginst5543 (U4887, STATE2_REG_3__SCAN_IN, U3336);
  nand ginst5544 (U4888, STATE2_REG_2__SCAN_IN, U4882);
  nand ginst5545 (U4889, U3629, U4886);
  nand ginst5546 (U4890, U2388, U2496);
  nand ginst5547 (U4891, U3307, U4890);
  nand ginst5548 (U4892, U3338, U4891);
  nand ginst5549 (U4893, STATE2_REG_2__SCAN_IN, U3339);
  nand ginst5550 (U4894, U4892, U4893);
  nand ginst5551 (U4895, U2415, U4878);
  nand ginst5552 (U4896, U2413, U2495);
  nand ginst5553 (U4897, U2412, U4877);
  nand ginst5554 (U4898, U2397, U4894);
  nand ginst5555 (U4899, INSTQUEUE_REG_9__7__SCAN_IN, U4889);
  nand ginst5556 (U4900, U2416, U4878);
  nand ginst5557 (U4901, U2411, U2495);
  nand ginst5558 (U4902, U2410, U4877);
  nand ginst5559 (U4903, U2396, U4894);
  nand ginst5560 (U4904, INSTQUEUE_REG_9__6__SCAN_IN, U4889);
  nand ginst5561 (U4905, U2420, U4878);
  nand ginst5562 (U4906, U2409, U2495);
  nand ginst5563 (U4907, U2408, U4877);
  nand ginst5564 (U4908, U2395, U4894);
  nand ginst5565 (U4909, INSTQUEUE_REG_9__5__SCAN_IN, U4889);
  nand ginst5566 (U4910, U2419, U4878);
  nand ginst5567 (U4911, U2407, U2495);
  nand ginst5568 (U4912, U2406, U4877);
  nand ginst5569 (U4913, U2394, U4894);
  nand ginst5570 (U4914, INSTQUEUE_REG_9__4__SCAN_IN, U4889);
  nand ginst5571 (U4915, U2418, U4878);
  nand ginst5572 (U4916, U2405, U2495);
  nand ginst5573 (U4917, U2404, U4877);
  nand ginst5574 (U4918, U2393, U4894);
  nand ginst5575 (U4919, INSTQUEUE_REG_9__3__SCAN_IN, U4889);
  nand ginst5576 (U4920, U2421, U4878);
  nand ginst5577 (U4921, U2403, U2495);
  nand ginst5578 (U4922, U2402, U4877);
  nand ginst5579 (U4923, U2392, U4894);
  nand ginst5580 (U4924, INSTQUEUE_REG_9__2__SCAN_IN, U4889);
  nand ginst5581 (U4925, U2414, U4878);
  nand ginst5582 (U4926, U2401, U2495);
  nand ginst5583 (U4927, U2400, U4877);
  nand ginst5584 (U4928, U2391, U4894);
  nand ginst5585 (U4929, INSTQUEUE_REG_9__1__SCAN_IN, U4889);
  nand ginst5586 (U4930, U2417, U4878);
  nand ginst5587 (U4931, U2399, U2495);
  nand ginst5588 (U4932, U2398, U4877);
  nand ginst5589 (U4933, U2390, U4894);
  nand ginst5590 (U4934, INSTQUEUE_REG_9__0__SCAN_IN, U4889);
  not ginst5591 (U4935, U3341);
  not ginst5592 (U4936, U3340);
  nand ginst5593 (U4937, U2440, U2445);
  not ginst5594 (U4938, U3342);
  not ginst5595 (U4939, U3226);
  nand ginst5596 (U4940, U2486, U4517);
  nand ginst5597 (U4941, U2358, U2498);
  nand ginst5598 (U4942, U3307, U4941);
  nand ginst5599 (U4943, U4938, U4942);
  nand ginst5600 (U4944, STATE2_REG_3__SCAN_IN, U3340);
  nand ginst5601 (U4945, STATE2_REG_2__SCAN_IN, U3226);
  nand ginst5602 (U4946, U3638, U4943);
  nand ginst5603 (U4947, U2388, U2498);
  nand ginst5604 (U4948, U3307, U4947);
  nand ginst5605 (U4949, U3342, U4948);
  nand ginst5606 (U4950, STATE2_REG_2__SCAN_IN, U4939);
  nand ginst5607 (U4951, U4949, U4950);
  nand ginst5608 (U4952, U2415, U4936);
  nand ginst5609 (U4953, U2413, U2497);
  nand ginst5610 (U4954, U2412, U4935);
  nand ginst5611 (U4955, U2397, U4951);
  nand ginst5612 (U4956, INSTQUEUE_REG_8__7__SCAN_IN, U4946);
  nand ginst5613 (U4957, U2416, U4936);
  nand ginst5614 (U4958, U2411, U2497);
  nand ginst5615 (U4959, U2410, U4935);
  nand ginst5616 (U4960, U2396, U4951);
  nand ginst5617 (U4961, INSTQUEUE_REG_8__6__SCAN_IN, U4946);
  nand ginst5618 (U4962, U2420, U4936);
  nand ginst5619 (U4963, U2409, U2497);
  nand ginst5620 (U4964, U2408, U4935);
  nand ginst5621 (U4965, U2395, U4951);
  nand ginst5622 (U4966, INSTQUEUE_REG_8__5__SCAN_IN, U4946);
  nand ginst5623 (U4967, U2419, U4936);
  nand ginst5624 (U4968, U2407, U2497);
  nand ginst5625 (U4969, U2406, U4935);
  nand ginst5626 (U4970, U2394, U4951);
  nand ginst5627 (U4971, INSTQUEUE_REG_8__4__SCAN_IN, U4946);
  nand ginst5628 (U4972, U2418, U4936);
  nand ginst5629 (U4973, U2405, U2497);
  nand ginst5630 (U4974, U2404, U4935);
  nand ginst5631 (U4975, U2393, U4951);
  nand ginst5632 (U4976, INSTQUEUE_REG_8__3__SCAN_IN, U4946);
  nand ginst5633 (U4977, U2421, U4936);
  nand ginst5634 (U4978, U2403, U2497);
  nand ginst5635 (U4979, U2402, U4935);
  nand ginst5636 (U4980, U2392, U4951);
  nand ginst5637 (U4981, INSTQUEUE_REG_8__2__SCAN_IN, U4946);
  nand ginst5638 (U4982, U2414, U4936);
  nand ginst5639 (U4983, U2401, U2497);
  nand ginst5640 (U4984, U2400, U4935);
  nand ginst5641 (U4985, U2391, U4951);
  nand ginst5642 (U4986, INSTQUEUE_REG_8__1__SCAN_IN, U4946);
  nand ginst5643 (U4987, U2417, U4936);
  nand ginst5644 (U4988, U2399, U2497);
  nand ginst5645 (U4989, U2398, U4935);
  nand ginst5646 (U4990, U2390, U4951);
  nand ginst5647 (U4991, INSTQUEUE_REG_8__0__SCAN_IN, U4946);
  not ginst5648 (U4992, U3346);
  nand ginst5649 (U4993, U2439, U2442);
  not ginst5650 (U4994, U3348);
  nand ginst5651 (U4995, U2433, U2436);
  not ginst5652 (U4996, U3349);
  nand ginst5653 (U4997, U2358, U2500);
  nand ginst5654 (U4998, U3307, U4997);
  nand ginst5655 (U4999, U4994, U4998);
  nand ginst5656 (U5000, STATE2_REG_3__SCAN_IN, U3343);
  nand ginst5657 (U5001, STATE2_REG_2__SCAN_IN, U4996);
  nand ginst5658 (U5002, U3647, U4999);
  nand ginst5659 (U5003, U2388, U2500);
  nand ginst5660 (U5004, U3307, U5003);
  nand ginst5661 (U5005, U3348, U5004);
  nand ginst5662 (U5006, STATE2_REG_2__SCAN_IN, U3349);
  nand ginst5663 (U5007, U5005, U5006);
  nand ginst5664 (U5008, U2415, U4525);
  nand ginst5665 (U5009, U2413, U4226);
  nand ginst5666 (U5010, U2412, U4992);
  nand ginst5667 (U5011, U2397, U5007);
  nand ginst5668 (U5012, INSTQUEUE_REG_7__7__SCAN_IN, U5002);
  nand ginst5669 (U5013, U2416, U4525);
  nand ginst5670 (U5014, U2411, U4226);
  nand ginst5671 (U5015, U2410, U4992);
  nand ginst5672 (U5016, U2396, U5007);
  nand ginst5673 (U5017, INSTQUEUE_REG_7__6__SCAN_IN, U5002);
  nand ginst5674 (U5018, U2420, U4525);
  nand ginst5675 (U5019, U2409, U4226);
  nand ginst5676 (U5020, U2408, U4992);
  nand ginst5677 (U5021, U2395, U5007);
  nand ginst5678 (U5022, INSTQUEUE_REG_7__5__SCAN_IN, U5002);
  nand ginst5679 (U5023, U2419, U4525);
  nand ginst5680 (U5024, U2407, U4226);
  nand ginst5681 (U5025, U2406, U4992);
  nand ginst5682 (U5026, U2394, U5007);
  nand ginst5683 (U5027, INSTQUEUE_REG_7__4__SCAN_IN, U5002);
  nand ginst5684 (U5028, U2418, U4525);
  nand ginst5685 (U5029, U2405, U4226);
  nand ginst5686 (U5030, U2404, U4992);
  nand ginst5687 (U5031, U2393, U5007);
  nand ginst5688 (U5032, INSTQUEUE_REG_7__3__SCAN_IN, U5002);
  nand ginst5689 (U5033, U2421, U4525);
  nand ginst5690 (U5034, U2403, U4226);
  nand ginst5691 (U5035, U2402, U4992);
  nand ginst5692 (U5036, U2392, U5007);
  nand ginst5693 (U5037, INSTQUEUE_REG_7__2__SCAN_IN, U5002);
  nand ginst5694 (U5038, U2414, U4525);
  nand ginst5695 (U5039, U2401, U4226);
  nand ginst5696 (U5040, U2400, U4992);
  nand ginst5697 (U5041, U2391, U5007);
  nand ginst5698 (U5042, INSTQUEUE_REG_7__1__SCAN_IN, U5002);
  nand ginst5699 (U5043, U2417, U4525);
  nand ginst5700 (U5044, U2399, U4226);
  nand ginst5701 (U5045, U2398, U4992);
  nand ginst5702 (U5046, U2390, U5007);
  nand ginst5703 (U5047, INSTQUEUE_REG_7__0__SCAN_IN, U5002);
  not ginst5704 (U5048, U3351);
  not ginst5705 (U5049, U3350);
  nand ginst5706 (U5050, U2439, U2443);
  not ginst5707 (U5051, U3352);
  not ginst5708 (U5052, U3227);
  nand ginst5709 (U5053, U2474, U4512);
  nand ginst5710 (U5054, U2358, U2502);
  nand ginst5711 (U5055, U3307, U5054);
  nand ginst5712 (U5056, U5051, U5055);
  nand ginst5713 (U5057, STATE2_REG_3__SCAN_IN, U3350);
  nand ginst5714 (U5058, STATE2_REG_2__SCAN_IN, U3227);
  nand ginst5715 (U5059, U3656, U5056);
  nand ginst5716 (U5060, U2388, U2502);
  nand ginst5717 (U5061, U3307, U5060);
  nand ginst5718 (U5062, U3352, U5061);
  nand ginst5719 (U5063, STATE2_REG_2__SCAN_IN, U5052);
  nand ginst5720 (U5064, U5062, U5063);
  nand ginst5721 (U5065, U2415, U5049);
  nand ginst5722 (U5066, U2413, U2501);
  nand ginst5723 (U5067, U2412, U5048);
  nand ginst5724 (U5068, U2397, U5064);
  nand ginst5725 (U5069, INSTQUEUE_REG_6__7__SCAN_IN, U5059);
  nand ginst5726 (U5070, U2416, U5049);
  nand ginst5727 (U5071, U2411, U2501);
  nand ginst5728 (U5072, U2410, U5048);
  nand ginst5729 (U5073, U2396, U5064);
  nand ginst5730 (U5074, INSTQUEUE_REG_6__6__SCAN_IN, U5059);
  nand ginst5731 (U5075, U2420, U5049);
  nand ginst5732 (U5076, U2409, U2501);
  nand ginst5733 (U5077, U2408, U5048);
  nand ginst5734 (U5078, U2395, U5064);
  nand ginst5735 (U5079, INSTQUEUE_REG_6__5__SCAN_IN, U5059);
  nand ginst5736 (U5080, U2419, U5049);
  nand ginst5737 (U5081, U2407, U2501);
  nand ginst5738 (U5082, U2406, U5048);
  nand ginst5739 (U5083, U2394, U5064);
  nand ginst5740 (U5084, INSTQUEUE_REG_6__4__SCAN_IN, U5059);
  nand ginst5741 (U5085, U2418, U5049);
  nand ginst5742 (U5086, U2405, U2501);
  nand ginst5743 (U5087, U2404, U5048);
  nand ginst5744 (U5088, U2393, U5064);
  nand ginst5745 (U5089, INSTQUEUE_REG_6__3__SCAN_IN, U5059);
  nand ginst5746 (U5090, U2421, U5049);
  nand ginst5747 (U5091, U2403, U2501);
  nand ginst5748 (U5092, U2402, U5048);
  nand ginst5749 (U5093, U2392, U5064);
  nand ginst5750 (U5094, INSTQUEUE_REG_6__2__SCAN_IN, U5059);
  nand ginst5751 (U5095, U2414, U5049);
  nand ginst5752 (U5096, U2401, U2501);
  nand ginst5753 (U5097, U2400, U5048);
  nand ginst5754 (U5098, U2391, U5064);
  nand ginst5755 (U5099, INSTQUEUE_REG_6__1__SCAN_IN, U5059);
  nand ginst5756 (U5100, U2417, U5049);
  nand ginst5757 (U5101, U2399, U2501);
  nand ginst5758 (U5102, U2398, U5048);
  nand ginst5759 (U5103, U2390, U5064);
  nand ginst5760 (U5104, INSTQUEUE_REG_6__0__SCAN_IN, U5059);
  not ginst5761 (U5105, U3354);
  not ginst5762 (U5106, U3353);
  nand ginst5763 (U5107, U2439, U2444);
  not ginst5764 (U5108, U3355);
  nand ginst5765 (U5109, U2433, U2437);
  not ginst5766 (U5110, U3356);
  nand ginst5767 (U5111, U2474, U4513);
  nand ginst5768 (U5112, U2358, U2504);
  nand ginst5769 (U5113, U3307, U5112);
  nand ginst5770 (U5114, U5108, U5113);
  nand ginst5771 (U5115, STATE2_REG_3__SCAN_IN, U3353);
  nand ginst5772 (U5116, STATE2_REG_2__SCAN_IN, U5110);
  nand ginst5773 (U5117, U3665, U5114);
  nand ginst5774 (U5118, U2388, U2504);
  nand ginst5775 (U5119, U3307, U5118);
  nand ginst5776 (U5120, U3355, U5119);
  nand ginst5777 (U5121, STATE2_REG_2__SCAN_IN, U3356);
  nand ginst5778 (U5122, U5120, U5121);
  nand ginst5779 (U5123, U2415, U5106);
  nand ginst5780 (U5124, U2413, U2503);
  nand ginst5781 (U5125, U2412, U5105);
  nand ginst5782 (U5126, U2397, U5122);
  nand ginst5783 (U5127, INSTQUEUE_REG_5__7__SCAN_IN, U5117);
  nand ginst5784 (U5128, U2416, U5106);
  nand ginst5785 (U5129, U2411, U2503);
  nand ginst5786 (U5130, U2410, U5105);
  nand ginst5787 (U5131, U2396, U5122);
  nand ginst5788 (U5132, INSTQUEUE_REG_5__6__SCAN_IN, U5117);
  nand ginst5789 (U5133, U2420, U5106);
  nand ginst5790 (U5134, U2409, U2503);
  nand ginst5791 (U5135, U2408, U5105);
  nand ginst5792 (U5136, U2395, U5122);
  nand ginst5793 (U5137, INSTQUEUE_REG_5__5__SCAN_IN, U5117);
  nand ginst5794 (U5138, U2419, U5106);
  nand ginst5795 (U5139, U2407, U2503);
  nand ginst5796 (U5140, U2406, U5105);
  nand ginst5797 (U5141, U2394, U5122);
  nand ginst5798 (U5142, INSTQUEUE_REG_5__4__SCAN_IN, U5117);
  nand ginst5799 (U5143, U2418, U5106);
  nand ginst5800 (U5144, U2405, U2503);
  nand ginst5801 (U5145, U2404, U5105);
  nand ginst5802 (U5146, U2393, U5122);
  nand ginst5803 (U5147, INSTQUEUE_REG_5__3__SCAN_IN, U5117);
  nand ginst5804 (U5148, U2421, U5106);
  nand ginst5805 (U5149, U2403, U2503);
  nand ginst5806 (U5150, U2402, U5105);
  nand ginst5807 (U5151, U2392, U5122);
  nand ginst5808 (U5152, INSTQUEUE_REG_5__2__SCAN_IN, U5117);
  nand ginst5809 (U5153, U2414, U5106);
  nand ginst5810 (U5154, U2401, U2503);
  nand ginst5811 (U5155, U2400, U5105);
  nand ginst5812 (U5156, U2391, U5122);
  nand ginst5813 (U5157, INSTQUEUE_REG_5__1__SCAN_IN, U5117);
  nand ginst5814 (U5158, U2417, U5106);
  nand ginst5815 (U5159, U2399, U2503);
  nand ginst5816 (U5160, U2398, U5105);
  nand ginst5817 (U5161, U2390, U5122);
  nand ginst5818 (U5162, INSTQUEUE_REG_5__0__SCAN_IN, U5117);
  not ginst5819 (U5163, U3358);
  not ginst5820 (U5164, U3357);
  nand ginst5821 (U5165, U2439, U2445);
  not ginst5822 (U5166, U3359);
  not ginst5823 (U5167, U3228);
  nand ginst5824 (U5168, U2474, U2486);
  nand ginst5825 (U5169, U2358, U2506);
  nand ginst5826 (U5170, U3307, U5169);
  nand ginst5827 (U5171, U5166, U5170);
  nand ginst5828 (U5172, STATE2_REG_3__SCAN_IN, U3357);
  nand ginst5829 (U5173, STATE2_REG_2__SCAN_IN, U3228);
  nand ginst5830 (U5174, U3674, U5171);
  nand ginst5831 (U5175, U2388, U2506);
  nand ginst5832 (U5176, U3307, U5175);
  nand ginst5833 (U5177, U3359, U5176);
  nand ginst5834 (U5178, STATE2_REG_2__SCAN_IN, U5167);
  nand ginst5835 (U5179, U5177, U5178);
  nand ginst5836 (U5180, U2415, U5164);
  nand ginst5837 (U5181, U2413, U2505);
  nand ginst5838 (U5182, U2412, U5163);
  nand ginst5839 (U5183, U2397, U5179);
  nand ginst5840 (U5184, INSTQUEUE_REG_4__7__SCAN_IN, U5174);
  nand ginst5841 (U5185, U2416, U5164);
  nand ginst5842 (U5186, U2411, U2505);
  nand ginst5843 (U5187, U2410, U5163);
  nand ginst5844 (U5188, U2396, U5179);
  nand ginst5845 (U5189, INSTQUEUE_REG_4__6__SCAN_IN, U5174);
  nand ginst5846 (U5190, U2420, U5164);
  nand ginst5847 (U5191, U2409, U2505);
  nand ginst5848 (U5192, U2408, U5163);
  nand ginst5849 (U5193, U2395, U5179);
  nand ginst5850 (U5194, INSTQUEUE_REG_4__5__SCAN_IN, U5174);
  nand ginst5851 (U5195, U2419, U5164);
  nand ginst5852 (U5196, U2407, U2505);
  nand ginst5853 (U5197, U2406, U5163);
  nand ginst5854 (U5198, U2394, U5179);
  nand ginst5855 (U5199, INSTQUEUE_REG_4__4__SCAN_IN, U5174);
  nand ginst5856 (U5200, U2418, U5164);
  nand ginst5857 (U5201, U2405, U2505);
  nand ginst5858 (U5202, U2404, U5163);
  nand ginst5859 (U5203, U2393, U5179);
  nand ginst5860 (U5204, INSTQUEUE_REG_4__3__SCAN_IN, U5174);
  nand ginst5861 (U5205, U2421, U5164);
  nand ginst5862 (U5206, U2403, U2505);
  nand ginst5863 (U5207, U2402, U5163);
  nand ginst5864 (U5208, U2392, U5179);
  nand ginst5865 (U5209, INSTQUEUE_REG_4__2__SCAN_IN, U5174);
  nand ginst5866 (U5210, U2414, U5164);
  nand ginst5867 (U5211, U2401, U2505);
  nand ginst5868 (U5212, U2400, U5163);
  nand ginst5869 (U5213, U2391, U5179);
  nand ginst5870 (U5214, INSTQUEUE_REG_4__1__SCAN_IN, U5174);
  nand ginst5871 (U5215, U2417, U5164);
  nand ginst5872 (U5216, U2399, U2505);
  nand ginst5873 (U5217, U2398, U5163);
  nand ginst5874 (U5218, U2390, U5179);
  nand ginst5875 (U5219, INSTQUEUE_REG_4__0__SCAN_IN, U5174);
  not ginst5876 (U5220, U3361);
  not ginst5877 (U5221, U3360);
  nand ginst5878 (U5222, U2441, U2442);
  not ginst5879 (U5223, U3362);
  nand ginst5880 (U5224, U2435, U2436);
  not ginst5881 (U5225, U3363);
  nand ginst5882 (U5226, U2508, U4516);
  nand ginst5883 (U5227, U2358, U2511);
  nand ginst5884 (U5228, U3307, U5227);
  nand ginst5885 (U5229, U5223, U5228);
  nand ginst5886 (U5230, STATE2_REG_3__SCAN_IN, U3360);
  nand ginst5887 (U5231, STATE2_REG_2__SCAN_IN, U5225);
  nand ginst5888 (U5232, U3683, U5229);
  nand ginst5889 (U5233, U2388, U2511);
  nand ginst5890 (U5234, U3307, U5233);
  nand ginst5891 (U5235, U3362, U5234);
  nand ginst5892 (U5236, STATE2_REG_2__SCAN_IN, U3363);
  nand ginst5893 (U5237, U5235, U5236);
  nand ginst5894 (U5238, U2415, U5221);
  nand ginst5895 (U5239, U2413, U2509);
  nand ginst5896 (U5240, U2412, U5220);
  nand ginst5897 (U5241, U2397, U5237);
  nand ginst5898 (U5242, INSTQUEUE_REG_3__7__SCAN_IN, U5232);
  nand ginst5899 (U5243, U2416, U5221);
  nand ginst5900 (U5244, U2411, U2509);
  nand ginst5901 (U5245, U2410, U5220);
  nand ginst5902 (U5246, U2396, U5237);
  nand ginst5903 (U5247, INSTQUEUE_REG_3__6__SCAN_IN, U5232);
  nand ginst5904 (U5248, U2420, U5221);
  nand ginst5905 (U5249, U2409, U2509);
  nand ginst5906 (U5250, U2408, U5220);
  nand ginst5907 (U5251, U2395, U5237);
  nand ginst5908 (U5252, INSTQUEUE_REG_3__5__SCAN_IN, U5232);
  nand ginst5909 (U5253, U2419, U5221);
  nand ginst5910 (U5254, U2407, U2509);
  nand ginst5911 (U5255, U2406, U5220);
  nand ginst5912 (U5256, U2394, U5237);
  nand ginst5913 (U5257, INSTQUEUE_REG_3__4__SCAN_IN, U5232);
  nand ginst5914 (U5258, U2418, U5221);
  nand ginst5915 (U5259, U2405, U2509);
  nand ginst5916 (U5260, U2404, U5220);
  nand ginst5917 (U5261, U2393, U5237);
  nand ginst5918 (U5262, INSTQUEUE_REG_3__3__SCAN_IN, U5232);
  nand ginst5919 (U5263, U2421, U5221);
  nand ginst5920 (U5264, U2403, U2509);
  nand ginst5921 (U5265, U2402, U5220);
  nand ginst5922 (U5266, U2392, U5237);
  nand ginst5923 (U5267, INSTQUEUE_REG_3__2__SCAN_IN, U5232);
  nand ginst5924 (U5268, U2414, U5221);
  nand ginst5925 (U5269, U2401, U2509);
  nand ginst5926 (U5270, U2400, U5220);
  nand ginst5927 (U5271, U2391, U5237);
  nand ginst5928 (U5272, INSTQUEUE_REG_3__1__SCAN_IN, U5232);
  nand ginst5929 (U5273, U2417, U5221);
  nand ginst5930 (U5274, U2399, U2509);
  nand ginst5931 (U5275, U2398, U5220);
  nand ginst5932 (U5276, U2390, U5237);
  nand ginst5933 (U5277, INSTQUEUE_REG_3__0__SCAN_IN, U5232);
  not ginst5934 (U5278, U3365);
  not ginst5935 (U5279, U3364);
  nand ginst5936 (U5280, U2441, U2443);
  not ginst5937 (U5281, U3366);
  not ginst5938 (U5282, U3229);
  nand ginst5939 (U5283, U2508, U4512);
  nand ginst5940 (U5284, U2358, U2513);
  nand ginst5941 (U5285, U3307, U5284);
  nand ginst5942 (U5286, U5281, U5285);
  nand ginst5943 (U5287, STATE2_REG_3__SCAN_IN, U3364);
  nand ginst5944 (U5288, STATE2_REG_2__SCAN_IN, U3229);
  nand ginst5945 (U5289, U3692, U5286);
  nand ginst5946 (U5290, U2388, U2513);
  nand ginst5947 (U5291, U3307, U5290);
  nand ginst5948 (U5292, U3366, U5291);
  nand ginst5949 (U5293, STATE2_REG_2__SCAN_IN, U5282);
  nand ginst5950 (U5294, U5292, U5293);
  nand ginst5951 (U5295, U2415, U5279);
  nand ginst5952 (U5296, U2413, U2512);
  nand ginst5953 (U5297, U2412, U5278);
  nand ginst5954 (U5298, U2397, U5294);
  nand ginst5955 (U5299, INSTQUEUE_REG_2__7__SCAN_IN, U5289);
  nand ginst5956 (U5300, U2416, U5279);
  nand ginst5957 (U5301, U2411, U2512);
  nand ginst5958 (U5302, U2410, U5278);
  nand ginst5959 (U5303, U2396, U5294);
  nand ginst5960 (U5304, INSTQUEUE_REG_2__6__SCAN_IN, U5289);
  nand ginst5961 (U5305, U2420, U5279);
  nand ginst5962 (U5306, U2409, U2512);
  nand ginst5963 (U5307, U2408, U5278);
  nand ginst5964 (U5308, U2395, U5294);
  nand ginst5965 (U5309, INSTQUEUE_REG_2__5__SCAN_IN, U5289);
  nand ginst5966 (U5310, U2419, U5279);
  nand ginst5967 (U5311, U2407, U2512);
  nand ginst5968 (U5312, U2406, U5278);
  nand ginst5969 (U5313, U2394, U5294);
  nand ginst5970 (U5314, INSTQUEUE_REG_2__4__SCAN_IN, U5289);
  nand ginst5971 (U5315, U2418, U5279);
  nand ginst5972 (U5316, U2405, U2512);
  nand ginst5973 (U5317, U2404, U5278);
  nand ginst5974 (U5318, U2393, U5294);
  nand ginst5975 (U5319, INSTQUEUE_REG_2__3__SCAN_IN, U5289);
  nand ginst5976 (U5320, U2421, U5279);
  nand ginst5977 (U5321, U2403, U2512);
  nand ginst5978 (U5322, U2402, U5278);
  nand ginst5979 (U5323, U2392, U5294);
  nand ginst5980 (U5324, INSTQUEUE_REG_2__2__SCAN_IN, U5289);
  nand ginst5981 (U5325, U2414, U5279);
  nand ginst5982 (U5326, U2401, U2512);
  nand ginst5983 (U5327, U2400, U5278);
  nand ginst5984 (U5328, U2391, U5294);
  nand ginst5985 (U5329, INSTQUEUE_REG_2__1__SCAN_IN, U5289);
  nand ginst5986 (U5330, U2417, U5279);
  nand ginst5987 (U5331, U2399, U2512);
  nand ginst5988 (U5332, U2398, U5278);
  nand ginst5989 (U5333, U2390, U5294);
  nand ginst5990 (U5334, INSTQUEUE_REG_2__0__SCAN_IN, U5289);
  not ginst5991 (U5335, U3368);
  not ginst5992 (U5336, U3367);
  nand ginst5993 (U5337, U2441, U2444);
  not ginst5994 (U5338, U3369);
  nand ginst5995 (U5339, U2435, U2437);
  not ginst5996 (U5340, U3370);
  nand ginst5997 (U5341, U2508, U4513);
  nand ginst5998 (U5342, U2358, U2515);
  nand ginst5999 (U5343, U3307, U5342);
  nand ginst6000 (U5344, U5338, U5343);
  nand ginst6001 (U5345, STATE2_REG_3__SCAN_IN, U3367);
  nand ginst6002 (U5346, STATE2_REG_2__SCAN_IN, U5340);
  nand ginst6003 (U5347, U3701, U5344);
  nand ginst6004 (U5348, U2388, U2515);
  nand ginst6005 (U5349, U3307, U5348);
  nand ginst6006 (U5350, U3369, U5349);
  nand ginst6007 (U5351, STATE2_REG_2__SCAN_IN, U3370);
  nand ginst6008 (U5352, U5350, U5351);
  nand ginst6009 (U5353, U2415, U5336);
  nand ginst6010 (U5354, U2413, U2514);
  nand ginst6011 (U5355, U2412, U5335);
  nand ginst6012 (U5356, U2397, U5352);
  nand ginst6013 (U5357, INSTQUEUE_REG_1__7__SCAN_IN, U5347);
  nand ginst6014 (U5358, U2416, U5336);
  nand ginst6015 (U5359, U2411, U2514);
  nand ginst6016 (U5360, U2410, U5335);
  nand ginst6017 (U5361, U2396, U5352);
  nand ginst6018 (U5362, INSTQUEUE_REG_1__6__SCAN_IN, U5347);
  nand ginst6019 (U5363, U2420, U5336);
  nand ginst6020 (U5364, U2409, U2514);
  nand ginst6021 (U5365, U2408, U5335);
  nand ginst6022 (U5366, U2395, U5352);
  nand ginst6023 (U5367, INSTQUEUE_REG_1__5__SCAN_IN, U5347);
  nand ginst6024 (U5368, U2419, U5336);
  nand ginst6025 (U5369, U2407, U2514);
  nand ginst6026 (U5370, U2406, U5335);
  nand ginst6027 (U5371, U2394, U5352);
  nand ginst6028 (U5372, INSTQUEUE_REG_1__4__SCAN_IN, U5347);
  nand ginst6029 (U5373, U2418, U5336);
  nand ginst6030 (U5374, U2405, U2514);
  nand ginst6031 (U5375, U2404, U5335);
  nand ginst6032 (U5376, U2393, U5352);
  nand ginst6033 (U5377, INSTQUEUE_REG_1__3__SCAN_IN, U5347);
  nand ginst6034 (U5378, U2421, U5336);
  nand ginst6035 (U5379, U2403, U2514);
  nand ginst6036 (U5380, U2402, U5335);
  nand ginst6037 (U5381, U2392, U5352);
  nand ginst6038 (U5382, INSTQUEUE_REG_1__2__SCAN_IN, U5347);
  nand ginst6039 (U5383, U2414, U5336);
  nand ginst6040 (U5384, U2401, U2514);
  nand ginst6041 (U5385, U2400, U5335);
  nand ginst6042 (U5386, U2391, U5352);
  nand ginst6043 (U5387, INSTQUEUE_REG_1__1__SCAN_IN, U5347);
  nand ginst6044 (U5388, U2417, U5336);
  nand ginst6045 (U5389, U2399, U2514);
  nand ginst6046 (U5390, U2398, U5335);
  nand ginst6047 (U5391, U2390, U5352);
  nand ginst6048 (U5392, INSTQUEUE_REG_1__0__SCAN_IN, U5347);
  not ginst6049 (U5393, U3372);
  not ginst6050 (U5394, U3371);
  nand ginst6051 (U5395, U2441, U2445);
  not ginst6052 (U5396, U3373);
  not ginst6053 (U5397, U3230);
  nand ginst6054 (U5398, U2486, U2508);
  nand ginst6055 (U5399, U2358, U2517);
  nand ginst6056 (U5400, U3307, U5399);
  nand ginst6057 (U5401, U5396, U5400);
  nand ginst6058 (U5402, STATE2_REG_3__SCAN_IN, U3371);
  nand ginst6059 (U5403, STATE2_REG_2__SCAN_IN, U3230);
  nand ginst6060 (U5404, U3710, U5401);
  nand ginst6061 (U5405, U2388, U2517);
  nand ginst6062 (U5406, U3307, U5405);
  nand ginst6063 (U5407, U3373, U5406);
  nand ginst6064 (U5408, STATE2_REG_2__SCAN_IN, U5397);
  nand ginst6065 (U5409, U5407, U5408);
  nand ginst6066 (U5410, U2415, U5394);
  nand ginst6067 (U5411, U2413, U2516);
  nand ginst6068 (U5412, U2412, U5393);
  nand ginst6069 (U5413, U2397, U5409);
  nand ginst6070 (U5414, INSTQUEUE_REG_0__7__SCAN_IN, U5404);
  nand ginst6071 (U5415, U2416, U5394);
  nand ginst6072 (U5416, U2411, U2516);
  nand ginst6073 (U5417, U2410, U5393);
  nand ginst6074 (U5418, U2396, U5409);
  nand ginst6075 (U5419, INSTQUEUE_REG_0__6__SCAN_IN, U5404);
  nand ginst6076 (U5420, U2420, U5394);
  nand ginst6077 (U5421, U2409, U2516);
  nand ginst6078 (U5422, U2408, U5393);
  nand ginst6079 (U5423, U2395, U5409);
  nand ginst6080 (U5424, INSTQUEUE_REG_0__5__SCAN_IN, U5404);
  nand ginst6081 (U5425, U2419, U5394);
  nand ginst6082 (U5426, U2407, U2516);
  nand ginst6083 (U5427, U2406, U5393);
  nand ginst6084 (U5428, U2394, U5409);
  nand ginst6085 (U5429, U2418, U5394);
  nand ginst6086 (U5430, U2405, U2516);
  nand ginst6087 (U5431, U2404, U5393);
  nand ginst6088 (U5432, U2393, U5409);
  nand ginst6089 (U5433, INSTQUEUE_REG_0__3__SCAN_IN, U5404);
  nand ginst6090 (U5434, U2421, U5394);
  nand ginst6091 (U5435, U2403, U2516);
  nand ginst6092 (U5436, U2402, U5393);
  nand ginst6093 (U5437, U2392, U5409);
  nand ginst6094 (U5438, INSTQUEUE_REG_0__2__SCAN_IN, U5404);
  nand ginst6095 (U5439, U2414, U5394);
  nand ginst6096 (U5440, U2401, U2516);
  nand ginst6097 (U5441, U2400, U5393);
  nand ginst6098 (U5442, U2391, U5409);
  nand ginst6099 (U5443, INSTQUEUE_REG_0__1__SCAN_IN, U5404);
  nand ginst6100 (U5444, U2417, U5394);
  nand ginst6101 (U5445, U2399, U2516);
  nand ginst6102 (U5446, U2398, U5393);
  nand ginst6103 (U5447, U2390, U5409);
  nand ginst6104 (U5448, INSTQUEUE_REG_0__0__SCAN_IN, U5404);
  not ginst6105 (U5449, U3410);
  nand ginst6106 (U5450, U3378, U3381, U4491);
  nand ginst6107 (U5451, U4161, U4388, U4448);
  not ginst6108 (U5452, U3231);
  nand ginst6109 (U5453, U3276, U4482);
  nand ginst6110 (U5454, U3270, U5452, U5453);
  nand ginst6111 (U5455, U2452, U3720);
  nand ginst6112 (U5456, U4196, U5450);
  nand ginst6113 (U5457, U3721, U7597);
  nand ginst6114 (U5458, GTE_485_U6, U3244, U4203);
  nand ginst6115 (U5459, U2449, U7482);
  nand ginst6116 (U5460, U4245, U4491);
  not ginst6117 (U5461, U4170);
  nand ginst6118 (U5462, U2368, U4170);
  nand ginst6119 (U5463, STATE2_REG_3__SCAN_IN, U3281);
  not ginst6120 (U5464, U4160);
  nand ginst6121 (U5465, INSTQUEUERD_ADDR_REG_2__SCAN_IN, INSTQUEUERD_ADDR_REG_1__SCAN_IN);
  nand ginst6122 (U5466, INSTQUEUERD_ADDR_REG_3__SCAN_IN, U5465);
  nand ginst6123 (U5467, INSTQUEUERD_ADDR_REG_1__SCAN_IN, U4369);
  not ginst6124 (U5468, U3429);
  nand ginst6125 (U5469, INSTQUEUERD_ADDR_REG_2__SCAN_IN, U3486);
  nand ginst6126 (U5470, INSTQUEUERD_ADDR_REG_3__SCAN_IN, U5469);
  not ginst6127 (U5471, U3425);
  nand ginst6128 (U5472, U3251, U3262);
  nand ginst6129 (U5473, INSTQUEUERD_ADDR_REG_3__SCAN_IN, U5472);
  nand ginst6130 (U5474, U2469, U3262);
  nand ginst6131 (U5475, U3277, U4482);
  nand ginst6132 (U5476, U2605, U4388);
  nand ginst6133 (U5477, U7482, U7691, U7692);
  nand ginst6134 (U5478, U4437, U5476);
  nand ginst6135 (U5479, U3381, U3396, U4388);
  nand ginst6136 (U5480, U4159, U5479);
  nand ginst6137 (U5481, U5480, U7617);
  nand ginst6138 (U5482, U4159, U4448);
  nand ginst6139 (U5483, U3382, U5482);
  nand ginst6140 (U5484, U4196, U5450);
  nand ginst6141 (U5485, U4245, U4491);
  nand ginst6142 (U5486, U3258, U5483);
  nand ginst6143 (U5487, U4482, U7695);
  nand ginst6144 (U5488, U3231, U4178);
  nand ginst6145 (U5489, U3279, U4205);
  nand ginst6146 (U5490, U3728, U5489);
  nand ginst6147 (U5491, R2182_U25, U7497);
  nand ginst6148 (U5492, U3425, U4206);
  nand ginst6149 (U5493, U3429, U4202);
  nand ginst6150 (U5494, U3735, U5491);
  nand ginst6151 (U5495, U3425, U4240);
  nand ginst6152 (U5496, U2427, U5494);
  nand ginst6153 (U5497, U5495, U5496);
  nand ginst6154 (U5498, INSTQUEUERD_ADDR_REG_2__SCAN_IN, U3262);
  not ginst6155 (U5499, U3388);
  nand ginst6156 (U5500, R2182_U42, U7497);
  nand ginst6157 (U5501, U3443, U4202);
  nand ginst6158 (U5502, U3737, U5500);
  nand ginst6159 (U5503, U2446, U3457);
  nand ginst6160 (U5504, U3388, U4240);
  nand ginst6161 (U5505, U2427, U5502);
  nand ginst6162 (U5506, U5503, U5504, U5505);
  not ginst6163 (U5507, U3389);
  nand ginst6164 (U5508, U2431, U4237);
  nand ginst6165 (U5509, U3279, U5508);
  nand ginst6166 (U5510, U5507, U5509);
  nand ginst6167 (U5511, R2182_U33, U7497);
  nand ginst6168 (U5512, U3252, U4202);
  nand ginst6169 (U5513, U3738, U5511);
  nand ginst6170 (U5514, U2446, U7700);
  nand ginst6171 (U5515, U4240, U5507);
  nand ginst6172 (U5516, U2427, U5513);
  nand ginst6173 (U5517, U5514, U5515, U5516);
  nand ginst6174 (U5518, R2182_U34, U7497);
  nand ginst6175 (U5519, U4163, U5518);
  nand ginst6176 (U5520, U3253, U4240);
  nand ginst6177 (U5521, U2427, U5519);
  nand ginst6178 (U5522, STATE2_REG_1__SCAN_IN, U7703);
  nand ginst6179 (U5523, U5520, U5521, U5522);
  nand ginst6180 (U5524, STATE2_REG_0__SCAN_IN, LT_589_U6, U2428);
  not ginst6181 (U5525, U3391);
  nand ginst6182 (U5526, STATE2_REG_1__SCAN_IN, U3283);
  nand ginst6183 (U5527, U3441, U4515);
  nand ginst6184 (U5528, U3345, U5527);
  nand ginst6185 (U5529, U3346, U5528);
  nand ginst6186 (U5530, U2388, U5529);
  nand ginst6187 (U5531, R2182_U25, U5526);
  nand ginst6188 (U5532, R2144_U8, U4214);
  nand ginst6189 (U5533, U3739, U5530);
  nand ginst6190 (U5534, U2388, U7721);
  nand ginst6191 (U5535, R2182_U42, U5526);
  nand ginst6192 (U5536, R2144_U49, U4214);
  nand ginst6193 (U5537, U3740, U5534);
  nand ginst6194 (U5538, U3313, U3320);
  nand ginst6195 (U5539, U2388, U5538);
  nand ginst6196 (U5540, R2182_U33, U5526);
  nand ginst6197 (U5541, R2144_U50, U4214);
  nand ginst6198 (U5542, U3741, U5539);
  nand ginst6199 (U5543, R2182_U34, U5526);
  nand ginst6200 (U5544, R2144_U43, U4197);
  nand ginst6201 (U5545, U4233, U5543, U5544);
  nand ginst6202 (U5546, U3259, U4465);
  nand ginst6203 (U5547, U2431, U4248);
  nand ginst6204 (U5548, U2518, U5547, U7730, U7731);
  nand ginst6205 (U5549, U4180, U4223, U4491);
  nand ginst6206 (U5550, U2368, U5548);
  nand ginst6207 (U5551, U3250, U4191);
  not ginst6208 (U5552, U3401);
  nand ginst6209 (U5553, U4196, U4250);
  nand ginst6210 (U5554, U2389, U4244);
  nand ginst6211 (U5555, U4238, U4254);
  nand ginst6212 (U5556, U4252, U4482);
  nand ginst6213 (U5557, U2519, U3746);
  nand ginst6214 (U5558, R2099_U86, U2380);
  nand ginst6215 (U5559, R2027_U5, U2378);
  nand ginst6216 (U5560, R2278_U17, U2377);
  nand ginst6217 (U5561, ADD_405_U4, U2375);
  nand ginst6218 (U5562, INSTADDRPOINTER_REG_0__SCAN_IN, U2374);
  nand ginst6219 (U5563, REIP_REG_0__SCAN_IN, U2370);
  nand ginst6220 (U5564, INSTADDRPOINTER_REG_0__SCAN_IN, U5552);
  nand ginst6221 (U5565, R2099_U87, U2380);
  nand ginst6222 (U5566, R2027_U71, U2378);
  nand ginst6223 (U5567, R2278_U42, U2377);
  nand ginst6224 (U5568, ADD_405_U81, U2375);
  nand ginst6225 (U5569, ADD_515_U4, U2374);
  nand ginst6226 (U5570, REIP_REG_1__SCAN_IN, U2370);
  nand ginst6227 (U5571, INSTADDRPOINTER_REG_1__SCAN_IN, U5552);
  nand ginst6228 (U5572, R2099_U138, U2380);
  nand ginst6229 (U5573, R2027_U60, U2378);
  nand ginst6230 (U5574, R2278_U101, U2377);
  nand ginst6231 (U5575, ADD_405_U5, U2375);
  nand ginst6232 (U5576, ADD_515_U71, U2374);
  nand ginst6233 (U5577, REIP_REG_2__SCAN_IN, U2370);
  nand ginst6234 (U5578, INSTADDRPOINTER_REG_2__SCAN_IN, U5552);
  nand ginst6235 (U5579, R2099_U42, U2380);
  nand ginst6236 (U5580, R2027_U57, U2378);
  nand ginst6237 (U5581, R2278_U92, U2377);
  nand ginst6238 (U5582, ADD_405_U93, U2375);
  nand ginst6239 (U5583, ADD_515_U68, U2374);
  nand ginst6240 (U5584, REIP_REG_3__SCAN_IN, U2370);
  nand ginst6241 (U5585, INSTADDRPOINTER_REG_3__SCAN_IN, U5552);
  nand ginst6242 (U5586, R2099_U41, U2380);
  nand ginst6243 (U5587, R2027_U56, U2378);
  nand ginst6244 (U5588, R2278_U89, U2377);
  nand ginst6245 (U5589, ADD_405_U68, U2375);
  nand ginst6246 (U5590, ADD_515_U67, U2374);
  nand ginst6247 (U5591, REIP_REG_4__SCAN_IN, U2370);
  nand ginst6248 (U5592, INSTADDRPOINTER_REG_4__SCAN_IN, U5552);
  nand ginst6249 (U5593, R2099_U40, U2380);
  nand ginst6250 (U5594, R2027_U55, U2378);
  nand ginst6251 (U5595, R2278_U86, U2377);
  nand ginst6252 (U5596, ADD_405_U67, U2375);
  nand ginst6253 (U5597, ADD_515_U66, U2374);
  nand ginst6254 (U5598, REIP_REG_5__SCAN_IN, U2370);
  nand ginst6255 (U5599, INSTADDRPOINTER_REG_5__SCAN_IN, U5552);
  nand ginst6256 (U5600, R2099_U39, U2380);
  nand ginst6257 (U5601, R2027_U54, U2378);
  nand ginst6258 (U5602, R2278_U83, U2377);
  nand ginst6259 (U5603, ADD_405_U66, U2375);
  nand ginst6260 (U5604, ADD_515_U65, U2374);
  nand ginst6261 (U5605, REIP_REG_6__SCAN_IN, U2370);
  nand ginst6262 (U5606, INSTADDRPOINTER_REG_6__SCAN_IN, U5552);
  nand ginst6263 (U5607, R2099_U38, U2380);
  nand ginst6264 (U5608, R2027_U53, U2378);
  nand ginst6265 (U5609, R2278_U80, U2377);
  nand ginst6266 (U5610, ADD_405_U65, U2375);
  nand ginst6267 (U5611, ADD_515_U64, U2374);
  nand ginst6268 (U5612, REIP_REG_7__SCAN_IN, U2370);
  nand ginst6269 (U5613, INSTADDRPOINTER_REG_7__SCAN_IN, U5552);
  nand ginst6270 (U5614, R2099_U37, U2380);
  nand ginst6271 (U5615, R2027_U52, U2378);
  nand ginst6272 (U5616, R2278_U77, U2377);
  nand ginst6273 (U5617, ADD_405_U64, U2375);
  nand ginst6274 (U5618, ADD_515_U63, U2374);
  nand ginst6275 (U5619, REIP_REG_8__SCAN_IN, U2370);
  nand ginst6276 (U5620, INSTADDRPOINTER_REG_8__SCAN_IN, U5552);
  nand ginst6277 (U5621, R2099_U36, U2380);
  nand ginst6278 (U5622, R2027_U51, U2378);
  nand ginst6279 (U5623, R2278_U74, U2377);
  nand ginst6280 (U5624, ADD_405_U63, U2375);
  nand ginst6281 (U5625, ADD_515_U62, U2374);
  nand ginst6282 (U5626, REIP_REG_9__SCAN_IN, U2370);
  nand ginst6283 (U5627, INSTADDRPOINTER_REG_9__SCAN_IN, U5552);
  nand ginst6284 (U5628, R2099_U85, U2380);
  nand ginst6285 (U5629, R2027_U81, U2378);
  nand ginst6286 (U5630, R2278_U160, U2377);
  nand ginst6287 (U5631, ADD_405_U91, U2375);
  nand ginst6288 (U5632, ADD_515_U91, U2374);
  nand ginst6289 (U5633, REIP_REG_10__SCAN_IN, U2370);
  nand ginst6290 (U5634, INSTADDRPOINTER_REG_10__SCAN_IN, U5552);
  nand ginst6291 (U5635, R2099_U84, U2380);
  nand ginst6292 (U5636, R2027_U80, U2378);
  nand ginst6293 (U5637, R2278_U157, U2377);
  nand ginst6294 (U5638, ADD_405_U90, U2375);
  nand ginst6295 (U5639, ADD_515_U90, U2374);
  nand ginst6296 (U5640, REIP_REG_11__SCAN_IN, U2370);
  nand ginst6297 (U5641, INSTADDRPOINTER_REG_11__SCAN_IN, U5552);
  nand ginst6298 (U5642, R2099_U83, U2380);
  nand ginst6299 (U5643, R2027_U79, U2378);
  nand ginst6300 (U5644, R2278_U154, U2377);
  nand ginst6301 (U5645, ADD_405_U89, U2375);
  nand ginst6302 (U5646, ADD_515_U89, U2374);
  nand ginst6303 (U5647, REIP_REG_12__SCAN_IN, U2370);
  nand ginst6304 (U5648, INSTADDRPOINTER_REG_12__SCAN_IN, U5552);
  nand ginst6305 (U5649, R2099_U82, U2380);
  nand ginst6306 (U5650, R2027_U78, U2378);
  nand ginst6307 (U5651, R2278_U151, U2377);
  nand ginst6308 (U5652, ADD_405_U88, U2375);
  nand ginst6309 (U5653, ADD_515_U88, U2374);
  nand ginst6310 (U5654, REIP_REG_13__SCAN_IN, U2370);
  nand ginst6311 (U5655, INSTADDRPOINTER_REG_13__SCAN_IN, U5552);
  nand ginst6312 (U5656, R2099_U81, U2380);
  nand ginst6313 (U5657, R2027_U77, U2378);
  nand ginst6314 (U5658, R2278_U148, U2377);
  nand ginst6315 (U5659, ADD_405_U87, U2375);
  nand ginst6316 (U5660, ADD_515_U87, U2374);
  nand ginst6317 (U5661, REIP_REG_14__SCAN_IN, U2370);
  nand ginst6318 (U5662, INSTADDRPOINTER_REG_14__SCAN_IN, U5552);
  nand ginst6319 (U5663, R2099_U80, U2380);
  nand ginst6320 (U5664, R2027_U76, U2378);
  nand ginst6321 (U5665, R2278_U145, U2377);
  nand ginst6322 (U5666, ADD_405_U86, U2375);
  nand ginst6323 (U5667, ADD_515_U86, U2374);
  nand ginst6324 (U5668, REIP_REG_15__SCAN_IN, U2370);
  nand ginst6325 (U5669, INSTADDRPOINTER_REG_15__SCAN_IN, U5552);
  nand ginst6326 (U5670, R2099_U79, U2380);
  nand ginst6327 (U5671, R2027_U75, U2378);
  nand ginst6328 (U5672, R2278_U142, U2377);
  nand ginst6329 (U5673, ADD_405_U85, U2375);
  nand ginst6330 (U5674, ADD_515_U85, U2374);
  nand ginst6331 (U5675, REIP_REG_16__SCAN_IN, U2370);
  nand ginst6332 (U5676, INSTADDRPOINTER_REG_16__SCAN_IN, U5552);
  nand ginst6333 (U5677, R2099_U78, U2380);
  nand ginst6334 (U5678, R2027_U74, U2378);
  nand ginst6335 (U5679, R2278_U139, U2377);
  nand ginst6336 (U5680, ADD_405_U84, U2375);
  nand ginst6337 (U5681, ADD_515_U84, U2374);
  nand ginst6338 (U5682, REIP_REG_17__SCAN_IN, U2370);
  nand ginst6339 (U5683, INSTADDRPOINTER_REG_17__SCAN_IN, U5552);
  nand ginst6340 (U5684, R2099_U77, U2380);
  nand ginst6341 (U5685, R2027_U73, U2378);
  nand ginst6342 (U5686, R2278_U136, U2377);
  nand ginst6343 (U5687, ADD_405_U83, U2375);
  nand ginst6344 (U5688, ADD_515_U83, U2374);
  nand ginst6345 (U5689, REIP_REG_18__SCAN_IN, U2370);
  nand ginst6346 (U5690, INSTADDRPOINTER_REG_18__SCAN_IN, U5552);
  nand ginst6347 (U5691, R2099_U76, U2380);
  nand ginst6348 (U5692, R2027_U72, U2378);
  nand ginst6349 (U5693, R2278_U133, U2377);
  nand ginst6350 (U5694, ADD_405_U82, U2375);
  nand ginst6351 (U5695, ADD_515_U82, U2374);
  nand ginst6352 (U5696, REIP_REG_19__SCAN_IN, U2370);
  nand ginst6353 (U5697, INSTADDRPOINTER_REG_19__SCAN_IN, U5552);
  nand ginst6354 (U5698, R2099_U75, U2380);
  nand ginst6355 (U5699, R2027_U70, U2378);
  nand ginst6356 (U5700, R2278_U129, U2377);
  nand ginst6357 (U5701, ADD_405_U80, U2375);
  nand ginst6358 (U5702, ADD_515_U81, U2374);
  nand ginst6359 (U5703, REIP_REG_20__SCAN_IN, U2370);
  nand ginst6360 (U5704, INSTADDRPOINTER_REG_20__SCAN_IN, U5552);
  nand ginst6361 (U5705, R2099_U74, U2380);
  nand ginst6362 (U5706, R2027_U69, U2378);
  nand ginst6363 (U5707, R2278_U126, U2377);
  nand ginst6364 (U5708, ADD_405_U79, U2375);
  nand ginst6365 (U5709, ADD_515_U80, U2374);
  nand ginst6366 (U5710, REIP_REG_21__SCAN_IN, U2370);
  nand ginst6367 (U5711, INSTADDRPOINTER_REG_21__SCAN_IN, U5552);
  nand ginst6368 (U5712, R2099_U73, U2380);
  nand ginst6369 (U5713, R2027_U68, U2378);
  nand ginst6370 (U5714, R2278_U123, U2377);
  nand ginst6371 (U5715, ADD_405_U78, U2375);
  nand ginst6372 (U5716, ADD_515_U79, U2374);
  nand ginst6373 (U5717, REIP_REG_22__SCAN_IN, U2370);
  nand ginst6374 (U5718, INSTADDRPOINTER_REG_22__SCAN_IN, U5552);
  nand ginst6375 (U5719, R2099_U72, U2380);
  nand ginst6376 (U5720, R2027_U67, U2378);
  nand ginst6377 (U5721, R2278_U120, U2377);
  nand ginst6378 (U5722, ADD_405_U77, U2375);
  nand ginst6379 (U5723, ADD_515_U78, U2374);
  nand ginst6380 (U5724, REIP_REG_23__SCAN_IN, U2370);
  nand ginst6381 (U5725, INSTADDRPOINTER_REG_23__SCAN_IN, U5552);
  nand ginst6382 (U5726, R2099_U71, U2380);
  nand ginst6383 (U5727, R2027_U66, U2378);
  nand ginst6384 (U5728, R2278_U117, U2377);
  nand ginst6385 (U5729, ADD_405_U76, U2375);
  nand ginst6386 (U5730, ADD_515_U77, U2374);
  nand ginst6387 (U5731, REIP_REG_24__SCAN_IN, U2370);
  nand ginst6388 (U5732, INSTADDRPOINTER_REG_24__SCAN_IN, U5552);
  nand ginst6389 (U5733, R2099_U70, U2380);
  nand ginst6390 (U5734, R2027_U65, U2378);
  nand ginst6391 (U5735, R2278_U114, U2377);
  nand ginst6392 (U5736, ADD_405_U75, U2375);
  nand ginst6393 (U5737, ADD_515_U76, U2374);
  nand ginst6394 (U5738, REIP_REG_25__SCAN_IN, U2370);
  nand ginst6395 (U5739, INSTADDRPOINTER_REG_25__SCAN_IN, U5552);
  nand ginst6396 (U5740, R2099_U69, U2380);
  nand ginst6397 (U5741, R2027_U64, U2378);
  nand ginst6398 (U5742, R2278_U111, U2377);
  nand ginst6399 (U5743, ADD_405_U74, U2375);
  nand ginst6400 (U5744, ADD_515_U75, U2374);
  nand ginst6401 (U5745, REIP_REG_26__SCAN_IN, U2370);
  nand ginst6402 (U5746, INSTADDRPOINTER_REG_26__SCAN_IN, U5552);
  nand ginst6403 (U5747, R2099_U68, U2380);
  nand ginst6404 (U5748, R2027_U63, U2378);
  nand ginst6405 (U5749, R2278_U108, U2377);
  nand ginst6406 (U5750, ADD_405_U73, U2375);
  nand ginst6407 (U5751, ADD_515_U74, U2374);
  nand ginst6408 (U5752, REIP_REG_27__SCAN_IN, U2370);
  nand ginst6409 (U5753, INSTADDRPOINTER_REG_27__SCAN_IN, U5552);
  nand ginst6410 (U5754, R2099_U67, U2380);
  nand ginst6411 (U5755, R2027_U62, U2378);
  nand ginst6412 (U5756, R2278_U105, U2377);
  nand ginst6413 (U5757, ADD_405_U72, U2375);
  nand ginst6414 (U5758, ADD_515_U73, U2374);
  nand ginst6415 (U5759, REIP_REG_28__SCAN_IN, U2370);
  nand ginst6416 (U5760, INSTADDRPOINTER_REG_28__SCAN_IN, U5552);
  nand ginst6417 (U5761, R2099_U66, U2380);
  nand ginst6418 (U5762, R2027_U61, U2378);
  nand ginst6419 (U5763, R2278_U103, U2377);
  nand ginst6420 (U5764, ADD_405_U71, U2375);
  nand ginst6421 (U5765, ADD_515_U72, U2374);
  nand ginst6422 (U5766, REIP_REG_29__SCAN_IN, U2370);
  nand ginst6423 (U5767, INSTADDRPOINTER_REG_29__SCAN_IN, U5552);
  nand ginst6424 (U5768, R2099_U65, U2380);
  nand ginst6425 (U5769, R2027_U59, U2378);
  nand ginst6426 (U5770, R2278_U98, U2377);
  nand ginst6427 (U5771, ADD_405_U70, U2375);
  nand ginst6428 (U5772, ADD_515_U70, U2374);
  nand ginst6429 (U5773, REIP_REG_30__SCAN_IN, U2370);
  nand ginst6430 (U5774, INSTADDRPOINTER_REG_30__SCAN_IN, U5552);
  nand ginst6431 (U5775, R2099_U64, U2380);
  nand ginst6432 (U5776, R2027_U58, U2378);
  nand ginst6433 (U5777, R2278_U96, U2377);
  nand ginst6434 (U5778, ADD_405_U69, U2375);
  nand ginst6435 (U5779, ADD_515_U69, U2374);
  nand ginst6436 (U5780, REIP_REG_31__SCAN_IN, U2370);
  nand ginst6437 (U5781, INSTADDRPOINTER_REG_31__SCAN_IN, U5552);
  nand ginst6438 (U5782, U3281, U4197);
  not ginst6439 (U5783, U3403);
  nand ginst6440 (U5784, STATE2_REG_2__SCAN_IN, U3281);
  nand ginst6441 (U5785, STATE2_REG_1__SCAN_IN, U3295);
  nand ginst6442 (U5786, U5784, U5785);
  nand ginst6443 (U5787, PHYADDRPOINTER_REG_0__SCAN_IN, U2376);
  nand ginst6444 (U5788, R2278_U17, U2372);
  nand ginst6445 (U5789, REIP_REG_0__SCAN_IN, U2365);
  nand ginst6446 (U5790, R2358_U82, U2364);
  nand ginst6447 (U5791, PHYADDRPOINTER_REG_0__SCAN_IN, U5783);
  nand ginst6448 (U5792, R2337_U5, U2376);
  nand ginst6449 (U5793, R2278_U42, U2372);
  nand ginst6450 (U5794, REIP_REG_1__SCAN_IN, U2365);
  nand ginst6451 (U5795, R2358_U112, U2364);
  nand ginst6452 (U5796, PHYADDRPOINTER_REG_1__SCAN_IN, U5783);
  nand ginst6453 (U5797, R2337_U60, U2376);
  nand ginst6454 (U5798, R2278_U101, U2372);
  nand ginst6455 (U5799, REIP_REG_2__SCAN_IN, U2365);
  nand ginst6456 (U5800, R2358_U19, U2364);
  nand ginst6457 (U5801, PHYADDRPOINTER_REG_2__SCAN_IN, U5783);
  nand ginst6458 (U5802, R2337_U57, U2376);
  nand ginst6459 (U5803, R2278_U92, U2372);
  nand ginst6460 (U5804, REIP_REG_3__SCAN_IN, U2365);
  nand ginst6461 (U5805, R2358_U20, U2364);
  nand ginst6462 (U5806, PHYADDRPOINTER_REG_3__SCAN_IN, U5783);
  nand ginst6463 (U5807, R2337_U56, U2376);
  nand ginst6464 (U5808, R2278_U89, U2372);
  nand ginst6465 (U5809, REIP_REG_4__SCAN_IN, U2365);
  nand ginst6466 (U5810, R2358_U90, U2364);
  nand ginst6467 (U5811, PHYADDRPOINTER_REG_4__SCAN_IN, U5783);
  nand ginst6468 (U5812, R2337_U55, U2376);
  nand ginst6469 (U5813, R2278_U86, U2372);
  nand ginst6470 (U5814, REIP_REG_5__SCAN_IN, U2365);
  nand ginst6471 (U5815, R2358_U88, U2364);
  nand ginst6472 (U5816, PHYADDRPOINTER_REG_5__SCAN_IN, U5783);
  nand ginst6473 (U5817, R2337_U54, U2376);
  nand ginst6474 (U5818, R2278_U83, U2372);
  nand ginst6475 (U5819, REIP_REG_6__SCAN_IN, U2365);
  nand ginst6476 (U5820, R2358_U86, U2364);
  nand ginst6477 (U5821, PHYADDRPOINTER_REG_6__SCAN_IN, U5783);
  nand ginst6478 (U5822, R2337_U53, U2376);
  nand ginst6479 (U5823, R2278_U80, U2372);
  nand ginst6480 (U5824, REIP_REG_7__SCAN_IN, U2365);
  nand ginst6481 (U5825, R2358_U21, U2364);
  nand ginst6482 (U5826, PHYADDRPOINTER_REG_7__SCAN_IN, U5783);
  nand ginst6483 (U5827, R2337_U52, U2376);
  nand ginst6484 (U5828, R2278_U77, U2372);
  nand ginst6485 (U5829, REIP_REG_8__SCAN_IN, U2365);
  nand ginst6486 (U5830, R2358_U85, U2364);
  nand ginst6487 (U5831, PHYADDRPOINTER_REG_8__SCAN_IN, U5783);
  nand ginst6488 (U5832, R2337_U51, U2376);
  nand ginst6489 (U5833, R2278_U74, U2372);
  nand ginst6490 (U5834, REIP_REG_9__SCAN_IN, U2365);
  nand ginst6491 (U5835, R2358_U83, U2364);
  nand ginst6492 (U5836, PHYADDRPOINTER_REG_9__SCAN_IN, U5783);
  nand ginst6493 (U5837, R2337_U80, U2376);
  nand ginst6494 (U5838, R2278_U160, U2372);
  nand ginst6495 (U5839, REIP_REG_10__SCAN_IN, U2365);
  nand ginst6496 (U5840, R2358_U14, U2364);
  nand ginst6497 (U5841, PHYADDRPOINTER_REG_10__SCAN_IN, U5783);
  nand ginst6498 (U5842, R2337_U79, U2376);
  nand ginst6499 (U5843, R2278_U157, U2372);
  nand ginst6500 (U5844, REIP_REG_11__SCAN_IN, U2365);
  nand ginst6501 (U5845, R2358_U15, U2364);
  nand ginst6502 (U5846, PHYADDRPOINTER_REG_11__SCAN_IN, U5783);
  nand ginst6503 (U5847, R2337_U78, U2376);
  nand ginst6504 (U5848, R2278_U154, U2372);
  nand ginst6505 (U5849, REIP_REG_12__SCAN_IN, U2365);
  nand ginst6506 (U5850, R2358_U122, U2364);
  nand ginst6507 (U5851, PHYADDRPOINTER_REG_12__SCAN_IN, U5783);
  nand ginst6508 (U5852, R2337_U77, U2376);
  nand ginst6509 (U5853, R2278_U151, U2372);
  nand ginst6510 (U5854, REIP_REG_13__SCAN_IN, U2365);
  nand ginst6511 (U5855, R2358_U120, U2364);
  nand ginst6512 (U5856, PHYADDRPOINTER_REG_13__SCAN_IN, U5783);
  nand ginst6513 (U5857, R2337_U76, U2376);
  nand ginst6514 (U5858, R2278_U148, U2372);
  nand ginst6515 (U5859, REIP_REG_14__SCAN_IN, U2365);
  nand ginst6516 (U5860, R2358_U119, U2364);
  nand ginst6517 (U5861, PHYADDRPOINTER_REG_14__SCAN_IN, U5783);
  nand ginst6518 (U5862, R2337_U75, U2376);
  nand ginst6519 (U5863, R2278_U145, U2372);
  nand ginst6520 (U5864, REIP_REG_15__SCAN_IN, U2365);
  nand ginst6521 (U5865, R2358_U16, U2364);
  nand ginst6522 (U5866, PHYADDRPOINTER_REG_15__SCAN_IN, U5783);
  nand ginst6523 (U5867, R2337_U74, U2376);
  nand ginst6524 (U5868, R2278_U142, U2372);
  nand ginst6525 (U5869, REIP_REG_16__SCAN_IN, U2365);
  nand ginst6526 (U5870, R2358_U17, U2364);
  nand ginst6527 (U5871, PHYADDRPOINTER_REG_16__SCAN_IN, U5783);
  nand ginst6528 (U5872, R2337_U73, U2376);
  nand ginst6529 (U5873, R2278_U139, U2372);
  nand ginst6530 (U5874, REIP_REG_17__SCAN_IN, U2365);
  nand ginst6531 (U5875, R2358_U118, U2364);
  nand ginst6532 (U5876, PHYADDRPOINTER_REG_17__SCAN_IN, U5783);
  nand ginst6533 (U5877, R2337_U72, U2376);
  nand ginst6534 (U5878, R2278_U136, U2372);
  nand ginst6535 (U5879, REIP_REG_18__SCAN_IN, U2365);
  nand ginst6536 (U5880, R2358_U116, U2364);
  nand ginst6537 (U5881, PHYADDRPOINTER_REG_18__SCAN_IN, U5783);
  nand ginst6538 (U5882, R2337_U71, U2376);
  nand ginst6539 (U5883, R2278_U133, U2372);
  nand ginst6540 (U5884, REIP_REG_19__SCAN_IN, U2365);
  nand ginst6541 (U5885, R2358_U114, U2364);
  nand ginst6542 (U5886, PHYADDRPOINTER_REG_19__SCAN_IN, U5783);
  nand ginst6543 (U5887, R2337_U70, U2376);
  nand ginst6544 (U5888, R2278_U129, U2372);
  nand ginst6545 (U5889, REIP_REG_20__SCAN_IN, U2365);
  nand ginst6546 (U5890, R2358_U110, U2364);
  nand ginst6547 (U5891, PHYADDRPOINTER_REG_20__SCAN_IN, U5783);
  nand ginst6548 (U5892, R2337_U69, U2376);
  nand ginst6549 (U5893, R2278_U126, U2372);
  nand ginst6550 (U5894, REIP_REG_21__SCAN_IN, U2365);
  nand ginst6551 (U5895, R2358_U18, U2364);
  nand ginst6552 (U5896, PHYADDRPOINTER_REG_21__SCAN_IN, U5783);
  nand ginst6553 (U5897, R2337_U68, U2376);
  nand ginst6554 (U5898, R2278_U123, U2372);
  nand ginst6555 (U5899, REIP_REG_22__SCAN_IN, U2365);
  nand ginst6556 (U5900, R2358_U109, U2364);
  nand ginst6557 (U5901, PHYADDRPOINTER_REG_22__SCAN_IN, U5783);
  nand ginst6558 (U5902, R2337_U67, U2376);
  nand ginst6559 (U5903, R2278_U120, U2372);
  nand ginst6560 (U5904, REIP_REG_23__SCAN_IN, U2365);
  nand ginst6561 (U5905, R2358_U107, U2364);
  nand ginst6562 (U5906, PHYADDRPOINTER_REG_23__SCAN_IN, U5783);
  nand ginst6563 (U5907, R2337_U66, U2376);
  nand ginst6564 (U5908, R2278_U117, U2372);
  nand ginst6565 (U5909, REIP_REG_24__SCAN_IN, U2365);
  nand ginst6566 (U5910, R2358_U105, U2364);
  nand ginst6567 (U5911, PHYADDRPOINTER_REG_24__SCAN_IN, U5783);
  nand ginst6568 (U5912, R2337_U65, U2376);
  nand ginst6569 (U5913, R2278_U114, U2372);
  nand ginst6570 (U5914, REIP_REG_25__SCAN_IN, U2365);
  nand ginst6571 (U5915, R2358_U103, U2364);
  nand ginst6572 (U5916, PHYADDRPOINTER_REG_25__SCAN_IN, U5783);
  nand ginst6573 (U5917, R2337_U64, U2376);
  nand ginst6574 (U5918, R2278_U111, U2372);
  nand ginst6575 (U5919, REIP_REG_26__SCAN_IN, U2365);
  nand ginst6576 (U5920, R2358_U101, U2364);
  nand ginst6577 (U5921, PHYADDRPOINTER_REG_26__SCAN_IN, U5783);
  nand ginst6578 (U5922, R2337_U63, U2376);
  nand ginst6579 (U5923, R2278_U108, U2372);
  nand ginst6580 (U5924, REIP_REG_27__SCAN_IN, U2365);
  nand ginst6581 (U5925, R2358_U99, U2364);
  nand ginst6582 (U5926, PHYADDRPOINTER_REG_27__SCAN_IN, U5783);
  nand ginst6583 (U5927, R2337_U62, U2376);
  nand ginst6584 (U5928, R2278_U105, U2372);
  nand ginst6585 (U5929, REIP_REG_28__SCAN_IN, U2365);
  nand ginst6586 (U5930, R2358_U97, U2364);
  nand ginst6587 (U5931, PHYADDRPOINTER_REG_28__SCAN_IN, U5783);
  nand ginst6588 (U5932, R2337_U61, U2376);
  nand ginst6589 (U5933, R2278_U103, U2372);
  nand ginst6590 (U5934, REIP_REG_29__SCAN_IN, U2365);
  nand ginst6591 (U5935, R2358_U95, U2364);
  nand ginst6592 (U5936, PHYADDRPOINTER_REG_29__SCAN_IN, U5783);
  nand ginst6593 (U5937, R2337_U59, U2376);
  nand ginst6594 (U5938, R2278_U98, U2372);
  nand ginst6595 (U5939, REIP_REG_30__SCAN_IN, U2365);
  nand ginst6596 (U5940, R2358_U93, U2364);
  nand ginst6597 (U5941, PHYADDRPOINTER_REG_30__SCAN_IN, U5783);
  nand ginst6598 (U5942, R2337_U58, U2376);
  nand ginst6599 (U5943, R2278_U96, U2372);
  nand ginst6600 (U5944, REIP_REG_31__SCAN_IN, U2365);
  nand ginst6601 (U5945, R2358_U91, U2364);
  nand ginst6602 (U5946, PHYADDRPOINTER_REG_31__SCAN_IN, U5783);
  nand ginst6603 (U5947, READY_N, U3269);
  nand ginst6604 (U5948, EAX_REG_15__SCAN_IN, U2382);
  nand ginst6605 (U5949, DATAI_15_, U2381);
  nand ginst6606 (U5950, U5948, U5949);
  nand ginst6607 (U5951, EAX_REG_14__SCAN_IN, U2382);
  nand ginst6608 (U5952, DATAI_14_, U2381);
  nand ginst6609 (U5953, U5951, U5952);
  nand ginst6610 (U5954, EAX_REG_13__SCAN_IN, U2382);
  nand ginst6611 (U5955, DATAI_13_, U2381);
  nand ginst6612 (U5956, U5954, U5955);
  nand ginst6613 (U5957, EAX_REG_12__SCAN_IN, U2382);
  nand ginst6614 (U5958, DATAI_12_, U2381);
  nand ginst6615 (U5959, U5957, U5958);
  nand ginst6616 (U5960, EAX_REG_11__SCAN_IN, U2382);
  nand ginst6617 (U5961, DATAI_11_, U2381);
  nand ginst6618 (U5962, U5960, U5961);
  nand ginst6619 (U5963, EAX_REG_10__SCAN_IN, U2382);
  nand ginst6620 (U5964, DATAI_10_, U2381);
  nand ginst6621 (U5965, U5963, U5964);
  nand ginst6622 (U5966, EAX_REG_9__SCAN_IN, U2382);
  nand ginst6623 (U5967, DATAI_9_, U2381);
  nand ginst6624 (U5968, U5966, U5967);
  nand ginst6625 (U5969, EAX_REG_8__SCAN_IN, U2382);
  nand ginst6626 (U5970, DATAI_8_, U2381);
  nand ginst6627 (U5971, U5969, U5970);
  nand ginst6628 (U5972, EAX_REG_7__SCAN_IN, U2382);
  nand ginst6629 (U5973, DATAI_7_, U2381);
  nand ginst6630 (U5974, U5972, U5973);
  nand ginst6631 (U5975, EAX_REG_6__SCAN_IN, U2382);
  nand ginst6632 (U5976, DATAI_6_, U2381);
  nand ginst6633 (U5977, U5975, U5976);
  nand ginst6634 (U5978, EAX_REG_5__SCAN_IN, U2382);
  nand ginst6635 (U5979, DATAI_5_, U2381);
  nand ginst6636 (U5980, U5978, U5979);
  nand ginst6637 (U5981, EAX_REG_4__SCAN_IN, U2382);
  nand ginst6638 (U5982, DATAI_4_, U2381);
  nand ginst6639 (U5983, U5981, U5982);
  nand ginst6640 (U5984, EAX_REG_3__SCAN_IN, U2382);
  nand ginst6641 (U5985, DATAI_3_, U2381);
  nand ginst6642 (U5986, U5984, U5985);
  nand ginst6643 (U5987, EAX_REG_2__SCAN_IN, U2382);
  nand ginst6644 (U5988, DATAI_2_, U2381);
  nand ginst6645 (U5989, U5987, U5988);
  nand ginst6646 (U5990, EAX_REG_1__SCAN_IN, U2382);
  nand ginst6647 (U5991, DATAI_1_, U2381);
  nand ginst6648 (U5992, U5990, U5991);
  nand ginst6649 (U5993, EAX_REG_0__SCAN_IN, U2382);
  nand ginst6650 (U5994, DATAI_0_, U2381);
  nand ginst6651 (U5995, U5993, U5994);
  nand ginst6652 (U5996, EAX_REG_30__SCAN_IN, U2382);
  nand ginst6653 (U5997, DATAI_14_, U2381);
  nand ginst6654 (U5998, U5996, U5997);
  nand ginst6655 (U5999, EAX_REG_29__SCAN_IN, U2382);
  nand ginst6656 (U6000, DATAI_13_, U2381);
  nand ginst6657 (U6001, U5999, U6000);
  nand ginst6658 (U6002, EAX_REG_28__SCAN_IN, U2382);
  nand ginst6659 (U6003, DATAI_12_, U2381);
  nand ginst6660 (U6004, U6002, U6003);
  nand ginst6661 (U6005, EAX_REG_27__SCAN_IN, U2382);
  nand ginst6662 (U6006, DATAI_11_, U2381);
  nand ginst6663 (U6007, U6005, U6006);
  nand ginst6664 (U6008, EAX_REG_26__SCAN_IN, U2382);
  nand ginst6665 (U6009, DATAI_10_, U2381);
  nand ginst6666 (U6010, U6008, U6009);
  nand ginst6667 (U6011, EAX_REG_25__SCAN_IN, U2382);
  nand ginst6668 (U6012, DATAI_9_, U2381);
  nand ginst6669 (U6013, U6011, U6012);
  nand ginst6670 (U6014, EAX_REG_24__SCAN_IN, U2382);
  nand ginst6671 (U6015, DATAI_8_, U2381);
  nand ginst6672 (U6016, U6014, U6015);
  nand ginst6673 (U6017, EAX_REG_23__SCAN_IN, U2382);
  nand ginst6674 (U6018, DATAI_7_, U2381);
  nand ginst6675 (U6019, U6017, U6018);
  nand ginst6676 (U6020, EAX_REG_22__SCAN_IN, U2382);
  nand ginst6677 (U6021, DATAI_6_, U2381);
  nand ginst6678 (U6022, U6020, U6021);
  nand ginst6679 (U6023, EAX_REG_21__SCAN_IN, U2382);
  nand ginst6680 (U6024, DATAI_5_, U2381);
  nand ginst6681 (U6025, U6023, U6024);
  nand ginst6682 (U6026, EAX_REG_20__SCAN_IN, U2382);
  nand ginst6683 (U6027, DATAI_4_, U2381);
  nand ginst6684 (U6028, U6026, U6027);
  nand ginst6685 (U6029, EAX_REG_19__SCAN_IN, U2382);
  nand ginst6686 (U6030, DATAI_3_, U2381);
  nand ginst6687 (U6031, U6029, U6030);
  nand ginst6688 (U6032, EAX_REG_18__SCAN_IN, U2382);
  nand ginst6689 (U6033, DATAI_2_, U2381);
  nand ginst6690 (U6034, U6032, U6033);
  nand ginst6691 (U6035, EAX_REG_17__SCAN_IN, U2382);
  nand ginst6692 (U6036, DATAI_1_, U2381);
  nand ginst6693 (U6037, U6035, U6036);
  nand ginst6694 (U6038, EAX_REG_16__SCAN_IN, U2382);
  nand ginst6695 (U6039, DATAI_0_, U2381);
  nand ginst6696 (U6040, U6038, U6039);
  nand ginst6697 (U6041, U4223, U4247, U7594);
  nand ginst6698 (U6042, U2428, U3281);
  not ginst6699 (U6043, U3404);
  nand ginst6700 (U6044, LWORD_REG_0__SCAN_IN, U2385);
  nand ginst6701 (U6045, EAX_REG_0__SCAN_IN, U2384);
  nand ginst6702 (U6046, DATAO_REG_0__SCAN_IN, U6043);
  nand ginst6703 (U6047, LWORD_REG_1__SCAN_IN, U2385);
  nand ginst6704 (U6048, EAX_REG_1__SCAN_IN, U2384);
  nand ginst6705 (U6049, DATAO_REG_1__SCAN_IN, U6043);
  nand ginst6706 (U6050, LWORD_REG_2__SCAN_IN, U2385);
  nand ginst6707 (U6051, EAX_REG_2__SCAN_IN, U2384);
  nand ginst6708 (U6052, DATAO_REG_2__SCAN_IN, U6043);
  nand ginst6709 (U6053, LWORD_REG_3__SCAN_IN, U2385);
  nand ginst6710 (U6054, EAX_REG_3__SCAN_IN, U2384);
  nand ginst6711 (U6055, DATAO_REG_3__SCAN_IN, U6043);
  nand ginst6712 (U6056, LWORD_REG_4__SCAN_IN, U2385);
  nand ginst6713 (U6057, EAX_REG_4__SCAN_IN, U2384);
  nand ginst6714 (U6058, DATAO_REG_4__SCAN_IN, U6043);
  nand ginst6715 (U6059, LWORD_REG_5__SCAN_IN, U2385);
  nand ginst6716 (U6060, EAX_REG_5__SCAN_IN, U2384);
  nand ginst6717 (U6061, DATAO_REG_5__SCAN_IN, U6043);
  nand ginst6718 (U6062, LWORD_REG_6__SCAN_IN, U2385);
  nand ginst6719 (U6063, EAX_REG_6__SCAN_IN, U2384);
  nand ginst6720 (U6064, DATAO_REG_6__SCAN_IN, U6043);
  nand ginst6721 (U6065, LWORD_REG_7__SCAN_IN, U2385);
  nand ginst6722 (U6066, EAX_REG_7__SCAN_IN, U2384);
  nand ginst6723 (U6067, DATAO_REG_7__SCAN_IN, U6043);
  nand ginst6724 (U6068, LWORD_REG_8__SCAN_IN, U2385);
  nand ginst6725 (U6069, EAX_REG_8__SCAN_IN, U2384);
  nand ginst6726 (U6070, DATAO_REG_8__SCAN_IN, U6043);
  nand ginst6727 (U6071, LWORD_REG_9__SCAN_IN, U2385);
  nand ginst6728 (U6072, EAX_REG_9__SCAN_IN, U2384);
  nand ginst6729 (U6073, DATAO_REG_9__SCAN_IN, U6043);
  nand ginst6730 (U6074, LWORD_REG_10__SCAN_IN, U2385);
  nand ginst6731 (U6075, EAX_REG_10__SCAN_IN, U2384);
  nand ginst6732 (U6076, DATAO_REG_10__SCAN_IN, U6043);
  nand ginst6733 (U6077, LWORD_REG_11__SCAN_IN, U2385);
  nand ginst6734 (U6078, EAX_REG_11__SCAN_IN, U2384);
  nand ginst6735 (U6079, DATAO_REG_11__SCAN_IN, U6043);
  nand ginst6736 (U6080, LWORD_REG_12__SCAN_IN, U2385);
  nand ginst6737 (U6081, EAX_REG_12__SCAN_IN, U2384);
  nand ginst6738 (U6082, DATAO_REG_12__SCAN_IN, U6043);
  nand ginst6739 (U6083, LWORD_REG_13__SCAN_IN, U2385);
  nand ginst6740 (U6084, EAX_REG_13__SCAN_IN, U2384);
  nand ginst6741 (U6085, DATAO_REG_13__SCAN_IN, U6043);
  nand ginst6742 (U6086, LWORD_REG_14__SCAN_IN, U2385);
  nand ginst6743 (U6087, EAX_REG_14__SCAN_IN, U2384);
  nand ginst6744 (U6088, DATAO_REG_14__SCAN_IN, U6043);
  nand ginst6745 (U6089, LWORD_REG_15__SCAN_IN, U2385);
  nand ginst6746 (U6090, EAX_REG_15__SCAN_IN, U2384);
  nand ginst6747 (U6091, DATAO_REG_15__SCAN_IN, U6043);
  nand ginst6748 (U6092, EAX_REG_16__SCAN_IN, U2424);
  nand ginst6749 (U6093, UWORD_REG_0__SCAN_IN, U2385);
  nand ginst6750 (U6094, DATAO_REG_16__SCAN_IN, U6043);
  nand ginst6751 (U6095, EAX_REG_17__SCAN_IN, U2424);
  nand ginst6752 (U6096, UWORD_REG_1__SCAN_IN, U2385);
  nand ginst6753 (U6097, DATAO_REG_17__SCAN_IN, U6043);
  nand ginst6754 (U6098, EAX_REG_18__SCAN_IN, U2424);
  nand ginst6755 (U6099, UWORD_REG_2__SCAN_IN, U2385);
  nand ginst6756 (U6100, DATAO_REG_18__SCAN_IN, U6043);
  nand ginst6757 (U6101, EAX_REG_19__SCAN_IN, U2424);
  nand ginst6758 (U6102, UWORD_REG_3__SCAN_IN, U2385);
  nand ginst6759 (U6103, DATAO_REG_19__SCAN_IN, U6043);
  nand ginst6760 (U6104, EAX_REG_20__SCAN_IN, U2424);
  nand ginst6761 (U6105, UWORD_REG_4__SCAN_IN, U2385);
  nand ginst6762 (U6106, DATAO_REG_20__SCAN_IN, U6043);
  nand ginst6763 (U6107, EAX_REG_21__SCAN_IN, U2424);
  nand ginst6764 (U6108, UWORD_REG_5__SCAN_IN, U2385);
  nand ginst6765 (U6109, DATAO_REG_21__SCAN_IN, U6043);
  nand ginst6766 (U6110, EAX_REG_22__SCAN_IN, U2424);
  nand ginst6767 (U6111, UWORD_REG_6__SCAN_IN, U2385);
  nand ginst6768 (U6112, DATAO_REG_22__SCAN_IN, U6043);
  nand ginst6769 (U6113, EAX_REG_23__SCAN_IN, U2424);
  nand ginst6770 (U6114, UWORD_REG_7__SCAN_IN, U2385);
  nand ginst6771 (U6115, DATAO_REG_23__SCAN_IN, U6043);
  nand ginst6772 (U6116, EAX_REG_24__SCAN_IN, U2424);
  nand ginst6773 (U6117, UWORD_REG_8__SCAN_IN, U2385);
  nand ginst6774 (U6118, DATAO_REG_24__SCAN_IN, U6043);
  nand ginst6775 (U6119, EAX_REG_25__SCAN_IN, U2424);
  nand ginst6776 (U6120, UWORD_REG_9__SCAN_IN, U2385);
  nand ginst6777 (U6121, DATAO_REG_25__SCAN_IN, U6043);
  nand ginst6778 (U6122, EAX_REG_26__SCAN_IN, U2424);
  nand ginst6779 (U6123, UWORD_REG_10__SCAN_IN, U2385);
  nand ginst6780 (U6124, DATAO_REG_26__SCAN_IN, U6043);
  nand ginst6781 (U6125, EAX_REG_27__SCAN_IN, U2424);
  nand ginst6782 (U6126, UWORD_REG_11__SCAN_IN, U2385);
  nand ginst6783 (U6127, DATAO_REG_27__SCAN_IN, U6043);
  nand ginst6784 (U6128, EAX_REG_28__SCAN_IN, U2424);
  nand ginst6785 (U6129, UWORD_REG_12__SCAN_IN, U2385);
  nand ginst6786 (U6130, DATAO_REG_28__SCAN_IN, U6043);
  nand ginst6787 (U6131, EAX_REG_29__SCAN_IN, U2424);
  nand ginst6788 (U6132, UWORD_REG_13__SCAN_IN, U2385);
  nand ginst6789 (U6133, DATAO_REG_29__SCAN_IN, U6043);
  nand ginst6790 (U6134, EAX_REG_30__SCAN_IN, U2424);
  nand ginst6791 (U6135, UWORD_REG_14__SCAN_IN, U2385);
  nand ginst6792 (U6136, DATAO_REG_30__SCAN_IN, U6043);
  nand ginst6793 (U6137, GTE_485_U6, U2447, U4182);
  nand ginst6794 (U6138, U4182, U4185, U4242);
  nand ginst6795 (U6139, R2167_U17, U3270, U4188);
  nand ginst6796 (U6140, U3244, U7491);
  nand ginst6797 (U6141, U3871, U6140);
  nand ginst6798 (U6142, DATAI_0_, U2422);
  nand ginst6799 (U6143, R2358_U82, U2386);
  nand ginst6800 (U6144, EAX_REG_0__SCAN_IN, U3411);
  nand ginst6801 (U6145, DATAI_1_, U2422);
  nand ginst6802 (U6146, R2358_U112, U2386);
  nand ginst6803 (U6147, EAX_REG_1__SCAN_IN, U3411);
  nand ginst6804 (U6148, DATAI_2_, U2422);
  nand ginst6805 (U6149, R2358_U19, U2386);
  nand ginst6806 (U6150, EAX_REG_2__SCAN_IN, U3411);
  nand ginst6807 (U6151, DATAI_3_, U2422);
  nand ginst6808 (U6152, R2358_U20, U2386);
  nand ginst6809 (U6153, EAX_REG_3__SCAN_IN, U3411);
  nand ginst6810 (U6154, DATAI_4_, U2422);
  nand ginst6811 (U6155, R2358_U90, U2386);
  nand ginst6812 (U6156, EAX_REG_4__SCAN_IN, U3411);
  nand ginst6813 (U6157, DATAI_5_, U2422);
  nand ginst6814 (U6158, R2358_U88, U2386);
  nand ginst6815 (U6159, EAX_REG_5__SCAN_IN, U3411);
  nand ginst6816 (U6160, DATAI_6_, U2422);
  nand ginst6817 (U6161, R2358_U86, U2386);
  nand ginst6818 (U6162, EAX_REG_6__SCAN_IN, U3411);
  nand ginst6819 (U6163, DATAI_7_, U2422);
  nand ginst6820 (U6164, R2358_U21, U2386);
  nand ginst6821 (U6165, EAX_REG_7__SCAN_IN, U3411);
  nand ginst6822 (U6166, DATAI_8_, U2422);
  nand ginst6823 (U6167, R2358_U85, U2386);
  nand ginst6824 (U6168, EAX_REG_8__SCAN_IN, U3411);
  nand ginst6825 (U6169, DATAI_9_, U2422);
  nand ginst6826 (U6170, R2358_U83, U2386);
  nand ginst6827 (U6171, EAX_REG_9__SCAN_IN, U3411);
  nand ginst6828 (U6172, DATAI_10_, U2422);
  nand ginst6829 (U6173, R2358_U14, U2386);
  nand ginst6830 (U6174, EAX_REG_10__SCAN_IN, U3411);
  nand ginst6831 (U6175, DATAI_11_, U2422);
  nand ginst6832 (U6176, R2358_U15, U2386);
  nand ginst6833 (U6177, EAX_REG_11__SCAN_IN, U3411);
  nand ginst6834 (U6178, DATAI_12_, U2422);
  nand ginst6835 (U6179, R2358_U122, U2386);
  nand ginst6836 (U6180, EAX_REG_12__SCAN_IN, U3411);
  nand ginst6837 (U6181, DATAI_13_, U2422);
  nand ginst6838 (U6182, R2358_U120, U2386);
  nand ginst6839 (U6183, EAX_REG_13__SCAN_IN, U3411);
  nand ginst6840 (U6184, DATAI_14_, U2422);
  nand ginst6841 (U6185, R2358_U119, U2386);
  nand ginst6842 (U6186, EAX_REG_14__SCAN_IN, U3411);
  nand ginst6843 (U6187, DATAI_15_, U2422);
  nand ginst6844 (U6188, R2358_U16, U2386);
  nand ginst6845 (U6189, EAX_REG_15__SCAN_IN, U3411);
  nand ginst6846 (U6190, DATAI_16_, U2423);
  nand ginst6847 (U6191, DATAI_0_, U2387);
  nand ginst6848 (U6192, R2358_U17, U2386);
  nand ginst6849 (U6193, EAX_REG_16__SCAN_IN, U3411);
  nand ginst6850 (U6194, DATAI_17_, U2423);
  nand ginst6851 (U6195, DATAI_1_, U2387);
  nand ginst6852 (U6196, R2358_U118, U2386);
  nand ginst6853 (U6197, EAX_REG_17__SCAN_IN, U3411);
  nand ginst6854 (U6198, DATAI_18_, U2423);
  nand ginst6855 (U6199, DATAI_2_, U2387);
  nand ginst6856 (U6200, R2358_U116, U2386);
  nand ginst6857 (U6201, EAX_REG_18__SCAN_IN, U3411);
  nand ginst6858 (U6202, DATAI_19_, U2423);
  nand ginst6859 (U6203, DATAI_3_, U2387);
  nand ginst6860 (U6204, R2358_U114, U2386);
  nand ginst6861 (U6205, EAX_REG_19__SCAN_IN, U3411);
  nand ginst6862 (U6206, DATAI_20_, U2423);
  nand ginst6863 (U6207, DATAI_4_, U2387);
  nand ginst6864 (U6208, R2358_U110, U2386);
  nand ginst6865 (U6209, EAX_REG_20__SCAN_IN, U3411);
  nand ginst6866 (U6210, DATAI_21_, U2423);
  nand ginst6867 (U6211, DATAI_5_, U2387);
  nand ginst6868 (U6212, R2358_U18, U2386);
  nand ginst6869 (U6213, EAX_REG_21__SCAN_IN, U3411);
  nand ginst6870 (U6214, DATAI_22_, U2423);
  nand ginst6871 (U6215, DATAI_6_, U2387);
  nand ginst6872 (U6216, R2358_U109, U2386);
  nand ginst6873 (U6217, EAX_REG_22__SCAN_IN, U3411);
  nand ginst6874 (U6218, DATAI_23_, U2423);
  nand ginst6875 (U6219, DATAI_7_, U2387);
  nand ginst6876 (U6220, R2358_U107, U2386);
  nand ginst6877 (U6221, EAX_REG_23__SCAN_IN, U3411);
  nand ginst6878 (U6222, DATAI_24_, U2423);
  nand ginst6879 (U6223, DATAI_8_, U2387);
  nand ginst6880 (U6224, R2358_U105, U2386);
  nand ginst6881 (U6225, EAX_REG_24__SCAN_IN, U3411);
  nand ginst6882 (U6226, DATAI_25_, U2423);
  nand ginst6883 (U6227, DATAI_9_, U2387);
  nand ginst6884 (U6228, R2358_U103, U2386);
  nand ginst6885 (U6229, EAX_REG_25__SCAN_IN, U3411);
  nand ginst6886 (U6230, DATAI_26_, U2423);
  nand ginst6887 (U6231, DATAI_10_, U2387);
  nand ginst6888 (U6232, R2358_U101, U2386);
  nand ginst6889 (U6233, EAX_REG_26__SCAN_IN, U3411);
  nand ginst6890 (U6234, DATAI_27_, U2423);
  nand ginst6891 (U6235, DATAI_11_, U2387);
  nand ginst6892 (U6236, R2358_U99, U2386);
  nand ginst6893 (U6237, EAX_REG_27__SCAN_IN, U3411);
  nand ginst6894 (U6238, DATAI_28_, U2423);
  nand ginst6895 (U6239, DATAI_12_, U2387);
  nand ginst6896 (U6240, R2358_U97, U2386);
  nand ginst6897 (U6241, EAX_REG_28__SCAN_IN, U3411);
  nand ginst6898 (U6242, DATAI_29_, U2423);
  nand ginst6899 (U6243, DATAI_13_, U2387);
  nand ginst6900 (U6244, R2358_U95, U2386);
  nand ginst6901 (U6245, EAX_REG_29__SCAN_IN, U3411);
  nand ginst6902 (U6246, DATAI_30_, U2423);
  nand ginst6903 (U6247, DATAI_14_, U2387);
  nand ginst6904 (U6248, R2358_U93, U2386);
  nand ginst6905 (U6249, EAX_REG_30__SCAN_IN, U3411);
  nand ginst6906 (U6250, DATAI_31_, U2423);
  nand ginst6907 (U6251, U3260, U4186);
  nand ginst6908 (U6252, U4193, U6251);
  nand ginst6909 (U6253, R2358_U82, U2383);
  nand ginst6910 (U6254, R2099_U86, U2371);
  nand ginst6911 (U6255, EBX_REG_0__SCAN_IN, U3413);
  nand ginst6912 (U6256, R2358_U112, U2383);
  nand ginst6913 (U6257, R2099_U87, U2371);
  nand ginst6914 (U6258, EBX_REG_1__SCAN_IN, U3413);
  nand ginst6915 (U6259, R2358_U19, U2383);
  nand ginst6916 (U6260, R2099_U138, U2371);
  nand ginst6917 (U6261, EBX_REG_2__SCAN_IN, U3413);
  nand ginst6918 (U6262, R2358_U20, U2383);
  nand ginst6919 (U6263, R2099_U42, U2371);
  nand ginst6920 (U6264, EBX_REG_3__SCAN_IN, U3413);
  nand ginst6921 (U6265, R2358_U90, U2383);
  nand ginst6922 (U6266, R2099_U41, U2371);
  nand ginst6923 (U6267, EBX_REG_4__SCAN_IN, U3413);
  nand ginst6924 (U6268, R2358_U88, U2383);
  nand ginst6925 (U6269, R2099_U40, U2371);
  nand ginst6926 (U6270, EBX_REG_5__SCAN_IN, U3413);
  nand ginst6927 (U6271, R2358_U86, U2383);
  nand ginst6928 (U6272, R2099_U39, U2371);
  nand ginst6929 (U6273, EBX_REG_6__SCAN_IN, U3413);
  nand ginst6930 (U6274, R2358_U21, U2383);
  nand ginst6931 (U6275, R2099_U38, U2371);
  nand ginst6932 (U6276, EBX_REG_7__SCAN_IN, U3413);
  nand ginst6933 (U6277, R2358_U85, U2383);
  nand ginst6934 (U6278, R2099_U37, U2371);
  nand ginst6935 (U6279, EBX_REG_8__SCAN_IN, U3413);
  nand ginst6936 (U6280, R2358_U83, U2383);
  nand ginst6937 (U6281, R2099_U36, U2371);
  nand ginst6938 (U6282, EBX_REG_9__SCAN_IN, U3413);
  nand ginst6939 (U6283, R2358_U14, U2383);
  nand ginst6940 (U6284, R2099_U85, U2371);
  nand ginst6941 (U6285, EBX_REG_10__SCAN_IN, U3413);
  nand ginst6942 (U6286, R2358_U15, U2383);
  nand ginst6943 (U6287, R2099_U84, U2371);
  nand ginst6944 (U6288, EBX_REG_11__SCAN_IN, U3413);
  nand ginst6945 (U6289, R2358_U122, U2383);
  nand ginst6946 (U6290, R2099_U83, U2371);
  nand ginst6947 (U6291, EBX_REG_12__SCAN_IN, U3413);
  nand ginst6948 (U6292, R2358_U120, U2383);
  nand ginst6949 (U6293, R2099_U82, U2371);
  nand ginst6950 (U6294, EBX_REG_13__SCAN_IN, U3413);
  nand ginst6951 (U6295, R2358_U119, U2383);
  nand ginst6952 (U6296, R2099_U81, U2371);
  nand ginst6953 (U6297, EBX_REG_14__SCAN_IN, U3413);
  nand ginst6954 (U6298, R2358_U16, U2383);
  nand ginst6955 (U6299, R2099_U80, U2371);
  nand ginst6956 (U6300, EBX_REG_15__SCAN_IN, U3413);
  nand ginst6957 (U6301, R2358_U17, U2383);
  nand ginst6958 (U6302, R2099_U79, U2371);
  nand ginst6959 (U6303, EBX_REG_16__SCAN_IN, U3413);
  nand ginst6960 (U6304, R2358_U118, U2383);
  nand ginst6961 (U6305, R2099_U78, U2371);
  nand ginst6962 (U6306, EBX_REG_17__SCAN_IN, U3413);
  nand ginst6963 (U6307, R2358_U116, U2383);
  nand ginst6964 (U6308, R2099_U77, U2371);
  nand ginst6965 (U6309, EBX_REG_18__SCAN_IN, U3413);
  nand ginst6966 (U6310, R2358_U114, U2383);
  nand ginst6967 (U6311, R2099_U76, U2371);
  nand ginst6968 (U6312, EBX_REG_19__SCAN_IN, U3413);
  nand ginst6969 (U6313, R2358_U110, U2383);
  nand ginst6970 (U6314, R2099_U75, U2371);
  nand ginst6971 (U6315, EBX_REG_20__SCAN_IN, U3413);
  nand ginst6972 (U6316, R2358_U18, U2383);
  nand ginst6973 (U6317, R2099_U74, U2371);
  nand ginst6974 (U6318, EBX_REG_21__SCAN_IN, U3413);
  nand ginst6975 (U6319, R2358_U109, U2383);
  nand ginst6976 (U6320, R2099_U73, U2371);
  nand ginst6977 (U6321, EBX_REG_22__SCAN_IN, U3413);
  nand ginst6978 (U6322, R2358_U107, U2383);
  nand ginst6979 (U6323, R2099_U72, U2371);
  nand ginst6980 (U6324, EBX_REG_23__SCAN_IN, U3413);
  nand ginst6981 (U6325, R2358_U105, U2383);
  nand ginst6982 (U6326, R2099_U71, U2371);
  nand ginst6983 (U6327, EBX_REG_24__SCAN_IN, U3413);
  nand ginst6984 (U6328, R2358_U103, U2383);
  nand ginst6985 (U6329, R2099_U70, U2371);
  nand ginst6986 (U6330, EBX_REG_25__SCAN_IN, U3413);
  nand ginst6987 (U6331, R2358_U101, U2383);
  nand ginst6988 (U6332, R2099_U69, U2371);
  nand ginst6989 (U6333, EBX_REG_26__SCAN_IN, U3413);
  nand ginst6990 (U6334, R2358_U99, U2383);
  nand ginst6991 (U6335, R2099_U68, U2371);
  nand ginst6992 (U6336, EBX_REG_27__SCAN_IN, U3413);
  nand ginst6993 (U6337, R2358_U97, U2383);
  nand ginst6994 (U6338, R2099_U67, U2371);
  nand ginst6995 (U6339, EBX_REG_28__SCAN_IN, U3413);
  nand ginst6996 (U6340, R2358_U95, U2383);
  nand ginst6997 (U6341, R2099_U66, U2371);
  nand ginst6998 (U6342, EBX_REG_29__SCAN_IN, U3413);
  nand ginst6999 (U6343, R2358_U93, U2383);
  nand ginst7000 (U6344, R2099_U65, U2371);
  nand ginst7001 (U6345, EBX_REG_30__SCAN_IN, U3413);
  nand ginst7002 (U6346, R2099_U64, U2371);
  nand ginst7003 (U6347, EBX_REG_31__SCAN_IN, U3413);
  nand ginst7004 (U6348, GTE_485_U6, U4192);
  nand ginst7005 (U6349, R2167_U17, U4190);
  nand ginst7006 (U6350, U3250, U4191);
  not ginst7007 (U6351, U3418);
  nand ginst7008 (U6352, STATE2_REG_2__SCAN_IN, U4237);
  nand ginst7009 (U6353, STATE2_REG_1__SCAN_IN, R2337_U58);
  nand ginst7010 (U6354, U6352, U6353);
  or ginst7011 (U6355, READY_N, STATEBS16_REG_SCAN_IN);
  nand ginst7012 (U6356, R2099_U86, U2604);
  nand ginst7013 (U6357, REIP_REG_0__SCAN_IN, U7473);
  nand ginst7014 (U6358, EBX_REG_0__SCAN_IN, U7472);
  nand ginst7015 (U6359, R2358_U82, U2429);
  nand ginst7016 (U6360, R2182_U34, U2426);
  nand ginst7017 (U6361, PHYADDRPOINTER_REG_0__SCAN_IN, U2373);
  nand ginst7018 (U6362, PHYADDRPOINTER_REG_0__SCAN_IN, U2366);
  nand ginst7019 (U6363, REIP_REG_0__SCAN_IN, U6351);
  nand ginst7020 (U6364, R2099_U87, U2604);
  nand ginst7021 (U6365, R2096_U4, U7473);
  nand ginst7022 (U6366, EBX_REG_1__SCAN_IN, U7472);
  nand ginst7023 (U6367, R2358_U112, U2429);
  nand ginst7024 (U6368, R2182_U33, U2426);
  nand ginst7025 (U6369, PHYADDRPOINTER_REG_1__SCAN_IN, U2373);
  nand ginst7026 (U6370, R2337_U5, U2366);
  nand ginst7027 (U6371, REIP_REG_1__SCAN_IN, U6351);
  nand ginst7028 (U6372, R2099_U138, U2604);
  nand ginst7029 (U6373, R2096_U71, U7473);
  nand ginst7030 (U6374, EBX_REG_2__SCAN_IN, U7472);
  nand ginst7031 (U6375, R2358_U19, U2429);
  nand ginst7032 (U6376, R2182_U42, U2426);
  nand ginst7033 (U6377, PHYADDRPOINTER_REG_2__SCAN_IN, U2373);
  nand ginst7034 (U6378, R2337_U60, U2366);
  nand ginst7035 (U6379, REIP_REG_2__SCAN_IN, U6351);
  nand ginst7036 (U6380, R2099_U42, U2604);
  nand ginst7037 (U6381, R2096_U68, U7473);
  nand ginst7038 (U6382, EBX_REG_3__SCAN_IN, U7472);
  nand ginst7039 (U6383, R2358_U20, U2429);
  nand ginst7040 (U6384, R2182_U25, U2426);
  nand ginst7041 (U6385, PHYADDRPOINTER_REG_3__SCAN_IN, U2373);
  nand ginst7042 (U6386, R2337_U57, U2366);
  nand ginst7043 (U6387, REIP_REG_3__SCAN_IN, U6351);
  nand ginst7044 (U6388, R2099_U41, U2604);
  nand ginst7045 (U6389, R2096_U67, U7473);
  nand ginst7046 (U6390, EBX_REG_4__SCAN_IN, U7472);
  nand ginst7047 (U6391, R2358_U90, U2429);
  nand ginst7048 (U6392, R2182_U24, U2426);
  nand ginst7049 (U6393, PHYADDRPOINTER_REG_4__SCAN_IN, U2373);
  nand ginst7050 (U6394, R2337_U56, U2366);
  nand ginst7051 (U6395, REIP_REG_4__SCAN_IN, U6351);
  nand ginst7052 (U6396, R2099_U40, U2604);
  nand ginst7053 (U6397, R2096_U66, U7473);
  nand ginst7054 (U6398, EBX_REG_5__SCAN_IN, U7472);
  nand ginst7055 (U6399, R2358_U88, U2429);
  nand ginst7056 (U6400, R2182_U5, U2426);
  nand ginst7057 (U6401, PHYADDRPOINTER_REG_5__SCAN_IN, U2373);
  nand ginst7058 (U6402, R2337_U55, U2366);
  nand ginst7059 (U6403, REIP_REG_5__SCAN_IN, U6351);
  nand ginst7060 (U6404, R2099_U39, U2604);
  nand ginst7061 (U6405, R2096_U65, U7473);
  nand ginst7062 (U6406, EBX_REG_6__SCAN_IN, U7472);
  nand ginst7063 (U6407, PHYADDRPOINTER_REG_6__SCAN_IN, U2373);
  nand ginst7064 (U6408, R2358_U86, U2367);
  nand ginst7065 (U6409, R2337_U54, U2366);
  nand ginst7066 (U6410, REIP_REG_6__SCAN_IN, U6351);
  nand ginst7067 (U6411, R2099_U38, U2604);
  nand ginst7068 (U6412, R2096_U64, U7473);
  nand ginst7069 (U6413, EBX_REG_7__SCAN_IN, U7472);
  nand ginst7070 (U6414, PHYADDRPOINTER_REG_7__SCAN_IN, U2373);
  nand ginst7071 (U6415, R2358_U21, U2367);
  nand ginst7072 (U6416, R2337_U53, U2366);
  nand ginst7073 (U6417, REIP_REG_7__SCAN_IN, U6351);
  nand ginst7074 (U6418, R2099_U37, U2604);
  nand ginst7075 (U6419, R2096_U63, U7473);
  nand ginst7076 (U6420, EBX_REG_8__SCAN_IN, U7472);
  nand ginst7077 (U6421, PHYADDRPOINTER_REG_8__SCAN_IN, U2373);
  nand ginst7078 (U6422, R2358_U85, U2367);
  nand ginst7079 (U6423, R2337_U52, U2366);
  nand ginst7080 (U6424, REIP_REG_8__SCAN_IN, U6351);
  nand ginst7081 (U6425, R2099_U36, U2604);
  nand ginst7082 (U6426, R2096_U62, U7473);
  nand ginst7083 (U6427, EBX_REG_9__SCAN_IN, U7472);
  nand ginst7084 (U6428, PHYADDRPOINTER_REG_9__SCAN_IN, U2373);
  nand ginst7085 (U6429, R2358_U83, U2367);
  nand ginst7086 (U6430, R2337_U51, U2366);
  nand ginst7087 (U6431, REIP_REG_9__SCAN_IN, U6351);
  nand ginst7088 (U6432, R2099_U85, U2604);
  nand ginst7089 (U6433, R2096_U91, U7473);
  nand ginst7090 (U6434, EBX_REG_10__SCAN_IN, U7472);
  nand ginst7091 (U6435, PHYADDRPOINTER_REG_10__SCAN_IN, U2373);
  nand ginst7092 (U6436, R2358_U14, U2367);
  nand ginst7093 (U6437, R2337_U80, U2366);
  nand ginst7094 (U6438, REIP_REG_10__SCAN_IN, U6351);
  nand ginst7095 (U6439, R2099_U84, U2604);
  nand ginst7096 (U6440, R2096_U90, U7473);
  nand ginst7097 (U6441, EBX_REG_11__SCAN_IN, U7472);
  nand ginst7098 (U6442, PHYADDRPOINTER_REG_11__SCAN_IN, U2373);
  nand ginst7099 (U6443, R2358_U15, U2367);
  nand ginst7100 (U6444, R2337_U79, U2366);
  nand ginst7101 (U6445, REIP_REG_11__SCAN_IN, U6351);
  nand ginst7102 (U6446, R2099_U83, U2604);
  nand ginst7103 (U6447, R2096_U89, U7473);
  nand ginst7104 (U6448, EBX_REG_12__SCAN_IN, U7472);
  nand ginst7105 (U6449, PHYADDRPOINTER_REG_12__SCAN_IN, U2373);
  nand ginst7106 (U6450, R2358_U122, U2367);
  nand ginst7107 (U6451, R2337_U78, U2366);
  nand ginst7108 (U6452, REIP_REG_12__SCAN_IN, U6351);
  nand ginst7109 (U6453, R2099_U82, U2604);
  nand ginst7110 (U6454, R2096_U88, U7473);
  nand ginst7111 (U6455, EBX_REG_13__SCAN_IN, U7472);
  nand ginst7112 (U6456, PHYADDRPOINTER_REG_13__SCAN_IN, U2373);
  nand ginst7113 (U6457, R2358_U120, U2367);
  nand ginst7114 (U6458, R2337_U77, U2366);
  nand ginst7115 (U6459, REIP_REG_13__SCAN_IN, U6351);
  nand ginst7116 (U6460, R2099_U81, U2604);
  nand ginst7117 (U6461, R2096_U87, U7473);
  nand ginst7118 (U6462, EBX_REG_14__SCAN_IN, U7472);
  nand ginst7119 (U6463, PHYADDRPOINTER_REG_14__SCAN_IN, U2373);
  nand ginst7120 (U6464, R2358_U119, U2367);
  nand ginst7121 (U6465, R2337_U76, U2366);
  nand ginst7122 (U6466, REIP_REG_14__SCAN_IN, U6351);
  nand ginst7123 (U6467, R2099_U80, U2604);
  nand ginst7124 (U6468, R2096_U86, U7473);
  nand ginst7125 (U6469, EBX_REG_15__SCAN_IN, U7472);
  nand ginst7126 (U6470, PHYADDRPOINTER_REG_15__SCAN_IN, U2373);
  nand ginst7127 (U6471, R2358_U16, U2367);
  nand ginst7128 (U6472, R2337_U75, U2366);
  nand ginst7129 (U6473, REIP_REG_15__SCAN_IN, U6351);
  nand ginst7130 (U6474, R2099_U79, U2604);
  nand ginst7131 (U6475, R2096_U85, U7473);
  nand ginst7132 (U6476, EBX_REG_16__SCAN_IN, U7472);
  nand ginst7133 (U6477, PHYADDRPOINTER_REG_16__SCAN_IN, U2373);
  nand ginst7134 (U6478, R2358_U17, U2367);
  nand ginst7135 (U6479, R2337_U74, U2366);
  nand ginst7136 (U6480, REIP_REG_16__SCAN_IN, U6351);
  nand ginst7137 (U6481, R2099_U78, U2604);
  nand ginst7138 (U6482, R2096_U84, U7473);
  nand ginst7139 (U6483, EBX_REG_17__SCAN_IN, U7472);
  nand ginst7140 (U6484, PHYADDRPOINTER_REG_17__SCAN_IN, U2373);
  nand ginst7141 (U6485, R2358_U118, U2367);
  nand ginst7142 (U6486, R2337_U73, U2366);
  nand ginst7143 (U6487, REIP_REG_17__SCAN_IN, U6351);
  nand ginst7144 (U6488, R2099_U77, U2604);
  nand ginst7145 (U6489, R2096_U83, U7473);
  nand ginst7146 (U6490, EBX_REG_18__SCAN_IN, U7472);
  nand ginst7147 (U6491, PHYADDRPOINTER_REG_18__SCAN_IN, U2373);
  nand ginst7148 (U6492, R2358_U116, U2367);
  nand ginst7149 (U6493, R2337_U72, U2366);
  nand ginst7150 (U6494, REIP_REG_18__SCAN_IN, U6351);
  nand ginst7151 (U6495, R2099_U76, U2604);
  nand ginst7152 (U6496, R2096_U82, U7473);
  nand ginst7153 (U6497, EBX_REG_19__SCAN_IN, U7472);
  nand ginst7154 (U6498, PHYADDRPOINTER_REG_19__SCAN_IN, U2373);
  nand ginst7155 (U6499, R2358_U114, U2367);
  nand ginst7156 (U6500, R2337_U71, U2366);
  nand ginst7157 (U6501, REIP_REG_19__SCAN_IN, U6351);
  nand ginst7158 (U6502, R2099_U75, U2604);
  nand ginst7159 (U6503, R2096_U81, U7473);
  nand ginst7160 (U6504, EBX_REG_20__SCAN_IN, U7472);
  nand ginst7161 (U6505, PHYADDRPOINTER_REG_20__SCAN_IN, U2373);
  nand ginst7162 (U6506, R2358_U110, U2367);
  nand ginst7163 (U6507, R2337_U70, U2366);
  nand ginst7164 (U6508, REIP_REG_20__SCAN_IN, U6351);
  nand ginst7165 (U6509, R2099_U74, U2604);
  nand ginst7166 (U6510, R2096_U80, U7473);
  nand ginst7167 (U6511, EBX_REG_21__SCAN_IN, U7472);
  nand ginst7168 (U6512, PHYADDRPOINTER_REG_21__SCAN_IN, U2373);
  nand ginst7169 (U6513, R2358_U18, U2367);
  nand ginst7170 (U6514, R2337_U69, U2366);
  nand ginst7171 (U6515, REIP_REG_21__SCAN_IN, U6351);
  nand ginst7172 (U6516, R2099_U73, U2604);
  nand ginst7173 (U6517, R2096_U79, U7473);
  nand ginst7174 (U6518, EBX_REG_22__SCAN_IN, U7472);
  nand ginst7175 (U6519, PHYADDRPOINTER_REG_22__SCAN_IN, U2373);
  nand ginst7176 (U6520, R2358_U109, U2367);
  nand ginst7177 (U6521, R2337_U68, U2366);
  nand ginst7178 (U6522, REIP_REG_22__SCAN_IN, U6351);
  nand ginst7179 (U6523, R2099_U72, U2604);
  nand ginst7180 (U6524, R2096_U78, U7473);
  nand ginst7181 (U6525, EBX_REG_23__SCAN_IN, U7472);
  nand ginst7182 (U6526, PHYADDRPOINTER_REG_23__SCAN_IN, U2373);
  nand ginst7183 (U6527, R2358_U107, U2367);
  nand ginst7184 (U6528, R2337_U67, U2366);
  nand ginst7185 (U6529, REIP_REG_23__SCAN_IN, U6351);
  nand ginst7186 (U6530, R2099_U71, U2604);
  nand ginst7187 (U6531, R2096_U77, U7473);
  nand ginst7188 (U6532, EBX_REG_24__SCAN_IN, U7472);
  nand ginst7189 (U6533, PHYADDRPOINTER_REG_24__SCAN_IN, U2373);
  nand ginst7190 (U6534, R2358_U105, U2367);
  nand ginst7191 (U6535, R2337_U66, U2366);
  nand ginst7192 (U6536, REIP_REG_24__SCAN_IN, U6351);
  nand ginst7193 (U6537, R2099_U70, U2604);
  nand ginst7194 (U6538, R2096_U76, U7473);
  nand ginst7195 (U6539, EBX_REG_25__SCAN_IN, U7472);
  nand ginst7196 (U6540, PHYADDRPOINTER_REG_25__SCAN_IN, U2373);
  nand ginst7197 (U6541, R2358_U103, U2367);
  nand ginst7198 (U6542, R2337_U65, U2366);
  nand ginst7199 (U6543, REIP_REG_25__SCAN_IN, U6351);
  nand ginst7200 (U6544, R2099_U69, U2604);
  nand ginst7201 (U6545, R2096_U75, U7473);
  nand ginst7202 (U6546, EBX_REG_26__SCAN_IN, U7472);
  nand ginst7203 (U6547, PHYADDRPOINTER_REG_26__SCAN_IN, U2373);
  nand ginst7204 (U6548, R2358_U101, U2367);
  nand ginst7205 (U6549, R2337_U64, U2366);
  nand ginst7206 (U6550, REIP_REG_26__SCAN_IN, U6351);
  nand ginst7207 (U6551, R2099_U68, U2604);
  nand ginst7208 (U6552, R2096_U74, U7473);
  nand ginst7209 (U6553, EBX_REG_27__SCAN_IN, U7472);
  nand ginst7210 (U6554, PHYADDRPOINTER_REG_27__SCAN_IN, U2373);
  nand ginst7211 (U6555, R2358_U99, U2367);
  nand ginst7212 (U6556, R2337_U63, U2366);
  nand ginst7213 (U6557, REIP_REG_27__SCAN_IN, U6351);
  nand ginst7214 (U6558, R2099_U67, U2604);
  nand ginst7215 (U6559, R2096_U73, U7473);
  nand ginst7216 (U6560, EBX_REG_28__SCAN_IN, U7472);
  nand ginst7217 (U6561, PHYADDRPOINTER_REG_28__SCAN_IN, U2373);
  nand ginst7218 (U6562, R2358_U97, U2367);
  nand ginst7219 (U6563, R2337_U62, U2366);
  nand ginst7220 (U6564, REIP_REG_28__SCAN_IN, U6351);
  nand ginst7221 (U6565, R2099_U66, U2604);
  nand ginst7222 (U6566, R2096_U72, U7473);
  nand ginst7223 (U6567, EBX_REG_29__SCAN_IN, U7472);
  nand ginst7224 (U6568, PHYADDRPOINTER_REG_29__SCAN_IN, U2373);
  nand ginst7225 (U6569, R2358_U95, U2367);
  nand ginst7226 (U6570, R2337_U61, U2366);
  nand ginst7227 (U6571, REIP_REG_29__SCAN_IN, U6351);
  nand ginst7228 (U6572, R2099_U65, U2604);
  nand ginst7229 (U6573, R2096_U70, U7473);
  nand ginst7230 (U6574, EBX_REG_30__SCAN_IN, U7472);
  nand ginst7231 (U6575, PHYADDRPOINTER_REG_30__SCAN_IN, U2373);
  nand ginst7232 (U6576, R2358_U93, U2367);
  nand ginst7233 (U6577, R2337_U59, U2366);
  nand ginst7234 (U6578, REIP_REG_30__SCAN_IN, U6351);
  nand ginst7235 (U6579, R2099_U64, U2604);
  nand ginst7236 (U6580, R2096_U69, U7473);
  nand ginst7237 (U6581, EBX_REG_31__SCAN_IN, U7472);
  nand ginst7238 (U6582, PHYADDRPOINTER_REG_31__SCAN_IN, U2373);
  nand ginst7239 (U6583, R2358_U91, U2367);
  nand ginst7240 (U6584, R2337_U58, U2366);
  nand ginst7241 (U6585, REIP_REG_31__SCAN_IN, U6351);
  nand ginst7242 (U6586, DATAWIDTH_REG_0__SCAN_IN, DATAWIDTH_REG_1__SCAN_IN);
  or ginst7243 (U6587, REIP_REG_0__SCAN_IN, REIP_REG_1__SCAN_IN);
  not ginst7244 (U6588, U4165);
  nand ginst7245 (U6589, FLUSH_REG_SCAN_IN, U4165);
  nand ginst7246 (U6590, U2428, U3954);
  not ginst7247 (U6591, U4168);
  nand ginst7248 (U6592, STATEBS16_REG_SCAN_IN, U4485);
  nand ginst7249 (U6593, U4196, U6592);
  nand ginst7250 (U6594, U3952, U6593);
  nand ginst7251 (U6595, STATE2_REG_0__SCAN_IN, U6594);
  nand ginst7252 (U6596, U3259, U4181);
  nand ginst7253 (U6597, U3953, U6595);
  nand ginst7254 (U6598, U2368, U2473);
  nand ginst7255 (U6599, CODEFETCH_REG_SCAN_IN, U6598);
  nand ginst7256 (U6600, STATE2_REG_0__SCAN_IN, U4243);
  nand ginst7257 (U6601, ADS_N_REG_SCAN_IN, STATE_REG_0__SCAN_IN);
  not ginst7258 (U6602, U4169);
  nand ginst7259 (U6603, U3278, U3956);
  nand ginst7260 (U6604, U3393, U3957, U4487);
  nand ginst7261 (U6605, MEMORYFETCH_REG_SCAN_IN, U6604);
  nand ginst7262 (U6606, INSTQUEUE_REG_15__7__SCAN_IN, U2544);
  nand ginst7263 (U6607, INSTQUEUE_REG_14__7__SCAN_IN, U2543);
  nand ginst7264 (U6608, INSTQUEUE_REG_13__7__SCAN_IN, U2542);
  nand ginst7265 (U6609, INSTQUEUE_REG_12__7__SCAN_IN, U2541);
  nand ginst7266 (U6610, INSTQUEUE_REG_11__7__SCAN_IN, U2539);
  nand ginst7267 (U6611, INSTQUEUE_REG_10__7__SCAN_IN, U2538);
  nand ginst7268 (U6612, INSTQUEUE_REG_9__7__SCAN_IN, U2537);
  nand ginst7269 (U6613, INSTQUEUE_REG_8__7__SCAN_IN, U2536);
  nand ginst7270 (U6614, INSTQUEUE_REG_7__7__SCAN_IN, U2534);
  nand ginst7271 (U6615, INSTQUEUE_REG_6__7__SCAN_IN, U2533);
  nand ginst7272 (U6616, INSTQUEUE_REG_5__7__SCAN_IN, U2532);
  nand ginst7273 (U6617, INSTQUEUE_REG_4__7__SCAN_IN, U2531);
  nand ginst7274 (U6618, INSTQUEUE_REG_3__7__SCAN_IN, U2529);
  nand ginst7275 (U6619, INSTQUEUE_REG_2__7__SCAN_IN, U2527);
  nand ginst7276 (U6620, INSTQUEUE_REG_1__7__SCAN_IN, U2525);
  nand ginst7277 (U6621, INSTQUEUE_REG_0__7__SCAN_IN, U2523);
  nand ginst7278 (U6622, INSTQUEUE_REG_15__6__SCAN_IN, U2544);
  nand ginst7279 (U6623, INSTQUEUE_REG_14__6__SCAN_IN, U2543);
  nand ginst7280 (U6624, INSTQUEUE_REG_13__6__SCAN_IN, U2542);
  nand ginst7281 (U6625, INSTQUEUE_REG_12__6__SCAN_IN, U2541);
  nand ginst7282 (U6626, INSTQUEUE_REG_11__6__SCAN_IN, U2539);
  nand ginst7283 (U6627, INSTQUEUE_REG_10__6__SCAN_IN, U2538);
  nand ginst7284 (U6628, INSTQUEUE_REG_9__6__SCAN_IN, U2537);
  nand ginst7285 (U6629, INSTQUEUE_REG_8__6__SCAN_IN, U2536);
  nand ginst7286 (U6630, INSTQUEUE_REG_7__6__SCAN_IN, U2534);
  nand ginst7287 (U6631, INSTQUEUE_REG_6__6__SCAN_IN, U2533);
  nand ginst7288 (U6632, INSTQUEUE_REG_5__6__SCAN_IN, U2532);
  nand ginst7289 (U6633, INSTQUEUE_REG_4__6__SCAN_IN, U2531);
  nand ginst7290 (U6634, INSTQUEUE_REG_3__6__SCAN_IN, U2529);
  nand ginst7291 (U6635, INSTQUEUE_REG_2__6__SCAN_IN, U2527);
  nand ginst7292 (U6636, INSTQUEUE_REG_1__6__SCAN_IN, U2525);
  nand ginst7293 (U6637, INSTQUEUE_REG_0__6__SCAN_IN, U2523);
  nand ginst7294 (U6638, INSTQUEUE_REG_15__5__SCAN_IN, U2544);
  nand ginst7295 (U6639, INSTQUEUE_REG_14__5__SCAN_IN, U2543);
  nand ginst7296 (U6640, INSTQUEUE_REG_13__5__SCAN_IN, U2542);
  nand ginst7297 (U6641, INSTQUEUE_REG_12__5__SCAN_IN, U2541);
  nand ginst7298 (U6642, INSTQUEUE_REG_11__5__SCAN_IN, U2539);
  nand ginst7299 (U6643, INSTQUEUE_REG_10__5__SCAN_IN, U2538);
  nand ginst7300 (U6644, INSTQUEUE_REG_9__5__SCAN_IN, U2537);
  nand ginst7301 (U6645, INSTQUEUE_REG_8__5__SCAN_IN, U2536);
  nand ginst7302 (U6646, INSTQUEUE_REG_7__5__SCAN_IN, U2534);
  nand ginst7303 (U6647, INSTQUEUE_REG_6__5__SCAN_IN, U2533);
  nand ginst7304 (U6648, INSTQUEUE_REG_5__5__SCAN_IN, U2532);
  nand ginst7305 (U6649, INSTQUEUE_REG_4__5__SCAN_IN, U2531);
  nand ginst7306 (U6650, INSTQUEUE_REG_3__5__SCAN_IN, U2529);
  nand ginst7307 (U6651, INSTQUEUE_REG_2__5__SCAN_IN, U2527);
  nand ginst7308 (U6652, INSTQUEUE_REG_1__5__SCAN_IN, U2525);
  nand ginst7309 (U6653, INSTQUEUE_REG_0__5__SCAN_IN, U2523);
  nand ginst7310 (U6654, INSTQUEUE_REG_15__4__SCAN_IN, U2544);
  nand ginst7311 (U6655, INSTQUEUE_REG_14__4__SCAN_IN, U2543);
  nand ginst7312 (U6656, INSTQUEUE_REG_13__4__SCAN_IN, U2542);
  nand ginst7313 (U6657, INSTQUEUE_REG_12__4__SCAN_IN, U2541);
  nand ginst7314 (U6658, INSTQUEUE_REG_11__4__SCAN_IN, U2539);
  nand ginst7315 (U6659, INSTQUEUE_REG_10__4__SCAN_IN, U2538);
  nand ginst7316 (U6660, INSTQUEUE_REG_9__4__SCAN_IN, U2537);
  nand ginst7317 (U6661, INSTQUEUE_REG_8__4__SCAN_IN, U2536);
  nand ginst7318 (U6662, INSTQUEUE_REG_7__4__SCAN_IN, U2534);
  nand ginst7319 (U6663, INSTQUEUE_REG_6__4__SCAN_IN, U2533);
  nand ginst7320 (U6664, INSTQUEUE_REG_5__4__SCAN_IN, U2532);
  nand ginst7321 (U6665, INSTQUEUE_REG_4__4__SCAN_IN, U2531);
  nand ginst7322 (U6666, INSTQUEUE_REG_3__4__SCAN_IN, U2529);
  nand ginst7323 (U6667, INSTQUEUE_REG_2__4__SCAN_IN, U2527);
  nand ginst7324 (U6668, INSTQUEUE_REG_1__4__SCAN_IN, U2525);
  nand ginst7325 (U6669, INSTQUEUE_REG_15__3__SCAN_IN, U2544);
  nand ginst7326 (U6670, INSTQUEUE_REG_14__3__SCAN_IN, U2543);
  nand ginst7327 (U6671, INSTQUEUE_REG_13__3__SCAN_IN, U2542);
  nand ginst7328 (U6672, INSTQUEUE_REG_12__3__SCAN_IN, U2541);
  nand ginst7329 (U6673, INSTQUEUE_REG_11__3__SCAN_IN, U2539);
  nand ginst7330 (U6674, INSTQUEUE_REG_10__3__SCAN_IN, U2538);
  nand ginst7331 (U6675, INSTQUEUE_REG_9__3__SCAN_IN, U2537);
  nand ginst7332 (U6676, INSTQUEUE_REG_8__3__SCAN_IN, U2536);
  nand ginst7333 (U6677, INSTQUEUE_REG_7__3__SCAN_IN, U2534);
  nand ginst7334 (U6678, INSTQUEUE_REG_6__3__SCAN_IN, U2533);
  nand ginst7335 (U6679, INSTQUEUE_REG_5__3__SCAN_IN, U2532);
  nand ginst7336 (U6680, INSTQUEUE_REG_4__3__SCAN_IN, U2531);
  nand ginst7337 (U6681, INSTQUEUE_REG_3__3__SCAN_IN, U2529);
  nand ginst7338 (U6682, INSTQUEUE_REG_2__3__SCAN_IN, U2527);
  nand ginst7339 (U6683, INSTQUEUE_REG_1__3__SCAN_IN, U2525);
  nand ginst7340 (U6684, INSTQUEUE_REG_0__3__SCAN_IN, U2523);
  nand ginst7341 (U6685, INSTQUEUE_REG_15__2__SCAN_IN, U2544);
  nand ginst7342 (U6686, INSTQUEUE_REG_14__2__SCAN_IN, U2543);
  nand ginst7343 (U6687, INSTQUEUE_REG_13__2__SCAN_IN, U2542);
  nand ginst7344 (U6688, INSTQUEUE_REG_12__2__SCAN_IN, U2541);
  nand ginst7345 (U6689, INSTQUEUE_REG_11__2__SCAN_IN, U2539);
  nand ginst7346 (U6690, INSTQUEUE_REG_10__2__SCAN_IN, U2538);
  nand ginst7347 (U6691, INSTQUEUE_REG_9__2__SCAN_IN, U2537);
  nand ginst7348 (U6692, INSTQUEUE_REG_8__2__SCAN_IN, U2536);
  nand ginst7349 (U6693, INSTQUEUE_REG_7__2__SCAN_IN, U2534);
  nand ginst7350 (U6694, INSTQUEUE_REG_6__2__SCAN_IN, U2533);
  nand ginst7351 (U6695, INSTQUEUE_REG_5__2__SCAN_IN, U2532);
  nand ginst7352 (U6696, INSTQUEUE_REG_4__2__SCAN_IN, U2531);
  nand ginst7353 (U6697, INSTQUEUE_REG_3__2__SCAN_IN, U2529);
  nand ginst7354 (U6698, INSTQUEUE_REG_2__2__SCAN_IN, U2527);
  nand ginst7355 (U6699, INSTQUEUE_REG_1__2__SCAN_IN, U2525);
  nand ginst7356 (U6700, INSTQUEUE_REG_0__2__SCAN_IN, U2523);
  nand ginst7357 (U6701, INSTQUEUE_REG_15__1__SCAN_IN, U2544);
  nand ginst7358 (U6702, INSTQUEUE_REG_14__1__SCAN_IN, U2543);
  nand ginst7359 (U6703, INSTQUEUE_REG_13__1__SCAN_IN, U2542);
  nand ginst7360 (U6704, INSTQUEUE_REG_12__1__SCAN_IN, U2541);
  nand ginst7361 (U6705, INSTQUEUE_REG_11__1__SCAN_IN, U2539);
  nand ginst7362 (U6706, INSTQUEUE_REG_10__1__SCAN_IN, U2538);
  nand ginst7363 (U6707, INSTQUEUE_REG_9__1__SCAN_IN, U2537);
  nand ginst7364 (U6708, INSTQUEUE_REG_8__1__SCAN_IN, U2536);
  nand ginst7365 (U6709, INSTQUEUE_REG_7__1__SCAN_IN, U2534);
  nand ginst7366 (U6710, INSTQUEUE_REG_6__1__SCAN_IN, U2533);
  nand ginst7367 (U6711, INSTQUEUE_REG_5__1__SCAN_IN, U2532);
  nand ginst7368 (U6712, INSTQUEUE_REG_4__1__SCAN_IN, U2531);
  nand ginst7369 (U6713, INSTQUEUE_REG_3__1__SCAN_IN, U2529);
  nand ginst7370 (U6714, INSTQUEUE_REG_2__1__SCAN_IN, U2527);
  nand ginst7371 (U6715, INSTQUEUE_REG_1__1__SCAN_IN, U2525);
  nand ginst7372 (U6716, INSTQUEUE_REG_0__1__SCAN_IN, U2523);
  nand ginst7373 (U6717, INSTQUEUE_REG_15__0__SCAN_IN, U2544);
  nand ginst7374 (U6718, INSTQUEUE_REG_14__0__SCAN_IN, U2543);
  nand ginst7375 (U6719, INSTQUEUE_REG_13__0__SCAN_IN, U2542);
  nand ginst7376 (U6720, INSTQUEUE_REG_12__0__SCAN_IN, U2541);
  nand ginst7377 (U6721, INSTQUEUE_REG_11__0__SCAN_IN, U2539);
  nand ginst7378 (U6722, INSTQUEUE_REG_10__0__SCAN_IN, U2538);
  nand ginst7379 (U6723, INSTQUEUE_REG_9__0__SCAN_IN, U2537);
  nand ginst7380 (U6724, INSTQUEUE_REG_8__0__SCAN_IN, U2536);
  nand ginst7381 (U6725, INSTQUEUE_REG_7__0__SCAN_IN, U2534);
  nand ginst7382 (U6726, INSTQUEUE_REG_6__0__SCAN_IN, U2533);
  nand ginst7383 (U6727, INSTQUEUE_REG_5__0__SCAN_IN, U2532);
  nand ginst7384 (U6728, INSTQUEUE_REG_4__0__SCAN_IN, U2531);
  nand ginst7385 (U6729, INSTQUEUE_REG_3__0__SCAN_IN, U2529);
  nand ginst7386 (U6730, INSTQUEUE_REG_2__0__SCAN_IN, U2527);
  nand ginst7387 (U6731, INSTQUEUE_REG_1__0__SCAN_IN, U2525);
  nand ginst7388 (U6732, INSTQUEUE_REG_0__0__SCAN_IN, U2523);
  nand ginst7389 (U6733, STATE2_REG_2__SCAN_IN, U4448);
  nand ginst7390 (U6734, U3399, U6733);
  nand ginst7391 (U6735, EAX_REG_9__SCAN_IN, U4176);
  nand ginst7392 (U6736, PHYADDRPOINTER_REG_9__SCAN_IN, U4175);
  nand ginst7393 (U6737, R2337_U51, U2352);
  nand ginst7394 (U6738, EAX_REG_8__SCAN_IN, U4176);
  nand ginst7395 (U6739, PHYADDRPOINTER_REG_8__SCAN_IN, U4175);
  nand ginst7396 (U6740, R2337_U52, U2352);
  nand ginst7397 (U6741, EAX_REG_7__SCAN_IN, U4176);
  nand ginst7398 (U6742, PHYADDRPOINTER_REG_7__SCAN_IN, U4175);
  nand ginst7399 (U6743, R2337_U53, U2352);
  nand ginst7400 (U6744, EAX_REG_6__SCAN_IN, U4176);
  nand ginst7401 (U6745, PHYADDRPOINTER_REG_6__SCAN_IN, U4175);
  nand ginst7402 (U6746, R2337_U54, U2352);
  nand ginst7403 (U6747, R2182_U5, U6734);
  nand ginst7404 (U6748, EAX_REG_5__SCAN_IN, U4176);
  nand ginst7405 (U6749, PHYADDRPOINTER_REG_5__SCAN_IN, U4175);
  nand ginst7406 (U6750, R2337_U55, U2352);
  nand ginst7407 (U6751, R2182_U24, U6734);
  nand ginst7408 (U6752, EAX_REG_4__SCAN_IN, U4176);
  nand ginst7409 (U6753, PHYADDRPOINTER_REG_4__SCAN_IN, U4175);
  nand ginst7410 (U6754, R2337_U56, U2352);
  nand ginst7411 (U6755, INSTQUEUERD_ADDR_REG_4__SCAN_IN, U2353);
  nand ginst7412 (U6756, EAX_REG_31__SCAN_IN, U4176);
  nand ginst7413 (U6757, PHYADDRPOINTER_REG_31__SCAN_IN, U4175);
  nand ginst7414 (U6758, R2337_U58, U2352);
  nand ginst7415 (U6759, R2182_U26, U6734);
  nand ginst7416 (U6760, EAX_REG_30__SCAN_IN, U4176);
  nand ginst7417 (U6761, PHYADDRPOINTER_REG_30__SCAN_IN, U4175);
  nand ginst7418 (U6762, R2337_U59, U2352);
  nand ginst7419 (U6763, R2182_U25, U6734);
  nand ginst7420 (U6764, EAX_REG_3__SCAN_IN, U4176);
  nand ginst7421 (U6765, PHYADDRPOINTER_REG_3__SCAN_IN, U4175);
  nand ginst7422 (U6766, R2337_U57, U2352);
  nand ginst7423 (U6767, INSTQUEUERD_ADDR_REG_3__SCAN_IN, U2353);
  nand ginst7424 (U6768, R2182_U27, U6734);
  nand ginst7425 (U6769, EAX_REG_29__SCAN_IN, U4176);
  nand ginst7426 (U6770, PHYADDRPOINTER_REG_29__SCAN_IN, U4175);
  nand ginst7427 (U6771, R2337_U61, U2352);
  nand ginst7428 (U6772, R2182_U28, U6734);
  nand ginst7429 (U6773, EAX_REG_28__SCAN_IN, U4176);
  nand ginst7430 (U6774, PHYADDRPOINTER_REG_28__SCAN_IN, U4175);
  nand ginst7431 (U6775, R2337_U62, U2352);
  nand ginst7432 (U6776, R2182_U29, U6734);
  nand ginst7433 (U6777, EAX_REG_27__SCAN_IN, U4176);
  nand ginst7434 (U6778, PHYADDRPOINTER_REG_27__SCAN_IN, U4175);
  nand ginst7435 (U6779, R2337_U63, U2352);
  nand ginst7436 (U6780, R2182_U30, U6734);
  nand ginst7437 (U6781, EAX_REG_26__SCAN_IN, U4176);
  nand ginst7438 (U6782, PHYADDRPOINTER_REG_26__SCAN_IN, U4175);
  nand ginst7439 (U6783, R2337_U64, U2352);
  nand ginst7440 (U6784, R2182_U31, U6734);
  nand ginst7441 (U6785, EAX_REG_25__SCAN_IN, U4176);
  nand ginst7442 (U6786, PHYADDRPOINTER_REG_25__SCAN_IN, U4175);
  nand ginst7443 (U6787, R2337_U65, U2352);
  nand ginst7444 (U6788, R2182_U32, U6734);
  nand ginst7445 (U6789, EAX_REG_24__SCAN_IN, U4176);
  nand ginst7446 (U6790, PHYADDRPOINTER_REG_24__SCAN_IN, U4175);
  nand ginst7447 (U6791, R2337_U66, U2352);
  nand ginst7448 (U6792, R2182_U6, U6734);
  nand ginst7449 (U6793, EAX_REG_23__SCAN_IN, U4176);
  nand ginst7450 (U6794, PHYADDRPOINTER_REG_23__SCAN_IN, U4175);
  nand ginst7451 (U6795, R2337_U67, U2352);
  nand ginst7452 (U6796, U2724, U6734);
  nand ginst7453 (U6797, EAX_REG_22__SCAN_IN, U4176);
  nand ginst7454 (U6798, PHYADDRPOINTER_REG_22__SCAN_IN, U4175);
  nand ginst7455 (U6799, R2337_U68, U2352);
  nand ginst7456 (U6800, U2725, U6734);
  nand ginst7457 (U6801, EAX_REG_21__SCAN_IN, U4176);
  nand ginst7458 (U6802, PHYADDRPOINTER_REG_21__SCAN_IN, U4175);
  nand ginst7459 (U6803, R2337_U69, U2352);
  nand ginst7460 (U6804, U2726, U6734);
  nand ginst7461 (U6805, EAX_REG_20__SCAN_IN, U4176);
  nand ginst7462 (U6806, PHYADDRPOINTER_REG_20__SCAN_IN, U4175);
  nand ginst7463 (U6807, R2337_U70, U2352);
  nand ginst7464 (U6808, R2182_U42, U6734);
  nand ginst7465 (U6809, EAX_REG_2__SCAN_IN, U4176);
  nand ginst7466 (U6810, PHYADDRPOINTER_REG_2__SCAN_IN, U4175);
  nand ginst7467 (U6811, R2337_U60, U2352);
  nand ginst7468 (U6812, INSTQUEUERD_ADDR_REG_2__SCAN_IN, U2353);
  nand ginst7469 (U6813, U2727, U6734);
  nand ginst7470 (U6814, EAX_REG_19__SCAN_IN, U4176);
  nand ginst7471 (U6815, PHYADDRPOINTER_REG_19__SCAN_IN, U4175);
  nand ginst7472 (U6816, R2337_U71, U2352);
  nand ginst7473 (U6817, U2728, U6734);
  nand ginst7474 (U6818, EAX_REG_18__SCAN_IN, U4176);
  nand ginst7475 (U6819, PHYADDRPOINTER_REG_18__SCAN_IN, U4175);
  nand ginst7476 (U6820, R2337_U72, U2352);
  nand ginst7477 (U6821, U2729, U6734);
  nand ginst7478 (U6822, EAX_REG_17__SCAN_IN, U4176);
  nand ginst7479 (U6823, PHYADDRPOINTER_REG_17__SCAN_IN, U4175);
  nand ginst7480 (U6824, R2337_U73, U2352);
  nand ginst7481 (U6825, U2730, U6734);
  nand ginst7482 (U6826, EAX_REG_16__SCAN_IN, U4176);
  nand ginst7483 (U6827, PHYADDRPOINTER_REG_16__SCAN_IN, U4175);
  nand ginst7484 (U6828, R2337_U74, U2352);
  nand ginst7485 (U6829, EAX_REG_15__SCAN_IN, U4176);
  nand ginst7486 (U6830, PHYADDRPOINTER_REG_15__SCAN_IN, U4175);
  nand ginst7487 (U6831, R2337_U75, U2352);
  nand ginst7488 (U6832, EAX_REG_14__SCAN_IN, U4176);
  nand ginst7489 (U6833, PHYADDRPOINTER_REG_14__SCAN_IN, U4175);
  nand ginst7490 (U6834, R2337_U76, U2352);
  nand ginst7491 (U6835, EAX_REG_13__SCAN_IN, U4176);
  nand ginst7492 (U6836, PHYADDRPOINTER_REG_13__SCAN_IN, U4175);
  nand ginst7493 (U6837, R2337_U77, U2352);
  nand ginst7494 (U6838, EAX_REG_12__SCAN_IN, U4176);
  nand ginst7495 (U6839, PHYADDRPOINTER_REG_12__SCAN_IN, U4175);
  nand ginst7496 (U6840, R2337_U78, U2352);
  nand ginst7497 (U6841, EAX_REG_11__SCAN_IN, U4176);
  nand ginst7498 (U6842, PHYADDRPOINTER_REG_11__SCAN_IN, U4175);
  nand ginst7499 (U6843, R2337_U79, U2352);
  nand ginst7500 (U6844, EAX_REG_10__SCAN_IN, U4176);
  nand ginst7501 (U6845, PHYADDRPOINTER_REG_10__SCAN_IN, U4175);
  nand ginst7502 (U6846, R2337_U80, U2352);
  nand ginst7503 (U6847, R2182_U33, U6734);
  nand ginst7504 (U6848, EAX_REG_1__SCAN_IN, U4176);
  nand ginst7505 (U6849, PHYADDRPOINTER_REG_1__SCAN_IN, U4175);
  nand ginst7506 (U6850, R2337_U5, U2352);
  nand ginst7507 (U6851, INSTQUEUERD_ADDR_REG_1__SCAN_IN, U2353);
  nand ginst7508 (U6852, R2182_U34, U6734);
  nand ginst7509 (U6853, EAX_REG_0__SCAN_IN, U4176);
  nand ginst7510 (U6854, PHYADDRPOINTER_REG_0__SCAN_IN, U4175);
  nand ginst7511 (U6855, PHYADDRPOINTER_REG_0__SCAN_IN, U2352);
  nand ginst7512 (U6856, INSTQUEUERD_ADDR_REG_0__SCAN_IN, U2353);
  nand ginst7513 (U6857, R2144_U49, U6734);
  nand ginst7514 (U6858, U3296, U3426, U4448);
  nand ginst7515 (U6859, R2144_U80, U4147);
  nand ginst7516 (U6860, ADD_371_U6, U4196);
  nand ginst7517 (U6861, R2144_U10, U4147);
  nand ginst7518 (U6862, ADD_371_U17, U4196);
  nand ginst7519 (U6863, R2144_U9, U4147);
  nand ginst7520 (U6864, ADD_371_U18, U4196);
  nand ginst7521 (U6865, R2144_U45, U4147);
  nand ginst7522 (U6866, ADD_371_U19, U4196);
  nand ginst7523 (U6867, R2144_U47, U4147);
  nand ginst7524 (U6868, ADD_371_U20, U4196);
  nand ginst7525 (U6869, R2144_U8, U4147);
  nand ginst7526 (U6870, ADD_371_U25, U4196);
  nand ginst7527 (U6871, R2144_U49, U4147);
  nand ginst7528 (U6872, ADD_371_U5, U4196);
  nand ginst7529 (U6873, U3270, U4482);
  nand ginst7530 (U6874, R2144_U50, U4147);
  nand ginst7531 (U6875, ADD_371_U21, U4196);
  nand ginst7532 (U6876, U2605, U3271);
  nand ginst7533 (U6877, R2144_U43, U4147);
  nand ginst7534 (U6878, ADD_371_U4, U4196);
  nand ginst7535 (U6879, U3270, U4482);
  nand ginst7536 (U6880, INSTQUEUE_REG_15__1__SCAN_IN, U2564);
  nand ginst7537 (U6881, INSTQUEUE_REG_14__1__SCAN_IN, U2563);
  nand ginst7538 (U6882, INSTQUEUE_REG_13__1__SCAN_IN, U2562);
  nand ginst7539 (U6883, INSTQUEUE_REG_12__1__SCAN_IN, U2561);
  nand ginst7540 (U6884, INSTQUEUE_REG_11__1__SCAN_IN, U2559);
  nand ginst7541 (U6885, INSTQUEUE_REG_10__1__SCAN_IN, U2558);
  nand ginst7542 (U6886, INSTQUEUE_REG_9__1__SCAN_IN, U2557);
  nand ginst7543 (U6887, INSTQUEUE_REG_8__1__SCAN_IN, U2556);
  nand ginst7544 (U6888, INSTQUEUE_REG_7__1__SCAN_IN, U2554);
  nand ginst7545 (U6889, INSTQUEUE_REG_6__1__SCAN_IN, U2553);
  nand ginst7546 (U6890, INSTQUEUE_REG_5__1__SCAN_IN, U2552);
  nand ginst7547 (U6891, INSTQUEUE_REG_4__1__SCAN_IN, U2551);
  nand ginst7548 (U6892, INSTQUEUE_REG_3__1__SCAN_IN, U2549);
  nand ginst7549 (U6893, INSTQUEUE_REG_2__1__SCAN_IN, U2548);
  nand ginst7550 (U6894, INSTQUEUE_REG_1__1__SCAN_IN, U2547);
  nand ginst7551 (U6895, INSTQUEUE_REG_0__1__SCAN_IN, U2546);
  nand ginst7552 (U6896, U4017, U4018, U4019, U4020);
  nand ginst7553 (U6897, U3392, U3405);
  nand ginst7554 (U6898, INSTQUEUE_REG_15__0__SCAN_IN, U2564);
  nand ginst7555 (U6899, INSTQUEUE_REG_14__0__SCAN_IN, U2563);
  nand ginst7556 (U6900, INSTQUEUE_REG_13__0__SCAN_IN, U2562);
  nand ginst7557 (U6901, INSTQUEUE_REG_12__0__SCAN_IN, U2561);
  nand ginst7558 (U6902, INSTQUEUE_REG_11__0__SCAN_IN, U2559);
  nand ginst7559 (U6903, INSTQUEUE_REG_10__0__SCAN_IN, U2558);
  nand ginst7560 (U6904, INSTQUEUE_REG_9__0__SCAN_IN, U2557);
  nand ginst7561 (U6905, INSTQUEUE_REG_8__0__SCAN_IN, U2556);
  nand ginst7562 (U6906, INSTQUEUE_REG_7__0__SCAN_IN, U2554);
  nand ginst7563 (U6907, INSTQUEUE_REG_6__0__SCAN_IN, U2553);
  nand ginst7564 (U6908, INSTQUEUE_REG_5__0__SCAN_IN, U2552);
  nand ginst7565 (U6909, INSTQUEUE_REG_4__0__SCAN_IN, U2551);
  nand ginst7566 (U6910, INSTQUEUE_REG_3__0__SCAN_IN, U2549);
  nand ginst7567 (U6911, INSTQUEUE_REG_2__0__SCAN_IN, U2548);
  nand ginst7568 (U6912, INSTQUEUE_REG_1__0__SCAN_IN, U2547);
  nand ginst7569 (U6913, INSTQUEUE_REG_0__0__SCAN_IN, U2546);
  nand ginst7570 (U6914, U4021, U4022, U4023, U4024);
  nand ginst7571 (U6915, U3221, U4195);
  nand ginst7572 (U6916, SUB_357_U8, U2355);
  nand ginst7573 (U6917, U3220, U4195);
  nand ginst7574 (U6918, SUB_357_U6, U2355);
  nand ginst7575 (U6919, U3219, U4195);
  nand ginst7576 (U6920, SUB_357_U9, U2355);
  nand ginst7577 (U6921, U3218, U4195);
  nand ginst7578 (U6922, SUB_357_U13, U2355);
  nand ginst7579 (U6923, U3217, U4195);
  nand ginst7580 (U6924, SUB_357_U11, U2355);
  nand ginst7581 (U6925, R2182_U25, U3281);
  nand ginst7582 (U6926, U3216, U4195);
  nand ginst7583 (U6927, SUB_357_U12, U2355);
  nand ginst7584 (U6928, R2182_U42, U3281);
  nand ginst7585 (U6929, INSTQUEUE_REG_15__7__SCAN_IN, U2564);
  nand ginst7586 (U6930, INSTQUEUE_REG_14__7__SCAN_IN, U2563);
  nand ginst7587 (U6931, INSTQUEUE_REG_13__7__SCAN_IN, U2562);
  nand ginst7588 (U6932, INSTQUEUE_REG_12__7__SCAN_IN, U2561);
  nand ginst7589 (U6933, INSTQUEUE_REG_11__7__SCAN_IN, U2559);
  nand ginst7590 (U6934, INSTQUEUE_REG_10__7__SCAN_IN, U2558);
  nand ginst7591 (U6935, INSTQUEUE_REG_9__7__SCAN_IN, U2557);
  nand ginst7592 (U6936, INSTQUEUE_REG_8__7__SCAN_IN, U2556);
  nand ginst7593 (U6937, INSTQUEUE_REG_7__7__SCAN_IN, U2554);
  nand ginst7594 (U6938, INSTQUEUE_REG_6__7__SCAN_IN, U2553);
  nand ginst7595 (U6939, INSTQUEUE_REG_5__7__SCAN_IN, U2552);
  nand ginst7596 (U6940, INSTQUEUE_REG_4__7__SCAN_IN, U2551);
  nand ginst7597 (U6941, INSTQUEUE_REG_3__7__SCAN_IN, U2549);
  nand ginst7598 (U6942, INSTQUEUE_REG_2__7__SCAN_IN, U2548);
  nand ginst7599 (U6943, INSTQUEUE_REG_1__7__SCAN_IN, U2547);
  nand ginst7600 (U6944, INSTQUEUE_REG_0__7__SCAN_IN, U2546);
  nand ginst7601 (U6945, U4025, U4026, U4027, U4028);
  nand ginst7602 (U6946, INSTQUEUE_REG_15__6__SCAN_IN, U2564);
  nand ginst7603 (U6947, INSTQUEUE_REG_14__6__SCAN_IN, U2563);
  nand ginst7604 (U6948, INSTQUEUE_REG_13__6__SCAN_IN, U2562);
  nand ginst7605 (U6949, INSTQUEUE_REG_12__6__SCAN_IN, U2561);
  nand ginst7606 (U6950, INSTQUEUE_REG_11__6__SCAN_IN, U2559);
  nand ginst7607 (U6951, INSTQUEUE_REG_10__6__SCAN_IN, U2558);
  nand ginst7608 (U6952, INSTQUEUE_REG_9__6__SCAN_IN, U2557);
  nand ginst7609 (U6953, INSTQUEUE_REG_8__6__SCAN_IN, U2556);
  nand ginst7610 (U6954, INSTQUEUE_REG_7__6__SCAN_IN, U2554);
  nand ginst7611 (U6955, INSTQUEUE_REG_6__6__SCAN_IN, U2553);
  nand ginst7612 (U6956, INSTQUEUE_REG_5__6__SCAN_IN, U2552);
  nand ginst7613 (U6957, INSTQUEUE_REG_4__6__SCAN_IN, U2551);
  nand ginst7614 (U6958, INSTQUEUE_REG_3__6__SCAN_IN, U2549);
  nand ginst7615 (U6959, INSTQUEUE_REG_2__6__SCAN_IN, U2548);
  nand ginst7616 (U6960, INSTQUEUE_REG_1__6__SCAN_IN, U2547);
  nand ginst7617 (U6961, INSTQUEUE_REG_0__6__SCAN_IN, U2546);
  nand ginst7618 (U6962, U4029, U4030, U4031, U4032);
  nand ginst7619 (U6963, INSTQUEUE_REG_15__5__SCAN_IN, U2564);
  nand ginst7620 (U6964, INSTQUEUE_REG_14__5__SCAN_IN, U2563);
  nand ginst7621 (U6965, INSTQUEUE_REG_13__5__SCAN_IN, U2562);
  nand ginst7622 (U6966, INSTQUEUE_REG_12__5__SCAN_IN, U2561);
  nand ginst7623 (U6967, INSTQUEUE_REG_11__5__SCAN_IN, U2559);
  nand ginst7624 (U6968, INSTQUEUE_REG_10__5__SCAN_IN, U2558);
  nand ginst7625 (U6969, INSTQUEUE_REG_9__5__SCAN_IN, U2557);
  nand ginst7626 (U6970, INSTQUEUE_REG_8__5__SCAN_IN, U2556);
  nand ginst7627 (U6971, INSTQUEUE_REG_7__5__SCAN_IN, U2554);
  nand ginst7628 (U6972, INSTQUEUE_REG_6__5__SCAN_IN, U2553);
  nand ginst7629 (U6973, INSTQUEUE_REG_5__5__SCAN_IN, U2552);
  nand ginst7630 (U6974, INSTQUEUE_REG_4__5__SCAN_IN, U2551);
  nand ginst7631 (U6975, INSTQUEUE_REG_3__5__SCAN_IN, U2549);
  nand ginst7632 (U6976, INSTQUEUE_REG_2__5__SCAN_IN, U2548);
  nand ginst7633 (U6977, INSTQUEUE_REG_1__5__SCAN_IN, U2547);
  nand ginst7634 (U6978, INSTQUEUE_REG_0__5__SCAN_IN, U2546);
  nand ginst7635 (U6979, U4033, U4034, U4035, U4036);
  nand ginst7636 (U6980, INSTQUEUE_REG_15__4__SCAN_IN, U2564);
  nand ginst7637 (U6981, INSTQUEUE_REG_14__4__SCAN_IN, U2563);
  nand ginst7638 (U6982, INSTQUEUE_REG_13__4__SCAN_IN, U2562);
  nand ginst7639 (U6983, INSTQUEUE_REG_12__4__SCAN_IN, U2561);
  nand ginst7640 (U6984, INSTQUEUE_REG_11__4__SCAN_IN, U2559);
  nand ginst7641 (U6985, INSTQUEUE_REG_10__4__SCAN_IN, U2558);
  nand ginst7642 (U6986, INSTQUEUE_REG_9__4__SCAN_IN, U2557);
  nand ginst7643 (U6987, INSTQUEUE_REG_8__4__SCAN_IN, U2556);
  nand ginst7644 (U6988, INSTQUEUE_REG_7__4__SCAN_IN, U2554);
  nand ginst7645 (U6989, INSTQUEUE_REG_6__4__SCAN_IN, U2553);
  nand ginst7646 (U6990, INSTQUEUE_REG_5__4__SCAN_IN, U2552);
  nand ginst7647 (U6991, INSTQUEUE_REG_4__4__SCAN_IN, U2551);
  nand ginst7648 (U6992, INSTQUEUE_REG_3__4__SCAN_IN, U2549);
  nand ginst7649 (U6993, INSTQUEUE_REG_2__4__SCAN_IN, U2548);
  nand ginst7650 (U6994, INSTQUEUE_REG_1__4__SCAN_IN, U2547);
  nand ginst7651 (U6995, INSTQUEUE_REG_15__3__SCAN_IN, U2564);
  nand ginst7652 (U6996, INSTQUEUE_REG_14__3__SCAN_IN, U2563);
  nand ginst7653 (U6997, INSTQUEUE_REG_13__3__SCAN_IN, U2562);
  nand ginst7654 (U6998, INSTQUEUE_REG_12__3__SCAN_IN, U2561);
  nand ginst7655 (U6999, INSTQUEUE_REG_11__3__SCAN_IN, U2559);
  nand ginst7656 (U7000, INSTQUEUE_REG_10__3__SCAN_IN, U2558);
  nand ginst7657 (U7001, INSTQUEUE_REG_9__3__SCAN_IN, U2557);
  nand ginst7658 (U7002, INSTQUEUE_REG_8__3__SCAN_IN, U2556);
  nand ginst7659 (U7003, INSTQUEUE_REG_7__3__SCAN_IN, U2554);
  nand ginst7660 (U7004, INSTQUEUE_REG_6__3__SCAN_IN, U2553);
  nand ginst7661 (U7005, INSTQUEUE_REG_5__3__SCAN_IN, U2552);
  nand ginst7662 (U7006, INSTQUEUE_REG_4__3__SCAN_IN, U2551);
  nand ginst7663 (U7007, INSTQUEUE_REG_3__3__SCAN_IN, U2549);
  nand ginst7664 (U7008, INSTQUEUE_REG_2__3__SCAN_IN, U2548);
  nand ginst7665 (U7009, INSTQUEUE_REG_1__3__SCAN_IN, U2547);
  nand ginst7666 (U7010, INSTQUEUE_REG_0__3__SCAN_IN, U2546);
  nand ginst7667 (U7011, U4041, U4042, U4043, U4044);
  nand ginst7668 (U7012, INSTQUEUE_REG_15__2__SCAN_IN, U2564);
  nand ginst7669 (U7013, INSTQUEUE_REG_14__2__SCAN_IN, U2563);
  nand ginst7670 (U7014, INSTQUEUE_REG_13__2__SCAN_IN, U2562);
  nand ginst7671 (U7015, INSTQUEUE_REG_12__2__SCAN_IN, U2561);
  nand ginst7672 (U7016, INSTQUEUE_REG_11__2__SCAN_IN, U2559);
  nand ginst7673 (U7017, INSTQUEUE_REG_10__2__SCAN_IN, U2558);
  nand ginst7674 (U7018, INSTQUEUE_REG_9__2__SCAN_IN, U2557);
  nand ginst7675 (U7019, INSTQUEUE_REG_8__2__SCAN_IN, U2556);
  nand ginst7676 (U7020, INSTQUEUE_REG_7__2__SCAN_IN, U2554);
  nand ginst7677 (U7021, INSTQUEUE_REG_6__2__SCAN_IN, U2553);
  nand ginst7678 (U7022, INSTQUEUE_REG_5__2__SCAN_IN, U2552);
  nand ginst7679 (U7023, INSTQUEUE_REG_4__2__SCAN_IN, U2551);
  nand ginst7680 (U7024, INSTQUEUE_REG_3__2__SCAN_IN, U2549);
  nand ginst7681 (U7025, INSTQUEUE_REG_2__2__SCAN_IN, U2548);
  nand ginst7682 (U7026, INSTQUEUE_REG_1__2__SCAN_IN, U2547);
  nand ginst7683 (U7027, INSTQUEUE_REG_0__2__SCAN_IN, U2546);
  nand ginst7684 (U7028, U4045, U4046, U4047, U4048);
  nand ginst7685 (U7029, U3215, U4195);
  nand ginst7686 (U7030, SUB_357_U7, U2355);
  nand ginst7687 (U7031, R2182_U33, U3281);
  nand ginst7688 (U7032, U3214, U4195);
  nand ginst7689 (U7033, SUB_357_U10, U2355);
  nand ginst7690 (U7034, R2182_U34, U3281);
  nand ginst7691 (U7035, U3221, U4194);
  nand ginst7692 (U7036, INSTQUEUE_REG_0__7__SCAN_IN, U4180);
  nand ginst7693 (U7037, U3220, U4194);
  nand ginst7694 (U7038, INSTQUEUE_REG_0__6__SCAN_IN, U4180);
  nand ginst7695 (U7039, U3219, U4194);
  nand ginst7696 (U7040, INSTQUEUE_REG_0__5__SCAN_IN, U4180);
  nand ginst7697 (U7041, U3218, U4194);
  nand ginst7698 (U7042, U3217, U4194);
  nand ginst7699 (U7043, INSTQUEUE_REG_0__3__SCAN_IN, U4180);
  nand ginst7700 (U7044, U3216, U4194);
  nand ginst7701 (U7045, INSTQUEUE_REG_0__2__SCAN_IN, U4180);
  nand ginst7702 (U7046, U3215, U4194);
  nand ginst7703 (U7047, INSTQUEUE_REG_0__1__SCAN_IN, U4180);
  nand ginst7704 (U7048, U3214, U4194);
  nand ginst7705 (U7049, U3221, U4388);
  nand ginst7706 (U7050, INSTQUEUE_REG_0__0__SCAN_IN, U4180);
  nand ginst7707 (U7051, U3414, U3415);
  nand ginst7708 (U7052, INSTQUEUERD_ADDR_REG_3__SCAN_IN, U3251);
  not ginst7709 (U7053, U3432);
  nand ginst7710 (U7054, INSTQUEUE_REG_8__7__SCAN_IN, U2582);
  nand ginst7711 (U7055, INSTQUEUE_REG_9__7__SCAN_IN, U2581);
  nand ginst7712 (U7056, INSTQUEUE_REG_10__7__SCAN_IN, U2580);
  nand ginst7713 (U7057, INSTQUEUE_REG_11__7__SCAN_IN, U2579);
  nand ginst7714 (U7058, INSTQUEUE_REG_12__7__SCAN_IN, U2577);
  nand ginst7715 (U7059, INSTQUEUE_REG_13__7__SCAN_IN, U2576);
  nand ginst7716 (U7060, INSTQUEUE_REG_14__7__SCAN_IN, U2575);
  nand ginst7717 (U7061, INSTQUEUE_REG_15__7__SCAN_IN, U2574);
  nand ginst7718 (U7062, INSTQUEUE_REG_0__7__SCAN_IN, U2573);
  nand ginst7719 (U7063, INSTQUEUE_REG_1__7__SCAN_IN, U2572);
  nand ginst7720 (U7064, INSTQUEUE_REG_2__7__SCAN_IN, U2571);
  nand ginst7721 (U7065, INSTQUEUE_REG_3__7__SCAN_IN, U2570);
  nand ginst7722 (U7066, INSTQUEUE_REG_4__7__SCAN_IN, U2568);
  nand ginst7723 (U7067, INSTQUEUE_REG_5__7__SCAN_IN, U2567);
  nand ginst7724 (U7068, INSTQUEUE_REG_6__7__SCAN_IN, U2566);
  nand ginst7725 (U7069, INSTQUEUE_REG_7__7__SCAN_IN, U2565);
  nand ginst7726 (U7070, U4051, U4052, U4053, U4054);
  nand ginst7727 (U7071, U3408, U3412);
  nand ginst7728 (U7072, U4061, U4179);
  nand ginst7729 (U7073, U3409, U7072);
  nand ginst7730 (U7074, U3265, U4491);
  not ginst7731 (U7075, U3232);
  nand ginst7732 (U7076, U3381, U4142, U4388, U4491);
  nand ginst7733 (U7077, STATE2_REG_0__SCAN_IN, U4177);
  nand ginst7734 (U7078, U3232, U4055);
  not ginst7735 (U7079, U3438);
  nand ginst7736 (U7080, U3438, U5480, U7617);
  nand ginst7737 (U7081, U4182, U7080);
  not ginst7738 (U7082, U3437);
  nand ginst7739 (U7083, INSTQUEUEWR_ADDR_REG_3__SCAN_IN, U3284);
  nand ginst7740 (U7084, INSTQUEUERD_ADDR_REG_3__SCAN_IN, U3437);
  nand ginst7741 (U7085, U3347, U4191);
  nand ginst7742 (U7086, INSTQUEUE_REG_8__6__SCAN_IN, U2582);
  nand ginst7743 (U7087, INSTQUEUE_REG_9__6__SCAN_IN, U2581);
  nand ginst7744 (U7088, INSTQUEUE_REG_10__6__SCAN_IN, U2580);
  nand ginst7745 (U7089, INSTQUEUE_REG_11__6__SCAN_IN, U2579);
  nand ginst7746 (U7090, INSTQUEUE_REG_12__6__SCAN_IN, U2577);
  nand ginst7747 (U7091, INSTQUEUE_REG_13__6__SCAN_IN, U2576);
  nand ginst7748 (U7092, INSTQUEUE_REG_14__6__SCAN_IN, U2575);
  nand ginst7749 (U7093, INSTQUEUE_REG_15__6__SCAN_IN, U2574);
  nand ginst7750 (U7094, INSTQUEUE_REG_0__6__SCAN_IN, U2573);
  nand ginst7751 (U7095, INSTQUEUE_REG_1__6__SCAN_IN, U2572);
  nand ginst7752 (U7096, INSTQUEUE_REG_2__6__SCAN_IN, U2571);
  nand ginst7753 (U7097, INSTQUEUE_REG_3__6__SCAN_IN, U2570);
  nand ginst7754 (U7098, INSTQUEUE_REG_4__6__SCAN_IN, U2568);
  nand ginst7755 (U7099, INSTQUEUE_REG_5__6__SCAN_IN, U2567);
  nand ginst7756 (U7100, INSTQUEUE_REG_6__6__SCAN_IN, U2566);
  nand ginst7757 (U7101, INSTQUEUE_REG_7__6__SCAN_IN, U2565);
  nand ginst7758 (U7102, U4067, U4068, U4069, U4070);
  nand ginst7759 (U7103, INSTQUEUE_REG_8__5__SCAN_IN, U2582);
  nand ginst7760 (U7104, INSTQUEUE_REG_9__5__SCAN_IN, U2581);
  nand ginst7761 (U7105, INSTQUEUE_REG_10__5__SCAN_IN, U2580);
  nand ginst7762 (U7106, INSTQUEUE_REG_11__5__SCAN_IN, U2579);
  nand ginst7763 (U7107, INSTQUEUE_REG_12__5__SCAN_IN, U2577);
  nand ginst7764 (U7108, INSTQUEUE_REG_13__5__SCAN_IN, U2576);
  nand ginst7765 (U7109, INSTQUEUE_REG_14__5__SCAN_IN, U2575);
  nand ginst7766 (U7110, INSTQUEUE_REG_15__5__SCAN_IN, U2574);
  nand ginst7767 (U7111, INSTQUEUE_REG_0__5__SCAN_IN, U2573);
  nand ginst7768 (U7112, INSTQUEUE_REG_1__5__SCAN_IN, U2572);
  nand ginst7769 (U7113, INSTQUEUE_REG_2__5__SCAN_IN, U2571);
  nand ginst7770 (U7114, INSTQUEUE_REG_3__5__SCAN_IN, U2570);
  nand ginst7771 (U7115, INSTQUEUE_REG_4__5__SCAN_IN, U2568);
  nand ginst7772 (U7116, INSTQUEUE_REG_5__5__SCAN_IN, U2567);
  nand ginst7773 (U7117, INSTQUEUE_REG_6__5__SCAN_IN, U2566);
  nand ginst7774 (U7118, INSTQUEUE_REG_7__5__SCAN_IN, U2565);
  nand ginst7775 (U7119, U4071, U4072, U4073, U4074);
  nand ginst7776 (U7120, INSTQUEUE_REG_8__4__SCAN_IN, U2582);
  nand ginst7777 (U7121, INSTQUEUE_REG_9__4__SCAN_IN, U2581);
  nand ginst7778 (U7122, INSTQUEUE_REG_10__4__SCAN_IN, U2580);
  nand ginst7779 (U7123, INSTQUEUE_REG_11__4__SCAN_IN, U2579);
  nand ginst7780 (U7124, INSTQUEUE_REG_12__4__SCAN_IN, U2577);
  nand ginst7781 (U7125, INSTQUEUE_REG_13__4__SCAN_IN, U2576);
  nand ginst7782 (U7126, INSTQUEUE_REG_14__4__SCAN_IN, U2575);
  nand ginst7783 (U7127, INSTQUEUE_REG_15__4__SCAN_IN, U2574);
  nand ginst7784 (U7128, INSTQUEUE_REG_1__4__SCAN_IN, U2572);
  nand ginst7785 (U7129, INSTQUEUE_REG_2__4__SCAN_IN, U2571);
  nand ginst7786 (U7130, INSTQUEUE_REG_3__4__SCAN_IN, U2570);
  nand ginst7787 (U7131, INSTQUEUE_REG_4__4__SCAN_IN, U2568);
  nand ginst7788 (U7132, INSTQUEUE_REG_5__4__SCAN_IN, U2567);
  nand ginst7789 (U7133, INSTQUEUE_REG_6__4__SCAN_IN, U2566);
  nand ginst7790 (U7134, INSTQUEUE_REG_7__4__SCAN_IN, U2565);
  nand ginst7791 (U7135, INSTQUEUE_REG_8__3__SCAN_IN, U2582);
  nand ginst7792 (U7136, INSTQUEUE_REG_9__3__SCAN_IN, U2581);
  nand ginst7793 (U7137, INSTQUEUE_REG_10__3__SCAN_IN, U2580);
  nand ginst7794 (U7138, INSTQUEUE_REG_11__3__SCAN_IN, U2579);
  nand ginst7795 (U7139, INSTQUEUE_REG_12__3__SCAN_IN, U2577);
  nand ginst7796 (U7140, INSTQUEUE_REG_13__3__SCAN_IN, U2576);
  nand ginst7797 (U7141, INSTQUEUE_REG_14__3__SCAN_IN, U2575);
  nand ginst7798 (U7142, INSTQUEUE_REG_15__3__SCAN_IN, U2574);
  nand ginst7799 (U7143, INSTQUEUE_REG_0__3__SCAN_IN, U2573);
  nand ginst7800 (U7144, INSTQUEUE_REG_1__3__SCAN_IN, U2572);
  nand ginst7801 (U7145, INSTQUEUE_REG_2__3__SCAN_IN, U2571);
  nand ginst7802 (U7146, INSTQUEUE_REG_3__3__SCAN_IN, U2570);
  nand ginst7803 (U7147, INSTQUEUE_REG_4__3__SCAN_IN, U2568);
  nand ginst7804 (U7148, INSTQUEUE_REG_5__3__SCAN_IN, U2567);
  nand ginst7805 (U7149, INSTQUEUE_REG_6__3__SCAN_IN, U2566);
  nand ginst7806 (U7150, INSTQUEUE_REG_7__3__SCAN_IN, U2565);
  nand ginst7807 (U7151, U4080, U4081, U4082, U4083);
  nand ginst7808 (U7152, INSTQUEUE_REG_8__2__SCAN_IN, U2582);
  nand ginst7809 (U7153, INSTQUEUE_REG_9__2__SCAN_IN, U2581);
  nand ginst7810 (U7154, INSTQUEUE_REG_10__2__SCAN_IN, U2580);
  nand ginst7811 (U7155, INSTQUEUE_REG_11__2__SCAN_IN, U2579);
  nand ginst7812 (U7156, INSTQUEUE_REG_12__2__SCAN_IN, U2577);
  nand ginst7813 (U7157, INSTQUEUE_REG_13__2__SCAN_IN, U2576);
  nand ginst7814 (U7158, INSTQUEUE_REG_14__2__SCAN_IN, U2575);
  nand ginst7815 (U7159, INSTQUEUE_REG_15__2__SCAN_IN, U2574);
  nand ginst7816 (U7160, INSTQUEUE_REG_0__2__SCAN_IN, U2573);
  nand ginst7817 (U7161, INSTQUEUE_REG_1__2__SCAN_IN, U2572);
  nand ginst7818 (U7162, INSTQUEUE_REG_2__2__SCAN_IN, U2571);
  nand ginst7819 (U7163, INSTQUEUE_REG_3__2__SCAN_IN, U2570);
  nand ginst7820 (U7164, INSTQUEUE_REG_4__2__SCAN_IN, U2568);
  nand ginst7821 (U7165, INSTQUEUE_REG_5__2__SCAN_IN, U2567);
  nand ginst7822 (U7166, INSTQUEUE_REG_6__2__SCAN_IN, U2566);
  nand ginst7823 (U7167, INSTQUEUE_REG_7__2__SCAN_IN, U2565);
  nand ginst7824 (U7168, U4084, U4085, U4086, U4087);
  nand ginst7825 (U7169, INSTQUEUE_REG_8__1__SCAN_IN, U2582);
  nand ginst7826 (U7170, INSTQUEUE_REG_9__1__SCAN_IN, U2581);
  nand ginst7827 (U7171, INSTQUEUE_REG_10__1__SCAN_IN, U2580);
  nand ginst7828 (U7172, INSTQUEUE_REG_11__1__SCAN_IN, U2579);
  nand ginst7829 (U7173, INSTQUEUE_REG_12__1__SCAN_IN, U2577);
  nand ginst7830 (U7174, INSTQUEUE_REG_13__1__SCAN_IN, U2576);
  nand ginst7831 (U7175, INSTQUEUE_REG_14__1__SCAN_IN, U2575);
  nand ginst7832 (U7176, INSTQUEUE_REG_15__1__SCAN_IN, U2574);
  nand ginst7833 (U7177, INSTQUEUE_REG_0__1__SCAN_IN, U2573);
  nand ginst7834 (U7178, INSTQUEUE_REG_1__1__SCAN_IN, U2572);
  nand ginst7835 (U7179, INSTQUEUE_REG_2__1__SCAN_IN, U2571);
  nand ginst7836 (U7180, INSTQUEUE_REG_3__1__SCAN_IN, U2570);
  nand ginst7837 (U7181, INSTQUEUE_REG_4__1__SCAN_IN, U2568);
  nand ginst7838 (U7182, INSTQUEUE_REG_5__1__SCAN_IN, U2567);
  nand ginst7839 (U7183, INSTQUEUE_REG_6__1__SCAN_IN, U2566);
  nand ginst7840 (U7184, INSTQUEUE_REG_7__1__SCAN_IN, U2565);
  nand ginst7841 (U7185, U4088, U4089, U4090, U4091);
  nand ginst7842 (U7186, INSTQUEUE_REG_8__0__SCAN_IN, U2582);
  nand ginst7843 (U7187, INSTQUEUE_REG_9__0__SCAN_IN, U2581);
  nand ginst7844 (U7188, INSTQUEUE_REG_10__0__SCAN_IN, U2580);
  nand ginst7845 (U7189, INSTQUEUE_REG_11__0__SCAN_IN, U2579);
  nand ginst7846 (U7190, INSTQUEUE_REG_12__0__SCAN_IN, U2577);
  nand ginst7847 (U7191, INSTQUEUE_REG_13__0__SCAN_IN, U2576);
  nand ginst7848 (U7192, INSTQUEUE_REG_14__0__SCAN_IN, U2575);
  nand ginst7849 (U7193, INSTQUEUE_REG_15__0__SCAN_IN, U2574);
  nand ginst7850 (U7194, INSTQUEUE_REG_0__0__SCAN_IN, U2573);
  nand ginst7851 (U7195, INSTQUEUE_REG_1__0__SCAN_IN, U2572);
  nand ginst7852 (U7196, INSTQUEUE_REG_2__0__SCAN_IN, U2571);
  nand ginst7853 (U7197, INSTQUEUE_REG_3__0__SCAN_IN, U2570);
  nand ginst7854 (U7198, INSTQUEUE_REG_4__0__SCAN_IN, U2568);
  nand ginst7855 (U7199, INSTQUEUE_REG_5__0__SCAN_IN, U2567);
  nand ginst7856 (U7200, INSTQUEUE_REG_6__0__SCAN_IN, U2566);
  nand ginst7857 (U7201, INSTQUEUE_REG_7__0__SCAN_IN, U2565);
  nand ginst7858 (U7202, U4092, U4093, U4094, U4095);
  nand ginst7859 (U7203, INSTQUEUEWR_ADDR_REG_2__SCAN_IN, U3284);
  nand ginst7860 (U7204, U3442, U4191);
  nand ginst7861 (U7205, INSTQUEUEWR_ADDR_REG_1__SCAN_IN, U3284);
  nand ginst7862 (U7206, U3222, U4191);
  not ginst7863 (U7207, U4171);
  nand ginst7864 (U7208, INSTQUEUE_REG_8__7__SCAN_IN, U2602);
  nand ginst7865 (U7209, INSTQUEUE_REG_9__7__SCAN_IN, U2601);
  nand ginst7866 (U7210, INSTQUEUE_REG_10__7__SCAN_IN, U2600);
  nand ginst7867 (U7211, INSTQUEUE_REG_11__7__SCAN_IN, U2599);
  nand ginst7868 (U7212, INSTQUEUE_REG_12__7__SCAN_IN, U2597);
  nand ginst7869 (U7213, INSTQUEUE_REG_13__7__SCAN_IN, U2596);
  nand ginst7870 (U7214, INSTQUEUE_REG_14__7__SCAN_IN, U2595);
  nand ginst7871 (U7215, INSTQUEUE_REG_15__7__SCAN_IN, U2594);
  nand ginst7872 (U7216, INSTQUEUE_REG_0__7__SCAN_IN, U2592);
  nand ginst7873 (U7217, INSTQUEUE_REG_1__7__SCAN_IN, U2591);
  nand ginst7874 (U7218, INSTQUEUE_REG_2__7__SCAN_IN, U2590);
  nand ginst7875 (U7219, INSTQUEUE_REG_3__7__SCAN_IN, U2589);
  nand ginst7876 (U7220, INSTQUEUE_REG_4__7__SCAN_IN, U2587);
  nand ginst7877 (U7221, INSTQUEUE_REG_5__7__SCAN_IN, U2586);
  nand ginst7878 (U7222, INSTQUEUE_REG_6__7__SCAN_IN, U2585);
  nand ginst7879 (U7223, INSTQUEUE_REG_7__7__SCAN_IN, U2584);
  nand ginst7880 (U7224, U4109, U4110, U4111, U4112);
  nand ginst7881 (U7225, INSTQUEUE_REG_8__6__SCAN_IN, U2602);
  nand ginst7882 (U7226, INSTQUEUE_REG_9__6__SCAN_IN, U2601);
  nand ginst7883 (U7227, INSTQUEUE_REG_10__6__SCAN_IN, U2600);
  nand ginst7884 (U7228, INSTQUEUE_REG_11__6__SCAN_IN, U2599);
  nand ginst7885 (U7229, INSTQUEUE_REG_12__6__SCAN_IN, U2597);
  nand ginst7886 (U7230, INSTQUEUE_REG_13__6__SCAN_IN, U2596);
  nand ginst7887 (U7231, INSTQUEUE_REG_14__6__SCAN_IN, U2595);
  nand ginst7888 (U7232, INSTQUEUE_REG_15__6__SCAN_IN, U2594);
  nand ginst7889 (U7233, INSTQUEUE_REG_0__6__SCAN_IN, U2592);
  nand ginst7890 (U7234, INSTQUEUE_REG_1__6__SCAN_IN, U2591);
  nand ginst7891 (U7235, INSTQUEUE_REG_2__6__SCAN_IN, U2590);
  nand ginst7892 (U7236, INSTQUEUE_REG_3__6__SCAN_IN, U2589);
  nand ginst7893 (U7237, INSTQUEUE_REG_4__6__SCAN_IN, U2587);
  nand ginst7894 (U7238, INSTQUEUE_REG_5__6__SCAN_IN, U2586);
  nand ginst7895 (U7239, INSTQUEUE_REG_6__6__SCAN_IN, U2585);
  nand ginst7896 (U7240, INSTQUEUE_REG_7__6__SCAN_IN, U2584);
  nand ginst7897 (U7241, U4113, U4114, U4115, U4116);
  nand ginst7898 (U7242, INSTQUEUE_REG_8__5__SCAN_IN, U2602);
  nand ginst7899 (U7243, INSTQUEUE_REG_9__5__SCAN_IN, U2601);
  nand ginst7900 (U7244, INSTQUEUE_REG_10__5__SCAN_IN, U2600);
  nand ginst7901 (U7245, INSTQUEUE_REG_11__5__SCAN_IN, U2599);
  nand ginst7902 (U7246, INSTQUEUE_REG_12__5__SCAN_IN, U2597);
  nand ginst7903 (U7247, INSTQUEUE_REG_13__5__SCAN_IN, U2596);
  nand ginst7904 (U7248, INSTQUEUE_REG_14__5__SCAN_IN, U2595);
  nand ginst7905 (U7249, INSTQUEUE_REG_15__5__SCAN_IN, U2594);
  nand ginst7906 (U7250, INSTQUEUE_REG_0__5__SCAN_IN, U2592);
  nand ginst7907 (U7251, INSTQUEUE_REG_1__5__SCAN_IN, U2591);
  nand ginst7908 (U7252, INSTQUEUE_REG_2__5__SCAN_IN, U2590);
  nand ginst7909 (U7253, INSTQUEUE_REG_3__5__SCAN_IN, U2589);
  nand ginst7910 (U7254, INSTQUEUE_REG_4__5__SCAN_IN, U2587);
  nand ginst7911 (U7255, INSTQUEUE_REG_5__5__SCAN_IN, U2586);
  nand ginst7912 (U7256, INSTQUEUE_REG_6__5__SCAN_IN, U2585);
  nand ginst7913 (U7257, INSTQUEUE_REG_7__5__SCAN_IN, U2584);
  nand ginst7914 (U7258, U4117, U4118, U4119, U4120);
  nand ginst7915 (U7259, INSTQUEUE_REG_8__4__SCAN_IN, U2602);
  nand ginst7916 (U7260, INSTQUEUE_REG_9__4__SCAN_IN, U2601);
  nand ginst7917 (U7261, INSTQUEUE_REG_10__4__SCAN_IN, U2600);
  nand ginst7918 (U7262, INSTQUEUE_REG_11__4__SCAN_IN, U2599);
  nand ginst7919 (U7263, INSTQUEUE_REG_12__4__SCAN_IN, U2597);
  nand ginst7920 (U7264, INSTQUEUE_REG_13__4__SCAN_IN, U2596);
  nand ginst7921 (U7265, INSTQUEUE_REG_14__4__SCAN_IN, U2595);
  nand ginst7922 (U7266, INSTQUEUE_REG_15__4__SCAN_IN, U2594);
  nand ginst7923 (U7267, INSTQUEUE_REG_1__4__SCAN_IN, U2591);
  nand ginst7924 (U7268, INSTQUEUE_REG_2__4__SCAN_IN, U2590);
  nand ginst7925 (U7269, INSTQUEUE_REG_3__4__SCAN_IN, U2589);
  nand ginst7926 (U7270, INSTQUEUE_REG_4__4__SCAN_IN, U2587);
  nand ginst7927 (U7271, INSTQUEUE_REG_5__4__SCAN_IN, U2586);
  nand ginst7928 (U7272, INSTQUEUE_REG_6__4__SCAN_IN, U2585);
  nand ginst7929 (U7273, INSTQUEUE_REG_7__4__SCAN_IN, U2584);
  nand ginst7930 (U7274, INSTQUEUE_REG_8__3__SCAN_IN, U2602);
  nand ginst7931 (U7275, INSTQUEUE_REG_9__3__SCAN_IN, U2601);
  nand ginst7932 (U7276, INSTQUEUE_REG_10__3__SCAN_IN, U2600);
  nand ginst7933 (U7277, INSTQUEUE_REG_11__3__SCAN_IN, U2599);
  nand ginst7934 (U7278, INSTQUEUE_REG_12__3__SCAN_IN, U2597);
  nand ginst7935 (U7279, INSTQUEUE_REG_13__3__SCAN_IN, U2596);
  nand ginst7936 (U7280, INSTQUEUE_REG_14__3__SCAN_IN, U2595);
  nand ginst7937 (U7281, INSTQUEUE_REG_15__3__SCAN_IN, U2594);
  nand ginst7938 (U7282, INSTQUEUE_REG_0__3__SCAN_IN, U2592);
  nand ginst7939 (U7283, INSTQUEUE_REG_1__3__SCAN_IN, U2591);
  nand ginst7940 (U7284, INSTQUEUE_REG_2__3__SCAN_IN, U2590);
  nand ginst7941 (U7285, INSTQUEUE_REG_3__3__SCAN_IN, U2589);
  nand ginst7942 (U7286, INSTQUEUE_REG_4__3__SCAN_IN, U2587);
  nand ginst7943 (U7287, INSTQUEUE_REG_5__3__SCAN_IN, U2586);
  nand ginst7944 (U7288, INSTQUEUE_REG_6__3__SCAN_IN, U2585);
  nand ginst7945 (U7289, INSTQUEUE_REG_7__3__SCAN_IN, U2584);
  nand ginst7946 (U7290, U4125, U4126, U4127, U4128);
  nand ginst7947 (U7291, INSTQUEUE_REG_8__2__SCAN_IN, U2602);
  nand ginst7948 (U7292, INSTQUEUE_REG_9__2__SCAN_IN, U2601);
  nand ginst7949 (U7293, INSTQUEUE_REG_10__2__SCAN_IN, U2600);
  nand ginst7950 (U7294, INSTQUEUE_REG_11__2__SCAN_IN, U2599);
  nand ginst7951 (U7295, INSTQUEUE_REG_12__2__SCAN_IN, U2597);
  nand ginst7952 (U7296, INSTQUEUE_REG_13__2__SCAN_IN, U2596);
  nand ginst7953 (U7297, INSTQUEUE_REG_14__2__SCAN_IN, U2595);
  nand ginst7954 (U7298, INSTQUEUE_REG_15__2__SCAN_IN, U2594);
  nand ginst7955 (U7299, INSTQUEUE_REG_0__2__SCAN_IN, U2592);
  nand ginst7956 (U7300, INSTQUEUE_REG_1__2__SCAN_IN, U2591);
  nand ginst7957 (U7301, INSTQUEUE_REG_2__2__SCAN_IN, U2590);
  nand ginst7958 (U7302, INSTQUEUE_REG_3__2__SCAN_IN, U2589);
  nand ginst7959 (U7303, INSTQUEUE_REG_4__2__SCAN_IN, U2587);
  nand ginst7960 (U7304, INSTQUEUE_REG_5__2__SCAN_IN, U2586);
  nand ginst7961 (U7305, INSTQUEUE_REG_6__2__SCAN_IN, U2585);
  nand ginst7962 (U7306, INSTQUEUE_REG_7__2__SCAN_IN, U2584);
  nand ginst7963 (U7307, U4129, U4130, U4131, U4132);
  nand ginst7964 (U7308, INSTQUEUE_REG_8__1__SCAN_IN, U2602);
  nand ginst7965 (U7309, INSTQUEUE_REG_9__1__SCAN_IN, U2601);
  nand ginst7966 (U7310, INSTQUEUE_REG_10__1__SCAN_IN, U2600);
  nand ginst7967 (U7311, INSTQUEUE_REG_11__1__SCAN_IN, U2599);
  nand ginst7968 (U7312, INSTQUEUE_REG_12__1__SCAN_IN, U2597);
  nand ginst7969 (U7313, INSTQUEUE_REG_13__1__SCAN_IN, U2596);
  nand ginst7970 (U7314, INSTQUEUE_REG_14__1__SCAN_IN, U2595);
  nand ginst7971 (U7315, INSTQUEUE_REG_15__1__SCAN_IN, U2594);
  nand ginst7972 (U7316, INSTQUEUE_REG_0__1__SCAN_IN, U2592);
  nand ginst7973 (U7317, INSTQUEUE_REG_1__1__SCAN_IN, U2591);
  nand ginst7974 (U7318, INSTQUEUE_REG_2__1__SCAN_IN, U2590);
  nand ginst7975 (U7319, INSTQUEUE_REG_3__1__SCAN_IN, U2589);
  nand ginst7976 (U7320, INSTQUEUE_REG_4__1__SCAN_IN, U2587);
  nand ginst7977 (U7321, INSTQUEUE_REG_5__1__SCAN_IN, U2586);
  nand ginst7978 (U7322, INSTQUEUE_REG_6__1__SCAN_IN, U2585);
  nand ginst7979 (U7323, INSTQUEUE_REG_7__1__SCAN_IN, U2584);
  nand ginst7980 (U7324, U4133, U4134, U4135, U4136);
  nand ginst7981 (U7325, INSTQUEUE_REG_8__0__SCAN_IN, U2602);
  nand ginst7982 (U7326, INSTQUEUE_REG_9__0__SCAN_IN, U2601);
  nand ginst7983 (U7327, INSTQUEUE_REG_10__0__SCAN_IN, U2600);
  nand ginst7984 (U7328, INSTQUEUE_REG_11__0__SCAN_IN, U2599);
  nand ginst7985 (U7329, INSTQUEUE_REG_12__0__SCAN_IN, U2597);
  nand ginst7986 (U7330, INSTQUEUE_REG_13__0__SCAN_IN, U2596);
  nand ginst7987 (U7331, INSTQUEUE_REG_14__0__SCAN_IN, U2595);
  nand ginst7988 (U7332, INSTQUEUE_REG_15__0__SCAN_IN, U2594);
  nand ginst7989 (U7333, INSTQUEUE_REG_0__0__SCAN_IN, U2592);
  nand ginst7990 (U7334, INSTQUEUE_REG_1__0__SCAN_IN, U2591);
  nand ginst7991 (U7335, INSTQUEUE_REG_2__0__SCAN_IN, U2590);
  nand ginst7992 (U7336, INSTQUEUE_REG_3__0__SCAN_IN, U2589);
  nand ginst7993 (U7337, INSTQUEUE_REG_4__0__SCAN_IN, U2587);
  nand ginst7994 (U7338, INSTQUEUE_REG_5__0__SCAN_IN, U2586);
  nand ginst7995 (U7339, INSTQUEUE_REG_6__0__SCAN_IN, U2585);
  nand ginst7996 (U7340, INSTQUEUE_REG_7__0__SCAN_IN, U2584);
  nand ginst7997 (U7341, U4137, U4138, U4139, U4140);
  nand ginst7998 (U7342, U2354, U4219, U4222);
  nand ginst7999 (U7343, U4141, U7075);
  nand ginst8000 (U7344, U3383, U3397);
  nand ginst8001 (U7345, U4222, U7344);
  nand ginst8002 (U7346, U2452, U4178);
  nand ginst8003 (U7347, U3258, U7343);
  nand ginst8004 (U7348, U4196, U7076);
  nand ginst8005 (U7349, U4148, U4196);
  nand ginst8006 (U7350, U2451, U4198);
  nand ginst8007 (U7351, U3407, U3421, U4183, U7349, U7350);
  nand ginst8008 (U7352, R2238_U6, U7351);
  nand ginst8009 (U7353, SUB_450_U6, U2354);
  nand ginst8010 (U7354, R2238_U19, U7351);
  nand ginst8011 (U7355, SUB_450_U19, U2354);
  nand ginst8012 (U7356, R2238_U20, U7351);
  nand ginst8013 (U7357, SUB_450_U20, U2354);
  nand ginst8014 (U7358, R2238_U21, U7351);
  nand ginst8015 (U7359, SUB_450_U21, U2354);
  nand ginst8016 (U7360, R2238_U22, U7351);
  nand ginst8017 (U7361, SUB_450_U22, U2354);
  nand ginst8018 (U7362, R2238_U7, U7351);
  nand ginst8019 (U7363, SUB_450_U7, U2354);
  nand ginst8020 (U7364, R2238_U19, U4180);
  nand ginst8021 (U7365, INSTQUEUERD_ADDR_REG_4__SCAN_IN, U3281);
  nand ginst8022 (U7366, R2238_U20, U4180);
  nand ginst8023 (U7367, INSTQUEUERD_ADDR_REG_3__SCAN_IN, U3281);
  nand ginst8024 (U7368, STATE2_REG_0__SCAN_IN, U4161);
  nand ginst8025 (U7369, U3407, U7368);
  nand ginst8026 (U7370, R2238_U21, U4180);
  nand ginst8027 (U7371, INSTQUEUERD_ADDR_REG_2__SCAN_IN, U3281);
  nand ginst8028 (U7372, U2450, U3258);
  nand ginst8029 (U7373, R2238_U22, U4180);
  nand ginst8030 (U7374, INSTQUEUERD_ADDR_REG_1__SCAN_IN, U3281);
  nand ginst8031 (U7375, U2451, U3271);
  nand ginst8032 (U7376, R2238_U7, U4180);
  nand ginst8033 (U7377, INSTQUEUERD_ADDR_REG_0__SCAN_IN, U3281);
  nand ginst8034 (U7378, U3277, U3380);
  nand ginst8035 (U7379, U3271, U3436);
  nand ginst8036 (U7380, INSTADDRPOINTER_REG_9__SCAN_IN, U7379);
  nand ginst8037 (U7381, EBX_REG_9__SCAN_IN, U7378);
  nand ginst8038 (U7382, INSTADDRPOINTER_REG_8__SCAN_IN, U7379);
  nand ginst8039 (U7383, EBX_REG_8__SCAN_IN, U7378);
  nand ginst8040 (U7384, INSTADDRPOINTER_REG_7__SCAN_IN, U7379);
  nand ginst8041 (U7385, EBX_REG_7__SCAN_IN, U7378);
  nand ginst8042 (U7386, INSTADDRPOINTER_REG_6__SCAN_IN, U7379);
  nand ginst8043 (U7387, EBX_REG_6__SCAN_IN, U7378);
  nand ginst8044 (U7388, INSTADDRPOINTER_REG_5__SCAN_IN, U7379);
  nand ginst8045 (U7389, EBX_REG_5__SCAN_IN, U7378);
  nand ginst8046 (U7390, INSTADDRPOINTER_REG_4__SCAN_IN, U7379);
  nand ginst8047 (U7391, EBX_REG_4__SCAN_IN, U7378);
  nand ginst8048 (U7392, INSTADDRPOINTER_REG_31__SCAN_IN, U7379);
  nand ginst8049 (U7393, EBX_REG_31__SCAN_IN, U7378);
  nand ginst8050 (U7394, INSTADDRPOINTER_REG_30__SCAN_IN, U7379);
  nand ginst8051 (U7395, EBX_REG_30__SCAN_IN, U7378);
  nand ginst8052 (U7396, INSTADDRPOINTER_REG_3__SCAN_IN, U7379);
  nand ginst8053 (U7397, EBX_REG_3__SCAN_IN, U7378);
  nand ginst8054 (U7398, INSTADDRPOINTER_REG_29__SCAN_IN, U7379);
  nand ginst8055 (U7399, EBX_REG_29__SCAN_IN, U7378);
  nand ginst8056 (U7400, INSTADDRPOINTER_REG_28__SCAN_IN, U7379);
  nand ginst8057 (U7401, EBX_REG_28__SCAN_IN, U7378);
  nand ginst8058 (U7402, INSTADDRPOINTER_REG_27__SCAN_IN, U7379);
  nand ginst8059 (U7403, EBX_REG_27__SCAN_IN, U7378);
  nand ginst8060 (U7404, INSTADDRPOINTER_REG_26__SCAN_IN, U7379);
  nand ginst8061 (U7405, EBX_REG_26__SCAN_IN, U7378);
  nand ginst8062 (U7406, INSTADDRPOINTER_REG_25__SCAN_IN, U7379);
  nand ginst8063 (U7407, EBX_REG_25__SCAN_IN, U7378);
  nand ginst8064 (U7408, INSTADDRPOINTER_REG_24__SCAN_IN, U7379);
  nand ginst8065 (U7409, EBX_REG_24__SCAN_IN, U7378);
  nand ginst8066 (U7410, INSTADDRPOINTER_REG_23__SCAN_IN, U7379);
  nand ginst8067 (U7411, EBX_REG_23__SCAN_IN, U7378);
  nand ginst8068 (U7412, INSTADDRPOINTER_REG_22__SCAN_IN, U7379);
  nand ginst8069 (U7413, EBX_REG_22__SCAN_IN, U7378);
  nand ginst8070 (U7414, INSTADDRPOINTER_REG_21__SCAN_IN, U7379);
  nand ginst8071 (U7415, EBX_REG_21__SCAN_IN, U7378);
  nand ginst8072 (U7416, INSTADDRPOINTER_REG_20__SCAN_IN, U7379);
  nand ginst8073 (U7417, EBX_REG_20__SCAN_IN, U7378);
  nand ginst8074 (U7418, INSTADDRPOINTER_REG_2__SCAN_IN, U7379);
  nand ginst8075 (U7419, EBX_REG_2__SCAN_IN, U7378);
  nand ginst8076 (U7420, INSTADDRPOINTER_REG_19__SCAN_IN, U7379);
  nand ginst8077 (U7421, EBX_REG_19__SCAN_IN, U7378);
  nand ginst8078 (U7422, INSTADDRPOINTER_REG_18__SCAN_IN, U7379);
  nand ginst8079 (U7423, EBX_REG_18__SCAN_IN, U7378);
  nand ginst8080 (U7424, INSTADDRPOINTER_REG_17__SCAN_IN, U7379);
  nand ginst8081 (U7425, EBX_REG_17__SCAN_IN, U7378);
  nand ginst8082 (U7426, INSTADDRPOINTER_REG_16__SCAN_IN, U7379);
  nand ginst8083 (U7427, EBX_REG_16__SCAN_IN, U7378);
  nand ginst8084 (U7428, INSTADDRPOINTER_REG_15__SCAN_IN, U7379);
  nand ginst8085 (U7429, EBX_REG_15__SCAN_IN, U7378);
  nand ginst8086 (U7430, INSTADDRPOINTER_REG_14__SCAN_IN, U7379);
  nand ginst8087 (U7431, EBX_REG_14__SCAN_IN, U7378);
  nand ginst8088 (U7432, INSTADDRPOINTER_REG_13__SCAN_IN, U7379);
  nand ginst8089 (U7433, EBX_REG_13__SCAN_IN, U7378);
  nand ginst8090 (U7434, INSTADDRPOINTER_REG_12__SCAN_IN, U7379);
  nand ginst8091 (U7435, EBX_REG_12__SCAN_IN, U7378);
  nand ginst8092 (U7436, INSTADDRPOINTER_REG_11__SCAN_IN, U7379);
  nand ginst8093 (U7437, EBX_REG_11__SCAN_IN, U7378);
  nand ginst8094 (U7438, INSTADDRPOINTER_REG_10__SCAN_IN, U7379);
  nand ginst8095 (U7439, EBX_REG_10__SCAN_IN, U7378);
  nand ginst8096 (U7440, INSTADDRPOINTER_REG_1__SCAN_IN, U7379);
  nand ginst8097 (U7441, EBX_REG_1__SCAN_IN, U7378);
  nand ginst8098 (U7442, INSTADDRPOINTER_REG_0__SCAN_IN, U7379);
  nand ginst8099 (U7443, EBX_REG_0__SCAN_IN, U7378);
  nand ginst8100 (U7444, U4465, U4484);
  nand ginst8101 (U7445, INSTQUEUERD_ADDR_REG_4__SCAN_IN, U2430);
  nand ginst8102 (U7446, U3249, U3476);
  nand ginst8103 (U7447, INSTQUEUERD_ADDR_REG_3__SCAN_IN, U2430);
  nand ginst8104 (U7448, U3249, U3477);
  nand ginst8105 (U7449, FLUSH_REG_SCAN_IN, U2446, U3457);
  nand ginst8106 (U7450, INSTQUEUERD_ADDR_REG_2__SCAN_IN, U2430);
  nand ginst8107 (U7451, U3249, U3478);
  nand ginst8108 (U7452, FLUSH_REG_SCAN_IN, U2446, U7700);
  nand ginst8109 (U7453, INSTQUEUERD_ADDR_REG_1__SCAN_IN, U2430);
  nand ginst8110 (U7454, U3249, U3479);
  nand ginst8111 (U7455, INSTQUEUERD_ADDR_REG_0__SCAN_IN, U2430);
  nand ginst8112 (U7456, STATE_REG_0__SCAN_IN, U4173);
  or ginst8113 (U7457, READY_N, STATE2_REG_2__SCAN_IN);
  nand ginst8114 (U7458, U4098, U7206);
  nand ginst8115 (U7459, U3409, U7072);
  nand ginst8116 (U7460, STATE2_REG_0__SCAN_IN, U4199);
  nand ginst8117 (U7461, STATE2_REG_0__SCAN_IN, U4200);
  nand ginst8118 (U7462, STATE2_REG_0__SCAN_IN, U4201);
  nand ginst8119 (U7463, STATE2_REG_0__SCAN_IN, U4224);
  nand ginst8120 (U7464, STATE2_REG_0__SCAN_IN, U4252);
  nand ginst8121 (U7465, STATE2_REG_0__SCAN_IN, U7620);
  nand ginst8122 (U7466, U2608, U3253);
  nand ginst8123 (U7467, U4105, U4106, U4108, U7081);
  nand ginst8124 (U7468, STATE2_REG_0__SCAN_IN, U7620);
  nand ginst8125 (U7469, U2379, U3416);
  nand ginst8126 (U7470, U2369, U6355);
  nand ginst8127 (U7471, U2369, U3876);
  nand ginst8128 (U7472, U4217, U7469, U7470);
  nand ginst8129 (U7473, U4218, U7471);
  nand ginst8130 (U7474, U4159, U4182, U5479);
  nand ginst8131 (U7475, U4182, U7079);
  nand ginst8132 (U7476, U3379, U4182);
  nand ginst8133 (U7477, STATE2_REG_0__SCAN_IN, U4224);
  nand ginst8134 (U7478, U4060, U7772, U7773);
  nand ginst8135 (U7479, U4096, U7204);
  nand ginst8136 (U7480, U4097, U7082);
  not ginst8137 (U7481, U3266);
  not ginst8138 (U7482, U3263);
  nand ginst8139 (U7483, U2607, U4056, U4057, U4058, U4059);
  nand ginst8140 (U7484, U3722, U7481);
  nand ginst8141 (U7485, U3723, U5457);
  nand ginst8142 (U7486, U2425, U7481);
  nand ginst8143 (U7487, U2425, U7481);
  nand ginst8144 (U7488, U6348, U6349, U7487);
  nand ginst8145 (U7489, R2167_U17, U7481);
  nand ginst8146 (U7490, R2167_U17, U4189, U7481);
  nand ginst8147 (U7491, U6137, U7490);
  nand ginst8148 (U7492, U7073, U7481);
  nand ginst8149 (U7493, U7459, U7481);
  nand ginst8150 (U7494, U4102, U4103, U4104);
  nand ginst8151 (U7495, U3747, U7481);
  nand ginst8152 (U7496, U3748, U3749, U5553);
  nand ginst8153 (U7497, U2519, U3734);
  nand ginst8154 (U7498, U5950, U7481);
  nand ginst8155 (U7499, U5953, U7481);
  nand ginst8156 (U7500, U5956, U7481);
  nand ginst8157 (U7501, U5959, U7481);
  nand ginst8158 (U7502, U5962, U7481);
  nand ginst8159 (U7503, U5965, U7481);
  nand ginst8160 (U7504, U5968, U7481);
  nand ginst8161 (U7505, U5971, U7481);
  nand ginst8162 (U7506, U5974, U7481);
  nand ginst8163 (U7507, U5977, U7481);
  nand ginst8164 (U7508, U5980, U7481);
  nand ginst8165 (U7509, U5983, U7481);
  nand ginst8166 (U7510, U5986, U7481);
  nand ginst8167 (U7511, U5989, U7481);
  nand ginst8168 (U7512, U5992, U7481);
  nand ginst8169 (U7513, U5995, U7481);
  nand ginst8170 (U7514, U5998, U7481);
  nand ginst8171 (U7515, U6001, U7481);
  nand ginst8172 (U7516, U6004, U7481);
  nand ginst8173 (U7517, U6007, U7481);
  nand ginst8174 (U7518, U6010, U7481);
  nand ginst8175 (U7519, U6013, U7481);
  nand ginst8176 (U7520, U6016, U7481);
  nand ginst8177 (U7521, U6019, U7481);
  nand ginst8178 (U7522, U6022, U7481);
  nand ginst8179 (U7523, U6025, U7481);
  nand ginst8180 (U7524, U6028, U7481);
  nand ginst8181 (U7525, U6031, U7481);
  nand ginst8182 (U7526, U6034, U7481);
  nand ginst8183 (U7527, U6037, U7481);
  nand ginst8184 (U7528, U6040, U7481);
  nand ginst8185 (U7529, U2357, U7481);
  nand ginst8186 (U7530, UWORD_REG_0__SCAN_IN, U7529);
  nand ginst8187 (U7531, U2357, U7481);
  nand ginst8188 (U7532, UWORD_REG_1__SCAN_IN, U7531);
  nand ginst8189 (U7533, U2357, U7481);
  nand ginst8190 (U7534, UWORD_REG_2__SCAN_IN, U7533);
  nand ginst8191 (U7535, U2357, U7481);
  nand ginst8192 (U7536, UWORD_REG_3__SCAN_IN, U7535);
  nand ginst8193 (U7537, U2357, U7481);
  nand ginst8194 (U7538, UWORD_REG_4__SCAN_IN, U7537);
  nand ginst8195 (U7539, U2357, U7481);
  nand ginst8196 (U7540, UWORD_REG_5__SCAN_IN, U7539);
  nand ginst8197 (U7541, U2357, U7481);
  nand ginst8198 (U7542, UWORD_REG_6__SCAN_IN, U7541);
  nand ginst8199 (U7543, U2357, U7481);
  nand ginst8200 (U7544, UWORD_REG_7__SCAN_IN, U7543);
  nand ginst8201 (U7545, U2357, U7481);
  nand ginst8202 (U7546, UWORD_REG_8__SCAN_IN, U7545);
  nand ginst8203 (U7547, U2357, U7481);
  nand ginst8204 (U7548, UWORD_REG_9__SCAN_IN, U7547);
  nand ginst8205 (U7549, U2357, U7481);
  nand ginst8206 (U7550, UWORD_REG_10__SCAN_IN, U7549);
  nand ginst8207 (U7551, U2357, U7481);
  nand ginst8208 (U7552, UWORD_REG_11__SCAN_IN, U7551);
  nand ginst8209 (U7553, U2357, U7481);
  nand ginst8210 (U7554, UWORD_REG_12__SCAN_IN, U7553);
  nand ginst8211 (U7555, U2357, U7481);
  nand ginst8212 (U7556, UWORD_REG_13__SCAN_IN, U7555);
  nand ginst8213 (U7557, U2357, U7481);
  nand ginst8214 (U7558, UWORD_REG_14__SCAN_IN, U7557);
  nand ginst8215 (U7559, U2357, U7481);
  nand ginst8216 (U7560, LWORD_REG_0__SCAN_IN, U7559);
  nand ginst8217 (U7561, U2357, U7481);
  nand ginst8218 (U7562, LWORD_REG_1__SCAN_IN, U7561);
  nand ginst8219 (U7563, U2357, U7481);
  nand ginst8220 (U7564, LWORD_REG_2__SCAN_IN, U7563);
  nand ginst8221 (U7565, U2357, U7481);
  nand ginst8222 (U7566, LWORD_REG_3__SCAN_IN, U7565);
  nand ginst8223 (U7567, U2357, U7481);
  nand ginst8224 (U7568, LWORD_REG_4__SCAN_IN, U7567);
  nand ginst8225 (U7569, U2357, U7481);
  nand ginst8226 (U7570, LWORD_REG_5__SCAN_IN, U7569);
  nand ginst8227 (U7571, U2357, U7481);
  nand ginst8228 (U7572, LWORD_REG_6__SCAN_IN, U7571);
  nand ginst8229 (U7573, U2357, U7481);
  nand ginst8230 (U7574, LWORD_REG_7__SCAN_IN, U7573);
  nand ginst8231 (U7575, U2357, U7481);
  nand ginst8232 (U7576, LWORD_REG_8__SCAN_IN, U7575);
  nand ginst8233 (U7577, U2357, U7481);
  nand ginst8234 (U7578, LWORD_REG_9__SCAN_IN, U7577);
  nand ginst8235 (U7579, U2357, U7481);
  nand ginst8236 (U7580, LWORD_REG_10__SCAN_IN, U7579);
  nand ginst8237 (U7581, U2357, U7481);
  nand ginst8238 (U7582, LWORD_REG_11__SCAN_IN, U7581);
  nand ginst8239 (U7583, U2357, U7481);
  nand ginst8240 (U7584, LWORD_REG_12__SCAN_IN, U7583);
  nand ginst8241 (U7585, U2357, U7481);
  nand ginst8242 (U7586, LWORD_REG_13__SCAN_IN, U7585);
  nand ginst8243 (U7587, U2357, U7481);
  nand ginst8244 (U7588, LWORD_REG_14__SCAN_IN, U7587);
  nand ginst8245 (U7589, U2357, U7481);
  nand ginst8246 (U7590, LWORD_REG_15__SCAN_IN, U7589);
  nand ginst8247 (U7591, U3556, U4247, U7481);
  nand ginst8248 (U7592, U3569, U7671, U7672);
  nand ginst8249 (U7593, U3855, U7481);
  nand ginst8250 (U7594, U3415, U7593);
  nand ginst8251 (U7595, U4196, U7481);
  nand ginst8252 (U7596, U3434, U7595);
  nand ginst8253 (U7597, U3266, U3387);
  nand ginst8254 (U7598, U3742, U7481);
  nand ginst8255 (U7599, U3743, U7598);
  nand ginst8256 (U7600, INSTQUEUE_REG_0__4__SCAN_IN, U5404);
  nand ginst8257 (U7601, INSTQUEUE_REG_0__4__SCAN_IN, U2523);
  nand ginst8258 (U7602, INSTQUEUE_REG_0__4__SCAN_IN, U2546);
  nand ginst8259 (U7603, U4037, U4038, U4039, U4040);
  nand ginst8260 (U7604, INSTQUEUE_REG_0__4__SCAN_IN, U4180);
  nand ginst8261 (U7605, INSTQUEUE_REG_0__4__SCAN_IN, U2573);
  nand ginst8262 (U7606, U4075, U4076, U4077, U4079);
  nand ginst8263 (U7607, INSTQUEUE_REG_0__4__SCAN_IN, U2592);
  nand ginst8264 (U7608, U4121, U4122, U4123, U4124);
  not ginst8265 (U7609, U3246);
  nand ginst8266 (U7610, U3248, U7609);
  nand ginst8267 (U7611, STATE_REG_1__SCAN_IN, U4346, U4349);
  nand ginst8268 (U7612, STATE_REG_2__SCAN_IN, U7456);
  nand ginst8269 (U7613, STATE_REG_1__SCAN_IN, U4346);
  nand ginst8270 (U7614, U4490, U4498);
  nand ginst8271 (U7615, U4159, U5475);
  nand ginst8272 (U7616, U3270, U3276);
  not ginst8273 (U7617, U3379);
  nand ginst8274 (U7618, U4196, U7478);
  nand ginst8275 (U7619, U4159, U5475);
  nand ginst8276 (U7620, U7618, U7619);
  nand ginst8277 (U7621, BE_N_REG_3__SCAN_IN, U3236);
  nand ginst8278 (U7622, BYTEENABLE_REG_3__SCAN_IN, U4209);
  nand ginst8279 (U7623, BE_N_REG_2__SCAN_IN, U3236);
  nand ginst8280 (U7624, BYTEENABLE_REG_2__SCAN_IN, U4209);
  nand ginst8281 (U7625, BE_N_REG_1__SCAN_IN, U3236);
  nand ginst8282 (U7626, BYTEENABLE_REG_1__SCAN_IN, U4209);
  nand ginst8283 (U7627, BE_N_REG_0__SCAN_IN, U3236);
  nand ginst8284 (U7628, BYTEENABLE_REG_0__SCAN_IN, U4209);
  nand ginst8285 (U7629, REQUESTPENDING_REG_SCAN_IN, STATE_REG_0__SCAN_IN, U3238);
  nand ginst8286 (U7630, STATE_REG_2__SCAN_IN, U3246);
  nand ginst8287 (U7631, U7629, U7630);
  nand ginst8288 (U7632, STATE_REG_1__SCAN_IN, U4349, U7612);
  nand ginst8289 (U7633, U3235, U7631);
  nand ginst8290 (U7634, STATE_REG_2__SCAN_IN, STATE_REG_0__SCAN_IN, U3247);
  nand ginst8291 (U7635, U3238, U4359);
  or ginst8292 (U7636, STATE_REG_1__SCAN_IN, STATE_REG_0__SCAN_IN);
  nand ginst8293 (U7637, STATE_REG_0__SCAN_IN, U4246);
  not ginst8294 (U7638, U3449);
  nand ginst8295 (U7639, DATAWIDTH_REG_0__SCAN_IN, U7638);
  nand ginst8296 (U7640, U3449, U3450);
  nand ginst8297 (U7641, U3449, U4364);
  nand ginst8298 (U7642, DATAWIDTH_REG_1__SCAN_IN, U7638);
  nand ginst8299 (U7643, U3252, U3528, U3529);
  nand ginst8300 (U7644, INSTQUEUE_REG_7__4__SCAN_IN, INSTQUEUERD_ADDR_REG_2__SCAN_IN, INSTQUEUERD_ADDR_REG_1__SCAN_IN, INSTQUEUERD_ADDR_REG_0__SCAN_IN, U3257);
  nand ginst8301 (U7645, INSTQUEUE_REG_5__4__SCAN_IN, INSTQUEUERD_ADDR_REG_2__SCAN_IN, INSTQUEUERD_ADDR_REG_0__SCAN_IN, U3252, U3257);
  nand ginst8302 (U7646, INSTQUEUE_REG_2__4__SCAN_IN, INSTQUEUERD_ADDR_REG_1__SCAN_IN, U3251, U3253, U3257);
  nand ginst8303 (U7647, U3257, U3530, U3531);
  nand ginst8304 (U7648, INSTQUEUERD_ADDR_REG_3__SCAN_IN, U3532, U3533);
  nand ginst8305 (U7649, U3252, U3534, U3535);
  nand ginst8306 (U7650, INSTQUEUERD_ADDR_REG_1__SCAN_IN, U3536, U3537);
  nand ginst8307 (U7651, U3253, U3538, U3539);
  nand ginst8308 (U7652, INSTQUEUE_REG_15__4__SCAN_IN, INSTQUEUERD_ADDR_REG_3__SCAN_IN, INSTQUEUERD_ADDR_REG_2__SCAN_IN, INSTQUEUERD_ADDR_REG_1__SCAN_IN, INSTQUEUERD_ADDR_REG_0__SCAN_IN);
  nand ginst8309 (U7653, INSTQUEUE_REG_0__4__SCAN_IN, U3251, U3252, U3253, U3257);
  nand ginst8310 (U7654, INSTQUEUE_REG_8__4__SCAN_IN, INSTQUEUERD_ADDR_REG_3__SCAN_IN, U3251, U3252, U3253);
  nand ginst8311 (U7655, INSTQUEUE_REG_10__4__SCAN_IN, INSTQUEUERD_ADDR_REG_3__SCAN_IN, INSTQUEUERD_ADDR_REG_1__SCAN_IN, U3251, U3253);
  nand ginst8312 (U7656, INSTQUEUERD_ADDR_REG_0__SCAN_IN, U3540, U3541);
  nand ginst8313 (U7657, INSTQUEUE_REG_3__4__SCAN_IN, INSTQUEUERD_ADDR_REG_1__SCAN_IN, INSTQUEUERD_ADDR_REG_0__SCAN_IN, U3251, U3257);
  nand ginst8314 (U7658, INSTQUEUE_REG_11__4__SCAN_IN, INSTQUEUERD_ADDR_REG_3__SCAN_IN, INSTQUEUERD_ADDR_REG_1__SCAN_IN, INSTQUEUERD_ADDR_REG_0__SCAN_IN, U3251);
  nand ginst8315 (U7659, INSTQUEUE_REG_3__5__SCAN_IN, INSTQUEUERD_ADDR_REG_1__SCAN_IN, INSTQUEUERD_ADDR_REG_0__SCAN_IN, U3251, U3257);
  nand ginst8316 (U7660, INSTQUEUERD_ADDR_REG_3__SCAN_IN, U3516, U3517);
  nand ginst8317 (U7661, INSTQUEUE_REG_9__6__SCAN_IN, INSTQUEUERD_ADDR_REG_3__SCAN_IN, INSTQUEUERD_ADDR_REG_0__SCAN_IN, U3251, U3252);
  nand ginst8318 (U7662, INSTQUEUERD_ADDR_REG_1__SCAN_IN, U3522, U3523);
  nand ginst8319 (U7663, INSTQUEUE_REG_10__6__SCAN_IN, INSTQUEUERD_ADDR_REG_3__SCAN_IN, INSTQUEUERD_ADDR_REG_1__SCAN_IN, U3251, U3253);
  nand ginst8320 (U7664, INSTQUEUE_REG_11__6__SCAN_IN, INSTQUEUERD_ADDR_REG_3__SCAN_IN, INSTQUEUERD_ADDR_REG_1__SCAN_IN, INSTQUEUERD_ADDR_REG_0__SCAN_IN, U3251);
  nand ginst8321 (U7665, INSTQUEUE_REG_0__6__SCAN_IN, U3251, U3252, U3253, U3257);
  nand ginst8322 (U7666, INSTQUEUE_REG_8__6__SCAN_IN, INSTQUEUERD_ADDR_REG_3__SCAN_IN, U3251, U3252, U3253);
  nand ginst8323 (U7667, U3424, U4482);
  nand ginst8324 (U7668, U3271, U7489);
  nand ginst8325 (U7669, R2167_U17, U4204);
  nand ginst8326 (U7670, U3260, U4494);
  nand ginst8327 (U7671, STATE2_REG_0__SCAN_IN, U4500);
  nand ginst8328 (U7672, U3281, U4501);
  nand ginst8329 (U7673, STATE2_REG_3__SCAN_IN, U3282);
  nand ginst8330 (U7674, U2428, U4502);
  or ginst8331 (U7675, STATEBS16_REG_SCAN_IN, STATE2_REG_0__SCAN_IN);
  nand ginst8332 (U7676, STATE2_REG_0__SCAN_IN, U7457);
  nand ginst8333 (U7677, STATE2_REG_0__SCAN_IN, U4510);
  nand ginst8334 (U7678, U3281, U4509, U7592);
  nand ginst8335 (U7679, R2144_U49, U3300);
  nand ginst8336 (U7680, U3298, U4516);
  not ginst8337 (U7681, U3441);
  nand ginst8338 (U7682, INSTQUEUEWR_ADDR_REG_2__SCAN_IN, U3292);
  nand ginst8339 (U7683, U3291, U4521);
  not ginst8340 (U7684, U3442);
  nand ginst8341 (U7685, U3260, U4204);
  nand ginst8342 (U7686, R2167_U17, U7485);
  nand ginst8343 (U7687, U4420, U5454);
  nand ginst8344 (U7688, U4159, U5455);
  nand ginst8345 (U7689, U3454, U4160);
  nand ginst8346 (U7690, INSTQUEUERD_ADDR_REG_4__SCAN_IN, U5464);
  nand ginst8347 (U7691, U3265, U4448);
  nand ginst8348 (U7692, U3264, U4403);
  nand ginst8349 (U7693, U3258, U3402);
  nand ginst8350 (U7694, U4465, U5481);
  nand ginst8351 (U7695, U7693, U7694);
  nand ginst8352 (U7696, INSTQUEUERD_ADDR_REG_3__SCAN_IN, U5464);
  nand ginst8353 (U7697, U4160, U5497);
  nand ginst8354 (U7698, INSTADDRPOINTER_REG_1__SCAN_IN, U4162);
  nand ginst8355 (U7699, INSTADDRPOINTER_REG_31__SCAN_IN, SUB_580_U6);
  not ginst8356 (U7700, U3457);
  nand ginst8357 (U7701, INSTADDRPOINTER_REG_0__SCAN_IN, U4162);
  nand ginst8358 (U7702, INSTADDRPOINTER_REG_0__SCAN_IN, INSTADDRPOINTER_REG_31__SCAN_IN);
  not ginst8359 (U7703, U3458);
  nand ginst8360 (U7704, U5489, U5499);
  nand ginst8361 (U7705, U3388, U4206);
  nand ginst8362 (U7706, INSTQUEUERD_ADDR_REG_1__SCAN_IN, U3251);
  nand ginst8363 (U7707, INSTQUEUERD_ADDR_REG_2__SCAN_IN, U3252);
  not ginst8364 (U7708, U3443);
  nand ginst8365 (U7709, INSTQUEUERD_ADDR_REG_2__SCAN_IN, U5464);
  nand ginst8366 (U7710, U4160, U5506);
  nand ginst8367 (U7711, INSTQUEUERD_ADDR_REG_1__SCAN_IN, U5464);
  nand ginst8368 (U7712, U4160, U5517);
  nand ginst8369 (U7713, INSTQUEUERD_ADDR_REG_0__SCAN_IN, U4202);
  nand ginst8370 (U7714, U3253, U5509);
  nand ginst8371 (U7715, INSTQUEUERD_ADDR_REG_0__SCAN_IN, U5464);
  nand ginst8372 (U7716, U4160, U5523);
  nand ginst8373 (U7717, INSTQUEUEWR_ADDR_REG_3__SCAN_IN, U5525);
  nand ginst8374 (U7718, U3391, U5533);
  nand ginst8375 (U7719, U4515, U7681);
  nand ginst8376 (U7720, U3301, U3441);
  nand ginst8377 (U7721, U7719, U7720);
  nand ginst8378 (U7722, INSTQUEUEWR_ADDR_REG_2__SCAN_IN, U5525);
  nand ginst8379 (U7723, U3391, U5537);
  nand ginst8380 (U7724, INSTQUEUEWR_ADDR_REG_1__SCAN_IN, U5525);
  nand ginst8381 (U7725, U3391, U5542);
  nand ginst8382 (U7726, INSTQUEUEWR_ADDR_REG_0__SCAN_IN, U5525);
  nand ginst8383 (U7727, U3391, U5545);
  nand ginst8384 (U7728, U3375, U4465);
  nand ginst8385 (U7729, U3258, U3268);
  nand ginst8386 (U7730, U3244, U4159, U7728, U7729);
  nand ginst8387 (U7731, R2167_U17, U4420, U7599);
  nand ginst8388 (U7732, EAX_REG_31__SCAN_IN, U3411);
  nand ginst8389 (U7733, U3466, U4211);
  nand ginst8390 (U7734, BYTEENABLE_REG_3__SCAN_IN, U3420);
  nand ginst8391 (U7735, U3467, U4208);
  or ginst8392 (U7736, DATAWIDTH_REG_0__SCAN_IN, DATAWIDTH_REG_1__SCAN_IN);
  nand ginst8393 (U7737, DATAWIDTH_REG_0__SCAN_IN, U3400);
  nand ginst8394 (U7738, U7736, U7737);
  nand ginst8395 (U7739, U3240, U7738);
  nand ginst8396 (U7740, REIP_REG_0__SCAN_IN, REIP_REG_1__SCAN_IN);
  nand ginst8397 (U7741, U7739, U7740);
  nand ginst8398 (U7742, BYTEENABLE_REG_2__SCAN_IN, U3420);
  nand ginst8399 (U7743, U4208, U7741);
  nand ginst8400 (U7744, BYTEENABLE_REG_1__SCAN_IN, U3420);
  nand ginst8401 (U7745, REIP_REG_1__SCAN_IN, U4208);
  nand ginst8402 (U7746, BYTEENABLE_REG_0__SCAN_IN, U3420);
  nand ginst8403 (U7747, U4208, U6587);
  nand ginst8404 (U7748, U3423, U4209);
  nand ginst8405 (U7749, W_R_N_REG_SCAN_IN, U3236);
  nand ginst8406 (U7750, MORE_REG_SCAN_IN, U4165);
  nand ginst8407 (U7751, U4225, U6588);
  nand ginst8408 (U7752, STATEBS16_REG_SCAN_IN, U7638);
  nand ginst8409 (U7753, BS16_N, U3449);
  nand ginst8410 (U7754, REQUESTPENDING_REG_SCAN_IN, U6591);
  nand ginst8411 (U7755, U4168, U6597);
  nand ginst8412 (U7756, U3422, U4209);
  nand ginst8413 (U7757, D_C_N_REG_SCAN_IN, U3236);
  nand ginst8414 (U7758, M_IO_N_REG_SCAN_IN, U3236);
  nand ginst8415 (U7759, MEMORYFETCH_REG_SCAN_IN, U4209);
  nand ginst8416 (U7760, READREQUEST_REG_SCAN_IN, U6602);
  nand ginst8417 (U7761, U4169, U6603);
  nand ginst8418 (U7762, U3475, U4170);
  nand ginst8419 (U7763, INSTQUEUERD_ADDR_REG_4__SCAN_IN, U5461);
  nand ginst8420 (U7764, INSTQUEUERD_ADDR_REG_3__SCAN_IN, U5461);
  nand ginst8421 (U7765, U4170, U5494);
  nand ginst8422 (U7766, INSTQUEUERD_ADDR_REG_2__SCAN_IN, U5461);
  nand ginst8423 (U7767, U4170, U5502);
  nand ginst8424 (U7768, INSTQUEUERD_ADDR_REG_1__SCAN_IN, U5461);
  nand ginst8425 (U7769, U4170, U5513);
  nand ginst8426 (U7770, INSTQUEUERD_ADDR_REG_0__SCAN_IN, U5461);
  nand ginst8427 (U7771, U4170, U5519);
  nand ginst8428 (U7772, U2605, U3264);
  nand ginst8429 (U7773, U4448, U7483);
  nand ginst8430 (U7774, U3288, U4191);
  nand ginst8431 (U7775, INSTQUEUEWR_ADDR_REG_0__SCAN_IN, U3284);
  nand ginst8432 (U7776, INSTQUEUERD_ADDR_REG_3__SCAN_IN, U4171);
  nand ginst8433 (U7777, U3257, U7207);
  not ginst8434 (U7778, U3444);
  nand ginst8435 (U7779, U3263, U3271);
  nand ginst8436 (U7780, U4482, U7695);
  nand ginst8437 (U7781, U3249, U3480);
  nand ginst8438 (U7782, FLUSH_REG_SCAN_IN, STATE2_REG_1__SCAN_IN, U7703);
  buf ginst8439 (W_R_N_REG_SCAN_IN_BUFF, W_R_N_REG_SCAN_IN);

endmodule

/*************** Perturb block ***************/
module Perturb (INSTQUEUE_REG_12__2__SCAN_IN, INSTQUEUE_REG_2__5__SCAN_IN, INSTQUEUE_REG_1__0__SCAN_IN, INSTQUEUE_REG_0__4__SCAN_IN, INSTADDRPOINTER_REG_21__SCAN_IN, INSTQUEUE_REG_9__5__SCAN_IN, INSTQUEUE_REG_1__1__SCAN_IN, INSTQUEUE_REG_2__1__SCAN_IN, INSTQUEUE_REG_12__0__SCAN_IN, INSTADDRPOINTER_REG_20__SCAN_IN, INSTQUEUEWR_ADDR_REG_1__SCAN_IN, INSTQUEUE_REG_10__0__SCAN_IN, INSTADDRPOINTER_REG_11__SCAN_IN, INSTADDRPOINTER_REG_2__SCAN_IN, INSTQUEUERD_ADDR_REG_1__SCAN_IN, INSTADDRPOINTER_REG_4__SCAN_IN, INSTQUEUE_REG_14__5__SCAN_IN, INSTQUEUE_REG_0__7__SCAN_IN, INSTQUEUE_REG_6__6__SCAN_IN, INSTQUEUE_REG_9__3__SCAN_IN, INSTQUEUE_REG_2__7__SCAN_IN, INSTQUEUE_REG_1__3__SCAN_IN, INSTQUEUE_REG_3__7__SCAN_IN, INSTQUEUE_REG_5__0__SCAN_IN, STATE2_REG_2__SCAN_IN, INSTQUEUE_REG_11__3__SCAN_IN, INSTQUEUE_REG_6__2__SCAN_IN, EBX_REG_5__SCAN_IN, INSTQUEUE_REG_12__5__SCAN_IN, INSTQUEUE_REG_5__7__SCAN_IN, INSTQUEUE_REG_12__7__SCAN_IN, INSTQUEUEWR_ADDR_REG_2__SCAN_IN, perturb_signal);

  input INSTQUEUE_REG_12__2__SCAN_IN, INSTQUEUE_REG_2__5__SCAN_IN, INSTQUEUE_REG_1__0__SCAN_IN, INSTQUEUE_REG_0__4__SCAN_IN, INSTADDRPOINTER_REG_21__SCAN_IN, INSTQUEUE_REG_9__5__SCAN_IN, INSTQUEUE_REG_1__1__SCAN_IN, INSTQUEUE_REG_2__1__SCAN_IN, INSTQUEUE_REG_12__0__SCAN_IN, INSTADDRPOINTER_REG_20__SCAN_IN, INSTQUEUEWR_ADDR_REG_1__SCAN_IN, INSTQUEUE_REG_10__0__SCAN_IN, INSTADDRPOINTER_REG_11__SCAN_IN, INSTADDRPOINTER_REG_2__SCAN_IN, INSTQUEUERD_ADDR_REG_1__SCAN_IN, INSTADDRPOINTER_REG_4__SCAN_IN, INSTQUEUE_REG_14__5__SCAN_IN, INSTQUEUE_REG_0__7__SCAN_IN, INSTQUEUE_REG_6__6__SCAN_IN, INSTQUEUE_REG_9__3__SCAN_IN, INSTQUEUE_REG_2__7__SCAN_IN, INSTQUEUE_REG_1__3__SCAN_IN, INSTQUEUE_REG_3__7__SCAN_IN, INSTQUEUE_REG_5__0__SCAN_IN, STATE2_REG_2__SCAN_IN, INSTQUEUE_REG_11__3__SCAN_IN, INSTQUEUE_REG_6__2__SCAN_IN, EBX_REG_5__SCAN_IN, INSTQUEUE_REG_12__5__SCAN_IN, INSTQUEUE_REG_5__7__SCAN_IN, INSTQUEUE_REG_12__7__SCAN_IN, INSTQUEUEWR_ADDR_REG_2__SCAN_IN;
  output perturb_signal;
  //SatHard key=10101101100011010101110000110110
  wire [31:0] sat_res_inputs;
  wire [31:0] keyvalue;
  assign sat_res_inputs[31:0] = {INSTQUEUE_REG_12__2__SCAN_IN, INSTQUEUE_REG_2__5__SCAN_IN, INSTQUEUE_REG_1__0__SCAN_IN, INSTQUEUE_REG_0__4__SCAN_IN, INSTADDRPOINTER_REG_21__SCAN_IN, INSTQUEUE_REG_9__5__SCAN_IN, INSTQUEUE_REG_1__1__SCAN_IN, INSTQUEUE_REG_2__1__SCAN_IN, INSTQUEUE_REG_12__0__SCAN_IN, INSTADDRPOINTER_REG_20__SCAN_IN, INSTQUEUEWR_ADDR_REG_1__SCAN_IN, INSTQUEUE_REG_10__0__SCAN_IN, INSTADDRPOINTER_REG_11__SCAN_IN, INSTADDRPOINTER_REG_2__SCAN_IN, INSTQUEUERD_ADDR_REG_1__SCAN_IN, INSTADDRPOINTER_REG_4__SCAN_IN, INSTQUEUE_REG_14__5__SCAN_IN, INSTQUEUE_REG_0__7__SCAN_IN, INSTQUEUE_REG_6__6__SCAN_IN, INSTQUEUE_REG_9__3__SCAN_IN, INSTQUEUE_REG_2__7__SCAN_IN, INSTQUEUE_REG_1__3__SCAN_IN, INSTQUEUE_REG_3__7__SCAN_IN, INSTQUEUE_REG_5__0__SCAN_IN, STATE2_REG_2__SCAN_IN, INSTQUEUE_REG_11__3__SCAN_IN, INSTQUEUE_REG_6__2__SCAN_IN, EBX_REG_5__SCAN_IN, INSTQUEUE_REG_12__5__SCAN_IN, INSTQUEUE_REG_5__7__SCAN_IN, INSTQUEUE_REG_12__7__SCAN_IN, INSTQUEUEWR_ADDR_REG_2__SCAN_IN};
  assign keyvalue[31:0] = 32'b10101101100011010101110000110110;

  integer ham_dist_peturb, idx;
  wire [31:0] diff;
  assign diff = sat_res_inputs ^ keyvalue;

  always@* begin
    ham_dist_peturb = 0;
    for(idx=0; idx<32; idx=idx+1) ham_dist_peturb = $signed($unsigned(ham_dist_peturb) + diff[idx]);
  end

  assign perturb_signal =  (ham_dist_peturb==4) ? 'b1 : 'b0;

endmodule
/*************** Perturb block ***************/

/*************** Restore block ***************/
module Restore (INSTQUEUE_REG_12__2__SCAN_IN, INSTQUEUE_REG_2__5__SCAN_IN, INSTQUEUE_REG_1__0__SCAN_IN, INSTQUEUE_REG_0__4__SCAN_IN, INSTADDRPOINTER_REG_21__SCAN_IN, INSTQUEUE_REG_9__5__SCAN_IN, INSTQUEUE_REG_1__1__SCAN_IN, INSTQUEUE_REG_2__1__SCAN_IN, INSTQUEUE_REG_12__0__SCAN_IN, INSTADDRPOINTER_REG_20__SCAN_IN, INSTQUEUEWR_ADDR_REG_1__SCAN_IN, INSTQUEUE_REG_10__0__SCAN_IN, INSTADDRPOINTER_REG_11__SCAN_IN, INSTADDRPOINTER_REG_2__SCAN_IN, INSTQUEUERD_ADDR_REG_1__SCAN_IN, INSTADDRPOINTER_REG_4__SCAN_IN, INSTQUEUE_REG_14__5__SCAN_IN, INSTQUEUE_REG_0__7__SCAN_IN, INSTQUEUE_REG_6__6__SCAN_IN, INSTQUEUE_REG_9__3__SCAN_IN, INSTQUEUE_REG_2__7__SCAN_IN, INSTQUEUE_REG_1__3__SCAN_IN, INSTQUEUE_REG_3__7__SCAN_IN, INSTQUEUE_REG_5__0__SCAN_IN, STATE2_REG_2__SCAN_IN, INSTQUEUE_REG_11__3__SCAN_IN, INSTQUEUE_REG_6__2__SCAN_IN, EBX_REG_5__SCAN_IN, INSTQUEUE_REG_12__5__SCAN_IN, INSTQUEUE_REG_5__7__SCAN_IN, INSTQUEUE_REG_12__7__SCAN_IN, INSTQUEUEWR_ADDR_REG_2__SCAN_IN, keyinput0, keyinput1, keyinput2, keyinput3, keyinput4, keyinput5, keyinput6, keyinput7, keyinput8, keyinput9, keyinput10, keyinput11, keyinput12, keyinput13, keyinput14, keyinput15, keyinput16, keyinput17, keyinput18, keyinput19, keyinput20, keyinput21, keyinput22, keyinput23, keyinput24, keyinput25, keyinput26, keyinput27, keyinput28, keyinput29, keyinput30, keyinput31, restore_signal);

  input INSTQUEUE_REG_12__2__SCAN_IN, INSTQUEUE_REG_2__5__SCAN_IN, INSTQUEUE_REG_1__0__SCAN_IN, INSTQUEUE_REG_0__4__SCAN_IN, INSTADDRPOINTER_REG_21__SCAN_IN, INSTQUEUE_REG_9__5__SCAN_IN, INSTQUEUE_REG_1__1__SCAN_IN, INSTQUEUE_REG_2__1__SCAN_IN, INSTQUEUE_REG_12__0__SCAN_IN, INSTADDRPOINTER_REG_20__SCAN_IN, INSTQUEUEWR_ADDR_REG_1__SCAN_IN, INSTQUEUE_REG_10__0__SCAN_IN, INSTADDRPOINTER_REG_11__SCAN_IN, INSTADDRPOINTER_REG_2__SCAN_IN, INSTQUEUERD_ADDR_REG_1__SCAN_IN, INSTADDRPOINTER_REG_4__SCAN_IN, INSTQUEUE_REG_14__5__SCAN_IN, INSTQUEUE_REG_0__7__SCAN_IN, INSTQUEUE_REG_6__6__SCAN_IN, INSTQUEUE_REG_9__3__SCAN_IN, INSTQUEUE_REG_2__7__SCAN_IN, INSTQUEUE_REG_1__3__SCAN_IN, INSTQUEUE_REG_3__7__SCAN_IN, INSTQUEUE_REG_5__0__SCAN_IN, STATE2_REG_2__SCAN_IN, INSTQUEUE_REG_11__3__SCAN_IN, INSTQUEUE_REG_6__2__SCAN_IN, EBX_REG_5__SCAN_IN, INSTQUEUE_REG_12__5__SCAN_IN, INSTQUEUE_REG_5__7__SCAN_IN, INSTQUEUE_REG_12__7__SCAN_IN, INSTQUEUEWR_ADDR_REG_2__SCAN_IN, keyinput0, keyinput1, keyinput2, keyinput3, keyinput4, keyinput5, keyinput6, keyinput7, keyinput8, keyinput9, keyinput10, keyinput11, keyinput12, keyinput13, keyinput14, keyinput15, keyinput16, keyinput17, keyinput18, keyinput19, keyinput20, keyinput21, keyinput22, keyinput23, keyinput24, keyinput25, keyinput26, keyinput27, keyinput28, keyinput29, keyinput30, keyinput31;
  output restore_signal;
  //SatHard key=10101101100011010101110000110110
  wire [31:0] sat_res_inputs;
  wire [31:0] keyinputs;
  assign sat_res_inputs[31:0] = {INSTQUEUE_REG_12__2__SCAN_IN, INSTQUEUE_REG_2__5__SCAN_IN, INSTQUEUE_REG_1__0__SCAN_IN, INSTQUEUE_REG_0__4__SCAN_IN, INSTADDRPOINTER_REG_21__SCAN_IN, INSTQUEUE_REG_9__5__SCAN_IN, INSTQUEUE_REG_1__1__SCAN_IN, INSTQUEUE_REG_2__1__SCAN_IN, INSTQUEUE_REG_12__0__SCAN_IN, INSTADDRPOINTER_REG_20__SCAN_IN, INSTQUEUEWR_ADDR_REG_1__SCAN_IN, INSTQUEUE_REG_10__0__SCAN_IN, INSTADDRPOINTER_REG_11__SCAN_IN, INSTADDRPOINTER_REG_2__SCAN_IN, INSTQUEUERD_ADDR_REG_1__SCAN_IN, INSTADDRPOINTER_REG_4__SCAN_IN, INSTQUEUE_REG_14__5__SCAN_IN, INSTQUEUE_REG_0__7__SCAN_IN, INSTQUEUE_REG_6__6__SCAN_IN, INSTQUEUE_REG_9__3__SCAN_IN, INSTQUEUE_REG_2__7__SCAN_IN, INSTQUEUE_REG_1__3__SCAN_IN, INSTQUEUE_REG_3__7__SCAN_IN, INSTQUEUE_REG_5__0__SCAN_IN, STATE2_REG_2__SCAN_IN, INSTQUEUE_REG_11__3__SCAN_IN, INSTQUEUE_REG_6__2__SCAN_IN, EBX_REG_5__SCAN_IN, INSTQUEUE_REG_12__5__SCAN_IN, INSTQUEUE_REG_5__7__SCAN_IN, INSTQUEUE_REG_12__7__SCAN_IN, INSTQUEUEWR_ADDR_REG_2__SCAN_IN};
  assign keyinputs[31:0] = {keyinput0, keyinput1, keyinput2, keyinput3, keyinput4, keyinput5, keyinput6, keyinput7, keyinput8, keyinput9, keyinput10, keyinput11, keyinput12, keyinput13, keyinput14, keyinput15, keyinput16, keyinput17, keyinput18, keyinput19, keyinput20, keyinput21, keyinput22, keyinput23, keyinput24, keyinput25, keyinput26, keyinput27, keyinput28, keyinput29, keyinput30, keyinput31};
  integer ham_dist_restore, idx;
  wire [31:0] diff;
  assign diff = sat_res_inputs ^ keyinputs;

  always@* begin
    ham_dist_restore = 0;
    for(idx=0; idx<32; idx=idx+1) ham_dist_restore = $signed($unsigned(ham_dist_restore) + diff[idx]);
  end

  assign restore_signal = (ham_dist_restore==4) ? 'b1 : 'b0;

endmodule
/*************** Restore block ***************/
