// Main module
module c3540(1, 13, 20, 33, 41, 45, 50, 58, 68, 77, 87, 97, 107, 116, 124, 125, 128, 132, 137, 143, 150, 159, 169, 179, 190, 200, 213, 222, 223, 226, 232, 238, 244, 250, 257, 264, 270, 274, 283, 294, 303, 311, 317, 322, 326, 329, 330, 343, 349, 350, 1713, 1947, 3195, 3833, 3987, 4028, 4145, 4589, 4667, 4815, 4944, 5002, 5045, 5047, 5078, 5102, 5120, 5121, 5192, 5231, 5360, 5361);

  input 1, 13, 20, 33, 41, 45, 50, 58, 68, 77, 87, 97, 107, 116, 124, 125, 128, 132, 137, 143, 150, 159, 169, 179, 190, 200, 213, 222, 223, 226, 232, 238, 244, 250, 257, 264, 270, 274, 283, 294, 303, 311, 317, 322, 326, 329, 330, 343, 349, 350;
  output 1713, 1947, 3195, 3833, 3987, 4028, 4145, 4589, 4667, 4815, 4944, 5002, 5045, 5047, 5078, 5102, 5120, 5121, 5192, 5231, 5360, 5361;
  wire 655, 665, 670, 679, 683, 686, 690, 699, 702, 706, 715, 724, 727, 736, 740, 749, 753, 763, 768, 769, 772, 779, 782, 786, 793, 794, 798, 803, 820, 821, 825, 829, 832, 835, 836, 839, 842, 845, 848, 851, 854, 858, 861, 864, 867, 870, 874, 877, 880, 883, 886, 889, 890, 891, 892, 895, 896, 913, 914, 915, 916, 917, 920, 923, 926, 929, 932, 935, 938, 941, 944, 947, 950, 953, 956, 959, 962, 965, 1067, 1117, 1179, 1196, 1197, 1202, 1219, 1250, 1251, 1252, 1253, 1254, 1255, 1256, 1257, 1258, 1259, 1260, 1261, 1262, 1263, 1264, 1267, 1268, 1271, 1272, 1273, 1276, 1279, 1298, 1302, 1306, 1315, 1322, 1325, 1328, 1331, 1334, 1337, 1338, 1339, 1340, 1343, 1344, 1345, 1346, 1347, 1348, 1349, 1350, 1351, 1352, 1353, 1358, 1363, 1366, 1369, 1384, 1401, 1402, 1403, 1404, 1405, 1406, 1407, 1408, 1409, 1426, 1427, 1452, 1459, 1460, 1461, 1464, 1467, 1468, 1469, 1470, 1471, 1474, 1475, 1478, 1481, 1484, 1487, 1490, 1493, 1496, 1499, 1502, 1505, 1507, 1508, 1509, 1510, 1511, 1512, 1520, 1562, 1579, 1580, 1581, 1582, 1583, 1584, 1585, 1586, 1587, 1588, 1589, 1590, 1591, 1592, 1593, 1594, 1595, 1596, 1597, 1598, 1599, 1600, 1643, 1644, 1645, 1646, 1647, 1648, 1649, 1650, 1667, 1670, 1673, 1674, 1675, 1676, 1677, 1678, 1679, 1680, 1691, 1692, 1693, 1694, 1714, 1715, 1718, 1721, 1722, 1725, 1726, 1727, 1728, 1729, 1730, 1731, 1735, 1736, 1737, 1738, 1747, 1756, 1761, 1764, 1765, 1766, 1767, 1768, 1769, 1770, 1787, 1788, 1789, 1790, 1791, 1792, 1793, 1794, 1795, 1796, 1797, 1798, 1799, 1800, 1801, 1802, 1803, 1806, 1809, 1812, 1815, 1818, 1821, 1824, 1833, 1842, 1843, 1844, 1845, 1846, 1847, 1848, 1849, 1850, 1851, 1852, 1853, 1854, 1855, 1856, 1857, 1858, 1859, 1860, 1861, 1862, 1863, 1864, 1869, 1870, 1873, 1874, 1875, 1878, 1879, 1880, 1883, 1884, 1885, 1888, 1889, 1890, 1893, 1894, 1895, 1898, 1899, 1900, 1903, 1904, 1905, 1908, 1909, 1912, 1913, 1917, 1922, 1926, 1930, 1933, 1936, 1939, 1940, 1941, 1942, 1943, 1944, 1945, 1946, 1960, 1961, 1966, 1981, 1982, 1983, 1986, 1987, 1988, 1989, 1990, 1991, 2022, 2023, 2024, 2025, 2026, 2027, 2028, 2029, 2030, 2031, 2032, 2033, 2034, 2035, 2036, 2037, 2038, 2043, 2052, 2057, 2068, 2073, 2078, 2083, 2088, 2093, 2098, 2103, 2121, 2122, 2123, 2124, 2125, 2126, 2127, 2128, 2133, 2134, 2135, 2136, 2137, 2138, 2139, 2141, 2142, 2143, 2144, 2145, 2146, 2147, 2148, 2149, 2150, 2151, 2152, 2153, 2154, 2155, 2156, 2157, 2158, 2175, 2178, 2179, 2180, 2181, 2183, 2184, 2185, 2188, 2191, 2194, 2197, 2200, 2203, 2206, 2209, 2210, 2211, 2212, 2221, 2230, 2231, 2232, 2233, 2234, 2235, 2236, 2237, 2238, 2239, 2240, 2241, 2242, 2243, 2244, 2245, 2270, 2277, 2282, 2287, 2294, 2299, 2304, 2307, 2310, 2313, 2316, 2319, 2322, 2325, 2328, 2331, 2334, 2341, 2342, 2347, 2348, 2349, 2350, 2351, 2352, 2353, 2354, 2355, 2374, 2375, 2376, 2379, 2398, 2417, 2418, 2419, 2420, 2421, 2422, 2425, 2426, 2427, 2430, 2431, 2432, 2435, 2436, 2437, 2438, 2439, 2440, 2443, 2444, 2445, 2448, 2449, 2450, 2467, 2468, 2469, 2470, 2471, 2474, 2475, 2476, 2477, 2478, 2481, 2482, 2483, 2486, 2487, 2488, 2497, 2506, 2515, 2524, 2533, 2542, 2551, 2560, 2569, 2578, 2587, 2596, 2605, 2614, 2623, 2632, 2633, 2634, 2635, 2636, 2637, 2638, 2639, 2640, 2641, 2642, 2643, 2644, 2645, 2646, 2647, 2648, 2652, 2656, 2659, 2662, 2666, 2670, 2673, 2677, 2681, 2684, 2688, 2692, 2697, 2702, 2706, 2710, 2715, 2719, 2723, 2728, 2729, 2730, 2731, 2732, 2733, 2734, 2735, 2736, 2737, 2738, 2739, 2740, 2741, 2742, 2743, 2744, 2745, 2746, 2748, 2749, 2750, 2751, 2754, 2755, 2756, 2757, 2758, 2761, 2764, 2768, 2769, 2898, 2899, 2900, 2901, 2962, 2966, 2967, 2970, 2973, 2977, 2980, 2984, 2985, 2986, 2987, 2988, 2989, 2990, 2991, 2992, 2993, 2994, 2995, 2996, 2997, 2998, 2999, 3000, 3001, 3002, 3003, 3004, 3005, 3006, 3007, 3008, 3009, 3010, 3011, 3012, 3013, 3014, 3015, 3016, 3017, 3018, 3019, 3020, 3021, 3022, 3023, 3024, 3025, 3026, 3027, 3028, 3029, 3030, 3031, 3032, 3033, 3034, 3035, 3036, 3037, 3038, 3039, 3040, 3041, 3042, 3043, 3044, 3045, 3046, 3047, 3048, 3049, 3050, 3051, 3052, 3053, 3054, 3055, 3056, 3057, 3058, 3059, 3060, 3061, 3062, 3063, 3064, 3065, 3066, 3067, 3068, 3069, 3070, 3071, 3072, 3073, 3074, 3075, 3076, 3077, 3078, 3079, 3080, 3081, 3082, 3083, 3084, 3085, 3086, 3087, 3088, 3089, 3090, 3091, 3092, 3093, 3094, 3095, 3096, 3097, 3098, 3099, 3100, 3101, 3102, 3103, 3104, 3105, 3106, 3107, 3108, 3109, 3110, 3111, 3112, 3115, 3118, 3119, 3122, 3125, 3128, 3131, 3134, 3135, 3138, 3141, 3142, 3145, 3148, 3149, 3152, 3155, 3158, 3161, 3164, 3165, 3168, 3171, 3172, 3175, 3178, 3181, 3184, 3187, 3190, 3191, 3192, 3193, 3194, 3196, 3206, 3207, 3208, 3209, 3210, 3211, 3212, 3213, 3214, 3215, 3216, 3217, 3218, 3219, 3220, 3221, 3222, 3223, 3224, 3225, 3226, 3227, 3228, 3229, 3230, 3231, 3232, 3233, 3234, 3235, 3236, 3237, 3238, 3239, 3240, 3241, 3242, 3243, 3244, 3245, 3246, 3247, 3248, 3249, 3250, 3251, 3252, 3253, 3254, 3255, 3256, 3257, 3258, 3259, 3260, 3261, 3262, 3263, 3264, 3265, 3266, 3267, 3268, 3269, 3270, 3271, 3272, 3273, 3274, 3275, 3276, 3277, 3278, 3279, 3280, 3281, 3282, 3283, 3284, 3285, 3286, 3287, 3288, 3289, 3290, 3291, 3292, 3293, 3294, 3295, 3296, 3297, 3298, 3299, 3300, 3301, 3302, 3303, 3304, 3305, 3306, 3307, 3308, 3309, 3310, 3311, 3312, 3313, 3314, 3315, 3316, 3317, 3318, 3319, 3320, 3321, 3322, 3323, 3324, 3325, 3326, 3327, 3328, 3329, 3330, 3331, 3332, 3333, 3334, 3383, 3384, 3387, 3388, 3389, 3390, 3391, 3392, 3393, 3394, 3395, 3396, 3397, 3398, 3399, 3400, 3401, 3402, 3403, 3404, 3405, 3406, 3407, 3410, 3413, 3414, 3415, 3419, 3423, 3426, 3429, 3430, 3431, 3434, 3437, 3438, 3439, 3442, 3445, 3446, 3447, 3451, 3455, 3458, 3461, 3462, 3463, 3466, 3469, 3470, 3471, 3472, 3475, 3478, 3481, 3484, 3487, 3490, 3493, 3496, 3499, 3502, 3505, 3508, 3511, 3514, 3517, 3520, 3523, 3534, 3535, 3536, 3537, 3538, 3539, 3540, 3541, 3542, 3543, 3544, 3545, 3546, 3547, 3548, 3549, 3550, 3551, 3552, 3557, 3568, 3573, 3578, 3589, 3594, 3605, 3626, 3627, 3628, 3629, 3630, 3631, 3632, 3633, 3634, 3635, 3636, 3637, 3638, 3639, 3640, 3641, 3642, 3643, 3644, 3645, 3648, 3651, 3652, 3653, 3654, 3657, 3658, 3661, 3662, 3663, 3664, 3667, 3670, 3671, 3672, 3673, 3676, 3677, 3680, 3681, 3682, 3685, 3686, 3687, 3688, 3689, 3690, 3693, 3694, 3695, 3696, 3697, 3700, 3703, 3704, 3705, 3706, 3707, 3708, 3711, 3712, 3713, 3714, 3715, 3716, 3717, 3718, 3719, 3720, 3721, 3731, 3734, 3740, 3743, 3753, 3756, 3762, 3765, 3766, 3773, 3774, 3775, 3776, 3777, 3778, 3779, 3780, 3786, 3789, 3800, 3803, 3809, 3812, 3815, 3818, 3821, 3824, 3827, 3830, 3834, 3835, 3838, 3845, 3850, 3855, 3858, 3861, 3865, 3868, 3884, 3885, 3894, 3895, 3898, 3899, 3906, 3911, 3912, 3913, 3916, 3917, 3920, 3921, 3924, 3925, 3926, 3930, 3931, 3932, 3935, 3936, 3937, 3940, 3947, 3948, 3950, 3953, 3956, 3959, 3962, 3965, 3968, 3971, 3974, 3977, 3980, 3983, 3992, 3996, 4013, 4029, 4030, 4031, 4032, 4033, 4034, 4035, 4042, 4043, 4044, 4045, 4046, 4047, 4048, 4049, 4050, 4051, 4052, 4053, 4054, 4055, 4056, 4057, 4058, 4059, 4062, 4065, 4066, 4067, 4070, 4073, 4074, 4075, 4076, 4077, 4078, 4079, 4080, 4085, 4086, 4088, 4090, 4091, 4094, 4098, 4101, 4104, 4105, 4106, 4107, 4108, 4109, 4110, 4111, 4112, 4113, 4114, 4115, 4116, 4119, 4122, 4123, 4126, 4127, 4128, 4139, 4142, 4146, 4147, 4148, 4149, 4150, 4151, 4152, 4153, 4154, 4161, 4167, 4174, 4182, 4186, 4189, 4190, 4191, 4192, 4193, 4194, 4195, 4196, 4197, 4200, 4203, 4209, 4213, 4218, 4223, 4238, 4239, 4241, 4242, 4247, 4251, 4252, 4253, 4254, 4255, 4256, 4257, 4258, 4283, 4284, 4287, 4291, 4295, 4296, 4299, 4303, 4304, 4305, 4310, 4316, 4317, 4318, 4319, 4322, 4325, 4326, 4327, 4328, 4329, 4330, 4331, 4335, 4338, 4341, 4344, 4347, 4350, 4353, 4356, 4359, 4362, 4365, 4368, 4371, 4376, 4377, 4387, 4390, 4393, 4398, 4413, 4416, 4421, 4427, 4430, 4435, 4442, 4443, 4446, 4447, 4448, 4452, 4458, 4461, 4462, 4463, 4464, 4465, 4468, 4472, 4475, 4479, 4484, 4486, 4487, 4491, 4493, 4496, 4497, 4498, 4503, 4506, 4507, 4508, 4509, 4510, 4511, 4515, 4526, 4527, 4528, 4529, 4530, 4531, 4534, 4537, 4540, 4545, 4549, 4552, 4555, 4558, 4559, 4562, 4563, 4564, 4568, 4569, 4572, 4573, 4576, 4581, 4584, 4587, 4588, 4593, 4596, 4597, 4599, 4602, 4603, 4608, 4613, 4616, 4619, 4623, 4628, 4629, 4630, 4635, 4636, 4640, 4641, 4642, 4643, 4644, 4647, 4650, 4656, 4659, 4664, 4668, 4669, 4670, 4673, 4674, 4675, 4676, 4677, 4678, 4679, 4687, 4688, 4691, 4694, 4697, 4700, 4704, 4705, 4706, 4707, 4708, 4711, 4716, 4717, 4721, 4722, 4726, 4727, 4730, 4733, 4740, 4743, 4747, 4748, 4749, 4750, 4753, 4754, 4755, 4756, 4757, 4769, 4772, 4775, 4778, 4786, 4787, 4788, 4789, 4794, 4797, 4800, 4805, 4808, 4812, 4816, 4817, 4818, 4822, 4823, 4826, 4829, 4830, 4831, 4838, 4844, 4847, 4850, 4854, 4859, 4860, 4868, 4870, 4872, 4873, 4876, 4880, 4885, 4889, 4895, 4896, 4897, 4898, 4899, 4900, 4901, 4902, 4904, 4905, 4906, 4907, 4913, 4916, 4920, 4921, 4924, 4925, 4926, 4928, 4929, 4930, 4931, 4937, 4940, 4946, 4949, 4950, 4951, 4952, 4953, 4954, 4957, 4964, 4965, 4968, 4969, 4970, 4973, 4978, 4979, 4980, 4981, 4982, 4983, 4984, 4985, 4988, 4991, 4996, 4999, 5007, 5010, 5013, 5018, 5021, 5026, 5029, 5030, 5039, 5042, 5046, 5050, 5055, 5058, 5061, 5066, 5070, 5080, 5085, 5094, 5095, 5097, 5103, 5108, 5109, 5110, 5111, 5114, 5117, 5122, 5125, 5128, 5133, 5136, 5139, 5145, 5151, 5154, 5159, 5160, 5163, 5166, 5173, 5174, 5177, 5182, 5183, 5184, 5188, 5193, 5196, 5197, 5198, 5199, 5201, 5203, 5205, 5209, 5212, 5215, 5217, 5219, 5220, 5221, 5222, 5223, 5224, 5225, 5228, 5232, 5233, 5234, 5235, 5236, 5240, 5242, 5243, 5245, 5246, 5250, 5253, 5254, 5257, 5258, 5261, 5266, 5269, 5277, 5278, 5279, 5283, 5284, 5285, 5286, 5289, 5292, 5295, 5298, 5303, 5306, 5309, 5312, 5313, 5322, 5323, 5324, 5327, 5332, 5335, 5340, 5341, 5344, 5345, 5348, 5349, 5350, 5351, 5352, 5353, 5354, 5355, 5356, 5357, 5358, 5359;

  and ginst1 (1067, 250, 768);
  or ginst2 (1117, 20, 820);
  or ginst3 (1179, 169, 895);
  not ginst4 (1196, 793);
  or ginst5 (1197, 1, 915);
  and ginst6 (1202, 913, 914);
  or ginst7 (1219, 1, 916);
  and ginst8 (1250, 842, 848, 854);
  nand ginst9 (1251, 226, 655);
  nand ginst10 (1252, 232, 670);
  nand ginst11 (1253, 238, 690);
  nand ginst12 (1254, 244, 706);
  nand ginst13 (1255, 250, 715);
  nand ginst14 (1256, 257, 727);
  nand ginst15 (1257, 264, 740);
  nand ginst16 (1258, 270, 753);
  not ginst17 (1259, 926);
  not ginst18 (1260, 929);
  not ginst19 (1261, 932);
  not ginst20 (1262, 935);
  nand ginst21 (1263, 679, 686);
  nand ginst22 (1264, 736, 749);
  nand ginst23 (1267, 683, 699);
  buf ginst24 (1268, 665);
  not ginst25 (1271, 953);
  not ginst26 (1272, 959);
  buf ginst27 (1273, 839);
  buf ginst28 (1276, 839);
  buf ginst29 (1279, 782);
  buf ginst30 (1298, 825);
  buf ginst31 (1302, 832);
  and ginst32 (1306, 779, 835);
  and ginst33 (1315, 779, 832, 836);
  and ginst34 (1322, 769, 836);
  and ginst35 (1325, 772, 786, 798);
  nand ginst36 (1328, 772, 786, 798);
  nand ginst37 (1331, 772, 786);
  buf ginst38 (1334, 874);
  nand ginst39 (1337, 45, 782, 794);
  nand ginst40 (1338, 842, 848, 854);
  not ginst41 (1339, 956);
  and ginst42 (1340, 861, 867, 870);
  nand ginst43 (1343, 861, 867, 870);
  not ginst44 (1344, 962);
  not ginst45 (1345, 803);
  not ginst46 (1346, 803);
  not ginst47 (1347, 803);
  not ginst48 (1348, 803);
  not ginst49 (1349, 803);
  not ginst50 (1350, 803);
  not ginst51 (1351, 803);
  not ginst52 (1352, 803);
  or ginst53 (1353, 883, 886);
  nor ginst54 (1358, 883, 886);
  buf ginst55 (1363, 892);
  not ginst56 (1366, 892);
  buf ginst57 (1369, 821);
  buf ginst58 (1384, 825);
  not ginst59 (1401, 896);
  not ginst60 (1402, 896);
  not ginst61 (1403, 896);
  not ginst62 (1404, 896);
  not ginst63 (1405, 896);
  not ginst64 (1406, 896);
  not ginst65 (1407, 896);
  not ginst66 (1408, 896);
  or ginst67 (1409, 1, 1196);
  not ginst68 (1426, 829);
  not ginst69 (1427, 829);
  and ginst70 (1452, 769, 782, 794);
  not ginst71 (1459, 917);
  not ginst72 (1460, 965);
  or ginst73 (1461, 920, 923);
  nor ginst74 (1464, 920, 923);
  not ginst75 (1467, 938);
  not ginst76 (1468, 941);
  not ginst77 (1469, 944);
  not ginst78 (1470, 947);
  buf ginst79 (1471, 679);
  not ginst80 (1474, 950);
  buf ginst81 (1475, 686);
  buf ginst82 (1478, 702);
  buf ginst83 (1481, 724);
  buf ginst84 (1484, 736);
  buf ginst85 (1487, 749);
  buf ginst86 (1490, 763);
  buf ginst87 (1493, 877);
  buf ginst88 (1496, 877);
  buf ginst89 (1499, 880);
  buf ginst90 (1502, 880);
  nand ginst91 (1505, 702, 1250);
  and ginst92 (1507, 1251, 1252, 1253, 1254);
  and ginst93 (1508, 1255, 1256, 1257, 1258);
  nand ginst94 (1509, 929, 1259);
  nand ginst95 (1510, 926, 1260);
  nand ginst96 (1511, 935, 1261);
  nand ginst97 (1512, 932, 1262);
  and ginst98 (1520, 655, 1263);
  and ginst99 (1562, 874, 1337);
  not ginst100 (1579, 1117);
  and ginst101 (1580, 803, 1117);
  and ginst102 (1581, 1338, 1345);
  not ginst103 (1582, 1117);
  and ginst104 (1583, 803, 1117);
  not ginst105 (1584, 1117);
  and ginst106 (1585, 803, 1117);
  and ginst107 (1586, 854, 1347);
  not ginst108 (1587, 1117);
  and ginst109 (1588, 803, 1117);
  and ginst110 (1589, 77, 1348);
  not ginst111 (1590, 1117);
  and ginst112 (1591, 803, 1117);
  and ginst113 (1592, 1343, 1349);
  not ginst114 (1593, 1117);
  and ginst115 (1594, 803, 1117);
  not ginst116 (1595, 1117);
  and ginst117 (1596, 803, 1117);
  and ginst118 (1597, 870, 1351);
  not ginst119 (1598, 1117);
  and ginst120 (1599, 803, 1117);
  and ginst121 (1600, 116, 1352);
  and ginst122 (1643, 222, 1401);
  and ginst123 (1644, 223, 1402);
  and ginst124 (1645, 226, 1403);
  and ginst125 (1646, 232, 1404);
  and ginst126 (1647, 238, 1405);
  and ginst127 (1648, 244, 1406);
  and ginst128 (1649, 250, 1407);
  and ginst129 (1650, 257, 1408);
  and ginst130 (1667, 1, 13, 1426);
  and ginst131 (1670, 1, 13, 1427);
  not ginst132 (1673, 1202);
  not ginst133 (1674, 1202);
  not ginst134 (1675, 1202);
  not ginst135 (1676, 1202);
  not ginst136 (1677, 1202);
  not ginst137 (1678, 1202);
  not ginst138 (1679, 1202);
  not ginst139 (1680, 1202);
  nand ginst140 (1691, 941, 1467);
  nand ginst141 (1692, 938, 1468);
  nand ginst142 (1693, 947, 1469);
  nand ginst143 (1694, 944, 1470);
  not ginst144 (1713, 1505);
  and ginst145 (1714, 87, 1264);
  nand ginst146 (1715, 1509, 1510);
  nand ginst147 (1718, 1511, 1512);
  nand ginst148 (1721, 1507, 1508);
  and ginst149 (1722, 763, 1340);
  nand ginst150 (1725, 763, 1340);
  not ginst151 (1726, 1268);
  nand ginst152 (1727, 1271, 1493);
  not ginst153 (1728, 1493);
  and ginst154 (1729, 683, 1268);
  nand ginst155 (1730, 1272, 1499);
  not ginst156 (1731, 1499);
  nand ginst157 (1735, 87, 1264);
  not ginst158 (1736, 1273);
  not ginst159 (1737, 1276);
  nand ginst160 (1738, 821, 1325);
  nand ginst161 (1747, 825, 1325);
  nand ginst162 (1756, 772, 798, 1279);
  nand ginst163 (1761, 772, 786, 798, 1302);
  nand ginst164 (1764, 1339, 1496);
  not ginst165 (1765, 1496);
  nand ginst166 (1766, 1344, 1502);
  not ginst167 (1767, 1502);
  not ginst168 (1768, 1328);
  not ginst169 (1769, 1334);
  not ginst170 (1770, 1331);
  and ginst171 (1787, 845, 1579);
  and ginst172 (1788, 150, 1580);
  and ginst173 (1789, 851, 1582);
  and ginst174 (1790, 159, 1583);
  and ginst175 (1791, 77, 1584);
  and ginst176 (1792, 50, 1585);
  and ginst177 (1793, 858, 1587);
  and ginst178 (1794, 845, 1588);
  and ginst179 (1795, 864, 1590);
  and ginst180 (1796, 851, 1591);
  and ginst181 (1797, 107, 1593);
  and ginst182 (1798, 77, 1594);
  and ginst183 (1799, 116, 1595);
  and ginst184 (1800, 858, 1596);
  and ginst185 (1801, 283, 1598);
  and ginst186 (1802, 864, 1599);
  and ginst187 (1803, 200, 1363);
  and ginst188 (1806, 889, 1363);
  and ginst189 (1809, 890, 1366);
  and ginst190 (1812, 891, 1366);
  nand ginst191 (1815, 1298, 1302);
  nand ginst192 (1818, 821, 1302);
  nand ginst193 (1821, 772, 1179, 1279);
  nand ginst194 (1824, 786, 794, 1298);
  nand ginst195 (1833, 786, 1298);
  not ginst196 (1842, 1369);
  not ginst197 (1843, 1369);
  not ginst198 (1844, 1369);
  not ginst199 (1845, 1369);
  not ginst200 (1846, 1369);
  not ginst201 (1847, 1369);
  not ginst202 (1848, 1369);
  not ginst203 (1849, 1384);
  and ginst204 (1850, 896, 1384);
  not ginst205 (1851, 1384);
  and ginst206 (1852, 896, 1384);
  not ginst207 (1853, 1384);
  and ginst208 (1854, 896, 1384);
  not ginst209 (1855, 1384);
  and ginst210 (1856, 896, 1384);
  not ginst211 (1857, 1384);
  and ginst212 (1858, 896, 1384);
  not ginst213 (1859, 1384);
  and ginst214 (1860, 896, 1384);
  not ginst215 (1861, 1384);
  and ginst216 (1862, 896, 1384);
  not ginst217 (1863, 1384);
  and ginst218 (1864, 896, 1384);
  and ginst219 (1869, 1202, 1409);
  nor ginst220 (1870, 50, 1409);
  not ginst221 (1873, 1306);
  and ginst222 (1874, 1202, 1409);
  nor ginst223 (1875, 58, 1409);
  not ginst224 (1878, 1306);
  and ginst225 (1879, 1202, 1409);
  nor ginst226 (1880, 68, 1409);
  not ginst227 (1883, 1306);
  and ginst228 (1884, 1202, 1409);
  nor ginst229 (1885, 77, 1409);
  not ginst230 (1888, 1306);
  and ginst231 (1889, 1202, 1409);
  nor ginst232 (1890, 87, 1409);
  not ginst233 (1893, 1322);
  and ginst234 (1894, 1202, 1409);
  nor ginst235 (1895, 97, 1409);
  not ginst236 (1898, 1315);
  and ginst237 (1899, 1202, 1409);
  nor ginst238 (1900, 107, 1409);
  not ginst239 (1903, 1315);
  and ginst240 (1904, 1202, 1409);
  nor ginst241 (1905, 116, 1409);
  not ginst242 (1908, 1315);
  and ginst243 (1909, 213, 1452);
  nand ginst244 (1912, 213, 1452);
  and ginst245 (1913, 213, 343, 1452);
  nand ginst246 (1917, 213, 343, 1452);
  and ginst247 (1922, 213, 343, 1452);
  nand ginst248 (1926, 213, 343, 1452);
  buf ginst249 (1930, 1464);
  nand ginst250 (1933, 1691, 1692);
  nand ginst251 (1936, 1693, 1694);
  not ginst252 (1939, 1471);
  nand ginst253 (1940, 1471, 1474);
  not ginst254 (1941, 1475);
  not ginst255 (1942, 1478);
  not ginst256 (1943, 1481);
  not ginst257 (1944, 1484);
  not ginst258 (1945, 1487);
  not ginst259 (1946, 1490);
  not ginst260 (1947, 1714);
  nand ginst261 (1960, 953, 1728);
  nand ginst262 (1961, 959, 1731);
  and ginst263 (1966, 1276, 1520);
  nand ginst264 (1981, 956, 1765);
  nand ginst265 (1982, 962, 1767);
  and ginst266 (1983, 1067, 1768);
  or ginst267 (1986, 1581, 1787, 1788);
  or ginst268 (1987, 1586, 1791, 1792);
  or ginst269 (1988, 1589, 1793, 1794);
  or ginst270 (1989, 1592, 1795, 1796);
  or ginst271 (1990, 1597, 1799, 1800);
  or ginst272 (1991, 1600, 1801, 1802);
  and ginst273 (2022, 77, 1849);
  and ginst274 (2023, 223, 1850);
  and ginst275 (2024, 87, 1851);
  and ginst276 (2025, 226, 1852);
  and ginst277 (2026, 97, 1853);
  and ginst278 (2027, 232, 1854);
  and ginst279 (2028, 107, 1855);
  and ginst280 (2029, 238, 1856);
  and ginst281 (2030, 116, 1857);
  and ginst282 (2031, 244, 1858);
  and ginst283 (2032, 283, 1859);
  and ginst284 (2033, 250, 1860);
  and ginst285 (2034, 294, 1861);
  and ginst286 (2035, 257, 1862);
  and ginst287 (2036, 303, 1863);
  and ginst288 (2037, 264, 1864);
  buf ginst289 (2038, 1667);
  not ginst290 (2043, 1667);
  buf ginst291 (2052, 1670);
  not ginst292 (2057, 1670);
  and ginst293 (2068, 50, 1197, 1869);
  and ginst294 (2073, 58, 1197, 1874);
  and ginst295 (2078, 68, 1197, 1879);
  and ginst296 (2083, 77, 1197, 1884);
  and ginst297 (2088, 87, 1219, 1889);
  and ginst298 (2093, 97, 1219, 1894);
  and ginst299 (2098, 107, 1219, 1899);
  and ginst300 (2103, 116, 1219, 1904);
  not ginst301 (2121, 1562);
  not ginst302 (2122, 1562);
  not ginst303 (2123, 1562);
  not ginst304 (2124, 1562);
  not ginst305 (2125, 1562);
  not ginst306 (2126, 1562);
  not ginst307 (2127, 1562);
  not ginst308 (2128, 1562);
  nand ginst309 (2133, 950, 1939);
  nand ginst310 (2134, 1478, 1941);
  nand ginst311 (2135, 1475, 1942);
  nand ginst312 (2136, 1484, 1943);
  nand ginst313 (2137, 1481, 1944);
  nand ginst314 (2138, 1490, 1945);
  nand ginst315 (2139, 1487, 1946);
  not ginst316 (2141, 1933);
  not ginst317 (2142, 1936);
  not ginst318 (2143, 1738);
  and ginst319 (2144, 1738, 1747);
  not ginst320 (2145, 1747);
  nand ginst321 (2146, 1727, 1960);
  nand ginst322 (2147, 1730, 1961);
  and ginst323 (2148, 58, 665, 1267, 1722);
  not ginst324 (2149, 1738);
  and ginst325 (2150, 1738, 1747);
  not ginst326 (2151, 1747);
  not ginst327 (2152, 1738);
  not ginst328 (2153, 1747);
  and ginst329 (2154, 1738, 1747);
  not ginst330 (2155, 1738);
  not ginst331 (2156, 1747);
  and ginst332 (2157, 1738, 1747);
  buf ginst333 (2158, 1761);
  buf ginst334 (2175, 1761);
  nand ginst335 (2178, 1764, 1981);
  nand ginst336 (2179, 1766, 1982);
  not ginst337 (2180, 1756);
  and ginst338 (2181, 1328, 1756);
  not ginst339 (2183, 1756);
  and ginst340 (2184, 1331, 1756);
  nand ginst341 (2185, 1358, 1812);
  nand ginst342 (2188, 1358, 1809);
  nand ginst343 (2191, 1353, 1812);
  nand ginst344 (2194, 1353, 1809);
  nand ginst345 (2197, 1358, 1806);
  nand ginst346 (2200, 1358, 1803);
  nand ginst347 (2203, 1353, 1806);
  nand ginst348 (2206, 1353, 1803);
  not ginst349 (2209, 1815);
  not ginst350 (2210, 1818);
  and ginst351 (2211, 1815, 1818);
  buf ginst352 (2212, 1821);
  buf ginst353 (2221, 1821);
  not ginst354 (2230, 1833);
  not ginst355 (2231, 1833);
  not ginst356 (2232, 1833);
  not ginst357 (2233, 1833);
  not ginst358 (2234, 1824);
  not ginst359 (2235, 1824);
  not ginst360 (2236, 1824);
  not ginst361 (2237, 1824);
  or ginst362 (2238, 1643, 2022, 2023);
  or ginst363 (2239, 1644, 2024, 2025);
  or ginst364 (2240, 1645, 2026, 2027);
  or ginst365 (2241, 1646, 2028, 2029);
  or ginst366 (2242, 1647, 2030, 2031);
  or ginst367 (2243, 1648, 2032, 2033);
  or ginst368 (2244, 1649, 2034, 2035);
  or ginst369 (2245, 1650, 2036, 2037);
  and ginst370 (2270, 1673, 1986);
  and ginst371 (2277, 1675, 1987);
  and ginst372 (2282, 1676, 1988);
  and ginst373 (2287, 1677, 1989);
  and ginst374 (2294, 1679, 1990);
  and ginst375 (2299, 1680, 1991);
  buf ginst376 (2304, 1917);
  and ginst377 (2307, 350, 1930);
  nand ginst378 (2310, 350, 1930);
  buf ginst379 (2313, 1715);
  buf ginst380 (2316, 1718);
  buf ginst381 (2319, 1715);
  buf ginst382 (2322, 1718);
  nand ginst383 (2325, 1940, 2133);
  nand ginst384 (2328, 2134, 2135);
  nand ginst385 (2331, 2136, 2137);
  nand ginst386 (2334, 2138, 2139);
  nand ginst387 (2341, 1936, 2141);
  nand ginst388 (2342, 1933, 2142);
  and ginst389 (2347, 724, 2144);
  and ginst390 (2348, 699, 1726, 2146);
  and ginst391 (2349, 753, 2147);
  and ginst392 (2350, 1273, 2148);
  and ginst393 (2351, 736, 2150);
  and ginst394 (2352, 1735, 2153);
  and ginst395 (2353, 763, 2154);
  and ginst396 (2354, 1725, 2156);
  and ginst397 (2355, 749, 2157);
  not ginst398 (2374, 2178);
  not ginst399 (2375, 2179);
  and ginst400 (2376, 1520, 2180);
  and ginst401 (2379, 1721, 2181);
  and ginst402 (2398, 665, 2211);
  and ginst403 (2417, 226, 1873, 2057);
  and ginst404 (2418, 274, 1306, 2057);
  and ginst405 (2419, 2052, 2238);
  and ginst406 (2420, 232, 1878, 2057);
  and ginst407 (2421, 274, 1306, 2057);
  and ginst408 (2422, 2052, 2239);
  and ginst409 (2425, 238, 1883, 2057);
  and ginst410 (2426, 274, 1306, 2057);
  and ginst411 (2427, 2052, 2240);
  and ginst412 (2430, 244, 1888, 2057);
  and ginst413 (2431, 274, 1306, 2057);
  and ginst414 (2432, 2052, 2241);
  and ginst415 (2435, 250, 1893, 2043);
  and ginst416 (2436, 274, 1322, 2043);
  and ginst417 (2437, 2038, 2242);
  and ginst418 (2438, 257, 1898, 2043);
  and ginst419 (2439, 274, 1315, 2043);
  and ginst420 (2440, 2038, 2243);
  and ginst421 (2443, 264, 1903, 2043);
  and ginst422 (2444, 274, 1315, 2043);
  and ginst423 (2445, 2038, 2244);
  and ginst424 (2448, 270, 1908, 2043);
  and ginst425 (2449, 274, 1315, 2043);
  and ginst426 (2450, 2038, 2245);
  not ginst427 (2467, 2313);
  not ginst428 (2468, 2316);
  not ginst429 (2469, 2319);
  not ginst430 (2470, 2322);
  nand ginst431 (2471, 2341, 2342);
  not ginst432 (2474, 2325);
  not ginst433 (2475, 2328);
  not ginst434 (2476, 2331);
  not ginst435 (2477, 2334);
  or ginst436 (2478, 1729, 2348);
  not ginst437 (2481, 2175);
  and ginst438 (2482, 1334, 2175);
  and ginst439 (2483, 2183, 2349);
  and ginst440 (2486, 1346, 2374);
  and ginst441 (2487, 1350, 2375);
  buf ginst442 (2488, 2185);
  buf ginst443 (2497, 2188);
  buf ginst444 (2506, 2191);
  buf ginst445 (2515, 2194);
  buf ginst446 (2524, 2197);
  buf ginst447 (2533, 2200);
  buf ginst448 (2542, 2203);
  buf ginst449 (2551, 2206);
  buf ginst450 (2560, 2185);
  buf ginst451 (2569, 2188);
  buf ginst452 (2578, 2191);
  buf ginst453 (2587, 2194);
  buf ginst454 (2596, 2197);
  buf ginst455 (2605, 2200);
  buf ginst456 (2614, 2203);
  buf ginst457 (2623, 2206);
  not ginst458 (2632, 2212);
  and ginst459 (2633, 1833, 2212);
  not ginst460 (2634, 2212);
  and ginst461 (2635, 1833, 2212);
  not ginst462 (2636, 2212);
  and ginst463 (2637, 1833, 2212);
  not ginst464 (2638, 2212);
  and ginst465 (2639, 1833, 2212);
  not ginst466 (2640, 2221);
  and ginst467 (2641, 1824, 2221);
  not ginst468 (2642, 2221);
  and ginst469 (2643, 1824, 2221);
  not ginst470 (2644, 2221);
  and ginst471 (2645, 1824, 2221);
  not ginst472 (2646, 2221);
  and ginst473 (2647, 1824, 2221);
  or ginst474 (2648, 1870, 2068, 2270);
  nor ginst475 (2652, 1870, 2068, 2270);
  or ginst476 (2656, 2417, 2418, 2419);
  or ginst477 (2659, 2420, 2421, 2422);
  or ginst478 (2662, 1880, 2078, 2277);
  nor ginst479 (2666, 1880, 2078, 2277);
  or ginst480 (2670, 2425, 2426, 2427);
  or ginst481 (2673, 1885, 2083, 2282);
  nor ginst482 (2677, 1885, 2083, 2282);
  or ginst483 (2681, 2430, 2431, 2432);
  or ginst484 (2684, 1890, 2088, 2287);
  nor ginst485 (2688, 1890, 2088, 2287);
  or ginst486 (2692, 2435, 2436, 2437);
  or ginst487 (2697, 2438, 2439, 2440);
  or ginst488 (2702, 1900, 2098, 2294);
  nor ginst489 (2706, 1900, 2098, 2294);
  or ginst490 (2710, 2443, 2444, 2445);
  or ginst491 (2715, 1905, 2103, 2299);
  nor ginst492 (2719, 1905, 2103, 2299);
  or ginst493 (2723, 2448, 2449, 2450);
  not ginst494 (2728, 2304);
  not ginst495 (2729, 2158);
  and ginst496 (2730, 1562, 2158);
  not ginst497 (2731, 2158);
  and ginst498 (2732, 1562, 2158);
  not ginst499 (2733, 2158);
  and ginst500 (2734, 1562, 2158);
  not ginst501 (2735, 2158);
  and ginst502 (2736, 1562, 2158);
  not ginst503 (2737, 2158);
  and ginst504 (2738, 1562, 2158);
  not ginst505 (2739, 2158);
  and ginst506 (2740, 1562, 2158);
  not ginst507 (2741, 2158);
  and ginst508 (2742, 1562, 2158);
  not ginst509 (2743, 2158);
  and ginst510 (2744, 1562, 2158);
  or ginst511 (2745, 1983, 2376, 2379);
  nor ginst512 (2746, 1983, 2376, 2379);
  nand ginst513 (2748, 2316, 2467);
  nand ginst514 (2749, 2313, 2468);
  nand ginst515 (2750, 2322, 2469);
  nand ginst516 (2751, 2319, 2470);
  nand ginst517 (2754, 2328, 2474);
  nand ginst518 (2755, 2325, 2475);
  nand ginst519 (2756, 2334, 2476);
  nand ginst520 (2757, 2331, 2477);
  and ginst521 (2758, 1520, 2481);
  and ginst522 (2761, 1722, 2482);
  and ginst523 (2764, 1770, 2478);
  or ginst524 (2768, 1789, 1790, 2486);
  or ginst525 (2769, 1797, 1798, 2487);
  and ginst526 (2898, 665, 2633);
  and ginst527 (2899, 679, 2635);
  and ginst528 (2900, 686, 2637);
  and ginst529 (2901, 702, 2639);
  not ginst530 (2962, 2746);
  nand ginst531 (2966, 2748, 2749);
  nand ginst532 (2967, 2750, 2751);
  buf ginst533 (2970, 2471);
  nand ginst534 (2973, 2754, 2755);
  nand ginst535 (2977, 2756, 2757);
  and ginst536 (2980, 2143, 2471);
  not ginst537 (2984, 2488);
  not ginst538 (2985, 2497);
  not ginst539 (2986, 2506);
  not ginst540 (2987, 2515);
  not ginst541 (2988, 2524);
  not ginst542 (2989, 2533);
  not ginst543 (2990, 2542);
  not ginst544 (2991, 2551);
  not ginst545 (2992, 2488);
  not ginst546 (2993, 2497);
  not ginst547 (2994, 2506);
  not ginst548 (2995, 2515);
  not ginst549 (2996, 2524);
  not ginst550 (2997, 2533);
  not ginst551 (2998, 2542);
  not ginst552 (2999, 2551);
  not ginst553 (3000, 2488);
  not ginst554 (3001, 2497);
  not ginst555 (3002, 2506);
  not ginst556 (3003, 2515);
  not ginst557 (3004, 2524);
  not ginst558 (3005, 2533);
  not ginst559 (3006, 2542);
  not ginst560 (3007, 2551);
  not ginst561 (3008, 2488);
  not ginst562 (3009, 2497);
  not ginst563 (3010, 2506);
  not ginst564 (3011, 2515);
  not ginst565 (3012, 2524);
  not ginst566 (3013, 2533);
  not ginst567 (3014, 2542);
  not ginst568 (3015, 2551);
  not ginst569 (3016, 2488);
  not ginst570 (3017, 2497);
  not ginst571 (3018, 2506);
  not ginst572 (3019, 2515);
  not ginst573 (3020, 2524);
  not ginst574 (3021, 2533);
  not ginst575 (3022, 2542);
  not ginst576 (3023, 2551);
  not ginst577 (3024, 2488);
  not ginst578 (3025, 2497);
  not ginst579 (3026, 2506);
  not ginst580 (3027, 2515);
  not ginst581 (3028, 2524);
  not ginst582 (3029, 2533);
  not ginst583 (3030, 2542);
  not ginst584 (3031, 2551);
  not ginst585 (3032, 2488);
  not ginst586 (3033, 2497);
  not ginst587 (3034, 2506);
  not ginst588 (3035, 2515);
  not ginst589 (3036, 2524);
  not ginst590 (3037, 2533);
  not ginst591 (3038, 2542);
  not ginst592 (3039, 2551);
  not ginst593 (3040, 2488);
  not ginst594 (3041, 2497);
  not ginst595 (3042, 2506);
  not ginst596 (3043, 2515);
  not ginst597 (3044, 2524);
  not ginst598 (3045, 2533);
  not ginst599 (3046, 2542);
  not ginst600 (3047, 2551);
  not ginst601 (3048, 2560);
  not ginst602 (3049, 2569);
  not ginst603 (3050, 2578);
  not ginst604 (3051, 2587);
  not ginst605 (3052, 2596);
  not ginst606 (3053, 2605);
  not ginst607 (3054, 2614);
  not ginst608 (3055, 2623);
  not ginst609 (3056, 2560);
  not ginst610 (3057, 2569);
  not ginst611 (3058, 2578);
  not ginst612 (3059, 2587);
  not ginst613 (3060, 2596);
  not ginst614 (3061, 2605);
  not ginst615 (3062, 2614);
  not ginst616 (3063, 2623);
  not ginst617 (3064, 2560);
  not ginst618 (3065, 2569);
  not ginst619 (3066, 2578);
  not ginst620 (3067, 2587);
  not ginst621 (3068, 2596);
  not ginst622 (3069, 2605);
  not ginst623 (3070, 2614);
  not ginst624 (3071, 2623);
  not ginst625 (3072, 2560);
  not ginst626 (3073, 2569);
  not ginst627 (3074, 2578);
  not ginst628 (3075, 2587);
  not ginst629 (3076, 2596);
  not ginst630 (3077, 2605);
  not ginst631 (3078, 2614);
  not ginst632 (3079, 2623);
  not ginst633 (3080, 2560);
  not ginst634 (3081, 2569);
  not ginst635 (3082, 2578);
  not ginst636 (3083, 2587);
  not ginst637 (3084, 2596);
  not ginst638 (3085, 2605);
  not ginst639 (3086, 2614);
  not ginst640 (3087, 2623);
  not ginst641 (3088, 2560);
  not ginst642 (3089, 2569);
  not ginst643 (3090, 2578);
  not ginst644 (3091, 2587);
  not ginst645 (3092, 2596);
  not ginst646 (3093, 2605);
  not ginst647 (3094, 2614);
  not ginst648 (3095, 2623);
  not ginst649 (3096, 2560);
  not ginst650 (3097, 2569);
  not ginst651 (3098, 2578);
  not ginst652 (3099, 2587);
  not ginst653 (3100, 2596);
  not ginst654 (3101, 2605);
  not ginst655 (3102, 2614);
  not ginst656 (3103, 2623);
  not ginst657 (3104, 2560);
  not ginst658 (3105, 2569);
  not ginst659 (3106, 2578);
  not ginst660 (3107, 2587);
  not ginst661 (3108, 2596);
  not ginst662 (3109, 2605);
  not ginst663 (3110, 2614);
  not ginst664 (3111, 2623);
  buf ginst665 (3112, 2656);
  not ginst666 (3115, 2656);
  not ginst667 (3118, 2652);
  and ginst668 (3119, 1674, 2768);
  buf ginst669 (3122, 2659);
  not ginst670 (3125, 2659);
  buf ginst671 (3128, 2670);
  not ginst672 (3131, 2670);
  not ginst673 (3134, 2666);
  buf ginst674 (3135, 2681);
  not ginst675 (3138, 2681);
  not ginst676 (3141, 2677);
  buf ginst677 (3142, 2692);
  not ginst678 (3145, 2692);
  not ginst679 (3148, 2688);
  and ginst680 (3149, 1678, 2769);
  buf ginst681 (3152, 2697);
  not ginst682 (3155, 2697);
  buf ginst683 (3158, 2710);
  not ginst684 (3161, 2710);
  not ginst685 (3164, 2706);
  buf ginst686 (3165, 2723);
  not ginst687 (3168, 2723);
  not ginst688 (3171, 2719);
  and ginst689 (3172, 1909, 2648);
  and ginst690 (3175, 1913, 2662);
  and ginst691 (3178, 1913, 2673);
  and ginst692 (3181, 1913, 2684);
  and ginst693 (3184, 1922, 2702);
  and ginst694 (3187, 1922, 2715);
  not ginst695 (3190, 2692);
  not ginst696 (3191, 2697);
  not ginst697 (3192, 2710);
  not ginst698 (3193, 2723);
  and ginst699 (3194, 1459, 2692, 2697, 2710, 2723);
  nand ginst700 (3195, 2745, 2962);
  not ginst701 (3196, 2966);
  or ginst702 (3206, 2145, 2347, 2980);
  and ginst703 (3207, 124, 2984);
  and ginst704 (3208, 159, 2985);
  and ginst705 (3209, 150, 2986);
  and ginst706 (3210, 143, 2987);
  and ginst707 (3211, 137, 2988);
  and ginst708 (3212, 132, 2989);
  and ginst709 (3213, 128, 2990);
  and ginst710 (3214, 125, 2991);
  and ginst711 (3215, 125, 2992);
  and ginst712 (3216, 655, 2993);
  and ginst713 (3217, 159, 2994);
  and ginst714 (3218, 150, 2995);
  and ginst715 (3219, 143, 2996);
  and ginst716 (3220, 137, 2997);
  and ginst717 (3221, 132, 2998);
  and ginst718 (3222, 128, 2999);
  and ginst719 (3223, 128, 3000);
  and ginst720 (3224, 670, 3001);
  and ginst721 (3225, 655, 3002);
  and ginst722 (3226, 159, 3003);
  and ginst723 (3227, 150, 3004);
  and ginst724 (3228, 143, 3005);
  and ginst725 (3229, 137, 3006);
  and ginst726 (3230, 132, 3007);
  and ginst727 (3231, 132, 3008);
  and ginst728 (3232, 690, 3009);
  and ginst729 (3233, 670, 3010);
  and ginst730 (3234, 655, 3011);
  and ginst731 (3235, 159, 3012);
  and ginst732 (3236, 150, 3013);
  and ginst733 (3237, 143, 3014);
  and ginst734 (3238, 137, 3015);
  and ginst735 (3239, 137, 3016);
  and ginst736 (3240, 706, 3017);
  and ginst737 (3241, 690, 3018);
  and ginst738 (3242, 670, 3019);
  and ginst739 (3243, 655, 3020);
  and ginst740 (3244, 159, 3021);
  and ginst741 (3245, 150, 3022);
  and ginst742 (3246, 143, 3023);
  and ginst743 (3247, 143, 3024);
  and ginst744 (3248, 715, 3025);
  and ginst745 (3249, 706, 3026);
  and ginst746 (3250, 690, 3027);
  and ginst747 (3251, 670, 3028);
  and ginst748 (3252, 655, 3029);
  and ginst749 (3253, 159, 3030);
  and ginst750 (3254, 150, 3031);
  and ginst751 (3255, 150, 3032);
  and ginst752 (3256, 727, 3033);
  and ginst753 (3257, 715, 3034);
  and ginst754 (3258, 706, 3035);
  and ginst755 (3259, 690, 3036);
  and ginst756 (3260, 670, 3037);
  and ginst757 (3261, 655, 3038);
  and ginst758 (3262, 159, 3039);
  and ginst759 (3263, 159, 3040);
  and ginst760 (3264, 740, 3041);
  and ginst761 (3265, 727, 3042);
  and ginst762 (3266, 715, 3043);
  and ginst763 (3267, 706, 3044);
  and ginst764 (3268, 690, 3045);
  and ginst765 (3269, 670, 3046);
  and ginst766 (3270, 655, 3047);
  and ginst767 (3271, 283, 3048);
  and ginst768 (3272, 670, 3049);
  and ginst769 (3273, 690, 3050);
  and ginst770 (3274, 706, 3051);
  and ginst771 (3275, 715, 3052);
  and ginst772 (3276, 727, 3053);
  and ginst773 (3277, 740, 3054);
  and ginst774 (3278, 753, 3055);
  and ginst775 (3279, 294, 3056);
  and ginst776 (3280, 690, 3057);
  and ginst777 (3281, 706, 3058);
  and ginst778 (3282, 715, 3059);
  and ginst779 (3283, 727, 3060);
  and ginst780 (3284, 740, 3061);
  and ginst781 (3285, 753, 3062);
  and ginst782 (3286, 283, 3063);
  and ginst783 (3287, 303, 3064);
  and ginst784 (3288, 706, 3065);
  and ginst785 (3289, 715, 3066);
  and ginst786 (3290, 727, 3067);
  and ginst787 (3291, 740, 3068);
  and ginst788 (3292, 753, 3069);
  and ginst789 (3293, 283, 3070);
  and ginst790 (3294, 294, 3071);
  and ginst791 (3295, 311, 3072);
  and ginst792 (3296, 715, 3073);
  and ginst793 (3297, 727, 3074);
  and ginst794 (3298, 740, 3075);
  and ginst795 (3299, 753, 3076);
  and ginst796 (3300, 283, 3077);
  and ginst797 (3301, 294, 3078);
  and ginst798 (3302, 303, 3079);
  and ginst799 (3303, 317, 3080);
  and ginst800 (3304, 727, 3081);
  and ginst801 (3305, 740, 3082);
  and ginst802 (3306, 753, 3083);
  and ginst803 (3307, 283, 3084);
  and ginst804 (3308, 294, 3085);
  and ginst805 (3309, 303, 3086);
  and ginst806 (3310, 311, 3087);
  and ginst807 (3311, 322, 3088);
  and ginst808 (3312, 740, 3089);
  and ginst809 (3313, 753, 3090);
  and ginst810 (3314, 283, 3091);
  and ginst811 (3315, 294, 3092);
  and ginst812 (3316, 303, 3093);
  and ginst813 (3317, 311, 3094);
  and ginst814 (3318, 317, 3095);
  and ginst815 (3319, 326, 3096);
  and ginst816 (3320, 753, 3097);
  and ginst817 (3321, 283, 3098);
  and ginst818 (3322, 294, 3099);
  and ginst819 (3323, 303, 3100);
  and ginst820 (3324, 311, 3101);
  and ginst821 (3325, 317, 3102);
  and ginst822 (3326, 322, 3103);
  and ginst823 (3327, 329, 3104);
  and ginst824 (3328, 283, 3105);
  and ginst825 (3329, 294, 3106);
  and ginst826 (3330, 303, 3107);
  and ginst827 (3331, 311, 3108);
  and ginst828 (3332, 317, 3109);
  and ginst829 (3333, 322, 3110);
  and ginst830 (3334, 326, 3111);
  and ginst831 (3383, 917, 3190, 3191, 3192, 3193);
  buf ginst832 (3384, 2977);
  and ginst833 (3387, 1736, 3196);
  and ginst834 (3388, 2149, 2977);
  and ginst835 (3389, 1737, 2973);
  nor ginst836 (3390, 3207, 3208, 3209, 3210, 3211, 3212, 3213, 3214);
  nor ginst837 (3391, 3215, 3216, 3217, 3218, 3219, 3220, 3221, 3222);
  nor ginst838 (3392, 3223, 3224, 3225, 3226, 3227, 3228, 3229, 3230);
  nor ginst839 (3393, 3231, 3232, 3233, 3234, 3235, 3236, 3237, 3238);
  nor ginst840 (3394, 3239, 3240, 3241, 3242, 3243, 3244, 3245, 3246);
  nor ginst841 (3395, 3247, 3248, 3249, 3250, 3251, 3252, 3253, 3254);
  nor ginst842 (3396, 3255, 3256, 3257, 3258, 3259, 3260, 3261, 3262);
  nor ginst843 (3397, 3263, 3264, 3265, 3266, 3267, 3268, 3269, 3270);
  nor ginst844 (3398, 3271, 3272, 3273, 3274, 3275, 3276, 3277, 3278);
  nor ginst845 (3399, 3279, 3280, 3281, 3282, 3283, 3284, 3285, 3286);
  nor ginst846 (3400, 3287, 3288, 3289, 3290, 3291, 3292, 3293, 3294);
  nor ginst847 (3401, 3295, 3296, 3297, 3298, 3299, 3300, 3301, 3302);
  nor ginst848 (3402, 3303, 3304, 3305, 3306, 3307, 3308, 3309, 3310);
  nor ginst849 (3403, 3311, 3312, 3313, 3314, 3315, 3316, 3317, 3318);
  nor ginst850 (3404, 3319, 3320, 3321, 3322, 3323, 3324, 3325, 3326);
  nor ginst851 (3405, 3327, 3328, 3329, 3330, 3331, 3332, 3333, 3334);
  and ginst852 (3406, 2641, 3206);
  and ginst853 (3407, 169, 2648, 3112);
  and ginst854 (3410, 179, 2648, 3115);
  and ginst855 (3413, 190, 2652, 3115);
  and ginst856 (3414, 200, 2652, 3112);
  or ginst857 (3415, 1875, 2073, 3119);
  nor ginst858 (3419, 1875, 2073, 3119);
  and ginst859 (3423, 169, 2662, 3128);
  and ginst860 (3426, 179, 2662, 3131);
  and ginst861 (3429, 190, 2666, 3131);
  and ginst862 (3430, 200, 2666, 3128);
  and ginst863 (3431, 169, 2673, 3135);
  and ginst864 (3434, 179, 2673, 3138);
  and ginst865 (3437, 190, 2677, 3138);
  and ginst866 (3438, 200, 2677, 3135);
  and ginst867 (3439, 169, 2684, 3142);
  and ginst868 (3442, 179, 2684, 3145);
  and ginst869 (3445, 190, 2688, 3145);
  and ginst870 (3446, 200, 2688, 3142);
  or ginst871 (3447, 1895, 2093, 3149);
  nor ginst872 (3451, 1895, 2093, 3149);
  and ginst873 (3455, 169, 2702, 3158);
  and ginst874 (3458, 179, 2702, 3161);
  and ginst875 (3461, 190, 2706, 3161);
  and ginst876 (3462, 200, 2706, 3158);
  and ginst877 (3463, 169, 2715, 3165);
  and ginst878 (3466, 179, 2715, 3168);
  and ginst879 (3469, 190, 2719, 3168);
  and ginst880 (3470, 200, 2719, 3165);
  or ginst881 (3471, 3194, 3383);
  buf ginst882 (3472, 2967);
  buf ginst883 (3475, 2970);
  buf ginst884 (3478, 2967);
  buf ginst885 (3481, 2970);
  buf ginst886 (3484, 2973);
  buf ginst887 (3487, 2973);
  buf ginst888 (3490, 3172);
  buf ginst889 (3493, 3172);
  buf ginst890 (3496, 3175);
  buf ginst891 (3499, 3175);
  buf ginst892 (3502, 3178);
  buf ginst893 (3505, 3178);
  buf ginst894 (3508, 3181);
  buf ginst895 (3511, 3181);
  buf ginst896 (3514, 3184);
  buf ginst897 (3517, 3184);
  buf ginst898 (3520, 3187);
  buf ginst899 (3523, 3187);
  nor ginst900 (3534, 2350, 3387);
  or ginst901 (3535, 2151, 2351, 3388);
  nor ginst902 (3536, 1966, 3389);
  and ginst903 (3537, 2209, 3390);
  and ginst904 (3538, 2210, 3398);
  and ginst905 (3539, 1842, 3391);
  and ginst906 (3540, 1369, 3399);
  and ginst907 (3541, 1843, 3392);
  and ginst908 (3542, 1369, 3400);
  and ginst909 (3543, 1844, 3393);
  and ginst910 (3544, 1369, 3401);
  and ginst911 (3545, 1845, 3394);
  and ginst912 (3546, 1369, 3402);
  and ginst913 (3547, 1846, 3395);
  and ginst914 (3548, 1369, 3403);
  and ginst915 (3549, 1847, 3396);
  and ginst916 (3550, 1369, 3404);
  and ginst917 (3551, 1848, 3397);
  and ginst918 (3552, 1369, 3405);
  or ginst919 (3557, 3118, 3413, 3414);
  or ginst920 (3568, 3134, 3429, 3430);
  or ginst921 (3573, 3141, 3437, 3438);
  or ginst922 (3578, 3148, 3445, 3446);
  or ginst923 (3589, 3164, 3461, 3462);
  or ginst924 (3594, 3171, 3469, 3470);
  and ginst925 (3605, 2728, 3471);
  not ginst926 (3626, 3478);
  not ginst927 (3627, 3481);
  not ginst928 (3628, 3487);
  not ginst929 (3629, 3484);
  not ginst930 (3630, 3472);
  not ginst931 (3631, 3475);
  and ginst932 (3632, 2152, 3536);
  and ginst933 (3633, 2155, 3534);
  or ginst934 (3634, 2398, 3537, 3538);
  or ginst935 (3635, 3539, 3540);
  or ginst936 (3636, 3541, 3542);
  or ginst937 (3637, 3543, 3544);
  or ginst938 (3638, 3545, 3546);
  or ginst939 (3639, 3547, 3548);
  or ginst940 (3640, 3549, 3550);
  or ginst941 (3641, 3551, 3552);
  and ginst942 (3642, 2643, 3535);
  or ginst943 (3643, 3407, 3410);
  nor ginst944 (3644, 3407, 3410);
  and ginst945 (3645, 169, 3122, 3415);
  and ginst946 (3648, 179, 3125, 3415);
  and ginst947 (3651, 190, 3125, 3419);
  and ginst948 (3652, 200, 3122, 3419);
  not ginst949 (3653, 3419);
  or ginst950 (3654, 3423, 3426);
  nor ginst951 (3657, 3423, 3426);
  or ginst952 (3658, 3431, 3434);
  nor ginst953 (3661, 3431, 3434);
  or ginst954 (3662, 3439, 3442);
  nor ginst955 (3663, 3439, 3442);
  and ginst956 (3664, 169, 3152, 3447);
  and ginst957 (3667, 179, 3155, 3447);
  and ginst958 (3670, 190, 3155, 3451);
  and ginst959 (3671, 200, 3152, 3451);
  not ginst960 (3672, 3451);
  or ginst961 (3673, 3455, 3458);
  nor ginst962 (3676, 3455, 3458);
  or ginst963 (3677, 3463, 3466);
  nor ginst964 (3680, 3463, 3466);
  not ginst965 (3681, 3493);
  and ginst966 (3682, 1909, 3415);
  not ginst967 (3685, 3496);
  not ginst968 (3686, 3499);
  not ginst969 (3687, 3502);
  not ginst970 (3688, 3505);
  not ginst971 (3689, 3511);
  and ginst972 (3690, 1922, 3447);
  not ginst973 (3693, 3517);
  not ginst974 (3694, 3520);
  not ginst975 (3695, 3523);
  not ginst976 (3696, 3514);
  buf ginst977 (3697, 3384);
  buf ginst978 (3700, 3384);
  not ginst979 (3703, 3490);
  not ginst980 (3704, 3508);
  nand ginst981 (3705, 3475, 3630);
  nand ginst982 (3706, 3472, 3631);
  nand ginst983 (3707, 3481, 3626);
  nand ginst984 (3708, 3478, 3627);
  or ginst985 (3711, 2352, 2353, 3632);
  or ginst986 (3712, 2354, 2355, 3633);
  and ginst987 (3713, 2632, 3634);
  and ginst988 (3714, 2634, 3635);
  and ginst989 (3715, 2636, 3636);
  and ginst990 (3716, 2638, 3637);
  and ginst991 (3717, 2640, 3638);
  and ginst992 (3718, 2642, 3639);
  and ginst993 (3719, 2644, 3640);
  and ginst994 (3720, 2646, 3641);
  and ginst995 (3721, 3557, 3644);
  or ginst996 (3731, 3651, 3652, 3653);
  and ginst997 (3734, 3568, 3657);
  and ginst998 (3740, 3573, 3661);
  and ginst999 (3743, 3578, 3663);
  or ginst1000 (3753, 3670, 3671, 3672);
  and ginst1001 (3756, 3589, 3676);
  and ginst1002 (3762, 3594, 3680);
  not ginst1003 (3765, 3643);
  not ginst1004 (3766, 3662);
  nand ginst1005 (3773, 3705, 3706);
  nand ginst1006 (3774, 3707, 3708);
  nand ginst1007 (3775, 3628, 3700);
  not ginst1008 (3776, 3700);
  nand ginst1009 (3777, 3629, 3697);
  not ginst1010 (3778, 3697);
  and ginst1011 (3779, 2645, 3712);
  and ginst1012 (3780, 2647, 3711);
  or ginst1013 (3786, 3645, 3648);
  nor ginst1014 (3789, 3645, 3648);
  or ginst1015 (3800, 3664, 3667);
  nor ginst1016 (3803, 3664, 3667);
  and ginst1017 (3809, 1917, 3654);
  and ginst1018 (3812, 1917, 3658);
  and ginst1019 (3815, 1926, 3673);
  and ginst1020 (3818, 1926, 3677);
  buf ginst1021 (3821, 3682);
  buf ginst1022 (3824, 3682);
  buf ginst1023 (3827, 3690);
  buf ginst1024 (3830, 3690);
  nand ginst1025 (3833, 3773, 3774);
  nand ginst1026 (3834, 3487, 3776);
  nand ginst1027 (3835, 3484, 3778);
  and ginst1028 (3838, 3731, 3789);
  and ginst1029 (3845, 3753, 3803);
  buf ginst1030 (3850, 3721);
  buf ginst1031 (3855, 3734);
  buf ginst1032 (3858, 3740);
  buf ginst1033 (3861, 3743);
  buf ginst1034 (3865, 3756);
  buf ginst1035 (3868, 3762);
  nand ginst1036 (3884, 3775, 3834);
  nand ginst1037 (3885, 3777, 3835);
  nand ginst1038 (3894, 3721, 3786);
  nand ginst1039 (3895, 3743, 3800);
  not ginst1040 (3898, 3821);
  not ginst1041 (3899, 3824);
  not ginst1042 (3906, 3830);
  not ginst1043 (3911, 3827);
  and ginst1044 (3912, 1912, 3786);
  buf ginst1045 (3913, 3812);
  and ginst1046 (3916, 1917, 3800);
  buf ginst1047 (3917, 3818);
  not ginst1048 (3920, 3809);
  buf ginst1049 (3921, 3818);
  not ginst1050 (3924, 3884);
  not ginst1051 (3925, 3885);
  and ginst1052 (3926, 3721, 3734, 3740, 3838);
  nand ginst1053 (3930, 3654, 3721, 3838);
  nand ginst1054 (3931, 3658, 3721, 3734, 3838);
  and ginst1055 (3932, 3743, 3756, 3762, 3845);
  nand ginst1056 (3935, 3673, 3743, 3845);
  nand ginst1057 (3936, 3677, 3743, 3756, 3845);
  buf ginst1058 (3937, 3838);
  buf ginst1059 (3940, 3845);
  not ginst1060 (3947, 3912);
  not ginst1061 (3948, 3916);
  buf ginst1062 (3950, 3850);
  buf ginst1063 (3953, 3850);
  buf ginst1064 (3956, 3855);
  buf ginst1065 (3959, 3855);
  buf ginst1066 (3962, 3858);
  buf ginst1067 (3965, 3858);
  buf ginst1068 (3968, 3861);
  buf ginst1069 (3971, 3861);
  buf ginst1070 (3974, 3865);
  buf ginst1071 (3977, 3865);
  buf ginst1072 (3980, 3868);
  buf ginst1073 (3983, 3868);
  nand ginst1074 (3987, 3924, 3925);
  nand ginst1075 (3992, 3765, 3894, 3930, 3931);
  nand ginst1076 (3996, 3766, 3895, 3935, 3936);
  not ginst1077 (4013, 3921);
  and ginst1078 (4028, 3926, 3932);
  nand ginst1079 (4029, 3681, 3953);
  nand ginst1080 (4030, 3686, 3959);
  nand ginst1081 (4031, 3688, 3965);
  nand ginst1082 (4032, 3689, 3971);
  nand ginst1083 (4033, 3693, 3977);
  nand ginst1084 (4034, 3695, 3983);
  buf ginst1085 (4035, 3926);
  not ginst1086 (4042, 3953);
  not ginst1087 (4043, 3956);
  nand ginst1088 (4044, 3685, 3956);
  not ginst1089 (4045, 3959);
  not ginst1090 (4046, 3962);
  nand ginst1091 (4047, 3687, 3962);
  not ginst1092 (4048, 3965);
  not ginst1093 (4049, 3971);
  not ginst1094 (4050, 3977);
  not ginst1095 (4051, 3980);
  nand ginst1096 (4052, 3694, 3980);
  not ginst1097 (4053, 3983);
  not ginst1098 (4054, 3974);
  nand ginst1099 (4055, 3696, 3974);
  and ginst1100 (4056, 2304, 3932);
  not ginst1101 (4057, 3950);
  nand ginst1102 (4058, 3703, 3950);
  buf ginst1103 (4059, 3937);
  buf ginst1104 (4062, 3937);
  not ginst1105 (4065, 3968);
  nand ginst1106 (4066, 3704, 3968);
  buf ginst1107 (4067, 3940);
  buf ginst1108 (4070, 3940);
  nand ginst1109 (4073, 3926, 3996);
  not ginst1110 (4074, 3992);
  nand ginst1111 (4075, 3493, 4042);
  nand ginst1112 (4076, 3499, 4045);
  nand ginst1113 (4077, 3505, 4048);
  nand ginst1114 (4078, 3511, 4049);
  nand ginst1115 (4079, 3517, 4050);
  nand ginst1116 (4080, 3523, 4053);
  nand ginst1117 (4085, 3496, 4043);
  nand ginst1118 (4086, 3502, 4046);
  nand ginst1119 (4088, 3520, 4051);
  nand ginst1120 (4090, 3514, 4054);
  and ginst1121 (4091, 1926, 3996);
  or ginst1122 (4094, 3605, 4056);
  nand ginst1123 (4098, 3490, 4057);
  nand ginst1124 (4101, 3508, 4065);
  and ginst1125 (4104, 4073, 4074);
  nand ginst1126 (4105, 4029, 4075);
  nand ginst1127 (4106, 3899, 4062);
  nand ginst1128 (4107, 4030, 4076);
  nand ginst1129 (4108, 4031, 4077);
  nand ginst1130 (4109, 4032, 4078);
  nand ginst1131 (4110, 3906, 4070);
  nand ginst1132 (4111, 4033, 4079);
  nand ginst1133 (4112, 4034, 4080);
  not ginst1134 (4113, 4059);
  nand ginst1135 (4114, 3898, 4059);
  not ginst1136 (4115, 4062);
  nand ginst1137 (4116, 4044, 4085);
  nand ginst1138 (4119, 4047, 4086);
  not ginst1139 (4122, 4070);
  nand ginst1140 (4123, 4052, 4088);
  not ginst1141 (4126, 4067);
  nand ginst1142 (4127, 3911, 4067);
  nand ginst1143 (4128, 4055, 4090);
  nand ginst1144 (4139, 4058, 4098);
  nand ginst1145 (4142, 4066, 4101);
  not ginst1146 (4145, 4104);
  not ginst1147 (4146, 4105);
  nand ginst1148 (4147, 3824, 4115);
  not ginst1149 (4148, 4107);
  not ginst1150 (4149, 4108);
  not ginst1151 (4150, 4109);
  nand ginst1152 (4151, 3830, 4122);
  not ginst1153 (4152, 4111);
  not ginst1154 (4153, 4112);
  nand ginst1155 (4154, 3821, 4113);
  nand ginst1156 (4161, 3827, 4126);
  buf ginst1157 (4167, 4091);
  buf ginst1158 (4174, 4094);
  buf ginst1159 (4182, 4091);
  and ginst1160 (4186, 330, 4094);
  and ginst1161 (4189, 2230, 4146);
  nand ginst1162 (4190, 4106, 4147);
  and ginst1163 (4191, 2232, 4148);
  and ginst1164 (4192, 2233, 4149);
  and ginst1165 (4193, 2234, 4150);
  nand ginst1166 (4194, 4110, 4151);
  and ginst1167 (4195, 2236, 4152);
  and ginst1168 (4196, 2237, 4153);
  nand ginst1169 (4197, 4114, 4154);
  buf ginst1170 (4200, 4116);
  buf ginst1171 (4203, 4116);
  buf ginst1172 (4209, 4119);
  buf ginst1173 (4213, 4119);
  nand ginst1174 (4218, 4127, 4161);
  buf ginst1175 (4223, 4123);
  and ginst1176 (4238, 3917, 4128);
  not ginst1177 (4239, 4139);
  not ginst1178 (4241, 4142);
  and ginst1179 (4242, 330, 4123);
  buf ginst1180 (4247, 4128);
  nor ginst1181 (4251, 2898, 3713, 4189);
  not ginst1182 (4252, 4190);
  nor ginst1183 (4253, 2900, 3715, 4191);
  nor ginst1184 (4254, 2901, 3716, 4192);
  nor ginst1185 (4255, 3406, 3717, 4193);
  not ginst1186 (4256, 4194);
  nor ginst1187 (4257, 3719, 3779, 4195);
  nor ginst1188 (4258, 3720, 3780, 4196);
  and ginst1189 (4283, 4035, 4167);
  and ginst1190 (4284, 4035, 4174);
  or ginst1191 (4287, 3815, 4238);
  not ginst1192 (4291, 4186);
  not ginst1193 (4295, 4167);
  buf ginst1194 (4296, 4167);
  not ginst1195 (4299, 4182);
  and ginst1196 (4303, 2231, 4252);
  and ginst1197 (4304, 2235, 4256);
  buf ginst1198 (4305, 4197);
  or ginst1199 (4310, 3992, 4283);
  and ginst1200 (4316, 4174, 4203, 4213);
  and ginst1201 (4317, 4174, 4209);
  and ginst1202 (4318, 4128, 4218, 4223);
  and ginst1203 (4319, 4128, 4223);
  and ginst1204 (4322, 4167, 4209);
  nand ginst1205 (4325, 3913, 4203);
  nand ginst1206 (4326, 4167, 4203, 4213);
  nand ginst1207 (4327, 3815, 4218);
  nand ginst1208 (4328, 3917, 4128, 4218);
  nand ginst1209 (4329, 4013, 4247);
  not ginst1210 (4330, 4247);
  and ginst1211 (4331, 330, 4094, 4295);
  and ginst1212 (4335, 2730, 4251);
  and ginst1213 (4338, 2734, 4253);
  and ginst1214 (4341, 2736, 4254);
  and ginst1215 (4344, 2738, 4255);
  and ginst1216 (4347, 2742, 4257);
  and ginst1217 (4350, 2744, 4258);
  buf ginst1218 (4353, 4197);
  buf ginst1219 (4356, 4203);
  buf ginst1220 (4359, 4209);
  buf ginst1221 (4362, 4218);
  buf ginst1222 (4365, 4242);
  buf ginst1223 (4368, 4242);
  and ginst1224 (4371, 4223, 4223);
  nor ginst1225 (4376, 2899, 3714, 4303);
  nor ginst1226 (4377, 3642, 3718, 4304);
  and ginst1227 (4387, 330, 4317);
  and ginst1228 (4390, 330, 4318);
  nand ginst1229 (4393, 3921, 4330);
  buf ginst1230 (4398, 4287);
  buf ginst1231 (4413, 4284);
  nand ginst1232 (4416, 3920, 4325, 4326);
  or ginst1233 (4421, 3812, 4322);
  nand ginst1234 (4427, 3948, 4327, 4328);
  buf ginst1235 (4430, 4287);
  and ginst1236 (4435, 330, 4316);
  or ginst1237 (4442, 4296, 4331);
  and ginst1238 (4443, 4174, 4203, 4213, 4305);
  nand ginst1239 (4446, 3809, 4305);
  nand ginst1240 (4447, 3913, 4200, 4305);
  nand ginst1241 (4448, 4167, 4200, 4213, 4305);
  not ginst1242 (4452, 4356);
  nand ginst1243 (4458, 4329, 4393);
  not ginst1244 (4461, 4365);
  not ginst1245 (4462, 4368);
  nand ginst1246 (4463, 1460, 4371);
  not ginst1247 (4464, 4371);
  buf ginst1248 (4465, 4310);
  nor ginst1249 (4468, 4296, 4331);
  and ginst1250 (4472, 2732, 4376);
  and ginst1251 (4475, 2740, 4377);
  buf ginst1252 (4479, 4310);
  not ginst1253 (4484, 4353);
  not ginst1254 (4486, 4359);
  nand ginst1255 (4487, 4299, 4359);
  not ginst1256 (4491, 4362);
  and ginst1257 (4493, 330, 4319);
  not ginst1258 (4496, 4398);
  and ginst1259 (4497, 4287, 4398);
  and ginst1260 (4498, 1769, 4442);
  nand ginst1261 (4503, 3947, 4446, 4447, 4448);
  not ginst1262 (4506, 4413);
  not ginst1263 (4507, 4435);
  not ginst1264 (4508, 4421);
  nand ginst1265 (4509, 4421, 4452);
  not ginst1266 (4510, 4427);
  nand ginst1267 (4511, 4241, 4427);
  nand ginst1268 (4515, 965, 4464);
  not ginst1269 (4526, 4416);
  nand ginst1270 (4527, 4416, 4484);
  nand ginst1271 (4528, 4182, 4486);
  not ginst1272 (4529, 4430);
  nand ginst1273 (4530, 4430, 4491);
  buf ginst1274 (4531, 4387);
  buf ginst1275 (4534, 4387);
  buf ginst1276 (4537, 4390);
  buf ginst1277 (4540, 4390);
  and ginst1278 (4545, 330, 4319, 4496);
  and ginst1279 (4549, 330, 4443);
  nand ginst1280 (4552, 4356, 4508);
  nand ginst1281 (4555, 4142, 4510);
  not ginst1282 (4558, 4493);
  nand ginst1283 (4559, 4463, 4515);
  not ginst1284 (4562, 4465);
  and ginst1285 (4563, 4310, 4465);
  buf ginst1286 (4564, 4468);
  not ginst1287 (4568, 4479);
  buf ginst1288 (4569, 4443);
  nand ginst1289 (4572, 4353, 4526);
  nand ginst1290 (4573, 4362, 4529);
  nand ginst1291 (4576, 4487, 4528);
  buf ginst1292 (4581, 4458);
  buf ginst1293 (4584, 4458);
  or ginst1294 (4587, 2758, 2761, 4498);
  nor ginst1295 (4588, 2758, 2761, 4498);
  or ginst1296 (4589, 4497, 4545);
  nand ginst1297 (4593, 4509, 4552);
  not ginst1298 (4596, 4531);
  not ginst1299 (4597, 4534);
  nand ginst1300 (4599, 4511, 4555);
  not ginst1301 (4602, 4537);
  not ginst1302 (4603, 4540);
  and ginst1303 (4608, 330, 4284, 4562);
  buf ginst1304 (4613, 4503);
  buf ginst1305 (4616, 4503);
  nand ginst1306 (4619, 4527, 4572);
  nand ginst1307 (4623, 4530, 4573);
  not ginst1308 (4628, 4588);
  nand ginst1309 (4629, 4506, 4569);
  not ginst1310 (4630, 4569);
  not ginst1311 (4635, 4576);
  nand ginst1312 (4636, 4291, 4576);
  not ginst1313 (4640, 4581);
  nand ginst1314 (4641, 4461, 4581);
  not ginst1315 (4642, 4584);
  nand ginst1316 (4643, 4462, 4584);
  nor ginst1317 (4644, 4563, 4608);
  and ginst1318 (4647, 2128, 4559);
  and ginst1319 (4650, 2743, 4559);
  buf ginst1320 (4656, 4549);
  buf ginst1321 (4659, 4549);
  buf ginst1322 (4664, 4564);
  and ginst1323 (4667, 4587, 4628);
  nand ginst1324 (4668, 4413, 4630);
  not ginst1325 (4669, 4616);
  nand ginst1326 (4670, 4239, 4616);
  not ginst1327 (4673, 4619);
  nand ginst1328 (4674, 4507, 4619);
  nand ginst1329 (4675, 4186, 4635);
  not ginst1330 (4676, 4623);
  nand ginst1331 (4677, 4558, 4623);
  nand ginst1332 (4678, 4365, 4640);
  nand ginst1333 (4679, 4368, 4642);
  not ginst1334 (4687, 4613);
  nand ginst1335 (4688, 4568, 4613);
  buf ginst1336 (4691, 4593);
  buf ginst1337 (4694, 4593);
  buf ginst1338 (4697, 4599);
  buf ginst1339 (4700, 4599);
  nand ginst1340 (4704, 4629, 4668);
  nand ginst1341 (4705, 4139, 4669);
  not ginst1342 (4706, 4656);
  not ginst1343 (4707, 4659);
  nand ginst1344 (4708, 4435, 4673);
  nand ginst1345 (4711, 4636, 4675);
  nand ginst1346 (4716, 4493, 4676);
  nand ginst1347 (4717, 4641, 4678);
  nand ginst1348 (4721, 4643, 4679);
  buf ginst1349 (4722, 4644);
  not ginst1350 (4726, 4664);
  or ginst1351 (4727, 4350, 4647, 4650);
  nor ginst1352 (4730, 4350, 4647, 4650);
  nand ginst1353 (4733, 4479, 4687);
  nand ginst1354 (4740, 4670, 4705);
  nand ginst1355 (4743, 4674, 4708);
  not ginst1356 (4747, 4691);
  nand ginst1357 (4748, 4596, 4691);
  not ginst1358 (4749, 4694);
  nand ginst1359 (4750, 4597, 4694);
  not ginst1360 (4753, 4697);
  nand ginst1361 (4754, 4602, 4697);
  not ginst1362 (4755, 4700);
  nand ginst1363 (4756, 4603, 4700);
  nand ginst1364 (4757, 4677, 4716);
  nand ginst1365 (4769, 4688, 4733);
  and ginst1366 (4772, 330, 4704);
  not ginst1367 (4775, 4721);
  not ginst1368 (4778, 4730);
  nand ginst1369 (4786, 4531, 4747);
  nand ginst1370 (4787, 4534, 4749);
  nand ginst1371 (4788, 4537, 4753);
  nand ginst1372 (4789, 4540, 4755);
  and ginst1373 (4794, 2124, 4711);
  and ginst1374 (4797, 2735, 4711);
  and ginst1375 (4800, 2127, 4717);
  buf ginst1376 (4805, 4722);
  and ginst1377 (4808, 4468, 4717);
  buf ginst1378 (4812, 4727);
  and ginst1379 (4815, 4727, 4778);
  not ginst1380 (4816, 4769);
  not ginst1381 (4817, 4772);
  nand ginst1382 (4818, 4748, 4786);
  nand ginst1383 (4822, 4750, 4787);
  nand ginst1384 (4823, 4754, 4788);
  nand ginst1385 (4826, 4756, 4789);
  nand ginst1386 (4829, 4726, 4775);
  not ginst1387 (4830, 4775);
  and ginst1388 (4831, 2122, 4743);
  and ginst1389 (4838, 2126, 4757);
  buf ginst1390 (4844, 4740);
  buf ginst1391 (4847, 4740);
  buf ginst1392 (4850, 4743);
  buf ginst1393 (4854, 4757);
  nand ginst1394 (4859, 4772, 4816);
  nand ginst1395 (4860, 4769, 4817);
  not ginst1396 (4868, 4826);
  not ginst1397 (4870, 4805);
  not ginst1398 (4872, 4808);
  nand ginst1399 (4873, 4664, 4830);
  or ginst1400 (4876, 4341, 4794, 4797);
  nor ginst1401 (4880, 4341, 4794, 4797);
  not ginst1402 (4885, 4812);
  not ginst1403 (4889, 4822);
  nand ginst1404 (4895, 4859, 4860);
  not ginst1405 (4896, 4844);
  nand ginst1406 (4897, 4706, 4844);
  not ginst1407 (4898, 4847);
  nand ginst1408 (4899, 4707, 4847);
  nor ginst1409 (4900, 4564, 4868);
  and ginst1410 (4901, 4564, 4717, 4757, 4823);
  not ginst1411 (4902, 4850);
  not ginst1412 (4904, 4854);
  nand ginst1413 (4905, 4854, 4872);
  nand ginst1414 (4906, 4829, 4873);
  and ginst1415 (4907, 2123, 4818);
  and ginst1416 (4913, 2125, 4823);
  and ginst1417 (4916, 4644, 4818);
  not ginst1418 (4920, 4880);
  and ginst1419 (4921, 2184, 4895);
  nand ginst1420 (4924, 4656, 4896);
  nand ginst1421 (4925, 4659, 4898);
  or ginst1422 (4926, 4900, 4901);
  nand ginst1423 (4928, 4870, 4889);
  not ginst1424 (4929, 4889);
  nand ginst1425 (4930, 4808, 4904);
  not ginst1426 (4931, 4906);
  buf ginst1427 (4937, 4876);
  buf ginst1428 (4940, 4876);
  and ginst1429 (4944, 4876, 4920);
  nand ginst1430 (4946, 4897, 4924);
  nand ginst1431 (4949, 4899, 4925);
  nand ginst1432 (4950, 4902, 4916);
  not ginst1433 (4951, 4916);
  nand ginst1434 (4952, 4805, 4929);
  nand ginst1435 (4953, 4905, 4930);
  and ginst1436 (4954, 2737, 4926);
  and ginst1437 (4957, 2741, 4931);
  or ginst1438 (4964, 2483, 2764, 4921);
  nor ginst1439 (4965, 2483, 2764, 4921);
  not ginst1440 (4968, 4949);
  nand ginst1441 (4969, 4850, 4951);
  nand ginst1442 (4970, 4928, 4952);
  and ginst1443 (4973, 2739, 4953);
  not ginst1444 (4978, 4937);
  not ginst1445 (4979, 4940);
  not ginst1446 (4980, 4965);
  nor ginst1447 (4981, 4722, 4968);
  and ginst1448 (4982, 4722, 4743, 4818, 4946);
  nand ginst1449 (4983, 4950, 4969);
  not ginst1450 (4984, 4970);
  and ginst1451 (4985, 2121, 4946);
  or ginst1452 (4988, 4344, 4913, 4954);
  nor ginst1453 (4991, 4344, 4913, 4954);
  or ginst1454 (4996, 4347, 4800, 4957);
  nor ginst1455 (4999, 4347, 4800, 4957);
  and ginst1456 (5002, 4964, 4980);
  or ginst1457 (5007, 4981, 4982);
  and ginst1458 (5010, 2731, 4983);
  and ginst1459 (5013, 2733, 4984);
  or ginst1460 (5018, 4475, 4838, 4973);
  nor ginst1461 (5021, 4475, 4838, 4973);
  not ginst1462 (5026, 4991);
  not ginst1463 (5029, 4999);
  and ginst1464 (5030, 2729, 5007);
  buf ginst1465 (5039, 4996);
  buf ginst1466 (5042, 4988);
  and ginst1467 (5045, 4988, 5026);
  not ginst1468 (5046, 5021);
  and ginst1469 (5047, 4996, 5029);
  or ginst1470 (5050, 4472, 4831, 5010);
  nor ginst1471 (5055, 4472, 4831, 5010);
  or ginst1472 (5058, 4338, 4907, 5013);
  nor ginst1473 (5061, 4338, 4907, 5013);
  and ginst1474 (5066, 4730, 4991, 4999, 5021);
  buf ginst1475 (5070, 5018);
  and ginst1476 (5078, 5018, 5046);
  or ginst1477 (5080, 4335, 4985, 5030);
  nor ginst1478 (5085, 4335, 4985, 5030);
  nand ginst1479 (5094, 4885, 5039);
  not ginst1480 (5095, 5039);
  not ginst1481 (5097, 5042);
  and ginst1482 (5102, 5050, 5050);
  not ginst1483 (5103, 5061);
  nand ginst1484 (5108, 4812, 5095);
  not ginst1485 (5109, 5070);
  nand ginst1486 (5110, 5070, 5097);
  buf ginst1487 (5111, 5058);
  and ginst1488 (5114, 1461, 5050);
  buf ginst1489 (5117, 5050);
  and ginst1490 (5120, 5080, 5080);
  and ginst1491 (5121, 5058, 5103);
  nand ginst1492 (5122, 5094, 5108);
  nand ginst1493 (5125, 5042, 5109);
  and ginst1494 (5128, 1461, 5080);
  and ginst1495 (5133, 4880, 5055, 5061, 5085);
  and ginst1496 (5136, 1464, 5055, 5085);
  buf ginst1497 (5139, 5080);
  nand ginst1498 (5145, 5110, 5125);
  buf ginst1499 (5151, 5111);
  buf ginst1500 (5154, 5111);
  not ginst1501 (5159, 5117);
  buf ginst1502 (5160, 5114);
  buf ginst1503 (5163, 5114);
  and ginst1504 (5166, 5066, 5133);
  and ginst1505 (5173, 5066, 5133);
  buf ginst1506 (5174, 5122);
  buf ginst1507 (5177, 5122);
  not ginst1508 (5182, 5139);
  nand ginst1509 (5183, 5139, 5159);
  buf ginst1510 (5184, 5128);
  buf ginst1511 (5188, 5128);
  not ginst1512 (5192, 5166);
  nor ginst1513 (5193, 5136, 5173);
  nand ginst1514 (5196, 4978, 5151);
  not ginst1515 (5197, 5151);
  nand ginst1516 (5198, 4979, 5154);
  not ginst1517 (5199, 5154);
  not ginst1518 (5201, 5160);
  not ginst1519 (5203, 5163);
  buf ginst1520 (5205, 5145);
  buf ginst1521 (5209, 5145);
  nand ginst1522 (5212, 5117, 5182);
  and ginst1523 (5215, 213, 5193);
  not ginst1524 (5217, 5174);
  not ginst1525 (5219, 5177);
  nand ginst1526 (5220, 4937, 5197);
  nand ginst1527 (5221, 4940, 5199);
  not ginst1528 (5222, 5184);
  nand ginst1529 (5223, 5184, 5201);
  nand ginst1530 (5224, 5188, 5203);
  not ginst1531 (5225, 5188);
  nand ginst1532 (5228, 5183, 5212);
  not ginst1533 (5231, 5215);
  nand ginst1534 (5232, 5205, 5217);
  not ginst1535 (5233, 5205);
  nand ginst1536 (5234, 5209, 5219);
  not ginst1537 (5235, 5209);
  nand ginst1538 (5236, 5196, 5220);
  nand ginst1539 (5240, 5198, 5221);
  nand ginst1540 (5242, 5160, 5222);
  nand ginst1541 (5243, 5163, 5225);
  nand ginst1542 (5245, 5174, 5233);
  nand ginst1543 (5246, 5177, 5235);
  not ginst1544 (5250, 5240);
  not ginst1545 (5253, 5228);
  nand ginst1546 (5254, 5223, 5242);
  nand ginst1547 (5257, 5224, 5243);
  nand ginst1548 (5258, 5232, 5245);
  nand ginst1549 (5261, 5234, 5246);
  not ginst1550 (5266, 5257);
  buf ginst1551 (5269, 5236);
  and ginst1552 (5277, 2307, 5236, 5254);
  and ginst1553 (5278, 2310, 5250, 5254);
  not ginst1554 (5279, 5261);
  not ginst1555 (5283, 5269);
  nand ginst1556 (5284, 5253, 5269);
  and ginst1557 (5285, 2310, 5236, 5266);
  and ginst1558 (5286, 2307, 5250, 5266);
  buf ginst1559 (5289, 5258);
  buf ginst1560 (5292, 5258);
  nand ginst1561 (5295, 5228, 5283);
  or ginst1562 (5298, 5277, 5278, 5285, 5286);
  buf ginst1563 (5303, 5279);
  buf ginst1564 (5306, 5279);
  nand ginst1565 (5309, 5284, 5295);
  not ginst1566 (5312, 5292);
  not ginst1567 (5313, 5289);
  not ginst1568 (5322, 5306);
  not ginst1569 (5323, 5303);
  buf ginst1570 (5324, 5298);
  buf ginst1571 (5327, 5298);
  buf ginst1572 (5332, 5309);
  buf ginst1573 (5335, 5309);
  nand ginst1574 (5340, 5323, 5324);
  nand ginst1575 (5341, 5322, 5327);
  not ginst1576 (5344, 5327);
  not ginst1577 (5345, 5324);
  nand ginst1578 (5348, 5313, 5332);
  nand ginst1579 (5349, 5312, 5335);
  nand ginst1580 (5350, 5303, 5345);
  nand ginst1581 (5351, 5306, 5344);
  not ginst1582 (5352, 5335);
  not ginst1583 (5353, 5332);
  nand ginst1584 (5354, 5289, 5353);
  nand ginst1585 (5355, 5292, 5352);
  nand ginst1586 (5356, 5340, 5350);
  nand ginst1587 (5357, 5341, 5351);
  nand ginst1588 (5358, 5348, 5354);
  nand ginst1589 (5359, 5349, 5355);
  and ginst1590 (5360, 5356, 5357);
  nand ginst1591 (5361, 5358, 5359);
  buf ginst1592 (655, 50);
  not ginst1593 (665, 50);
  buf ginst1594 (670, 58);
  not ginst1595 (679, 58);
  buf ginst1596 (683, 68);
  not ginst1597 (686, 68);
  buf ginst1598 (690, 68);
  buf ginst1599 (699, 77);
  not ginst1600 (702, 77);
  buf ginst1601 (706, 77);
  buf ginst1602 (715, 87);
  not ginst1603 (724, 87);
  buf ginst1604 (727, 97);
  not ginst1605 (736, 97);
  buf ginst1606 (740, 107);
  not ginst1607 (749, 107);
  buf ginst1608 (753, 116);
  not ginst1609 (763, 116);
  or ginst1610 (768, 257, 264);
  not ginst1611 (769, 1);
  buf ginst1612 (772, 1);
  not ginst1613 (779, 1);
  buf ginst1614 (782, 13);
  not ginst1615 (786, 13);
  and ginst1616 (793, 13, 20);
  not ginst1617 (794, 20);
  buf ginst1618 (798, 20);
  not ginst1619 (803, 20);
  not ginst1620 (820, 33);
  buf ginst1621 (821, 33);
  not ginst1622 (825, 33);
  and ginst1623 (829, 33, 41);
  not ginst1624 (832, 41);
  or ginst1625 (835, 41, 45);
  buf ginst1626 (836, 45);
  not ginst1627 (839, 45);
  not ginst1628 (842, 50);
  buf ginst1629 (845, 58);
  not ginst1630 (848, 58);
  buf ginst1631 (851, 68);
  not ginst1632 (854, 68);
  buf ginst1633 (858, 87);
  not ginst1634 (861, 87);
  buf ginst1635 (864, 97);
  not ginst1636 (867, 97);
  not ginst1637 (870, 107);
  buf ginst1638 (874, 1);
  buf ginst1639 (877, 68);
  buf ginst1640 (880, 107);
  not ginst1641 (883, 20);
  buf ginst1642 (886, 190);
  not ginst1643 (889, 200);
  and ginst1644 (890, 20, 200);
  nand ginst1645 (891, 20, 200);
  and ginst1646 (892, 20, 179);
  not ginst1647 (895, 20);
  or ginst1648 (896, 33, 349);
  nand ginst1649 (913, 1, 13);
  nand ginst1650 (914, 1, 20, 33);
  not ginst1651 (915, 20);
  not ginst1652 (916, 33);
  buf ginst1653 (917, 179);
  not ginst1654 (920, 213);
  buf ginst1655 (923, 343);
  buf ginst1656 (926, 226);
  buf ginst1657 (929, 232);
  buf ginst1658 (932, 238);
  buf ginst1659 (935, 244);
  buf ginst1660 (938, 250);
  buf ginst1661 (941, 257);
  buf ginst1662 (944, 264);
  buf ginst1663 (947, 270);
  buf ginst1664 (950, 50);
  buf ginst1665 (953, 58);
  buf ginst1666 (956, 58);
  buf ginst1667 (959, 97);
  buf ginst1668 (962, 97);
  buf ginst1669 (965, 330);

endmodule
