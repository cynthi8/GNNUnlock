//key=01101100100010100011000101110110
// Main module
module c2670_SFLL-HD(0)_32_1(i_1, i_2, i_3, i_4, i_5, i_6, i_7, i_8, i_11, i_14, i_15, i_16, i_19, i_20, i_21, i_22, i_23, i_24, i_25, i_26, i_27, i_28, i_29, i_32, i_33, i_34, i_35, i_36, i_37, i_40, i_43, i_44, i_47, i_48, i_49, i_50, i_51, i_52, i_53, i_54, i_55, i_56, i_57, i_60, i_61, i_62, i_63, i_64, i_65, i_66, i_67, i_68, i_69, i_72, i_73, i_74, i_75, i_76, i_77, i_78, i_79, i_80, i_81, i_82, i_85, i_86, i_87, i_88, i_89, i_90, i_91, i_92, i_93, i_94, i_95, i_96, i_99, i_100, i_101, i_102, i_103, i_104, i_105, i_106, i_107, i_108, i_111, i_112, i_113, i_114, i_115, i_116, i_117, i_118, i_119, i_120, i_123, i_124, i_125, i_126, i_127, i_128, i_129, i_130, i_131, i_132, i_135, i_136, i_137, i_138, i_139, i_140, i_141, i_142, i_143, i_144, i_145, i_146, i_147, i_148, i_149, i_150, i_151, i_152, i_153, i_154, i_155, i_156, i_157, i_158, i_159, i_160, i_161, i_162, i_163, i_164, i_165, i_166, i_167, i_168, i_169, i_170, i_171, i_172, i_173, i_174, i_175, i_176, i_177, i_178, i_179, i_180, i_181, i_182, i_183, i_184, i_185, i_186, i_187, i_188, i_189, i_190, i_191, i_192, i_193, i_194, i_195, i_196, i_197, i_198, i_199, i_200, i_201, i_202, i_203, i_204, i_205, i_206, i_207, i_208, i_209, i_210, i_211, i_212, i_213, i_214, i_215, i_216, i_217, i_218, i_219, i_224, i_227, i_230, i_231, i_234, i_237, i_241, i_246, i_253, i_256, i_259, i_262, i_263, i_266, i_269, i_272, i_275, i_278, i_281, i_284, i_287, i_290, i_294, i_297, i_301, i_305, i_309, i_313, i_316, i_319, i_322, i_325, i_328, i_331, i_334, i_337, i_340, i_343, i_346, i_349, i_352, i_355, keyinput0, keyinput1, keyinput2, keyinput3, keyinput4, keyinput5, keyinput6, keyinput7, keyinput8, keyinput9, keyinput10, keyinput11, keyinput12, keyinput13, keyinput14, keyinput15, keyinput16, keyinput17, keyinput18, keyinput19, keyinput20, keyinput21, keyinput22, keyinput23, keyinput24, keyinput25, keyinput26, keyinput27, keyinput28, keyinput29, keyinput30, keyinput31, i_143, i_144, i_145, i_146, i_147, i_148, i_149, i_150, i_151, i_152, i_153, i_154, i_155, i_156, i_157, i_158, i_159, i_160, i_161, i_162, i_163, i_164, i_165, i_166, i_167, i_168, i_169, i_170, i_171, i_172, i_173, i_174, i_175, i_176, i_177, i_178, i_179, i_180, i_181, i_182, i_183, i_184, i_185, i_186, i_187, i_188, i_189, i_190, i_191, i_192, i_193, i_194, i_195, i_196, i_197, i_198, i_199, i_200, i_201, i_202, i_203, i_204, i_205, i_206, i_207, i_208, i_209, i_210, i_211, i_212, i_213, i_214, i_215, i_216, i_217, i_218, i_398, i_400, i_401, i_419, i_420, i_456, i_457, i_458, i_487, i_488, i_489, i_490, i_491, i_492, i_493, i_494, i_792, i_799, i_805, i_1026, i_1028, i_1029, i_1269, i_1277, i_1448, i_1726, i_1816, i_1817, i_1818, i_1819, i_1820, i_1821, i_1969, i_1970, i_1971, i_2010, i_2012, i_2014, i_2016, i_2018, i_2020, i_2022, i_2387, i_2388, i_2389, i_2390, i_2496, i_2643, i_2644, i_2891, i_2925, i_2970, i_2971, i_3038, i_3079, i_3546, i_3671, i_3803, i_3804, i_3809, i_3851, i_3875, i_3881, i_3882);

  input i_1, i_2, i_3, i_4, i_5, i_6, i_7, i_8, i_11, i_14, i_15, i_16, i_19, i_20, i_21, i_22, i_23, i_24, i_25, i_26, i_27, i_28, i_29, i_32, i_33, i_34, i_35, i_36, i_37, i_40, i_43, i_44, i_47, i_48, i_49, i_50, i_51, i_52, i_53, i_54, i_55, i_56, i_57, i_60, i_61, i_62, i_63, i_64, i_65, i_66, i_67, i_68, i_69, i_72, i_73, i_74, i_75, i_76, i_77, i_78, i_79, i_80, i_81, i_82, i_85, i_86, i_87, i_88, i_89, i_90, i_91, i_92, i_93, i_94, i_95, i_96, i_99, i_100, i_101, i_102, i_103, i_104, i_105, i_106, i_107, i_108, i_111, i_112, i_113, i_114, i_115, i_116, i_117, i_118, i_119, i_120, i_123, i_124, i_125, i_126, i_127, i_128, i_129, i_130, i_131, i_132, i_135, i_136, i_137, i_138, i_139, i_140, i_141, i_142, i_143, i_144, i_145, i_146, i_147, i_148, i_149, i_150, i_151, i_152, i_153, i_154, i_155, i_156, i_157, i_158, i_159, i_160, i_161, i_162, i_163, i_164, i_165, i_166, i_167, i_168, i_169, i_170, i_171, i_172, i_173, i_174, i_175, i_176, i_177, i_178, i_179, i_180, i_181, i_182, i_183, i_184, i_185, i_186, i_187, i_188, i_189, i_190, i_191, i_192, i_193, i_194, i_195, i_196, i_197, i_198, i_199, i_200, i_201, i_202, i_203, i_204, i_205, i_206, i_207, i_208, i_209, i_210, i_211, i_212, i_213, i_214, i_215, i_216, i_217, i_218, i_219, i_224, i_227, i_230, i_231, i_234, i_237, i_241, i_246, i_253, i_256, i_259, i_262, i_263, i_266, i_269, i_272, i_275, i_278, i_281, i_284, i_287, i_290, i_294, i_297, i_301, i_305, i_309, i_313, i_316, i_319, i_322, i_325, i_328, i_331, i_334, i_337, i_340, i_343, i_346, i_349, i_352, i_355, keyinput0, keyinput1, keyinput2, keyinput3, keyinput4, keyinput5, keyinput6, keyinput7, keyinput8, keyinput9, keyinput10, keyinput11, keyinput12, keyinput13, keyinput14, keyinput15, keyinput16, keyinput17, keyinput18, keyinput19, keyinput20, keyinput21, keyinput22, keyinput23, keyinput24, keyinput25, keyinput26, keyinput27, keyinput28, keyinput29, keyinput30, keyinput31;
  output i_143, i_144, i_145, i_146, i_147, i_148, i_149, i_150, i_151, i_152, i_153, i_154, i_155, i_156, i_157, i_158, i_159, i_160, i_161, i_162, i_163, i_164, i_165, i_166, i_167, i_168, i_169, i_170, i_171, i_172, i_173, i_174, i_175, i_176, i_177, i_178, i_179, i_180, i_181, i_182, i_183, i_184, i_185, i_186, i_187, i_188, i_189, i_190, i_191, i_192, i_193, i_194, i_195, i_196, i_197, i_198, i_199, i_200, i_201, i_202, i_203, i_204, i_205, i_206, i_207, i_208, i_209, i_210, i_211, i_212, i_213, i_214, i_215, i_216, i_217, i_218, i_398, i_400, i_401, i_419, i_420, i_456, i_457, i_458, i_487, i_488, i_489, i_490, i_491, i_492, i_493, i_494, i_792, i_799, i_805, i_1026, i_1028, i_1029, i_1269, i_1277, i_1448, i_1726, i_1816, i_1817, i_1818, i_1819, i_1820, i_1821, i_1969, i_1970, i_1971, i_2010, i_2012, i_2014, i_2016, i_2018, i_2020, i_2022, i_2387, i_2388, i_2389, i_2390, i_2496, i_2643, i_2644, i_2891, i_2925, i_2970, i_2971, i_3038, i_3079, i_3546, i_3671, i_3803, i_3804, i_3809, i_3851, i_3875, i_3881, i_3882;
  wire i_1027, i_1032, i_1033, i_1034, i_1037, i_1042, i_1053, i_1064, i_1065, i_1066, i_1067, i_1068, i_1069, i_1070, i_1075, i_1086, i_1097, i_1098, i_1099, i_1100, i_1101, i_1102, i_1113, i_1124, i_1125, i_1126, i_1127, i_1128, i_1129, i_1133, i_1137, i_1140, i_1141, i_1142, i_1143, i_1144, i_1145, i_1146, i_1157, i_1168, i_1169, i_1170, i_1171, i_1172, i_1173, i_1178, i_1184, i_1185, i_1186, i_1187, i_1188, i_1189, i_1190, i_1195, i_1200, i_1205, i_1210, i_1211, i_1212, i_1213, i_1214, i_1215, i_1216, i_1219, i_1222, i_1225, i_1228, i_1231, i_1234, i_1237, i_1240, i_1243, i_1246, i_1249, i_1250, i_1251, i_1254, i_1257, i_1260, i_1263, i_1266, i_1275, i_1276, i_1302, i_1351, i_1352, i_1353, i_1354, i_1355, i_1395, i_1396, i_1397, i_1398, i_1399, i_1422, i_1423, i_1424, i_1425, i_1426, i_1427, i_1440, i_1441, i_1449, i_1450, i_1451, i_1452, i_1453, i_1454, i_1455, i_1456, i_1457, i_1458, i_1459, i_1460, i_1461, i_1462, i_1463, i_1464, i_1465, i_1466, i_1467, i_1468, i_1469, i_1470, i_1471, i_1472, i_1473, i_1474, i_1475, i_1476, i_1477, i_1478, i_1479, i_1480, i_1481, i_1482, i_1483, i_1484, i_1485, i_1486, i_1487, i_1488, i_1489, i_1490, i_1491, i_1492, i_1493, i_1494, i_1495, i_1496, i_1499, i_1502, i_1506, i_1510, i_1513, i_1516, i_1519, i_1520, i_1521, i_1522, i_1523, i_1524, i_1525, i_1526, i_1527, i_1528, i_1529, i_1530, i_1531, i_1532, i_1533, i_1534, i_1535, i_1536, i_1537, i_1538, i_1539, i_1540, i_1541, i_1542, i_1543, i_1544, i_1545, i_1546, i_1547, i_1548, i_1549, i_1550, i_1551, i_1552, i_1553, i_1557, i_1561, i_1564, i_1565, i_1566, i_1567, i_1568, i_1569, i_1570, i_1571, i_1572, i_1573, i_1574, i_1575, i_1576, i_1577, i_1578, i_1581, i_1582, i_1585, i_1588, i_1591, i_1596, i_1600, i_1606, i_1612, i_1615, i_1619, i_1624, i_1628, i_1631, i_1634, i_1637, i_1642, i_1647, i_1651, i_1656, i_1676, i_1681, i_1686, i_1690, i_1708, i_1770, i_1773, i_1776, i_1777, i_1778, i_1781, i_1784, i_1785, i_1795, i_1798, i_1801, i_1804, i_1807, i_1808, i_1809, i_1810, i_1811, i_1813, i_1814, i_1815, i_1822, i_1823, i_1824, i_1827, i_1830, i_1831, i_1832, i_1833, i_1836, i_1841, i_1848, i_1852, i_1856, i_1863, i_1870, i_1875, i_1880, i_1885, i_1888, i_1891, i_1894, i_1897, i_1908, i_1909, i_1910, i_1911, i_1912, i_1913, i_1914, i_1915, i_1916, i_1917, i_1918, i_1919, i_1928, i_1929, i_1930, i_1931, i_1932, i_1933, i_1934, i_1935, i_1936, i_1939, i_1940, i_1941, i_1942, i_1945, i_1948, i_1951, i_1954, i_1957, i_1960, i_1963, i_1966, i_2028, i_2029, i_2030, i_2031, i_2032, i_2033, i_2034, i_2040, i_2041, i_2042, i_2043, i_2046, i_2049, i_2052, i_2055, i_2058, i_2061, i_2064, i_2067, i_2070, i_2073, i_2076, i_2079, i_2095, i_2098, i_2101, i_2104, i_2107, i_2110, i_2113, i_2119, i_2120, i_2125, i_2126, i_2127, i_2128, i_2135, i_2141, i_2144, i_2147, i_2150, i_2153, i_2154, i_2155, i_2156, i_2157, i_2158, i_2171, i_2172, i_2173, i_2174, i_2175, i_2176, i_2177, i_2178, i_2185, i_2188, i_2191, i_2194, i_2197, i_2200, i_2201, i_2204, i_2207, i_2210, i_2213, i_2216, i_2219, i_2234, i_2235, i_2236, i_2237, i_2250, i_2266, i_2269, i_2291, i_2294, i_2297, i_2298, i_2300, i_2301, i_2302, i_2303, i_2304, i_2305, i_2306, i_2307, i_2308, i_2309, i_2310, i_2311, i_2312, i_2313, i_2314, i_2315, i_2316, i_2317, i_2318, i_2319, i_2320, i_2321, i_2322, i_2323, i_2324, i_2325, i_2326, i_2327, i_2328, i_2329, i_2330, i_2331, i_2332, i_2333, i_2334, i_2335, i_2336, i_2337, i_2338, i_2339, i_2340, i_2354, i_2355, i_2356, i_2357, i_2358, i_2359, i_2364, i_2365, i_2366, i_2367, i_2368, i_2372, i_2373, i_2374, i_2375, i_2376, i_2377, i_2382, i_2386, i_2391, i_2395, i_2400, i_2403, i_2406, i_2407, i_2408, i_2409, i_2410, i_2411, i_2412, i_2413, i_2414, i_2415, i_2416, i_2417, i_2421, i_2425, i_2428, i_2429, i_2430, i_2431, i_2432, i_2433, i_2434, i_2437, i_2440, i_2443, i_2446, i_2449, i_2452, i_2453, i_2454, i_2457, i_2460, i_2463, i_2466, i_2469, i_2472, i_2475, i_2478, i_2481, i_2484, i_2487, i_2490, i_2493, i_2503, i_2504, i_2510, i_2511, i_2521, i_2528, i_2531, i_2534, i_2537, i_2540, i_2544, i_2545, i_2546, i_2547, i_2548, i_2549, i_2550, i_2551, i_2552, i_2553, i_2563, i_2564, i_2565, i_2566, i_2567, i_2568, i_2579, i_2603, i_2607, i_2608, i_2609, i_2610, i_2611, i_2612, i_2613, i_2617, i_2618, i_2619, i_2620, i_2621, i_2624, i_2628, i_2629, i_2630, i_2631, i_2632, i_2633, i_2634, i_2635, i_2636, i_2638, i_2645, i_2646, i_2652, i_2655, i_2656, i_2659, i_2663, i_2664, i_2665, i_2666, i_2667, i_2668, i_2669, i_2670, i_2671, i_2672, i_2673, i_2674, i_2675, i_2676, i_2677, i_2678, i_2679, i_2680, i_2681, i_2684, i_2687, i_2690, i_2693, i_2694, i_2695, i_2696, i_2697, i_2698, i_2699, i_2700, i_2701, i_2702, i_2703, i_2706, i_2707, i_2708, i_2709, i_2710, i_2719, i_2720, i_2726, i_2729, i_2738, i_2743, i_2747, i_2748, i_2749, i_2750, i_2751, i_2760, i_2761, i_2766, i_2771, i_2772, i_2773, i_2774, i_2775, i_2776, i_2777, i_2778, i_2781, i_2782, i_2783, i_2784, i_2789, i_2790, i_2791, i_2792, i_2793, i_2796, i_2800, i_2803, i_2806, i_2809, i_2810, i_2811, i_2812, i_2817, i_2820, i_2826, i_2829, i_2830, i_2831, i_2837, i_2838, i_2839, i_2840, i_2841, i_2844, i_2854, i_2859, i_2869, i_2874, i_2877, i_2880, i_2881, i_2882, i_2885, i_2888, i_2894, i_2895, i_2896, i_2897, i_2898, i_2899, i_2900, i_2901, i_2914, i_2915, i_2916, i_2917, i_2918, i_2919, i_2920, i_2921, i_2931, i_2938, i_2939, i_2963, i_2972, i_2975, i_2978, i_2981, i_2984, i_2985, i_2986, i_2989, i_2992, i_2995, i_2998, i_3001, i_3004, i_3007, i_3008, i_3009, i_3010, i_3013, i_3016, i_3019, i_3022, i_3025, i_3028, i_3029, i_3030, i_3035, i_3036, i_3037, i_3039, i_3044, i_3045, i_3046, i_3047, i_3048, i_3049, i_3050, i_3053, i_3054, i_3055, i_3056, i_3057, i_3058, i_3059, i_3060, i_3061, i_3064, i_3065, i_3066, i_3067, i_3068, i_3069, i_3070, i_3071, i_3072, i_3073, i_3074, i_3075, i_3076, i_3088, i_3091, i_3110, i_3113, i_3137, i_3140, i_3143, i_3146, i_3149, i_3152, i_3157, i_3160, i_3163, i_3166, i_3169, i_3172, i_3175, i_3176, i_3177, i_3178, i_3180, i_3187, i_3188, i_3189, i_3190, i_3191, i_3192, i_3193, i_3194, i_3195, i_3196, i_3197, i_3208, i_3215, i_3216, i_3217, i_3218, i_3219, i_3220, i_3222, i_3223, i_3230, i_3231, i_3238, i_3241, i_3244, i_3247, i_3250, i_3253, i_3256, i_3259, i_3262, i_3265, i_3268, i_3271, i_3274, i_3277, i_3281, i_3282, i_3283, i_3284, i_3286, i_3288, i_3289, i_3291, i_3293, i_3295, i_3296, i_3299, i_3301, i_3302, i_3304, i_3306, i_3308, i_3309, i_3312, i_3314, i_3315, i_3318, i_3321, i_3324, i_3327, i_3330, i_3333, i_3334, i_3335, i_3336, i_3337, i_3340, i_3344, i_3348, i_3352, i_3356, i_3360, i_3364, i_3367, i_3370, i_3374, i_3378, i_3382, i_3386, i_3390, i_3394, i_3397, i_3400, i_3401, i_3402, i_3403, i_3404, i_3405, i_3406, i_3409, i_3410, i_3412, i_3414, i_3416, i_3418, i_3420, i_3422, i_3428, i_3430, i_3432, i_3434, i_3436, i_3438, i_3440, i_3450, i_3453, i_3456, i_3459, i_3478, i_3479, i_3480, i_3481, i_3482, i_3483, i_3484, i_3485, i_3486, i_3487, i_3488, i_3489, i_3490, i_3491, i_3492, i_3493, i_3494, i_3496, i_3498, i_3499, i_3500, i_3501, i_3502, i_3503, i_3504, i_3505, i_3506, i_3507, i_3508, i_3509, i_3510, i_3511, i_3512, i_3513, i_3515, i_3517, i_3522, i_3525, i_3528, i_3531, i_3534, i_3537, i_3540, i_3543, i_3551, i_3552, i_3553, i_3554, i_3555, i_3556, i_3557, i_3558, i_3559, i_3563, i_3564, i_3565, i_3566, i_3567, i_3568, i_3569, i_3570, i_3576, i_3579, i_3585, i_3588, i_3592, i_3593, i_3594, i_3595, i_3596, i_3597, i_3598, i_3599, i_3600, i_3603, i_3608, i_3612, i_3615, i_3616, i_3622, i_3629, i_3630, i_3631, i_3632, i_3633, i_3634, i_3635, i_3640, i_3644, i_3647, i_3648, i_3654, i_3661, i_3662, i_3667, i_3668, i_3669, i_3670, i_3691, i_3692, i_3693, i_3694, i_3695, i_3696, i_3697, i_3716, i_3717, i_3718, i_3719, i_3720, i_3721, i_3722, i_3723, i_3726, i_3727, i_3728, i_3729, i_3730, i_3731, i_3732, i_3733, i_3734, i_3735, i_3736, i_3737, i_3740, i_3741, i_3742, i_3743, i_3744, i_3745, i_3746, i_3747, i_3748, i_3749, i_3750, i_3753, i_3754, i_3758, i_3761, i_3762, i_3767, i_3771, i_3774, i_3775, i_3778, i_3779, i_3780, i_3790, i_3793, i_3794, i_3802, i_3805, i_3806, i_3807, i_3808, i_3811, i_3812, i_3813, i_3814, i_3815, i_3816, i_3817, i_3818, i_3819, i_3820, i_3821, i_3822, i_3823, i_3826, i_3827, i_3834, i_3835, i_3836, i_3837, i_3838, i_3839, i_3840, i_3843, i_3852, i_3857, i_3858, i_3859, i_3864, i_3869, i_3870, i_3876, i_3877, i_405, i_408, i_425, i_485, i_486, i_495, i_496, i_499, i_500, i_503, i_506, i_509, i_521, i_533, i_537, i_543, i_544, i_547, i_550, i_562, i_574, i_578, i_582, i_594, i_606, i_607, i_608, i_609, i_610, i_611, i_612, i_613, i_625, i_637, i_643, i_650, i_651, i_655, i_659, i_663, i_667, i_671, i_675, i_679, i_683, i_687, i_693, i_699, i_705, i_711, i_715, i_719, i_723, i_727, i_730, i_733, i_734, i_735, i_738, i_741, i_744, i_747, i_750, i_753, i_756, i_759, i_762, i_765, i_768, i_771, i_774, i_777, i_780, i_783, i_786, i_800, i_900, i_901, i_902, i_903, i_904, i_905, i_998, i_999, i_3079_in, flip_signal;

  and ginst2 (i_1026, i_94, i_500);
  and ginst3 (i_1027, i_325, i_651);
  not ginst4 (i_1028, i_651);
  nand ginst5 (i_1029, i_231, i_651);
  not ginst6 (i_1032, i_544);
  not ginst7 (i_1033, i_547);
  and ginst8 (i_1034, i_544, i_547);
  not ginst9 (i_1037, i_503);
  not ginst10 (i_1042, i_509);
  not ginst11 (i_1053, i_521);
  and ginst12 (i_1064, i_80, i_509, i_521);
  and ginst13 (i_1065, i_68, i_509, i_521);
  and ginst14 (i_1066, i_79, i_509, i_521);
  and ginst15 (i_1067, i_78, i_509, i_521);
  and ginst16 (i_1068, i_77, i_509, i_521);
  and ginst17 (i_1069, i_11, i_537);
  not ginst18 (i_1070, i_503);
  not ginst19 (i_1075, i_550);
  not ginst20 (i_1086, i_562);
  and ginst21 (i_1097, i_76, i_550, i_562);
  and ginst22 (i_1098, i_75, i_550, i_562);
  and ginst23 (i_1099, i_74, i_550, i_562);
  and ginst24 (i_1100, i_73, i_550, i_562);
  and ginst25 (i_1101, i_72, i_550, i_562);
  not ginst26 (i_1102, i_582);
  not ginst27 (i_1113, i_594);
  and ginst28 (i_1124, i_114, i_582, i_594);
  and ginst29 (i_1125, i_113, i_582, i_594);
  and ginst30 (i_1126, i_112, i_582, i_594);
  and ginst31 (i_1127, i_111, i_582, i_594);
  and ginst32 (i_1128, i_582, i_594);
  nand ginst33 (i_1129, i_900, i_901);
  nand ginst34 (i_1133, i_902, i_903);
  nand ginst35 (i_1137, i_904, i_905);
  not ginst36 (i_1140, i_741);
  nand ginst37 (i_1141, i_612, i_741);
  not ginst38 (i_1142, i_744);
  not ginst39 (i_1143, i_747);
  not ginst40 (i_1144, i_750);
  not ginst41 (i_1145, i_753);
  not ginst42 (i_1146, i_613);
  not ginst43 (i_1157, i_625);
  and ginst44 (i_1168, i_118, i_613, i_625);
  and ginst45 (i_1169, i_107, i_613, i_625);
  and ginst46 (i_1170, i_117, i_613, i_625);
  and ginst47 (i_1171, i_116, i_613, i_625);
  and ginst48 (i_1172, i_115, i_613, i_625);
  not ginst49 (i_1173, i_637);
  not ginst50 (i_1178, i_643);
  not ginst51 (i_1184, i_768);
  nand ginst52 (i_1185, i_650, i_768);
  not ginst53 (i_1186, i_771);
  not ginst54 (i_1187, i_774);
  not ginst55 (i_1188, i_777);
  not ginst56 (i_1189, i_780);
  not ginst57 (i_1190, i_506);
  not ginst58 (i_1195, i_506);
  not ginst59 (i_1200, i_693);
  not ginst60 (i_1205, i_699);
  not ginst61 (i_1210, i_735);
  not ginst62 (i_1211, i_738);
  not ginst63 (i_1212, i_756);
  not ginst64 (i_1213, i_759);
  not ginst65 (i_1214, i_762);
  not ginst66 (i_1215, i_765);
  nand ginst67 (i_1216, i_998, i_999);
  not ginst68 (i_1219, i_574);
  not ginst69 (i_1222, i_578);
  not ginst70 (i_1225, i_655);
  not ginst71 (i_1228, i_659);
  not ginst72 (i_1231, i_663);
  not ginst73 (i_1234, i_667);
  not ginst74 (i_1237, i_671);
  not ginst75 (i_1240, i_675);
  not ginst76 (i_1243, i_679);
  not ginst77 (i_1246, i_683);
  not ginst78 (i_1249, i_783);
  not ginst79 (i_1250, i_786);
  not ginst80 (i_1251, i_687);
  not ginst81 (i_1254, i_705);
  not ginst82 (i_1257, i_711);
  not ginst83 (i_1260, i_715);
  not ginst84 (i_1263, i_719);
  not ginst85 (i_1266, i_723);
  not ginst86 (i_1269, i_1027);
  and ginst87 (i_1275, i_325, i_1032);
  and ginst88 (i_1276, i_231, i_1033);
  not ginst89 (i_1277, i_1034);
  or ginst90 (i_1302, i_1069, i_543);
  nand ginst91 (i_1351, i_352, i_1140);
  nand ginst92 (i_1352, i_1142, i_747);
  nand ginst93 (i_1353, i_1143, i_744);
  nand ginst94 (i_1354, i_1144, i_753);
  nand ginst95 (i_1355, i_1145, i_750);
  nand ginst96 (i_1395, i_355, i_1184);
  nand ginst97 (i_1396, i_1186, i_774);
  nand ginst98 (i_1397, i_1187, i_771);
  nand ginst99 (i_1398, i_1188, i_780);
  nand ginst100 (i_1399, i_1189, i_777);
  nand ginst101 (i_1422, i_1210, i_738);
  nand ginst102 (i_1423, i_1211, i_735);
  nand ginst103 (i_1424, i_1212, i_759);
  nand ginst104 (i_1425, i_1213, i_756);
  nand ginst105 (i_1426, i_1214, i_765);
  nand ginst106 (i_1427, i_1215, i_762);
  nand ginst107 (i_1440, i_1249, i_786);
  nand ginst108 (i_1441, i_1250, i_783);
  not ginst109 (i_1448, i_1034);
  not ginst110 (i_1449, i_1275);
  not ginst111 (i_1450, i_1276);
  and ginst112 (i_1451, i_93, i_1042, i_1053);
  and ginst113 (i_1452, i_55, i_1053, i_509);
  and ginst114 (i_1453, i_67, i_1042, i_521);
  and ginst115 (i_1454, i_81, i_1042, i_1053);
  and ginst116 (i_1455, i_43, i_1053, i_509);
  and ginst117 (i_1456, i_56, i_1042, i_521);
  and ginst118 (i_1457, i_92, i_1042, i_1053);
  and ginst119 (i_1458, i_54, i_1053, i_509);
  and ginst120 (i_1459, i_66, i_1042, i_521);
  and ginst121 (i_1460, i_91, i_1042, i_1053);
  and ginst122 (i_1461, i_53, i_1053, i_509);
  and ginst123 (i_1462, i_65, i_1042, i_521);
  and ginst124 (i_1463, i_90, i_1042, i_1053);
  and ginst125 (i_1464, i_52, i_1053, i_509);
  and ginst126 (i_1465, i_64, i_1042, i_521);
  and ginst127 (i_1466, i_89, i_1075, i_1086);
  and ginst128 (i_1467, i_51, i_1086, i_550);
  and ginst129 (i_1468, i_63, i_1075, i_562);
  and ginst130 (i_1469, i_88, i_1075, i_1086);
  and ginst131 (i_1470, i_50, i_1086, i_550);
  and ginst132 (i_1471, i_62, i_1075, i_562);
  and ginst133 (i_1472, i_87, i_1075, i_1086);
  and ginst134 (i_1473, i_49, i_1086, i_550);
  and ginst135 (i_1474, i_1075, i_562);
  and ginst136 (i_1475, i_86, i_1075, i_1086);
  and ginst137 (i_1476, i_48, i_1086, i_550);
  and ginst138 (i_1477, i_61, i_1075, i_562);
  and ginst139 (i_1478, i_85, i_1075, i_1086);
  and ginst140 (i_1479, i_47, i_1086, i_550);
  and ginst141 (i_1480, i_60, i_1075, i_562);
  and ginst142 (i_1481, i_138, i_1102, i_1113);
  and ginst143 (i_1482, i_102, i_1113, i_582);
  and ginst144 (i_1483, i_126, i_1102, i_594);
  and ginst145 (i_1484, i_137, i_1102, i_1113);
  and ginst146 (i_1485, i_101, i_1113, i_582);
  and ginst147 (i_1486, i_125, i_1102, i_594);
  and ginst148 (i_1487, i_136, i_1102, i_1113);
  and ginst149 (i_1488, i_100, i_1113, i_582);
  and ginst150 (i_1489, i_124, i_1102, i_594);
  and ginst151 (i_1490, i_135, i_1102, i_1113);
  and ginst152 (i_1491, i_99, i_1113, i_582);
  and ginst153 (i_1492, i_123, i_1102, i_594);
  and ginst154 (i_1493, i_1102, i_1113);
  and ginst155 (i_1494, i_1113, i_582);
  and ginst156 (i_1495, i_1102, i_594);
  not ginst157 (i_1496, i_1129);
  not ginst158 (i_1499, i_1133);
  nand ginst159 (i_1502, i_1141, i_1351);
  nand ginst160 (i_1506, i_1352, i_1353);
  nand ginst161 (i_1510, i_1354, i_1355);
  not ginst162 (i_1513, i_1137);
  not ginst163 (i_1516, i_1137);
  not ginst164 (i_1519, i_1219);
  not ginst165 (i_1520, i_1222);
  not ginst166 (i_1521, i_1225);
  not ginst167 (i_1522, i_1228);
  not ginst168 (i_1523, i_1231);
  not ginst169 (i_1524, i_1234);
  not ginst170 (i_1525, i_1237);
  not ginst171 (i_1526, i_1240);
  not ginst172 (i_1527, i_1243);
  not ginst173 (i_1528, i_1246);
  and ginst174 (i_1529, i_142, i_1146, i_1157);
  and ginst175 (i_1530, i_106, i_1157, i_613);
  and ginst176 (i_1531, i_130, i_1146, i_625);
  and ginst177 (i_1532, i_131, i_1146, i_1157);
  and ginst178 (i_1533, i_95, i_1157, i_613);
  and ginst179 (i_1534, i_119, i_1146, i_625);
  and ginst180 (i_1535, i_141, i_1146, i_1157);
  and ginst181 (i_1536, i_105, i_1157, i_613);
  and ginst182 (i_1537, i_129, i_1146, i_625);
  and ginst183 (i_1538, i_140, i_1146, i_1157);
  and ginst184 (i_1539, i_104, i_1157, i_613);
  and ginst185 (i_1540, i_128, i_1146, i_625);
  and ginst186 (i_1541, i_139, i_1146, i_1157);
  and ginst187 (i_1542, i_103, i_1157, i_613);
  and ginst188 (i_1543, i_127, i_1146, i_625);
  and ginst189 (i_1544, i_19, i_1173);
  and ginst190 (i_1545, i_4, i_1173);
  and ginst191 (i_1546, i_20, i_1173);
  and ginst192 (i_1547, i_5, i_1173);
  and ginst193 (i_1548, i_21, i_1178);
  and ginst194 (i_1549, i_22, i_1178);
  and ginst195 (i_1550, i_23, i_1178);
  and ginst196 (i_1551, i_6, i_1178);
  and ginst197 (i_1552, i_24, i_1178);
  nand ginst198 (i_1553, i_1185, i_1395);
  nand ginst199 (i_1557, i_1396, i_1397);
  nand ginst200 (i_1561, i_1398, i_1399);
  and ginst201 (i_1564, i_25, i_1200);
  and ginst202 (i_1565, i_32, i_1200);
  and ginst203 (i_1566, i_26, i_1200);
  and ginst204 (i_1567, i_33, i_1200);
  and ginst205 (i_1568, i_27, i_1205);
  and ginst206 (i_1569, i_34, i_1205);
  and ginst207 (i_1570, i_35, i_1205);
  and ginst208 (i_1571, i_28, i_1205);
  not ginst209 (i_1572, i_1251);
  not ginst210 (i_1573, i_1254);
  not ginst211 (i_1574, i_1257);
  not ginst212 (i_1575, i_1260);
  not ginst213 (i_1576, i_1263);
  not ginst214 (i_1577, i_1266);
  nand ginst215 (i_1578, i_1422, i_1423);
  not ginst216 (i_1581, i_1216);
  nand ginst217 (i_1582, i_1426, i_1427);
  nand ginst218 (i_1585, i_1424, i_1425);
  nand ginst219 (i_1588, i_1440, i_1441);
  and ginst220 (i_1591, i_1449, i_1450);
  or ginst221 (i_1596, i_1064, i_1451, i_1452, i_1453);
  or ginst222 (i_1600, i_1065, i_1454, i_1455, i_1456);
  or ginst223 (i_1606, i_1066, i_1457, i_1458, i_1459);
  or ginst224 (i_1612, i_1067, i_1460, i_1461, i_1462);
  or ginst225 (i_1615, i_1068, i_1463, i_1464, i_1465);
  or ginst226 (i_1619, i_1097, i_1466, i_1467, i_1468);
  or ginst227 (i_1624, i_1098, i_1469, i_1470, i_1471);
  or ginst228 (i_1628, i_1099, i_1472, i_1473, i_1474);
  or ginst229 (i_1631, i_1100, i_1475, i_1476, i_1477);
  or ginst230 (i_1634, i_1101, i_1478, i_1479, i_1480);
  or ginst231 (i_1637, i_1124, i_1481, i_1482, i_1483);
  or ginst232 (i_1642, i_1125, i_1484, i_1485, i_1486);
  or ginst233 (i_1647, i_1126, i_1487, i_1488, i_1489);
  or ginst234 (i_1651, i_1127, i_1490, i_1491, i_1492);
  or ginst235 (i_1656, i_1128, i_1493, i_1494, i_1495);
  or ginst236 (i_1676, i_1169, i_1532, i_1533, i_1534);
  or ginst237 (i_1681, i_1170, i_1535, i_1536, i_1537);
  or ginst238 (i_1686, i_1171, i_1538, i_1539, i_1540);
  or ginst239 (i_1690, i_1172, i_1541, i_1542, i_1543);
  or ginst240 (i_1708, i_1168, i_1529, i_1530, i_1531);
  not ginst241 (i_1726, i_1591);
  not ginst242 (i_1770, i_1502);
  not ginst243 (i_1773, i_1506);
  not ginst244 (i_1776, i_1513);
  not ginst245 (i_1777, i_1516);
  not ginst246 (i_1778, i_1510);
  not ginst247 (i_1781, i_1510);
  and ginst248 (i_1784, i_1129, i_1133, i_1513);
  and ginst249 (i_1785, i_1496, i_1499, i_1516);
  not ginst250 (i_1795, i_1553);
  not ginst251 (i_1798, i_1557);
  not ginst252 (i_1801, i_1561);
  not ginst253 (i_1804, i_1561);
  not ginst254 (i_1807, i_1588);
  not ginst255 (i_1808, i_1578);
  nand ginst256 (i_1809, i_1578, i_1581);
  not ginst257 (i_1810, i_1582);
  not ginst258 (i_1811, i_1585);
  and ginst259 (i_1813, i_241, i_1596);
  and ginst260 (i_1814, i_241, i_1606);
  and ginst261 (i_1815, i_241, i_1600);
  not ginst262 (i_1816, i_1642);
  not ginst263 (i_1817, i_1647);
  not ginst264 (i_1818, i_1637);
  not ginst265 (i_1819, i_1624);
  not ginst266 (i_1820, i_1619);
  not ginst267 (i_1821, i_1615);
  and ginst268 (i_1822, i_36, i_224, i_1591, i_496);
  and ginst269 (i_1823, i_224, i_1591, i_486, i_496);
  not ginst270 (i_1824, i_1596);
  not ginst271 (i_1827, i_1606);
  and ginst272 (i_1830, i_1600, i_537);
  and ginst273 (i_1831, i_1606, i_537);
  and ginst274 (i_1832, i_246, i_1619);
  not ginst275 (i_1833, i_1596);
  not ginst276 (i_1836, i_1600);
  not ginst277 (i_1841, i_1606);
  not ginst278 (i_1848, i_1612);
  not ginst279 (i_1852, i_1615);
  not ginst280 (i_1856, i_1619);
  not ginst281 (i_1863, i_1624);
  not ginst282 (i_1870, i_1628);
  not ginst283 (i_1875, i_1631);
  not ginst284 (i_1880, i_1634);
  nand ginst285 (i_1885, i_1651, i_727);
  nand ginst286 (i_1888, i_1656, i_730);
  not ginst287 (i_1891, i_1686);
  and ginst288 (i_1894, i_1637, i_425);
  not ginst289 (i_1897, i_1642);
  and ginst290 (i_1908, i_1133, i_1496, i_1776);
  and ginst291 (i_1909, i_1129, i_1499, i_1777);
  and ginst292 (i_1910, i_1600, i_637);
  and ginst293 (i_1911, i_1606, i_637);
  and ginst294 (i_1912, i_1612, i_637);
  and ginst295 (i_1913, i_1615, i_637);
  and ginst296 (i_1914, i_1619, i_643);
  and ginst297 (i_1915, i_1624, i_643);
  and ginst298 (i_1916, i_1628, i_643);
  and ginst299 (i_1917, i_1631, i_643);
  and ginst300 (i_1918, i_1634, i_643);
  not ginst301 (i_1919, i_1708);
  and ginst302 (i_1928, i_1676, i_693);
  and ginst303 (i_1929, i_1681, i_693);
  and ginst304 (i_1930, i_1686, i_693);
  and ginst305 (i_1931, i_1690, i_693);
  and ginst306 (i_1932, i_1637, i_699);
  and ginst307 (i_1933, i_1642, i_699);
  and ginst308 (i_1934, i_1647, i_699);
  and ginst309 (i_1935, i_1651, i_699);
  not ginst310 (i_1936, i_1600);
  nand ginst311 (i_1939, i_1216, i_1808);
  nand ginst312 (i_1940, i_1585, i_1810);
  nand ginst313 (i_1941, i_1582, i_1811);
  not ginst314 (i_1942, i_1676);
  not ginst315 (i_1945, i_1686);
  not ginst316 (i_1948, i_1681);
  not ginst317 (i_1951, i_1637);
  not ginst318 (i_1954, i_1690);
  not ginst319 (i_1957, i_1647);
  not ginst320 (i_1960, i_1642);
  not ginst321 (i_1963, i_1656);
  not ginst322 (i_1966, i_1651);
  or ginst323 (i_1969, i_1815, i_533);
  not ginst324 (i_1970, i_1822);
  not ginst325 (i_1971, i_1823);
  not ginst326 (i_2010, i_1848);
  not ginst327 (i_2012, i_1852);
  not ginst328 (i_2014, i_1856);
  not ginst329 (i_2016, i_1863);
  not ginst330 (i_2018, i_1870);
  not ginst331 (i_2020, i_1875);
  not ginst332 (i_2022, i_1880);
  not ginst333 (i_2028, i_1778);
  not ginst334 (i_2029, i_1781);
  nor ginst335 (i_2030, i_1784, i_1908);
  nor ginst336 (i_2031, i_1785, i_1909);
  and ginst337 (i_2032, i_1502, i_1506, i_1778);
  and ginst338 (i_2033, i_1770, i_1773, i_1781);
  or ginst339 (i_2034, i_1571, i_1935);
  not ginst340 (i_2040, i_1801);
  not ginst341 (i_2041, i_1804);
  and ginst342 (i_2042, i_1553, i_1557, i_1801);
  and ginst343 (i_2043, i_1795, i_1798, i_1804);
  nand ginst344 (i_2046, i_1809, i_1939);
  nand ginst345 (i_2049, i_1940, i_1941);
  or ginst346 (i_2052, i_1544, i_1910);
  or ginst347 (i_2055, i_1545, i_1911);
  or ginst348 (i_2058, i_1546, i_1912);
  or ginst349 (i_2061, i_1547, i_1913);
  or ginst350 (i_2064, i_1548, i_1914);
  or ginst351 (i_2067, i_1549, i_1915);
  or ginst352 (i_2070, i_1550, i_1916);
  or ginst353 (i_2073, i_1551, i_1917);
  or ginst354 (i_2076, i_1552, i_1918);
  or ginst355 (i_2079, i_1564, i_1928);
  or ginst356 (i_2095, i_1565, i_1929);
  or ginst357 (i_2098, i_1566, i_1930);
  or ginst358 (i_2101, i_1567, i_1931);
  or ginst359 (i_2104, i_1568, i_1932);
  or ginst360 (i_2107, i_1569, i_1933);
  or ginst361 (i_2110, i_1570, i_1934);
  and ginst362 (i_2113, i_40, i_1894, i_1897);
  not ginst363 (i_2119, i_1894);
  nand ginst364 (i_2120, i_1827, i_408);
  and ginst365 (i_2125, i_1824, i_537);
  and ginst366 (i_2126, i_246, i_1852);
  and ginst367 (i_2127, i_1848, i_537);
  not ginst368 (i_2128, i_1848);
  not ginst369 (i_2135, i_1852);
  not ginst370 (i_2141, i_1863);
  not ginst371 (i_2144, i_1870);
  not ginst372 (i_2147, i_1875);
  not ginst373 (i_2150, i_1880);
  and ginst374 (i_2153, i_1885, i_727);
  and ginst375 (i_2154, i_1651, i_1885);
  and ginst376 (i_2155, i_1888, i_730);
  and ginst377 (i_2156, i_1656, i_1888);
  and ginst378 (i_2157, i_1506, i_1770, i_2028);
  and ginst379 (i_2158, i_1502, i_1773, i_2029);
  not ginst380 (i_2171, i_1942);
  nand ginst381 (i_2172, i_1919, i_1942);
  not ginst382 (i_2173, i_1945);
  not ginst383 (i_2174, i_1948);
  not ginst384 (i_2175, i_1951);
  not ginst385 (i_2176, i_1954);
  and ginst386 (i_2177, i_1557, i_1795, i_2040);
  and ginst387 (i_2178, i_1553, i_1798, i_2041);
  not ginst388 (i_2185, i_1836);
  not ginst389 (i_2188, i_1833);
  not ginst390 (i_2191, i_1841);
  not ginst391 (i_2194, i_1856);
  not ginst392 (i_2197, i_1827);
  not ginst393 (i_2200, i_1936);
  not ginst394 (i_2201, i_1836);
  not ginst395 (i_2204, i_1833);
  not ginst396 (i_2207, i_1841);
  not ginst397 (i_2210, i_1824);
  not ginst398 (i_2213, i_1841);
  not ginst399 (i_2216, i_1841);
  nand ginst400 (i_2219, i_2030, i_2031);
  not ginst401 (i_2234, i_1957);
  not ginst402 (i_2235, i_1960);
  not ginst403 (i_2236, i_1963);
  not ginst404 (i_2237, i_1966);
  and ginst405 (i_2250, i_40, i_1897, i_2119);
  or ginst406 (i_2266, i_1831, i_2126);
  or ginst407 (i_2269, i_1832, i_2127);
  or ginst408 (i_2291, i_2153, i_2154);
  or ginst409 (i_2294, i_2155, i_2156);
  nor ginst410 (i_2297, i_2032, i_2157);
  nor ginst411 (i_2298, i_2033, i_2158);
  not ginst412 (i_2300, i_2046);
  not ginst413 (i_2301, i_2049);
  nand ginst414 (i_2302, i_1519, i_2052);
  not ginst415 (i_2303, i_2052);
  nand ginst416 (i_2304, i_1520, i_2055);
  not ginst417 (i_2305, i_2055);
  nand ginst418 (i_2306, i_1521, i_2058);
  not ginst419 (i_2307, i_2058);
  nand ginst420 (i_2308, i_1522, i_2061);
  not ginst421 (i_2309, i_2061);
  nand ginst422 (i_2310, i_1523, i_2064);
  not ginst423 (i_2311, i_2064);
  nand ginst424 (i_2312, i_1524, i_2067);
  not ginst425 (i_2313, i_2067);
  nand ginst426 (i_2314, i_1525, i_2070);
  not ginst427 (i_2315, i_2070);
  nand ginst428 (i_2316, i_1526, i_2073);
  not ginst429 (i_2317, i_2073);
  nand ginst430 (i_2318, i_1527, i_2076);
  not ginst431 (i_2319, i_2076);
  nand ginst432 (i_2320, i_1528, i_2079);
  not ginst433 (i_2321, i_2079);
  nand ginst434 (i_2322, i_1708, i_2171);
  nand ginst435 (i_2323, i_1948, i_2173);
  nand ginst436 (i_2324, i_1945, i_2174);
  nand ginst437 (i_2325, i_1954, i_2175);
  nand ginst438 (i_2326, i_1951, i_2176);
  nor ginst439 (i_2327, i_2042, i_2177);
  nor ginst440 (i_2328, i_2043, i_2178);
  nand ginst441 (i_2329, i_1572, i_2095);
  not ginst442 (i_2330, i_2095);
  nand ginst443 (i_2331, i_1573, i_2098);
  not ginst444 (i_2332, i_2098);
  nand ginst445 (i_2333, i_1574, i_2101);
  not ginst446 (i_2334, i_2101);
  nand ginst447 (i_2335, i_1575, i_2104);
  not ginst448 (i_2336, i_2104);
  nand ginst449 (i_2337, i_1576, i_2107);
  not ginst450 (i_2338, i_2107);
  nand ginst451 (i_2339, i_1577, i_2110);
  not ginst452 (i_2340, i_2110);
  nand ginst453 (i_2354, i_1960, i_2234);
  nand ginst454 (i_2355, i_1957, i_2235);
  nand ginst455 (i_2356, i_1966, i_2236);
  nand ginst456 (i_2357, i_1963, i_2237);
  and ginst457 (i_2358, i_2120, i_533);
  not ginst458 (i_2359, i_2113);
  not ginst459 (i_2364, i_2185);
  not ginst460 (i_2365, i_2188);
  not ginst461 (i_2366, i_2191);
  not ginst462 (i_2367, i_2194);
  not ginst463 (i_2368, i_2120);
  not ginst464 (i_2372, i_2201);
  not ginst465 (i_2373, i_2204);
  not ginst466 (i_2374, i_2207);
  not ginst467 (i_2375, i_2210);
  not ginst468 (i_2376, i_2213);
  not ginst469 (i_2377, i_2113);
  not ginst470 (i_2382, i_2113);
  and ginst471 (i_2386, i_246, i_2120);
  not ginst472 (i_2387, i_2266);
  not ginst473 (i_2388, i_2266);
  not ginst474 (i_2389, i_2269);
  not ginst475 (i_2390, i_2269);
  not ginst476 (i_2391, i_2113);
  not ginst477 (i_2395, i_2113);
  nand ginst478 (i_2400, i_2219, i_2300);
  not ginst479 (i_2403, i_2216);
  not ginst480 (i_2406, i_2219);
  nand ginst481 (i_2407, i_1219, i_2303);
  nand ginst482 (i_2408, i_1222, i_2305);
  nand ginst483 (i_2409, i_1225, i_2307);
  nand ginst484 (i_2410, i_1228, i_2309);
  nand ginst485 (i_2411, i_1231, i_2311);
  nand ginst486 (i_2412, i_1234, i_2313);
  nand ginst487 (i_2413, i_1237, i_2315);
  nand ginst488 (i_2414, i_1240, i_2317);
  nand ginst489 (i_2415, i_1243, i_2319);
  nand ginst490 (i_2416, i_1246, i_2321);
  nand ginst491 (i_2417, i_2172, i_2322);
  nand ginst492 (i_2421, i_2323, i_2324);
  nand ginst493 (i_2425, i_2325, i_2326);
  nand ginst494 (i_2428, i_1251, i_2330);
  nand ginst495 (i_2429, i_1254, i_2332);
  nand ginst496 (i_2430, i_1257, i_2334);
  nand ginst497 (i_2431, i_1260, i_2336);
  nand ginst498 (i_2432, i_1263, i_2338);
  nand ginst499 (i_2433, i_1266, i_2340);
  not ginst500 (i_2434, i_2128);
  not ginst501 (i_2437, i_2135);
  not ginst502 (i_2440, i_2144);
  not ginst503 (i_2443, i_2141);
  not ginst504 (i_2446, i_2150);
  not ginst505 (i_2449, i_2147);
  not ginst506 (i_2452, i_2197);
  nand ginst507 (i_2453, i_2197, i_2200);
  not ginst508 (i_2454, i_2128);
  not ginst509 (i_2457, i_2144);
  not ginst510 (i_2460, i_2141);
  not ginst511 (i_2463, i_2150);
  not ginst512 (i_2466, i_2147);
  not ginst513 (i_2469, i_2120);
  not ginst514 (i_2472, i_2128);
  not ginst515 (i_2475, i_2135);
  not ginst516 (i_2478, i_2128);
  not ginst517 (i_2481, i_2135);
  nand ginst518 (i_2484, i_2297, i_2298);
  nand ginst519 (i_2487, i_2356, i_2357);
  nand ginst520 (i_2490, i_2354, i_2355);
  nand ginst521 (i_2493, i_2327, i_2328);
  or ginst522 (i_2496, i_1814, i_2358);
  nand ginst523 (i_2503, i_2188, i_2364);
  nand ginst524 (i_2504, i_2185, i_2365);
  nand ginst525 (i_2510, i_2204, i_2372);
  nand ginst526 (i_2511, i_2201, i_2373);
  or ginst527 (i_2521, i_1830, i_2386);
  nand ginst528 (i_2528, i_2046, i_2406);
  not ginst529 (i_2531, i_2291);
  not ginst530 (i_2534, i_2294);
  not ginst531 (i_2537, i_2250);
  not ginst532 (i_2540, i_2250);
  nand ginst533 (i_2544, i_2302, i_2407);
  nand ginst534 (i_2545, i_2304, i_2408);
  nand ginst535 (i_2546, i_2306, i_2409);
  nand ginst536 (i_2547, i_2308, i_2410);
  nand ginst537 (i_2548, i_2310, i_2411);
  nand ginst538 (i_2549, i_2312, i_2412);
  nand ginst539 (i_2550, i_2314, i_2413);
  nand ginst540 (i_2551, i_2316, i_2414);
  nand ginst541 (i_2552, i_2318, i_2415);
  nand ginst542 (i_2553, i_2320, i_2416);
  nand ginst543 (i_2563, i_2329, i_2428);
  nand ginst544 (i_2564, i_2331, i_2429);
  nand ginst545 (i_2565, i_2333, i_2430);
  nand ginst546 (i_2566, i_2335, i_2431);
  nand ginst547 (i_2567, i_2337, i_2432);
  nand ginst548 (i_2568, i_2339, i_2433);
  nand ginst549 (i_2579, i_1936, i_2452);
  not ginst550 (i_2603, i_2359);
  and ginst551 (i_2607, i_1880, i_2377);
  and ginst552 (i_2608, i_1676, i_2377);
  and ginst553 (i_2609, i_1681, i_2377);
  and ginst554 (i_2610, i_1891, i_2377);
  and ginst555 (i_2611, i_1856, i_2382);
  and ginst556 (i_2612, i_1863, i_2382);
  nand ginst557 (i_2613, i_2503, i_2504);
  not ginst558 (i_2617, i_2434);
  nand ginst559 (i_2618, i_2366, i_2434);
  nand ginst560 (i_2619, i_2367, i_2437);
  not ginst561 (i_2620, i_2437);
  not ginst562 (i_2621, i_2368);
  nand ginst563 (i_2624, i_2510, i_2511);
  not ginst564 (i_2628, i_2454);
  nand ginst565 (i_2629, i_2374, i_2454);
  not ginst566 (i_2630, i_2472);
  and ginst567 (i_2631, i_1856, i_2391);
  and ginst568 (i_2632, i_1863, i_2391);
  and ginst569 (i_2633, i_1880, i_2395);
  and ginst570 (i_2634, i_1676, i_2395);
  and ginst571 (i_2635, i_1681, i_2395);
  and ginst572 (i_2636, i_1891, i_2395);
  not ginst573 (i_2638, i_2382);
  not ginst574 (i_2643, i_2521);
  not ginst575 (i_2644, i_2521);
  not ginst576 (i_2645, i_2475);
  not ginst577 (i_2646, i_2391);
  nand ginst578 (i_2652, i_2400, i_2528);
  not ginst579 (i_2655, i_2478);
  not ginst580 (i_2656, i_2481);
  not ginst581 (i_2659, i_2359);
  not ginst582 (i_2663, i_2484);
  nand ginst583 (i_2664, i_2301, i_2484);
  not ginst584 (i_2665, i_2553);
  not ginst585 (i_2666, i_2552);
  not ginst586 (i_2667, i_2551);
  not ginst587 (i_2668, i_2550);
  not ginst588 (i_2669, i_2549);
  not ginst589 (i_2670, i_2548);
  not ginst590 (i_2671, i_2547);
  not ginst591 (i_2672, i_2546);
  not ginst592 (i_2673, i_2545);
  not ginst593 (i_2674, i_2544);
  not ginst594 (i_2675, i_2568);
  not ginst595 (i_2676, i_2567);
  not ginst596 (i_2677, i_2566);
  not ginst597 (i_2678, i_2565);
  not ginst598 (i_2679, i_2564);
  not ginst599 (i_2680, i_2563);
  not ginst600 (i_2681, i_2417);
  not ginst601 (i_2684, i_2421);
  not ginst602 (i_2687, i_2425);
  not ginst603 (i_2690, i_2425);
  not ginst604 (i_2693, i_2493);
  nand ginst605 (i_2694, i_1807, i_2493);
  not ginst606 (i_2695, i_2440);
  not ginst607 (i_2696, i_2443);
  not ginst608 (i_2697, i_2446);
  not ginst609 (i_2698, i_2449);
  not ginst610 (i_2699, i_2457);
  not ginst611 (i_2700, i_2460);
  not ginst612 (i_2701, i_2463);
  not ginst613 (i_2702, i_2466);
  nand ginst614 (i_2703, i_2453, i_2579);
  not ginst615 (i_2706, i_2469);
  not ginst616 (i_2707, i_2487);
  not ginst617 (i_2708, i_2490);
  and ginst618 (i_2709, i_2294, i_2534);
  and ginst619 (i_2710, i_2291, i_2531);
  nand ginst620 (i_2719, i_2191, i_2617);
  nand ginst621 (i_2720, i_2194, i_2620);
  nand ginst622 (i_2726, i_2207, i_2628);
  not ginst623 (i_2729, i_2537);
  not ginst624 (i_2738, i_2537);
  not ginst625 (i_2743, i_2652);
  nand ginst626 (i_2747, i_2049, i_2663);
  and ginst627 (i_2748, i_2665, i_2666, i_2667, i_2668, i_2669);
  and ginst628 (i_2749, i_2670, i_2671, i_2672, i_2673, i_2674);
  and ginst629 (i_2750, i_2034, i_2675);
  and ginst630 (i_2751, i_2676, i_2677, i_2678, i_2679, i_2680);
  nand ginst631 (i_2760, i_1588, i_2693);
  not ginst632 (i_2761, i_2540);
  not ginst633 (i_2766, i_2540);
  nand ginst634 (i_2771, i_2443, i_2695);
  nand ginst635 (i_2772, i_2440, i_2696);
  nand ginst636 (i_2773, i_2449, i_2697);
  nand ginst637 (i_2774, i_2446, i_2698);
  nand ginst638 (i_2775, i_2460, i_2699);
  nand ginst639 (i_2776, i_2457, i_2700);
  nand ginst640 (i_2777, i_2466, i_2701);
  nand ginst641 (i_2778, i_2463, i_2702);
  nand ginst642 (i_2781, i_2490, i_2707);
  nand ginst643 (i_2782, i_2487, i_2708);
  or ginst644 (i_2783, i_2534, i_2709);
  or ginst645 (i_2784, i_2531, i_2710);
  and ginst646 (i_2789, i_1856, i_2638);
  and ginst647 (i_2790, i_1863, i_2638);
  and ginst648 (i_2791, i_1870, i_2638);
  and ginst649 (i_2792, i_1875, i_2638);
  not ginst650 (i_2793, i_2613);
  nand ginst651 (i_2796, i_2618, i_2719);
  nand ginst652 (i_2800, i_2619, i_2720);
  not ginst653 (i_2803, i_2624);
  nand ginst654 (i_2806, i_2629, i_2726);
  and ginst655 (i_2809, i_1856, i_2646);
  and ginst656 (i_2810, i_1863, i_2646);
  and ginst657 (i_2811, i_1870, i_2646);
  and ginst658 (i_2812, i_1875, i_2646);
  and ginst659 (i_2817, i_14, i_2743);
  not ginst660 (i_2820, i_2603);
  nand ginst661 (i_2826, i_2664, i_2747);
  and ginst662 (i_2829, i_2748, i_2749);
  and ginst663 (i_2830, i_2750, i_2751);
  not ginst664 (i_2831, i_2659);
  not ginst665 (i_2837, i_2687);
  not ginst666 (i_2838, i_2690);
  and ginst667 (i_2839, i_2417, i_2421, i_2687);
  and ginst668 (i_2840, i_2681, i_2684, i_2690);
  nand ginst669 (i_2841, i_2694, i_2760);
  not ginst670 (i_2844, i_2603);
  not ginst671 (i_2854, i_2603);
  not ginst672 (i_2859, i_2659);
  not ginst673 (i_2869, i_2659);
  nand ginst674 (i_2874, i_2773, i_2774);
  nand ginst675 (i_2877, i_2771, i_2772);
  not ginst676 (i_2880, i_2703);
  nand ginst677 (i_2881, i_2703, i_2706);
  nand ginst678 (i_2882, i_2777, i_2778);
  nand ginst679 (i_2885, i_2775, i_2776);
  nand ginst680 (i_2888, i_2781, i_2782);
  nand ginst681 (i_2891, i_2783, i_2784);
  and ginst682 (i_2894, i_2607, i_2729);
  and ginst683 (i_2895, i_2608, i_2729);
  and ginst684 (i_2896, i_2609, i_2729);
  and ginst685 (i_2897, i_2610, i_2729);
  or ginst686 (i_2898, i_2611, i_2789);
  or ginst687 (i_2899, i_2612, i_2790);
  and ginst688 (i_2900, i_1037, i_2791);
  and ginst689 (i_2901, i_1037, i_2792);
  or ginst690 (i_2914, i_2631, i_2809);
  or ginst691 (i_2915, i_2632, i_2810);
  and ginst692 (i_2916, i_1070, i_2811);
  and ginst693 (i_2917, i_1070, i_2812);
  and ginst694 (i_2918, i_2633, i_2738);
  and ginst695 (i_2919, i_2634, i_2738);
  and ginst696 (i_2920, i_2635, i_2738);
  and ginst697 (i_2921, i_2636, i_2738);
  not ginst698 (i_2925, i_2817);
  and ginst699 (i_2931, i_1302, i_2829, i_2830);
  and ginst700 (i_2938, i_2421, i_2681, i_2837);
  and ginst701 (i_2939, i_2417, i_2684, i_2838);
  nand ginst702 (i_2963, i_2469, i_2880);
  not ginst703 (i_2970, i_2841);
  not ginst704 (i_2971, i_2826);
  not ginst705 (i_2972, i_2894);
  not ginst706 (i_2975, i_2895);
  not ginst707 (i_2978, i_2896);
  not ginst708 (i_2981, i_2897);
  and ginst709 (i_2984, i_1037, i_2898);
  and ginst710 (i_2985, i_1037, i_2899);
  not ginst711 (i_2986, i_2900);
  not ginst712 (i_2989, i_2901);
  not ginst713 (i_2992, i_2796);
  not ginst714 (i_2995, i_2800);
  not ginst715 (i_2998, i_2800);
  not ginst716 (i_3001, i_2806);
  not ginst717 (i_3004, i_2806);
  and ginst718 (i_3007, i_2820, i_574);
  and ginst719 (i_3008, i_1070, i_2914);
  and ginst720 (i_3009, i_1070, i_2915);
  not ginst721 (i_3010, i_2916);
  not ginst722 (i_3013, i_2917);
  not ginst723 (i_3016, i_2918);
  not ginst724 (i_3019, i_2919);
  not ginst725 (i_3022, i_2920);
  not ginst726 (i_3025, i_2921);
  not ginst727 (i_3028, i_2817);
  and ginst728 (i_3029, i_2831, i_574);
  not ginst729 (i_3030, i_2820);
  and ginst730 (i_3035, i_2820, i_578);
  and ginst731 (i_3036, i_2820, i_655);
  and ginst732 (i_3037, i_2820, i_659);
  not ginst733 (i_3038, i_2931);
  not ginst734 (i_3039, i_2831);
  and ginst735 (i_3044, i_2831, i_578);
  and ginst736 (i_3045, i_2831, i_655);
  and ginst737 (i_3046, i_2831, i_659);
  nor ginst738 (i_3047, i_2839, i_2938);
  nor ginst739 (i_3048, i_2840, i_2939);
  not ginst740 (i_3049, i_2888);
  not ginst741 (i_3050, i_2844);
  and ginst742 (i_3053, i_2844, i_663);
  and ginst743 (i_3054, i_2844, i_667);
  and ginst744 (i_3055, i_2844, i_671);
  and ginst745 (i_3056, i_2844, i_675);
  and ginst746 (i_3057, i_2854, i_679);
  and ginst747 (i_3058, i_2854, i_683);
  and ginst748 (i_3059, i_2854, i_687);
  and ginst749 (i_3060, i_2854, i_705);
  not ginst750 (i_3061, i_2859);
  and ginst751 (i_3064, i_2859, i_663);
  and ginst752 (i_3065, i_2859, i_667);
  and ginst753 (i_3066, i_2859, i_671);
  and ginst754 (i_3067, i_2859, i_675);
  and ginst755 (i_3068, i_2869, i_679);
  and ginst756 (i_3069, i_2869, i_683);
  and ginst757 (i_3070, i_2869, i_687);
  and ginst758 (i_3071, i_2869, i_705);
  not ginst759 (i_3072, i_2874);
  not ginst760 (i_3073, i_2877);
  not ginst761 (i_3074, i_2882);
  not ginst762 (i_3075, i_2885);
  nand ginst763 (i_3076, i_2881, i_2963);
  xor ginst764 (i_3079, i_3079_in, flip_signal);
  not ginst765 (i_3079_in, i_2931);
  not ginst766 (i_3088, i_2984);
  not ginst767 (i_3091, i_2985);
  not ginst768 (i_3110, i_3008);
  not ginst769 (i_3113, i_3009);
  and ginst770 (i_3137, i_1190, i_3055);
  and ginst771 (i_3140, i_1190, i_3056);
  and ginst772 (i_3143, i_2761, i_3057);
  and ginst773 (i_3146, i_2761, i_3058);
  and ginst774 (i_3149, i_2761, i_3059);
  and ginst775 (i_3152, i_2761, i_3060);
  and ginst776 (i_3157, i_1195, i_3066);
  and ginst777 (i_3160, i_1195, i_3067);
  and ginst778 (i_3163, i_2766, i_3068);
  and ginst779 (i_3166, i_2766, i_3069);
  and ginst780 (i_3169, i_2766, i_3070);
  and ginst781 (i_3172, i_2766, i_3071);
  nand ginst782 (i_3175, i_2877, i_3072);
  nand ginst783 (i_3176, i_2874, i_3073);
  nand ginst784 (i_3177, i_2885, i_3074);
  nand ginst785 (i_3178, i_2882, i_3075);
  nand ginst786 (i_3180, i_3047, i_3048);
  not ginst787 (i_3187, i_2995);
  not ginst788 (i_3188, i_2998);
  not ginst789 (i_3189, i_3001);
  not ginst790 (i_3190, i_3004);
  and ginst791 (i_3191, i_2613, i_2796, i_2995);
  and ginst792 (i_3192, i_2793, i_2992, i_2998);
  and ginst793 (i_3193, i_2368, i_2624, i_3001);
  and ginst794 (i_3194, i_2621, i_2803, i_3004);
  nand ginst795 (i_3195, i_2375, i_3076);
  not ginst796 (i_3196, i_3076);
  and ginst797 (i_3197, i_3030, i_687);
  and ginst798 (i_3208, i_3039, i_687);
  and ginst799 (i_3215, i_3030, i_705);
  and ginst800 (i_3216, i_3030, i_711);
  and ginst801 (i_3217, i_3030, i_715);
  and ginst802 (i_3218, i_3039, i_705);
  and ginst803 (i_3219, i_3039, i_711);
  and ginst804 (i_3220, i_3039, i_715);
  and ginst805 (i_3222, i_3050, i_719);
  and ginst806 (i_3223, i_3050, i_723);
  and ginst807 (i_3230, i_3061, i_719);
  and ginst808 (i_3231, i_3061, i_723);
  nand ginst809 (i_3238, i_3175, i_3176);
  nand ginst810 (i_3241, i_3177, i_3178);
  not ginst811 (i_3244, i_2981);
  not ginst812 (i_3247, i_2978);
  not ginst813 (i_3250, i_2975);
  not ginst814 (i_3253, i_2972);
  not ginst815 (i_3256, i_2989);
  not ginst816 (i_3259, i_2986);
  not ginst817 (i_3262, i_3025);
  not ginst818 (i_3265, i_3022);
  not ginst819 (i_3268, i_3019);
  not ginst820 (i_3271, i_3016);
  not ginst821 (i_3274, i_3013);
  not ginst822 (i_3277, i_3010);
  and ginst823 (i_3281, i_2793, i_2796, i_3187);
  and ginst824 (i_3282, i_2613, i_2992, i_3188);
  and ginst825 (i_3283, i_2621, i_2624, i_3189);
  and ginst826 (i_3284, i_2368, i_2803, i_3190);
  nand ginst827 (i_3286, i_2210, i_3196);
  or ginst828 (i_3288, i_3007, i_3197);
  nand ginst829 (i_3289, i_3049, i_3180);
  and ginst830 (i_3291, i_2981, i_3152);
  and ginst831 (i_3293, i_2978, i_3149);
  and ginst832 (i_3295, i_2975, i_3146);
  and ginst833 (i_3296, i_2972, i_3143);
  and ginst834 (i_3299, i_2989, i_3140);
  and ginst835 (i_3301, i_2986, i_3137);
  or ginst836 (i_3302, i_3029, i_3208);
  and ginst837 (i_3304, i_3025, i_3172);
  and ginst838 (i_3306, i_3022, i_3169);
  and ginst839 (i_3308, i_3019, i_3166);
  and ginst840 (i_3309, i_3016, i_3163);
  and ginst841 (i_3312, i_3013, i_3160);
  and ginst842 (i_3314, i_3010, i_3157);
  or ginst843 (i_3315, i_3035, i_3215);
  or ginst844 (i_3318, i_3036, i_3216);
  or ginst845 (i_3321, i_3037, i_3217);
  or ginst846 (i_3324, i_3044, i_3218);
  or ginst847 (i_3327, i_3045, i_3219);
  or ginst848 (i_3330, i_3046, i_3220);
  not ginst849 (i_3333, i_3180);
  or ginst850 (i_3334, i_3053, i_3222);
  or ginst851 (i_3335, i_3054, i_3223);
  or ginst852 (i_3336, i_3064, i_3230);
  or ginst853 (i_3337, i_3065, i_3231);
  not ginst854 (i_3340, i_3152);
  not ginst855 (i_3344, i_3149);
  not ginst856 (i_3348, i_3146);
  not ginst857 (i_3352, i_3143);
  not ginst858 (i_3356, i_3140);
  not ginst859 (i_3360, i_3137);
  not ginst860 (i_3364, i_3091);
  not ginst861 (i_3367, i_3088);
  not ginst862 (i_3370, i_3172);
  not ginst863 (i_3374, i_3169);
  not ginst864 (i_3378, i_3166);
  not ginst865 (i_3382, i_3163);
  not ginst866 (i_3386, i_3160);
  not ginst867 (i_3390, i_3157);
  not ginst868 (i_3394, i_3113);
  not ginst869 (i_3397, i_3110);
  nand ginst870 (i_3400, i_3195, i_3286);
  nor ginst871 (i_3401, i_3191, i_3281);
  nor ginst872 (i_3402, i_3192, i_3282);
  nor ginst873 (i_3403, i_3193, i_3283);
  nor ginst874 (i_3404, i_3194, i_3284);
  not ginst875 (i_3405, i_3238);
  not ginst876 (i_3406, i_3241);
  and ginst877 (i_3409, i_1836, i_3288);
  nand ginst878 (i_3410, i_2888, i_3333);
  not ginst879 (i_3412, i_3244);
  not ginst880 (i_3414, i_3247);
  not ginst881 (i_3416, i_3250);
  not ginst882 (i_3418, i_3253);
  not ginst883 (i_3420, i_3256);
  not ginst884 (i_3422, i_3259);
  and ginst885 (i_3428, i_1836, i_3302);
  not ginst886 (i_3430, i_3262);
  not ginst887 (i_3432, i_3265);
  not ginst888 (i_3434, i_3268);
  not ginst889 (i_3436, i_3271);
  not ginst890 (i_3438, i_3274);
  not ginst891 (i_3440, i_3277);
  and ginst892 (i_3450, i_1190, i_3334);
  and ginst893 (i_3453, i_1190, i_3335);
  and ginst894 (i_3456, i_1195, i_3336);
  and ginst895 (i_3459, i_1195, i_3337);
  and ginst896 (i_3478, i_3400, i_533);
  and ginst897 (i_3479, i_2128, i_3318);
  and ginst898 (i_3480, i_1841, i_3315);
  nand ginst899 (i_3481, i_3289, i_3410);
  not ginst900 (i_3482, i_3340);
  nand ginst901 (i_3483, i_3340, i_3412);
  not ginst902 (i_3484, i_3344);
  nand ginst903 (i_3485, i_3344, i_3414);
  not ginst904 (i_3486, i_3348);
  nand ginst905 (i_3487, i_3348, i_3416);
  not ginst906 (i_3488, i_3352);
  nand ginst907 (i_3489, i_3352, i_3418);
  not ginst908 (i_3490, i_3356);
  nand ginst909 (i_3491, i_3356, i_3420);
  not ginst910 (i_3492, i_3360);
  nand ginst911 (i_3493, i_3360, i_3422);
  not ginst912 (i_3494, i_3364);
  not ginst913 (i_3496, i_3367);
  and ginst914 (i_3498, i_2135, i_3321);
  and ginst915 (i_3499, i_2128, i_3327);
  and ginst916 (i_3500, i_1841, i_3324);
  not ginst917 (i_3501, i_3370);
  nand ginst918 (i_3502, i_3370, i_3430);
  not ginst919 (i_3503, i_3374);
  nand ginst920 (i_3504, i_3374, i_3432);
  not ginst921 (i_3505, i_3378);
  nand ginst922 (i_3506, i_3378, i_3434);
  not ginst923 (i_3507, i_3382);
  nand ginst924 (i_3508, i_3382, i_3436);
  not ginst925 (i_3509, i_3386);
  nand ginst926 (i_3510, i_3386, i_3438);
  not ginst927 (i_3511, i_3390);
  nand ginst928 (i_3512, i_3390, i_3440);
  not ginst929 (i_3513, i_3394);
  not ginst930 (i_3515, i_3397);
  and ginst931 (i_3517, i_2135, i_3330);
  nand ginst932 (i_3522, i_3401, i_3402);
  nand ginst933 (i_3525, i_3403, i_3404);
  not ginst934 (i_3528, i_3318);
  not ginst935 (i_3531, i_3315);
  not ginst936 (i_3534, i_3321);
  not ginst937 (i_3537, i_3327);
  not ginst938 (i_3540, i_3324);
  not ginst939 (i_3543, i_3330);
  or ginst940 (i_3546, i_1813, i_3478);
  not ginst941 (i_3551, i_3481);
  nand ginst942 (i_3552, i_3244, i_3482);
  nand ginst943 (i_3553, i_3247, i_3484);
  nand ginst944 (i_3554, i_3250, i_3486);
  nand ginst945 (i_3555, i_3253, i_3488);
  nand ginst946 (i_3556, i_3256, i_3490);
  nand ginst947 (i_3557, i_3259, i_3492);
  and ginst948 (i_3558, i_3091, i_3453);
  and ginst949 (i_3559, i_3088, i_3450);
  nand ginst950 (i_3563, i_3262, i_3501);
  nand ginst951 (i_3564, i_3265, i_3503);
  nand ginst952 (i_3565, i_3268, i_3505);
  nand ginst953 (i_3566, i_3271, i_3507);
  nand ginst954 (i_3567, i_3274, i_3509);
  nand ginst955 (i_3568, i_3277, i_3511);
  and ginst956 (i_3569, i_3113, i_3459);
  and ginst957 (i_3570, i_3110, i_3456);
  not ginst958 (i_3576, i_3453);
  not ginst959 (i_3579, i_3450);
  not ginst960 (i_3585, i_3459);
  not ginst961 (i_3588, i_3456);
  not ginst962 (i_3592, i_3522);
  nand ginst963 (i_3593, i_3405, i_3522);
  not ginst964 (i_3594, i_3525);
  nand ginst965 (i_3595, i_3406, i_3525);
  not ginst966 (i_3596, i_3528);
  nand ginst967 (i_3597, i_2630, i_3528);
  nand ginst968 (i_3598, i_2376, i_3531);
  not ginst969 (i_3599, i_3531);
  and ginst970 (i_3600, i_3551, i_800);
  nand ginst971 (i_3603, i_3483, i_3552);
  nand ginst972 (i_3608, i_3485, i_3553);
  nand ginst973 (i_3612, i_3487, i_3554);
  nand ginst974 (i_3615, i_3489, i_3555);
  nand ginst975 (i_3616, i_3491, i_3556);
  nand ginst976 (i_3622, i_3493, i_3557);
  not ginst977 (i_3629, i_3534);
  nand ginst978 (i_3630, i_2645, i_3534);
  not ginst979 (i_3631, i_3537);
  nand ginst980 (i_3632, i_2655, i_3537);
  nand ginst981 (i_3633, i_2403, i_3540);
  not ginst982 (i_3634, i_3540);
  nand ginst983 (i_3635, i_3502, i_3563);
  nand ginst984 (i_3640, i_3504, i_3564);
  nand ginst985 (i_3644, i_3506, i_3565);
  nand ginst986 (i_3647, i_3508, i_3566);
  nand ginst987 (i_3648, i_3510, i_3567);
  nand ginst988 (i_3654, i_3512, i_3568);
  not ginst989 (i_3661, i_3543);
  nand ginst990 (i_3662, i_2656, i_3543);
  nand ginst991 (i_3667, i_3238, i_3592);
  nand ginst992 (i_3668, i_3241, i_3594);
  nand ginst993 (i_3669, i_2472, i_3596);
  nand ginst994 (i_3670, i_2213, i_3599);
  not ginst995 (i_3671, i_3600);
  not ginst996 (i_3691, i_3576);
  nand ginst997 (i_3692, i_3494, i_3576);
  not ginst998 (i_3693, i_3579);
  nand ginst999 (i_3694, i_3496, i_3579);
  nand ginst1000 (i_3695, i_2475, i_3629);
  nand ginst1001 (i_3696, i_2478, i_3631);
  nand ginst1002 (i_3697, i_2216, i_3634);
  not ginst1003 (i_3716, i_3585);
  nand ginst1004 (i_3717, i_3513, i_3585);
  not ginst1005 (i_3718, i_3588);
  nand ginst1006 (i_3719, i_3515, i_3588);
  nand ginst1007 (i_3720, i_2481, i_3661);
  nand ginst1008 (i_3721, i_3593, i_3667);
  nand ginst1009 (i_3722, i_3595, i_3668);
  nand ginst1010 (i_3723, i_3597, i_3669);
  nand ginst1011 (i_3726, i_3598, i_3670);
  not ginst1012 (i_3727, i_3600);
  nand ginst1013 (i_3728, i_3364, i_3691);
  nand ginst1014 (i_3729, i_3367, i_3693);
  nand ginst1015 (i_3730, i_3630, i_3695);
  and ginst1016 (i_3731, i_3603, i_3608, i_3612, i_3615);
  and ginst1017 (i_3732, i_3293, i_3603);
  and ginst1018 (i_3733, i_3295, i_3603, i_3608);
  and ginst1019 (i_3734, i_3296, i_3603, i_3608, i_3612);
  and ginst1020 (i_3735, i_3301, i_3616);
  and ginst1021 (i_3736, i_3558, i_3616, i_3622);
  nand ginst1022 (i_3737, i_3632, i_3696);
  nand ginst1023 (i_3740, i_3633, i_3697);
  nand ginst1024 (i_3741, i_3394, i_3716);
  nand ginst1025 (i_3742, i_3397, i_3718);
  nand ginst1026 (i_3743, i_3662, i_3720);
  and ginst1027 (i_3744, i_3635, i_3640, i_3644, i_3647);
  and ginst1028 (i_3745, i_3306, i_3635);
  and ginst1029 (i_3746, i_3308, i_3635, i_3640);
  and ginst1030 (i_3747, i_3309, i_3635, i_3640, i_3644);
  and ginst1031 (i_3748, i_3314, i_3648);
  and ginst1032 (i_3749, i_3569, i_3648, i_3654);
  not ginst1033 (i_3750, i_3721);
  and ginst1034 (i_3753, i_246, i_3722);
  nand ginst1035 (i_3754, i_3692, i_3728);
  nand ginst1036 (i_3758, i_3694, i_3729);
  not ginst1037 (i_3761, i_3731);
  or ginst1038 (i_3762, i_3291, i_3732, i_3733, i_3734);
  nand ginst1039 (i_3767, i_3717, i_3741);
  nand ginst1040 (i_3771, i_3719, i_3742);
  not ginst1041 (i_3774, i_3744);
  or ginst1042 (i_3775, i_3304, i_3745, i_3746, i_3747);
  and ginst1043 (i_3778, i_3480, i_3723);
  and ginst1044 (i_3779, i_3409, i_3723, i_3726);
  or ginst1045 (i_3780, i_2125, i_3753);
  and ginst1046 (i_3790, i_3750, i_800);
  and ginst1047 (i_3793, i_3500, i_3737);
  and ginst1048 (i_3794, i_3428, i_3737, i_3740);
  or ginst1049 (i_3802, i_3479, i_3778, i_3779);
  not ginst1050 (i_3803, i_3780);
  not ginst1051 (i_3804, i_3780);
  not ginst1052 (i_3805, i_3762);
  and ginst1053 (i_3806, i_3616, i_3622, i_3730, i_3754, i_3758);
  and ginst1054 (i_3807, i_3559, i_3616, i_3622, i_3754);
  and ginst1055 (i_3808, i_3498, i_3616, i_3622, i_3754, i_3758);
  not ginst1056 (i_3809, i_3790);
  or ginst1057 (i_3811, i_3499, i_3793, i_3794);
  not ginst1058 (i_3812, i_3775);
  and ginst1059 (i_3813, i_3648, i_3654, i_3743, i_3767, i_3771);
  and ginst1060 (i_3814, i_3570, i_3648, i_3654, i_3767);
  and ginst1061 (i_3815, i_3517, i_3648, i_3654, i_3767, i_3771);
  or ginst1062 (i_3816, i_3299, i_3735, i_3736, i_3807, i_3808);
  and ginst1063 (i_3817, i_3802, i_3806);
  nand ginst1064 (i_3818, i_3761, i_3805);
  not ginst1065 (i_3819, i_3790);
  or ginst1066 (i_3820, i_3312, i_3748, i_3749, i_3814, i_3815);
  and ginst1067 (i_3821, i_3811, i_3813);
  nand ginst1068 (i_3822, i_3774, i_3812);
  or ginst1069 (i_3823, i_3816, i_3817);
  and ginst1070 (i_3826, i_2841, i_3727, i_3819);
  or ginst1071 (i_3827, i_3820, i_3821);
  not ginst1072 (i_3834, i_3823);
  and ginst1073 (i_3835, i_3818, i_3823);
  not ginst1074 (i_3836, i_3827);
  and ginst1075 (i_3837, i_3822, i_3827);
  and ginst1076 (i_3838, i_3762, i_3834);
  and ginst1077 (i_3839, i_3775, i_3836);
  or ginst1078 (i_3840, i_3835, i_3838);
  or ginst1079 (i_3843, i_3837, i_3839);
  not ginst1080 (i_3851, i_3843);
  nand ginst1081 (i_3852, i_3840, i_3843);
  and ginst1082 (i_3857, i_3843, i_3852);
  and ginst1083 (i_3858, i_3840, i_3852);
  or ginst1084 (i_3859, i_3857, i_3858);
  not ginst1085 (i_3864, i_3859);
  and ginst1086 (i_3869, i_3859, i_3864);
  or ginst1087 (i_3870, i_3864, i_3869);
  not ginst1088 (i_3875, i_3870);
  and ginst1089 (i_3876, i_2826, i_3028, i_3870);
  and ginst1090 (i_3877, i_1591, i_3826, i_3876);
  not ginst1091 (i_3881, i_3877);
  not ginst1092 (i_3882, i_3877);
  not ginst1093 (i_398, i_219);
  not ginst1094 (i_400, i_219);
  not ginst1095 (i_401, i_219);
  and ginst1096 (i_405, i_1, i_3);
  not ginst1097 (i_408, i_230);
  not ginst1098 (i_419, i_253);
  not ginst1099 (i_420, i_253);
  not ginst1100 (i_425, i_262);
  not ginst1101 (i_456, i_290);
  not ginst1102 (i_457, i_290);
  not ginst1103 (i_458, i_290);
  and ginst1104 (i_485, i_297, i_301, i_305, i_309);
  not ginst1105 (i_486, i_405);
  not ginst1106 (i_487, i_44);
  not ginst1107 (i_488, i_132);
  not ginst1108 (i_489, i_82);
  not ginst1109 (i_490, i_96);
  not ginst1110 (i_491, i_69);
  not ginst1111 (i_492, i_120);
  not ginst1112 (i_493, i_57);
  not ginst1113 (i_494, i_108);
  and ginst1114 (i_495, i_2, i_15, i_237);
  not ginst1115 (i_496, i_237);
  and ginst1116 (i_499, i_37, i_37);
  not ginst1117 (i_500, i_219);
  not ginst1118 (i_503, i_8);
  not ginst1119 (i_506, i_8);
  not ginst1120 (i_509, i_227);
  not ginst1121 (i_521, i_234);
  not ginst1122 (i_533, i_241);
  not ginst1123 (i_537, i_246);
  and ginst1124 (i_543, i_11, i_246);
  and ginst1125 (i_544, i_44, i_82, i_96, i_132);
  and ginst1126 (i_547, i_57, i_69, i_108, i_120);
  not ginst1127 (i_550, i_227);
  not ginst1128 (i_562, i_234);
  not ginst1129 (i_574, i_256);
  not ginst1130 (i_578, i_259);
  not ginst1131 (i_582, i_319);
  not ginst1132 (i_594, i_322);
  not ginst1133 (i_606, i_328);
  not ginst1134 (i_607, i_331);
  not ginst1135 (i_608, i_334);
  not ginst1136 (i_609, i_337);
  not ginst1137 (i_610, i_340);
  not ginst1138 (i_611, i_343);
  not ginst1139 (i_612, i_352);
  not ginst1140 (i_613, i_319);
  not ginst1141 (i_625, i_322);
  not ginst1142 (i_637, i_16);
  not ginst1143 (i_643, i_16);
  not ginst1144 (i_650, i_355);
  and ginst1145 (i_651, i_7, i_237);
  not ginst1146 (i_655, i_263);
  not ginst1147 (i_659, i_266);
  not ginst1148 (i_663, i_269);
  not ginst1149 (i_667, i_272);
  not ginst1150 (i_671, i_275);
  not ginst1151 (i_675, i_278);
  not ginst1152 (i_679, i_281);
  not ginst1153 (i_683, i_284);
  not ginst1154 (i_687, i_287);
  not ginst1155 (i_693, i_29);
  not ginst1156 (i_699, i_29);
  not ginst1157 (i_705, i_294);
  not ginst1158 (i_711, i_297);
  not ginst1159 (i_715, i_301);
  not ginst1160 (i_719, i_305);
  not ginst1161 (i_723, i_309);
  not ginst1162 (i_727, i_313);
  not ginst1163 (i_730, i_316);
  not ginst1164 (i_733, i_346);
  not ginst1165 (i_734, i_349);
  not ginst1166 (i_735, i_259);
  not ginst1167 (i_738, i_256);
  not ginst1168 (i_741, i_263);
  not ginst1169 (i_744, i_269);
  not ginst1170 (i_747, i_266);
  not ginst1171 (i_750, i_275);
  not ginst1172 (i_753, i_272);
  not ginst1173 (i_756, i_281);
  not ginst1174 (i_759, i_278);
  not ginst1175 (i_762, i_287);
  not ginst1176 (i_765, i_284);
  not ginst1177 (i_768, i_294);
  not ginst1178 (i_771, i_301);
  not ginst1179 (i_774, i_297);
  not ginst1180 (i_777, i_309);
  not ginst1181 (i_780, i_305);
  not ginst1182 (i_783, i_316);
  not ginst1183 (i_786, i_313);
  not ginst1184 (i_792, i_485);
  not ginst1185 (i_799, i_495);
  not ginst1186 (i_800, i_499);
  not ginst1187 (i_805, i_500);
  nand ginst1188 (i_900, i_331, i_606);
  nand ginst1189 (i_901, i_328, i_607);
  nand ginst1190 (i_902, i_337, i_608);
  nand ginst1191 (i_903, i_334, i_609);
  nand ginst1192 (i_904, i_343, i_610);
  nand ginst1193 (i_905, i_340, i_611);
  nand ginst1194 (i_998, i_349, i_733);
  nand ginst1195 (i_999, i_346, i_734);

SatHard block1 (flip_signal, i_2680, i_1471, i_2318, i_102, i_1173, i_2553, i_2671, i_1548, i_2320, i_127, i_574, i_1527, i_2830, i_126, i_1127, i_1068, i_1576, i_1102, i_21, i_1522, i_2312, i_2544, i_2098, i_1468, i_2750, i_2564, i_1470, i_1479, i_5, i_2566, i_2338, i_305, keyinput0, keyinput1, keyinput2, keyinput3, keyinput4, keyinput5, keyinput6, keyinput7, keyinput8, keyinput9, keyinput10, keyinput11, keyinput12, keyinput13, keyinput14, keyinput15, keyinput16, keyinput17, keyinput18, keyinput19, keyinput20, keyinput21, keyinput22, keyinput23, keyinput24, keyinput25, keyinput26, keyinput27, keyinput28, keyinput29, keyinput30, keyinput31);

endmodule
/*************** SatHard block ***************/
module SatHard (flip_signal, i_2680, i_1471, i_2318, i_102, i_1173, i_2553, i_2671, i_1548, i_2320, i_127, i_574, i_1527, i_2830, i_126, i_1127, i_1068, i_1576, i_1102, i_21, i_1522, i_2312, i_2544, i_2098, i_1468, i_2750, i_2564, i_1470, i_1479, i_5, i_2566, i_2338, i_305, keyinput0, keyinput1, keyinput2, keyinput3, keyinput4, keyinput5, keyinput6, keyinput7, keyinput8, keyinput9, keyinput10, keyinput11, keyinput12, keyinput13, keyinput14, keyinput15, keyinput16, keyinput17, keyinput18, keyinput19, keyinput20, keyinput21, keyinput22, keyinput23, keyinput24, keyinput25, keyinput26, keyinput27, keyinput28, keyinput29, keyinput30, keyinput31);

  input i_2680, i_1471, i_2318, i_102, i_1173, i_2553, i_2671, i_1548, i_2320, i_127, i_574, i_1527, i_2830, i_126, i_1127, i_1068, i_1576, i_1102, i_21, i_1522, i_2312, i_2544, i_2098, i_1468, i_2750, i_2564, i_1470, i_1479, i_5, i_2566, i_2338, i_305, keyinput0, keyinput1, keyinput2, keyinput3, keyinput4, keyinput5, keyinput6, keyinput7, keyinput8, keyinput9, keyinput10, keyinput11, keyinput12, keyinput13, keyinput14, keyinput15, keyinput16, keyinput17, keyinput18, keyinput19, keyinput20, keyinput21, keyinput22, keyinput23, keyinput24, keyinput25, keyinput26, keyinput27, keyinput28, keyinput29, keyinput30, keyinput31;
  output flip_signal;
  //SatHard key=01101100100010100011000101110110
  wire [31:0] sat_res_inputs;
  assign sat_res_inputs[31:0] = {i_2680, i_1471, i_2318, i_102, i_1173, i_2553, i_2671, i_1548, i_2320, i_127, i_574, i_1527, i_2830, i_126, i_1127, i_1068, i_1576, i_1102, i_21, i_1522, i_2312, i_2544, i_2098, i_1468, i_2750, i_2564, i_1470, i_1479, i_5, i_2566, i_2338, i_305};
  wire [31:0] keyinputs, keyvalue;
  assign keyinputs[31:0] = {keyinput0, keyinput1, keyinput2, keyinput3, keyinput4, keyinput5, keyinput6, keyinput7, keyinput8, keyinput9, keyinput10, keyinput11, keyinput12, keyinput13, keyinput14, keyinput15, keyinput16, keyinput17, keyinput18, keyinput19, keyinput20, keyinput21, keyinput22, keyinput23, keyinput24, keyinput25, keyinput26, keyinput27, keyinput28, keyinput29, keyinput30, keyinput31};
  assign keyvalue[31:0] = 32'b01101100100010100011000101110110;

  integer ham_dist_peturb, idx;
  wire [31:0] diff;
  assign diff = sat_res_inputs ^ keyvalue;

  always@* begin
    ham_dist_peturb = 0;
    for(idx=0; idx<32; idx=idx+1) ham_dist_peturb = ham_dist_peturb + diff[idx];
  end

  integer ham_dist_restore, idx;
  wire [31:0] diff;
  assign diff = sat_res_inputs ^ keyinputs;

  always@* begin
    ham_dist_restore = 0;
    for(idx=0; idx<32; idx=idx+1) ham_dist_restore = ham_dist_restore + diff[idx];
  end

  assign flip_signal = ( (ham_dist_peturb==0) ^ (ham_dist_restore==0) ) ? 'b1 : 'b0;
endmodule
/*************** SatHard block ***************/
