// Main module
module c5315(1, 4, 11, 14, 17, 20, 23, 24, 25, 26, 27, 31, 34, 37, 40, 43, 46, 49, 52, 53, 54, 61, 64, 67, 70, 73, 76, 79, 80, 81, 82, 83, 86, 87, 88, 91, 94, 97, 100, 103, 106, 109, 112, 113, 114, 115, 116, 117, 118, 119, 120, 121, 122, 123, 126, 127, 128, 129, 130, 131, 132, 135, 136, 137, 140, 141, 145, 146, 149, 152, 155, 158, 161, 164, 167, 170, 173, 176, 179, 182, 185, 188, 191, 194, 197, 200, 203, 206, 209, 210, 217, 218, 225, 226, 233, 234, 241, 242, 245, 248, 251, 254, 257, 264, 265, 272, 273, 280, 281, 288, 289, 292, 293, 299, 302, 307, 308, 315, 316, 323, 324, 331, 332, 335, 338, 341, 348, 351, 358, 361, 366, 369, 372, 373, 374, 386, 389, 400, 411, 422, 435, 446, 457, 468, 479, 490, 503, 514, 523, 534, 545, 549, 552, 556, 559, 562, 566, 571, 574, 577, 580, 583, 588, 591, 592, 595, 596, 597, 598, 599, 603, 607, 610, 613, 616, 619, 625, 631, 709, 816, 1066, 1137, 1138, 1139, 1140, 1141, 1142, 1143, 1144, 1145, 1147, 1152, 1153, 1154, 1155, 1972, 2054, 2060, 2061, 2139, 2142, 2309, 2387, 2527, 2584, 2590, 2623, 3357, 3358, 3359, 3360, 3604, 3613, 4272, 4275, 4278, 4279, 4737, 4738, 4739, 4740, 5240, 5388, 6641, 6643, 6646, 6648, 6716, 6877, 6924, 6925, 6926, 6927, 7015, 7363, 7365, 7432, 7449, 7465, 7466, 7467, 7469, 7470, 7471, 7472, 7473, 7474, 7476, 7503, 7504, 7506, 7511, 7515, 7516, 7517, 7518, 7519, 7520, 7521, 7522, 7600, 7601, 7602, 7603, 7604, 7605, 7606, 7607, 7626, 7698, 7699, 7700, 7701, 7702, 7703, 7704, 7705, 7706, 7707, 7735, 7736, 7737, 7738, 7739, 7740, 7741, 7742, 7754, 7755, 7756, 7757, 7758, 7759, 7760, 7761, 8075, 8076, 8123, 8124, 8127, 8128);

  input 1, 4, 11, 14, 17, 20, 23, 24, 25, 26, 27, 31, 34, 37, 40, 43, 46, 49, 52, 53, 54, 61, 64, 67, 70, 73, 76, 79, 80, 81, 82, 83, 86, 87, 88, 91, 94, 97, 100, 103, 106, 109, 112, 113, 114, 115, 116, 117, 118, 119, 120, 121, 122, 123, 126, 127, 128, 129, 130, 131, 132, 135, 136, 137, 140, 141, 145, 146, 149, 152, 155, 158, 161, 164, 167, 170, 173, 176, 179, 182, 185, 188, 191, 194, 197, 200, 203, 206, 209, 210, 217, 218, 225, 226, 233, 234, 241, 242, 245, 248, 251, 254, 257, 264, 265, 272, 273, 280, 281, 288, 289, 292, 293, 299, 302, 307, 308, 315, 316, 323, 324, 331, 332, 335, 338, 341, 348, 351, 358, 361, 366, 369, 372, 373, 374, 386, 389, 400, 411, 422, 435, 446, 457, 468, 479, 490, 503, 514, 523, 534, 545, 549, 552, 556, 559, 562, 566, 571, 574, 577, 580, 583, 588, 591, 592, 595, 596, 597, 598, 599, 603, 607, 610, 613, 616, 619, 625, 631;
  output 709, 816, 1066, 1137, 1138, 1139, 1140, 1141, 1142, 1143, 1144, 1145, 1147, 1152, 1153, 1154, 1155, 1972, 2054, 2060, 2061, 2139, 2142, 2309, 2387, 2527, 2584, 2590, 2623, 3357, 3358, 3359, 3360, 3604, 3613, 4272, 4275, 4278, 4279, 4737, 4738, 4739, 4740, 5240, 5388, 6641, 6643, 6646, 6648, 6716, 6877, 6924, 6925, 6926, 6927, 7015, 7363, 7365, 7432, 7449, 7465, 7466, 7467, 7469, 7470, 7471, 7472, 7473, 7474, 7476, 7503, 7504, 7506, 7511, 7515, 7516, 7517, 7518, 7519, 7520, 7521, 7522, 7600, 7601, 7602, 7603, 7604, 7605, 7606, 7607, 7626, 7698, 7699, 7700, 7701, 7702, 7703, 7704, 7705, 7706, 7707, 7735, 7736, 7737, 7738, 7739, 7740, 7741, 7742, 7754, 7755, 7756, 7757, 7758, 7759, 7760, 7761, 8075, 8076, 8123, 8124, 8127, 8128;
  wire 1042, 1043, 1067, 1080, 1092, 1104, 1146, 1148, 1149, 1150, 1151, 1156, 1157, 1161, 1173, 1185, 1197, 1209, 1213, 1216, 1219, 1223, 1235, 1247, 1259, 1271, 1280, 1292, 1303, 1315, 1327, 1339, 1351, 1363, 1375, 1378, 1381, 1384, 1387, 1390, 1393, 1396, 1415, 1418, 1421, 1424, 1427, 1430, 1433, 1436, 1455, 1462, 1469, 1475, 1479, 1482, 1492, 1495, 1498, 1501, 1504, 1507, 1510, 1513, 1516, 1519, 1522, 1525, 1542, 1545, 1548, 1551, 1554, 1557, 1560, 1563, 1566, 1573, 1580, 1583, 1588, 1594, 1597, 1600, 1603, 1606, 1609, 1612, 1615, 1618, 1621, 1624, 1627, 1630, 1633, 1636, 1639, 1642, 1645, 1648, 1651, 1654, 1657, 1660, 1663, 1675, 1685, 1697, 1709, 1721, 1727, 1731, 1743, 1755, 1758, 1761, 1769, 1777, 1785, 1793, 1800, 1807, 1814, 1821, 1824, 1827, 1830, 1833, 1836, 1839, 1842, 1845, 1848, 1851, 1854, 1857, 1860, 1863, 1866, 1869, 1872, 1875, 1878, 1881, 1884, 1887, 1890, 1893, 1896, 1899, 1902, 1905, 1908, 1911, 1914, 1917, 1920, 1923, 1926, 1929, 1932, 1935, 1938, 1941, 1944, 1947, 1950, 1953, 1956, 1959, 1962, 1965, 1968, 2349, 2350, 2585, 2586, 2587, 2588, 2589, 2591, 2592, 2593, 2594, 2595, 2596, 2597, 2598, 2599, 2600, 2601, 2602, 2603, 2604, 2605, 2606, 2607, 2608, 2609, 2610, 2611, 2612, 2613, 2614, 2615, 2616, 2617, 2618, 2619, 2620, 2621, 2622, 2624, 2625, 2626, 2627, 2628, 2629, 2630, 2631, 2632, 2633, 2634, 2635, 2636, 2637, 2638, 2639, 2640, 2641, 2642, 2643, 2644, 2645, 2646, 2647, 2653, 2664, 2675, 2681, 2692, 2703, 2704, 2709, 2710, 2711, 2712, 2713, 2714, 2715, 2716, 2717, 2718, 2719, 2720, 2721, 2722, 2728, 2739, 2750, 2756, 2767, 2778, 2779, 2790, 2801, 2812, 2823, 2824, 2825, 2826, 2827, 2828, 2829, 2830, 2831, 2832, 2833, 2834, 2835, 2836, 2837, 2838, 2839, 2840, 2841, 2842, 2843, 2844, 2845, 2846, 2847, 2848, 2849, 2850, 2851, 2852, 2853, 2854, 2855, 2861, 2867, 2868, 2869, 2870, 2871, 2872, 2873, 2874, 2875, 2876, 2877, 2882, 2891, 2901, 2902, 2903, 2904, 2905, 2906, 2907, 2908, 2909, 2910, 2911, 2912, 2913, 2914, 2915, 2916, 2917, 2918, 2919, 2920, 2921, 2922, 2923, 2924, 2925, 2926, 2927, 2928, 2929, 2930, 2931, 2932, 2933, 2934, 2935, 2936, 2937, 2938, 2939, 2940, 2941, 2942, 2948, 2954, 2955, 2956, 2957, 2958, 2959, 2960, 2961, 2962, 2963, 2964, 2969, 2970, 2971, 2972, 2973, 2974, 2975, 2976, 2977, 2978, 2979, 2980, 2981, 2982, 2983, 2984, 2985, 2986, 2987, 2988, 2989, 2990, 2991, 2992, 2993, 2994, 2995, 2996, 2997, 2998, 2999, 3000, 3003, 3006, 3007, 3010, 3013, 3014, 3015, 3016, 3017, 3018, 3019, 3020, 3021, 3022, 3023, 3024, 3025, 3026, 3027, 3028, 3029, 3030, 3031, 3032, 3033, 3034, 3035, 3038, 3041, 3052, 3063, 3068, 3071, 3072, 3073, 3074, 3075, 3086, 3097, 3108, 3119, 3130, 3141, 3142, 3143, 3144, 3145, 3146, 3147, 3158, 3169, 3180, 3191, 3194, 3195, 3196, 3197, 3198, 3199, 3200, 3203, 3401, 3402, 3403, 3404, 3405, 3406, 3407, 3408, 3409, 3410, 3411, 3412, 3413, 3414, 3415, 3416, 3444, 3445, 3446, 3447, 3448, 3449, 3450, 3451, 3452, 3453, 3454, 3455, 3456, 3459, 3460, 3461, 3462, 3463, 3464, 3465, 3466, 3481, 3482, 3483, 3484, 3485, 3486, 3487, 3488, 3489, 3490, 3491, 3492, 3493, 3502, 3503, 3504, 3505, 3506, 3507, 3508, 3509, 3510, 3511, 3512, 3513, 3514, 3515, 3558, 3559, 3560, 3561, 3562, 3563, 3605, 3606, 3607, 3608, 3609, 3610, 3614, 3615, 3616, 3617, 3618, 3619, 3620, 3621, 3622, 3623, 3624, 3625, 3626, 3627, 3628, 3629, 3630, 3631, 3632, 3633, 3634, 3635, 3636, 3637, 3638, 3639, 3640, 3641, 3642, 3643, 3644, 3645, 3646, 3647, 3648, 3649, 3650, 3651, 3652, 3653, 3654, 3655, 3656, 3657, 3658, 3659, 3660, 3661, 3662, 3663, 3664, 3665, 3666, 3667, 3668, 3669, 3670, 3671, 3672, 3673, 3674, 3675, 3676, 3677, 3678, 3679, 3680, 3681, 3682, 3683, 3684, 3685, 3686, 3687, 3688, 3689, 3691, 3700, 3701, 3702, 3703, 3704, 3705, 3708, 3709, 3710, 3711, 3712, 3713, 3715, 3716, 3717, 3718, 3719, 3720, 3721, 3722, 3723, 3724, 3725, 3726, 3727, 3728, 3729, 3730, 3731, 3732, 3738, 3739, 3740, 3741, 3742, 3743, 3744, 3745, 3746, 3747, 3748, 3749, 3750, 3751, 3752, 3753, 3754, 3755, 3756, 3757, 3758, 3759, 3760, 3761, 3762, 3763, 3764, 3765, 3766, 3767, 3768, 3769, 3770, 3771, 3775, 3779, 3780, 3781, 3782, 3783, 3784, 3785, 3786, 3787, 3788, 3789, 3793, 3797, 3800, 3801, 3802, 3803, 3804, 3805, 3806, 3807, 3808, 3809, 3810, 3813, 3816, 3819, 3822, 3823, 3824, 3827, 3828, 3829, 3830, 3831, 3834, 3835, 3836, 3837, 3838, 3839, 3840, 3841, 3842, 3849, 3855, 3861, 3867, 3873, 3881, 3887, 3893, 3908, 3909, 3911, 3914, 3915, 3916, 3917, 3918, 3919, 3920, 3921, 3927, 3933, 3942, 3948, 3956, 3962, 3968, 3975, 3976, 3977, 3978, 3979, 3980, 3981, 3982, 3983, 3984, 3987, 3988, 3989, 3990, 3991, 3998, 4008, 4011, 4021, 4024, 4027, 4031, 4032, 4033, 4034, 4035, 4036, 4037, 4038, 4039, 4040, 4041, 4042, 4067, 4080, 4088, 4091, 4094, 4097, 4100, 4103, 4106, 4109, 4144, 4147, 4150, 4153, 4156, 4159, 4183, 4184, 4185, 4186, 4188, 4191, 4196, 4197, 4198, 4199, 4200, 4203, 4206, 4209, 4212, 4215, 4219, 4223, 4224, 4225, 4228, 4231, 4234, 4237, 4240, 4243, 4246, 4249, 4252, 4255, 4258, 4263, 4264, 4267, 4268, 4269, 4270, 4271, 4273, 4274, 4276, 4277, 4280, 4284, 4290, 4297, 4298, 4301, 4305, 4310, 4316, 4320, 4325, 4331, 4332, 4336, 4342, 4349, 4357, 4364, 4375, 4379, 4385, 4392, 4396, 4400, 4405, 4412, 4418, 4425, 4436, 4440, 4445, 4451, 4456, 4462, 4469, 4477, 4512, 4515, 4516, 4521, 4523, 4524, 4532, 4547, 4548, 4551, 4554, 4557, 4560, 4563, 4566, 4569, 4572, 4575, 4578, 4581, 4584, 4587, 4590, 4593, 4596, 4599, 4602, 4605, 4608, 4611, 4614, 4617, 4621, 4624, 4627, 4630, 4633, 4637, 4640, 4643, 4646, 4649, 4652, 4655, 4658, 4662, 4665, 4668, 4671, 4674, 4677, 4680, 4683, 4686, 4689, 4692, 4695, 4698, 4701, 4702, 4720, 4721, 4724, 4725, 4726, 4727, 4728, 4729, 4730, 4731, 4732, 4733, 4734, 4735, 4736, 4741, 4855, 4856, 4908, 4909, 4939, 4942, 4947, 4953, 4954, 4955, 4956, 4957, 4958, 4959, 4960, 4961, 4965, 4966, 4967, 4968, 4972, 4973, 4974, 4975, 4976, 4977, 4978, 4979, 4980, 4981, 4982, 4983, 4984, 4985, 4986, 4987, 5049, 5052, 5053, 5054, 5055, 5056, 5057, 5058, 5059, 5060, 5061, 5062, 5063, 5065, 5066, 5067, 5068, 5069, 5070, 5071, 5072, 5073, 5074, 5075, 5076, 5077, 5078, 5079, 5080, 5081, 5082, 5083, 5084, 5085, 5086, 5087, 5088, 5089, 5090, 5091, 5092, 5093, 5094, 5095, 5096, 5097, 5098, 5099, 5100, 5101, 5102, 5103, 5104, 5105, 5106, 5107, 5108, 5109, 5110, 5111, 5112, 5113, 5114, 5115, 5116, 5117, 5118, 5119, 5120, 5121, 5122, 5123, 5124, 5125, 5126, 5127, 5128, 5129, 5130, 5131, 5132, 5133, 5135, 5136, 5137, 5138, 5139, 5140, 5141, 5142, 5143, 5144, 5145, 5146, 5147, 5148, 5150, 5153, 5154, 5155, 5156, 5157, 5160, 5161, 5162, 5163, 5164, 5165, 5166, 5169, 5172, 5173, 5176, 5177, 5180, 5183, 5186, 5189, 5192, 5195, 5198, 5199, 5202, 5205, 5208, 5211, 5214, 5217, 5220, 5223, 5224, 5225, 5226, 5227, 5228, 5229, 5230, 5232, 5233, 5234, 5235, 5236, 5239, 5241, 5242, 5243, 5244, 5245, 5246, 5247, 5248, 5249, 5250, 5252, 5253, 5254, 5255, 5256, 5257, 5258, 5259, 5260, 5261, 5262, 5263, 5264, 5274, 5275, 5282, 5283, 5284, 5298, 5299, 5300, 5303, 5304, 5305, 5306, 5307, 5308, 5309, 5310, 5311, 5312, 5315, 5319, 5324, 5328, 5331, 5332, 5346, 5363, 5364, 5365, 5366, 5367, 5368, 5369, 5370, 5371, 5374, 5377, 5382, 5385, 5389, 5396, 5407, 5418, 5424, 5431, 5441, 5452, 5462, 5469, 5470, 5477, 5488, 5498, 5506, 5520, 5536, 5549, 5555, 5562, 5573, 5579, 5595, 5606, 5616, 5617, 5618, 5619, 5620, 5621, 5622, 5624, 5634, 5655, 5671, 5684, 5690, 5691, 5692, 5696, 5700, 5703, 5707, 5711, 5726, 5727, 5728, 5730, 5731, 5732, 5733, 5734, 5735, 5736, 5739, 5742, 5745, 5755, 5756, 5954, 5955, 5956, 6005, 6006, 6023, 6024, 6025, 6028, 6031, 6034, 6037, 6040, 6044, 6045, 6048, 6051, 6054, 6065, 6066, 6067, 6068, 6069, 6071, 6072, 6073, 6074, 6075, 6076, 6077, 6078, 6079, 6080, 6083, 6084, 6085, 6086, 6087, 6088, 6089, 6090, 6091, 6094, 6095, 6096, 6097, 6098, 6099, 6100, 6101, 6102, 6103, 6104, 6105, 6106, 6107, 6108, 6111, 6112, 6113, 6114, 6115, 6116, 6117, 6120, 6121, 6122, 6123, 6124, 6125, 6126, 6127, 6128, 6129, 6130, 6131, 6132, 6133, 6134, 6135, 6136, 6137, 6138, 6139, 6140, 6143, 6144, 6145, 6146, 6147, 6148, 6149, 6152, 6153, 6154, 6155, 6156, 6157, 6158, 6159, 6160, 6161, 6162, 6163, 6164, 6168, 6171, 6172, 6173, 6174, 6175, 6178, 6179, 6180, 6181, 6182, 6183, 6184, 6185, 6186, 6187, 6188, 6189, 6190, 6191, 6192, 6193, 6194, 6197, 6200, 6203, 6206, 6209, 6212, 6215, 6218, 6221, 6234, 6235, 6238, 6241, 6244, 6247, 6250, 6253, 6256, 6259, 6262, 6265, 6268, 6271, 6274, 6277, 6280, 6283, 6286, 6289, 6292, 6295, 6298, 6301, 6304, 6307, 6310, 6313, 6316, 6319, 6322, 6325, 6328, 6331, 6335, 6338, 6341, 6344, 6347, 6350, 6353, 6356, 6359, 6364, 6367, 6370, 6373, 6374, 6375, 6376, 6377, 6378, 6382, 6386, 6388, 6392, 6397, 6411, 6415, 6419, 6427, 6434, 6437, 6441, 6445, 6448, 6449, 6466, 6469, 6470, 6471, 6472, 6473, 6474, 6475, 6476, 6477, 6478, 6482, 6486, 6490, 6494, 6500, 6504, 6508, 6512, 6516, 6526, 6536, 6539, 6553, 6556, 6566, 6569, 6572, 6575, 6580, 6584, 6587, 6592, 6599, 6606, 6609, 6619, 6622, 6630, 6631, 6632, 6633, 6634, 6637, 6640, 6650, 6651, 6653, 6655, 6657, 6659, 6660, 6661, 6662, 6663, 6664, 6666, 6668, 6670, 6672, 6675, 6680, 6681, 6682, 6683, 6689, 6690, 6691, 6692, 6693, 6695, 6698, 6699, 6700, 6703, 6708, 6709, 6710, 6711, 6712, 6713, 6714, 6715, 6718, 6719, 6720, 6721, 6722, 6724, 6739, 6740, 6741, 6744, 6745, 6746, 6751, 6752, 6753, 6754, 6755, 6760, 6761, 6762, 6772, 6773, 6776, 6777, 6782, 6783, 6784, 6785, 6790, 6791, 6792, 6795, 6801, 6802, 6803, 6804, 6805, 6806, 6807, 6808, 6809, 6810, 6811, 6812, 6813, 6814, 6815, 6816, 6817, 6823, 6824, 6825, 6826, 6827, 6828, 6829, 6830, 6831, 6834, 6835, 6836, 6837, 6838, 6839, 6840, 6841, 6842, 6843, 6844, 6850, 6851, 6852, 6853, 6854, 6855, 6856, 6857, 6860, 6861, 6862, 6863, 6866, 6872, 6873, 6874, 6875, 6876, 6879, 6880, 6881, 6884, 6885, 6888, 6889, 6890, 6891, 6894, 6895, 6896, 6897, 6900, 6901, 6904, 6905, 6908, 6909, 6912, 6913, 6914, 6915, 6916, 6919, 6922, 6923, 6930, 6932, 6935, 6936, 6937, 6938, 6939, 6940, 6946, 6947, 6948, 6949, 6953, 6954, 6955, 6956, 6957, 6958, 6964, 6965, 6966, 6967, 6973, 6974, 6975, 6976, 6977, 6978, 6979, 6987, 6990, 6999, 7002, 7003, 7006, 7011, 7012, 7013, 7016, 7018, 7019, 7020, 7021, 7022, 7023, 7028, 7031, 7034, 7037, 7040, 7041, 7044, 7045, 7046, 7047, 7048, 7049, 7054, 7057, 7060, 7064, 7065, 7072, 7073, 7074, 7075, 7076, 7079, 7080, 7083, 7084, 7085, 7086, 7087, 7088, 7089, 7090, 7093, 7094, 7097, 7101, 7105, 7110, 7114, 7115, 7116, 7125, 7126, 7127, 7130, 7131, 7139, 7140, 7141, 7146, 7147, 7149, 7150, 7151, 7152, 7153, 7158, 7159, 7160, 7166, 7167, 7168, 7169, 7170, 7171, 7172, 7173, 7174, 7175, 7176, 7177, 7178, 7179, 7180, 7181, 7182, 7183, 7184, 7185, 7186, 7187, 7188, 7189, 7190, 7196, 7197, 7198, 7204, 7205, 7206, 7207, 7208, 7209, 7212, 7215, 7216, 7217, 7218, 7219, 7222, 7225, 7228, 7229, 7236, 7239, 7242, 7245, 7250, 7257, 7260, 7263, 7268, 7269, 7270, 7276, 7282, 7288, 7294, 7300, 7301, 7304, 7310, 7320, 7321, 7328, 7338, 7339, 7340, 7341, 7342, 7349, 7357, 7364, 7394, 7397, 7402, 7405, 7406, 7407, 7408, 7409, 7412, 7415, 7416, 7417, 7418, 7419, 7420, 7421, 7424, 7425, 7426, 7427, 7428, 7429, 7430, 7431, 7433, 7434, 7435, 7436, 7437, 7438, 7439, 7440, 7441, 7442, 7443, 7444, 7445, 7446, 7447, 7448, 7450, 7451, 7452, 7453, 7454, 7455, 7456, 7457, 7458, 7459, 7460, 7461, 7462, 7463, 7464, 7468, 7479, 7481, 7482, 7483, 7484, 7485, 7486, 7487, 7488, 7489, 7492, 7493, 7498, 7499, 7500, 7505, 7507, 7508, 7509, 7510, 7512, 7513, 7514, 7525, 7526, 7527, 7528, 7529, 7530, 7531, 7537, 7543, 7549, 7555, 7561, 7567, 7573, 7579, 7582, 7585, 7586, 7587, 7588, 7589, 7592, 7595, 7598, 7599, 7624, 7625, 7631, 7636, 7657, 7658, 7665, 7666, 7667, 7668, 7669, 7670, 7671, 7672, 7673, 7674, 7675, 7676, 7677, 7678, 7679, 7680, 7681, 7682, 7683, 7684, 7685, 7686, 7687, 7688, 7689, 7690, 7691, 7692, 7693, 7694, 7695, 7696, 7697, 7708, 7709, 7710, 7711, 7712, 7715, 7718, 7719, 7720, 7721, 7722, 7723, 7724, 7727, 7728, 7729, 7730, 7731, 7732, 7733, 7734, 7743, 7744, 7749, 7750, 7751, 7762, 7765, 7768, 7769, 7770, 7771, 7772, 7775, 7778, 7781, 7782, 7787, 7788, 7795, 7796, 7797, 7798, 7799, 7800, 7803, 7806, 7807, 7808, 7809, 7810, 7811, 7812, 7815, 7816, 7821, 7822, 7823, 7826, 7829, 7832, 7833, 7834, 7835, 7836, 7839, 7842, 7845, 7846, 7851, 7852, 7859, 7860, 7861, 7862, 7863, 7864, 7867, 7870, 7871, 7872, 7873, 7874, 7875, 7876, 7879, 7880, 7885, 7886, 7887, 7890, 7893, 7896, 7897, 7898, 7899, 7900, 7903, 7906, 7909, 7910, 7917, 7918, 7923, 7924, 7925, 7926, 7927, 7928, 7929, 7930, 7931, 7932, 7935, 7938, 7939, 7940, 7943, 7944, 7945, 7946, 7951, 7954, 7957, 7960, 7963, 7966, 7967, 7968, 7969, 7970, 7973, 7974, 7984, 7985, 7987, 7988, 7989, 7990, 7991, 7992, 7993, 7994, 7995, 7996, 7997, 7998, 8001, 8004, 8009, 8013, 8017, 8020, 8021, 8022, 8023, 8025, 8026, 8027, 8031, 8032, 8033, 8034, 8035, 8036, 8037, 8038, 8039, 8040, 8041, 8042, 8043, 8044, 8045, 8048, 8055, 8056, 8057, 8058, 8059, 8060, 8061, 8064, 8071, 8072, 8073, 8074, 8077, 8078, 8079, 8082, 8089, 8090, 8091, 8092, 8093, 8096, 8099, 8102, 8113, 8114, 8115, 8116, 8117, 8118, 8119, 8120, 8121, 8122, 8125, 8126;

  and ginst1 (1042, 135, 631);
  not ginst2 (1043, 591);
  buf ginst3 (1066, 592);
  not ginst4 (1067, 595);
  not ginst5 (1080, 596);
  not ginst6 (1092, 597);
  not ginst7 (1104, 598);
  not ginst8 (1137, 545);
  not ginst9 (1138, 348);
  not ginst10 (1139, 366);
  and ginst11 (1140, 552, 562);
  not ginst12 (1141, 549);
  not ginst13 (1142, 545);
  not ginst14 (1143, 545);
  not ginst15 (1144, 338);
  not ginst16 (1145, 358);
  nand ginst17 (1146, 373, 1);
  and ginst18 (1147, 141, 145);
  not ginst19 (1148, 592);
  not ginst20 (1149, 1042);
  and ginst21 (1150, 1043, 27);
  and ginst22 (1151, 386, 556);
  not ginst23 (1152, 245);
  not ginst24 (1153, 552);
  not ginst25 (1154, 562);
  not ginst26 (1155, 559);
  and ginst27 (1156, 386, 559, 556, 552);
  not ginst28 (1157, 566);
  buf ginst29 (1161, 571);
  buf ginst30 (1173, 574);
  buf ginst31 (1185, 571);
  buf ginst32 (1197, 574);
  buf ginst33 (1209, 137);
  buf ginst34 (1213, 137);
  buf ginst35 (1216, 141);
  not ginst36 (1219, 583);
  buf ginst37 (1223, 577);
  buf ginst38 (1235, 580);
  buf ginst39 (1247, 577);
  buf ginst40 (1259, 580);
  buf ginst41 (1271, 254);
  buf ginst42 (1280, 251);
  buf ginst43 (1292, 251);
  buf ginst44 (1303, 248);
  buf ginst45 (1315, 248);
  buf ginst46 (1327, 610);
  buf ginst47 (1339, 607);
  buf ginst48 (1351, 613);
  buf ginst49 (1363, 616);
  buf ginst50 (1375, 210);
  buf ginst51 (1378, 210);
  buf ginst52 (1381, 218);
  buf ginst53 (1384, 218);
  buf ginst54 (1387, 226);
  buf ginst55 (1390, 226);
  buf ginst56 (1393, 234);
  buf ginst57 (1396, 234);
  buf ginst58 (1415, 257);
  buf ginst59 (1418, 257);
  buf ginst60 (1421, 265);
  buf ginst61 (1424, 265);
  buf ginst62 (1427, 273);
  buf ginst63 (1430, 273);
  buf ginst64 (1433, 281);
  buf ginst65 (1436, 281);
  buf ginst66 (1455, 335);
  buf ginst67 (1462, 335);
  buf ginst68 (1469, 206);
  and ginst69 (1475, 27, 31);
  buf ginst70 (1479, 1);
  buf ginst71 (1482, 588);
  buf ginst72 (1492, 293);
  buf ginst73 (1495, 302);
  buf ginst74 (1498, 308);
  buf ginst75 (1501, 308);
  buf ginst76 (1504, 316);
  buf ginst77 (1507, 316);
  buf ginst78 (1510, 324);
  buf ginst79 (1513, 324);
  buf ginst80 (1516, 341);
  buf ginst81 (1519, 341);
  buf ginst82 (1522, 351);
  buf ginst83 (1525, 351);
  buf ginst84 (1542, 257);
  buf ginst85 (1545, 257);
  buf ginst86 (1548, 265);
  buf ginst87 (1551, 265);
  buf ginst88 (1554, 273);
  buf ginst89 (1557, 273);
  buf ginst90 (1560, 281);
  buf ginst91 (1563, 281);
  buf ginst92 (1566, 332);
  buf ginst93 (1573, 332);
  buf ginst94 (1580, 549);
  and ginst95 (1583, 31, 27);
  not ginst96 (1588, 588);
  buf ginst97 (1594, 324);
  buf ginst98 (1597, 324);
  buf ginst99 (1600, 341);
  buf ginst100 (1603, 341);
  buf ginst101 (1606, 351);
  buf ginst102 (1609, 351);
  buf ginst103 (1612, 293);
  buf ginst104 (1615, 302);
  buf ginst105 (1618, 308);
  buf ginst106 (1621, 308);
  buf ginst107 (1624, 316);
  buf ginst108 (1627, 316);
  buf ginst109 (1630, 361);
  buf ginst110 (1633, 361);
  buf ginst111 (1636, 210);
  buf ginst112 (1639, 210);
  buf ginst113 (1642, 218);
  buf ginst114 (1645, 218);
  buf ginst115 (1648, 226);
  buf ginst116 (1651, 226);
  buf ginst117 (1654, 234);
  buf ginst118 (1657, 234);
  not ginst119 (1660, 324);
  buf ginst120 (1663, 242);
  buf ginst121 (1675, 242);
  buf ginst122 (1685, 254);
  buf ginst123 (1697, 610);
  buf ginst124 (1709, 607);
  buf ginst125 (1721, 625);
  buf ginst126 (1727, 619);
  buf ginst127 (1731, 613);
  buf ginst128 (1743, 616);
  not ginst129 (1755, 599);
  not ginst130 (1758, 603);
  buf ginst131 (1761, 619);
  buf ginst132 (1769, 625);
  buf ginst133 (1777, 619);
  buf ginst134 (1785, 625);
  buf ginst135 (1793, 619);
  buf ginst136 (1800, 625);
  buf ginst137 (1807, 619);
  buf ginst138 (1814, 625);
  buf ginst139 (1821, 299);
  buf ginst140 (1824, 446);
  buf ginst141 (1827, 457);
  buf ginst142 (1830, 468);
  buf ginst143 (1833, 422);
  buf ginst144 (1836, 435);
  buf ginst145 (1839, 389);
  buf ginst146 (1842, 400);
  buf ginst147 (1845, 411);
  buf ginst148 (1848, 374);
  buf ginst149 (1851, 4);
  buf ginst150 (1854, 446);
  buf ginst151 (1857, 457);
  buf ginst152 (1860, 468);
  buf ginst153 (1863, 435);
  buf ginst154 (1866, 389);
  buf ginst155 (1869, 400);
  buf ginst156 (1872, 411);
  buf ginst157 (1875, 422);
  buf ginst158 (1878, 374);
  buf ginst159 (1881, 479);
  buf ginst160 (1884, 490);
  buf ginst161 (1887, 503);
  buf ginst162 (1890, 514);
  buf ginst163 (1893, 523);
  buf ginst164 (1896, 534);
  buf ginst165 (1899, 54);
  buf ginst166 (1902, 479);
  buf ginst167 (1905, 503);
  buf ginst168 (1908, 514);
  buf ginst169 (1911, 523);
  buf ginst170 (1914, 534);
  buf ginst171 (1917, 490);
  buf ginst172 (1920, 361);
  buf ginst173 (1923, 369);
  buf ginst174 (1926, 341);
  buf ginst175 (1929, 351);
  buf ginst176 (1932, 308);
  buf ginst177 (1935, 316);
  buf ginst178 (1938, 293);
  buf ginst179 (1941, 302);
  buf ginst180 (1944, 281);
  buf ginst181 (1947, 289);
  buf ginst182 (1950, 265);
  buf ginst183 (1953, 273);
  buf ginst184 (1956, 234);
  buf ginst185 (1959, 257);
  buf ginst186 (1962, 218);
  buf ginst187 (1965, 226);
  buf ginst188 (1968, 210);
  not ginst189 (1972, 1146);
  and ginst190 (2054, 136, 1148);
  not ginst191 (2060, 1150);
  not ginst192 (2061, 1151);
  buf ginst193 (2139, 1209);
  buf ginst194 (2142, 1216);
  buf ginst195 (2309, 1479);
  and ginst196 (2349, 1104, 514);
  or ginst197 (2350, 1067, 514);
  buf ginst198 (2387, 1580);
  buf ginst199 (2527, 1821);
  not ginst200 (2584, 1580);
  and ginst201 (2585, 170, 1161, 1173);
  and ginst202 (2586, 173, 1161, 1173);
  and ginst203 (2587, 167, 1161, 1173);
  and ginst204 (2588, 164, 1161, 1173);
  and ginst205 (2589, 161, 1161, 1173);
  nand ginst206 (2590, 1475, 140);
  and ginst207 (2591, 185, 1185, 1197);
  and ginst208 (2592, 158, 1185, 1197);
  and ginst209 (2593, 152, 1185, 1197);
  and ginst210 (2594, 146, 1185, 1197);
  and ginst211 (2595, 170, 1223, 1235);
  and ginst212 (2596, 173, 1223, 1235);
  and ginst213 (2597, 167, 1223, 1235);
  and ginst214 (2598, 164, 1223, 1235);
  and ginst215 (2599, 161, 1223, 1235);
  and ginst216 (2600, 185, 1247, 1259);
  and ginst217 (2601, 158, 1247, 1259);
  and ginst218 (2602, 152, 1247, 1259);
  and ginst219 (2603, 146, 1247, 1259);
  and ginst220 (2604, 106, 1731, 1743);
  and ginst221 (2605, 61, 1327, 1339);
  and ginst222 (2606, 106, 1697, 1709);
  and ginst223 (2607, 49, 1697, 1709);
  and ginst224 (2608, 103, 1697, 1709);
  and ginst225 (2609, 40, 1697, 1709);
  and ginst226 (2610, 37, 1697, 1709);
  and ginst227 (2611, 20, 1327, 1339);
  and ginst228 (2612, 17, 1327, 1339);
  and ginst229 (2613, 70, 1327, 1339);
  and ginst230 (2614, 64, 1327, 1339);
  and ginst231 (2615, 49, 1731, 1743);
  and ginst232 (2616, 103, 1731, 1743);
  and ginst233 (2617, 40, 1731, 1743);
  and ginst234 (2618, 37, 1731, 1743);
  and ginst235 (2619, 20, 1351, 1363);
  and ginst236 (2620, 17, 1351, 1363);
  and ginst237 (2621, 70, 1351, 1363);
  and ginst238 (2622, 64, 1351, 1363);
  not ginst239 (2623, 1475);
  and ginst240 (2624, 123, 1758, 599);
  and ginst241 (2625, 1777, 1785);
  and ginst242 (2626, 61, 1351, 1363);
  and ginst243 (2627, 1761, 1769);
  not ginst244 (2628, 1824);
  not ginst245 (2629, 1827);
  not ginst246 (2630, 1830);
  not ginst247 (2631, 1833);
  not ginst248 (2632, 1836);
  not ginst249 (2633, 1839);
  not ginst250 (2634, 1842);
  not ginst251 (2635, 1845);
  not ginst252 (2636, 1848);
  not ginst253 (2637, 1851);
  not ginst254 (2638, 1854);
  not ginst255 (2639, 1857);
  not ginst256 (2640, 1860);
  not ginst257 (2641, 1863);
  not ginst258 (2642, 1866);
  not ginst259 (2643, 1869);
  not ginst260 (2644, 1872);
  not ginst261 (2645, 1875);
  not ginst262 (2646, 1878);
  buf ginst263 (2647, 1209);
  not ginst264 (2653, 1161);
  not ginst265 (2664, 1173);
  buf ginst266 (2675, 1209);
  not ginst267 (2681, 1185);
  not ginst268 (2692, 1197);
  and ginst269 (2703, 179, 1185, 1197);
  buf ginst270 (2704, 1479);
  not ginst271 (2709, 1881);
  not ginst272 (2710, 1884);
  not ginst273 (2711, 1887);
  not ginst274 (2712, 1890);
  not ginst275 (2713, 1893);
  not ginst276 (2714, 1896);
  not ginst277 (2715, 1899);
  not ginst278 (2716, 1902);
  not ginst279 (2717, 1905);
  not ginst280 (2718, 1908);
  not ginst281 (2719, 1911);
  not ginst282 (2720, 1914);
  not ginst283 (2721, 1917);
  buf ginst284 (2722, 1213);
  not ginst285 (2728, 1223);
  not ginst286 (2739, 1235);
  buf ginst287 (2750, 1213);
  not ginst288 (2756, 1247);
  not ginst289 (2767, 1259);
  and ginst290 (2778, 179, 1247, 1259);
  not ginst291 (2779, 1327);
  not ginst292 (2790, 1339);
  not ginst293 (2801, 1351);
  not ginst294 (2812, 1363);
  not ginst295 (2823, 1375);
  not ginst296 (2824, 1378);
  not ginst297 (2825, 1381);
  not ginst298 (2826, 1384);
  not ginst299 (2827, 1387);
  not ginst300 (2828, 1390);
  not ginst301 (2829, 1393);
  not ginst302 (2830, 1396);
  and ginst303 (2831, 1104, 457, 1378);
  and ginst304 (2832, 1104, 468, 1384);
  and ginst305 (2833, 1104, 422, 1390);
  and ginst306 (2834, 1104, 435, 1396);
  and ginst307 (2835, 1067, 1375);
  and ginst308 (2836, 1067, 1381);
  and ginst309 (2837, 1067, 1387);
  and ginst310 (2838, 1067, 1393);
  not ginst311 (2839, 1415);
  not ginst312 (2840, 1418);
  not ginst313 (2841, 1421);
  not ginst314 (2842, 1424);
  not ginst315 (2843, 1427);
  not ginst316 (2844, 1430);
  not ginst317 (2845, 1433);
  not ginst318 (2846, 1436);
  and ginst319 (2847, 1104, 389, 1418);
  and ginst320 (2848, 1104, 400, 1424);
  and ginst321 (2849, 1104, 411, 1430);
  and ginst322 (2850, 1104, 374, 1436);
  and ginst323 (2851, 1067, 1415);
  and ginst324 (2852, 1067, 1421);
  and ginst325 (2853, 1067, 1427);
  and ginst326 (2854, 1067, 1433);
  not ginst327 (2855, 1455);
  not ginst328 (2861, 1462);
  and ginst329 (2867, 292, 1455);
  and ginst330 (2868, 288, 1455);
  and ginst331 (2869, 280, 1455);
  and ginst332 (2870, 272, 1455);
  and ginst333 (2871, 264, 1455);
  and ginst334 (2872, 241, 1462);
  and ginst335 (2873, 233, 1462);
  and ginst336 (2874, 225, 1462);
  and ginst337 (2875, 217, 1462);
  and ginst338 (2876, 209, 1462);
  buf ginst339 (2877, 1216);
  not ginst340 (2882, 1482);
  not ginst341 (2891, 1475);
  not ginst342 (2901, 1492);
  not ginst343 (2902, 1495);
  not ginst344 (2903, 1498);
  not ginst345 (2904, 1501);
  not ginst346 (2905, 1504);
  not ginst347 (2906, 1507);
  and ginst348 (2907, 1303, 1495);
  and ginst349 (2908, 1303, 479, 1501);
  and ginst350 (2909, 1303, 490, 1507);
  and ginst351 (2910, 1663, 1492);
  and ginst352 (2911, 1663, 1498);
  and ginst353 (2912, 1663, 1504);
  not ginst354 (2913, 1510);
  not ginst355 (2914, 1513);
  not ginst356 (2915, 1516);
  not ginst357 (2916, 1519);
  not ginst358 (2917, 1522);
  not ginst359 (2918, 1525);
  and ginst360 (2919, 1104, 503, 1513);
  not ginst361 (2920, 2349);
  and ginst362 (2921, 1104, 523, 1519);
  and ginst363 (2922, 1104, 534, 1525);
  and ginst364 (2923, 1067, 1510);
  and ginst365 (2924, 1067, 1516);
  and ginst366 (2925, 1067, 1522);
  not ginst367 (2926, 1542);
  not ginst368 (2927, 1545);
  not ginst369 (2928, 1548);
  not ginst370 (2929, 1551);
  not ginst371 (2930, 1554);
  not ginst372 (2931, 1557);
  not ginst373 (2932, 1560);
  not ginst374 (2933, 1563);
  and ginst375 (2934, 1303, 389, 1545);
  and ginst376 (2935, 1303, 400, 1551);
  and ginst377 (2936, 1303, 411, 1557);
  and ginst378 (2937, 1303, 374, 1563);
  and ginst379 (2938, 1663, 1542);
  and ginst380 (2939, 1663, 1548);
  and ginst381 (2940, 1663, 1554);
  and ginst382 (2941, 1663, 1560);
  not ginst383 (2942, 1566);
  not ginst384 (2948, 1573);
  and ginst385 (2954, 372, 1566);
  and ginst386 (2955, 366, 1566);
  and ginst387 (2956, 358, 1566);
  and ginst388 (2957, 348, 1566);
  and ginst389 (2958, 338, 1566);
  and ginst390 (2959, 331, 1573);
  and ginst391 (2960, 323, 1573);
  and ginst392 (2961, 315, 1573);
  and ginst393 (2962, 307, 1573);
  and ginst394 (2963, 299, 1573);
  not ginst395 (2964, 1588);
  and ginst396 (2969, 83, 1588);
  and ginst397 (2970, 86, 1588);
  and ginst398 (2971, 88, 1588);
  and ginst399 (2972, 88, 1588);
  not ginst400 (2973, 1594);
  not ginst401 (2974, 1597);
  not ginst402 (2975, 1600);
  not ginst403 (2976, 1603);
  not ginst404 (2977, 1606);
  not ginst405 (2978, 1609);
  and ginst406 (2979, 1315, 503, 1597);
  and ginst407 (2980, 1315, 514);
  and ginst408 (2981, 1315, 523, 1603);
  and ginst409 (2982, 1315, 534, 1609);
  and ginst410 (2983, 1675, 1594);
  or ginst411 (2984, 1675, 514);
  and ginst412 (2985, 1675, 1600);
  and ginst413 (2986, 1675, 1606);
  not ginst414 (2987, 1612);
  not ginst415 (2988, 1615);
  not ginst416 (2989, 1618);
  not ginst417 (2990, 1621);
  not ginst418 (2991, 1624);
  not ginst419 (2992, 1627);
  and ginst420 (2993, 1315, 1615);
  and ginst421 (2994, 1315, 479, 1621);
  and ginst422 (2995, 1315, 490, 1627);
  and ginst423 (2996, 1675, 1612);
  and ginst424 (2997, 1675, 1618);
  and ginst425 (2998, 1675, 1624);
  not ginst426 (2999, 1630);
  buf ginst427 (3000, 1469);
  buf ginst428 (3003, 1469);
  not ginst429 (3006, 1633);
  buf ginst430 (3007, 1469);
  buf ginst431 (3010, 1469);
  and ginst432 (3013, 1315, 1630);
  and ginst433 (3014, 1315, 1633);
  not ginst434 (3015, 1636);
  not ginst435 (3016, 1639);
  not ginst436 (3017, 1642);
  not ginst437 (3018, 1645);
  not ginst438 (3019, 1648);
  not ginst439 (3020, 1651);
  not ginst440 (3021, 1654);
  not ginst441 (3022, 1657);
  and ginst442 (3023, 1303, 457, 1639);
  and ginst443 (3024, 1303, 468, 1645);
  and ginst444 (3025, 1303, 422, 1651);
  and ginst445 (3026, 1303, 435, 1657);
  and ginst446 (3027, 1663, 1636);
  and ginst447 (3028, 1663, 1642);
  and ginst448 (3029, 1663, 1648);
  and ginst449 (3030, 1663, 1654);
  not ginst450 (3031, 1920);
  not ginst451 (3032, 1923);
  not ginst452 (3033, 1926);
  not ginst453 (3034, 1929);
  buf ginst454 (3035, 1660);
  buf ginst455 (3038, 1660);
  not ginst456 (3041, 1697);
  not ginst457 (3052, 1709);
  not ginst458 (3063, 1721);
  not ginst459 (3068, 1727);
  and ginst460 (3071, 97, 1721);
  and ginst461 (3072, 94, 1721);
  and ginst462 (3073, 97, 1721);
  and ginst463 (3074, 94, 1721);
  not ginst464 (3075, 1731);
  not ginst465 (3086, 1743);
  not ginst466 (3097, 1761);
  not ginst467 (3108, 1769);
  not ginst468 (3119, 1777);
  not ginst469 (3130, 1785);
  not ginst470 (3141, 1944);
  not ginst471 (3142, 1947);
  not ginst472 (3143, 1950);
  not ginst473 (3144, 1953);
  not ginst474 (3145, 1956);
  not ginst475 (3146, 1959);
  not ginst476 (3147, 1793);
  not ginst477 (3158, 1800);
  not ginst478 (3169, 1807);
  not ginst479 (3180, 1814);
  buf ginst480 (3191, 1821);
  not ginst481 (3194, 1932);
  not ginst482 (3195, 1935);
  not ginst483 (3196, 1938);
  not ginst484 (3197, 1941);
  not ginst485 (3198, 1962);
  not ginst486 (3199, 1965);
  buf ginst487 (3200, 1469);
  not ginst488 (3203, 1968);
  buf ginst489 (3357, 2704);
  buf ginst490 (3358, 2704);
  buf ginst491 (3359, 2704);
  buf ginst492 (3360, 2704);
  and ginst493 (3401, 457, 1092, 2824);
  and ginst494 (3402, 468, 1092, 2826);
  and ginst495 (3403, 422, 1092, 2828);
  and ginst496 (3404, 435, 1092, 2830);
  and ginst497 (3405, 1080, 2823);
  and ginst498 (3406, 1080, 2825);
  and ginst499 (3407, 1080, 2827);
  and ginst500 (3408, 1080, 2829);
  and ginst501 (3409, 389, 1092, 2840);
  and ginst502 (3410, 400, 1092, 2842);
  and ginst503 (3411, 411, 1092, 2844);
  and ginst504 (3412, 374, 1092, 2846);
  and ginst505 (3413, 1080, 2839);
  and ginst506 (3414, 1080, 2841);
  and ginst507 (3415, 1080, 2843);
  and ginst508 (3416, 1080, 2845);
  and ginst509 (3444, 1280, 2902);
  and ginst510 (3445, 479, 1280, 2904);
  and ginst511 (3446, 490, 1280, 2906);
  and ginst512 (3447, 1685, 2901);
  and ginst513 (3448, 1685, 2903);
  and ginst514 (3449, 1685, 2905);
  and ginst515 (3450, 503, 1092, 2914);
  and ginst516 (3451, 523, 1092, 2916);
  and ginst517 (3452, 534, 1092, 2918);
  and ginst518 (3453, 1080, 2913);
  and ginst519 (3454, 1080, 2915);
  and ginst520 (3455, 1080, 2917);
  and ginst521 (3456, 2920, 2350);
  and ginst522 (3459, 389, 1280, 2927);
  and ginst523 (3460, 400, 1280, 2929);
  and ginst524 (3461, 411, 1280, 2931);
  and ginst525 (3462, 374, 1280, 2933);
  and ginst526 (3463, 1685, 2926);
  and ginst527 (3464, 1685, 2928);
  and ginst528 (3465, 1685, 2930);
  and ginst529 (3466, 1685, 2932);
  and ginst530 (3481, 503, 1292, 2974);
  not ginst531 (3482, 2980);
  and ginst532 (3483, 523, 1292, 2976);
  and ginst533 (3484, 534, 1292, 2978);
  and ginst534 (3485, 1271, 2973);
  and ginst535 (3486, 1271, 2975);
  and ginst536 (3487, 1271, 2977);
  and ginst537 (3488, 1292, 2988);
  and ginst538 (3489, 479, 1292, 2990);
  and ginst539 (3490, 490, 1292, 2992);
  and ginst540 (3491, 1271, 2987);
  and ginst541 (3492, 1271, 2989);
  and ginst542 (3493, 1271, 2991);
  and ginst543 (3502, 1292, 2999);
  and ginst544 (3503, 1292, 3006);
  and ginst545 (3504, 457, 1280, 3016);
  and ginst546 (3505, 468, 1280, 3018);
  and ginst547 (3506, 422, 1280, 3020);
  and ginst548 (3507, 435, 1280, 3022);
  and ginst549 (3508, 1685, 3015);
  and ginst550 (3509, 1685, 3017);
  and ginst551 (3510, 1685, 3019);
  and ginst552 (3511, 1685, 3021);
  nand ginst553 (3512, 1923, 3031);
  nand ginst554 (3513, 1920, 3032);
  nand ginst555 (3514, 1929, 3033);
  nand ginst556 (3515, 1926, 3034);
  nand ginst557 (3558, 1947, 3141);
  nand ginst558 (3559, 1944, 3142);
  nand ginst559 (3560, 1953, 3143);
  nand ginst560 (3561, 1950, 3144);
  nand ginst561 (3562, 1959, 3145);
  nand ginst562 (3563, 1956, 3146);
  buf ginst563 (3604, 3191);
  nand ginst564 (3605, 1935, 3194);
  nand ginst565 (3606, 1932, 3195);
  nand ginst566 (3607, 1941, 3196);
  nand ginst567 (3608, 1938, 3197);
  nand ginst568 (3609, 1965, 3198);
  nand ginst569 (3610, 1962, 3199);
  not ginst570 (3613, 3191);
  and ginst571 (3614, 2882, 2891);
  and ginst572 (3615, 1482, 2891);
  and ginst573 (3616, 200, 2653, 1173);
  and ginst574 (3617, 203, 2653, 1173);
  and ginst575 (3618, 197, 2653, 1173);
  and ginst576 (3619, 194, 2653, 1173);
  and ginst577 (3620, 191, 2653, 1173);
  and ginst578 (3621, 182, 2681, 1197);
  and ginst579 (3622, 188, 2681, 1197);
  and ginst580 (3623, 155, 2681, 1197);
  and ginst581 (3624, 149, 2681, 1197);
  and ginst582 (3625, 2882, 2891);
  and ginst583 (3626, 1482, 2891);
  and ginst584 (3627, 200, 2728, 1235);
  and ginst585 (3628, 203, 2728, 1235);
  and ginst586 (3629, 197, 2728, 1235);
  and ginst587 (3630, 194, 2728, 1235);
  and ginst588 (3631, 191, 2728, 1235);
  and ginst589 (3632, 182, 2756, 1259);
  and ginst590 (3633, 188, 2756, 1259);
  and ginst591 (3634, 155, 2756, 1259);
  and ginst592 (3635, 149, 2756, 1259);
  and ginst593 (3636, 2882, 2891);
  and ginst594 (3637, 1482, 2891);
  and ginst595 (3638, 109, 3075, 1743);
  and ginst596 (3639, 2882, 2891);
  and ginst597 (3640, 1482, 2891);
  and ginst598 (3641, 11, 2779, 1339);
  and ginst599 (3642, 109, 3041, 1709);
  and ginst600 (3643, 46, 3041, 1709);
  and ginst601 (3644, 100, 3041, 1709);
  and ginst602 (3645, 91, 3041, 1709);
  and ginst603 (3646, 43, 3041, 1709);
  and ginst604 (3647, 76, 2779, 1339);
  and ginst605 (3648, 73, 2779, 1339);
  and ginst606 (3649, 67, 2779, 1339);
  and ginst607 (3650, 14, 2779, 1339);
  and ginst608 (3651, 46, 3075, 1743);
  and ginst609 (3652, 100, 3075, 1743);
  and ginst610 (3653, 91, 3075, 1743);
  and ginst611 (3654, 43, 3075, 1743);
  and ginst612 (3655, 76, 2801, 1363);
  and ginst613 (3656, 73, 2801, 1363);
  and ginst614 (3657, 67, 2801, 1363);
  and ginst615 (3658, 14, 2801, 1363);
  and ginst616 (3659, 120, 3119, 1785);
  and ginst617 (3660, 11, 2801, 1363);
  and ginst618 (3661, 118, 3097, 1769);
  and ginst619 (3662, 176, 2681, 1197);
  and ginst620 (3663, 176, 2756, 1259);
  or ginst621 (3664, 2831, 3401);
  or ginst622 (3665, 2832, 3402);
  or ginst623 (3666, 2833, 3403);
  or ginst624 (3667, 2834, 3404);
  or ginst625 (3668, 2835, 3405, 457);
  or ginst626 (3669, 2836, 3406, 468);
  or ginst627 (3670, 2837, 3407, 422);
  or ginst628 (3671, 2838, 3408, 435);
  or ginst629 (3672, 2847, 3409);
  or ginst630 (3673, 2848, 3410);
  or ginst631 (3674, 2849, 3411);
  or ginst632 (3675, 2850, 3412);
  or ginst633 (3676, 2851, 3413, 389);
  or ginst634 (3677, 2852, 3414, 400);
  or ginst635 (3678, 2853, 3415, 411);
  or ginst636 (3679, 2854, 3416, 374);
  and ginst637 (3680, 289, 2855);
  and ginst638 (3681, 281, 2855);
  and ginst639 (3682, 273, 2855);
  and ginst640 (3683, 265, 2855);
  and ginst641 (3684, 257, 2855);
  and ginst642 (3685, 234, 2861);
  and ginst643 (3686, 226, 2861);
  and ginst644 (3687, 218, 2861);
  and ginst645 (3688, 210, 2861);
  and ginst646 (3689, 206, 2861);
  not ginst647 (3691, 2891);
  or ginst648 (3700, 2907, 3444);
  or ginst649 (3701, 2908, 3445);
  or ginst650 (3702, 2909, 3446);
  or ginst651 (3703, 2911, 3448, 479);
  or ginst652 (3704, 2912, 3449, 490);
  or ginst653 (3705, 2910, 3447);
  or ginst654 (3708, 2919, 3450);
  or ginst655 (3709, 2921, 3451);
  or ginst656 (3710, 2922, 3452);
  or ginst657 (3711, 2923, 3453, 503);
  or ginst658 (3712, 2924, 3454, 523);
  or ginst659 (3713, 2925, 3455, 534);
  or ginst660 (3715, 2934, 3459);
  or ginst661 (3716, 2935, 3460);
  or ginst662 (3717, 2936, 3461);
  or ginst663 (3718, 2937, 3462);
  or ginst664 (3719, 2938, 3463, 389);
  or ginst665 (3720, 2939, 3464, 400);
  or ginst666 (3721, 2940, 3465, 411);
  or ginst667 (3722, 2941, 3466, 374);
  and ginst668 (3723, 369, 2942);
  and ginst669 (3724, 361, 2942);
  and ginst670 (3725, 351, 2942);
  and ginst671 (3726, 341, 2942);
  and ginst672 (3727, 324, 2948);
  and ginst673 (3728, 316, 2948);
  and ginst674 (3729, 308, 2948);
  and ginst675 (3730, 302, 2948);
  and ginst676 (3731, 293, 2948);
  or ginst677 (3732, 2942, 2958);
  and ginst678 (3738, 83, 2964);
  and ginst679 (3739, 87, 2964);
  and ginst680 (3740, 34, 2964);
  and ginst681 (3741, 34, 2964);
  or ginst682 (3742, 2979, 3481);
  or ginst683 (3743, 2981, 3483);
  or ginst684 (3744, 2982, 3484);
  or ginst685 (3745, 2983, 3485, 503);
  or ginst686 (3746, 2985, 3486, 523);
  or ginst687 (3747, 2986, 3487, 534);
  or ginst688 (3748, 2993, 3488);
  or ginst689 (3749, 2994, 3489);
  or ginst690 (3750, 2995, 3490);
  or ginst691 (3751, 2997, 3492, 479);
  or ginst692 (3752, 2998, 3493, 490);
  not ginst693 (3753, 3000);
  not ginst694 (3754, 3003);
  not ginst695 (3755, 3007);
  not ginst696 (3756, 3010);
  or ginst697 (3757, 3013, 3502);
  and ginst698 (3758, 1315, 446, 3003);
  or ginst699 (3759, 3014, 3503);
  and ginst700 (3760, 1315, 446, 3010);
  and ginst701 (3761, 1675, 3000);
  and ginst702 (3762, 1675, 3007);
  or ginst703 (3763, 3023, 3504);
  or ginst704 (3764, 3024, 3505);
  or ginst705 (3765, 3025, 3506);
  or ginst706 (3766, 3026, 3507);
  or ginst707 (3767, 3027, 3508, 457);
  or ginst708 (3768, 3028, 3509, 468);
  or ginst709 (3769, 3029, 3510, 422);
  or ginst710 (3770, 3030, 3511, 435);
  nand ginst711 (3771, 3512, 3513);
  nand ginst712 (3775, 3514, 3515);
  not ginst713 (3779, 3035);
  not ginst714 (3780, 3038);
  and ginst715 (3781, 117, 3097, 1769);
  and ginst716 (3782, 126, 3097, 1769);
  and ginst717 (3783, 127, 3097, 1769);
  and ginst718 (3784, 128, 3097, 1769);
  and ginst719 (3785, 131, 3119, 1785);
  and ginst720 (3786, 129, 3119, 1785);
  and ginst721 (3787, 119, 3119, 1785);
  and ginst722 (3788, 130, 3119, 1785);
  nand ginst723 (3789, 3558, 3559);
  nand ginst724 (3793, 3560, 3561);
  nand ginst725 (3797, 3562, 3563);
  and ginst726 (3800, 122, 3147, 1800);
  and ginst727 (3801, 113, 3147, 1800);
  and ginst728 (3802, 53, 3147, 1800);
  and ginst729 (3803, 114, 3147, 1800);
  and ginst730 (3804, 115, 3147, 1800);
  and ginst731 (3805, 52, 3169, 1814);
  and ginst732 (3806, 112, 3169, 1814);
  and ginst733 (3807, 116, 3169, 1814);
  and ginst734 (3808, 121, 3169, 1814);
  and ginst735 (3809, 123, 3169, 1814);
  nand ginst736 (3810, 3607, 3608);
  nand ginst737 (3813, 3605, 3606);
  and ginst738 (3816, 3482, 2984);
  or ginst739 (3819, 2996, 3491);
  not ginst740 (3822, 3200);
  nand ginst741 (3823, 3200, 3203);
  nand ginst742 (3824, 3609, 3610);
  not ginst743 (3827, 3456);
  or ginst744 (3828, 3739, 2970);
  or ginst745 (3829, 3740, 2971);
  or ginst746 (3830, 3741, 2972);
  or ginst747 (3831, 3738, 2969);
  not ginst748 (3834, 3664);
  not ginst749 (3835, 3665);
  not ginst750 (3836, 3666);
  not ginst751 (3837, 3667);
  not ginst752 (3838, 3672);
  not ginst753 (3839, 3673);
  not ginst754 (3840, 3674);
  not ginst755 (3841, 3675);
  or ginst756 (3842, 3681, 2868);
  or ginst757 (3849, 3682, 2869);
  or ginst758 (3855, 3683, 2870);
  or ginst759 (3861, 3684, 2871);
  or ginst760 (3867, 3685, 2872);
  or ginst761 (3873, 3686, 2873);
  or ginst762 (3881, 3687, 2874);
  or ginst763 (3887, 3688, 2875);
  or ginst764 (3893, 3689, 2876);
  not ginst765 (3908, 3701);
  not ginst766 (3909, 3702);
  not ginst767 (3911, 3700);
  not ginst768 (3914, 3708);
  not ginst769 (3915, 3709);
  not ginst770 (3916, 3710);
  not ginst771 (3917, 3715);
  not ginst772 (3918, 3716);
  not ginst773 (3919, 3717);
  not ginst774 (3920, 3718);
  or ginst775 (3921, 3724, 2955);
  or ginst776 (3927, 3725, 2956);
  or ginst777 (3933, 3726, 2957);
  or ginst778 (3942, 3727, 2959);
  or ginst779 (3948, 3728, 2960);
  or ginst780 (3956, 3729, 2961);
  or ginst781 (3962, 3730, 2962);
  or ginst782 (3968, 3731, 2963);
  not ginst783 (3975, 3742);
  not ginst784 (3976, 3743);
  not ginst785 (3977, 3744);
  not ginst786 (3978, 3749);
  not ginst787 (3979, 3750);
  and ginst788 (3980, 446, 1292, 3754);
  and ginst789 (3981, 446, 1292, 3756);
  and ginst790 (3982, 1271, 3753);
  and ginst791 (3983, 1271, 3755);
  not ginst792 (3984, 3757);
  not ginst793 (3987, 3759);
  not ginst794 (3988, 3763);
  not ginst795 (3989, 3764);
  not ginst796 (3990, 3765);
  not ginst797 (3991, 3766);
  and ginst798 (3998, 3456, 3119, 3130);
  or ginst799 (4008, 3723, 2954);
  or ginst800 (4011, 3680, 2867);
  not ginst801 (4021, 3748);
  nand ginst802 (4024, 1968, 3822);
  not ginst803 (4027, 3705);
  and ginst804 (4031, 3828, 1583);
  and ginst805 (4032, 24, 2882, 3691);
  and ginst806 (4033, 25, 1482, 3691);
  and ginst807 (4034, 26, 2882, 3691);
  and ginst808 (4035, 81, 1482, 3691);
  and ginst809 (4036, 3829, 1583);
  and ginst810 (4037, 79, 2882, 3691);
  and ginst811 (4038, 23, 1482, 3691);
  and ginst812 (4039, 82, 2882, 3691);
  and ginst813 (4040, 80, 1482, 3691);
  and ginst814 (4041, 3830, 1583);
  and ginst815 (4042, 3831, 1583);
  and ginst816 (4067, 3732, 514);
  and ginst817 (4080, 514, 3732);
  and ginst818 (4088, 3834, 3668);
  and ginst819 (4091, 3835, 3669);
  and ginst820 (4094, 3836, 3670);
  and ginst821 (4097, 3837, 3671);
  and ginst822 (4100, 3838, 3676);
  and ginst823 (4103, 3839, 3677);
  and ginst824 (4106, 3840, 3678);
  and ginst825 (4109, 3841, 3679);
  and ginst826 (4144, 3908, 3703);
  and ginst827 (4147, 3909, 3704);
  buf ginst828 (4150, 3705);
  and ginst829 (4153, 3914, 3711);
  and ginst830 (4156, 3915, 3712);
  and ginst831 (4159, 3916, 3713);
  or ginst832 (4183, 3758, 3980);
  or ginst833 (4184, 3760, 3981);
  or ginst834 (4185, 3761, 3982, 446);
  or ginst835 (4186, 3762, 3983, 446);
  not ginst836 (4188, 3771);
  not ginst837 (4191, 3775);
  and ginst838 (4196, 3775, 3771, 3035);
  and ginst839 (4197, 3987, 3119, 3130);
  and ginst840 (4198, 3920, 3722);
  not ginst841 (4199, 3816);
  not ginst842 (4200, 3789);
  not ginst843 (4203, 3793);
  buf ginst844 (4206, 3797);
  buf ginst845 (4209, 3797);
  buf ginst846 (4212, 3732);
  buf ginst847 (4215, 3732);
  buf ginst848 (4219, 3732);
  not ginst849 (4223, 3810);
  not ginst850 (4224, 3813);
  and ginst851 (4225, 3918, 3720);
  and ginst852 (4228, 3919, 3721);
  and ginst853 (4231, 3991, 3770);
  and ginst854 (4234, 3917, 3719);
  and ginst855 (4237, 3989, 3768);
  and ginst856 (4240, 3990, 3769);
  and ginst857 (4243, 3988, 3767);
  and ginst858 (4246, 3976, 3746);
  and ginst859 (4249, 3977, 3747);
  and ginst860 (4252, 3975, 3745);
  and ginst861 (4255, 3978, 3751);
  and ginst862 (4258, 3979, 3752);
  not ginst863 (4263, 3819);
  nand ginst864 (4264, 4024, 3823);
  not ginst865 (4267, 3824);
  and ginst866 (4268, 446, 3893);
  not ginst867 (4269, 3911);
  not ginst868 (4270, 3984);
  and ginst869 (4271, 3893, 446);
  not ginst870 (4272, 4031);
  or ginst871 (4273, 4032, 4033, 3614, 3615);
  or ginst872 (4274, 4034, 4035, 3625, 3626);
  not ginst873 (4275, 4036);
  or ginst874 (4276, 4037, 4038, 3636, 3637);
  or ginst875 (4277, 4039, 4040, 3639, 3640);
  not ginst876 (4278, 4041);
  not ginst877 (4279, 4042);
  and ginst878 (4280, 3887, 457);
  and ginst879 (4284, 3881, 468);
  and ginst880 (4290, 422, 3873);
  and ginst881 (4297, 3867, 435);
  and ginst882 (4298, 3861, 389);
  and ginst883 (4301, 3855, 400);
  and ginst884 (4305, 3849, 411);
  and ginst885 (4310, 3842, 374);
  and ginst886 (4316, 457, 3887);
  and ginst887 (4320, 468, 3881);
  and ginst888 (4325, 422, 3873);
  and ginst889 (4331, 435, 3867);
  and ginst890 (4332, 389, 3861);
  and ginst891 (4336, 400, 3855);
  and ginst892 (4342, 411, 3849);
  and ginst893 (4349, 374, 3842);
  not ginst894 (4357, 3968);
  not ginst895 (4364, 3962);
  buf ginst896 (4375, 3962);
  and ginst897 (4379, 3956, 479);
  and ginst898 (4385, 490, 3948);
  and ginst899 (4392, 3942, 503);
  and ginst900 (4396, 3933, 523);
  and ginst901 (4400, 3927, 534);
  not ginst902 (4405, 3921);
  buf ginst903 (4412, 3921);
  not ginst904 (4418, 3968);
  not ginst905 (4425, 3962);
  buf ginst906 (4436, 3962);
  and ginst907 (4440, 479, 3956);
  and ginst908 (4445, 490, 3948);
  and ginst909 (4451, 503, 3942);
  and ginst910 (4456, 523, 3933);
  and ginst911 (4462, 534, 3927);
  buf ginst912 (4469, 3921);
  not ginst913 (4477, 3921);
  buf ginst914 (4512, 3968);
  not ginst915 (4515, 4183);
  not ginst916 (4516, 4184);
  not ginst917 (4521, 4008);
  not ginst918 (4523, 4011);
  not ginst919 (4524, 4198);
  not ginst920 (4532, 3984);
  and ginst921 (4547, 3911, 3169, 3180);
  buf ginst922 (4548, 3893);
  buf ginst923 (4551, 3887);
  buf ginst924 (4554, 3881);
  buf ginst925 (4557, 3873);
  buf ginst926 (4560, 3867);
  buf ginst927 (4563, 3861);
  buf ginst928 (4566, 3855);
  buf ginst929 (4569, 3849);
  buf ginst930 (4572, 3842);
  nor ginst931 (4575, 422, 3873);
  buf ginst932 (4578, 3893);
  buf ginst933 (4581, 3887);
  buf ginst934 (4584, 3881);
  buf ginst935 (4587, 3867);
  buf ginst936 (4590, 3861);
  buf ginst937 (4593, 3855);
  buf ginst938 (4596, 3849);
  buf ginst939 (4599, 3873);
  buf ginst940 (4602, 3842);
  nor ginst941 (4605, 422, 3873);
  nor ginst942 (4608, 374, 3842);
  buf ginst943 (4611, 3956);
  buf ginst944 (4614, 3948);
  buf ginst945 (4617, 3942);
  buf ginst946 (4621, 3933);
  buf ginst947 (4624, 3927);
  nor ginst948 (4627, 490, 3948);
  buf ginst949 (4630, 3956);
  buf ginst950 (4633, 3942);
  buf ginst951 (4637, 3933);
  buf ginst952 (4640, 3927);
  buf ginst953 (4643, 3948);
  nor ginst954 (4646, 490, 3948);
  buf ginst955 (4649, 3927);
  buf ginst956 (4652, 3933);
  buf ginst957 (4655, 3921);
  buf ginst958 (4658, 3942);
  buf ginst959 (4662, 3956);
  buf ginst960 (4665, 3948);
  buf ginst961 (4668, 3968);
  buf ginst962 (4671, 3962);
  buf ginst963 (4674, 3873);
  buf ginst964 (4677, 3867);
  buf ginst965 (4680, 3887);
  buf ginst966 (4683, 3881);
  buf ginst967 (4686, 3893);
  buf ginst968 (4689, 3849);
  buf ginst969 (4692, 3842);
  buf ginst970 (4695, 3861);
  buf ginst971 (4698, 3855);
  nand ginst972 (4701, 3813, 4223);
  nand ginst973 (4702, 3810, 4224);
  not ginst974 (4720, 4021);
  nand ginst975 (4721, 4021, 4263);
  not ginst976 (4724, 4147);
  not ginst977 (4725, 4144);
  not ginst978 (4726, 4159);
  not ginst979 (4727, 4156);
  not ginst980 (4728, 4153);
  not ginst981 (4729, 4097);
  not ginst982 (4730, 4094);
  not ginst983 (4731, 4091);
  not ginst984 (4732, 4088);
  not ginst985 (4733, 4109);
  not ginst986 (4734, 4106);
  not ginst987 (4735, 4103);
  not ginst988 (4736, 4100);
  and ginst989 (4737, 4273, 2877);
  and ginst990 (4738, 4274, 2877);
  and ginst991 (4739, 4276, 2877);
  and ginst992 (4740, 4277, 2877);
  and ginst993 (4741, 4150, 1758, 1755);
  not ginst994 (4855, 4212);
  nand ginst995 (4856, 4212, 2712);
  nand ginst996 (4908, 4215, 2718);
  not ginst997 (4909, 4215);
  and ginst998 (4939, 4515, 4185);
  and ginst999 (4942, 4516, 4186);
  not ginst1000 (4947, 4219);
  and ginst1001 (4953, 4188, 3775, 3779);
  and ginst1002 (4954, 3771, 4191, 3780);
  and ginst1003 (4955, 4191, 4188, 3038);
  and ginst1004 (4956, 4109, 3097, 3108);
  and ginst1005 (4957, 4106, 3097, 3108);
  and ginst1006 (4958, 4103, 3097, 3108);
  and ginst1007 (4959, 4100, 3097, 3108);
  and ginst1008 (4960, 4159, 3119, 3130);
  and ginst1009 (4961, 4156, 3119, 3130);
  not ginst1010 (4965, 4225);
  not ginst1011 (4966, 4228);
  not ginst1012 (4967, 4231);
  not ginst1013 (4968, 4234);
  not ginst1014 (4972, 4246);
  not ginst1015 (4973, 4249);
  not ginst1016 (4974, 4252);
  nand ginst1017 (4975, 4252, 4199);
  not ginst1018 (4976, 4206);
  not ginst1019 (4977, 4209);
  and ginst1020 (4978, 3793, 3789, 4206);
  and ginst1021 (4979, 4203, 4200, 4209);
  and ginst1022 (4980, 4097, 3147, 3158);
  and ginst1023 (4981, 4094, 3147, 3158);
  and ginst1024 (4982, 4091, 3147, 3158);
  and ginst1025 (4983, 4088, 3147, 3158);
  and ginst1026 (4984, 4153, 3169, 3180);
  and ginst1027 (4985, 4147, 3169, 3180);
  and ginst1028 (4986, 4144, 3169, 3180);
  and ginst1029 (4987, 4150, 3169, 3180);
  nand ginst1030 (5049, 4701, 4702);
  not ginst1031 (5052, 4237);
  not ginst1032 (5053, 4240);
  not ginst1033 (5054, 4243);
  not ginst1034 (5055, 4255);
  not ginst1035 (5056, 4258);
  nand ginst1036 (5057, 3819, 4720);
  not ginst1037 (5058, 4264);
  nand ginst1038 (5059, 4264, 4267);
  and ginst1039 (5060, 4724, 4725, 4269, 4027);
  and ginst1040 (5061, 4726, 4727, 3827, 4728);
  and ginst1041 (5062, 4729, 4730, 4731, 4732);
  and ginst1042 (5063, 4733, 4734, 4735, 4736);
  and ginst1043 (5065, 4357, 4375);
  and ginst1044 (5066, 4364, 4357, 4379);
  and ginst1045 (5067, 4418, 4436);
  and ginst1046 (5068, 4425, 4418, 4440);
  not ginst1047 (5069, 4548);
  nand ginst1048 (5070, 4548, 2628);
  not ginst1049 (5071, 4551);
  nand ginst1050 (5072, 4551, 2629);
  not ginst1051 (5073, 4554);
  nand ginst1052 (5074, 4554, 2630);
  not ginst1053 (5075, 4557);
  nand ginst1054 (5076, 4557, 2631);
  not ginst1055 (5077, 4560);
  nand ginst1056 (5078, 4560, 2632);
  not ginst1057 (5079, 4563);
  nand ginst1058 (5080, 4563, 2633);
  not ginst1059 (5081, 4566);
  nand ginst1060 (5082, 4566, 2634);
  not ginst1061 (5083, 4569);
  nand ginst1062 (5084, 4569, 2635);
  not ginst1063 (5085, 4572);
  nand ginst1064 (5086, 4572, 2636);
  not ginst1065 (5087, 4575);
  nand ginst1066 (5088, 4578, 2638);
  not ginst1067 (5089, 4578);
  nand ginst1068 (5090, 4581, 2639);
  not ginst1069 (5091, 4581);
  nand ginst1070 (5092, 4584, 2640);
  not ginst1071 (5093, 4584);
  nand ginst1072 (5094, 4587, 2641);
  not ginst1073 (5095, 4587);
  nand ginst1074 (5096, 4590, 2642);
  not ginst1075 (5097, 4590);
  nand ginst1076 (5098, 4593, 2643);
  not ginst1077 (5099, 4593);
  nand ginst1078 (5100, 4596, 2644);
  not ginst1079 (5101, 4596);
  nand ginst1080 (5102, 4599, 2645);
  not ginst1081 (5103, 4599);
  nand ginst1082 (5104, 4602, 2646);
  not ginst1083 (5105, 4602);
  not ginst1084 (5106, 4611);
  nand ginst1085 (5107, 4611, 2709);
  not ginst1086 (5108, 4614);
  nand ginst1087 (5109, 4614, 2710);
  not ginst1088 (5110, 4617);
  nand ginst1089 (5111, 4617, 2711);
  nand ginst1090 (5112, 1890, 4855);
  not ginst1091 (5113, 4621);
  nand ginst1092 (5114, 4621, 2713);
  not ginst1093 (5115, 4624);
  nand ginst1094 (5116, 4624, 2714);
  and ginst1095 (5117, 4364, 4379);
  and ginst1096 (5118, 4364, 4379);
  and ginst1097 (5119, 54, 4405);
  not ginst1098 (5120, 4627);
  nand ginst1099 (5121, 4630, 2716);
  not ginst1100 (5122, 4630);
  nand ginst1101 (5123, 4633, 2717);
  not ginst1102 (5124, 4633);
  nand ginst1103 (5125, 1908, 4909);
  nand ginst1104 (5126, 4637, 2719);
  not ginst1105 (5127, 4637);
  nand ginst1106 (5128, 4640, 2720);
  not ginst1107 (5129, 4640);
  nand ginst1108 (5130, 4643, 2721);
  not ginst1109 (5131, 4643);
  and ginst1110 (5132, 4425, 4440);
  and ginst1111 (5133, 4425, 4440);
  not ginst1112 (5135, 4649);
  not ginst1113 (5136, 4652);
  nand ginst1114 (5137, 4655, 4521);
  not ginst1115 (5138, 4655);
  not ginst1116 (5139, 4658);
  nand ginst1117 (5140, 4658, 4947);
  not ginst1118 (5141, 4674);
  not ginst1119 (5142, 4677);
  not ginst1120 (5143, 4680);
  not ginst1121 (5144, 4683);
  nand ginst1122 (5145, 4686, 4523);
  not ginst1123 (5146, 4686);
  nor ginst1124 (5147, 4953, 4196);
  nor ginst1125 (5148, 4954, 4955);
  not ginst1126 (5150, 4524);
  nand ginst1127 (5153, 4228, 4965);
  nand ginst1128 (5154, 4225, 4966);
  nand ginst1129 (5155, 4234, 4967);
  nand ginst1130 (5156, 4231, 4968);
  not ginst1131 (5157, 4532);
  nand ginst1132 (5160, 4249, 4972);
  nand ginst1133 (5161, 4246, 4973);
  nand ginst1134 (5162, 3816, 4974);
  and ginst1135 (5163, 4200, 3793, 4976);
  and ginst1136 (5164, 3789, 4203, 4977);
  and ginst1137 (5165, 4942, 3147, 3158);
  not ginst1138 (5166, 4512);
  buf ginst1139 (5169, 4290);
  not ginst1140 (5172, 4605);
  buf ginst1141 (5173, 4325);
  not ginst1142 (5176, 4608);
  buf ginst1143 (5177, 4349);
  buf ginst1144 (5180, 4405);
  buf ginst1145 (5183, 4357);
  buf ginst1146 (5186, 4357);
  buf ginst1147 (5189, 4364);
  buf ginst1148 (5192, 4364);
  buf ginst1149 (5195, 4385);
  not ginst1150 (5198, 4646);
  buf ginst1151 (5199, 4418);
  buf ginst1152 (5202, 4425);
  buf ginst1153 (5205, 4445);
  buf ginst1154 (5208, 4418);
  buf ginst1155 (5211, 4425);
  buf ginst1156 (5214, 4477);
  buf ginst1157 (5217, 4469);
  buf ginst1158 (5220, 4477);
  not ginst1159 (5223, 4662);
  not ginst1160 (5224, 4665);
  not ginst1161 (5225, 4668);
  not ginst1162 (5226, 4671);
  not ginst1163 (5227, 4689);
  not ginst1164 (5228, 4692);
  not ginst1165 (5229, 4695);
  not ginst1166 (5230, 4698);
  nand ginst1167 (5232, 4240, 5052);
  nand ginst1168 (5233, 4237, 5053);
  nand ginst1169 (5234, 4258, 5055);
  nand ginst1170 (5235, 4255, 5056);
  nand ginst1171 (5236, 4721, 5057);
  nand ginst1172 (5239, 3824, 5058);
  and ginst1173 (5240, 5060, 5061, 4270);
  not ginst1174 (5241, 4939);
  nand ginst1175 (5242, 1824, 5069);
  nand ginst1176 (5243, 1827, 5071);
  nand ginst1177 (5244, 1830, 5073);
  nand ginst1178 (5245, 1833, 5075);
  nand ginst1179 (5246, 1836, 5077);
  nand ginst1180 (5247, 1839, 5079);
  nand ginst1181 (5248, 1842, 5081);
  nand ginst1182 (5249, 1845, 5083);
  nand ginst1183 (5250, 1848, 5085);
  nand ginst1184 (5252, 1854, 5089);
  nand ginst1185 (5253, 1857, 5091);
  nand ginst1186 (5254, 1860, 5093);
  nand ginst1187 (5255, 1863, 5095);
  nand ginst1188 (5256, 1866, 5097);
  nand ginst1189 (5257, 1869, 5099);
  nand ginst1190 (5258, 1872, 5101);
  nand ginst1191 (5259, 1875, 5103);
  nand ginst1192 (5260, 1878, 5105);
  nand ginst1193 (5261, 1881, 5106);
  nand ginst1194 (5262, 1884, 5108);
  nand ginst1195 (5263, 1887, 5110);
  nand ginst1196 (5264, 5112, 4856);
  nand ginst1197 (5274, 1893, 5113);
  nand ginst1198 (5275, 1896, 5115);
  nand ginst1199 (5282, 1902, 5122);
  nand ginst1200 (5283, 1905, 5124);
  nand ginst1201 (5284, 4908, 5125);
  nand ginst1202 (5298, 1911, 5127);
  nand ginst1203 (5299, 1914, 5129);
  nand ginst1204 (5300, 1917, 5131);
  nand ginst1205 (5303, 4652, 5135);
  nand ginst1206 (5304, 4649, 5136);
  nand ginst1207 (5305, 4008, 5138);
  nand ginst1208 (5306, 4219, 5139);
  nand ginst1209 (5307, 4677, 5141);
  nand ginst1210 (5308, 4674, 5142);
  nand ginst1211 (5309, 4683, 5143);
  nand ginst1212 (5310, 4680, 5144);
  nand ginst1213 (5311, 4011, 5146);
  not ginst1214 (5312, 5049);
  nand ginst1215 (5315, 5153, 5154);
  nand ginst1216 (5319, 5155, 5156);
  nand ginst1217 (5324, 5160, 5161);
  nand ginst1218 (5328, 5162, 4975);
  nor ginst1219 (5331, 5163, 4978);
  nor ginst1220 (5332, 5164, 4979);
  or ginst1221 (5346, 4412, 5119);
  nand ginst1222 (5363, 4665, 5223);
  nand ginst1223 (5364, 4662, 5224);
  nand ginst1224 (5365, 4671, 5225);
  nand ginst1225 (5366, 4668, 5226);
  nand ginst1226 (5367, 4692, 5227);
  nand ginst1227 (5368, 4689, 5228);
  nand ginst1228 (5369, 4698, 5229);
  nand ginst1229 (5370, 4695, 5230);
  nand ginst1230 (5371, 5148, 5147);
  buf ginst1231 (5374, 4939);
  nand ginst1232 (5377, 5232, 5233);
  nand ginst1233 (5382, 5234, 5235);
  nand ginst1234 (5385, 5239, 5059);
  and ginst1235 (5388, 5062, 5063, 5241);
  nand ginst1236 (5389, 5242, 5070);
  nand ginst1237 (5396, 5243, 5072);
  nand ginst1238 (5407, 5244, 5074);
  nand ginst1239 (5418, 5245, 5076);
  nand ginst1240 (5424, 5246, 5078);
  nand ginst1241 (5431, 5247, 5080);
  nand ginst1242 (5441, 5248, 5082);
  nand ginst1243 (5452, 5249, 5084);
  nand ginst1244 (5462, 5250, 5086);
  not ginst1245 (5469, 5169);
  nand ginst1246 (5470, 5088, 5252);
  nand ginst1247 (5477, 5090, 5253);
  nand ginst1248 (5488, 5092, 5254);
  nand ginst1249 (5498, 5094, 5255);
  nand ginst1250 (5506, 5096, 5256);
  nand ginst1251 (5520, 5098, 5257);
  nand ginst1252 (5536, 5100, 5258);
  nand ginst1253 (5549, 5102, 5259);
  nand ginst1254 (5555, 5104, 5260);
  nand ginst1255 (5562, 5261, 5107);
  nand ginst1256 (5573, 5262, 5109);
  nand ginst1257 (5579, 5263, 5111);
  nand ginst1258 (5595, 5274, 5114);
  nand ginst1259 (5606, 5275, 5116);
  nand ginst1260 (5616, 5180, 2715);
  not ginst1261 (5617, 5180);
  not ginst1262 (5618, 5183);
  not ginst1263 (5619, 5186);
  not ginst1264 (5620, 5189);
  not ginst1265 (5621, 5192);
  not ginst1266 (5622, 5195);
  nand ginst1267 (5624, 5121, 5282);
  nand ginst1268 (5634, 5123, 5283);
  nand ginst1269 (5655, 5126, 5298);
  nand ginst1270 (5671, 5128, 5299);
  nand ginst1271 (5684, 5130, 5300);
  not ginst1272 (5690, 5202);
  not ginst1273 (5691, 5211);
  nand ginst1274 (5692, 5303, 5304);
  nand ginst1275 (5696, 5137, 5305);
  nand ginst1276 (5700, 5306, 5140);
  nand ginst1277 (5703, 5307, 5308);
  nand ginst1278 (5707, 5309, 5310);
  nand ginst1279 (5711, 5145, 5311);
  and ginst1280 (5726, 5166, 4512);
  not ginst1281 (5727, 5173);
  not ginst1282 (5728, 5177);
  not ginst1283 (5730, 5199);
  not ginst1284 (5731, 5205);
  not ginst1285 (5732, 5208);
  not ginst1286 (5733, 5214);
  not ginst1287 (5734, 5217);
  not ginst1288 (5735, 5220);
  nand ginst1289 (5736, 5365, 5366);
  nand ginst1290 (5739, 5363, 5364);
  nand ginst1291 (5742, 5369, 5370);
  nand ginst1292 (5745, 5367, 5368);
  not ginst1293 (5755, 5236);
  nand ginst1294 (5756, 5332, 5331);
  and ginst1295 (5954, 5264, 4396);
  nand ginst1296 (5955, 1899, 5617);
  not ginst1297 (5956, 5346);
  and ginst1298 (6005, 5284, 4456);
  and ginst1299 (6006, 5284, 4456);
  not ginst1300 (6023, 5371);
  nand ginst1301 (6024, 5371, 5312);
  not ginst1302 (6025, 5315);
  not ginst1303 (6028, 5324);
  buf ginst1304 (6031, 5319);
  buf ginst1305 (6034, 5319);
  buf ginst1306 (6037, 5328);
  buf ginst1307 (6040, 5328);
  not ginst1308 (6044, 5385);
  or ginst1309 (6045, 5166, 5726);
  buf ginst1310 (6048, 5264);
  buf ginst1311 (6051, 5284);
  buf ginst1312 (6054, 5284);
  not ginst1313 (6065, 5374);
  nand ginst1314 (6066, 5374, 5054);
  not ginst1315 (6067, 5377);
  not ginst1316 (6068, 5382);
  nand ginst1317 (6069, 5382, 5755);
  and ginst1318 (6071, 5470, 4316);
  and ginst1319 (6072, 5477, 5470, 4320);
  and ginst1320 (6073, 5488, 5470, 4325, 5477);
  and ginst1321 (6074, 5562, 4357, 4385, 4364);
  and ginst1322 (6075, 5389, 4280);
  and ginst1323 (6076, 5396, 5389, 4284);
  and ginst1324 (6077, 5407, 5389, 4290, 5396);
  and ginst1325 (6078, 5624, 4418, 4445, 4425);
  not ginst1326 (6079, 5418);
  and ginst1327 (6080, 5396, 5418, 5407, 5389);
  and ginst1328 (6083, 5396, 4284);
  and ginst1329 (6084, 5407, 4290, 5396);
  and ginst1330 (6085, 5418, 5407, 5396);
  and ginst1331 (6086, 5396, 4284);
  and ginst1332 (6087, 4290, 5407, 5396);
  and ginst1333 (6088, 5407, 4290);
  and ginst1334 (6089, 5418, 5407);
  and ginst1335 (6090, 5407, 4290);
  and ginst1336 (6091, 5431, 5462, 5441, 5424, 5452);
  and ginst1337 (6094, 5424, 4298);
  and ginst1338 (6095, 5431, 5424, 4301);
  and ginst1339 (6096, 5441, 5424, 4305, 5431);
  and ginst1340 (6097, 5452, 5441, 5424, 4310, 5431);
  and ginst1341 (6098, 5431, 4301);
  and ginst1342 (6099, 5441, 4305, 5431);
  and ginst1343 (6100, 5452, 5441, 4310, 5431);
  and ginst1344 (6101, 4, 5462, 5441, 5452, 5431);
  and ginst1345 (6102, 4305, 5441);
  and ginst1346 (6103, 5452, 5441, 4310);
  and ginst1347 (6104, 4, 5462, 5441, 5452);
  and ginst1348 (6105, 5452, 4310);
  and ginst1349 (6106, 4, 5462, 5452);
  and ginst1350 (6107, 4, 5462);
  and ginst1351 (6108, 5549, 5488, 5477, 5470);
  and ginst1352 (6111, 5477, 4320);
  and ginst1353 (6112, 5488, 4325, 5477);
  and ginst1354 (6113, 5549, 5488, 5477);
  and ginst1355 (6114, 5477, 4320);
  and ginst1356 (6115, 5488, 4325, 5477);
  and ginst1357 (6116, 5488, 4325);
  and ginst1358 (6117, 5555, 5536, 5520, 5506, 5498);
  and ginst1359 (6120, 5498, 4332);
  and ginst1360 (6121, 5506, 5498, 4336);
  and ginst1361 (6122, 5520, 5498, 4342, 5506);
  and ginst1362 (6123, 5536, 5520, 5498, 4349, 5506);
  and ginst1363 (6124, 5506, 4336);
  and ginst1364 (6125, 5520, 4342, 5506);
  and ginst1365 (6126, 5536, 5520, 4349, 5506);
  and ginst1366 (6127, 5555, 5520, 5506, 5536);
  and ginst1367 (6128, 5506, 4336);
  and ginst1368 (6129, 5520, 4342, 5506);
  and ginst1369 (6130, 5536, 5520, 4349, 5506);
  and ginst1370 (6131, 5520, 4342);
  and ginst1371 (6132, 5536, 5520, 4349);
  and ginst1372 (6133, 5555, 5520, 5536);
  and ginst1373 (6134, 5520, 4342);
  and ginst1374 (6135, 5536, 5520, 4349);
  and ginst1375 (6136, 5536, 4349);
  and ginst1376 (6137, 5549, 5488);
  and ginst1377 (6138, 5555, 5536);
  not ginst1378 (6139, 5573);
  and ginst1379 (6140, 4364, 5573, 5562, 4357);
  and ginst1380 (6143, 5562, 4385, 4364);
  and ginst1381 (6144, 5573, 5562, 4364);
  and ginst1382 (6145, 4385, 5562, 4364);
  and ginst1383 (6146, 5562, 4385);
  and ginst1384 (6147, 5573, 5562);
  and ginst1385 (6148, 5562, 4385);
  and ginst1386 (6149, 5264, 4405, 5595, 5579, 5606);
  and ginst1387 (6152, 5579, 4067);
  and ginst1388 (6153, 5264, 5579, 4396);
  and ginst1389 (6154, 5595, 5579, 4400, 5264);
  and ginst1390 (6155, 5606, 5595, 5579, 4412, 5264);
  and ginst1391 (6156, 5595, 4400, 5264);
  and ginst1392 (6157, 5606, 5595, 4412, 5264);
  and ginst1393 (6158, 54, 4405, 5595, 5606, 5264);
  and ginst1394 (6159, 4400, 5595);
  and ginst1395 (6160, 5606, 5595, 4412);
  and ginst1396 (6161, 54, 4405, 5595, 5606);
  and ginst1397 (6162, 5606, 4412);
  and ginst1398 (6163, 54, 4405, 5606);
  nand ginst1399 (6164, 5616, 5955);
  and ginst1400 (6168, 5684, 5624, 4425, 4418);
  and ginst1401 (6171, 5624, 4445, 4425);
  and ginst1402 (6172, 5684, 5624, 4425);
  and ginst1403 (6173, 5624, 4445, 4425);
  and ginst1404 (6174, 5624, 4445);
  and ginst1405 (6175, 4477, 5671, 5655, 5284, 5634);
  and ginst1406 (6178, 5634, 4080);
  and ginst1407 (6179, 5284, 5634, 4456);
  and ginst1408 (6180, 5655, 5634, 4462, 5284);
  and ginst1409 (6181, 5671, 5655, 5634, 4469, 5284);
  and ginst1410 (6182, 5655, 4462, 5284);
  and ginst1411 (6183, 5671, 5655, 4469, 5284);
  and ginst1412 (6184, 4477, 5655, 5284, 5671);
  and ginst1413 (6185, 5655, 4462, 5284);
  and ginst1414 (6186, 5671, 5655, 4469, 5284);
  and ginst1415 (6187, 5655, 4462);
  and ginst1416 (6188, 5671, 5655, 4469);
  and ginst1417 (6189, 4477, 5655, 5671);
  and ginst1418 (6190, 5655, 4462);
  and ginst1419 (6191, 5671, 5655, 4469);
  and ginst1420 (6192, 5671, 4469);
  and ginst1421 (6193, 5684, 5624);
  and ginst1422 (6194, 4477, 5671);
  not ginst1423 (6197, 5692);
  not ginst1424 (6200, 5696);
  not ginst1425 (6203, 5703);
  not ginst1426 (6206, 5707);
  buf ginst1427 (6209, 5700);
  buf ginst1428 (6212, 5700);
  buf ginst1429 (6215, 5711);
  buf ginst1430 (6218, 5711);
  nand ginst1431 (6221, 5049, 6023);
  not ginst1432 (6234, 5756);
  nand ginst1433 (6235, 5756, 6044);
  buf ginst1434 (6238, 5462);
  buf ginst1435 (6241, 5389);
  buf ginst1436 (6244, 5389);
  buf ginst1437 (6247, 5396);
  buf ginst1438 (6250, 5396);
  buf ginst1439 (6253, 5407);
  buf ginst1440 (6256, 5407);
  buf ginst1441 (6259, 5424);
  buf ginst1442 (6262, 5431);
  buf ginst1443 (6265, 5441);
  buf ginst1444 (6268, 5452);
  buf ginst1445 (6271, 5549);
  buf ginst1446 (6274, 5488);
  buf ginst1447 (6277, 5470);
  buf ginst1448 (6280, 5477);
  buf ginst1449 (6283, 5549);
  buf ginst1450 (6286, 5488);
  buf ginst1451 (6289, 5470);
  buf ginst1452 (6292, 5477);
  buf ginst1453 (6295, 5555);
  buf ginst1454 (6298, 5536);
  buf ginst1455 (6301, 5498);
  buf ginst1456 (6304, 5520);
  buf ginst1457 (6307, 5506);
  buf ginst1458 (6310, 5506);
  buf ginst1459 (6313, 5555);
  buf ginst1460 (6316, 5536);
  buf ginst1461 (6319, 5498);
  buf ginst1462 (6322, 5520);
  buf ginst1463 (6325, 5562);
  buf ginst1464 (6328, 5562);
  buf ginst1465 (6331, 5579);
  buf ginst1466 (6335, 5595);
  buf ginst1467 (6338, 5606);
  buf ginst1468 (6341, 5684);
  buf ginst1469 (6344, 5624);
  buf ginst1470 (6347, 5684);
  buf ginst1471 (6350, 5624);
  buf ginst1472 (6353, 5671);
  buf ginst1473 (6356, 5634);
  buf ginst1474 (6359, 5655);
  buf ginst1475 (6364, 5671);
  buf ginst1476 (6367, 5634);
  buf ginst1477 (6370, 5655);
  not ginst1478 (6373, 5736);
  not ginst1479 (6374, 5739);
  not ginst1480 (6375, 5742);
  not ginst1481 (6376, 5745);
  nand ginst1482 (6377, 4243, 6065);
  nand ginst1483 (6378, 5236, 6068);
  or ginst1484 (6382, 4268, 6071, 6072, 6073);
  or ginst1485 (6386, 3968, 5065, 5066, 6074);
  or ginst1486 (6388, 4271, 6075, 6076, 6077);
  or ginst1487 (6392, 3968, 5067, 5068, 6078);
  or ginst1488 (6397, 4297, 6094, 6095, 6096, 6097);
  or ginst1489 (6411, 4320, 6116);
  or ginst1490 (6415, 4331, 6120, 6121, 6122, 6123);
  or ginst1491 (6419, 4342, 6136);
  or ginst1492 (6427, 4392, 6152, 6153, 6154, 6155);
  not ginst1493 (6434, 6048);
  or ginst1494 (6437, 4440, 6174);
  or ginst1495 (6441, 4451, 6178, 6179, 6180, 6181);
  or ginst1496 (6445, 4462, 6192);
  not ginst1497 (6448, 6051);
  not ginst1498 (6449, 6054);
  nand ginst1499 (6466, 6221, 6024);
  not ginst1500 (6469, 6031);
  not ginst1501 (6470, 6034);
  not ginst1502 (6471, 6037);
  not ginst1503 (6472, 6040);
  and ginst1504 (6473, 5315, 4524, 6031);
  and ginst1505 (6474, 6025, 5150, 6034);
  and ginst1506 (6475, 5324, 4532, 6037);
  and ginst1507 (6476, 6028, 5157, 6040);
  nand ginst1508 (6477, 5385, 6234);
  nand ginst1509 (6478, 6045, 132);
  or ginst1510 (6482, 4280, 6083, 6084, 6085);
  nor ginst1511 (6486, 4280, 6086, 6087);
  or ginst1512 (6490, 4284, 6088, 6089);
  nor ginst1513 (6494, 4284, 6090);
  or ginst1514 (6500, 4298, 6098, 6099, 6100, 6101);
  or ginst1515 (6504, 4301, 6102, 6103, 6104);
  or ginst1516 (6508, 4305, 6105, 6106);
  or ginst1517 (6512, 4310, 6107);
  or ginst1518 (6516, 4316, 6111, 6112, 6113);
  nor ginst1519 (6526, 4316, 6114, 6115);
  or ginst1520 (6536, 4336, 6131, 6132, 6133);
  or ginst1521 (6539, 4332, 6124, 6125, 6126, 6127);
  nor ginst1522 (6553, 4336, 6134, 6135);
  nor ginst1523 (6556, 4332, 6128, 6129, 6130);
  or ginst1524 (6566, 4375, 5117, 6143, 6144);
  nor ginst1525 (6569, 4375, 5118, 6145);
  or ginst1526 (6572, 4379, 6146, 6147);
  nor ginst1527 (6575, 4379, 6148);
  or ginst1528 (6580, 4067, 5954, 6156, 6157, 6158);
  or ginst1529 (6584, 4396, 6159, 6160, 6161);
  or ginst1530 (6587, 4400, 6162, 6163);
  or ginst1531 (6592, 4436, 5132, 6171, 6172);
  nor ginst1532 (6599, 4436, 5133, 6173);
  or ginst1533 (6606, 4456, 6187, 6188, 6189);
  or ginst1534 (6609, 4080, 6005, 6182, 6183, 6184);
  nor ginst1535 (6619, 4456, 6190, 6191);
  nor ginst1536 (6622, 4080, 6006, 6185, 6186);
  nand ginst1537 (6630, 5739, 6373);
  nand ginst1538 (6631, 5736, 6374);
  nand ginst1539 (6632, 5745, 6375);
  nand ginst1540 (6633, 5742, 6376);
  nand ginst1541 (6634, 6377, 6066);
  nand ginst1542 (6637, 6069, 6378);
  not ginst1543 (6640, 6164);
  and ginst1544 (6641, 6108, 6117);
  and ginst1545 (6643, 6140, 6149);
  and ginst1546 (6646, 6168, 6175);
  and ginst1547 (6648, 6080, 6091);
  nand ginst1548 (6650, 6238, 2637);
  not ginst1549 (6651, 6238);
  not ginst1550 (6653, 6241);
  not ginst1551 (6655, 6244);
  not ginst1552 (6657, 6247);
  not ginst1553 (6659, 6250);
  nand ginst1554 (6660, 6253, 5087);
  not ginst1555 (6661, 6253);
  nand ginst1556 (6662, 6256, 5469);
  not ginst1557 (6663, 6256);
  and ginst1558 (6664, 6091, 4);
  not ginst1559 (6666, 6259);
  not ginst1560 (6668, 6262);
  not ginst1561 (6670, 6265);
  not ginst1562 (6672, 6268);
  not ginst1563 (6675, 6117);
  not ginst1564 (6680, 6280);
  not ginst1565 (6681, 6292);
  not ginst1566 (6682, 6307);
  not ginst1567 (6683, 6310);
  nand ginst1568 (6689, 6325, 5120);
  not ginst1569 (6690, 6325);
  nand ginst1570 (6691, 6328, 5622);
  not ginst1571 (6692, 6328);
  and ginst1572 (6693, 6149, 54);
  not ginst1573 (6695, 6331);
  not ginst1574 (6698, 6335);
  nand ginst1575 (6699, 6338, 5956);
  not ginst1576 (6700, 6338);
  not ginst1577 (6703, 6175);
  not ginst1578 (6708, 6209);
  not ginst1579 (6709, 6212);
  not ginst1580 (6710, 6215);
  not ginst1581 (6711, 6218);
  and ginst1582 (6712, 5696, 5692, 6209);
  and ginst1583 (6713, 6200, 6197, 6212);
  and ginst1584 (6714, 5707, 5703, 6215);
  and ginst1585 (6715, 6206, 6203, 6218);
  buf ginst1586 (6716, 6466);
  and ginst1587 (6718, 6164, 1777, 3130);
  and ginst1588 (6719, 5150, 5315, 6469);
  and ginst1589 (6720, 4524, 6025, 6470);
  and ginst1590 (6721, 5157, 5324, 6471);
  and ginst1591 (6722, 4532, 6028, 6472);
  nand ginst1592 (6724, 6477, 6235);
  not ginst1593 (6739, 6271);
  not ginst1594 (6740, 6274);
  not ginst1595 (6741, 6277);
  not ginst1596 (6744, 6283);
  not ginst1597 (6745, 6286);
  not ginst1598 (6746, 6289);
  not ginst1599 (6751, 6295);
  not ginst1600 (6752, 6298);
  not ginst1601 (6753, 6301);
  not ginst1602 (6754, 6304);
  not ginst1603 (6755, 6322);
  not ginst1604 (6760, 6313);
  not ginst1605 (6761, 6316);
  not ginst1606 (6762, 6319);
  not ginst1607 (6772, 6341);
  not ginst1608 (6773, 6344);
  not ginst1609 (6776, 6347);
  not ginst1610 (6777, 6350);
  not ginst1611 (6782, 6353);
  not ginst1612 (6783, 6356);
  not ginst1613 (6784, 6359);
  not ginst1614 (6785, 6370);
  not ginst1615 (6790, 6364);
  not ginst1616 (6791, 6367);
  nand ginst1617 (6792, 6630, 6631);
  nand ginst1618 (6795, 6632, 6633);
  and ginst1619 (6801, 6108, 6415);
  and ginst1620 (6802, 6427, 6140);
  and ginst1621 (6803, 6397, 6080);
  and ginst1622 (6804, 6168, 6441);
  not ginst1623 (6805, 6466);
  nand ginst1624 (6806, 1851, 6651);
  not ginst1625 (6807, 6482);
  nand ginst1626 (6808, 6482, 6653);
  not ginst1627 (6809, 6486);
  nand ginst1628 (6810, 6486, 6655);
  not ginst1629 (6811, 6490);
  nand ginst1630 (6812, 6490, 6657);
  not ginst1631 (6813, 6494);
  nand ginst1632 (6814, 6494, 6659);
  nand ginst1633 (6815, 4575, 6661);
  nand ginst1634 (6816, 5169, 6663);
  or ginst1635 (6817, 6397, 6664);
  not ginst1636 (6823, 6500);
  nand ginst1637 (6824, 6500, 6666);
  not ginst1638 (6825, 6504);
  nand ginst1639 (6826, 6504, 6668);
  not ginst1640 (6827, 6508);
  nand ginst1641 (6828, 6508, 6670);
  not ginst1642 (6829, 6512);
  nand ginst1643 (6830, 6512, 6672);
  not ginst1644 (6831, 6415);
  not ginst1645 (6834, 6566);
  nand ginst1646 (6835, 6566, 5618);
  not ginst1647 (6836, 6569);
  nand ginst1648 (6837, 6569, 5619);
  not ginst1649 (6838, 6572);
  nand ginst1650 (6839, 6572, 5620);
  not ginst1651 (6840, 6575);
  nand ginst1652 (6841, 6575, 5621);
  nand ginst1653 (6842, 4627, 6690);
  nand ginst1654 (6843, 5195, 6692);
  or ginst1655 (6844, 6427, 6693);
  not ginst1656 (6850, 6580);
  nand ginst1657 (6851, 6580, 6695);
  not ginst1658 (6852, 6584);
  nand ginst1659 (6853, 6584, 6434);
  not ginst1660 (6854, 6587);
  nand ginst1661 (6855, 6587, 6698);
  nand ginst1662 (6856, 5346, 6700);
  not ginst1663 (6857, 6441);
  and ginst1664 (6860, 6197, 5696, 6708);
  and ginst1665 (6861, 5692, 6200, 6709);
  and ginst1666 (6862, 6203, 5707, 6710);
  and ginst1667 (6863, 5703, 6206, 6711);
  or ginst1668 (6866, 4197, 6718, 3785);
  nor ginst1669 (6872, 6719, 6473);
  nor ginst1670 (6873, 6720, 6474);
  nor ginst1671 (6874, 6721, 6475);
  nor ginst1672 (6875, 6722, 6476);
  not ginst1673 (6876, 6637);
  buf ginst1674 (6877, 6724);
  and ginst1675 (6879, 6045, 6478);
  and ginst1676 (6880, 6478, 132);
  or ginst1677 (6881, 6411, 6137);
  not ginst1678 (6884, 6516);
  not ginst1679 (6885, 6411);
  not ginst1680 (6888, 6526);
  not ginst1681 (6889, 6536);
  nand ginst1682 (6890, 6536, 5176);
  or ginst1683 (6891, 6419, 6138);
  not ginst1684 (6894, 6539);
  not ginst1685 (6895, 6553);
  nand ginst1686 (6896, 6553, 5728);
  not ginst1687 (6897, 6419);
  not ginst1688 (6900, 6556);
  or ginst1689 (6901, 6437, 6193);
  not ginst1690 (6904, 6592);
  not ginst1691 (6905, 6437);
  not ginst1692 (6908, 6599);
  or ginst1693 (6909, 6445, 6194);
  not ginst1694 (6912, 6606);
  not ginst1695 (6913, 6609);
  not ginst1696 (6914, 6619);
  nand ginst1697 (6915, 6619, 5734);
  not ginst1698 (6916, 6445);
  not ginst1699 (6919, 6622);
  not ginst1700 (6922, 6634);
  nand ginst1701 (6923, 6634, 6067);
  or ginst1702 (6924, 6382, 6801);
  or ginst1703 (6925, 6386, 6802);
  or ginst1704 (6926, 6388, 6803);
  or ginst1705 (6927, 6392, 6804);
  not ginst1706 (6930, 6724);
  nand ginst1707 (6932, 6650, 6806);
  nand ginst1708 (6935, 6241, 6807);
  nand ginst1709 (6936, 6244, 6809);
  nand ginst1710 (6937, 6247, 6811);
  nand ginst1711 (6938, 6250, 6813);
  nand ginst1712 (6939, 6660, 6815);
  nand ginst1713 (6940, 6662, 6816);
  nand ginst1714 (6946, 6259, 6823);
  nand ginst1715 (6947, 6262, 6825);
  nand ginst1716 (6948, 6265, 6827);
  nand ginst1717 (6949, 6268, 6829);
  nand ginst1718 (6953, 5183, 6834);
  nand ginst1719 (6954, 5186, 6836);
  nand ginst1720 (6955, 5189, 6838);
  nand ginst1721 (6956, 5192, 6840);
  nand ginst1722 (6957, 6689, 6842);
  nand ginst1723 (6958, 6691, 6843);
  nand ginst1724 (6964, 6331, 6850);
  nand ginst1725 (6965, 6048, 6852);
  nand ginst1726 (6966, 6335, 6854);
  nand ginst1727 (6967, 6699, 6856);
  nor ginst1728 (6973, 6860, 6712);
  nor ginst1729 (6974, 6861, 6713);
  nor ginst1730 (6975, 6862, 6714);
  nor ginst1731 (6976, 6863, 6715);
  not ginst1732 (6977, 6792);
  not ginst1733 (6978, 6795);
  or ginst1734 (6979, 6879, 6880);
  nand ginst1735 (6987, 4608, 6889);
  nand ginst1736 (6990, 5177, 6895);
  nand ginst1737 (6999, 5217, 6914);
  nand ginst1738 (7002, 5377, 6922);
  nand ginst1739 (7003, 6873, 6872);
  nand ginst1740 (7006, 6875, 6874);
  and ginst1741 (7011, 6866, 2681, 2692);
  and ginst1742 (7012, 6866, 2756, 2767);
  and ginst1743 (7013, 6866, 2779, 2790);
  not ginst1744 (7015, 6866);
  and ginst1745 (7016, 6866, 2801, 2812);
  nand ginst1746 (7018, 6935, 6808);
  nand ginst1747 (7019, 6936, 6810);
  nand ginst1748 (7020, 6937, 6812);
  nand ginst1749 (7021, 6938, 6814);
  not ginst1750 (7022, 6939);
  not ginst1751 (7023, 6817);
  nand ginst1752 (7028, 6946, 6824);
  nand ginst1753 (7031, 6947, 6826);
  nand ginst1754 (7034, 6948, 6828);
  nand ginst1755 (7037, 6949, 6830);
  and ginst1756 (7040, 6817, 6079);
  and ginst1757 (7041, 6831, 6675);
  nand ginst1758 (7044, 6953, 6835);
  nand ginst1759 (7045, 6954, 6837);
  nand ginst1760 (7046, 6955, 6839);
  nand ginst1761 (7047, 6956, 6841);
  not ginst1762 (7048, 6957);
  not ginst1763 (7049, 6844);
  nand ginst1764 (7054, 6964, 6851);
  nand ginst1765 (7057, 6965, 6853);
  nand ginst1766 (7060, 6966, 6855);
  and ginst1767 (7064, 6844, 6139);
  and ginst1768 (7065, 6857, 6703);
  not ginst1769 (7072, 6881);
  nand ginst1770 (7073, 6881, 5172);
  not ginst1771 (7074, 6885);
  nand ginst1772 (7075, 6885, 5727);
  nand ginst1773 (7076, 6890, 6987);
  not ginst1774 (7079, 6891);
  nand ginst1775 (7080, 6896, 6990);
  not ginst1776 (7083, 6897);
  not ginst1777 (7084, 6901);
  nand ginst1778 (7085, 6901, 5198);
  not ginst1779 (7086, 6905);
  nand ginst1780 (7087, 6905, 5731);
  not ginst1781 (7088, 6909);
  nand ginst1782 (7089, 6909, 6912);
  buf ginst1783 (709, 141);
  nand ginst1784 (7090, 6915, 6999);
  not ginst1785 (7093, 6916);
  nand ginst1786 (7094, 6974, 6973);
  nand ginst1787 (7097, 6976, 6975);
  nand ginst1788 (7101, 7002, 6923);
  not ginst1789 (7105, 6932);
  not ginst1790 (7110, 6967);
  and ginst1791 (7114, 6979, 603, 1755);
  not ginst1792 (7115, 7019);
  not ginst1793 (7116, 7021);
  and ginst1794 (7125, 6817, 7018);
  and ginst1795 (7126, 6817, 7020);
  and ginst1796 (7127, 6817, 7022);
  not ginst1797 (7130, 7045);
  not ginst1798 (7131, 7047);
  and ginst1799 (7139, 6844, 7044);
  and ginst1800 (7140, 6844, 7046);
  and ginst1801 (7141, 6844, 7048);
  and ginst1802 (7146, 6932, 1761, 3108);
  and ginst1803 (7147, 6967, 1777, 3130);
  not ginst1804 (7149, 7003);
  not ginst1805 (7150, 7006);
  nand ginst1806 (7151, 7006, 6876);
  nand ginst1807 (7152, 4605, 7072);
  nand ginst1808 (7153, 5173, 7074);
  nand ginst1809 (7158, 4646, 7084);
  nand ginst1810 (7159, 5205, 7086);
  nand ginst1811 (7160, 6606, 7088);
  not ginst1812 (7166, 7037);
  not ginst1813 (7167, 7034);
  not ginst1814 (7168, 7031);
  not ginst1815 (7169, 7028);
  not ginst1816 (7170, 7060);
  not ginst1817 (7171, 7057);
  not ginst1818 (7172, 7054);
  and ginst1819 (7173, 7115, 7023);
  and ginst1820 (7174, 7116, 7023);
  and ginst1821 (7175, 6940, 7023);
  and ginst1822 (7176, 5418, 7023);
  not ginst1823 (7177, 7041);
  and ginst1824 (7178, 7130, 7049);
  and ginst1825 (7179, 7131, 7049);
  and ginst1826 (7180, 6958, 7049);
  and ginst1827 (7181, 5573, 7049);
  not ginst1828 (7182, 7065);
  not ginst1829 (7183, 7094);
  nand ginst1830 (7184, 7094, 6977);
  not ginst1831 (7185, 7097);
  nand ginst1832 (7186, 7097, 6978);
  and ginst1833 (7187, 7037, 1761, 3108);
  and ginst1834 (7188, 7034, 1761, 3108);
  and ginst1835 (7189, 7031, 1761, 3108);
  or ginst1836 (7190, 4956, 7146, 3781);
  and ginst1837 (7196, 7060, 1777, 3130);
  and ginst1838 (7197, 7057, 1777, 3130);
  or ginst1839 (7198, 4960, 7147, 3786);
  nand ginst1840 (7204, 7101, 7149);
  not ginst1841 (7205, 7101);
  nand ginst1842 (7206, 6637, 7150);
  and ginst1843 (7207, 7028, 1793, 3158);
  and ginst1844 (7208, 7054, 1807, 3180);
  nand ginst1845 (7209, 7073, 7152);
  nand ginst1846 (7212, 7075, 7153);
  not ginst1847 (7215, 7076);
  nand ginst1848 (7216, 7076, 7079);
  not ginst1849 (7217, 7080);
  nand ginst1850 (7218, 7080, 7083);
  nand ginst1851 (7219, 7085, 7158);
  nand ginst1852 (7222, 7087, 7159);
  nand ginst1853 (7225, 7089, 7160);
  not ginst1854 (7228, 7090);
  nand ginst1855 (7229, 7090, 7093);
  or ginst1856 (7236, 7173, 7125);
  or ginst1857 (7239, 7174, 7126);
  or ginst1858 (7242, 7175, 7127);
  or ginst1859 (7245, 7176, 7040);
  or ginst1860 (7250, 7178, 7139);
  or ginst1861 (7257, 7179, 7140);
  or ginst1862 (7260, 7180, 7141);
  or ginst1863 (7263, 7181, 7064);
  nand ginst1864 (7268, 6792, 7183);
  nand ginst1865 (7269, 6795, 7185);
  or ginst1866 (7270, 4957, 7187, 3782);
  or ginst1867 (7276, 4958, 7188, 3783);
  or ginst1868 (7282, 4959, 7189, 3784);
  or ginst1869 (7288, 4961, 7196, 3787);
  or ginst1870 (7294, 3998, 7197, 3788);
  nand ginst1871 (7300, 7003, 7205);
  nand ginst1872 (7301, 7206, 7151);
  or ginst1873 (7304, 4980, 7207, 3800);
  or ginst1874 (7310, 4984, 7208, 3805);
  nand ginst1875 (7320, 6891, 7215);
  nand ginst1876 (7321, 6897, 7217);
  nand ginst1877 (7328, 6916, 7228);
  and ginst1878 (7338, 7190, 1185, 2692);
  and ginst1879 (7339, 7198, 2681, 2692);
  and ginst1880 (7340, 7190, 1247, 2767);
  and ginst1881 (7341, 7198, 2756, 2767);
  and ginst1882 (7342, 7190, 1327, 2790);
  and ginst1883 (7349, 7198, 2779, 2790);
  and ginst1884 (7357, 7198, 2801, 2812);
  not ginst1885 (7363, 7198);
  and ginst1886 (7364, 7190, 1351, 2812);
  not ginst1887 (7365, 7190);
  nand ginst1888 (7394, 7268, 7184);
  nand ginst1889 (7397, 7269, 7186);
  nand ginst1890 (7402, 7204, 7300);
  not ginst1891 (7405, 7209);
  nand ginst1892 (7406, 7209, 6884);
  not ginst1893 (7407, 7212);
  nand ginst1894 (7408, 7212, 6888);
  nand ginst1895 (7409, 7320, 7216);
  nand ginst1896 (7412, 7321, 7218);
  not ginst1897 (7415, 7219);
  nand ginst1898 (7416, 7219, 6904);
  not ginst1899 (7417, 7222);
  nand ginst1900 (7418, 7222, 6908);
  not ginst1901 (7419, 7225);
  nand ginst1902 (7420, 7225, 6913);
  nand ginst1903 (7421, 7328, 7229);
  not ginst1904 (7424, 7245);
  not ginst1905 (7425, 7242);
  not ginst1906 (7426, 7239);
  not ginst1907 (7427, 7236);
  not ginst1908 (7428, 7263);
  not ginst1909 (7429, 7260);
  not ginst1910 (7430, 7257);
  not ginst1911 (7431, 7250);
  not ginst1912 (7432, 7250);
  and ginst1913 (7433, 7310, 2653, 2664);
  and ginst1914 (7434, 7304, 1161, 2664);
  or ginst1915 (7435, 7011, 7338, 3621, 2591);
  and ginst1916 (7436, 7270, 1185, 2692);
  and ginst1917 (7437, 7288, 2681, 2692);
  and ginst1918 (7438, 7276, 1185, 2692);
  and ginst1919 (7439, 7294, 2681, 2692);
  and ginst1920 (7440, 7282, 1185, 2692);
  and ginst1921 (7441, 7310, 2728, 2739);
  and ginst1922 (7442, 7304, 1223, 2739);
  or ginst1923 (7443, 7012, 7340, 3632, 2600);
  and ginst1924 (7444, 7270, 1247, 2767);
  and ginst1925 (7445, 7288, 2756, 2767);
  and ginst1926 (7446, 7276, 1247, 2767);
  and ginst1927 (7447, 7294, 2756, 2767);
  and ginst1928 (7448, 7282, 1247, 2767);
  or ginst1929 (7449, 7013, 7342, 3641, 2605);
  and ginst1930 (7450, 7310, 3041, 3052);
  and ginst1931 (7451, 7304, 1697, 3052);
  and ginst1932 (7452, 7294, 2779, 2790);
  and ginst1933 (7453, 7282, 1327, 2790);
  and ginst1934 (7454, 7288, 2779, 2790);
  and ginst1935 (7455, 7276, 1327, 2790);
  and ginst1936 (7456, 7270, 1327, 2790);
  and ginst1937 (7457, 7310, 3075, 3086);
  and ginst1938 (7458, 7304, 1731, 3086);
  and ginst1939 (7459, 7294, 2801, 2812);
  and ginst1940 (7460, 7282, 1351, 2812);
  and ginst1941 (7461, 7288, 2801, 2812);
  and ginst1942 (7462, 7276, 1351, 2812);
  and ginst1943 (7463, 7270, 1351, 2812);
  and ginst1944 (7464, 7250, 603, 599);
  not ginst1945 (7465, 7310);
  not ginst1946 (7466, 7294);
  not ginst1947 (7467, 7288);
  not ginst1948 (7468, 7301);
  or ginst1949 (7469, 7016, 7364, 3660, 2626);
  not ginst1950 (7470, 7304);
  not ginst1951 (7471, 7282);
  not ginst1952 (7472, 7276);
  not ginst1953 (7473, 7270);
  buf ginst1954 (7474, 7394);
  buf ginst1955 (7476, 7397);
  and ginst1956 (7479, 7301, 3068);
  and ginst1957 (7481, 7245, 1793, 3158);
  and ginst1958 (7482, 7242, 1793, 3158);
  and ginst1959 (7483, 7239, 1793, 3158);
  and ginst1960 (7484, 7236, 1793, 3158);
  and ginst1961 (7485, 7263, 1807, 3180);
  and ginst1962 (7486, 7260, 1807, 3180);
  and ginst1963 (7487, 7257, 1807, 3180);
  and ginst1964 (7488, 7250, 1807, 3180);
  nand ginst1965 (7489, 6979, 7250);
  nand ginst1966 (7492, 6516, 7405);
  nand ginst1967 (7493, 6526, 7407);
  nand ginst1968 (7498, 6592, 7415);
  nand ginst1969 (7499, 6599, 7417);
  nand ginst1970 (7500, 6609, 7419);
  and ginst1971 (7503, 7105, 7166, 7167, 7168, 7169, 7424, 7425, 7426, 7427);
  and ginst1972 (7504, 6640, 7110, 7170, 7171, 7172, 7428, 7429, 7430, 7431);
  or ginst1973 (7505, 7433, 7434, 3616, 2585);
  and ginst1974 (7506, 7435, 2675);
  or ginst1975 (7507, 7339, 7436, 3622, 2592);
  or ginst1976 (7508, 7437, 7438, 3623, 2593);
  or ginst1977 (7509, 7439, 7440, 3624, 2594);
  or ginst1978 (7510, 7441, 7442, 3627, 2595);
  and ginst1979 (7511, 7443, 2750);
  or ginst1980 (7512, 7341, 7444, 3633, 2601);
  or ginst1981 (7513, 7445, 7446, 3634, 2602);
  or ginst1982 (7514, 7447, 7448, 3635, 2603);
  or ginst1983 (7515, 7450, 7451, 3646, 2610);
  or ginst1984 (7516, 7452, 7453, 3647, 2611);
  or ginst1985 (7517, 7454, 7455, 3648, 2612);
  or ginst1986 (7518, 7349, 7456, 3649, 2613);
  or ginst1987 (7519, 7457, 7458, 3654, 2618);
  or ginst1988 (7520, 7459, 7460, 3655, 2619);
  or ginst1989 (7521, 7461, 7462, 3656, 2620);
  or ginst1990 (7522, 7357, 7463, 3657, 2621);
  or ginst1991 (7525, 4741, 7114, 2624, 7464);
  and ginst1992 (7526, 7468, 3119, 3130);
  not ginst1993 (7527, 7394);
  not ginst1994 (7528, 7397);
  not ginst1995 (7529, 7402);
  and ginst1996 (7530, 7402, 3068);
  or ginst1997 (7531, 4981, 7481, 3801);
  or ginst1998 (7537, 4982, 7482, 3802);
  or ginst1999 (7543, 4983, 7483, 3803);
  or ginst2000 (7549, 5165, 7484, 3804);
  or ginst2001 (7555, 4985, 7485, 3806);
  or ginst2002 (7561, 4986, 7486, 3807);
  or ginst2003 (7567, 4547, 7487, 3808);
  or ginst2004 (7573, 4987, 7488, 3809);
  nand ginst2005 (7579, 7492, 7406);
  nand ginst2006 (7582, 7493, 7408);
  not ginst2007 (7585, 7409);
  nand ginst2008 (7586, 7409, 6894);
  not ginst2009 (7587, 7412);
  nand ginst2010 (7588, 7412, 6900);
  nand ginst2011 (7589, 7498, 7416);
  nand ginst2012 (7592, 7499, 7418);
  nand ginst2013 (7595, 7500, 7420);
  not ginst2014 (7598, 7421);
  nand ginst2015 (7599, 7421, 6919);
  and ginst2016 (7600, 7505, 2647);
  and ginst2017 (7601, 7507, 2675);
  and ginst2018 (7602, 7508, 2675);
  and ginst2019 (7603, 7509, 2675);
  and ginst2020 (7604, 7510, 2722);
  and ginst2021 (7605, 7512, 2750);
  and ginst2022 (7606, 7513, 2750);
  and ginst2023 (7607, 7514, 2750);
  and ginst2024 (7624, 6979, 7489);
  and ginst2025 (7625, 7489, 7250);
  and ginst2026 (7626, 1149, 7525);
  and ginst2027 (7631, 562, 7527, 7528, 6805, 6930);
  and ginst2028 (7636, 7529, 3097, 3108);
  nand ginst2029 (7657, 6539, 7585);
  nand ginst2030 (7658, 6556, 7587);
  nand ginst2031 (7665, 6622, 7598);
  and ginst2032 (7666, 7555, 2653, 2664);
  and ginst2033 (7667, 7531, 1161, 2664);
  and ginst2034 (7668, 7561, 2653, 2664);
  and ginst2035 (7669, 7537, 1161, 2664);
  and ginst2036 (7670, 7567, 2653, 2664);
  and ginst2037 (7671, 7543, 1161, 2664);
  and ginst2038 (7672, 7573, 2653, 2664);
  and ginst2039 (7673, 7549, 1161, 2664);
  and ginst2040 (7674, 7555, 2728, 2739);
  and ginst2041 (7675, 7531, 1223, 2739);
  and ginst2042 (7676, 7561, 2728, 2739);
  and ginst2043 (7677, 7537, 1223, 2739);
  and ginst2044 (7678, 7567, 2728, 2739);
  and ginst2045 (7679, 7543, 1223, 2739);
  and ginst2046 (7680, 7573, 2728, 2739);
  and ginst2047 (7681, 7549, 1223, 2739);
  and ginst2048 (7682, 7573, 3075, 3086);
  and ginst2049 (7683, 7549, 1731, 3086);
  and ginst2050 (7684, 7573, 3041, 3052);
  and ginst2051 (7685, 7549, 1697, 3052);
  and ginst2052 (7686, 7567, 3041, 3052);
  and ginst2053 (7687, 7543, 1697, 3052);
  and ginst2054 (7688, 7561, 3041, 3052);
  and ginst2055 (7689, 7537, 1697, 3052);
  and ginst2056 (7690, 7555, 3041, 3052);
  and ginst2057 (7691, 7531, 1697, 3052);
  and ginst2058 (7692, 7567, 3075, 3086);
  and ginst2059 (7693, 7543, 1731, 3086);
  and ginst2060 (7694, 7561, 3075, 3086);
  and ginst2061 (7695, 7537, 1731, 3086);
  and ginst2062 (7696, 7555, 3075, 3086);
  and ginst2063 (7697, 7531, 1731, 3086);
  or ginst2064 (7698, 7624, 7625);
  not ginst2065 (7699, 7573);
  not ginst2066 (7700, 7567);
  not ginst2067 (7701, 7561);
  not ginst2068 (7702, 7555);
  and ginst2069 (7703, 1156, 7631, 245);
  not ginst2070 (7704, 7549);
  not ginst2071 (7705, 7543);
  not ginst2072 (7706, 7537);
  not ginst2073 (7707, 7531);
  not ginst2074 (7708, 7579);
  nand ginst2075 (7709, 7579, 6739);
  not ginst2076 (7710, 7582);
  nand ginst2077 (7711, 7582, 6744);
  nand ginst2078 (7712, 7657, 7586);
  nand ginst2079 (7715, 7658, 7588);
  not ginst2080 (7718, 7589);
  nand ginst2081 (7719, 7589, 6772);
  not ginst2082 (7720, 7592);
  nand ginst2083 (7721, 7592, 6776);
  not ginst2084 (7722, 7595);
  nand ginst2085 (7723, 7595, 5733);
  nand ginst2086 (7724, 7665, 7599);
  or ginst2087 (7727, 7666, 7667, 3617, 2586);
  or ginst2088 (7728, 7668, 7669, 3618, 2587);
  or ginst2089 (7729, 7670, 7671, 3619, 2588);
  or ginst2090 (7730, 7672, 7673, 3620, 2589);
  or ginst2091 (7731, 7674, 7675, 3628, 2596);
  or ginst2092 (7732, 7676, 7677, 3629, 2597);
  or ginst2093 (7733, 7678, 7679, 3630, 2598);
  or ginst2094 (7734, 7680, 7681, 3631, 2599);
  or ginst2095 (7735, 7682, 7683, 3638, 2604);
  or ginst2096 (7736, 7684, 7685, 3642, 2606);
  or ginst2097 (7737, 7686, 7687, 3643, 2607);
  or ginst2098 (7738, 7688, 7689, 3644, 2608);
  or ginst2099 (7739, 7690, 7691, 3645, 2609);
  or ginst2100 (7740, 7692, 7693, 3651, 2615);
  or ginst2101 (7741, 7694, 7695, 3652, 2616);
  or ginst2102 (7742, 7696, 7697, 3653, 2617);
  nand ginst2103 (7743, 6271, 7708);
  nand ginst2104 (7744, 6283, 7710);
  nand ginst2105 (7749, 6341, 7718);
  nand ginst2106 (7750, 6347, 7720);
  nand ginst2107 (7751, 5214, 7722);
  and ginst2108 (7754, 7727, 2647);
  and ginst2109 (7755, 7728, 2647);
  and ginst2110 (7756, 7729, 2647);
  and ginst2111 (7757, 7730, 2647);
  and ginst2112 (7758, 7731, 2722);
  and ginst2113 (7759, 7732, 2722);
  and ginst2114 (7760, 7733, 2722);
  and ginst2115 (7761, 7734, 2722);
  nand ginst2116 (7762, 7743, 7709);
  nand ginst2117 (7765, 7744, 7711);
  not ginst2118 (7768, 7712);
  nand ginst2119 (7769, 7712, 6751);
  not ginst2120 (7770, 7715);
  nand ginst2121 (7771, 7715, 6760);
  nand ginst2122 (7772, 7749, 7719);
  nand ginst2123 (7775, 7750, 7721);
  nand ginst2124 (7778, 7751, 7723);
  not ginst2125 (7781, 7724);
  nand ginst2126 (7782, 7724, 5735);
  nand ginst2127 (7787, 6295, 7768);
  nand ginst2128 (7788, 6313, 7770);
  nand ginst2129 (7795, 5220, 7781);
  not ginst2130 (7796, 7762);
  nand ginst2131 (7797, 7762, 6740);
  not ginst2132 (7798, 7765);
  nand ginst2133 (7799, 7765, 6745);
  nand ginst2134 (7800, 7787, 7769);
  nand ginst2135 (7803, 7788, 7771);
  not ginst2136 (7806, 7772);
  nand ginst2137 (7807, 7772, 6773);
  not ginst2138 (7808, 7775);
  nand ginst2139 (7809, 7775, 6777);
  not ginst2140 (7810, 7778);
  nand ginst2141 (7811, 7778, 6782);
  nand ginst2142 (7812, 7795, 7782);
  nand ginst2143 (7815, 6274, 7796);
  nand ginst2144 (7816, 6286, 7798);
  nand ginst2145 (7821, 6344, 7806);
  nand ginst2146 (7822, 6350, 7808);
  nand ginst2147 (7823, 6353, 7810);
  nand ginst2148 (7826, 7815, 7797);
  nand ginst2149 (7829, 7816, 7799);
  not ginst2150 (7832, 7800);
  nand ginst2151 (7833, 7800, 6752);
  not ginst2152 (7834, 7803);
  nand ginst2153 (7835, 7803, 6761);
  nand ginst2154 (7836, 7821, 7807);
  nand ginst2155 (7839, 7822, 7809);
  nand ginst2156 (7842, 7823, 7811);
  not ginst2157 (7845, 7812);
  nand ginst2158 (7846, 7812, 6790);
  nand ginst2159 (7851, 6298, 7832);
  nand ginst2160 (7852, 6316, 7834);
  nand ginst2161 (7859, 6364, 7845);
  not ginst2162 (7860, 7826);
  nand ginst2163 (7861, 7826, 6741);
  not ginst2164 (7862, 7829);
  nand ginst2165 (7863, 7829, 6746);
  nand ginst2166 (7864, 7851, 7833);
  nand ginst2167 (7867, 7852, 7835);
  not ginst2168 (7870, 7836);
  nand ginst2169 (7871, 7836, 5730);
  not ginst2170 (7872, 7839);
  nand ginst2171 (7873, 7839, 5732);
  not ginst2172 (7874, 7842);
  nand ginst2173 (7875, 7842, 6783);
  nand ginst2174 (7876, 7859, 7846);
  nand ginst2175 (7879, 6277, 7860);
  nand ginst2176 (7880, 6289, 7862);
  nand ginst2177 (7885, 5199, 7870);
  nand ginst2178 (7886, 5208, 7872);
  nand ginst2179 (7887, 6356, 7874);
  nand ginst2180 (7890, 7879, 7861);
  nand ginst2181 (7893, 7880, 7863);
  not ginst2182 (7896, 7864);
  nand ginst2183 (7897, 7864, 6753);
  not ginst2184 (7898, 7867);
  nand ginst2185 (7899, 7867, 6762);
  nand ginst2186 (7900, 7885, 7871);
  nand ginst2187 (7903, 7886, 7873);
  nand ginst2188 (7906, 7887, 7875);
  not ginst2189 (7909, 7876);
  nand ginst2190 (7910, 7876, 6791);
  nand ginst2191 (7917, 6301, 7896);
  nand ginst2192 (7918, 6319, 7898);
  nand ginst2193 (7923, 6367, 7909);
  not ginst2194 (7924, 7890);
  nand ginst2195 (7925, 7890, 6680);
  not ginst2196 (7926, 7893);
  nand ginst2197 (7927, 7893, 6681);
  not ginst2198 (7928, 7900);
  nand ginst2199 (7929, 7900, 5690);
  not ginst2200 (7930, 7903);
  nand ginst2201 (7931, 7903, 5691);
  nand ginst2202 (7932, 7917, 7897);
  nand ginst2203 (7935, 7918, 7899);
  not ginst2204 (7938, 7906);
  nand ginst2205 (7939, 7906, 6784);
  nand ginst2206 (7940, 7923, 7910);
  nand ginst2207 (7943, 6280, 7924);
  nand ginst2208 (7944, 6292, 7926);
  nand ginst2209 (7945, 5202, 7928);
  nand ginst2210 (7946, 5211, 7930);
  nand ginst2211 (7951, 6359, 7938);
  nand ginst2212 (7954, 7943, 7925);
  nand ginst2213 (7957, 7944, 7927);
  nand ginst2214 (7960, 7945, 7929);
  nand ginst2215 (7963, 7946, 7931);
  not ginst2216 (7966, 7932);
  nand ginst2217 (7967, 7932, 6754);
  not ginst2218 (7968, 7935);
  nand ginst2219 (7969, 7935, 6755);
  nand ginst2220 (7970, 7951, 7939);
  not ginst2221 (7973, 7940);
  nand ginst2222 (7974, 7940, 6785);
  nand ginst2223 (7984, 6304, 7966);
  nand ginst2224 (7985, 6322, 7968);
  nand ginst2225 (7987, 6370, 7973);
  and ginst2226 (7988, 7957, 6831, 1157);
  and ginst2227 (7989, 7954, 6415, 1157);
  and ginst2228 (7990, 7957, 7041, 566);
  and ginst2229 (7991, 7954, 7177, 566);
  not ginst2230 (7992, 7970);
  nand ginst2231 (7993, 7970, 6448);
  and ginst2232 (7994, 7963, 6857, 1219);
  and ginst2233 (7995, 7960, 6441, 1219);
  and ginst2234 (7996, 7963, 7065, 583);
  and ginst2235 (7997, 7960, 7182, 583);
  nand ginst2236 (7998, 7984, 7967);
  nand ginst2237 (8001, 7985, 7969);
  nand ginst2238 (8004, 7987, 7974);
  nand ginst2239 (8009, 6051, 7992);
  or ginst2240 (8013, 7988, 7989, 7990, 7991);
  or ginst2241 (8017, 7994, 7995, 7996, 7997);
  not ginst2242 (8020, 7998);
  nand ginst2243 (8021, 7998, 6682);
  not ginst2244 (8022, 8001);
  nand ginst2245 (8023, 8001, 6683);
  nand ginst2246 (8025, 8009, 7993);
  not ginst2247 (8026, 8004);
  nand ginst2248 (8027, 8004, 6449);
  nand ginst2249 (8031, 6307, 8020);
  nand ginst2250 (8032, 6310, 8022);
  not ginst2251 (8033, 8013);
  nand ginst2252 (8034, 6054, 8026);
  and ginst2253 (8035, 583, 8025);
  not ginst2254 (8036, 8017);
  nand ginst2255 (8037, 8031, 8021);
  nand ginst2256 (8038, 8032, 8023);
  nand ginst2257 (8039, 8034, 8027);
  not ginst2258 (8040, 8038);
  and ginst2259 (8041, 566, 8037);
  not ginst2260 (8042, 8039);
  and ginst2261 (8043, 8040, 1157);
  and ginst2262 (8044, 8042, 1219);
  or ginst2263 (8045, 8043, 8041);
  or ginst2264 (8048, 8044, 8035);
  nand ginst2265 (8055, 8045, 8033);
  not ginst2266 (8056, 8045);
  nand ginst2267 (8057, 8048, 8036);
  not ginst2268 (8058, 8048);
  nand ginst2269 (8059, 8013, 8056);
  nand ginst2270 (8060, 8017, 8058);
  nand ginst2271 (8061, 8055, 8059);
  nand ginst2272 (8064, 8057, 8060);
  and ginst2273 (8071, 8064, 1777, 3130);
  and ginst2274 (8072, 8061, 1761, 3108);
  not ginst2275 (8073, 8061);
  not ginst2276 (8074, 8064);
  or ginst2277 (8075, 7526, 8071, 3659, 2625);
  or ginst2278 (8076, 7636, 8072, 3661, 2627);
  and ginst2279 (8077, 8073, 1727);
  and ginst2280 (8078, 8074, 1727);
  or ginst2281 (8079, 7530, 8077);
  or ginst2282 (8082, 7479, 8078);
  and ginst2283 (8089, 8079, 3063);
  and ginst2284 (8090, 8082, 3063);
  and ginst2285 (8091, 8079, 3063);
  and ginst2286 (8092, 8082, 3063);
  or ginst2287 (8093, 8089, 3071);
  or ginst2288 (8096, 8090, 3072);
  or ginst2289 (8099, 8091, 3073);
  or ginst2290 (8102, 8092, 3074);
  and ginst2291 (8113, 8102, 2779, 2790);
  and ginst2292 (8114, 8099, 1327, 2790);
  and ginst2293 (8115, 8102, 2801, 2812);
  and ginst2294 (8116, 8099, 1351, 2812);
  and ginst2295 (8117, 8096, 2681, 2692);
  and ginst2296 (8118, 8093, 1185, 2692);
  and ginst2297 (8119, 8096, 2756, 2767);
  and ginst2298 (8120, 8093, 1247, 2767);
  or ginst2299 (8121, 8117, 8118, 3662, 2703);
  or ginst2300 (8122, 8119, 8120, 3663, 2778);
  or ginst2301 (8123, 8113, 8114, 3650, 2614);
  or ginst2302 (8124, 8115, 8116, 3658, 2622);
  and ginst2303 (8125, 8121, 2675);
  and ginst2304 (8126, 8122, 2750);
  not ginst2305 (8127, 8125);
  not ginst2306 (8128, 8126);
  buf ginst2307 (816, 293);

endmodule
