// Main module
module c3540(N1, N13, N20, N33, N41, N45, N50, N58, N68, N77, N87, N97, N107, N116, N124, N125, N128, N132, N137, N143, N150, N159, N169, N179, N190, N200, N213, N222, N223, N226, N232, N238, N244, N250, N257, N264, N270, N274, N283, N294, N303, N311, N317, N322, N326, N329, N330, N343, N349, N350, N1713, N1947, N3195, N3833, N3987, N4028, N4145, N4589, N4667, N4815, N4944, N5002, N5045, N5047, N5078, N5102, N5120, N5121, N5192, N5231, N5360, N5361);

  input N1, N13, N20, N33, N41, N45, N50, N58, N68, N77, N87, N97, N107, N116, N124, N125, N128, N132, N137, N143, N150, N159, N169, N179, N190, N200, N213, N222, N223, N226, N232, N238, N244, N250, N257, N264, N270, N274, N283, N294, N303, N311, N317, N322, N326, N329, N330, N343, N349, N350;
  output N1713, N1947, N3195, N3833, N3987, N4028, N4145, N4589, N4667, N4815, N4944, N5002, N5045, N5047, N5078, N5102, N5120, N5121, N5192, N5231, N5360, N5361;
  wire N655, N665, N670, N679, N683, N686, N690, N699, N702, N706, N715, N724, N727, N736, N740, N749, N753, N763, N768, N769, N772, N779, N782, N786, N793, N794, N798, N803, N820, N821, N825, N829, N832, N835, N836, N839, N842, N845, N848, N851, N854, N858, N861, N864, N867, N870, N874, N877, N880, N883, N886, N889, N890, N891, N892, N895, N896, N913, N914, N915, N916, N917, N920, N923, N926, N929, N932, N935, N938, N941, N944, N947, N950, N953, N956, N959, N962, N965, N1067, N1117, N1179, N1196, N1197, N1202, N1219, N1250, N1251, N1252, N1253, N1254, N1255, N1256, N1257, N1258, N1259, N1260, N1261, N1262, N1263, N1264, N1267, N1268, N1271, N1272, N1273, N1276, N1279, N1298, N1302, N1306, N1315, N1322, N1325, N1328, N1331, N1334, N1337, N1338, N1339, N1340, N1343, N1344, N1345, N1346, N1347, N1348, N1349, N1350, N1351, N1352, N1353, N1358, N1363, N1366, N1369, N1384, N1401, N1402, N1403, N1404, N1405, N1406, N1407, N1408, N1409, N1426, N1427, N1452, N1459, N1460, N1461, N1464, N1467, N1468, N1469, N1470, N1471, N1474, N1475, N1478, N1481, N1484, N1487, N1490, N1493, N1496, N1499, N1502, N1505, N1507, N1508, N1509, N1510, N1511, N1512, N1520, N1562, N1579, N1580, N1581, N1582, N1583, N1584, N1585, N1586, N1587, N1588, N1589, N1590, N1591, N1592, N1593, N1594, N1595, N1596, N1597, N1598, N1599, N1600, N1643, N1644, N1645, N1646, N1647, N1648, N1649, N1650, N1667, N1670, N1673, N1674, N1675, N1676, N1677, N1678, N1679, N1680, N1691, N1692, N1693, N1694, N1714, N1715, N1718, N1721, N1722, N1725, N1726, N1727, N1728, N1729, N1730, N1731, N1735, N1736, N1737, N1738, N1747, N1756, N1761, N1764, N1765, N1766, N1767, N1768, N1769, N1770, N1787, N1788, N1789, N1790, N1791, N1792, N1793, N1794, N1795, N1796, N1797, N1798, N1799, N1800, N1801, N1802, N1803, N1806, N1809, N1812, N1815, N1818, N1821, N1824, N1833, N1842, N1843, N1844, N1845, N1846, N1847, N1848, N1849, N1850, N1851, N1852, N1853, N1854, N1855, N1856, N1857, N1858, N1859, N1860, N1861, N1862, N1863, N1864, N1869, N1870, N1873, N1874, N1875, N1878, N1879, N1880, N1883, N1884, N1885, N1888, N1889, N1890, N1893, N1894, N1895, N1898, N1899, N1900, N1903, N1904, N1905, N1908, N1909, N1912, N1913, N1917, N1922, N1926, N1930, N1933, N1936, N1939, N1940, N1941, N1942, N1943, N1944, N1945, N1946, N1960, N1961, N1966, N1981, N1982, N1983, N1986, N1987, N1988, N1989, N1990, N1991, N2022, N2023, N2024, N2025, N2026, N2027, N2028, N2029, N2030, N2031, N2032, N2033, N2034, N2035, N2036, N2037, N2038, N2043, N2052, N2057, N2068, N2073, N2078, N2083, N2088, N2093, N2098, N2103, N2121, N2122, N2123, N2124, N2125, N2126, N2127, N2128, N2133, N2134, N2135, N2136, N2137, N2138, N2139, N2141, N2142, N2143, N2144, N2145, N2146, N2147, N2148, N2149, N2150, N2151, N2152, N2153, N2154, N2155, N2156, N2157, N2158, N2175, N2178, N2179, N2180, N2181, N2183, N2184, N2185, N2188, N2191, N2194, N2197, N2200, N2203, N2206, N2209, N2210, N2211, N2212, N2221, N2230, N2231, N2232, N2233, N2234, N2235, N2236, N2237, N2238, N2239, N2240, N2241, N2242, N2243, N2244, N2245, N2270, N2277, N2282, N2287, N2294, N2299, N2304, N2307, N2310, N2313, N2316, N2319, N2322, N2325, N2328, N2331, N2334, N2341, N2342, N2347, N2348, N2349, N2350, N2351, N2352, N2353, N2354, N2355, N2374, N2375, N2376, N2379, N2398, N2417, N2418, N2419, N2420, N2421, N2422, N2425, N2426, N2427, N2430, N2431, N2432, N2435, N2436, N2437, N2438, N2439, N2440, N2443, N2444, N2445, N2448, N2449, N2450, N2467, N2468, N2469, N2470, N2471, N2474, N2475, N2476, N2477, N2478, N2481, N2482, N2483, N2486, N2487, N2488, N2497, N2506, N2515, N2524, N2533, N2542, N2551, N2560, N2569, N2578, N2587, N2596, N2605, N2614, N2623, N2632, N2633, N2634, N2635, N2636, N2637, N2638, N2639, N2640, N2641, N2642, N2643, N2644, N2645, N2646, N2647, N2648, N2652, N2656, N2659, N2662, N2666, N2670, N2673, N2677, N2681, N2684, N2688, N2692, N2697, N2702, N2706, N2710, N2715, N2719, N2723, N2728, N2729, N2730, N2731, N2732, N2733, N2734, N2735, N2736, N2737, N2738, N2739, N2740, N2741, N2742, N2743, N2744, N2745, N2746, N2748, N2749, N2750, N2751, N2754, N2755, N2756, N2757, N2758, N2761, N2764, N2768, N2769, N2898, N2899, N2900, N2901, N2962, N2966, N2967, N2970, N2973, N2977, N2980, N2984, N2985, N2986, N2987, N2988, N2989, N2990, N2991, N2992, N2993, N2994, N2995, N2996, N2997, N2998, N2999, N3000, N3001, N3002, N3003, N3004, N3005, N3006, N3007, N3008, N3009, N3010, N3011, N3012, N3013, N3014, N3015, N3016, N3017, N3018, N3019, N3020, N3021, N3022, N3023, N3024, N3025, N3026, N3027, N3028, N3029, N3030, N3031, N3032, N3033, N3034, N3035, N3036, N3037, N3038, N3039, N3040, N3041, N3042, N3043, N3044, N3045, N3046, N3047, N3048, N3049, N3050, N3051, N3052, N3053, N3054, N3055, N3056, N3057, N3058, N3059, N3060, N3061, N3062, N3063, N3064, N3065, N3066, N3067, N3068, N3069, N3070, N3071, N3072, N3073, N3074, N3075, N3076, N3077, N3078, N3079, N3080, N3081, N3082, N3083, N3084, N3085, N3086, N3087, N3088, N3089, N3090, N3091, N3092, N3093, N3094, N3095, N3096, N3097, N3098, N3099, N3100, N3101, N3102, N3103, N3104, N3105, N3106, N3107, N3108, N3109, N3110, N3111, N3112, N3115, N3118, N3119, N3122, N3125, N3128, N3131, N3134, N3135, N3138, N3141, N3142, N3145, N3148, N3149, N3152, N3155, N3158, N3161, N3164, N3165, N3168, N3171, N3172, N3175, N3178, N3181, N3184, N3187, N3190, N3191, N3192, N3193, N3194, N3196, N3206, N3207, N3208, N3209, N3210, N3211, N3212, N3213, N3214, N3215, N3216, N3217, N3218, N3219, N3220, N3221, N3222, N3223, N3224, N3225, N3226, N3227, N3228, N3229, N3230, N3231, N3232, N3233, N3234, N3235, N3236, N3237, N3238, N3239, N3240, N3241, N3242, N3243, N3244, N3245, N3246, N3247, N3248, N3249, N3250, N3251, N3252, N3253, N3254, N3255, N3256, N3257, N3258, N3259, N3260, N3261, N3262, N3263, N3264, N3265, N3266, N3267, N3268, N3269, N3270, N3271, N3272, N3273, N3274, N3275, N3276, N3277, N3278, N3279, N3280, N3281, N3282, N3283, N3284, N3285, N3286, N3287, N3288, N3289, N3290, N3291, N3292, N3293, N3294, N3295, N3296, N3297, N3298, N3299, N3300, N3301, N3302, N3303, N3304, N3305, N3306, N3307, N3308, N3309, N3310, N3311, N3312, N3313, N3314, N3315, N3316, N3317, N3318, N3319, N3320, N3321, N3322, N3323, N3324, N3325, N3326, N3327, N3328, N3329, N3330, N3331, N3332, N3333, N3334, N3383, N3384, N3387, N3388, N3389, N3390, N3391, N3392, N3393, N3394, N3395, N3396, N3397, N3398, N3399, N3400, N3401, N3402, N3403, N3404, N3405, N3406, N3407, N3410, N3413, N3414, N3415, N3419, N3423, N3426, N3429, N3430, N3431, N3434, N3437, N3438, N3439, N3442, N3445, N3446, N3447, N3451, N3455, N3458, N3461, N3462, N3463, N3466, N3469, N3470, N3471, N3472, N3475, N3478, N3481, N3484, N3487, N3490, N3493, N3496, N3499, N3502, N3505, N3508, N3511, N3514, N3517, N3520, N3523, N3534, N3535, N3536, N3537, N3538, N3539, N3540, N3541, N3542, N3543, N3544, N3545, N3546, N3547, N3548, N3549, N3550, N3551, N3552, N3557, N3568, N3573, N3578, N3589, N3594, N3605, N3626, N3627, N3628, N3629, N3630, N3631, N3632, N3633, N3634, N3635, N3636, N3637, N3638, N3639, N3640, N3641, N3642, N3643, N3644, N3645, N3648, N3651, N3652, N3653, N3654, N3657, N3658, N3661, N3662, N3663, N3664, N3667, N3670, N3671, N3672, N3673, N3676, N3677, N3680, N3681, N3682, N3685, N3686, N3687, N3688, N3689, N3690, N3693, N3694, N3695, N3696, N3697, N3700, N3703, N3704, N3705, N3706, N3707, N3708, N3711, N3712, N3713, N3714, N3715, N3716, N3717, N3718, N3719, N3720, N3721, N3731, N3734, N3740, N3743, N3753, N3756, N3762, N3765, N3766, N3773, N3774, N3775, N3776, N3777, N3778, N3779, N3780, N3786, N3789, N3800, N3803, N3809, N3812, N3815, N3818, N3821, N3824, N3827, N3830, N3834, N3835, N3838, N3845, N3850, N3855, N3858, N3861, N3865, N3868, N3884, N3885, N3894, N3895, N3898, N3899, N3906, N3911, N3912, N3913, N3916, N3917, N3920, N3921, N3924, N3925, N3926, N3930, N3931, N3932, N3935, N3936, N3937, N3940, N3947, N3948, N3950, N3953, N3956, N3959, N3962, N3965, N3968, N3971, N3974, N3977, N3980, N3983, N3992, N3996, N4013, N4029, N4030, N4031, N4032, N4033, N4034, N4035, N4042, N4043, N4044, N4045, N4046, N4047, N4048, N4049, N4050, N4051, N4052, N4053, N4054, N4055, N4056, N4057, N4058, N4059, N4062, N4065, N4066, N4067, N4070, N4073, N4074, N4075, N4076, N4077, N4078, N4079, N4080, N4085, N4086, N4088, N4090, N4091, N4094, N4098, N4101, N4104, N4105, N4106, N4107, N4108, N4109, N4110, N4111, N4112, N4113, N4114, N4115, N4116, N4119, N4122, N4123, N4126, N4127, N4128, N4139, N4142, N4146, N4147, N4148, N4149, N4150, N4151, N4152, N4153, N4154, N4161, N4167, N4174, N4182, N4186, N4189, N4190, N4191, N4192, N4193, N4194, N4195, N4196, N4197, N4200, N4203, N4209, N4213, N4218, N4223, N4238, N4239, N4241, N4242, N4247, N4251, N4252, N4253, N4254, N4255, N4256, N4257, N4258, N4283, N4284, N4287, N4291, N4295, N4296, N4299, N4303, N4304, N4305, N4310, N4316, N4317, N4318, N4319, N4322, N4325, N4326, N4327, N4328, N4329, N4330, N4331, N4335, N4338, N4341, N4344, N4347, N4350, N4353, N4356, N4359, N4362, N4365, N4368, N4371, N4376, N4377, N4387, N4390, N4393, N4398, N4413, N4416, N4421, N4427, N4430, N4435, N4442, N4443, N4446, N4447, N4448, N4452, N4458, N4461, N4462, N4463, N4464, N4465, N4468, N4472, N4475, N4479, N4484, N4486, N4487, N4491, N4493, N4496, N4497, N4498, N4503, N4506, N4507, N4508, N4509, N4510, N4511, N4515, N4526, N4527, N4528, N4529, N4530, N4531, N4534, N4537, N4540, N4545, N4549, N4552, N4555, N4558, N4559, N4562, N4563, N4564, N4568, N4569, N4572, N4573, N4576, N4581, N4584, N4587, N4588, N4593, N4596, N4597, N4599, N4602, N4603, N4608, N4613, N4616, N4619, N4623, N4628, N4629, N4630, N4635, N4636, N4640, N4641, N4642, N4643, N4644, N4647, N4650, N4656, N4659, N4664, N4668, N4669, N4670, N4673, N4674, N4675, N4676, N4677, N4678, N4679, N4687, N4688, N4691, N4694, N4697, N4700, N4704, N4705, N4706, N4707, N4708, N4711, N4716, N4717, N4721, N4722, N4726, N4727, N4730, N4733, N4740, N4743, N4747, N4748, N4749, N4750, N4753, N4754, N4755, N4756, N4757, N4769, N4772, N4775, N4778, N4786, N4787, N4788, N4789, N4794, N4797, N4800, N4805, N4808, N4812, N4816, N4817, N4818, N4822, N4823, N4826, N4829, N4830, N4831, N4838, N4844, N4847, N4850, N4854, N4859, N4860, N4868, N4870, N4872, N4873, N4876, N4880, N4885, N4889, N4895, N4896, N4897, N4898, N4899, N4900, N4901, N4902, N4904, N4905, N4906, N4907, N4913, N4916, N4920, N4921, N4924, N4925, N4926, N4928, N4929, N4930, N4931, N4937, N4940, N4946, N4949, N4950, N4951, N4952, N4953, N4954, N4957, N4964, N4965, N4968, N4969, N4970, N4973, N4978, N4979, N4980, N4981, N4982, N4983, N4984, N4985, N4988, N4991, N4996, N4999, N5007, N5010, N5013, N5018, N5021, N5026, N5029, N5030, N5039, N5042, N5046, N5050, N5055, N5058, N5061, N5066, N5070, N5080, N5085, N5094, N5095, N5097, N5103, N5108, N5109, N5110, N5111, N5114, N5117, N5122, N5125, N5128, N5133, N5136, N5139, N5145, N5151, N5154, N5159, N5160, N5163, N5166, N5173, N5174, N5177, N5182, N5183, N5184, N5188, N5193, N5196, N5197, N5198, N5199, N5201, N5203, N5205, N5209, N5212, N5215, N5217, N5219, N5220, N5221, N5222, N5223, N5224, N5225, N5228, N5232, N5233, N5234, N5235, N5236, N5240, N5242, N5243, N5245, N5246, N5250, N5253, N5254, N5257, N5258, N5261, N5266, N5269, N5277, N5278, N5279, N5283, N5284, N5285, N5286, N5289, N5292, N5295, N5298, N5303, N5306, N5309, N5312, N5313, N5322, N5323, N5324, N5327, N5332, N5335, N5340, N5341, N5344, N5345, N5348, N5349, N5350, N5351, N5352, N5353, N5354, N5355, N5356, N5357, N5358, N5359;

  and ginst1 (N1067, N768, N250);
  or ginst2 (N1117, N820, N20);
  or ginst3 (N1179, N895, N169);
  not ginst4 (N1196, N793);
  or ginst5 (N1197, N915, N1);
  and ginst6 (N1202, N913, N914);
  or ginst7 (N1219, N916, N1);
  and ginst8 (N1250, N842, N848, N854);
  nand ginst9 (N1251, N655, N226);
  nand ginst10 (N1252, N670, N232);
  nand ginst11 (N1253, N690, N238);
  nand ginst12 (N1254, N706, N244);
  nand ginst13 (N1255, N715, N250);
  nand ginst14 (N1256, N727, N257);
  nand ginst15 (N1257, N740, N264);
  nand ginst16 (N1258, N753, N270);
  not ginst17 (N1259, N926);
  not ginst18 (N1260, N929);
  not ginst19 (N1261, N932);
  not ginst20 (N1262, N935);
  nand ginst21 (N1263, N679, N686);
  nand ginst22 (N1264, N736, N749);
  nand ginst23 (N1267, N683, N699);
  buf ginst24 (N1268, N665);
  not ginst25 (N1271, N953);
  not ginst26 (N1272, N959);
  buf ginst27 (N1273, N839);
  buf ginst28 (N1276, N839);
  buf ginst29 (N1279, N782);
  buf ginst30 (N1298, N825);
  buf ginst31 (N1302, N832);
  and ginst32 (N1306, N779, N835);
  and ginst33 (N1315, N779, N832, N836);
  and ginst34 (N1322, N769, N836);
  and ginst35 (N1325, N772, N786, N798);
  nand ginst36 (N1328, N772, N786, N798);
  nand ginst37 (N1331, N772, N786);
  buf ginst38 (N1334, N874);
  nand ginst39 (N1337, N782, N794, N45);
  nand ginst40 (N1338, N842, N848, N854);
  not ginst41 (N1339, N956);
  and ginst42 (N1340, N861, N867, N870);
  nand ginst43 (N1343, N861, N867, N870);
  not ginst44 (N1344, N962);
  not ginst45 (N1345, N803);
  not ginst46 (N1346, N803);
  not ginst47 (N1347, N803);
  not ginst48 (N1348, N803);
  not ginst49 (N1349, N803);
  not ginst50 (N1350, N803);
  not ginst51 (N1351, N803);
  not ginst52 (N1352, N803);
  or ginst53 (N1353, N883, N886);
  nor ginst54 (N1358, N883, N886);
  buf ginst55 (N1363, N892);
  not ginst56 (N1366, N892);
  buf ginst57 (N1369, N821);
  buf ginst58 (N1384, N825);
  not ginst59 (N1401, N896);
  not ginst60 (N1402, N896);
  not ginst61 (N1403, N896);
  not ginst62 (N1404, N896);
  not ginst63 (N1405, N896);
  not ginst64 (N1406, N896);
  not ginst65 (N1407, N896);
  not ginst66 (N1408, N896);
  or ginst67 (N1409, N1196, N1);
  not ginst68 (N1426, N829);
  not ginst69 (N1427, N829);
  and ginst70 (N1452, N769, N782, N794);
  not ginst71 (N1459, N917);
  not ginst72 (N1460, N965);
  or ginst73 (N1461, N920, N923);
  nor ginst74 (N1464, N920, N923);
  not ginst75 (N1467, N938);
  not ginst76 (N1468, N941);
  not ginst77 (N1469, N944);
  not ginst78 (N1470, N947);
  buf ginst79 (N1471, N679);
  not ginst80 (N1474, N950);
  buf ginst81 (N1475, N686);
  buf ginst82 (N1478, N702);
  buf ginst83 (N1481, N724);
  buf ginst84 (N1484, N736);
  buf ginst85 (N1487, N749);
  buf ginst86 (N1490, N763);
  buf ginst87 (N1493, N877);
  buf ginst88 (N1496, N877);
  buf ginst89 (N1499, N880);
  buf ginst90 (N1502, N880);
  nand ginst91 (N1505, N702, N1250);
  and ginst92 (N1507, N1251, N1252, N1253, N1254);
  and ginst93 (N1508, N1255, N1256, N1257, N1258);
  nand ginst94 (N1509, N929, N1259);
  nand ginst95 (N1510, N926, N1260);
  nand ginst96 (N1511, N935, N1261);
  nand ginst97 (N1512, N932, N1262);
  and ginst98 (N1520, N655, N1263);
  and ginst99 (N1562, N874, N1337);
  not ginst100 (N1579, N1117);
  and ginst101 (N1580, N803, N1117);
  and ginst102 (N1581, N1338, N1345);
  not ginst103 (N1582, N1117);
  and ginst104 (N1583, N803, N1117);
  not ginst105 (N1584, N1117);
  and ginst106 (N1585, N803, N1117);
  and ginst107 (N1586, N854, N1347);
  not ginst108 (N1587, N1117);
  and ginst109 (N1588, N803, N1117);
  and ginst110 (N1589, N1348, N77);
  not ginst111 (N1590, N1117);
  and ginst112 (N1591, N803, N1117);
  and ginst113 (N1592, N1343, N1349);
  not ginst114 (N1593, N1117);
  and ginst115 (N1594, N803, N1117);
  not ginst116 (N1595, N1117);
  and ginst117 (N1596, N803, N1117);
  and ginst118 (N1597, N870, N1351);
  not ginst119 (N1598, N1117);
  and ginst120 (N1599, N803, N1117);
  and ginst121 (N1600, N1352, N116);
  and ginst122 (N1643, N1401, N222);
  and ginst123 (N1644, N1402, N223);
  and ginst124 (N1645, N1403, N226);
  and ginst125 (N1646, N1404, N232);
  and ginst126 (N1647, N1405, N238);
  and ginst127 (N1648, N1406, N244);
  and ginst128 (N1649, N1407, N250);
  and ginst129 (N1650, N1408, N257);
  and ginst130 (N1667, N1426, N1, N13);
  and ginst131 (N1670, N1427, N1, N13);
  not ginst132 (N1673, N1202);
  not ginst133 (N1674, N1202);
  not ginst134 (N1675, N1202);
  not ginst135 (N1676, N1202);
  not ginst136 (N1677, N1202);
  not ginst137 (N1678, N1202);
  not ginst138 (N1679, N1202);
  not ginst139 (N1680, N1202);
  nand ginst140 (N1691, N941, N1467);
  nand ginst141 (N1692, N938, N1468);
  nand ginst142 (N1693, N947, N1469);
  nand ginst143 (N1694, N944, N1470);
  not ginst144 (N1713, N1505);
  and ginst145 (N1714, N1264, N87);
  nand ginst146 (N1715, N1509, N1510);
  nand ginst147 (N1718, N1511, N1512);
  nand ginst148 (N1721, N1507, N1508);
  and ginst149 (N1722, N763, N1340);
  nand ginst150 (N1725, N763, N1340);
  not ginst151 (N1726, N1268);
  nand ginst152 (N1727, N1271, N1493);
  not ginst153 (N1728, N1493);
  and ginst154 (N1729, N683, N1268);
  nand ginst155 (N1730, N1272, N1499);
  not ginst156 (N1731, N1499);
  nand ginst157 (N1735, N1264, N87);
  not ginst158 (N1736, N1273);
  not ginst159 (N1737, N1276);
  nand ginst160 (N1738, N821, N1325);
  nand ginst161 (N1747, N825, N1325);
  nand ginst162 (N1756, N772, N798, N1279);
  nand ginst163 (N1761, N772, N786, N798, N1302);
  nand ginst164 (N1764, N1339, N1496);
  not ginst165 (N1765, N1496);
  nand ginst166 (N1766, N1344, N1502);
  not ginst167 (N1767, N1502);
  not ginst168 (N1768, N1328);
  not ginst169 (N1769, N1334);
  not ginst170 (N1770, N1331);
  and ginst171 (N1787, N845, N1579);
  and ginst172 (N1788, N1580, N150);
  and ginst173 (N1789, N851, N1582);
  and ginst174 (N1790, N1583, N159);
  and ginst175 (N1791, N1584, N77);
  and ginst176 (N1792, N1585, N50);
  and ginst177 (N1793, N858, N1587);
  and ginst178 (N1794, N845, N1588);
  and ginst179 (N1795, N864, N1590);
  and ginst180 (N1796, N851, N1591);
  and ginst181 (N1797, N1593, N107);
  and ginst182 (N1798, N1594, N77);
  and ginst183 (N1799, N1595, N116);
  and ginst184 (N1800, N858, N1596);
  and ginst185 (N1801, N1598, N283);
  and ginst186 (N1802, N864, N1599);
  and ginst187 (N1803, N1363, N200);
  and ginst188 (N1806, N889, N1363);
  and ginst189 (N1809, N890, N1366);
  and ginst190 (N1812, N891, N1366);
  nand ginst191 (N1815, N1298, N1302);
  nand ginst192 (N1818, N821, N1302);
  nand ginst193 (N1821, N772, N1179, N1279);
  nand ginst194 (N1824, N786, N794, N1298);
  nand ginst195 (N1833, N786, N1298);
  not ginst196 (N1842, N1369);
  not ginst197 (N1843, N1369);
  not ginst198 (N1844, N1369);
  not ginst199 (N1845, N1369);
  not ginst200 (N1846, N1369);
  not ginst201 (N1847, N1369);
  not ginst202 (N1848, N1369);
  not ginst203 (N1849, N1384);
  and ginst204 (N1850, N896, N1384);
  not ginst205 (N1851, N1384);
  and ginst206 (N1852, N896, N1384);
  not ginst207 (N1853, N1384);
  and ginst208 (N1854, N896, N1384);
  not ginst209 (N1855, N1384);
  and ginst210 (N1856, N896, N1384);
  not ginst211 (N1857, N1384);
  and ginst212 (N1858, N896, N1384);
  not ginst213 (N1859, N1384);
  and ginst214 (N1860, N896, N1384);
  not ginst215 (N1861, N1384);
  and ginst216 (N1862, N896, N1384);
  not ginst217 (N1863, N1384);
  and ginst218 (N1864, N896, N1384);
  and ginst219 (N1869, N1202, N1409);
  nor ginst220 (N1870, N1409, N50);
  not ginst221 (N1873, N1306);
  and ginst222 (N1874, N1202, N1409);
  nor ginst223 (N1875, N1409, N58);
  not ginst224 (N1878, N1306);
  and ginst225 (N1879, N1202, N1409);
  nor ginst226 (N1880, N1409, N68);
  not ginst227 (N1883, N1306);
  and ginst228 (N1884, N1202, N1409);
  nor ginst229 (N1885, N1409, N77);
  not ginst230 (N1888, N1306);
  and ginst231 (N1889, N1202, N1409);
  nor ginst232 (N1890, N1409, N87);
  not ginst233 (N1893, N1322);
  and ginst234 (N1894, N1202, N1409);
  nor ginst235 (N1895, N1409, N97);
  not ginst236 (N1898, N1315);
  and ginst237 (N1899, N1202, N1409);
  nor ginst238 (N1900, N1409, N107);
  not ginst239 (N1903, N1315);
  and ginst240 (N1904, N1202, N1409);
  nor ginst241 (N1905, N1409, N116);
  not ginst242 (N1908, N1315);
  and ginst243 (N1909, N1452, N213);
  nand ginst244 (N1912, N1452, N213);
  and ginst245 (N1913, N1452, N213, N343);
  nand ginst246 (N1917, N1452, N213, N343);
  and ginst247 (N1922, N1452, N213, N343);
  nand ginst248 (N1926, N1452, N213, N343);
  buf ginst249 (N1930, N1464);
  nand ginst250 (N1933, N1691, N1692);
  nand ginst251 (N1936, N1693, N1694);
  not ginst252 (N1939, N1471);
  nand ginst253 (N1940, N1471, N1474);
  not ginst254 (N1941, N1475);
  not ginst255 (N1942, N1478);
  not ginst256 (N1943, N1481);
  not ginst257 (N1944, N1484);
  not ginst258 (N1945, N1487);
  not ginst259 (N1946, N1490);
  not ginst260 (N1947, N1714);
  nand ginst261 (N1960, N953, N1728);
  nand ginst262 (N1961, N959, N1731);
  and ginst263 (N1966, N1276, N1520);
  nand ginst264 (N1981, N956, N1765);
  nand ginst265 (N1982, N962, N1767);
  and ginst266 (N1983, N1067, N1768);
  or ginst267 (N1986, N1581, N1787, N1788);
  or ginst268 (N1987, N1586, N1791, N1792);
  or ginst269 (N1988, N1589, N1793, N1794);
  or ginst270 (N1989, N1592, N1795, N1796);
  or ginst271 (N1990, N1597, N1799, N1800);
  or ginst272 (N1991, N1600, N1801, N1802);
  and ginst273 (N2022, N1849, N77);
  and ginst274 (N2023, N1850, N223);
  and ginst275 (N2024, N1851, N87);
  and ginst276 (N2025, N1852, N226);
  and ginst277 (N2026, N1853, N97);
  and ginst278 (N2027, N1854, N232);
  and ginst279 (N2028, N1855, N107);
  and ginst280 (N2029, N1856, N238);
  and ginst281 (N2030, N1857, N116);
  and ginst282 (N2031, N1858, N244);
  and ginst283 (N2032, N1859, N283);
  and ginst284 (N2033, N1860, N250);
  and ginst285 (N2034, N1861, N294);
  and ginst286 (N2035, N1862, N257);
  and ginst287 (N2036, N1863, N303);
  and ginst288 (N2037, N1864, N264);
  buf ginst289 (N2038, N1667);
  not ginst290 (N2043, N1667);
  buf ginst291 (N2052, N1670);
  not ginst292 (N2057, N1670);
  and ginst293 (N2068, N1197, N1869, N50);
  and ginst294 (N2073, N1197, N1874, N58);
  and ginst295 (N2078, N1197, N1879, N68);
  and ginst296 (N2083, N1197, N1884, N77);
  and ginst297 (N2088, N1219, N1889, N87);
  and ginst298 (N2093, N1219, N1894, N97);
  and ginst299 (N2098, N1219, N1899, N107);
  and ginst300 (N2103, N1219, N1904, N116);
  not ginst301 (N2121, N1562);
  not ginst302 (N2122, N1562);
  not ginst303 (N2123, N1562);
  not ginst304 (N2124, N1562);
  not ginst305 (N2125, N1562);
  not ginst306 (N2126, N1562);
  not ginst307 (N2127, N1562);
  not ginst308 (N2128, N1562);
  nand ginst309 (N2133, N950, N1939);
  nand ginst310 (N2134, N1478, N1941);
  nand ginst311 (N2135, N1475, N1942);
  nand ginst312 (N2136, N1484, N1943);
  nand ginst313 (N2137, N1481, N1944);
  nand ginst314 (N2138, N1490, N1945);
  nand ginst315 (N2139, N1487, N1946);
  not ginst316 (N2141, N1933);
  not ginst317 (N2142, N1936);
  not ginst318 (N2143, N1738);
  and ginst319 (N2144, N1738, N1747);
  not ginst320 (N2145, N1747);
  nand ginst321 (N2146, N1727, N1960);
  nand ginst322 (N2147, N1730, N1961);
  and ginst323 (N2148, N665, N1267, N1722, N58);
  not ginst324 (N2149, N1738);
  and ginst325 (N2150, N1738, N1747);
  not ginst326 (N2151, N1747);
  not ginst327 (N2152, N1738);
  not ginst328 (N2153, N1747);
  and ginst329 (N2154, N1738, N1747);
  not ginst330 (N2155, N1738);
  not ginst331 (N2156, N1747);
  and ginst332 (N2157, N1738, N1747);
  buf ginst333 (N2158, N1761);
  buf ginst334 (N2175, N1761);
  nand ginst335 (N2178, N1764, N1981);
  nand ginst336 (N2179, N1766, N1982);
  not ginst337 (N2180, N1756);
  and ginst338 (N2181, N1328, N1756);
  not ginst339 (N2183, N1756);
  and ginst340 (N2184, N1331, N1756);
  nand ginst341 (N2185, N1358, N1812);
  nand ginst342 (N2188, N1358, N1809);
  nand ginst343 (N2191, N1353, N1812);
  nand ginst344 (N2194, N1353, N1809);
  nand ginst345 (N2197, N1358, N1806);
  nand ginst346 (N2200, N1358, N1803);
  nand ginst347 (N2203, N1353, N1806);
  nand ginst348 (N2206, N1353, N1803);
  not ginst349 (N2209, N1815);
  not ginst350 (N2210, N1818);
  and ginst351 (N2211, N1815, N1818);
  buf ginst352 (N2212, N1821);
  buf ginst353 (N2221, N1821);
  not ginst354 (N2230, N1833);
  not ginst355 (N2231, N1833);
  not ginst356 (N2232, N1833);
  not ginst357 (N2233, N1833);
  not ginst358 (N2234, N1824);
  not ginst359 (N2235, N1824);
  not ginst360 (N2236, N1824);
  not ginst361 (N2237, N1824);
  or ginst362 (N2238, N1643, N2022, N2023);
  or ginst363 (N2239, N1644, N2024, N2025);
  or ginst364 (N2240, N1645, N2026, N2027);
  or ginst365 (N2241, N1646, N2028, N2029);
  or ginst366 (N2242, N1647, N2030, N2031);
  or ginst367 (N2243, N1648, N2032, N2033);
  or ginst368 (N2244, N1649, N2034, N2035);
  or ginst369 (N2245, N1650, N2036, N2037);
  and ginst370 (N2270, N1673, N1986);
  and ginst371 (N2277, N1675, N1987);
  and ginst372 (N2282, N1676, N1988);
  and ginst373 (N2287, N1677, N1989);
  and ginst374 (N2294, N1679, N1990);
  and ginst375 (N2299, N1680, N1991);
  buf ginst376 (N2304, N1917);
  and ginst377 (N2307, N1930, N350);
  nand ginst378 (N2310, N1930, N350);
  buf ginst379 (N2313, N1715);
  buf ginst380 (N2316, N1718);
  buf ginst381 (N2319, N1715);
  buf ginst382 (N2322, N1718);
  nand ginst383 (N2325, N1940, N2133);
  nand ginst384 (N2328, N2134, N2135);
  nand ginst385 (N2331, N2136, N2137);
  nand ginst386 (N2334, N2138, N2139);
  nand ginst387 (N2341, N1936, N2141);
  nand ginst388 (N2342, N1933, N2142);
  and ginst389 (N2347, N724, N2144);
  and ginst390 (N2348, N699, N1726, N2146);
  and ginst391 (N2349, N753, N2147);
  and ginst392 (N2350, N1273, N2148);
  and ginst393 (N2351, N736, N2150);
  and ginst394 (N2352, N1735, N2153);
  and ginst395 (N2353, N763, N2154);
  and ginst396 (N2354, N1725, N2156);
  and ginst397 (N2355, N749, N2157);
  not ginst398 (N2374, N2178);
  not ginst399 (N2375, N2179);
  and ginst400 (N2376, N1520, N2180);
  and ginst401 (N2379, N1721, N2181);
  and ginst402 (N2398, N665, N2211);
  and ginst403 (N2417, N1873, N2057, N226);
  and ginst404 (N2418, N1306, N2057, N274);
  and ginst405 (N2419, N2052, N2238);
  and ginst406 (N2420, N1878, N2057, N232);
  and ginst407 (N2421, N1306, N2057, N274);
  and ginst408 (N2422, N2052, N2239);
  and ginst409 (N2425, N1883, N2057, N238);
  and ginst410 (N2426, N1306, N2057, N274);
  and ginst411 (N2427, N2052, N2240);
  and ginst412 (N2430, N1888, N2057, N244);
  and ginst413 (N2431, N1306, N2057, N274);
  and ginst414 (N2432, N2052, N2241);
  and ginst415 (N2435, N1893, N2043, N250);
  and ginst416 (N2436, N1322, N2043, N274);
  and ginst417 (N2437, N2038, N2242);
  and ginst418 (N2438, N1898, N2043, N257);
  and ginst419 (N2439, N1315, N2043, N274);
  and ginst420 (N2440, N2038, N2243);
  and ginst421 (N2443, N1903, N2043, N264);
  and ginst422 (N2444, N1315, N2043, N274);
  and ginst423 (N2445, N2038, N2244);
  and ginst424 (N2448, N1908, N2043, N270);
  and ginst425 (N2449, N1315, N2043, N274);
  and ginst426 (N2450, N2038, N2245);
  not ginst427 (N2467, N2313);
  not ginst428 (N2468, N2316);
  not ginst429 (N2469, N2319);
  not ginst430 (N2470, N2322);
  nand ginst431 (N2471, N2341, N2342);
  not ginst432 (N2474, N2325);
  not ginst433 (N2475, N2328);
  not ginst434 (N2476, N2331);
  not ginst435 (N2477, N2334);
  or ginst436 (N2478, N1729, N2348);
  not ginst437 (N2481, N2175);
  and ginst438 (N2482, N1334, N2175);
  and ginst439 (N2483, N2183, N2349);
  and ginst440 (N2486, N1346, N2374);
  and ginst441 (N2487, N1350, N2375);
  buf ginst442 (N2488, N2185);
  buf ginst443 (N2497, N2188);
  buf ginst444 (N2506, N2191);
  buf ginst445 (N2515, N2194);
  buf ginst446 (N2524, N2197);
  buf ginst447 (N2533, N2200);
  buf ginst448 (N2542, N2203);
  buf ginst449 (N2551, N2206);
  buf ginst450 (N2560, N2185);
  buf ginst451 (N2569, N2188);
  buf ginst452 (N2578, N2191);
  buf ginst453 (N2587, N2194);
  buf ginst454 (N2596, N2197);
  buf ginst455 (N2605, N2200);
  buf ginst456 (N2614, N2203);
  buf ginst457 (N2623, N2206);
  not ginst458 (N2632, N2212);
  and ginst459 (N2633, N1833, N2212);
  not ginst460 (N2634, N2212);
  and ginst461 (N2635, N1833, N2212);
  not ginst462 (N2636, N2212);
  and ginst463 (N2637, N1833, N2212);
  not ginst464 (N2638, N2212);
  and ginst465 (N2639, N1833, N2212);
  not ginst466 (N2640, N2221);
  and ginst467 (N2641, N1824, N2221);
  not ginst468 (N2642, N2221);
  and ginst469 (N2643, N1824, N2221);
  not ginst470 (N2644, N2221);
  and ginst471 (N2645, N1824, N2221);
  not ginst472 (N2646, N2221);
  and ginst473 (N2647, N1824, N2221);
  or ginst474 (N2648, N1870, N2068, N2270);
  nor ginst475 (N2652, N1870, N2068, N2270);
  or ginst476 (N2656, N2417, N2418, N2419);
  or ginst477 (N2659, N2420, N2421, N2422);
  or ginst478 (N2662, N1880, N2078, N2277);
  nor ginst479 (N2666, N1880, N2078, N2277);
  or ginst480 (N2670, N2425, N2426, N2427);
  or ginst481 (N2673, N1885, N2083, N2282);
  nor ginst482 (N2677, N1885, N2083, N2282);
  or ginst483 (N2681, N2430, N2431, N2432);
  or ginst484 (N2684, N1890, N2088, N2287);
  nor ginst485 (N2688, N1890, N2088, N2287);
  or ginst486 (N2692, N2435, N2436, N2437);
  or ginst487 (N2697, N2438, N2439, N2440);
  or ginst488 (N2702, N1900, N2098, N2294);
  nor ginst489 (N2706, N1900, N2098, N2294);
  or ginst490 (N2710, N2443, N2444, N2445);
  or ginst491 (N2715, N1905, N2103, N2299);
  nor ginst492 (N2719, N1905, N2103, N2299);
  or ginst493 (N2723, N2448, N2449, N2450);
  not ginst494 (N2728, N2304);
  not ginst495 (N2729, N2158);
  and ginst496 (N2730, N1562, N2158);
  not ginst497 (N2731, N2158);
  and ginst498 (N2732, N1562, N2158);
  not ginst499 (N2733, N2158);
  and ginst500 (N2734, N1562, N2158);
  not ginst501 (N2735, N2158);
  and ginst502 (N2736, N1562, N2158);
  not ginst503 (N2737, N2158);
  and ginst504 (N2738, N1562, N2158);
  not ginst505 (N2739, N2158);
  and ginst506 (N2740, N1562, N2158);
  not ginst507 (N2741, N2158);
  and ginst508 (N2742, N1562, N2158);
  not ginst509 (N2743, N2158);
  and ginst510 (N2744, N1562, N2158);
  or ginst511 (N2745, N1983, N2376, N2379);
  nor ginst512 (N2746, N1983, N2376, N2379);
  nand ginst513 (N2748, N2316, N2467);
  nand ginst514 (N2749, N2313, N2468);
  nand ginst515 (N2750, N2322, N2469);
  nand ginst516 (N2751, N2319, N2470);
  nand ginst517 (N2754, N2328, N2474);
  nand ginst518 (N2755, N2325, N2475);
  nand ginst519 (N2756, N2334, N2476);
  nand ginst520 (N2757, N2331, N2477);
  and ginst521 (N2758, N1520, N2481);
  and ginst522 (N2761, N1722, N2482);
  and ginst523 (N2764, N1770, N2478);
  or ginst524 (N2768, N1789, N1790, N2486);
  or ginst525 (N2769, N1797, N1798, N2487);
  and ginst526 (N2898, N665, N2633);
  and ginst527 (N2899, N679, N2635);
  and ginst528 (N2900, N686, N2637);
  and ginst529 (N2901, N702, N2639);
  not ginst530 (N2962, N2746);
  nand ginst531 (N2966, N2748, N2749);
  nand ginst532 (N2967, N2750, N2751);
  buf ginst533 (N2970, N2471);
  nand ginst534 (N2973, N2754, N2755);
  nand ginst535 (N2977, N2756, N2757);
  and ginst536 (N2980, N2143, N2471);
  not ginst537 (N2984, N2488);
  not ginst538 (N2985, N2497);
  not ginst539 (N2986, N2506);
  not ginst540 (N2987, N2515);
  not ginst541 (N2988, N2524);
  not ginst542 (N2989, N2533);
  not ginst543 (N2990, N2542);
  not ginst544 (N2991, N2551);
  not ginst545 (N2992, N2488);
  not ginst546 (N2993, N2497);
  not ginst547 (N2994, N2506);
  not ginst548 (N2995, N2515);
  not ginst549 (N2996, N2524);
  not ginst550 (N2997, N2533);
  not ginst551 (N2998, N2542);
  not ginst552 (N2999, N2551);
  not ginst553 (N3000, N2488);
  not ginst554 (N3001, N2497);
  not ginst555 (N3002, N2506);
  not ginst556 (N3003, N2515);
  not ginst557 (N3004, N2524);
  not ginst558 (N3005, N2533);
  not ginst559 (N3006, N2542);
  not ginst560 (N3007, N2551);
  not ginst561 (N3008, N2488);
  not ginst562 (N3009, N2497);
  not ginst563 (N3010, N2506);
  not ginst564 (N3011, N2515);
  not ginst565 (N3012, N2524);
  not ginst566 (N3013, N2533);
  not ginst567 (N3014, N2542);
  not ginst568 (N3015, N2551);
  not ginst569 (N3016, N2488);
  not ginst570 (N3017, N2497);
  not ginst571 (N3018, N2506);
  not ginst572 (N3019, N2515);
  not ginst573 (N3020, N2524);
  not ginst574 (N3021, N2533);
  not ginst575 (N3022, N2542);
  not ginst576 (N3023, N2551);
  not ginst577 (N3024, N2488);
  not ginst578 (N3025, N2497);
  not ginst579 (N3026, N2506);
  not ginst580 (N3027, N2515);
  not ginst581 (N3028, N2524);
  not ginst582 (N3029, N2533);
  not ginst583 (N3030, N2542);
  not ginst584 (N3031, N2551);
  not ginst585 (N3032, N2488);
  not ginst586 (N3033, N2497);
  not ginst587 (N3034, N2506);
  not ginst588 (N3035, N2515);
  not ginst589 (N3036, N2524);
  not ginst590 (N3037, N2533);
  not ginst591 (N3038, N2542);
  not ginst592 (N3039, N2551);
  not ginst593 (N3040, N2488);
  not ginst594 (N3041, N2497);
  not ginst595 (N3042, N2506);
  not ginst596 (N3043, N2515);
  not ginst597 (N3044, N2524);
  not ginst598 (N3045, N2533);
  not ginst599 (N3046, N2542);
  not ginst600 (N3047, N2551);
  not ginst601 (N3048, N2560);
  not ginst602 (N3049, N2569);
  not ginst603 (N3050, N2578);
  not ginst604 (N3051, N2587);
  not ginst605 (N3052, N2596);
  not ginst606 (N3053, N2605);
  not ginst607 (N3054, N2614);
  not ginst608 (N3055, N2623);
  not ginst609 (N3056, N2560);
  not ginst610 (N3057, N2569);
  not ginst611 (N3058, N2578);
  not ginst612 (N3059, N2587);
  not ginst613 (N3060, N2596);
  not ginst614 (N3061, N2605);
  not ginst615 (N3062, N2614);
  not ginst616 (N3063, N2623);
  not ginst617 (N3064, N2560);
  not ginst618 (N3065, N2569);
  not ginst619 (N3066, N2578);
  not ginst620 (N3067, N2587);
  not ginst621 (N3068, N2596);
  not ginst622 (N3069, N2605);
  not ginst623 (N3070, N2614);
  not ginst624 (N3071, N2623);
  not ginst625 (N3072, N2560);
  not ginst626 (N3073, N2569);
  not ginst627 (N3074, N2578);
  not ginst628 (N3075, N2587);
  not ginst629 (N3076, N2596);
  not ginst630 (N3077, N2605);
  not ginst631 (N3078, N2614);
  not ginst632 (N3079, N2623);
  not ginst633 (N3080, N2560);
  not ginst634 (N3081, N2569);
  not ginst635 (N3082, N2578);
  not ginst636 (N3083, N2587);
  not ginst637 (N3084, N2596);
  not ginst638 (N3085, N2605);
  not ginst639 (N3086, N2614);
  not ginst640 (N3087, N2623);
  not ginst641 (N3088, N2560);
  not ginst642 (N3089, N2569);
  not ginst643 (N3090, N2578);
  not ginst644 (N3091, N2587);
  not ginst645 (N3092, N2596);
  not ginst646 (N3093, N2605);
  not ginst647 (N3094, N2614);
  not ginst648 (N3095, N2623);
  not ginst649 (N3096, N2560);
  not ginst650 (N3097, N2569);
  not ginst651 (N3098, N2578);
  not ginst652 (N3099, N2587);
  not ginst653 (N3100, N2596);
  not ginst654 (N3101, N2605);
  not ginst655 (N3102, N2614);
  not ginst656 (N3103, N2623);
  not ginst657 (N3104, N2560);
  not ginst658 (N3105, N2569);
  not ginst659 (N3106, N2578);
  not ginst660 (N3107, N2587);
  not ginst661 (N3108, N2596);
  not ginst662 (N3109, N2605);
  not ginst663 (N3110, N2614);
  not ginst664 (N3111, N2623);
  buf ginst665 (N3112, N2656);
  not ginst666 (N3115, N2656);
  not ginst667 (N3118, N2652);
  and ginst668 (N3119, N1674, N2768);
  buf ginst669 (N3122, N2659);
  not ginst670 (N3125, N2659);
  buf ginst671 (N3128, N2670);
  not ginst672 (N3131, N2670);
  not ginst673 (N3134, N2666);
  buf ginst674 (N3135, N2681);
  not ginst675 (N3138, N2681);
  not ginst676 (N3141, N2677);
  buf ginst677 (N3142, N2692);
  not ginst678 (N3145, N2692);
  not ginst679 (N3148, N2688);
  and ginst680 (N3149, N1678, N2769);
  buf ginst681 (N3152, N2697);
  not ginst682 (N3155, N2697);
  buf ginst683 (N3158, N2710);
  not ginst684 (N3161, N2710);
  not ginst685 (N3164, N2706);
  buf ginst686 (N3165, N2723);
  not ginst687 (N3168, N2723);
  not ginst688 (N3171, N2719);
  and ginst689 (N3172, N1909, N2648);
  and ginst690 (N3175, N1913, N2662);
  and ginst691 (N3178, N1913, N2673);
  and ginst692 (N3181, N1913, N2684);
  and ginst693 (N3184, N1922, N2702);
  and ginst694 (N3187, N1922, N2715);
  not ginst695 (N3190, N2692);
  not ginst696 (N3191, N2697);
  not ginst697 (N3192, N2710);
  not ginst698 (N3193, N2723);
  and ginst699 (N3194, N1459, N2692, N2697, N2710, N2723);
  nand ginst700 (N3195, N2745, N2962);
  not ginst701 (N3196, N2966);
  or ginst702 (N3206, N2145, N2347, N2980);
  and ginst703 (N3207, N2984, N124);
  and ginst704 (N3208, N2985, N159);
  and ginst705 (N3209, N2986, N150);
  and ginst706 (N3210, N2987, N143);
  and ginst707 (N3211, N2988, N137);
  and ginst708 (N3212, N2989, N132);
  and ginst709 (N3213, N2990, N128);
  and ginst710 (N3214, N2991, N125);
  and ginst711 (N3215, N2992, N125);
  and ginst712 (N3216, N655, N2993);
  and ginst713 (N3217, N2994, N159);
  and ginst714 (N3218, N2995, N150);
  and ginst715 (N3219, N2996, N143);
  and ginst716 (N3220, N2997, N137);
  and ginst717 (N3221, N2998, N132);
  and ginst718 (N3222, N2999, N128);
  and ginst719 (N3223, N3000, N128);
  and ginst720 (N3224, N670, N3001);
  and ginst721 (N3225, N655, N3002);
  and ginst722 (N3226, N3003, N159);
  and ginst723 (N3227, N3004, N150);
  and ginst724 (N3228, N3005, N143);
  and ginst725 (N3229, N3006, N137);
  and ginst726 (N3230, N3007, N132);
  and ginst727 (N3231, N3008, N132);
  and ginst728 (N3232, N690, N3009);
  and ginst729 (N3233, N670, N3010);
  and ginst730 (N3234, N655, N3011);
  and ginst731 (N3235, N3012, N159);
  and ginst732 (N3236, N3013, N150);
  and ginst733 (N3237, N3014, N143);
  and ginst734 (N3238, N3015, N137);
  and ginst735 (N3239, N3016, N137);
  and ginst736 (N3240, N706, N3017);
  and ginst737 (N3241, N690, N3018);
  and ginst738 (N3242, N670, N3019);
  and ginst739 (N3243, N655, N3020);
  and ginst740 (N3244, N3021, N159);
  and ginst741 (N3245, N3022, N150);
  and ginst742 (N3246, N3023, N143);
  and ginst743 (N3247, N3024, N143);
  and ginst744 (N3248, N715, N3025);
  and ginst745 (N3249, N706, N3026);
  and ginst746 (N3250, N690, N3027);
  and ginst747 (N3251, N670, N3028);
  and ginst748 (N3252, N655, N3029);
  and ginst749 (N3253, N3030, N159);
  and ginst750 (N3254, N3031, N150);
  and ginst751 (N3255, N3032, N150);
  and ginst752 (N3256, N727, N3033);
  and ginst753 (N3257, N715, N3034);
  and ginst754 (N3258, N706, N3035);
  and ginst755 (N3259, N690, N3036);
  and ginst756 (N3260, N670, N3037);
  and ginst757 (N3261, N655, N3038);
  and ginst758 (N3262, N3039, N159);
  and ginst759 (N3263, N3040, N159);
  and ginst760 (N3264, N740, N3041);
  and ginst761 (N3265, N727, N3042);
  and ginst762 (N3266, N715, N3043);
  and ginst763 (N3267, N706, N3044);
  and ginst764 (N3268, N690, N3045);
  and ginst765 (N3269, N670, N3046);
  and ginst766 (N3270, N655, N3047);
  and ginst767 (N3271, N3048, N283);
  and ginst768 (N3272, N670, N3049);
  and ginst769 (N3273, N690, N3050);
  and ginst770 (N3274, N706, N3051);
  and ginst771 (N3275, N715, N3052);
  and ginst772 (N3276, N727, N3053);
  and ginst773 (N3277, N740, N3054);
  and ginst774 (N3278, N753, N3055);
  and ginst775 (N3279, N3056, N294);
  and ginst776 (N3280, N690, N3057);
  and ginst777 (N3281, N706, N3058);
  and ginst778 (N3282, N715, N3059);
  and ginst779 (N3283, N727, N3060);
  and ginst780 (N3284, N740, N3061);
  and ginst781 (N3285, N753, N3062);
  and ginst782 (N3286, N3063, N283);
  and ginst783 (N3287, N3064, N303);
  and ginst784 (N3288, N706, N3065);
  and ginst785 (N3289, N715, N3066);
  and ginst786 (N3290, N727, N3067);
  and ginst787 (N3291, N740, N3068);
  and ginst788 (N3292, N753, N3069);
  and ginst789 (N3293, N3070, N283);
  and ginst790 (N3294, N3071, N294);
  and ginst791 (N3295, N3072, N311);
  and ginst792 (N3296, N715, N3073);
  and ginst793 (N3297, N727, N3074);
  and ginst794 (N3298, N740, N3075);
  and ginst795 (N3299, N753, N3076);
  and ginst796 (N3300, N3077, N283);
  and ginst797 (N3301, N3078, N294);
  and ginst798 (N3302, N3079, N303);
  and ginst799 (N3303, N3080, N317);
  and ginst800 (N3304, N727, N3081);
  and ginst801 (N3305, N740, N3082);
  and ginst802 (N3306, N753, N3083);
  and ginst803 (N3307, N3084, N283);
  and ginst804 (N3308, N3085, N294);
  and ginst805 (N3309, N3086, N303);
  and ginst806 (N3310, N3087, N311);
  and ginst807 (N3311, N3088, N322);
  and ginst808 (N3312, N740, N3089);
  and ginst809 (N3313, N753, N3090);
  and ginst810 (N3314, N3091, N283);
  and ginst811 (N3315, N3092, N294);
  and ginst812 (N3316, N3093, N303);
  and ginst813 (N3317, N3094, N311);
  and ginst814 (N3318, N3095, N317);
  and ginst815 (N3319, N3096, N326);
  and ginst816 (N3320, N753, N3097);
  and ginst817 (N3321, N3098, N283);
  and ginst818 (N3322, N3099, N294);
  and ginst819 (N3323, N3100, N303);
  and ginst820 (N3324, N3101, N311);
  and ginst821 (N3325, N3102, N317);
  and ginst822 (N3326, N3103, N322);
  and ginst823 (N3327, N3104, N329);
  and ginst824 (N3328, N3105, N283);
  and ginst825 (N3329, N3106, N294);
  and ginst826 (N3330, N3107, N303);
  and ginst827 (N3331, N3108, N311);
  and ginst828 (N3332, N3109, N317);
  and ginst829 (N3333, N3110, N322);
  and ginst830 (N3334, N3111, N326);
  and ginst831 (N3383, N917, N3190, N3191, N3192, N3193);
  buf ginst832 (N3384, N2977);
  and ginst833 (N3387, N1736, N3196);
  and ginst834 (N3388, N2149, N2977);
  and ginst835 (N3389, N1737, N2973);
  nor ginst836 (N3390, N3207, N3208, N3209, N3210, N3211, N3212, N3213, N3214);
  nor ginst837 (N3391, N3215, N3216, N3217, N3218, N3219, N3220, N3221, N3222);
  nor ginst838 (N3392, N3223, N3224, N3225, N3226, N3227, N3228, N3229, N3230);
  nor ginst839 (N3393, N3231, N3232, N3233, N3234, N3235, N3236, N3237, N3238);
  nor ginst840 (N3394, N3239, N3240, N3241, N3242, N3243, N3244, N3245, N3246);
  nor ginst841 (N3395, N3247, N3248, N3249, N3250, N3251, N3252, N3253, N3254);
  nor ginst842 (N3396, N3255, N3256, N3257, N3258, N3259, N3260, N3261, N3262);
  nor ginst843 (N3397, N3263, N3264, N3265, N3266, N3267, N3268, N3269, N3270);
  nor ginst844 (N3398, N3271, N3272, N3273, N3274, N3275, N3276, N3277, N3278);
  nor ginst845 (N3399, N3279, N3280, N3281, N3282, N3283, N3284, N3285, N3286);
  nor ginst846 (N3400, N3287, N3288, N3289, N3290, N3291, N3292, N3293, N3294);
  nor ginst847 (N3401, N3295, N3296, N3297, N3298, N3299, N3300, N3301, N3302);
  nor ginst848 (N3402, N3303, N3304, N3305, N3306, N3307, N3308, N3309, N3310);
  nor ginst849 (N3403, N3311, N3312, N3313, N3314, N3315, N3316, N3317, N3318);
  nor ginst850 (N3404, N3319, N3320, N3321, N3322, N3323, N3324, N3325, N3326);
  nor ginst851 (N3405, N3327, N3328, N3329, N3330, N3331, N3332, N3333, N3334);
  and ginst852 (N3406, N2641, N3206);
  and ginst853 (N3407, N2648, N3112, N169);
  and ginst854 (N3410, N2648, N3115, N179);
  and ginst855 (N3413, N2652, N3115, N190);
  and ginst856 (N3414, N2652, N3112, N200);
  or ginst857 (N3415, N1875, N2073, N3119);
  nor ginst858 (N3419, N1875, N2073, N3119);
  and ginst859 (N3423, N2662, N3128, N169);
  and ginst860 (N3426, N2662, N3131, N179);
  and ginst861 (N3429, N2666, N3131, N190);
  and ginst862 (N3430, N2666, N3128, N200);
  and ginst863 (N3431, N2673, N3135, N169);
  and ginst864 (N3434, N2673, N3138, N179);
  and ginst865 (N3437, N2677, N3138, N190);
  and ginst866 (N3438, N2677, N3135, N200);
  and ginst867 (N3439, N2684, N3142, N169);
  and ginst868 (N3442, N2684, N3145, N179);
  and ginst869 (N3445, N2688, N3145, N190);
  and ginst870 (N3446, N2688, N3142, N200);
  or ginst871 (N3447, N1895, N2093, N3149);
  nor ginst872 (N3451, N1895, N2093, N3149);
  and ginst873 (N3455, N2702, N3158, N169);
  and ginst874 (N3458, N2702, N3161, N179);
  and ginst875 (N3461, N2706, N3161, N190);
  and ginst876 (N3462, N2706, N3158, N200);
  and ginst877 (N3463, N2715, N3165, N169);
  and ginst878 (N3466, N2715, N3168, N179);
  and ginst879 (N3469, N2719, N3168, N190);
  and ginst880 (N3470, N2719, N3165, N200);
  or ginst881 (N3471, N3194, N3383);
  buf ginst882 (N3472, N2967);
  buf ginst883 (N3475, N2970);
  buf ginst884 (N3478, N2967);
  buf ginst885 (N3481, N2970);
  buf ginst886 (N3484, N2973);
  buf ginst887 (N3487, N2973);
  buf ginst888 (N3490, N3172);
  buf ginst889 (N3493, N3172);
  buf ginst890 (N3496, N3175);
  buf ginst891 (N3499, N3175);
  buf ginst892 (N3502, N3178);
  buf ginst893 (N3505, N3178);
  buf ginst894 (N3508, N3181);
  buf ginst895 (N3511, N3181);
  buf ginst896 (N3514, N3184);
  buf ginst897 (N3517, N3184);
  buf ginst898 (N3520, N3187);
  buf ginst899 (N3523, N3187);
  nor ginst900 (N3534, N2350, N3387);
  or ginst901 (N3535, N2151, N2351, N3388);
  nor ginst902 (N3536, N1966, N3389);
  and ginst903 (N3537, N2209, N3390);
  and ginst904 (N3538, N2210, N3398);
  and ginst905 (N3539, N1842, N3391);
  and ginst906 (N3540, N1369, N3399);
  and ginst907 (N3541, N1843, N3392);
  and ginst908 (N3542, N1369, N3400);
  and ginst909 (N3543, N1844, N3393);
  and ginst910 (N3544, N1369, N3401);
  and ginst911 (N3545, N1845, N3394);
  and ginst912 (N3546, N1369, N3402);
  and ginst913 (N3547, N1846, N3395);
  and ginst914 (N3548, N1369, N3403);
  and ginst915 (N3549, N1847, N3396);
  and ginst916 (N3550, N1369, N3404);
  and ginst917 (N3551, N1848, N3397);
  and ginst918 (N3552, N1369, N3405);
  or ginst919 (N3557, N3118, N3413, N3414);
  or ginst920 (N3568, N3134, N3429, N3430);
  or ginst921 (N3573, N3141, N3437, N3438);
  or ginst922 (N3578, N3148, N3445, N3446);
  or ginst923 (N3589, N3164, N3461, N3462);
  or ginst924 (N3594, N3171, N3469, N3470);
  and ginst925 (N3605, N2728, N3471);
  not ginst926 (N3626, N3478);
  not ginst927 (N3627, N3481);
  not ginst928 (N3628, N3487);
  not ginst929 (N3629, N3484);
  not ginst930 (N3630, N3472);
  not ginst931 (N3631, N3475);
  and ginst932 (N3632, N2152, N3536);
  and ginst933 (N3633, N2155, N3534);
  or ginst934 (N3634, N2398, N3537, N3538);
  or ginst935 (N3635, N3539, N3540);
  or ginst936 (N3636, N3541, N3542);
  or ginst937 (N3637, N3543, N3544);
  or ginst938 (N3638, N3545, N3546);
  or ginst939 (N3639, N3547, N3548);
  or ginst940 (N3640, N3549, N3550);
  or ginst941 (N3641, N3551, N3552);
  and ginst942 (N3642, N2643, N3535);
  or ginst943 (N3643, N3407, N3410);
  nor ginst944 (N3644, N3407, N3410);
  and ginst945 (N3645, N3122, N3415, N169);
  and ginst946 (N3648, N3125, N3415, N179);
  and ginst947 (N3651, N3125, N3419, N190);
  and ginst948 (N3652, N3122, N3419, N200);
  not ginst949 (N3653, N3419);
  or ginst950 (N3654, N3423, N3426);
  nor ginst951 (N3657, N3423, N3426);
  or ginst952 (N3658, N3431, N3434);
  nor ginst953 (N3661, N3431, N3434);
  or ginst954 (N3662, N3439, N3442);
  nor ginst955 (N3663, N3439, N3442);
  and ginst956 (N3664, N3152, N3447, N169);
  and ginst957 (N3667, N3155, N3447, N179);
  and ginst958 (N3670, N3155, N3451, N190);
  and ginst959 (N3671, N3152, N3451, N200);
  not ginst960 (N3672, N3451);
  or ginst961 (N3673, N3455, N3458);
  nor ginst962 (N3676, N3455, N3458);
  or ginst963 (N3677, N3463, N3466);
  nor ginst964 (N3680, N3463, N3466);
  not ginst965 (N3681, N3493);
  and ginst966 (N3682, N1909, N3415);
  not ginst967 (N3685, N3496);
  not ginst968 (N3686, N3499);
  not ginst969 (N3687, N3502);
  not ginst970 (N3688, N3505);
  not ginst971 (N3689, N3511);
  and ginst972 (N3690, N1922, N3447);
  not ginst973 (N3693, N3517);
  not ginst974 (N3694, N3520);
  not ginst975 (N3695, N3523);
  not ginst976 (N3696, N3514);
  buf ginst977 (N3697, N3384);
  buf ginst978 (N3700, N3384);
  not ginst979 (N3703, N3490);
  not ginst980 (N3704, N3508);
  nand ginst981 (N3705, N3475, N3630);
  nand ginst982 (N3706, N3472, N3631);
  nand ginst983 (N3707, N3481, N3626);
  nand ginst984 (N3708, N3478, N3627);
  or ginst985 (N3711, N2352, N2353, N3632);
  or ginst986 (N3712, N2354, N2355, N3633);
  and ginst987 (N3713, N2632, N3634);
  and ginst988 (N3714, N2634, N3635);
  and ginst989 (N3715, N2636, N3636);
  and ginst990 (N3716, N2638, N3637);
  and ginst991 (N3717, N2640, N3638);
  and ginst992 (N3718, N2642, N3639);
  and ginst993 (N3719, N2644, N3640);
  and ginst994 (N3720, N2646, N3641);
  and ginst995 (N3721, N3557, N3644);
  or ginst996 (N3731, N3651, N3652, N3653);
  and ginst997 (N3734, N3568, N3657);
  and ginst998 (N3740, N3573, N3661);
  and ginst999 (N3743, N3578, N3663);
  or ginst1000 (N3753, N3670, N3671, N3672);
  and ginst1001 (N3756, N3589, N3676);
  and ginst1002 (N3762, N3594, N3680);
  not ginst1003 (N3765, N3643);
  not ginst1004 (N3766, N3662);
  nand ginst1005 (N3773, N3705, N3706);
  nand ginst1006 (N3774, N3707, N3708);
  nand ginst1007 (N3775, N3628, N3700);
  not ginst1008 (N3776, N3700);
  nand ginst1009 (N3777, N3629, N3697);
  not ginst1010 (N3778, N3697);
  and ginst1011 (N3779, N2645, N3712);
  and ginst1012 (N3780, N2647, N3711);
  or ginst1013 (N3786, N3645, N3648);
  nor ginst1014 (N3789, N3645, N3648);
  or ginst1015 (N3800, N3664, N3667);
  nor ginst1016 (N3803, N3664, N3667);
  and ginst1017 (N3809, N1917, N3654);
  and ginst1018 (N3812, N1917, N3658);
  and ginst1019 (N3815, N1926, N3673);
  and ginst1020 (N3818, N1926, N3677);
  buf ginst1021 (N3821, N3682);
  buf ginst1022 (N3824, N3682);
  buf ginst1023 (N3827, N3690);
  buf ginst1024 (N3830, N3690);
  nand ginst1025 (N3833, N3773, N3774);
  nand ginst1026 (N3834, N3487, N3776);
  nand ginst1027 (N3835, N3484, N3778);
  and ginst1028 (N3838, N3731, N3789);
  and ginst1029 (N3845, N3753, N3803);
  buf ginst1030 (N3850, N3721);
  buf ginst1031 (N3855, N3734);
  buf ginst1032 (N3858, N3740);
  buf ginst1033 (N3861, N3743);
  buf ginst1034 (N3865, N3756);
  buf ginst1035 (N3868, N3762);
  nand ginst1036 (N3884, N3775, N3834);
  nand ginst1037 (N3885, N3777, N3835);
  nand ginst1038 (N3894, N3721, N3786);
  nand ginst1039 (N3895, N3743, N3800);
  not ginst1040 (N3898, N3821);
  not ginst1041 (N3899, N3824);
  not ginst1042 (N3906, N3830);
  not ginst1043 (N3911, N3827);
  and ginst1044 (N3912, N1912, N3786);
  buf ginst1045 (N3913, N3812);
  and ginst1046 (N3916, N1917, N3800);
  buf ginst1047 (N3917, N3818);
  not ginst1048 (N3920, N3809);
  buf ginst1049 (N3921, N3818);
  not ginst1050 (N3924, N3884);
  not ginst1051 (N3925, N3885);
  and ginst1052 (N3926, N3721, N3734, N3740, N3838);
  nand ginst1053 (N3930, N3654, N3721, N3838);
  nand ginst1054 (N3931, N3658, N3721, N3734, N3838);
  and ginst1055 (N3932, N3743, N3756, N3762, N3845);
  nand ginst1056 (N3935, N3673, N3743, N3845);
  nand ginst1057 (N3936, N3677, N3743, N3756, N3845);
  buf ginst1058 (N3937, N3838);
  buf ginst1059 (N3940, N3845);
  not ginst1060 (N3947, N3912);
  not ginst1061 (N3948, N3916);
  buf ginst1062 (N3950, N3850);
  buf ginst1063 (N3953, N3850);
  buf ginst1064 (N3956, N3855);
  buf ginst1065 (N3959, N3855);
  buf ginst1066 (N3962, N3858);
  buf ginst1067 (N3965, N3858);
  buf ginst1068 (N3968, N3861);
  buf ginst1069 (N3971, N3861);
  buf ginst1070 (N3974, N3865);
  buf ginst1071 (N3977, N3865);
  buf ginst1072 (N3980, N3868);
  buf ginst1073 (N3983, N3868);
  nand ginst1074 (N3987, N3924, N3925);
  nand ginst1075 (N3992, N3765, N3894, N3930, N3931);
  nand ginst1076 (N3996, N3766, N3895, N3935, N3936);
  not ginst1077 (N4013, N3921);
  and ginst1078 (N4028, N3926, N3932);
  nand ginst1079 (N4029, N3681, N3953);
  nand ginst1080 (N4030, N3686, N3959);
  nand ginst1081 (N4031, N3688, N3965);
  nand ginst1082 (N4032, N3689, N3971);
  nand ginst1083 (N4033, N3693, N3977);
  nand ginst1084 (N4034, N3695, N3983);
  buf ginst1085 (N4035, N3926);
  not ginst1086 (N4042, N3953);
  not ginst1087 (N4043, N3956);
  nand ginst1088 (N4044, N3685, N3956);
  not ginst1089 (N4045, N3959);
  not ginst1090 (N4046, N3962);
  nand ginst1091 (N4047, N3687, N3962);
  not ginst1092 (N4048, N3965);
  not ginst1093 (N4049, N3971);
  not ginst1094 (N4050, N3977);
  not ginst1095 (N4051, N3980);
  nand ginst1096 (N4052, N3694, N3980);
  not ginst1097 (N4053, N3983);
  not ginst1098 (N4054, N3974);
  nand ginst1099 (N4055, N3696, N3974);
  and ginst1100 (N4056, N2304, N3932);
  not ginst1101 (N4057, N3950);
  nand ginst1102 (N4058, N3703, N3950);
  buf ginst1103 (N4059, N3937);
  buf ginst1104 (N4062, N3937);
  not ginst1105 (N4065, N3968);
  nand ginst1106 (N4066, N3704, N3968);
  buf ginst1107 (N4067, N3940);
  buf ginst1108 (N4070, N3940);
  nand ginst1109 (N4073, N3926, N3996);
  not ginst1110 (N4074, N3992);
  nand ginst1111 (N4075, N3493, N4042);
  nand ginst1112 (N4076, N3499, N4045);
  nand ginst1113 (N4077, N3505, N4048);
  nand ginst1114 (N4078, N3511, N4049);
  nand ginst1115 (N4079, N3517, N4050);
  nand ginst1116 (N4080, N3523, N4053);
  nand ginst1117 (N4085, N3496, N4043);
  nand ginst1118 (N4086, N3502, N4046);
  nand ginst1119 (N4088, N3520, N4051);
  nand ginst1120 (N4090, N3514, N4054);
  and ginst1121 (N4091, N1926, N3996);
  or ginst1122 (N4094, N3605, N4056);
  nand ginst1123 (N4098, N3490, N4057);
  nand ginst1124 (N4101, N3508, N4065);
  and ginst1125 (N4104, N4073, N4074);
  nand ginst1126 (N4105, N4029, N4075);
  nand ginst1127 (N4106, N3899, N4062);
  nand ginst1128 (N4107, N4030, N4076);
  nand ginst1129 (N4108, N4031, N4077);
  nand ginst1130 (N4109, N4032, N4078);
  nand ginst1131 (N4110, N3906, N4070);
  nand ginst1132 (N4111, N4033, N4079);
  nand ginst1133 (N4112, N4034, N4080);
  not ginst1134 (N4113, N4059);
  nand ginst1135 (N4114, N3898, N4059);
  not ginst1136 (N4115, N4062);
  nand ginst1137 (N4116, N4044, N4085);
  nand ginst1138 (N4119, N4047, N4086);
  not ginst1139 (N4122, N4070);
  nand ginst1140 (N4123, N4052, N4088);
  not ginst1141 (N4126, N4067);
  nand ginst1142 (N4127, N3911, N4067);
  nand ginst1143 (N4128, N4055, N4090);
  nand ginst1144 (N4139, N4058, N4098);
  nand ginst1145 (N4142, N4066, N4101);
  not ginst1146 (N4145, N4104);
  not ginst1147 (N4146, N4105);
  nand ginst1148 (N4147, N3824, N4115);
  not ginst1149 (N4148, N4107);
  not ginst1150 (N4149, N4108);
  not ginst1151 (N4150, N4109);
  nand ginst1152 (N4151, N3830, N4122);
  not ginst1153 (N4152, N4111);
  not ginst1154 (N4153, N4112);
  nand ginst1155 (N4154, N3821, N4113);
  nand ginst1156 (N4161, N3827, N4126);
  buf ginst1157 (N4167, N4091);
  buf ginst1158 (N4174, N4094);
  buf ginst1159 (N4182, N4091);
  and ginst1160 (N4186, N4094, N330);
  and ginst1161 (N4189, N2230, N4146);
  nand ginst1162 (N4190, N4106, N4147);
  and ginst1163 (N4191, N2232, N4148);
  and ginst1164 (N4192, N2233, N4149);
  and ginst1165 (N4193, N2234, N4150);
  nand ginst1166 (N4194, N4110, N4151);
  and ginst1167 (N4195, N2236, N4152);
  and ginst1168 (N4196, N2237, N4153);
  nand ginst1169 (N4197, N4114, N4154);
  buf ginst1170 (N4200, N4116);
  buf ginst1171 (N4203, N4116);
  buf ginst1172 (N4209, N4119);
  buf ginst1173 (N4213, N4119);
  nand ginst1174 (N4218, N4127, N4161);
  buf ginst1175 (N4223, N4123);
  and ginst1176 (N4238, N3917, N4128);
  not ginst1177 (N4239, N4139);
  not ginst1178 (N4241, N4142);
  and ginst1179 (N4242, N4123, N330);
  buf ginst1180 (N4247, N4128);
  nor ginst1181 (N4251, N2898, N3713, N4189);
  not ginst1182 (N4252, N4190);
  nor ginst1183 (N4253, N2900, N3715, N4191);
  nor ginst1184 (N4254, N2901, N3716, N4192);
  nor ginst1185 (N4255, N3406, N3717, N4193);
  not ginst1186 (N4256, N4194);
  nor ginst1187 (N4257, N3719, N3779, N4195);
  nor ginst1188 (N4258, N3720, N3780, N4196);
  and ginst1189 (N4283, N4035, N4167);
  and ginst1190 (N4284, N4035, N4174);
  or ginst1191 (N4287, N3815, N4238);
  not ginst1192 (N4291, N4186);
  not ginst1193 (N4295, N4167);
  buf ginst1194 (N4296, N4167);
  not ginst1195 (N4299, N4182);
  and ginst1196 (N4303, N2231, N4252);
  and ginst1197 (N4304, N2235, N4256);
  buf ginst1198 (N4305, N4197);
  or ginst1199 (N4310, N3992, N4283);
  and ginst1200 (N4316, N4174, N4203, N4213);
  and ginst1201 (N4317, N4174, N4209);
  and ginst1202 (N4318, N4128, N4218, N4223);
  and ginst1203 (N4319, N4128, N4223);
  and ginst1204 (N4322, N4167, N4209);
  nand ginst1205 (N4325, N3913, N4203);
  nand ginst1206 (N4326, N4167, N4203, N4213);
  nand ginst1207 (N4327, N3815, N4218);
  nand ginst1208 (N4328, N3917, N4128, N4218);
  nand ginst1209 (N4329, N4013, N4247);
  not ginst1210 (N4330, N4247);
  and ginst1211 (N4331, N4094, N4295, N330);
  and ginst1212 (N4335, N2730, N4251);
  and ginst1213 (N4338, N2734, N4253);
  and ginst1214 (N4341, N2736, N4254);
  and ginst1215 (N4344, N2738, N4255);
  and ginst1216 (N4347, N2742, N4257);
  and ginst1217 (N4350, N2744, N4258);
  buf ginst1218 (N4353, N4197);
  buf ginst1219 (N4356, N4203);
  buf ginst1220 (N4359, N4209);
  buf ginst1221 (N4362, N4218);
  buf ginst1222 (N4365, N4242);
  buf ginst1223 (N4368, N4242);
  and ginst1224 (N4371, N4223, N4223);
  nor ginst1225 (N4376, N2899, N3714, N4303);
  nor ginst1226 (N4377, N3642, N3718, N4304);
  and ginst1227 (N4387, N4317, N330);
  and ginst1228 (N4390, N4318, N330);
  nand ginst1229 (N4393, N3921, N4330);
  buf ginst1230 (N4398, N4287);
  buf ginst1231 (N4413, N4284);
  nand ginst1232 (N4416, N3920, N4325, N4326);
  or ginst1233 (N4421, N3812, N4322);
  nand ginst1234 (N4427, N3948, N4327, N4328);
  buf ginst1235 (N4430, N4287);
  and ginst1236 (N4435, N4316, N330);
  or ginst1237 (N4442, N4296, N4331);
  and ginst1238 (N4443, N4174, N4203, N4213, N4305);
  nand ginst1239 (N4446, N3809, N4305);
  nand ginst1240 (N4447, N3913, N4200, N4305);
  nand ginst1241 (N4448, N4167, N4200, N4213, N4305);
  not ginst1242 (N4452, N4356);
  nand ginst1243 (N4458, N4329, N4393);
  not ginst1244 (N4461, N4365);
  not ginst1245 (N4462, N4368);
  nand ginst1246 (N4463, N1460, N4371);
  not ginst1247 (N4464, N4371);
  buf ginst1248 (N4465, N4310);
  nor ginst1249 (N4468, N4296, N4331);
  and ginst1250 (N4472, N2732, N4376);
  and ginst1251 (N4475, N2740, N4377);
  buf ginst1252 (N4479, N4310);
  not ginst1253 (N4484, N4353);
  not ginst1254 (N4486, N4359);
  nand ginst1255 (N4487, N4299, N4359);
  not ginst1256 (N4491, N4362);
  and ginst1257 (N4493, N4319, N330);
  not ginst1258 (N4496, N4398);
  and ginst1259 (N4497, N4287, N4398);
  and ginst1260 (N4498, N1769, N4442);
  nand ginst1261 (N4503, N3947, N4446, N4447, N4448);
  not ginst1262 (N4506, N4413);
  not ginst1263 (N4507, N4435);
  not ginst1264 (N4508, N4421);
  nand ginst1265 (N4509, N4421, N4452);
  not ginst1266 (N4510, N4427);
  nand ginst1267 (N4511, N4241, N4427);
  nand ginst1268 (N4515, N965, N4464);
  not ginst1269 (N4526, N4416);
  nand ginst1270 (N4527, N4416, N4484);
  nand ginst1271 (N4528, N4182, N4486);
  not ginst1272 (N4529, N4430);
  nand ginst1273 (N4530, N4430, N4491);
  buf ginst1274 (N4531, N4387);
  buf ginst1275 (N4534, N4387);
  buf ginst1276 (N4537, N4390);
  buf ginst1277 (N4540, N4390);
  and ginst1278 (N4545, N4319, N4496, N330);
  and ginst1279 (N4549, N4443, N330);
  nand ginst1280 (N4552, N4356, N4508);
  nand ginst1281 (N4555, N4142, N4510);
  not ginst1282 (N4558, N4493);
  nand ginst1283 (N4559, N4463, N4515);
  not ginst1284 (N4562, N4465);
  and ginst1285 (N4563, N4310, N4465);
  buf ginst1286 (N4564, N4468);
  not ginst1287 (N4568, N4479);
  buf ginst1288 (N4569, N4443);
  nand ginst1289 (N4572, N4353, N4526);
  nand ginst1290 (N4573, N4362, N4529);
  nand ginst1291 (N4576, N4487, N4528);
  buf ginst1292 (N4581, N4458);
  buf ginst1293 (N4584, N4458);
  or ginst1294 (N4587, N2758, N2761, N4498);
  nor ginst1295 (N4588, N2758, N2761, N4498);
  or ginst1296 (N4589, N4497, N4545);
  nand ginst1297 (N4593, N4509, N4552);
  not ginst1298 (N4596, N4531);
  not ginst1299 (N4597, N4534);
  nand ginst1300 (N4599, N4511, N4555);
  not ginst1301 (N4602, N4537);
  not ginst1302 (N4603, N4540);
  and ginst1303 (N4608, N4284, N4562, N330);
  buf ginst1304 (N4613, N4503);
  buf ginst1305 (N4616, N4503);
  nand ginst1306 (N4619, N4527, N4572);
  nand ginst1307 (N4623, N4530, N4573);
  not ginst1308 (N4628, N4588);
  nand ginst1309 (N4629, N4506, N4569);
  not ginst1310 (N4630, N4569);
  not ginst1311 (N4635, N4576);
  nand ginst1312 (N4636, N4291, N4576);
  not ginst1313 (N4640, N4581);
  nand ginst1314 (N4641, N4461, N4581);
  not ginst1315 (N4642, N4584);
  nand ginst1316 (N4643, N4462, N4584);
  nor ginst1317 (N4644, N4563, N4608);
  and ginst1318 (N4647, N2128, N4559);
  and ginst1319 (N4650, N2743, N4559);
  buf ginst1320 (N4656, N4549);
  buf ginst1321 (N4659, N4549);
  buf ginst1322 (N4664, N4564);
  and ginst1323 (N4667, N4587, N4628);
  nand ginst1324 (N4668, N4413, N4630);
  not ginst1325 (N4669, N4616);
  nand ginst1326 (N4670, N4239, N4616);
  not ginst1327 (N4673, N4619);
  nand ginst1328 (N4674, N4507, N4619);
  nand ginst1329 (N4675, N4186, N4635);
  not ginst1330 (N4676, N4623);
  nand ginst1331 (N4677, N4558, N4623);
  nand ginst1332 (N4678, N4365, N4640);
  nand ginst1333 (N4679, N4368, N4642);
  not ginst1334 (N4687, N4613);
  nand ginst1335 (N4688, N4568, N4613);
  buf ginst1336 (N4691, N4593);
  buf ginst1337 (N4694, N4593);
  buf ginst1338 (N4697, N4599);
  buf ginst1339 (N4700, N4599);
  nand ginst1340 (N4704, N4629, N4668);
  nand ginst1341 (N4705, N4139, N4669);
  not ginst1342 (N4706, N4656);
  not ginst1343 (N4707, N4659);
  nand ginst1344 (N4708, N4435, N4673);
  nand ginst1345 (N4711, N4636, N4675);
  nand ginst1346 (N4716, N4493, N4676);
  nand ginst1347 (N4717, N4641, N4678);
  nand ginst1348 (N4721, N4643, N4679);
  buf ginst1349 (N4722, N4644);
  not ginst1350 (N4726, N4664);
  or ginst1351 (N4727, N4350, N4647, N4650);
  nor ginst1352 (N4730, N4350, N4647, N4650);
  nand ginst1353 (N4733, N4479, N4687);
  nand ginst1354 (N4740, N4670, N4705);
  nand ginst1355 (N4743, N4674, N4708);
  not ginst1356 (N4747, N4691);
  nand ginst1357 (N4748, N4596, N4691);
  not ginst1358 (N4749, N4694);
  nand ginst1359 (N4750, N4597, N4694);
  not ginst1360 (N4753, N4697);
  nand ginst1361 (N4754, N4602, N4697);
  not ginst1362 (N4755, N4700);
  nand ginst1363 (N4756, N4603, N4700);
  nand ginst1364 (N4757, N4677, N4716);
  nand ginst1365 (N4769, N4688, N4733);
  and ginst1366 (N4772, N4704, N330);
  not ginst1367 (N4775, N4721);
  not ginst1368 (N4778, N4730);
  nand ginst1369 (N4786, N4531, N4747);
  nand ginst1370 (N4787, N4534, N4749);
  nand ginst1371 (N4788, N4537, N4753);
  nand ginst1372 (N4789, N4540, N4755);
  and ginst1373 (N4794, N2124, N4711);
  and ginst1374 (N4797, N2735, N4711);
  and ginst1375 (N4800, N2127, N4717);
  buf ginst1376 (N4805, N4722);
  and ginst1377 (N4808, N4468, N4717);
  buf ginst1378 (N4812, N4727);
  and ginst1379 (N4815, N4727, N4778);
  not ginst1380 (N4816, N4769);
  not ginst1381 (N4817, N4772);
  nand ginst1382 (N4818, N4748, N4786);
  nand ginst1383 (N4822, N4750, N4787);
  nand ginst1384 (N4823, N4754, N4788);
  nand ginst1385 (N4826, N4756, N4789);
  nand ginst1386 (N4829, N4726, N4775);
  not ginst1387 (N4830, N4775);
  and ginst1388 (N4831, N2122, N4743);
  and ginst1389 (N4838, N2126, N4757);
  buf ginst1390 (N4844, N4740);
  buf ginst1391 (N4847, N4740);
  buf ginst1392 (N4850, N4743);
  buf ginst1393 (N4854, N4757);
  nand ginst1394 (N4859, N4772, N4816);
  nand ginst1395 (N4860, N4769, N4817);
  not ginst1396 (N4868, N4826);
  not ginst1397 (N4870, N4805);
  not ginst1398 (N4872, N4808);
  nand ginst1399 (N4873, N4664, N4830);
  or ginst1400 (N4876, N4341, N4794, N4797);
  nor ginst1401 (N4880, N4341, N4794, N4797);
  not ginst1402 (N4885, N4812);
  not ginst1403 (N4889, N4822);
  nand ginst1404 (N4895, N4859, N4860);
  not ginst1405 (N4896, N4844);
  nand ginst1406 (N4897, N4706, N4844);
  not ginst1407 (N4898, N4847);
  nand ginst1408 (N4899, N4707, N4847);
  nor ginst1409 (N4900, N4564, N4868);
  and ginst1410 (N4901, N4564, N4717, N4757, N4823);
  not ginst1411 (N4902, N4850);
  not ginst1412 (N4904, N4854);
  nand ginst1413 (N4905, N4854, N4872);
  nand ginst1414 (N4906, N4829, N4873);
  and ginst1415 (N4907, N2123, N4818);
  and ginst1416 (N4913, N2125, N4823);
  and ginst1417 (N4916, N4644, N4818);
  not ginst1418 (N4920, N4880);
  and ginst1419 (N4921, N2184, N4895);
  nand ginst1420 (N4924, N4656, N4896);
  nand ginst1421 (N4925, N4659, N4898);
  or ginst1422 (N4926, N4900, N4901);
  nand ginst1423 (N4928, N4870, N4889);
  not ginst1424 (N4929, N4889);
  nand ginst1425 (N4930, N4808, N4904);
  not ginst1426 (N4931, N4906);
  buf ginst1427 (N4937, N4876);
  buf ginst1428 (N4940, N4876);
  and ginst1429 (N4944, N4876, N4920);
  nand ginst1430 (N4946, N4897, N4924);
  nand ginst1431 (N4949, N4899, N4925);
  nand ginst1432 (N4950, N4902, N4916);
  not ginst1433 (N4951, N4916);
  nand ginst1434 (N4952, N4805, N4929);
  nand ginst1435 (N4953, N4905, N4930);
  and ginst1436 (N4954, N2737, N4926);
  and ginst1437 (N4957, N2741, N4931);
  or ginst1438 (N4964, N2483, N2764, N4921);
  nor ginst1439 (N4965, N2483, N2764, N4921);
  not ginst1440 (N4968, N4949);
  nand ginst1441 (N4969, N4850, N4951);
  nand ginst1442 (N4970, N4928, N4952);
  and ginst1443 (N4973, N2739, N4953);
  not ginst1444 (N4978, N4937);
  not ginst1445 (N4979, N4940);
  not ginst1446 (N4980, N4965);
  nor ginst1447 (N4981, N4722, N4968);
  and ginst1448 (N4982, N4722, N4743, N4818, N4946);
  nand ginst1449 (N4983, N4950, N4969);
  not ginst1450 (N4984, N4970);
  and ginst1451 (N4985, N2121, N4946);
  or ginst1452 (N4988, N4344, N4913, N4954);
  nor ginst1453 (N4991, N4344, N4913, N4954);
  or ginst1454 (N4996, N4347, N4800, N4957);
  nor ginst1455 (N4999, N4347, N4800, N4957);
  and ginst1456 (N5002, N4964, N4980);
  or ginst1457 (N5007, N4981, N4982);
  and ginst1458 (N5010, N2731, N4983);
  and ginst1459 (N5013, N2733, N4984);
  or ginst1460 (N5018, N4475, N4838, N4973);
  nor ginst1461 (N5021, N4475, N4838, N4973);
  not ginst1462 (N5026, N4991);
  not ginst1463 (N5029, N4999);
  and ginst1464 (N5030, N2729, N5007);
  buf ginst1465 (N5039, N4996);
  buf ginst1466 (N5042, N4988);
  and ginst1467 (N5045, N4988, N5026);
  not ginst1468 (N5046, N5021);
  and ginst1469 (N5047, N4996, N5029);
  or ginst1470 (N5050, N4472, N4831, N5010);
  nor ginst1471 (N5055, N4472, N4831, N5010);
  or ginst1472 (N5058, N4338, N4907, N5013);
  nor ginst1473 (N5061, N4338, N4907, N5013);
  and ginst1474 (N5066, N4730, N4991, N4999, N5021);
  buf ginst1475 (N5070, N5018);
  and ginst1476 (N5078, N5018, N5046);
  or ginst1477 (N5080, N4335, N4985, N5030);
  nor ginst1478 (N5085, N4335, N4985, N5030);
  nand ginst1479 (N5094, N4885, N5039);
  not ginst1480 (N5095, N5039);
  not ginst1481 (N5097, N5042);
  and ginst1482 (N5102, N5050, N5050);
  not ginst1483 (N5103, N5061);
  nand ginst1484 (N5108, N4812, N5095);
  not ginst1485 (N5109, N5070);
  nand ginst1486 (N5110, N5070, N5097);
  buf ginst1487 (N5111, N5058);
  and ginst1488 (N5114, N1461, N5050);
  buf ginst1489 (N5117, N5050);
  and ginst1490 (N5120, N5080, N5080);
  and ginst1491 (N5121, N5058, N5103);
  nand ginst1492 (N5122, N5094, N5108);
  nand ginst1493 (N5125, N5042, N5109);
  and ginst1494 (N5128, N1461, N5080);
  and ginst1495 (N5133, N4880, N5055, N5061, N5085);
  and ginst1496 (N5136, N1464, N5055, N5085);
  buf ginst1497 (N5139, N5080);
  nand ginst1498 (N5145, N5110, N5125);
  buf ginst1499 (N5151, N5111);
  buf ginst1500 (N5154, N5111);
  not ginst1501 (N5159, N5117);
  buf ginst1502 (N5160, N5114);
  buf ginst1503 (N5163, N5114);
  and ginst1504 (N5166, N5066, N5133);
  and ginst1505 (N5173, N5066, N5133);
  buf ginst1506 (N5174, N5122);
  buf ginst1507 (N5177, N5122);
  not ginst1508 (N5182, N5139);
  nand ginst1509 (N5183, N5139, N5159);
  buf ginst1510 (N5184, N5128);
  buf ginst1511 (N5188, N5128);
  not ginst1512 (N5192, N5166);
  nor ginst1513 (N5193, N5136, N5173);
  nand ginst1514 (N5196, N4978, N5151);
  not ginst1515 (N5197, N5151);
  nand ginst1516 (N5198, N4979, N5154);
  not ginst1517 (N5199, N5154);
  not ginst1518 (N5201, N5160);
  not ginst1519 (N5203, N5163);
  buf ginst1520 (N5205, N5145);
  buf ginst1521 (N5209, N5145);
  nand ginst1522 (N5212, N5117, N5182);
  and ginst1523 (N5215, N5193, N213);
  not ginst1524 (N5217, N5174);
  not ginst1525 (N5219, N5177);
  nand ginst1526 (N5220, N4937, N5197);
  nand ginst1527 (N5221, N4940, N5199);
  not ginst1528 (N5222, N5184);
  nand ginst1529 (N5223, N5184, N5201);
  nand ginst1530 (N5224, N5188, N5203);
  not ginst1531 (N5225, N5188);
  nand ginst1532 (N5228, N5183, N5212);
  not ginst1533 (N5231, N5215);
  nand ginst1534 (N5232, N5205, N5217);
  not ginst1535 (N5233, N5205);
  nand ginst1536 (N5234, N5209, N5219);
  not ginst1537 (N5235, N5209);
  nand ginst1538 (N5236, N5196, N5220);
  nand ginst1539 (N5240, N5198, N5221);
  nand ginst1540 (N5242, N5160, N5222);
  nand ginst1541 (N5243, N5163, N5225);
  nand ginst1542 (N5245, N5174, N5233);
  nand ginst1543 (N5246, N5177, N5235);
  not ginst1544 (N5250, N5240);
  not ginst1545 (N5253, N5228);
  nand ginst1546 (N5254, N5223, N5242);
  nand ginst1547 (N5257, N5224, N5243);
  nand ginst1548 (N5258, N5232, N5245);
  nand ginst1549 (N5261, N5234, N5246);
  not ginst1550 (N5266, N5257);
  buf ginst1551 (N5269, N5236);
  and ginst1552 (N5277, N2307, N5236, N5254);
  and ginst1553 (N5278, N2310, N5250, N5254);
  not ginst1554 (N5279, N5261);
  not ginst1555 (N5283, N5269);
  nand ginst1556 (N5284, N5253, N5269);
  and ginst1557 (N5285, N2310, N5236, N5266);
  and ginst1558 (N5286, N2307, N5250, N5266);
  buf ginst1559 (N5289, N5258);
  buf ginst1560 (N5292, N5258);
  nand ginst1561 (N5295, N5228, N5283);
  or ginst1562 (N5298, N5277, N5278, N5285, N5286);
  buf ginst1563 (N5303, N5279);
  buf ginst1564 (N5306, N5279);
  nand ginst1565 (N5309, N5284, N5295);
  not ginst1566 (N5312, N5292);
  not ginst1567 (N5313, N5289);
  not ginst1568 (N5322, N5306);
  not ginst1569 (N5323, N5303);
  buf ginst1570 (N5324, N5298);
  buf ginst1571 (N5327, N5298);
  buf ginst1572 (N5332, N5309);
  buf ginst1573 (N5335, N5309);
  nand ginst1574 (N5340, N5323, N5324);
  nand ginst1575 (N5341, N5322, N5327);
  not ginst1576 (N5344, N5327);
  not ginst1577 (N5345, N5324);
  nand ginst1578 (N5348, N5313, N5332);
  nand ginst1579 (N5349, N5312, N5335);
  nand ginst1580 (N5350, N5303, N5345);
  nand ginst1581 (N5351, N5306, N5344);
  not ginst1582 (N5352, N5335);
  not ginst1583 (N5353, N5332);
  nand ginst1584 (N5354, N5289, N5353);
  nand ginst1585 (N5355, N5292, N5352);
  nand ginst1586 (N5356, N5340, N5350);
  nand ginst1587 (N5357, N5341, N5351);
  nand ginst1588 (N5358, N5348, N5354);
  nand ginst1589 (N5359, N5349, N5355);
  and ginst1590 (N5360, N5356, N5357);
  nand ginst1591 (N5361, N5358, N5359);
  buf ginst1592 (N655, N50);
  not ginst1593 (N665, N50);
  buf ginst1594 (N670, N58);
  not ginst1595 (N679, N58);
  buf ginst1596 (N683, N68);
  not ginst1597 (N686, N68);
  buf ginst1598 (N690, N68);
  buf ginst1599 (N699, N77);
  not ginst1600 (N702, N77);
  buf ginst1601 (N706, N77);
  buf ginst1602 (N715, N87);
  not ginst1603 (N724, N87);
  buf ginst1604 (N727, N97);
  not ginst1605 (N736, N97);
  buf ginst1606 (N740, N107);
  not ginst1607 (N749, N107);
  buf ginst1608 (N753, N116);
  not ginst1609 (N763, N116);
  or ginst1610 (N768, N257, N264);
  not ginst1611 (N769, N1);
  buf ginst1612 (N772, N1);
  not ginst1613 (N779, N1);
  buf ginst1614 (N782, N13);
  not ginst1615 (N786, N13);
  and ginst1616 (N793, N13, N20);
  not ginst1617 (N794, N20);
  buf ginst1618 (N798, N20);
  not ginst1619 (N803, N20);
  not ginst1620 (N820, N33);
  buf ginst1621 (N821, N33);
  not ginst1622 (N825, N33);
  and ginst1623 (N829, N33, N41);
  not ginst1624 (N832, N41);
  or ginst1625 (N835, N41, N45);
  buf ginst1626 (N836, N45);
  not ginst1627 (N839, N45);
  not ginst1628 (N842, N50);
  buf ginst1629 (N845, N58);
  not ginst1630 (N848, N58);
  buf ginst1631 (N851, N68);
  not ginst1632 (N854, N68);
  buf ginst1633 (N858, N87);
  not ginst1634 (N861, N87);
  buf ginst1635 (N864, N97);
  not ginst1636 (N867, N97);
  not ginst1637 (N870, N107);
  buf ginst1638 (N874, N1);
  buf ginst1639 (N877, N68);
  buf ginst1640 (N880, N107);
  not ginst1641 (N883, N20);
  buf ginst1642 (N886, N190);
  not ginst1643 (N889, N200);
  and ginst1644 (N890, N20, N200);
  nand ginst1645 (N891, N20, N200);
  and ginst1646 (N892, N20, N179);
  not ginst1647 (N895, N20);
  or ginst1648 (N896, N33, N349);
  nand ginst1649 (N913, N1, N13);
  nand ginst1650 (N914, N1, N20, N33);
  not ginst1651 (N915, N20);
  not ginst1652 (N916, N33);
  buf ginst1653 (N917, N179);
  not ginst1654 (N920, N213);
  buf ginst1655 (N923, N343);
  buf ginst1656 (N926, N226);
  buf ginst1657 (N929, N232);
  buf ginst1658 (N932, N238);
  buf ginst1659 (N935, N244);
  buf ginst1660 (N938, N250);
  buf ginst1661 (N941, N257);
  buf ginst1662 (N944, N264);
  buf ginst1663 (N947, N270);
  buf ginst1664 (N950, N50);
  buf ginst1665 (N953, N58);
  buf ginst1666 (N956, N58);
  buf ginst1667 (N959, N97);
  buf ginst1668 (N962, N97);
  buf ginst1669 (N965, N330);

endmodule
