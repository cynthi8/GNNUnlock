//key=0010100010100000110110101110100100110001101011001100011000111001
// Main module
module b17_C_SFLL-HD(2)_64_2(P1_MEMORYFETCH_REG_SCAN_IN, DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, DATAI_27_, DATAI_26_, DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, DATAI_21_, DATAI_20_, DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, DATAI_15_, DATAI_14_, DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, DATAI_9_, DATAI_8_, DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, DATAI_2_, DATAI_1_, DATAI_0_, HOLD, NA, BS16, READY1, READY2, P1_READREQUEST_REG_SCAN_IN, P1_ADS_N_REG_SCAN_IN, P1_CODEFETCH_REG_SCAN_IN, P1_M_IO_N_REG_SCAN_IN, P1_D_C_N_REG_SCAN_IN, P1_REQUESTPENDING_REG_SCAN_IN, P1_STATEBS16_REG_SCAN_IN, P1_MORE_REG_SCAN_IN, P1_FLUSH_REG_SCAN_IN, P1_W_R_N_REG_SCAN_IN, P1_BYTEENABLE_REG_0__SCAN_IN, P1_BYTEENABLE_REG_1__SCAN_IN, P1_BYTEENABLE_REG_2__SCAN_IN, P1_BYTEENABLE_REG_3__SCAN_IN, P1_REIP_REG_31__SCAN_IN, P1_REIP_REG_30__SCAN_IN, P1_REIP_REG_29__SCAN_IN, P1_REIP_REG_28__SCAN_IN, P1_REIP_REG_27__SCAN_IN, P1_REIP_REG_26__SCAN_IN, P1_REIP_REG_25__SCAN_IN, P1_REIP_REG_24__SCAN_IN, P1_REIP_REG_23__SCAN_IN, P1_REIP_REG_22__SCAN_IN, P1_REIP_REG_21__SCAN_IN, P1_REIP_REG_20__SCAN_IN, P1_REIP_REG_19__SCAN_IN, P1_REIP_REG_18__SCAN_IN, P1_REIP_REG_17__SCAN_IN, P1_REIP_REG_16__SCAN_IN, P1_REIP_REG_15__SCAN_IN, P1_REIP_REG_14__SCAN_IN, P1_REIP_REG_13__SCAN_IN, P1_REIP_REG_12__SCAN_IN, P1_REIP_REG_11__SCAN_IN, P1_REIP_REG_10__SCAN_IN, P1_REIP_REG_9__SCAN_IN, P1_REIP_REG_8__SCAN_IN, P1_REIP_REG_7__SCAN_IN, P1_REIP_REG_6__SCAN_IN, P1_REIP_REG_5__SCAN_IN, P1_REIP_REG_4__SCAN_IN, P1_REIP_REG_3__SCAN_IN, P1_REIP_REG_2__SCAN_IN, P1_REIP_REG_1__SCAN_IN, P1_REIP_REG_0__SCAN_IN, P1_EBX_REG_31__SCAN_IN, P1_EBX_REG_30__SCAN_IN, P1_EBX_REG_29__SCAN_IN, P1_EBX_REG_28__SCAN_IN, P1_EBX_REG_27__SCAN_IN, P1_EBX_REG_26__SCAN_IN, P1_EBX_REG_25__SCAN_IN, P1_EBX_REG_24__SCAN_IN, P1_EBX_REG_23__SCAN_IN, P1_EBX_REG_22__SCAN_IN, P1_EBX_REG_21__SCAN_IN, P1_EBX_REG_20__SCAN_IN, P1_EBX_REG_19__SCAN_IN, P1_EBX_REG_18__SCAN_IN, P1_EBX_REG_17__SCAN_IN, P1_EBX_REG_16__SCAN_IN, P1_EBX_REG_15__SCAN_IN, P1_EBX_REG_14__SCAN_IN, P1_EBX_REG_13__SCAN_IN, P1_EBX_REG_12__SCAN_IN, P1_EBX_REG_11__SCAN_IN, P1_EBX_REG_10__SCAN_IN, P1_EBX_REG_9__SCAN_IN, P1_EBX_REG_8__SCAN_IN, P1_EBX_REG_7__SCAN_IN, P1_EBX_REG_6__SCAN_IN, P1_EBX_REG_5__SCAN_IN, P1_EBX_REG_4__SCAN_IN, P1_EBX_REG_3__SCAN_IN, P1_EBX_REG_2__SCAN_IN, P1_EBX_REG_1__SCAN_IN, P1_EBX_REG_0__SCAN_IN, P1_EAX_REG_31__SCAN_IN, P1_EAX_REG_30__SCAN_IN, P1_EAX_REG_29__SCAN_IN, P1_EAX_REG_28__SCAN_IN, P1_EAX_REG_27__SCAN_IN, P1_EAX_REG_26__SCAN_IN, P1_EAX_REG_25__SCAN_IN, P1_EAX_REG_24__SCAN_IN, P1_EAX_REG_23__SCAN_IN, P1_EAX_REG_22__SCAN_IN, P1_EAX_REG_21__SCAN_IN, P1_EAX_REG_20__SCAN_IN, P1_EAX_REG_19__SCAN_IN, P1_EAX_REG_18__SCAN_IN, P1_EAX_REG_17__SCAN_IN, P1_EAX_REG_16__SCAN_IN, P1_EAX_REG_15__SCAN_IN, P1_EAX_REG_14__SCAN_IN, P1_EAX_REG_13__SCAN_IN, P1_EAX_REG_12__SCAN_IN, P1_EAX_REG_11__SCAN_IN, P1_EAX_REG_10__SCAN_IN, P1_EAX_REG_9__SCAN_IN, P1_EAX_REG_8__SCAN_IN, P1_EAX_REG_7__SCAN_IN, P1_EAX_REG_6__SCAN_IN, P1_EAX_REG_5__SCAN_IN, P1_EAX_REG_4__SCAN_IN, P1_EAX_REG_3__SCAN_IN, P1_EAX_REG_2__SCAN_IN, P1_EAX_REG_1__SCAN_IN, P1_EAX_REG_0__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_0__SCAN_IN, P1_UWORD_REG_0__SCAN_IN, P1_UWORD_REG_1__SCAN_IN, P1_UWORD_REG_2__SCAN_IN, P1_UWORD_REG_3__SCAN_IN, P1_UWORD_REG_4__SCAN_IN, P1_UWORD_REG_5__SCAN_IN, P1_UWORD_REG_6__SCAN_IN, P1_UWORD_REG_7__SCAN_IN, P1_UWORD_REG_8__SCAN_IN, P1_UWORD_REG_9__SCAN_IN, P1_UWORD_REG_10__SCAN_IN, P1_UWORD_REG_11__SCAN_IN, P1_UWORD_REG_12__SCAN_IN, P1_UWORD_REG_13__SCAN_IN, P1_UWORD_REG_14__SCAN_IN, P1_LWORD_REG_0__SCAN_IN, P1_LWORD_REG_1__SCAN_IN, P1_LWORD_REG_2__SCAN_IN, P1_LWORD_REG_3__SCAN_IN, P1_LWORD_REG_4__SCAN_IN, P1_LWORD_REG_5__SCAN_IN, P1_LWORD_REG_6__SCAN_IN, P1_LWORD_REG_7__SCAN_IN, P1_LWORD_REG_8__SCAN_IN, P1_LWORD_REG_9__SCAN_IN, P1_LWORD_REG_10__SCAN_IN, P1_LWORD_REG_11__SCAN_IN, P1_LWORD_REG_12__SCAN_IN, P1_LWORD_REG_13__SCAN_IN, P1_LWORD_REG_14__SCAN_IN, P1_LWORD_REG_15__SCAN_IN, P1_PHYADDRPOINTER_REG_31__SCAN_IN, P1_PHYADDRPOINTER_REG_30__SCAN_IN, P1_PHYADDRPOINTER_REG_29__SCAN_IN, P1_PHYADDRPOINTER_REG_28__SCAN_IN, P1_PHYADDRPOINTER_REG_27__SCAN_IN, P1_PHYADDRPOINTER_REG_26__SCAN_IN, P1_PHYADDRPOINTER_REG_25__SCAN_IN, P1_PHYADDRPOINTER_REG_24__SCAN_IN, P1_PHYADDRPOINTER_REG_23__SCAN_IN, P1_PHYADDRPOINTER_REG_22__SCAN_IN, P1_PHYADDRPOINTER_REG_21__SCAN_IN, P1_PHYADDRPOINTER_REG_20__SCAN_IN, P1_PHYADDRPOINTER_REG_19__SCAN_IN, P1_PHYADDRPOINTER_REG_18__SCAN_IN, P1_PHYADDRPOINTER_REG_17__SCAN_IN, P1_PHYADDRPOINTER_REG_16__SCAN_IN, P1_PHYADDRPOINTER_REG_15__SCAN_IN, P1_PHYADDRPOINTER_REG_14__SCAN_IN, P1_PHYADDRPOINTER_REG_13__SCAN_IN, P1_PHYADDRPOINTER_REG_12__SCAN_IN, P1_PHYADDRPOINTER_REG_11__SCAN_IN, P1_PHYADDRPOINTER_REG_10__SCAN_IN, P1_PHYADDRPOINTER_REG_9__SCAN_IN, P1_PHYADDRPOINTER_REG_8__SCAN_IN, P1_PHYADDRPOINTER_REG_7__SCAN_IN, P1_PHYADDRPOINTER_REG_6__SCAN_IN, P1_PHYADDRPOINTER_REG_5__SCAN_IN, P1_PHYADDRPOINTER_REG_4__SCAN_IN, P1_PHYADDRPOINTER_REG_3__SCAN_IN, P1_PHYADDRPOINTER_REG_2__SCAN_IN, P1_PHYADDRPOINTER_REG_1__SCAN_IN, P1_PHYADDRPOINTER_REG_0__SCAN_IN, P1_INSTADDRPOINTER_REG_31__SCAN_IN, P1_INSTADDRPOINTER_REG_30__SCAN_IN, P1_INSTADDRPOINTER_REG_29__SCAN_IN, P1_INSTADDRPOINTER_REG_28__SCAN_IN, P1_INSTADDRPOINTER_REG_27__SCAN_IN, P1_INSTADDRPOINTER_REG_26__SCAN_IN, P1_INSTADDRPOINTER_REG_25__SCAN_IN, P1_INSTADDRPOINTER_REG_24__SCAN_IN, P1_INSTADDRPOINTER_REG_23__SCAN_IN, P1_INSTADDRPOINTER_REG_22__SCAN_IN, P1_INSTADDRPOINTER_REG_21__SCAN_IN, P1_INSTADDRPOINTER_REG_20__SCAN_IN, P1_INSTADDRPOINTER_REG_19__SCAN_IN, P1_INSTADDRPOINTER_REG_18__SCAN_IN, P1_INSTADDRPOINTER_REG_17__SCAN_IN, P1_INSTADDRPOINTER_REG_16__SCAN_IN, P1_INSTADDRPOINTER_REG_15__SCAN_IN, P1_INSTADDRPOINTER_REG_14__SCAN_IN, P1_INSTADDRPOINTER_REG_13__SCAN_IN, P1_INSTADDRPOINTER_REG_12__SCAN_IN, P1_INSTADDRPOINTER_REG_11__SCAN_IN, P1_INSTADDRPOINTER_REG_10__SCAN_IN, P1_INSTADDRPOINTER_REG_9__SCAN_IN, P1_INSTADDRPOINTER_REG_8__SCAN_IN, P1_INSTADDRPOINTER_REG_7__SCAN_IN, P1_INSTADDRPOINTER_REG_6__SCAN_IN, P1_INSTADDRPOINTER_REG_5__SCAN_IN, P1_INSTADDRPOINTER_REG_4__SCAN_IN, P1_INSTADDRPOINTER_REG_3__SCAN_IN, P1_INSTADDRPOINTER_REG_2__SCAN_IN, P1_INSTADDRPOINTER_REG_1__SCAN_IN, P1_INSTADDRPOINTER_REG_0__SCAN_IN, P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN, P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN, P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN, P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN, P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN, P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN, P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN, P1_INSTQUEUE_REG_0__0__SCAN_IN, P1_INSTQUEUE_REG_0__1__SCAN_IN, P1_INSTQUEUE_REG_0__2__SCAN_IN, P1_INSTQUEUE_REG_0__3__SCAN_IN, P1_INSTQUEUE_REG_0__4__SCAN_IN, P1_INSTQUEUE_REG_0__5__SCAN_IN, P1_INSTQUEUE_REG_0__6__SCAN_IN, P1_INSTQUEUE_REG_0__7__SCAN_IN, P1_INSTQUEUE_REG_1__0__SCAN_IN, P1_INSTQUEUE_REG_1__1__SCAN_IN, P1_INSTQUEUE_REG_1__2__SCAN_IN, P1_INSTQUEUE_REG_1__3__SCAN_IN, P1_INSTQUEUE_REG_1__4__SCAN_IN, P1_INSTQUEUE_REG_1__5__SCAN_IN, P1_INSTQUEUE_REG_1__6__SCAN_IN, P1_INSTQUEUE_REG_1__7__SCAN_IN, P1_INSTQUEUE_REG_2__0__SCAN_IN, P1_INSTQUEUE_REG_2__1__SCAN_IN, P1_INSTQUEUE_REG_2__2__SCAN_IN, P1_INSTQUEUE_REG_2__3__SCAN_IN, P1_INSTQUEUE_REG_2__4__SCAN_IN, P1_INSTQUEUE_REG_2__5__SCAN_IN, P1_INSTQUEUE_REG_2__6__SCAN_IN, P1_INSTQUEUE_REG_2__7__SCAN_IN, P1_INSTQUEUE_REG_3__0__SCAN_IN, P1_INSTQUEUE_REG_3__1__SCAN_IN, P1_INSTQUEUE_REG_3__2__SCAN_IN, P1_INSTQUEUE_REG_3__3__SCAN_IN, P1_INSTQUEUE_REG_3__4__SCAN_IN, P1_INSTQUEUE_REG_3__5__SCAN_IN, P1_INSTQUEUE_REG_3__6__SCAN_IN, P1_INSTQUEUE_REG_3__7__SCAN_IN, P1_INSTQUEUE_REG_4__0__SCAN_IN, BUF1_REG_0__SCAN_IN, BUF1_REG_1__SCAN_IN, BUF1_REG_2__SCAN_IN, BUF1_REG_3__SCAN_IN, BUF1_REG_4__SCAN_IN, BUF1_REG_5__SCAN_IN, BUF1_REG_6__SCAN_IN, BUF1_REG_7__SCAN_IN, BUF1_REG_8__SCAN_IN, BUF1_REG_9__SCAN_IN, BUF1_REG_10__SCAN_IN, BUF1_REG_11__SCAN_IN, BUF1_REG_12__SCAN_IN, BUF1_REG_13__SCAN_IN, BUF1_REG_14__SCAN_IN, BUF1_REG_15__SCAN_IN, BUF1_REG_16__SCAN_IN, BUF1_REG_17__SCAN_IN, BUF1_REG_18__SCAN_IN, BUF1_REG_19__SCAN_IN, BUF1_REG_20__SCAN_IN, BUF1_REG_21__SCAN_IN, BUF1_REG_22__SCAN_IN, BUF1_REG_23__SCAN_IN, BUF1_REG_24__SCAN_IN, BUF1_REG_25__SCAN_IN, BUF1_REG_26__SCAN_IN, BUF1_REG_27__SCAN_IN, BUF1_REG_28__SCAN_IN, BUF1_REG_29__SCAN_IN, BUF1_REG_30__SCAN_IN, BUF1_REG_31__SCAN_IN, BUF2_REG_0__SCAN_IN, BUF2_REG_1__SCAN_IN, BUF2_REG_2__SCAN_IN, BUF2_REG_3__SCAN_IN, BUF2_REG_4__SCAN_IN, BUF2_REG_5__SCAN_IN, BUF2_REG_6__SCAN_IN, BUF2_REG_7__SCAN_IN, BUF2_REG_8__SCAN_IN, BUF2_REG_9__SCAN_IN, BUF2_REG_10__SCAN_IN, BUF2_REG_11__SCAN_IN, BUF2_REG_12__SCAN_IN, BUF2_REG_13__SCAN_IN, BUF2_REG_14__SCAN_IN, BUF2_REG_15__SCAN_IN, BUF2_REG_16__SCAN_IN, BUF2_REG_17__SCAN_IN, BUF2_REG_18__SCAN_IN, BUF2_REG_19__SCAN_IN, BUF2_REG_20__SCAN_IN, BUF2_REG_21__SCAN_IN, BUF2_REG_22__SCAN_IN, BUF2_REG_23__SCAN_IN, BUF2_REG_24__SCAN_IN, BUF2_REG_25__SCAN_IN, BUF2_REG_26__SCAN_IN, BUF2_REG_27__SCAN_IN, BUF2_REG_28__SCAN_IN, BUF2_REG_29__SCAN_IN, BUF2_REG_30__SCAN_IN, BUF2_REG_31__SCAN_IN, READY12_REG_SCAN_IN, READY21_REG_SCAN_IN, READY22_REG_SCAN_IN, READY11_REG_SCAN_IN, P3_BE_N_REG_3__SCAN_IN, P3_BE_N_REG_2__SCAN_IN, P3_BE_N_REG_1__SCAN_IN, P3_BE_N_REG_0__SCAN_IN, P3_ADDRESS_REG_29__SCAN_IN, P3_ADDRESS_REG_28__SCAN_IN, P3_ADDRESS_REG_27__SCAN_IN, P3_ADDRESS_REG_26__SCAN_IN, P3_ADDRESS_REG_25__SCAN_IN, P3_ADDRESS_REG_24__SCAN_IN, P3_ADDRESS_REG_23__SCAN_IN, P3_ADDRESS_REG_22__SCAN_IN, P3_ADDRESS_REG_21__SCAN_IN, P3_ADDRESS_REG_20__SCAN_IN, P3_ADDRESS_REG_19__SCAN_IN, P3_ADDRESS_REG_18__SCAN_IN, P3_ADDRESS_REG_17__SCAN_IN, P3_ADDRESS_REG_16__SCAN_IN, P3_ADDRESS_REG_15__SCAN_IN, P3_ADDRESS_REG_14__SCAN_IN, P3_ADDRESS_REG_13__SCAN_IN, P3_ADDRESS_REG_12__SCAN_IN, P3_ADDRESS_REG_11__SCAN_IN, P3_ADDRESS_REG_10__SCAN_IN, P3_ADDRESS_REG_9__SCAN_IN, P3_ADDRESS_REG_8__SCAN_IN, P3_ADDRESS_REG_7__SCAN_IN, P3_ADDRESS_REG_6__SCAN_IN, P3_ADDRESS_REG_5__SCAN_IN, P3_ADDRESS_REG_4__SCAN_IN, P3_ADDRESS_REG_3__SCAN_IN, P3_ADDRESS_REG_2__SCAN_IN, P3_ADDRESS_REG_1__SCAN_IN, P3_ADDRESS_REG_0__SCAN_IN, P3_STATE_REG_2__SCAN_IN, P3_STATE_REG_1__SCAN_IN, P3_STATE_REG_0__SCAN_IN, P3_DATAWIDTH_REG_0__SCAN_IN, P3_DATAWIDTH_REG_1__SCAN_IN, P3_DATAWIDTH_REG_2__SCAN_IN, P3_DATAWIDTH_REG_3__SCAN_IN, P3_DATAWIDTH_REG_4__SCAN_IN, P3_DATAWIDTH_REG_5__SCAN_IN, P3_DATAWIDTH_REG_6__SCAN_IN, P3_DATAWIDTH_REG_7__SCAN_IN, P3_DATAWIDTH_REG_8__SCAN_IN, P3_DATAWIDTH_REG_9__SCAN_IN, P3_DATAWIDTH_REG_10__SCAN_IN, P3_DATAWIDTH_REG_11__SCAN_IN, P3_DATAWIDTH_REG_12__SCAN_IN, P3_DATAWIDTH_REG_13__SCAN_IN, P3_DATAWIDTH_REG_14__SCAN_IN, P3_DATAWIDTH_REG_15__SCAN_IN, P3_DATAWIDTH_REG_16__SCAN_IN, P3_DATAWIDTH_REG_17__SCAN_IN, P3_DATAWIDTH_REG_18__SCAN_IN, P3_DATAWIDTH_REG_19__SCAN_IN, P3_DATAWIDTH_REG_20__SCAN_IN, P3_DATAWIDTH_REG_21__SCAN_IN, P3_DATAWIDTH_REG_22__SCAN_IN, P3_DATAWIDTH_REG_23__SCAN_IN, P3_DATAWIDTH_REG_24__SCAN_IN, P3_DATAWIDTH_REG_25__SCAN_IN, P3_DATAWIDTH_REG_26__SCAN_IN, P3_DATAWIDTH_REG_27__SCAN_IN, P3_DATAWIDTH_REG_28__SCAN_IN, P3_DATAWIDTH_REG_29__SCAN_IN, P3_DATAWIDTH_REG_30__SCAN_IN, P3_DATAWIDTH_REG_31__SCAN_IN, P3_STATE2_REG_3__SCAN_IN, P3_STATE2_REG_2__SCAN_IN, P3_STATE2_REG_1__SCAN_IN, P3_STATE2_REG_0__SCAN_IN, P3_INSTQUEUE_REG_15__7__SCAN_IN, P3_INSTQUEUE_REG_15__6__SCAN_IN, P3_INSTQUEUE_REG_15__5__SCAN_IN, P3_INSTQUEUE_REG_15__4__SCAN_IN, P3_INSTQUEUE_REG_15__3__SCAN_IN, P3_INSTQUEUE_REG_15__2__SCAN_IN, P3_INSTQUEUE_REG_15__1__SCAN_IN, P3_INSTQUEUE_REG_15__0__SCAN_IN, P3_INSTQUEUE_REG_14__7__SCAN_IN, P3_INSTQUEUE_REG_14__6__SCAN_IN, P3_INSTQUEUE_REG_14__5__SCAN_IN, P3_INSTQUEUE_REG_14__4__SCAN_IN, P3_INSTQUEUE_REG_14__3__SCAN_IN, P3_INSTQUEUE_REG_14__2__SCAN_IN, P3_INSTQUEUE_REG_14__1__SCAN_IN, P3_INSTQUEUE_REG_14__0__SCAN_IN, P3_INSTQUEUE_REG_13__7__SCAN_IN, P3_INSTQUEUE_REG_13__6__SCAN_IN, P3_INSTQUEUE_REG_13__5__SCAN_IN, P3_INSTQUEUE_REG_13__4__SCAN_IN, P3_INSTQUEUE_REG_13__3__SCAN_IN, P3_INSTQUEUE_REG_13__2__SCAN_IN, P3_INSTQUEUE_REG_13__1__SCAN_IN, P3_INSTQUEUE_REG_13__0__SCAN_IN, P3_INSTQUEUE_REG_12__7__SCAN_IN, P3_INSTQUEUE_REG_12__6__SCAN_IN, P3_INSTQUEUE_REG_12__5__SCAN_IN, P3_INSTQUEUE_REG_12__4__SCAN_IN, P3_INSTQUEUE_REG_12__3__SCAN_IN, P3_INSTQUEUE_REG_12__2__SCAN_IN, P3_INSTQUEUE_REG_12__1__SCAN_IN, P3_INSTQUEUE_REG_12__0__SCAN_IN, P3_INSTQUEUE_REG_11__7__SCAN_IN, P3_INSTQUEUE_REG_11__6__SCAN_IN, P3_INSTQUEUE_REG_11__5__SCAN_IN, P3_INSTQUEUE_REG_11__4__SCAN_IN, P3_INSTQUEUE_REG_11__3__SCAN_IN, P3_INSTQUEUE_REG_11__2__SCAN_IN, P3_INSTQUEUE_REG_11__1__SCAN_IN, P3_INSTQUEUE_REG_11__0__SCAN_IN, P3_INSTQUEUE_REG_10__7__SCAN_IN, P3_INSTQUEUE_REG_10__6__SCAN_IN, P3_INSTQUEUE_REG_10__5__SCAN_IN, P3_INSTQUEUE_REG_10__4__SCAN_IN, P3_INSTQUEUE_REG_10__3__SCAN_IN, P3_INSTQUEUE_REG_10__2__SCAN_IN, P3_INSTQUEUE_REG_10__1__SCAN_IN, P3_INSTQUEUE_REG_10__0__SCAN_IN, P3_INSTQUEUE_REG_9__7__SCAN_IN, P3_INSTQUEUE_REG_9__6__SCAN_IN, P3_INSTQUEUE_REG_9__5__SCAN_IN, P3_INSTQUEUE_REG_9__4__SCAN_IN, P3_INSTQUEUE_REG_9__3__SCAN_IN, P3_INSTQUEUE_REG_9__2__SCAN_IN, P3_INSTQUEUE_REG_9__1__SCAN_IN, P3_INSTQUEUE_REG_9__0__SCAN_IN, P3_INSTQUEUE_REG_8__7__SCAN_IN, P3_INSTQUEUE_REG_8__6__SCAN_IN, P3_INSTQUEUE_REG_8__5__SCAN_IN, P3_INSTQUEUE_REG_8__4__SCAN_IN, P3_INSTQUEUE_REG_8__3__SCAN_IN, P3_INSTQUEUE_REG_8__2__SCAN_IN, P3_INSTQUEUE_REG_8__1__SCAN_IN, P3_INSTQUEUE_REG_8__0__SCAN_IN, P3_INSTQUEUE_REG_7__7__SCAN_IN, P3_INSTQUEUE_REG_7__6__SCAN_IN, P3_INSTQUEUE_REG_7__5__SCAN_IN, P3_INSTQUEUE_REG_7__4__SCAN_IN, P3_INSTQUEUE_REG_7__3__SCAN_IN, P3_INSTQUEUE_REG_7__2__SCAN_IN, P3_INSTQUEUE_REG_7__1__SCAN_IN, P3_INSTQUEUE_REG_7__0__SCAN_IN, P3_INSTQUEUE_REG_6__7__SCAN_IN, P3_INSTQUEUE_REG_6__6__SCAN_IN, P3_INSTQUEUE_REG_6__5__SCAN_IN, P3_INSTQUEUE_REG_6__4__SCAN_IN, P3_INSTQUEUE_REG_6__3__SCAN_IN, P3_INSTQUEUE_REG_6__2__SCAN_IN, P3_INSTQUEUE_REG_6__1__SCAN_IN, P3_INSTQUEUE_REG_6__0__SCAN_IN, P3_INSTQUEUE_REG_5__7__SCAN_IN, P3_INSTQUEUE_REG_5__6__SCAN_IN, P3_INSTQUEUE_REG_5__5__SCAN_IN, P3_INSTQUEUE_REG_5__4__SCAN_IN, P3_INSTQUEUE_REG_5__3__SCAN_IN, P3_INSTQUEUE_REG_5__2__SCAN_IN, P3_INSTQUEUE_REG_5__1__SCAN_IN, P3_INSTQUEUE_REG_5__0__SCAN_IN, P3_INSTQUEUE_REG_4__7__SCAN_IN, P3_INSTQUEUE_REG_4__6__SCAN_IN, P3_INSTQUEUE_REG_4__5__SCAN_IN, P3_INSTQUEUE_REG_4__4__SCAN_IN, P3_INSTQUEUE_REG_4__3__SCAN_IN, P3_INSTQUEUE_REG_4__2__SCAN_IN, P3_INSTQUEUE_REG_4__1__SCAN_IN, P3_INSTQUEUE_REG_4__0__SCAN_IN, P3_INSTQUEUE_REG_3__7__SCAN_IN, P3_INSTQUEUE_REG_3__6__SCAN_IN, P3_INSTQUEUE_REG_3__5__SCAN_IN, P3_INSTQUEUE_REG_3__4__SCAN_IN, P3_INSTQUEUE_REG_3__3__SCAN_IN, P3_INSTQUEUE_REG_3__2__SCAN_IN, P3_INSTQUEUE_REG_3__1__SCAN_IN, P3_INSTQUEUE_REG_3__0__SCAN_IN, P3_INSTQUEUE_REG_2__7__SCAN_IN, P3_INSTQUEUE_REG_2__6__SCAN_IN, P3_INSTQUEUE_REG_2__5__SCAN_IN, P3_INSTQUEUE_REG_2__4__SCAN_IN, P3_INSTQUEUE_REG_2__3__SCAN_IN, P3_INSTQUEUE_REG_2__2__SCAN_IN, P3_INSTQUEUE_REG_2__1__SCAN_IN, P3_INSTQUEUE_REG_2__0__SCAN_IN, P3_INSTQUEUE_REG_1__7__SCAN_IN, P3_INSTQUEUE_REG_1__6__SCAN_IN, P3_INSTQUEUE_REG_1__5__SCAN_IN, P3_INSTQUEUE_REG_1__4__SCAN_IN, P3_INSTQUEUE_REG_1__3__SCAN_IN, P3_INSTQUEUE_REG_1__2__SCAN_IN, P3_INSTQUEUE_REG_1__1__SCAN_IN, P3_INSTQUEUE_REG_1__0__SCAN_IN, P3_INSTQUEUE_REG_0__7__SCAN_IN, P3_INSTQUEUE_REG_0__6__SCAN_IN, P3_INSTQUEUE_REG_0__5__SCAN_IN, P3_INSTQUEUE_REG_0__4__SCAN_IN, P3_INSTQUEUE_REG_0__3__SCAN_IN, P3_INSTQUEUE_REG_0__2__SCAN_IN, P3_INSTQUEUE_REG_0__1__SCAN_IN, P3_INSTQUEUE_REG_0__0__SCAN_IN, P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN, P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN, P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN, P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN, P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN, P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN, P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN, P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P3_INSTADDRPOINTER_REG_0__SCAN_IN, P3_INSTADDRPOINTER_REG_1__SCAN_IN, P3_INSTADDRPOINTER_REG_2__SCAN_IN, P3_INSTADDRPOINTER_REG_3__SCAN_IN, P3_INSTADDRPOINTER_REG_4__SCAN_IN, P3_INSTADDRPOINTER_REG_5__SCAN_IN, P3_INSTADDRPOINTER_REG_6__SCAN_IN, P3_INSTADDRPOINTER_REG_7__SCAN_IN, P3_INSTADDRPOINTER_REG_8__SCAN_IN, P3_INSTADDRPOINTER_REG_9__SCAN_IN, P3_INSTADDRPOINTER_REG_10__SCAN_IN, P3_INSTADDRPOINTER_REG_11__SCAN_IN, P3_INSTADDRPOINTER_REG_12__SCAN_IN, P3_INSTADDRPOINTER_REG_13__SCAN_IN, P3_INSTADDRPOINTER_REG_14__SCAN_IN, P3_INSTADDRPOINTER_REG_15__SCAN_IN, P3_INSTADDRPOINTER_REG_16__SCAN_IN, P3_INSTADDRPOINTER_REG_17__SCAN_IN, P3_INSTADDRPOINTER_REG_18__SCAN_IN, P3_INSTADDRPOINTER_REG_19__SCAN_IN, P3_INSTADDRPOINTER_REG_20__SCAN_IN, P3_INSTADDRPOINTER_REG_21__SCAN_IN, P3_INSTADDRPOINTER_REG_22__SCAN_IN, P3_INSTADDRPOINTER_REG_23__SCAN_IN, P3_INSTADDRPOINTER_REG_24__SCAN_IN, P3_INSTADDRPOINTER_REG_25__SCAN_IN, P3_INSTADDRPOINTER_REG_26__SCAN_IN, P3_INSTADDRPOINTER_REG_27__SCAN_IN, P3_INSTADDRPOINTER_REG_28__SCAN_IN, P3_INSTADDRPOINTER_REG_29__SCAN_IN, P3_INSTADDRPOINTER_REG_30__SCAN_IN, P3_INSTADDRPOINTER_REG_31__SCAN_IN, P3_PHYADDRPOINTER_REG_0__SCAN_IN, P3_PHYADDRPOINTER_REG_1__SCAN_IN, P3_PHYADDRPOINTER_REG_2__SCAN_IN, P3_PHYADDRPOINTER_REG_3__SCAN_IN, P3_PHYADDRPOINTER_REG_4__SCAN_IN, P3_PHYADDRPOINTER_REG_5__SCAN_IN, P3_PHYADDRPOINTER_REG_6__SCAN_IN, P3_PHYADDRPOINTER_REG_7__SCAN_IN, P3_PHYADDRPOINTER_REG_8__SCAN_IN, P3_PHYADDRPOINTER_REG_9__SCAN_IN, P3_PHYADDRPOINTER_REG_10__SCAN_IN, P3_PHYADDRPOINTER_REG_11__SCAN_IN, P3_PHYADDRPOINTER_REG_12__SCAN_IN, P3_PHYADDRPOINTER_REG_13__SCAN_IN, P3_PHYADDRPOINTER_REG_14__SCAN_IN, P3_PHYADDRPOINTER_REG_15__SCAN_IN, P3_PHYADDRPOINTER_REG_16__SCAN_IN, P3_PHYADDRPOINTER_REG_17__SCAN_IN, P3_PHYADDRPOINTER_REG_18__SCAN_IN, P3_PHYADDRPOINTER_REG_19__SCAN_IN, P3_PHYADDRPOINTER_REG_20__SCAN_IN, P3_PHYADDRPOINTER_REG_21__SCAN_IN, P3_PHYADDRPOINTER_REG_22__SCAN_IN, P3_PHYADDRPOINTER_REG_23__SCAN_IN, P3_PHYADDRPOINTER_REG_24__SCAN_IN, P3_PHYADDRPOINTER_REG_25__SCAN_IN, P3_PHYADDRPOINTER_REG_26__SCAN_IN, P3_PHYADDRPOINTER_REG_27__SCAN_IN, P3_PHYADDRPOINTER_REG_28__SCAN_IN, P3_PHYADDRPOINTER_REG_29__SCAN_IN, P3_PHYADDRPOINTER_REG_30__SCAN_IN, P3_PHYADDRPOINTER_REG_31__SCAN_IN, P3_LWORD_REG_15__SCAN_IN, P3_LWORD_REG_14__SCAN_IN, P3_LWORD_REG_13__SCAN_IN, P3_LWORD_REG_12__SCAN_IN, P3_LWORD_REG_11__SCAN_IN, P3_LWORD_REG_10__SCAN_IN, P3_LWORD_REG_9__SCAN_IN, P3_LWORD_REG_8__SCAN_IN, P3_LWORD_REG_7__SCAN_IN, P3_LWORD_REG_6__SCAN_IN, P3_LWORD_REG_5__SCAN_IN, P3_LWORD_REG_4__SCAN_IN, P3_LWORD_REG_3__SCAN_IN, P3_LWORD_REG_2__SCAN_IN, P3_LWORD_REG_1__SCAN_IN, P3_LWORD_REG_0__SCAN_IN, P3_UWORD_REG_14__SCAN_IN, P3_UWORD_REG_13__SCAN_IN, P3_UWORD_REG_12__SCAN_IN, P3_UWORD_REG_11__SCAN_IN, P3_UWORD_REG_10__SCAN_IN, P3_UWORD_REG_9__SCAN_IN, P3_UWORD_REG_8__SCAN_IN, P3_UWORD_REG_7__SCAN_IN, P3_UWORD_REG_6__SCAN_IN, P3_UWORD_REG_5__SCAN_IN, P3_UWORD_REG_4__SCAN_IN, P3_UWORD_REG_3__SCAN_IN, P3_UWORD_REG_2__SCAN_IN, P3_UWORD_REG_1__SCAN_IN, P3_UWORD_REG_0__SCAN_IN, P3_DATAO_REG_0__SCAN_IN, P3_DATAO_REG_1__SCAN_IN, P3_DATAO_REG_2__SCAN_IN, P3_DATAO_REG_3__SCAN_IN, P3_DATAO_REG_4__SCAN_IN, P3_DATAO_REG_5__SCAN_IN, P3_DATAO_REG_6__SCAN_IN, P3_DATAO_REG_7__SCAN_IN, P3_DATAO_REG_8__SCAN_IN, P3_DATAO_REG_9__SCAN_IN, P3_DATAO_REG_10__SCAN_IN, P3_DATAO_REG_11__SCAN_IN, P3_DATAO_REG_12__SCAN_IN, P3_DATAO_REG_13__SCAN_IN, P3_DATAO_REG_14__SCAN_IN, P3_DATAO_REG_15__SCAN_IN, P3_DATAO_REG_16__SCAN_IN, P3_DATAO_REG_17__SCAN_IN, P3_DATAO_REG_18__SCAN_IN, P3_DATAO_REG_19__SCAN_IN, P3_DATAO_REG_20__SCAN_IN, P3_DATAO_REG_21__SCAN_IN, P3_DATAO_REG_22__SCAN_IN, P3_DATAO_REG_23__SCAN_IN, P3_DATAO_REG_24__SCAN_IN, P3_DATAO_REG_25__SCAN_IN, P3_DATAO_REG_26__SCAN_IN, P3_DATAO_REG_27__SCAN_IN, P3_DATAO_REG_28__SCAN_IN, P3_DATAO_REG_29__SCAN_IN, P3_DATAO_REG_30__SCAN_IN, P3_DATAO_REG_31__SCAN_IN, P3_EAX_REG_0__SCAN_IN, P3_EAX_REG_1__SCAN_IN, P3_EAX_REG_2__SCAN_IN, P3_EAX_REG_3__SCAN_IN, P3_EAX_REG_4__SCAN_IN, P3_EAX_REG_5__SCAN_IN, P3_EAX_REG_6__SCAN_IN, P3_EAX_REG_7__SCAN_IN, P3_EAX_REG_8__SCAN_IN, P3_EAX_REG_9__SCAN_IN, P3_EAX_REG_10__SCAN_IN, P3_EAX_REG_11__SCAN_IN, P3_EAX_REG_12__SCAN_IN, P3_EAX_REG_13__SCAN_IN, P3_EAX_REG_14__SCAN_IN, P3_EAX_REG_15__SCAN_IN, P3_EAX_REG_16__SCAN_IN, P3_EAX_REG_17__SCAN_IN, P3_EAX_REG_18__SCAN_IN, P3_EAX_REG_19__SCAN_IN, P3_EAX_REG_20__SCAN_IN, P3_EAX_REG_21__SCAN_IN, P3_EAX_REG_22__SCAN_IN, P3_EAX_REG_23__SCAN_IN, P3_EAX_REG_24__SCAN_IN, P3_EAX_REG_25__SCAN_IN, P3_EAX_REG_26__SCAN_IN, P3_EAX_REG_27__SCAN_IN, P3_EAX_REG_28__SCAN_IN, P3_EAX_REG_29__SCAN_IN, P3_EAX_REG_30__SCAN_IN, P3_EAX_REG_31__SCAN_IN, P3_EBX_REG_0__SCAN_IN, P3_EBX_REG_1__SCAN_IN, P3_EBX_REG_2__SCAN_IN, P3_EBX_REG_3__SCAN_IN, P3_EBX_REG_4__SCAN_IN, P3_EBX_REG_5__SCAN_IN, P3_EBX_REG_6__SCAN_IN, P3_EBX_REG_7__SCAN_IN, P3_EBX_REG_8__SCAN_IN, P3_EBX_REG_9__SCAN_IN, P3_EBX_REG_10__SCAN_IN, P3_EBX_REG_11__SCAN_IN, P3_EBX_REG_12__SCAN_IN, P3_EBX_REG_13__SCAN_IN, P3_EBX_REG_14__SCAN_IN, P3_EBX_REG_15__SCAN_IN, P3_EBX_REG_16__SCAN_IN, P3_EBX_REG_17__SCAN_IN, P3_EBX_REG_18__SCAN_IN, P3_EBX_REG_19__SCAN_IN, P3_EBX_REG_20__SCAN_IN, P3_EBX_REG_21__SCAN_IN, P3_EBX_REG_22__SCAN_IN, P3_EBX_REG_23__SCAN_IN, P3_EBX_REG_24__SCAN_IN, P3_EBX_REG_25__SCAN_IN, P3_EBX_REG_26__SCAN_IN, P3_EBX_REG_27__SCAN_IN, P3_EBX_REG_28__SCAN_IN, P3_EBX_REG_29__SCAN_IN, P3_EBX_REG_30__SCAN_IN, P3_EBX_REG_31__SCAN_IN, P3_REIP_REG_0__SCAN_IN, P3_REIP_REG_1__SCAN_IN, P3_REIP_REG_2__SCAN_IN, P3_REIP_REG_3__SCAN_IN, P3_REIP_REG_4__SCAN_IN, P3_REIP_REG_5__SCAN_IN, P3_REIP_REG_6__SCAN_IN, P3_REIP_REG_7__SCAN_IN, P3_REIP_REG_8__SCAN_IN, P3_REIP_REG_9__SCAN_IN, P3_REIP_REG_10__SCAN_IN, P3_REIP_REG_11__SCAN_IN, P3_REIP_REG_12__SCAN_IN, P3_REIP_REG_13__SCAN_IN, P3_REIP_REG_14__SCAN_IN, P3_REIP_REG_15__SCAN_IN, P3_REIP_REG_16__SCAN_IN, P3_REIP_REG_17__SCAN_IN, P3_REIP_REG_18__SCAN_IN, P3_REIP_REG_19__SCAN_IN, P3_REIP_REG_20__SCAN_IN, P3_REIP_REG_21__SCAN_IN, P3_REIP_REG_22__SCAN_IN, P3_REIP_REG_23__SCAN_IN, P3_REIP_REG_24__SCAN_IN, P3_REIP_REG_25__SCAN_IN, P3_REIP_REG_26__SCAN_IN, P3_REIP_REG_27__SCAN_IN, P3_REIP_REG_28__SCAN_IN, P3_REIP_REG_29__SCAN_IN, P3_REIP_REG_30__SCAN_IN, P3_REIP_REG_31__SCAN_IN, P3_BYTEENABLE_REG_3__SCAN_IN, P3_BYTEENABLE_REG_2__SCAN_IN, P3_BYTEENABLE_REG_1__SCAN_IN, P3_BYTEENABLE_REG_0__SCAN_IN, P3_W_R_N_REG_SCAN_IN, P3_FLUSH_REG_SCAN_IN, P3_MORE_REG_SCAN_IN, P3_STATEBS16_REG_SCAN_IN, P3_REQUESTPENDING_REG_SCAN_IN, P3_D_C_N_REG_SCAN_IN, P3_M_IO_N_REG_SCAN_IN, P3_CODEFETCH_REG_SCAN_IN, P3_ADS_N_REG_SCAN_IN, P3_READREQUEST_REG_SCAN_IN, P3_MEMORYFETCH_REG_SCAN_IN, P2_BE_N_REG_3__SCAN_IN, P2_BE_N_REG_2__SCAN_IN, P2_BE_N_REG_1__SCAN_IN, P2_BE_N_REG_0__SCAN_IN, P2_ADDRESS_REG_29__SCAN_IN, P2_ADDRESS_REG_28__SCAN_IN, P2_ADDRESS_REG_27__SCAN_IN, P2_ADDRESS_REG_26__SCAN_IN, P2_ADDRESS_REG_25__SCAN_IN, P2_ADDRESS_REG_24__SCAN_IN, P2_ADDRESS_REG_23__SCAN_IN, P2_ADDRESS_REG_22__SCAN_IN, P2_ADDRESS_REG_21__SCAN_IN, P2_ADDRESS_REG_20__SCAN_IN, P2_ADDRESS_REG_19__SCAN_IN, P2_ADDRESS_REG_18__SCAN_IN, P2_ADDRESS_REG_17__SCAN_IN, P2_ADDRESS_REG_16__SCAN_IN, P2_ADDRESS_REG_15__SCAN_IN, P2_ADDRESS_REG_14__SCAN_IN, P2_ADDRESS_REG_13__SCAN_IN, P2_ADDRESS_REG_12__SCAN_IN, P2_ADDRESS_REG_11__SCAN_IN, P2_ADDRESS_REG_10__SCAN_IN, P2_ADDRESS_REG_9__SCAN_IN, P2_ADDRESS_REG_8__SCAN_IN, P2_ADDRESS_REG_7__SCAN_IN, P2_ADDRESS_REG_6__SCAN_IN, P2_ADDRESS_REG_5__SCAN_IN, P2_ADDRESS_REG_4__SCAN_IN, P2_ADDRESS_REG_3__SCAN_IN, P2_ADDRESS_REG_2__SCAN_IN, P2_ADDRESS_REG_1__SCAN_IN, P2_ADDRESS_REG_0__SCAN_IN, P2_STATE_REG_2__SCAN_IN, P2_STATE_REG_1__SCAN_IN, P2_STATE_REG_0__SCAN_IN, P2_DATAWIDTH_REG_0__SCAN_IN, P2_DATAWIDTH_REG_1__SCAN_IN, P2_DATAWIDTH_REG_2__SCAN_IN, P2_DATAWIDTH_REG_3__SCAN_IN, P2_DATAWIDTH_REG_4__SCAN_IN, P2_DATAWIDTH_REG_5__SCAN_IN, P2_DATAWIDTH_REG_6__SCAN_IN, P2_DATAWIDTH_REG_7__SCAN_IN, P2_DATAWIDTH_REG_8__SCAN_IN, P2_DATAWIDTH_REG_9__SCAN_IN, P2_DATAWIDTH_REG_10__SCAN_IN, P2_DATAWIDTH_REG_11__SCAN_IN, P2_DATAWIDTH_REG_12__SCAN_IN, P2_DATAWIDTH_REG_13__SCAN_IN, P2_DATAWIDTH_REG_14__SCAN_IN, P2_DATAWIDTH_REG_15__SCAN_IN, P2_DATAWIDTH_REG_16__SCAN_IN, P2_DATAWIDTH_REG_17__SCAN_IN, P2_DATAWIDTH_REG_18__SCAN_IN, P2_DATAWIDTH_REG_19__SCAN_IN, P2_DATAWIDTH_REG_20__SCAN_IN, P2_DATAWIDTH_REG_21__SCAN_IN, P2_DATAWIDTH_REG_22__SCAN_IN, P2_DATAWIDTH_REG_23__SCAN_IN, P2_DATAWIDTH_REG_24__SCAN_IN, P2_DATAWIDTH_REG_25__SCAN_IN, P2_DATAWIDTH_REG_26__SCAN_IN, P2_DATAWIDTH_REG_27__SCAN_IN, P2_DATAWIDTH_REG_28__SCAN_IN, P2_DATAWIDTH_REG_29__SCAN_IN, P2_DATAWIDTH_REG_30__SCAN_IN, P2_DATAWIDTH_REG_31__SCAN_IN, P2_STATE2_REG_3__SCAN_IN, P2_STATE2_REG_2__SCAN_IN, P2_STATE2_REG_1__SCAN_IN, P2_STATE2_REG_0__SCAN_IN, P2_INSTQUEUE_REG_15__7__SCAN_IN, P2_INSTQUEUE_REG_15__6__SCAN_IN, P2_INSTQUEUE_REG_15__5__SCAN_IN, P2_INSTQUEUE_REG_15__4__SCAN_IN, P2_INSTQUEUE_REG_15__3__SCAN_IN, P2_INSTQUEUE_REG_15__2__SCAN_IN, P2_INSTQUEUE_REG_15__1__SCAN_IN, P2_INSTQUEUE_REG_15__0__SCAN_IN, P2_INSTQUEUE_REG_14__7__SCAN_IN, P2_INSTQUEUE_REG_14__6__SCAN_IN, P2_INSTQUEUE_REG_14__5__SCAN_IN, P2_INSTQUEUE_REG_14__4__SCAN_IN, P2_INSTQUEUE_REG_14__3__SCAN_IN, P2_INSTQUEUE_REG_14__2__SCAN_IN, P2_INSTQUEUE_REG_14__1__SCAN_IN, P2_INSTQUEUE_REG_14__0__SCAN_IN, P2_INSTQUEUE_REG_13__7__SCAN_IN, P2_INSTQUEUE_REG_13__6__SCAN_IN, P2_INSTQUEUE_REG_13__5__SCAN_IN, P2_INSTQUEUE_REG_13__4__SCAN_IN, P2_INSTQUEUE_REG_13__3__SCAN_IN, P2_INSTQUEUE_REG_13__2__SCAN_IN, P2_INSTQUEUE_REG_13__1__SCAN_IN, P2_INSTQUEUE_REG_13__0__SCAN_IN, P2_INSTQUEUE_REG_12__7__SCAN_IN, P2_INSTQUEUE_REG_12__6__SCAN_IN, P2_INSTQUEUE_REG_12__5__SCAN_IN, P2_INSTQUEUE_REG_12__4__SCAN_IN, P2_INSTQUEUE_REG_12__3__SCAN_IN, P2_INSTQUEUE_REG_12__2__SCAN_IN, P2_INSTQUEUE_REG_12__1__SCAN_IN, P2_INSTQUEUE_REG_12__0__SCAN_IN, P2_INSTQUEUE_REG_11__7__SCAN_IN, P2_INSTQUEUE_REG_11__6__SCAN_IN, P2_INSTQUEUE_REG_11__5__SCAN_IN, P2_INSTQUEUE_REG_11__4__SCAN_IN, P2_INSTQUEUE_REG_11__3__SCAN_IN, P2_INSTQUEUE_REG_11__2__SCAN_IN, P2_INSTQUEUE_REG_11__1__SCAN_IN, P2_INSTQUEUE_REG_11__0__SCAN_IN, P2_INSTQUEUE_REG_10__7__SCAN_IN, P2_INSTQUEUE_REG_10__6__SCAN_IN, P2_INSTQUEUE_REG_10__5__SCAN_IN, P2_INSTQUEUE_REG_10__4__SCAN_IN, P2_INSTQUEUE_REG_10__3__SCAN_IN, P2_INSTQUEUE_REG_10__2__SCAN_IN, P2_INSTQUEUE_REG_10__1__SCAN_IN, P2_INSTQUEUE_REG_10__0__SCAN_IN, P2_INSTQUEUE_REG_9__7__SCAN_IN, P2_INSTQUEUE_REG_9__6__SCAN_IN, P2_INSTQUEUE_REG_9__5__SCAN_IN, P2_INSTQUEUE_REG_9__4__SCAN_IN, P2_INSTQUEUE_REG_9__3__SCAN_IN, P2_INSTQUEUE_REG_9__2__SCAN_IN, P2_INSTQUEUE_REG_9__1__SCAN_IN, P2_INSTQUEUE_REG_9__0__SCAN_IN, P2_INSTQUEUE_REG_8__7__SCAN_IN, P2_INSTQUEUE_REG_8__6__SCAN_IN, P2_INSTQUEUE_REG_8__5__SCAN_IN, P2_INSTQUEUE_REG_8__4__SCAN_IN, P2_INSTQUEUE_REG_8__3__SCAN_IN, P2_INSTQUEUE_REG_8__2__SCAN_IN, P2_INSTQUEUE_REG_8__1__SCAN_IN, P2_INSTQUEUE_REG_8__0__SCAN_IN, P2_INSTQUEUE_REG_7__7__SCAN_IN, P2_INSTQUEUE_REG_7__6__SCAN_IN, P2_INSTQUEUE_REG_7__5__SCAN_IN, P2_INSTQUEUE_REG_7__4__SCAN_IN, P2_INSTQUEUE_REG_7__3__SCAN_IN, P2_INSTQUEUE_REG_7__2__SCAN_IN, P2_INSTQUEUE_REG_7__1__SCAN_IN, P2_INSTQUEUE_REG_7__0__SCAN_IN, P2_INSTQUEUE_REG_6__7__SCAN_IN, P2_INSTQUEUE_REG_6__6__SCAN_IN, P2_INSTQUEUE_REG_6__5__SCAN_IN, P2_INSTQUEUE_REG_6__4__SCAN_IN, P2_INSTQUEUE_REG_6__3__SCAN_IN, P2_INSTQUEUE_REG_6__2__SCAN_IN, P2_INSTQUEUE_REG_6__1__SCAN_IN, P2_INSTQUEUE_REG_6__0__SCAN_IN, P2_INSTQUEUE_REG_5__7__SCAN_IN, P2_INSTQUEUE_REG_5__6__SCAN_IN, P2_INSTQUEUE_REG_5__5__SCAN_IN, P2_INSTQUEUE_REG_5__4__SCAN_IN, P2_INSTQUEUE_REG_5__3__SCAN_IN, P2_INSTQUEUE_REG_5__2__SCAN_IN, P2_INSTQUEUE_REG_5__1__SCAN_IN, P2_INSTQUEUE_REG_5__0__SCAN_IN, P2_INSTQUEUE_REG_4__7__SCAN_IN, P2_INSTQUEUE_REG_4__6__SCAN_IN, P2_INSTQUEUE_REG_4__5__SCAN_IN, P2_INSTQUEUE_REG_4__4__SCAN_IN, P2_INSTQUEUE_REG_4__3__SCAN_IN, P2_INSTQUEUE_REG_4__2__SCAN_IN, P2_INSTQUEUE_REG_4__1__SCAN_IN, P2_INSTQUEUE_REG_4__0__SCAN_IN, P2_INSTQUEUE_REG_3__7__SCAN_IN, P2_INSTQUEUE_REG_3__6__SCAN_IN, P2_INSTQUEUE_REG_3__5__SCAN_IN, P2_INSTQUEUE_REG_3__4__SCAN_IN, P2_INSTQUEUE_REG_3__3__SCAN_IN, P2_INSTQUEUE_REG_3__2__SCAN_IN, P2_INSTQUEUE_REG_3__1__SCAN_IN, P2_INSTQUEUE_REG_3__0__SCAN_IN, P2_INSTQUEUE_REG_2__7__SCAN_IN, P2_INSTQUEUE_REG_2__6__SCAN_IN, P2_INSTQUEUE_REG_2__5__SCAN_IN, P2_INSTQUEUE_REG_2__4__SCAN_IN, P2_INSTQUEUE_REG_2__3__SCAN_IN, P2_INSTQUEUE_REG_2__2__SCAN_IN, P2_INSTQUEUE_REG_2__1__SCAN_IN, P2_INSTQUEUE_REG_2__0__SCAN_IN, P2_INSTQUEUE_REG_1__7__SCAN_IN, P2_INSTQUEUE_REG_1__6__SCAN_IN, P2_INSTQUEUE_REG_1__5__SCAN_IN, P2_INSTQUEUE_REG_1__4__SCAN_IN, P2_INSTQUEUE_REG_1__3__SCAN_IN, P2_INSTQUEUE_REG_1__2__SCAN_IN, P2_INSTQUEUE_REG_1__1__SCAN_IN, P2_INSTQUEUE_REG_1__0__SCAN_IN, P2_INSTQUEUE_REG_0__7__SCAN_IN, P2_INSTQUEUE_REG_0__6__SCAN_IN, P2_INSTQUEUE_REG_0__5__SCAN_IN, P2_INSTQUEUE_REG_0__4__SCAN_IN, P2_INSTQUEUE_REG_0__3__SCAN_IN, P2_INSTQUEUE_REG_0__2__SCAN_IN, P2_INSTQUEUE_REG_0__1__SCAN_IN, P2_INSTQUEUE_REG_0__0__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN, P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN, P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN, P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN, P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN, P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P2_INSTADDRPOINTER_REG_0__SCAN_IN, P2_INSTADDRPOINTER_REG_1__SCAN_IN, P2_INSTADDRPOINTER_REG_2__SCAN_IN, P2_INSTADDRPOINTER_REG_3__SCAN_IN, P2_INSTADDRPOINTER_REG_4__SCAN_IN, P2_INSTADDRPOINTER_REG_5__SCAN_IN, P2_INSTADDRPOINTER_REG_6__SCAN_IN, P2_INSTADDRPOINTER_REG_7__SCAN_IN, P2_INSTADDRPOINTER_REG_8__SCAN_IN, P2_INSTADDRPOINTER_REG_9__SCAN_IN, P2_INSTADDRPOINTER_REG_10__SCAN_IN, P2_INSTADDRPOINTER_REG_11__SCAN_IN, P2_INSTADDRPOINTER_REG_12__SCAN_IN, P2_INSTADDRPOINTER_REG_13__SCAN_IN, P2_INSTADDRPOINTER_REG_14__SCAN_IN, P2_INSTADDRPOINTER_REG_15__SCAN_IN, P2_INSTADDRPOINTER_REG_16__SCAN_IN, P2_INSTADDRPOINTER_REG_17__SCAN_IN, P2_INSTADDRPOINTER_REG_18__SCAN_IN, P2_INSTADDRPOINTER_REG_19__SCAN_IN, P2_INSTADDRPOINTER_REG_20__SCAN_IN, P2_INSTADDRPOINTER_REG_21__SCAN_IN, P2_INSTADDRPOINTER_REG_22__SCAN_IN, P2_INSTADDRPOINTER_REG_23__SCAN_IN, P2_INSTADDRPOINTER_REG_24__SCAN_IN, P2_INSTADDRPOINTER_REG_25__SCAN_IN, P2_INSTADDRPOINTER_REG_26__SCAN_IN, P2_INSTADDRPOINTER_REG_27__SCAN_IN, P2_INSTADDRPOINTER_REG_28__SCAN_IN, P2_INSTADDRPOINTER_REG_29__SCAN_IN, P2_INSTADDRPOINTER_REG_30__SCAN_IN, P2_INSTADDRPOINTER_REG_31__SCAN_IN, P2_PHYADDRPOINTER_REG_0__SCAN_IN, P2_PHYADDRPOINTER_REG_1__SCAN_IN, P2_PHYADDRPOINTER_REG_2__SCAN_IN, P2_PHYADDRPOINTER_REG_3__SCAN_IN, P2_PHYADDRPOINTER_REG_4__SCAN_IN, P2_PHYADDRPOINTER_REG_5__SCAN_IN, P2_PHYADDRPOINTER_REG_6__SCAN_IN, P2_PHYADDRPOINTER_REG_7__SCAN_IN, P2_PHYADDRPOINTER_REG_8__SCAN_IN, P2_PHYADDRPOINTER_REG_9__SCAN_IN, P2_PHYADDRPOINTER_REG_10__SCAN_IN, P2_PHYADDRPOINTER_REG_11__SCAN_IN, P2_PHYADDRPOINTER_REG_12__SCAN_IN, P2_PHYADDRPOINTER_REG_13__SCAN_IN, P2_PHYADDRPOINTER_REG_14__SCAN_IN, P2_PHYADDRPOINTER_REG_15__SCAN_IN, P2_PHYADDRPOINTER_REG_16__SCAN_IN, P2_PHYADDRPOINTER_REG_17__SCAN_IN, P2_PHYADDRPOINTER_REG_18__SCAN_IN, P2_PHYADDRPOINTER_REG_19__SCAN_IN, P2_PHYADDRPOINTER_REG_20__SCAN_IN, P2_PHYADDRPOINTER_REG_21__SCAN_IN, P2_PHYADDRPOINTER_REG_22__SCAN_IN, P2_PHYADDRPOINTER_REG_23__SCAN_IN, P2_PHYADDRPOINTER_REG_24__SCAN_IN, P2_PHYADDRPOINTER_REG_25__SCAN_IN, P2_PHYADDRPOINTER_REG_26__SCAN_IN, P2_PHYADDRPOINTER_REG_27__SCAN_IN, P2_PHYADDRPOINTER_REG_28__SCAN_IN, P2_PHYADDRPOINTER_REG_29__SCAN_IN, P2_PHYADDRPOINTER_REG_30__SCAN_IN, P2_PHYADDRPOINTER_REG_31__SCAN_IN, P2_LWORD_REG_15__SCAN_IN, P2_LWORD_REG_14__SCAN_IN, P2_LWORD_REG_13__SCAN_IN, P2_LWORD_REG_12__SCAN_IN, P2_LWORD_REG_11__SCAN_IN, P2_LWORD_REG_10__SCAN_IN, P2_LWORD_REG_9__SCAN_IN, P2_LWORD_REG_8__SCAN_IN, P2_LWORD_REG_7__SCAN_IN, P2_LWORD_REG_6__SCAN_IN, P2_LWORD_REG_5__SCAN_IN, P2_LWORD_REG_4__SCAN_IN, P2_LWORD_REG_3__SCAN_IN, P2_LWORD_REG_2__SCAN_IN, P2_LWORD_REG_1__SCAN_IN, P2_LWORD_REG_0__SCAN_IN, P2_UWORD_REG_14__SCAN_IN, P2_UWORD_REG_13__SCAN_IN, P2_UWORD_REG_12__SCAN_IN, P2_UWORD_REG_11__SCAN_IN, P2_UWORD_REG_10__SCAN_IN, P2_UWORD_REG_9__SCAN_IN, P2_UWORD_REG_8__SCAN_IN, P2_UWORD_REG_7__SCAN_IN, P2_UWORD_REG_6__SCAN_IN, P2_UWORD_REG_5__SCAN_IN, P2_UWORD_REG_4__SCAN_IN, P2_UWORD_REG_3__SCAN_IN, P2_UWORD_REG_2__SCAN_IN, P2_UWORD_REG_1__SCAN_IN, P2_UWORD_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN, P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN, P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN, P2_DATAO_REG_5__SCAN_IN, P2_DATAO_REG_6__SCAN_IN, P2_DATAO_REG_7__SCAN_IN, P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_9__SCAN_IN, P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_11__SCAN_IN, P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_13__SCAN_IN, P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_15__SCAN_IN, P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_17__SCAN_IN, P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_19__SCAN_IN, P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_21__SCAN_IN, P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_23__SCAN_IN, P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_25__SCAN_IN, P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_27__SCAN_IN, P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_29__SCAN_IN, P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_31__SCAN_IN, P2_EAX_REG_0__SCAN_IN, P2_EAX_REG_1__SCAN_IN, P2_EAX_REG_2__SCAN_IN, P2_EAX_REG_3__SCAN_IN, P2_EAX_REG_4__SCAN_IN, P2_EAX_REG_5__SCAN_IN, P2_EAX_REG_6__SCAN_IN, P2_EAX_REG_7__SCAN_IN, P2_EAX_REG_8__SCAN_IN, P2_EAX_REG_9__SCAN_IN, P2_EAX_REG_10__SCAN_IN, P2_EAX_REG_11__SCAN_IN, P2_EAX_REG_12__SCAN_IN, P2_EAX_REG_13__SCAN_IN, P2_EAX_REG_14__SCAN_IN, P2_EAX_REG_15__SCAN_IN, P2_EAX_REG_16__SCAN_IN, P2_EAX_REG_17__SCAN_IN, P2_EAX_REG_18__SCAN_IN, P2_EAX_REG_19__SCAN_IN, P2_EAX_REG_20__SCAN_IN, P2_EAX_REG_21__SCAN_IN, P2_EAX_REG_22__SCAN_IN, P2_EAX_REG_23__SCAN_IN, P2_EAX_REG_24__SCAN_IN, P2_EAX_REG_25__SCAN_IN, P2_EAX_REG_26__SCAN_IN, P2_EAX_REG_27__SCAN_IN, P2_EAX_REG_28__SCAN_IN, P2_EAX_REG_29__SCAN_IN, P2_EAX_REG_30__SCAN_IN, P2_EAX_REG_31__SCAN_IN, P2_EBX_REG_0__SCAN_IN, P2_EBX_REG_1__SCAN_IN, P2_EBX_REG_2__SCAN_IN, P2_EBX_REG_3__SCAN_IN, P2_EBX_REG_4__SCAN_IN, P2_EBX_REG_5__SCAN_IN, P2_EBX_REG_6__SCAN_IN, P2_EBX_REG_7__SCAN_IN, P2_EBX_REG_8__SCAN_IN, P2_EBX_REG_9__SCAN_IN, P2_EBX_REG_10__SCAN_IN, P2_EBX_REG_11__SCAN_IN, P2_EBX_REG_12__SCAN_IN, P2_EBX_REG_13__SCAN_IN, P2_EBX_REG_14__SCAN_IN, P2_EBX_REG_15__SCAN_IN, P2_EBX_REG_16__SCAN_IN, P2_EBX_REG_17__SCAN_IN, P2_EBX_REG_18__SCAN_IN, P2_EBX_REG_19__SCAN_IN, P2_EBX_REG_20__SCAN_IN, P2_EBX_REG_21__SCAN_IN, P2_EBX_REG_22__SCAN_IN, P2_EBX_REG_23__SCAN_IN, P2_EBX_REG_24__SCAN_IN, P2_EBX_REG_25__SCAN_IN, P2_EBX_REG_26__SCAN_IN, P2_EBX_REG_27__SCAN_IN, P2_EBX_REG_28__SCAN_IN, P2_EBX_REG_29__SCAN_IN, P2_EBX_REG_30__SCAN_IN, P2_EBX_REG_31__SCAN_IN, P2_REIP_REG_0__SCAN_IN, P2_REIP_REG_1__SCAN_IN, P2_REIP_REG_2__SCAN_IN, P2_REIP_REG_3__SCAN_IN, P2_REIP_REG_4__SCAN_IN, P2_REIP_REG_5__SCAN_IN, P2_REIP_REG_6__SCAN_IN, P2_REIP_REG_7__SCAN_IN, P2_REIP_REG_8__SCAN_IN, P2_REIP_REG_9__SCAN_IN, P2_REIP_REG_10__SCAN_IN, P2_REIP_REG_11__SCAN_IN, P2_REIP_REG_12__SCAN_IN, P2_REIP_REG_13__SCAN_IN, P2_REIP_REG_14__SCAN_IN, P2_REIP_REG_15__SCAN_IN, P2_REIP_REG_16__SCAN_IN, P2_REIP_REG_17__SCAN_IN, P2_REIP_REG_18__SCAN_IN, P2_REIP_REG_19__SCAN_IN, P2_REIP_REG_20__SCAN_IN, P2_REIP_REG_21__SCAN_IN, P2_REIP_REG_22__SCAN_IN, P2_REIP_REG_23__SCAN_IN, P2_REIP_REG_24__SCAN_IN, P2_REIP_REG_25__SCAN_IN, P2_REIP_REG_26__SCAN_IN, P2_REIP_REG_27__SCAN_IN, P2_REIP_REG_28__SCAN_IN, P2_REIP_REG_29__SCAN_IN, P2_REIP_REG_30__SCAN_IN, P2_REIP_REG_31__SCAN_IN, P2_BYTEENABLE_REG_3__SCAN_IN, P2_BYTEENABLE_REG_2__SCAN_IN, P2_BYTEENABLE_REG_1__SCAN_IN, P2_BYTEENABLE_REG_0__SCAN_IN, P2_W_R_N_REG_SCAN_IN, P2_FLUSH_REG_SCAN_IN, P2_MORE_REG_SCAN_IN, P2_STATEBS16_REG_SCAN_IN, P2_REQUESTPENDING_REG_SCAN_IN, P2_D_C_N_REG_SCAN_IN, P2_M_IO_N_REG_SCAN_IN, P2_CODEFETCH_REG_SCAN_IN, P2_ADS_N_REG_SCAN_IN, P2_READREQUEST_REG_SCAN_IN, P2_MEMORYFETCH_REG_SCAN_IN, P1_BE_N_REG_3__SCAN_IN, P1_BE_N_REG_2__SCAN_IN, P1_BE_N_REG_1__SCAN_IN, P1_BE_N_REG_0__SCAN_IN, P1_ADDRESS_REG_29__SCAN_IN, P1_ADDRESS_REG_28__SCAN_IN, P1_ADDRESS_REG_27__SCAN_IN, P1_ADDRESS_REG_26__SCAN_IN, P1_ADDRESS_REG_25__SCAN_IN, P1_ADDRESS_REG_24__SCAN_IN, P1_ADDRESS_REG_23__SCAN_IN, P1_ADDRESS_REG_22__SCAN_IN, P1_ADDRESS_REG_21__SCAN_IN, P1_ADDRESS_REG_20__SCAN_IN, P1_ADDRESS_REG_19__SCAN_IN, P1_ADDRESS_REG_18__SCAN_IN, P1_ADDRESS_REG_17__SCAN_IN, P1_ADDRESS_REG_16__SCAN_IN, P1_ADDRESS_REG_15__SCAN_IN, P1_ADDRESS_REG_14__SCAN_IN, P1_ADDRESS_REG_13__SCAN_IN, P1_ADDRESS_REG_12__SCAN_IN, P1_ADDRESS_REG_11__SCAN_IN, P1_ADDRESS_REG_10__SCAN_IN, P1_ADDRESS_REG_9__SCAN_IN, P1_ADDRESS_REG_8__SCAN_IN, P1_ADDRESS_REG_7__SCAN_IN, P1_ADDRESS_REG_6__SCAN_IN, P1_ADDRESS_REG_5__SCAN_IN, P1_ADDRESS_REG_4__SCAN_IN, P1_ADDRESS_REG_3__SCAN_IN, P1_ADDRESS_REG_2__SCAN_IN, P1_ADDRESS_REG_1__SCAN_IN, P1_ADDRESS_REG_0__SCAN_IN, P1_STATE_REG_2__SCAN_IN, P1_STATE_REG_1__SCAN_IN, P1_STATE_REG_0__SCAN_IN, P1_DATAWIDTH_REG_0__SCAN_IN, P1_DATAWIDTH_REG_1__SCAN_IN, P1_DATAWIDTH_REG_2__SCAN_IN, P1_DATAWIDTH_REG_3__SCAN_IN, P1_DATAWIDTH_REG_4__SCAN_IN, P1_DATAWIDTH_REG_5__SCAN_IN, P1_DATAWIDTH_REG_6__SCAN_IN, P1_DATAWIDTH_REG_7__SCAN_IN, P1_DATAWIDTH_REG_8__SCAN_IN, P1_DATAWIDTH_REG_9__SCAN_IN, P1_DATAWIDTH_REG_10__SCAN_IN, P1_DATAWIDTH_REG_11__SCAN_IN, P1_DATAWIDTH_REG_12__SCAN_IN, P1_DATAWIDTH_REG_13__SCAN_IN, P1_DATAWIDTH_REG_14__SCAN_IN, P1_DATAWIDTH_REG_15__SCAN_IN, P1_DATAWIDTH_REG_16__SCAN_IN, P1_DATAWIDTH_REG_17__SCAN_IN, P1_DATAWIDTH_REG_18__SCAN_IN, P1_DATAWIDTH_REG_19__SCAN_IN, P1_DATAWIDTH_REG_20__SCAN_IN, P1_DATAWIDTH_REG_21__SCAN_IN, P1_DATAWIDTH_REG_22__SCAN_IN, P1_DATAWIDTH_REG_23__SCAN_IN, P1_DATAWIDTH_REG_24__SCAN_IN, P1_DATAWIDTH_REG_25__SCAN_IN, P1_DATAWIDTH_REG_26__SCAN_IN, P1_DATAWIDTH_REG_27__SCAN_IN, P1_DATAWIDTH_REG_28__SCAN_IN, P1_DATAWIDTH_REG_29__SCAN_IN, P1_DATAWIDTH_REG_30__SCAN_IN, P1_DATAWIDTH_REG_31__SCAN_IN, P1_STATE2_REG_3__SCAN_IN, P1_STATE2_REG_2__SCAN_IN, P1_STATE2_REG_1__SCAN_IN, P1_STATE2_REG_0__SCAN_IN, P1_INSTQUEUE_REG_15__7__SCAN_IN, P1_INSTQUEUE_REG_15__6__SCAN_IN, P1_INSTQUEUE_REG_15__5__SCAN_IN, P1_INSTQUEUE_REG_15__4__SCAN_IN, P1_INSTQUEUE_REG_15__3__SCAN_IN, P1_INSTQUEUE_REG_15__2__SCAN_IN, P1_INSTQUEUE_REG_15__1__SCAN_IN, P1_INSTQUEUE_REG_15__0__SCAN_IN, P1_INSTQUEUE_REG_14__7__SCAN_IN, P1_INSTQUEUE_REG_14__6__SCAN_IN, P1_INSTQUEUE_REG_14__5__SCAN_IN, P1_INSTQUEUE_REG_14__4__SCAN_IN, P1_INSTQUEUE_REG_14__3__SCAN_IN, P1_INSTQUEUE_REG_14__2__SCAN_IN, P1_INSTQUEUE_REG_14__1__SCAN_IN, P1_INSTQUEUE_REG_14__0__SCAN_IN, P1_INSTQUEUE_REG_13__7__SCAN_IN, P1_INSTQUEUE_REG_13__6__SCAN_IN, P1_INSTQUEUE_REG_13__5__SCAN_IN, P1_INSTQUEUE_REG_13__4__SCAN_IN, P1_INSTQUEUE_REG_13__3__SCAN_IN, P1_INSTQUEUE_REG_13__2__SCAN_IN, P1_INSTQUEUE_REG_13__1__SCAN_IN, P1_INSTQUEUE_REG_13__0__SCAN_IN, P1_INSTQUEUE_REG_12__7__SCAN_IN, P1_INSTQUEUE_REG_12__6__SCAN_IN, P1_INSTQUEUE_REG_12__5__SCAN_IN, P1_INSTQUEUE_REG_12__4__SCAN_IN, P1_INSTQUEUE_REG_12__3__SCAN_IN, P1_INSTQUEUE_REG_12__2__SCAN_IN, P1_INSTQUEUE_REG_12__1__SCAN_IN, P1_INSTQUEUE_REG_12__0__SCAN_IN, P1_INSTQUEUE_REG_11__7__SCAN_IN, P1_INSTQUEUE_REG_11__6__SCAN_IN, P1_INSTQUEUE_REG_11__5__SCAN_IN, P1_INSTQUEUE_REG_11__4__SCAN_IN, P1_INSTQUEUE_REG_11__3__SCAN_IN, P1_INSTQUEUE_REG_11__2__SCAN_IN, P1_INSTQUEUE_REG_11__1__SCAN_IN, P1_INSTQUEUE_REG_11__0__SCAN_IN, P1_INSTQUEUE_REG_10__7__SCAN_IN, P1_INSTQUEUE_REG_10__6__SCAN_IN, P1_INSTQUEUE_REG_10__5__SCAN_IN, P1_INSTQUEUE_REG_10__4__SCAN_IN, P1_INSTQUEUE_REG_10__3__SCAN_IN, P1_INSTQUEUE_REG_10__2__SCAN_IN, P1_INSTQUEUE_REG_10__1__SCAN_IN, P1_INSTQUEUE_REG_10__0__SCAN_IN, P1_INSTQUEUE_REG_9__7__SCAN_IN, P1_INSTQUEUE_REG_9__6__SCAN_IN, P1_INSTQUEUE_REG_9__5__SCAN_IN, P1_INSTQUEUE_REG_9__4__SCAN_IN, P1_INSTQUEUE_REG_9__3__SCAN_IN, P1_INSTQUEUE_REG_9__2__SCAN_IN, P1_INSTQUEUE_REG_9__1__SCAN_IN, P1_INSTQUEUE_REG_9__0__SCAN_IN, P1_INSTQUEUE_REG_8__7__SCAN_IN, P1_INSTQUEUE_REG_8__6__SCAN_IN, P1_INSTQUEUE_REG_8__5__SCAN_IN, P1_INSTQUEUE_REG_8__4__SCAN_IN, P1_INSTQUEUE_REG_8__3__SCAN_IN, P1_INSTQUEUE_REG_8__2__SCAN_IN, P1_INSTQUEUE_REG_8__1__SCAN_IN, P1_INSTQUEUE_REG_8__0__SCAN_IN, P1_INSTQUEUE_REG_7__7__SCAN_IN, P1_INSTQUEUE_REG_7__6__SCAN_IN, P1_INSTQUEUE_REG_7__5__SCAN_IN, P1_INSTQUEUE_REG_7__4__SCAN_IN, P1_INSTQUEUE_REG_7__3__SCAN_IN, P1_INSTQUEUE_REG_7__2__SCAN_IN, P1_INSTQUEUE_REG_7__1__SCAN_IN, P1_INSTQUEUE_REG_7__0__SCAN_IN, P1_INSTQUEUE_REG_6__7__SCAN_IN, P1_INSTQUEUE_REG_6__6__SCAN_IN, P1_INSTQUEUE_REG_6__5__SCAN_IN, P1_INSTQUEUE_REG_6__4__SCAN_IN, P1_INSTQUEUE_REG_6__3__SCAN_IN, P1_INSTQUEUE_REG_6__2__SCAN_IN, P1_INSTQUEUE_REG_6__1__SCAN_IN, P1_INSTQUEUE_REG_6__0__SCAN_IN, P1_INSTQUEUE_REG_5__7__SCAN_IN, P1_INSTQUEUE_REG_5__6__SCAN_IN, P1_INSTQUEUE_REG_5__5__SCAN_IN, P1_INSTQUEUE_REG_5__4__SCAN_IN, P1_INSTQUEUE_REG_5__3__SCAN_IN, P1_INSTQUEUE_REG_5__2__SCAN_IN, P1_INSTQUEUE_REG_5__1__SCAN_IN, P1_INSTQUEUE_REG_5__0__SCAN_IN, P1_INSTQUEUE_REG_4__7__SCAN_IN, P1_INSTQUEUE_REG_4__6__SCAN_IN, P1_INSTQUEUE_REG_4__5__SCAN_IN, P1_INSTQUEUE_REG_4__4__SCAN_IN, P1_INSTQUEUE_REG_4__3__SCAN_IN, P1_INSTQUEUE_REG_4__2__SCAN_IN, P1_INSTQUEUE_REG_4__1__SCAN_IN, keyinput0, keyinput1, keyinput2, keyinput3, keyinput4, keyinput5, keyinput6, keyinput7, keyinput8, keyinput9, keyinput10, keyinput11, keyinput12, keyinput13, keyinput14, keyinput15, keyinput16, keyinput17, keyinput18, keyinput19, keyinput20, keyinput21, keyinput22, keyinput23, keyinput24, keyinput25, keyinput26, keyinput27, keyinput28, keyinput29, keyinput30, keyinput31, keyinput32, keyinput33, keyinput34, keyinput35, keyinput36, keyinput37, keyinput38, keyinput39, keyinput40, keyinput41, keyinput42, keyinput43, keyinput44, keyinput45, keyinput46, keyinput47, keyinput48, keyinput49, keyinput50, keyinput51, keyinput52, keyinput53, keyinput54, keyinput55, keyinput56, keyinput57, keyinput58, keyinput59, keyinput60, keyinput61, keyinput62, keyinput63, P3_DATAO_REG_31__SCAN_IN, P3_DATAO_REG_30__SCAN_IN, P3_DATAO_REG_29__SCAN_IN, P3_DATAO_REG_28__SCAN_IN, P3_DATAO_REG_27__SCAN_IN, P3_DATAO_REG_26__SCAN_IN, P3_DATAO_REG_25__SCAN_IN, P3_DATAO_REG_24__SCAN_IN, P3_DATAO_REG_23__SCAN_IN, P3_DATAO_REG_22__SCAN_IN, P3_DATAO_REG_21__SCAN_IN, P3_DATAO_REG_20__SCAN_IN, P3_DATAO_REG_19__SCAN_IN, P3_DATAO_REG_18__SCAN_IN, P3_DATAO_REG_17__SCAN_IN, P3_DATAO_REG_16__SCAN_IN, P3_DATAO_REG_15__SCAN_IN, P3_DATAO_REG_14__SCAN_IN, P3_DATAO_REG_13__SCAN_IN, P3_DATAO_REG_12__SCAN_IN, P3_DATAO_REG_11__SCAN_IN, P3_DATAO_REG_10__SCAN_IN, P3_DATAO_REG_9__SCAN_IN, P3_DATAO_REG_8__SCAN_IN, P3_DATAO_REG_7__SCAN_IN, P3_DATAO_REG_6__SCAN_IN, P3_DATAO_REG_5__SCAN_IN, P3_DATAO_REG_4__SCAN_IN, P3_DATAO_REG_3__SCAN_IN, P3_DATAO_REG_2__SCAN_IN, P3_DATAO_REG_1__SCAN_IN, P3_DATAO_REG_0__SCAN_IN, P1_ADDRESS_REG_29__SCAN_IN, P1_ADDRESS_REG_28__SCAN_IN, P1_ADDRESS_REG_27__SCAN_IN, P1_ADDRESS_REG_26__SCAN_IN, P1_ADDRESS_REG_25__SCAN_IN, P1_ADDRESS_REG_24__SCAN_IN, P1_ADDRESS_REG_23__SCAN_IN, P1_ADDRESS_REG_22__SCAN_IN, P1_ADDRESS_REG_21__SCAN_IN, P1_ADDRESS_REG_20__SCAN_IN, P1_ADDRESS_REG_19__SCAN_IN, P1_ADDRESS_REG_18__SCAN_IN, P1_ADDRESS_REG_17__SCAN_IN, P1_ADDRESS_REG_16__SCAN_IN, P1_ADDRESS_REG_15__SCAN_IN, P1_ADDRESS_REG_14__SCAN_IN, P1_ADDRESS_REG_13__SCAN_IN, P1_ADDRESS_REG_12__SCAN_IN, P1_ADDRESS_REG_11__SCAN_IN, P1_ADDRESS_REG_10__SCAN_IN, P1_ADDRESS_REG_9__SCAN_IN, P1_ADDRESS_REG_8__SCAN_IN, P1_ADDRESS_REG_7__SCAN_IN, P1_ADDRESS_REG_6__SCAN_IN, P1_ADDRESS_REG_5__SCAN_IN, P1_ADDRESS_REG_4__SCAN_IN, P1_ADDRESS_REG_3__SCAN_IN, P1_ADDRESS_REG_2__SCAN_IN, P1_ADDRESS_REG_1__SCAN_IN, P1_ADDRESS_REG_0__SCAN_IN, U355, U356, U357, U358, U359, U360, U361, U362, U363, U364, U366, U367, U368, U369, U370, U371, U372, U373, U374, U375, U347, U348, U349, U350, U351, U352, U353, U354, U365, U376, P3_W_R_N_REG_SCAN_IN, P3_D_C_N_REG_SCAN_IN, P3_M_IO_N_REG_SCAN_IN, P1_ADS_N_REG_SCAN_IN, P3_ADS_N_REG_SCAN_IN, U247, U246, U245, U244, U243, U242, U241, U240, U239, U238, U237, U236, U235, U234, U233, U232, U231, U230, U229, U228, U227, U226, U225, U224, U223, U222, U221, U220, U219, U218, U217, U216, U251, U252, U253, U254, U255, U256, U257, U258, U259, U260, U261, U262, U263, U264, U265, U266, U267, U268, U269, U270, U271, U272, U273, U274, U275, U276, U277, U278, U279, U280, U281, U282, U212, U215, U213, U214, P3_U3274, P3_U3275, P3_U3276, P3_U3277, P3_U3061, P3_U3060, P3_U3059, P3_U3058, P3_U3057, P3_U3056, P3_U3055, P3_U3054, P3_U3053, P3_U3052, P3_U3051, P3_U3050, P3_U3049, P3_U3048, P3_U3047, P3_U3046, P3_U3045, P3_U3044, P3_U3043, P3_U3042, P3_U3041, P3_U3040, P3_U3039, P3_U3038, P3_U3037, P3_U3036, P3_U3035, P3_U3034, P3_U3033, P3_U3032, P3_U3031, P3_U3030, P3_U3029, P3_U3280, P3_U3281, P3_U3028, P3_U3027, P3_U3026, P3_U3025, P3_U3024, P3_U3023, P3_U3022, P3_U3021, P3_U3020, P3_U3019, P3_U3018, P3_U3017, P3_U3016, P3_U3015, P3_U3014, P3_U3013, P3_U3012, P3_U3011, P3_U3010, P3_U3009, P3_U3008, P3_U3007, P3_U3006, P3_U3005, P3_U3004, P3_U3003, P3_U3002, P3_U3001, P3_U3000, P3_U2999, P3_U3282, P3_U2998, P3_U2997, P3_U2996, P3_U2995, P3_U2994, P3_U2993, P3_U2992, P3_U2991, P3_U2990, P3_U2989, P3_U2988, P3_U2987, P3_U2986, P3_U2985, P3_U2984, P3_U2983, P3_U2982, P3_U2981, P3_U2980, P3_U2979, P3_U2978, P3_U2977, P3_U2976, P3_U2975, P3_U2974, P3_U2973, P3_U2972, P3_U2971, P3_U2970, P3_U2969, P3_U2968, P3_U2967, P3_U2966, P3_U2965, P3_U2964, P3_U2963, P3_U2962, P3_U2961, P3_U2960, P3_U2959, P3_U2958, P3_U2957, P3_U2956, P3_U2955, P3_U2954, P3_U2953, P3_U2952, P3_U2951, P3_U2950, P3_U2949, P3_U2948, P3_U2947, P3_U2946, P3_U2945, P3_U2944, P3_U2943, P3_U2942, P3_U2941, P3_U2940, P3_U2939, P3_U2938, P3_U2937, P3_U2936, P3_U2935, P3_U2934, P3_U2933, P3_U2932, P3_U2931, P3_U2930, P3_U2929, P3_U2928, P3_U2927, P3_U2926, P3_U2925, P3_U2924, P3_U2923, P3_U2922, P3_U2921, P3_U2920, P3_U2919, P3_U2918, P3_U2917, P3_U2916, P3_U2915, P3_U2914, P3_U2913, P3_U2912, P3_U2911, P3_U2910, P3_U2909, P3_U2908, P3_U2907, P3_U2906, P3_U2905, P3_U2904, P3_U2903, P3_U2902, P3_U2901, P3_U2900, P3_U2899, P3_U2898, P3_U2897, P3_U2896, P3_U2895, P3_U2894, P3_U2893, P3_U2892, P3_U2891, P3_U2890, P3_U2889, P3_U2888, P3_U2887, P3_U2886, P3_U2885, P3_U2884, P3_U2883, P3_U2882, P3_U2881, P3_U2880, P3_U2879, P3_U2878, P3_U2877, P3_U2876, P3_U2875, P3_U2874, P3_U2873, P3_U2872, P3_U2871, P3_U2870, P3_U2869, P3_U2868, P3_U3284, P3_U3285, P3_U3288, P3_U3289, P3_U3290, P3_U2867, P3_U2866, P3_U2865, P3_U2864, P3_U2863, P3_U2862, P3_U2861, P3_U2860, P3_U2859, P3_U2858, P3_U2857, P3_U2856, P3_U2855, P3_U2854, P3_U2853, P3_U2852, P3_U2851, P3_U2850, P3_U2849, P3_U2848, P3_U2847, P3_U2846, P3_U2845, P3_U2844, P3_U2843, P3_U2842, P3_U2841, P3_U2840, P3_U2839, P3_U2838, P3_U2837, P3_U2836, P3_U2835, P3_U2834, P3_U2833, P3_U2832, P3_U2831, P3_U2830, P3_U2829, P3_U2828, P3_U2827, P3_U2826, P3_U2825, P3_U2824, P3_U2823, P3_U2822, P3_U2821, P3_U2820, P3_U2819, P3_U2818, P3_U2817, P3_U2816, P3_U2815, P3_U2814, P3_U2813, P3_U2812, P3_U2811, P3_U2810, P3_U2809, P3_U2808, P3_U2807, P3_U2806, P3_U2805, P3_U2804, P3_U2803, P3_U2802, P3_U2801, P3_U2800, P3_U2799, P3_U2798, P3_U2797, P3_U2796, P3_U2795, P3_U2794, P3_U2793, P3_U2792, P3_U2791, P3_U2790, P3_U2789, P3_U2788, P3_U2787, P3_U2786, P3_U2785, P3_U2784, P3_U2783, P3_U2782, P3_U2781, P3_U2780, P3_U2779, P3_U2778, P3_U2777, P3_U2776, P3_U2775, P3_U2774, P3_U2773, P3_U2772, P3_U2771, P3_U2770, P3_U2769, P3_U2768, P3_U2767, P3_U2766, P3_U2765, P3_U2764, P3_U2763, P3_U2762, P3_U2761, P3_U2760, P3_U2759, P3_U2758, P3_U2757, P3_U2756, P3_U2755, P3_U2754, P3_U2753, P3_U2752, P3_U2751, P3_U2750, P3_U2749, P3_U2748, P3_U2747, P3_U2746, P3_U2745, P3_U2744, P3_U2743, P3_U2742, P3_U2741, P3_U2740, P3_U2739, P3_U2738, P3_U2737, P3_U2736, P3_U2735, P3_U2734, P3_U2733, P3_U2732, P3_U2731, P3_U2730, P3_U2729, P3_U2728, P3_U2727, P3_U2726, P3_U2725, P3_U2724, P3_U2723, P3_U2722, P3_U2721, P3_U2720, P3_U2719, P3_U2718, P3_U2717, P3_U2716, P3_U2715, P3_U2714, P3_U2713, P3_U2712, P3_U2711, P3_U2710, P3_U2709, P3_U2708, P3_U2707, P3_U2706, P3_U2705, P3_U2704, P3_U2703, P3_U2702, P3_U2701, P3_U2700, P3_U2699, P3_U2698, P3_U2697, P3_U2696, P3_U2695, P3_U2694, P3_U2693, P3_U2692, P3_U2691, P3_U2690, P3_U2689, P3_U2688, P3_U2687, P3_U2686, P3_U2685, P3_U2684, P3_U2683, P3_U2682, P3_U2681, P3_U2680, P3_U2679, P3_U2678, P3_U2677, P3_U2676, P3_U2675, P3_U2674, P3_U2673, P3_U2672, P3_U2671, P3_U2670, P3_U2669, P3_U2668, P3_U2667, P3_U2666, P3_U2665, P3_U2664, P3_U2663, P3_U2662, P3_U2661, P3_U2660, P3_U2659, P3_U2658, P3_U2657, P3_U2656, P3_U2655, P3_U2654, P3_U2653, P3_U2652, P3_U2651, P3_U2650, P3_U2649, P3_U2648, P3_U2647, P3_U2646, P3_U2645, P3_U2644, P3_U2643, P3_U2642, P3_U2641, P3_U2640, P3_U2639, P3_U3292, P3_U2638, P3_U3293, P3_U3294, P3_U2637, P3_U3295, P3_U2636, P3_U3296, P3_U2635, P3_U3297, P3_U2634, P3_U2633, P3_U3298, P3_U3299, P2_U3585, P2_U3586, P2_U3587, P2_U3588, P2_U3241, P2_U3240, P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234, P2_U3233, P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227, P2_U3226, P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220, P2_U3219, P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3214, P2_U3213, P2_U3212, P2_U3211, P2_U3210, P2_U3209, P2_U3591, P2_U3592, P2_U3208, P2_U3207, P2_U3206, P2_U3205, P2_U3204, P2_U3203, P2_U3202, P2_U3201, P2_U3200, P2_U3199, P2_U3198, P2_U3197, P2_U3196, P2_U3195, P2_U3194, P2_U3193, P2_U3192, P2_U3191, P2_U3190, P2_U3189, P2_U3188, P2_U3187, P2_U3186, P2_U3185, P2_U3184, P2_U3183, P2_U3182, P2_U3181, P2_U3180, P2_U3179, P2_U3593, P2_U3178, P2_U3177, P2_U3176, P2_U3175, P2_U3174, P2_U3173, P2_U3172, P2_U3171, P2_U3170, P2_U3169, P2_U3168, P2_U3167, P2_U3166, P2_U3165, P2_U3164, P2_U3163, P2_U3162, P2_U3161, P2_U3160, P2_U3159, P2_U3158, P2_U3157, P2_U3156, P2_U3155, P2_U3154, P2_U3153, P2_U3152, P2_U3151, P2_U3150, P2_U3149, P2_U3148, P2_U3147, P2_U3146, P2_U3145, P2_U3144, P2_U3143, P2_U3142, P2_U3141, P2_U3140, P2_U3139, P2_U3138, P2_U3137, P2_U3136, P2_U3135, P2_U3134, P2_U3133, P2_U3132, P2_U3131, P2_U3130, P2_U3129, P2_U3128, P2_U3127, P2_U3126, P2_U3125, P2_U3124, P2_U3123, P2_U3122, P2_U3121, P2_U3120, P2_U3119, P2_U3118, P2_U3117, P2_U3116, P2_U3115, P2_U3114, P2_U3113, P2_U3112, P2_U3111, P2_U3110, P2_U3109, P2_U3108, P2_U3107, P2_U3106, P2_U3105, P2_U3104, P2_U3103, P2_U3102, P2_U3101, P2_U3100, P2_U3099, P2_U3098, P2_U3097, P2_U3096, P2_U3095, P2_U3094, P2_U3093, P2_U3092, P2_U3091, P2_U3090, P2_U3089, P2_U3088, P2_U3087, P2_U3086, P2_U3085, P2_U3084, P2_U3083, P2_U3082, P2_U3081, P2_U3080, P2_U3079, P2_U3078, P2_U3077, P2_U3076, P2_U3075, P2_U3074, P2_U3073, P2_U3072, P2_U3071, P2_U3070, P2_U3069, P2_U3068, P2_U3067, P2_U3066, P2_U3065, P2_U3064, P2_U3063, P2_U3062, P2_U3061, P2_U3060, P2_U3059, P2_U3058, P2_U3057, P2_U3056, P2_U3055, P2_U3054, P2_U3053, P2_U3052, P2_U3051, P2_U3050, P2_U3049, P2_U3048, P2_U3595, P2_U3596, P2_U3599, P2_U3600, P2_U3601, P2_U3047, P2_U3602, P2_U3603, P2_U3604, P2_U3605, P2_U3046, P2_U3045, P2_U3044, P2_U3043, P2_U3042, P2_U3041, P2_U3040, P2_U3039, P2_U3038, P2_U3037, P2_U3036, P2_U3035, P2_U3034, P2_U3033, P2_U3032, P2_U3031, P2_U3030, P2_U3029, P2_U3028, P2_U3027, P2_U3026, P2_U3025, P2_U3024, P2_U3023, P2_U3022, P2_U3021, P2_U3020, P2_U3019, P2_U3018, P2_U3017, P2_U3016, P2_U3015, P2_U3014, P2_U3013, P2_U3012, P2_U3011, P2_U3010, P2_U3009, P2_U3008, P2_U3007, P2_U3006, P2_U3005, P2_U3004, P2_U3003, P2_U3002, P2_U3001, P2_U3000, P2_U2999, P2_U2998, P2_U2997, P2_U2996, P2_U2995, P2_U2994, P2_U2993, P2_U2992, P2_U2991, P2_U2990, P2_U2989, P2_U2988, P2_U2987, P2_U2986, P2_U2985, P2_U2984, P2_U2983, P2_U2982, P2_U2981, P2_U2980, P2_U2979, P2_U2978, P2_U2977, P2_U2976, P2_U2975, P2_U2974, P2_U2973, P2_U2972, P2_U2971, P2_U2970, P2_U2969, P2_U2968, P2_U2967, P2_U2966, P2_U2965, P2_U2964, P2_U2963, P2_U2962, P2_U2961, P2_U2960, P2_U2959, P2_U2958, P2_U2957, P2_U2956, P2_U2955, P2_U2954, P2_U2953, P2_U2952, P2_U2951, P2_U2950, P2_U2949, P2_U2948, P2_U2947, P2_U2946, P2_U2945, P2_U2944, P2_U2943, P2_U2942, P2_U2941, P2_U2940, P2_U2939, P2_U2938, P2_U2937, P2_U2936, P2_U2935, P2_U2934, P2_U2933, P2_U2932, P2_U2931, P2_U2930, P2_U2929, P2_U2928, P2_U2927, P2_U2926, P2_U2925, P2_U2924, P2_U2923, P2_U2922, P2_U2921, P2_U2920, P2_U2919, P2_U2918, P2_U2917, P2_U2916, P2_U2915, P2_U2914, P2_U2913, P2_U2912, P2_U2911, P2_U2910, P2_U2909, P2_U2908, P2_U2907, P2_U2906, P2_U2905, P2_U2904, P2_U2903, P2_U2902, P2_U2901, P2_U2900, P2_U2899, P2_U2898, P2_U2897, P2_U2896, P2_U2895, P2_U2894, P2_U2893, P2_U2892, P2_U2891, P2_U2890, P2_U2889, P2_U2888, P2_U2887, P2_U2886, P2_U2885, P2_U2884, P2_U2883, P2_U2882, P2_U2881, P2_U2880, P2_U2879, P2_U2878, P2_U2877, P2_U2876, P2_U2875, P2_U2874, P2_U2873, P2_U2872, P2_U2871, P2_U2870, P2_U2869, P2_U2868, P2_U2867, P2_U2866, P2_U2865, P2_U2864, P2_U2863, P2_U2862, P2_U2861, P2_U2860, P2_U2859, P2_U2858, P2_U2857, P2_U2856, P2_U2855, P2_U2854, P2_U2853, P2_U2852, P2_U2851, P2_U2850, P2_U2849, P2_U2848, P2_U2847, P2_U2846, P2_U2845, P2_U2844, P2_U2843, P2_U2842, P2_U2841, P2_U2840, P2_U2839, P2_U2838, P2_U2837, P2_U2836, P2_U2835, P2_U2834, P2_U2833, P2_U2832, P2_U2831, P2_U2830, P2_U2829, P2_U2828, P2_U2827, P2_U2826, P2_U2825, P2_U2824, P2_U2823, P2_U2822, P2_U2821, P2_U2820, P2_U3608, P2_U2819, P2_U3609, P2_U2818, P2_U3610, P2_U2817, P2_U3611, P2_U2816, P2_U2815, P2_U3612, P2_U2814, P1_U3458, P1_U3459, P1_U3460, P1_U3461, P1_U3226, P1_U3225, P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218, P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3212, P1_U3211, P1_U3210, P1_U3209, P1_U3208, P1_U3207, P1_U3206, P1_U3205, P1_U3204, P1_U3203, P1_U3202, P1_U3201, P1_U3200, P1_U3199, P1_U3198, P1_U3197, P1_U3196, P1_U3195, P1_U3194, P1_U3464, P1_U3465, P1_U3193, P1_U3192, P1_U3191, P1_U3190, P1_U3189, P1_U3188, P1_U3187, P1_U3186, P1_U3185, P1_U3184, P1_U3183, P1_U3182, P1_U3181, P1_U3180, P1_U3179, P1_U3178, P1_U3177, P1_U3176, P1_U3175, P1_U3174, P1_U3173, P1_U3172, P1_U3171, P1_U3170, P1_U3169, P1_U3168, P1_U3167, P1_U3166, P1_U3165, P1_U3164, P1_U3466, P1_U3163, P1_U3162, P1_U3161, P1_U3160, P1_U3159, P1_U3158, P1_U3157, P1_U3156, P1_U3155, P1_U3154, P1_U3153, P1_U3152, P1_U3151, P1_U3150, P1_U3149, P1_U3148, P1_U3147, P1_U3146, P1_U3145, P1_U3144, P1_U3143, P1_U3142, P1_U3141, P1_U3140, P1_U3139, P1_U3138, P1_U3137, P1_U3136, P1_U3135, P1_U3134, P1_U3133, P1_U3132, P1_U3131, P1_U3130, P1_U3129, P1_U3128, P1_U3127, P1_U3126, P1_U3125, P1_U3124, P1_U3123, P1_U3122, P1_U3121, P1_U3120, P1_U3119, P1_U3118, P1_U3117, P1_U3116, P1_U3115, P1_U3114, P1_U3113, P1_U3112, P1_U3111, P1_U3110, P1_U3109, P1_U3108, P1_U3107, P1_U3106, P1_U3105, P1_U3104, P1_U3103, P1_U3102, P1_U3101, P1_U3100, P1_U3099, P1_U3098, P1_U3097, P1_U3096, P1_U3095, P1_U3094, P1_U3093, P1_U3092, P1_U3091, P1_U3090, P1_U3089, P1_U3088, P1_U3087, P1_U3086, P1_U3085, P1_U3084, P1_U3083, P1_U3082, P1_U3081, P1_U3080, P1_U3079, P1_U3078, P1_U3077, P1_U3076, P1_U3075, P1_U3074, P1_U3073, P1_U3072, P1_U3071, P1_U3070, P1_U3069, P1_U3068, P1_U3067, P1_U3066, P1_U3065, P1_U3064, P1_U3063, P1_U3062, P1_U3061, P1_U3060, P1_U3059, P1_U3058, P1_U3057, P1_U3056, P1_U3055, P1_U3054, P1_U3053, P1_U3052, P1_U3051, P1_U3050, P1_U3049, P1_U3048, P1_U3047, P1_U3046, P1_U3045, P1_U3044, P1_U3043, P1_U3042, P1_U3041, P1_U3040, P1_U3039, P1_U3038, P1_U3037, P1_U3036, P1_U3035, P1_U3034, P1_U3033, P1_U3468, P1_U3469, P1_U3472, P1_U3473, P1_U3474, P1_U3032, P1_U3475, P1_U3476, P1_U3477, P1_U3478, P1_U3031, P1_U3030, P1_U3029, P1_U3028, P1_U3027, P1_U3026, P1_U3025, P1_U3024, P1_U3023, P1_U3022, P1_U3021, P1_U3020, P1_U3019, P1_U3018, P1_U3017, P1_U3016, P1_U3015, P1_U3014, P1_U3013, P1_U3012, P1_U3011, P1_U3010, P1_U3009, P1_U3008, P1_U3007, P1_U3006, P1_U3005, P1_U3004, P1_U3003, P1_U3002, P1_U3001, P1_U3000, P1_U2999, P1_U2998, P1_U2997, P1_U2996, P1_U2995, P1_U2994, P1_U2993, P1_U2992, P1_U2991, P1_U2990, P1_U2989, P1_U2988, P1_U2987, P1_U2986, P1_U2985, P1_U2984, P1_U2983, P1_U2982, P1_U2981, P1_U2980, P1_U2979, P1_U2978, P1_U2977, P1_U2976, P1_U2975, P1_U2974, P1_U2973, P1_U2972, P1_U2971, P1_U2970, P1_U2969, P1_U2968, P1_U2967, P1_U2966, P1_U2965, P1_U2964, P1_U2963, P1_U2962, P1_U2961, P1_U2960, P1_U2959, P1_U2958, P1_U2957, P1_U2956, P1_U2955, P1_U2954, P1_U2953, P1_U2952, P1_U2951, P1_U2950, P1_U2949, P1_U2948, P1_U2947, P1_U2946, P1_U2945, P1_U2944, P1_U2943, P1_U2942, P1_U2941, P1_U2940, P1_U2939, P1_U2938, P1_U2937, P1_U2936, P1_U2935, P1_U2934, P1_U2933, P1_U2932, P1_U2931, P1_U2930, P1_U2929, P1_U2928, P1_U2927, P1_U2926, P1_U2925, P1_U2924, P1_U2923, P1_U2922, P1_U2921, P1_U2920, P1_U2919, P1_U2918, P1_U2917, P1_U2916, P1_U2915, P1_U2914, P1_U2913, P1_U2912, P1_U2911, P1_U2910, P1_U2909, P1_U2908, P1_U2907, P1_U2906, P1_U2905, P1_U2904, P1_U2903, P1_U2902, P1_U2901, P1_U2900, P1_U2899, P1_U2898, P1_U2897, P1_U2896, P1_U2895, P1_U2894, P1_U2893, P1_U2892, P1_U2891, P1_U2890, P1_U2889, P1_U2888, P1_U2887, P1_U2886, P1_U2885, P1_U2884, P1_U2883, P1_U2882, P1_U2881, P1_U2880, P1_U2879, P1_U2878, P1_U2877, P1_U2876, P1_U2875, P1_U2874, P1_U2873, P1_U2872, P1_U2871, P1_U2870, P1_U2869, P1_U2868, P1_U2867, P1_U2866, P1_U2865, P1_U2864, P1_U2863, P1_U2862, P1_U2861, P1_U2860, P1_U2859, P1_U2858, P1_U2857, P1_U2856, P1_U2855, P1_U2854, P1_U2853, P1_U2852, P1_U2851, P1_U2850, P1_U2849, P1_U2848, P1_U2847, P1_U2846, P1_U2845, P1_U2844, P1_U2843, P1_U2842, P1_U2841, P1_U2840, P1_U2839, P1_U2838, P1_U2837, P1_U2836, P1_U2835, P1_U2834, P1_U2833, P1_U2832, P1_U2831, P1_U2830, P1_U2829, P1_U2828, P1_U2827, P1_U2826, P1_U2825, P1_U2824, P1_U2823, P1_U2822, P1_U2821, P1_U2820, P1_U2819, P1_U2818, P1_U2817, P1_U2816, P1_U2815, P1_U2814, P1_U2813, P1_U2812, P1_U2811, P1_U2810, P1_U2809, P1_U2808, P1_U3481, P1_U2807, P1_U3482, P1_U3483, P1_U2806, P1_U3484, P1_U2805, P1_U3485, P1_U2804, P1_U3486, P1_U2803, P1_U2802, P1_U3487, P1_U2801);

  input P1_MEMORYFETCH_REG_SCAN_IN, DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, DATAI_27_, DATAI_26_, DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, DATAI_21_, DATAI_20_, DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, DATAI_15_, DATAI_14_, DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, DATAI_9_, DATAI_8_, DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, DATAI_2_, DATAI_1_, DATAI_0_, HOLD, NA, BS16, READY1, READY2, P1_READREQUEST_REG_SCAN_IN, P1_ADS_N_REG_SCAN_IN, P1_CODEFETCH_REG_SCAN_IN, P1_M_IO_N_REG_SCAN_IN, P1_D_C_N_REG_SCAN_IN, P1_REQUESTPENDING_REG_SCAN_IN, P1_STATEBS16_REG_SCAN_IN, P1_MORE_REG_SCAN_IN, P1_FLUSH_REG_SCAN_IN, P1_W_R_N_REG_SCAN_IN, P1_BYTEENABLE_REG_0__SCAN_IN, P1_BYTEENABLE_REG_1__SCAN_IN, P1_BYTEENABLE_REG_2__SCAN_IN, P1_BYTEENABLE_REG_3__SCAN_IN, P1_REIP_REG_31__SCAN_IN, P1_REIP_REG_30__SCAN_IN, P1_REIP_REG_29__SCAN_IN, P1_REIP_REG_28__SCAN_IN, P1_REIP_REG_27__SCAN_IN, P1_REIP_REG_26__SCAN_IN, P1_REIP_REG_25__SCAN_IN, P1_REIP_REG_24__SCAN_IN, P1_REIP_REG_23__SCAN_IN, P1_REIP_REG_22__SCAN_IN, P1_REIP_REG_21__SCAN_IN, P1_REIP_REG_20__SCAN_IN, P1_REIP_REG_19__SCAN_IN, P1_REIP_REG_18__SCAN_IN, P1_REIP_REG_17__SCAN_IN, P1_REIP_REG_16__SCAN_IN, P1_REIP_REG_15__SCAN_IN, P1_REIP_REG_14__SCAN_IN, P1_REIP_REG_13__SCAN_IN, P1_REIP_REG_12__SCAN_IN, P1_REIP_REG_11__SCAN_IN, P1_REIP_REG_10__SCAN_IN, P1_REIP_REG_9__SCAN_IN, P1_REIP_REG_8__SCAN_IN, P1_REIP_REG_7__SCAN_IN, P1_REIP_REG_6__SCAN_IN, P1_REIP_REG_5__SCAN_IN, P1_REIP_REG_4__SCAN_IN, P1_REIP_REG_3__SCAN_IN, P1_REIP_REG_2__SCAN_IN, P1_REIP_REG_1__SCAN_IN, P1_REIP_REG_0__SCAN_IN, P1_EBX_REG_31__SCAN_IN, P1_EBX_REG_30__SCAN_IN, P1_EBX_REG_29__SCAN_IN, P1_EBX_REG_28__SCAN_IN, P1_EBX_REG_27__SCAN_IN, P1_EBX_REG_26__SCAN_IN, P1_EBX_REG_25__SCAN_IN, P1_EBX_REG_24__SCAN_IN, P1_EBX_REG_23__SCAN_IN, P1_EBX_REG_22__SCAN_IN, P1_EBX_REG_21__SCAN_IN, P1_EBX_REG_20__SCAN_IN, P1_EBX_REG_19__SCAN_IN, P1_EBX_REG_18__SCAN_IN, P1_EBX_REG_17__SCAN_IN, P1_EBX_REG_16__SCAN_IN, P1_EBX_REG_15__SCAN_IN, P1_EBX_REG_14__SCAN_IN, P1_EBX_REG_13__SCAN_IN, P1_EBX_REG_12__SCAN_IN, P1_EBX_REG_11__SCAN_IN, P1_EBX_REG_10__SCAN_IN, P1_EBX_REG_9__SCAN_IN, P1_EBX_REG_8__SCAN_IN, P1_EBX_REG_7__SCAN_IN, P1_EBX_REG_6__SCAN_IN, P1_EBX_REG_5__SCAN_IN, P1_EBX_REG_4__SCAN_IN, P1_EBX_REG_3__SCAN_IN, P1_EBX_REG_2__SCAN_IN, P1_EBX_REG_1__SCAN_IN, P1_EBX_REG_0__SCAN_IN, P1_EAX_REG_31__SCAN_IN, P1_EAX_REG_30__SCAN_IN, P1_EAX_REG_29__SCAN_IN, P1_EAX_REG_28__SCAN_IN, P1_EAX_REG_27__SCAN_IN, P1_EAX_REG_26__SCAN_IN, P1_EAX_REG_25__SCAN_IN, P1_EAX_REG_24__SCAN_IN, P1_EAX_REG_23__SCAN_IN, P1_EAX_REG_22__SCAN_IN, P1_EAX_REG_21__SCAN_IN, P1_EAX_REG_20__SCAN_IN, P1_EAX_REG_19__SCAN_IN, P1_EAX_REG_18__SCAN_IN, P1_EAX_REG_17__SCAN_IN, P1_EAX_REG_16__SCAN_IN, P1_EAX_REG_15__SCAN_IN, P1_EAX_REG_14__SCAN_IN, P1_EAX_REG_13__SCAN_IN, P1_EAX_REG_12__SCAN_IN, P1_EAX_REG_11__SCAN_IN, P1_EAX_REG_10__SCAN_IN, P1_EAX_REG_9__SCAN_IN, P1_EAX_REG_8__SCAN_IN, P1_EAX_REG_7__SCAN_IN, P1_EAX_REG_6__SCAN_IN, P1_EAX_REG_5__SCAN_IN, P1_EAX_REG_4__SCAN_IN, P1_EAX_REG_3__SCAN_IN, P1_EAX_REG_2__SCAN_IN, P1_EAX_REG_1__SCAN_IN, P1_EAX_REG_0__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_0__SCAN_IN, P1_UWORD_REG_0__SCAN_IN, P1_UWORD_REG_1__SCAN_IN, P1_UWORD_REG_2__SCAN_IN, P1_UWORD_REG_3__SCAN_IN, P1_UWORD_REG_4__SCAN_IN, P1_UWORD_REG_5__SCAN_IN, P1_UWORD_REG_6__SCAN_IN, P1_UWORD_REG_7__SCAN_IN, P1_UWORD_REG_8__SCAN_IN, P1_UWORD_REG_9__SCAN_IN, P1_UWORD_REG_10__SCAN_IN, P1_UWORD_REG_11__SCAN_IN, P1_UWORD_REG_12__SCAN_IN, P1_UWORD_REG_13__SCAN_IN, P1_UWORD_REG_14__SCAN_IN, P1_LWORD_REG_0__SCAN_IN, P1_LWORD_REG_1__SCAN_IN, P1_LWORD_REG_2__SCAN_IN, P1_LWORD_REG_3__SCAN_IN, P1_LWORD_REG_4__SCAN_IN, P1_LWORD_REG_5__SCAN_IN, P1_LWORD_REG_6__SCAN_IN, P1_LWORD_REG_7__SCAN_IN, P1_LWORD_REG_8__SCAN_IN, P1_LWORD_REG_9__SCAN_IN, P1_LWORD_REG_10__SCAN_IN, P1_LWORD_REG_11__SCAN_IN, P1_LWORD_REG_12__SCAN_IN, P1_LWORD_REG_13__SCAN_IN, P1_LWORD_REG_14__SCAN_IN, P1_LWORD_REG_15__SCAN_IN, P1_PHYADDRPOINTER_REG_31__SCAN_IN, P1_PHYADDRPOINTER_REG_30__SCAN_IN, P1_PHYADDRPOINTER_REG_29__SCAN_IN, P1_PHYADDRPOINTER_REG_28__SCAN_IN, P1_PHYADDRPOINTER_REG_27__SCAN_IN, P1_PHYADDRPOINTER_REG_26__SCAN_IN, P1_PHYADDRPOINTER_REG_25__SCAN_IN, P1_PHYADDRPOINTER_REG_24__SCAN_IN, P1_PHYADDRPOINTER_REG_23__SCAN_IN, P1_PHYADDRPOINTER_REG_22__SCAN_IN, P1_PHYADDRPOINTER_REG_21__SCAN_IN, P1_PHYADDRPOINTER_REG_20__SCAN_IN, P1_PHYADDRPOINTER_REG_19__SCAN_IN, P1_PHYADDRPOINTER_REG_18__SCAN_IN, P1_PHYADDRPOINTER_REG_17__SCAN_IN, P1_PHYADDRPOINTER_REG_16__SCAN_IN, P1_PHYADDRPOINTER_REG_15__SCAN_IN, P1_PHYADDRPOINTER_REG_14__SCAN_IN, P1_PHYADDRPOINTER_REG_13__SCAN_IN, P1_PHYADDRPOINTER_REG_12__SCAN_IN, P1_PHYADDRPOINTER_REG_11__SCAN_IN, P1_PHYADDRPOINTER_REG_10__SCAN_IN, P1_PHYADDRPOINTER_REG_9__SCAN_IN, P1_PHYADDRPOINTER_REG_8__SCAN_IN, P1_PHYADDRPOINTER_REG_7__SCAN_IN, P1_PHYADDRPOINTER_REG_6__SCAN_IN, P1_PHYADDRPOINTER_REG_5__SCAN_IN, P1_PHYADDRPOINTER_REG_4__SCAN_IN, P1_PHYADDRPOINTER_REG_3__SCAN_IN, P1_PHYADDRPOINTER_REG_2__SCAN_IN, P1_PHYADDRPOINTER_REG_1__SCAN_IN, P1_PHYADDRPOINTER_REG_0__SCAN_IN, P1_INSTADDRPOINTER_REG_31__SCAN_IN, P1_INSTADDRPOINTER_REG_30__SCAN_IN, P1_INSTADDRPOINTER_REG_29__SCAN_IN, P1_INSTADDRPOINTER_REG_28__SCAN_IN, P1_INSTADDRPOINTER_REG_27__SCAN_IN, P1_INSTADDRPOINTER_REG_26__SCAN_IN, P1_INSTADDRPOINTER_REG_25__SCAN_IN, P1_INSTADDRPOINTER_REG_24__SCAN_IN, P1_INSTADDRPOINTER_REG_23__SCAN_IN, P1_INSTADDRPOINTER_REG_22__SCAN_IN, P1_INSTADDRPOINTER_REG_21__SCAN_IN, P1_INSTADDRPOINTER_REG_20__SCAN_IN, P1_INSTADDRPOINTER_REG_19__SCAN_IN, P1_INSTADDRPOINTER_REG_18__SCAN_IN, P1_INSTADDRPOINTER_REG_17__SCAN_IN, P1_INSTADDRPOINTER_REG_16__SCAN_IN, P1_INSTADDRPOINTER_REG_15__SCAN_IN, P1_INSTADDRPOINTER_REG_14__SCAN_IN, P1_INSTADDRPOINTER_REG_13__SCAN_IN, P1_INSTADDRPOINTER_REG_12__SCAN_IN, P1_INSTADDRPOINTER_REG_11__SCAN_IN, P1_INSTADDRPOINTER_REG_10__SCAN_IN, P1_INSTADDRPOINTER_REG_9__SCAN_IN, P1_INSTADDRPOINTER_REG_8__SCAN_IN, P1_INSTADDRPOINTER_REG_7__SCAN_IN, P1_INSTADDRPOINTER_REG_6__SCAN_IN, P1_INSTADDRPOINTER_REG_5__SCAN_IN, P1_INSTADDRPOINTER_REG_4__SCAN_IN, P1_INSTADDRPOINTER_REG_3__SCAN_IN, P1_INSTADDRPOINTER_REG_2__SCAN_IN, P1_INSTADDRPOINTER_REG_1__SCAN_IN, P1_INSTADDRPOINTER_REG_0__SCAN_IN, P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN, P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN, P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN, P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN, P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN, P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN, P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN, P1_INSTQUEUE_REG_0__0__SCAN_IN, P1_INSTQUEUE_REG_0__1__SCAN_IN, P1_INSTQUEUE_REG_0__2__SCAN_IN, P1_INSTQUEUE_REG_0__3__SCAN_IN, P1_INSTQUEUE_REG_0__4__SCAN_IN, P1_INSTQUEUE_REG_0__5__SCAN_IN, P1_INSTQUEUE_REG_0__6__SCAN_IN, P1_INSTQUEUE_REG_0__7__SCAN_IN, P1_INSTQUEUE_REG_1__0__SCAN_IN, P1_INSTQUEUE_REG_1__1__SCAN_IN, P1_INSTQUEUE_REG_1__2__SCAN_IN, P1_INSTQUEUE_REG_1__3__SCAN_IN, P1_INSTQUEUE_REG_1__4__SCAN_IN, P1_INSTQUEUE_REG_1__5__SCAN_IN, P1_INSTQUEUE_REG_1__6__SCAN_IN, P1_INSTQUEUE_REG_1__7__SCAN_IN, P1_INSTQUEUE_REG_2__0__SCAN_IN, P1_INSTQUEUE_REG_2__1__SCAN_IN, P1_INSTQUEUE_REG_2__2__SCAN_IN, P1_INSTQUEUE_REG_2__3__SCAN_IN, P1_INSTQUEUE_REG_2__4__SCAN_IN, P1_INSTQUEUE_REG_2__5__SCAN_IN, P1_INSTQUEUE_REG_2__6__SCAN_IN, P1_INSTQUEUE_REG_2__7__SCAN_IN, P1_INSTQUEUE_REG_3__0__SCAN_IN, P1_INSTQUEUE_REG_3__1__SCAN_IN, P1_INSTQUEUE_REG_3__2__SCAN_IN, P1_INSTQUEUE_REG_3__3__SCAN_IN, P1_INSTQUEUE_REG_3__4__SCAN_IN, P1_INSTQUEUE_REG_3__5__SCAN_IN, P1_INSTQUEUE_REG_3__6__SCAN_IN, P1_INSTQUEUE_REG_3__7__SCAN_IN, P1_INSTQUEUE_REG_4__0__SCAN_IN, BUF1_REG_0__SCAN_IN, BUF1_REG_1__SCAN_IN, BUF1_REG_2__SCAN_IN, BUF1_REG_3__SCAN_IN, BUF1_REG_4__SCAN_IN, BUF1_REG_5__SCAN_IN, BUF1_REG_6__SCAN_IN, BUF1_REG_7__SCAN_IN, BUF1_REG_8__SCAN_IN, BUF1_REG_9__SCAN_IN, BUF1_REG_10__SCAN_IN, BUF1_REG_11__SCAN_IN, BUF1_REG_12__SCAN_IN, BUF1_REG_13__SCAN_IN, BUF1_REG_14__SCAN_IN, BUF1_REG_15__SCAN_IN, BUF1_REG_16__SCAN_IN, BUF1_REG_17__SCAN_IN, BUF1_REG_18__SCAN_IN, BUF1_REG_19__SCAN_IN, BUF1_REG_20__SCAN_IN, BUF1_REG_21__SCAN_IN, BUF1_REG_22__SCAN_IN, BUF1_REG_23__SCAN_IN, BUF1_REG_24__SCAN_IN, BUF1_REG_25__SCAN_IN, BUF1_REG_26__SCAN_IN, BUF1_REG_27__SCAN_IN, BUF1_REG_28__SCAN_IN, BUF1_REG_29__SCAN_IN, BUF1_REG_30__SCAN_IN, BUF1_REG_31__SCAN_IN, BUF2_REG_0__SCAN_IN, BUF2_REG_1__SCAN_IN, BUF2_REG_2__SCAN_IN, BUF2_REG_3__SCAN_IN, BUF2_REG_4__SCAN_IN, BUF2_REG_5__SCAN_IN, BUF2_REG_6__SCAN_IN, BUF2_REG_7__SCAN_IN, BUF2_REG_8__SCAN_IN, BUF2_REG_9__SCAN_IN, BUF2_REG_10__SCAN_IN, BUF2_REG_11__SCAN_IN, BUF2_REG_12__SCAN_IN, BUF2_REG_13__SCAN_IN, BUF2_REG_14__SCAN_IN, BUF2_REG_15__SCAN_IN, BUF2_REG_16__SCAN_IN, BUF2_REG_17__SCAN_IN, BUF2_REG_18__SCAN_IN, BUF2_REG_19__SCAN_IN, BUF2_REG_20__SCAN_IN, BUF2_REG_21__SCAN_IN, BUF2_REG_22__SCAN_IN, BUF2_REG_23__SCAN_IN, BUF2_REG_24__SCAN_IN, BUF2_REG_25__SCAN_IN, BUF2_REG_26__SCAN_IN, BUF2_REG_27__SCAN_IN, BUF2_REG_28__SCAN_IN, BUF2_REG_29__SCAN_IN, BUF2_REG_30__SCAN_IN, BUF2_REG_31__SCAN_IN, READY12_REG_SCAN_IN, READY21_REG_SCAN_IN, READY22_REG_SCAN_IN, READY11_REG_SCAN_IN, P3_BE_N_REG_3__SCAN_IN, P3_BE_N_REG_2__SCAN_IN, P3_BE_N_REG_1__SCAN_IN, P3_BE_N_REG_0__SCAN_IN, P3_ADDRESS_REG_29__SCAN_IN, P3_ADDRESS_REG_28__SCAN_IN, P3_ADDRESS_REG_27__SCAN_IN, P3_ADDRESS_REG_26__SCAN_IN, P3_ADDRESS_REG_25__SCAN_IN, P3_ADDRESS_REG_24__SCAN_IN, P3_ADDRESS_REG_23__SCAN_IN, P3_ADDRESS_REG_22__SCAN_IN, P3_ADDRESS_REG_21__SCAN_IN, P3_ADDRESS_REG_20__SCAN_IN, P3_ADDRESS_REG_19__SCAN_IN, P3_ADDRESS_REG_18__SCAN_IN, P3_ADDRESS_REG_17__SCAN_IN, P3_ADDRESS_REG_16__SCAN_IN, P3_ADDRESS_REG_15__SCAN_IN, P3_ADDRESS_REG_14__SCAN_IN, P3_ADDRESS_REG_13__SCAN_IN, P3_ADDRESS_REG_12__SCAN_IN, P3_ADDRESS_REG_11__SCAN_IN, P3_ADDRESS_REG_10__SCAN_IN, P3_ADDRESS_REG_9__SCAN_IN, P3_ADDRESS_REG_8__SCAN_IN, P3_ADDRESS_REG_7__SCAN_IN, P3_ADDRESS_REG_6__SCAN_IN, P3_ADDRESS_REG_5__SCAN_IN, P3_ADDRESS_REG_4__SCAN_IN, P3_ADDRESS_REG_3__SCAN_IN, P3_ADDRESS_REG_2__SCAN_IN, P3_ADDRESS_REG_1__SCAN_IN, P3_ADDRESS_REG_0__SCAN_IN, P3_STATE_REG_2__SCAN_IN, P3_STATE_REG_1__SCAN_IN, P3_STATE_REG_0__SCAN_IN, P3_DATAWIDTH_REG_0__SCAN_IN, P3_DATAWIDTH_REG_1__SCAN_IN, P3_DATAWIDTH_REG_2__SCAN_IN, P3_DATAWIDTH_REG_3__SCAN_IN, P3_DATAWIDTH_REG_4__SCAN_IN, P3_DATAWIDTH_REG_5__SCAN_IN, P3_DATAWIDTH_REG_6__SCAN_IN, P3_DATAWIDTH_REG_7__SCAN_IN, P3_DATAWIDTH_REG_8__SCAN_IN, P3_DATAWIDTH_REG_9__SCAN_IN, P3_DATAWIDTH_REG_10__SCAN_IN, P3_DATAWIDTH_REG_11__SCAN_IN, P3_DATAWIDTH_REG_12__SCAN_IN, P3_DATAWIDTH_REG_13__SCAN_IN, P3_DATAWIDTH_REG_14__SCAN_IN, P3_DATAWIDTH_REG_15__SCAN_IN, P3_DATAWIDTH_REG_16__SCAN_IN, P3_DATAWIDTH_REG_17__SCAN_IN, P3_DATAWIDTH_REG_18__SCAN_IN, P3_DATAWIDTH_REG_19__SCAN_IN, P3_DATAWIDTH_REG_20__SCAN_IN, P3_DATAWIDTH_REG_21__SCAN_IN, P3_DATAWIDTH_REG_22__SCAN_IN, P3_DATAWIDTH_REG_23__SCAN_IN, P3_DATAWIDTH_REG_24__SCAN_IN, P3_DATAWIDTH_REG_25__SCAN_IN, P3_DATAWIDTH_REG_26__SCAN_IN, P3_DATAWIDTH_REG_27__SCAN_IN, P3_DATAWIDTH_REG_28__SCAN_IN, P3_DATAWIDTH_REG_29__SCAN_IN, P3_DATAWIDTH_REG_30__SCAN_IN, P3_DATAWIDTH_REG_31__SCAN_IN, P3_STATE2_REG_3__SCAN_IN, P3_STATE2_REG_2__SCAN_IN, P3_STATE2_REG_1__SCAN_IN, P3_STATE2_REG_0__SCAN_IN, P3_INSTQUEUE_REG_15__7__SCAN_IN, P3_INSTQUEUE_REG_15__6__SCAN_IN, P3_INSTQUEUE_REG_15__5__SCAN_IN, P3_INSTQUEUE_REG_15__4__SCAN_IN, P3_INSTQUEUE_REG_15__3__SCAN_IN, P3_INSTQUEUE_REG_15__2__SCAN_IN, P3_INSTQUEUE_REG_15__1__SCAN_IN, P3_INSTQUEUE_REG_15__0__SCAN_IN, P3_INSTQUEUE_REG_14__7__SCAN_IN, P3_INSTQUEUE_REG_14__6__SCAN_IN, P3_INSTQUEUE_REG_14__5__SCAN_IN, P3_INSTQUEUE_REG_14__4__SCAN_IN, P3_INSTQUEUE_REG_14__3__SCAN_IN, P3_INSTQUEUE_REG_14__2__SCAN_IN, P3_INSTQUEUE_REG_14__1__SCAN_IN, P3_INSTQUEUE_REG_14__0__SCAN_IN, P3_INSTQUEUE_REG_13__7__SCAN_IN, P3_INSTQUEUE_REG_13__6__SCAN_IN, P3_INSTQUEUE_REG_13__5__SCAN_IN, P3_INSTQUEUE_REG_13__4__SCAN_IN, P3_INSTQUEUE_REG_13__3__SCAN_IN, P3_INSTQUEUE_REG_13__2__SCAN_IN, P3_INSTQUEUE_REG_13__1__SCAN_IN, P3_INSTQUEUE_REG_13__0__SCAN_IN, P3_INSTQUEUE_REG_12__7__SCAN_IN, P3_INSTQUEUE_REG_12__6__SCAN_IN, P3_INSTQUEUE_REG_12__5__SCAN_IN, P3_INSTQUEUE_REG_12__4__SCAN_IN, P3_INSTQUEUE_REG_12__3__SCAN_IN, P3_INSTQUEUE_REG_12__2__SCAN_IN, P3_INSTQUEUE_REG_12__1__SCAN_IN, P3_INSTQUEUE_REG_12__0__SCAN_IN, P3_INSTQUEUE_REG_11__7__SCAN_IN, P3_INSTQUEUE_REG_11__6__SCAN_IN, P3_INSTQUEUE_REG_11__5__SCAN_IN, P3_INSTQUEUE_REG_11__4__SCAN_IN, P3_INSTQUEUE_REG_11__3__SCAN_IN, P3_INSTQUEUE_REG_11__2__SCAN_IN, P3_INSTQUEUE_REG_11__1__SCAN_IN, P3_INSTQUEUE_REG_11__0__SCAN_IN, P3_INSTQUEUE_REG_10__7__SCAN_IN, P3_INSTQUEUE_REG_10__6__SCAN_IN, P3_INSTQUEUE_REG_10__5__SCAN_IN, P3_INSTQUEUE_REG_10__4__SCAN_IN, P3_INSTQUEUE_REG_10__3__SCAN_IN, P3_INSTQUEUE_REG_10__2__SCAN_IN, P3_INSTQUEUE_REG_10__1__SCAN_IN, P3_INSTQUEUE_REG_10__0__SCAN_IN, P3_INSTQUEUE_REG_9__7__SCAN_IN, P3_INSTQUEUE_REG_9__6__SCAN_IN, P3_INSTQUEUE_REG_9__5__SCAN_IN, P3_INSTQUEUE_REG_9__4__SCAN_IN, P3_INSTQUEUE_REG_9__3__SCAN_IN, P3_INSTQUEUE_REG_9__2__SCAN_IN, P3_INSTQUEUE_REG_9__1__SCAN_IN, P3_INSTQUEUE_REG_9__0__SCAN_IN, P3_INSTQUEUE_REG_8__7__SCAN_IN, P3_INSTQUEUE_REG_8__6__SCAN_IN, P3_INSTQUEUE_REG_8__5__SCAN_IN, P3_INSTQUEUE_REG_8__4__SCAN_IN, P3_INSTQUEUE_REG_8__3__SCAN_IN, P3_INSTQUEUE_REG_8__2__SCAN_IN, P3_INSTQUEUE_REG_8__1__SCAN_IN, P3_INSTQUEUE_REG_8__0__SCAN_IN, P3_INSTQUEUE_REG_7__7__SCAN_IN, P3_INSTQUEUE_REG_7__6__SCAN_IN, P3_INSTQUEUE_REG_7__5__SCAN_IN, P3_INSTQUEUE_REG_7__4__SCAN_IN, P3_INSTQUEUE_REG_7__3__SCAN_IN, P3_INSTQUEUE_REG_7__2__SCAN_IN, P3_INSTQUEUE_REG_7__1__SCAN_IN, P3_INSTQUEUE_REG_7__0__SCAN_IN, P3_INSTQUEUE_REG_6__7__SCAN_IN, P3_INSTQUEUE_REG_6__6__SCAN_IN, P3_INSTQUEUE_REG_6__5__SCAN_IN, P3_INSTQUEUE_REG_6__4__SCAN_IN, P3_INSTQUEUE_REG_6__3__SCAN_IN, P3_INSTQUEUE_REG_6__2__SCAN_IN, P3_INSTQUEUE_REG_6__1__SCAN_IN, P3_INSTQUEUE_REG_6__0__SCAN_IN, P3_INSTQUEUE_REG_5__7__SCAN_IN, P3_INSTQUEUE_REG_5__6__SCAN_IN, P3_INSTQUEUE_REG_5__5__SCAN_IN, P3_INSTQUEUE_REG_5__4__SCAN_IN, P3_INSTQUEUE_REG_5__3__SCAN_IN, P3_INSTQUEUE_REG_5__2__SCAN_IN, P3_INSTQUEUE_REG_5__1__SCAN_IN, P3_INSTQUEUE_REG_5__0__SCAN_IN, P3_INSTQUEUE_REG_4__7__SCAN_IN, P3_INSTQUEUE_REG_4__6__SCAN_IN, P3_INSTQUEUE_REG_4__5__SCAN_IN, P3_INSTQUEUE_REG_4__4__SCAN_IN, P3_INSTQUEUE_REG_4__3__SCAN_IN, P3_INSTQUEUE_REG_4__2__SCAN_IN, P3_INSTQUEUE_REG_4__1__SCAN_IN, P3_INSTQUEUE_REG_4__0__SCAN_IN, P3_INSTQUEUE_REG_3__7__SCAN_IN, P3_INSTQUEUE_REG_3__6__SCAN_IN, P3_INSTQUEUE_REG_3__5__SCAN_IN, P3_INSTQUEUE_REG_3__4__SCAN_IN, P3_INSTQUEUE_REG_3__3__SCAN_IN, P3_INSTQUEUE_REG_3__2__SCAN_IN, P3_INSTQUEUE_REG_3__1__SCAN_IN, P3_INSTQUEUE_REG_3__0__SCAN_IN, P3_INSTQUEUE_REG_2__7__SCAN_IN, P3_INSTQUEUE_REG_2__6__SCAN_IN, P3_INSTQUEUE_REG_2__5__SCAN_IN, P3_INSTQUEUE_REG_2__4__SCAN_IN, P3_INSTQUEUE_REG_2__3__SCAN_IN, P3_INSTQUEUE_REG_2__2__SCAN_IN, P3_INSTQUEUE_REG_2__1__SCAN_IN, P3_INSTQUEUE_REG_2__0__SCAN_IN, P3_INSTQUEUE_REG_1__7__SCAN_IN, P3_INSTQUEUE_REG_1__6__SCAN_IN, P3_INSTQUEUE_REG_1__5__SCAN_IN, P3_INSTQUEUE_REG_1__4__SCAN_IN, P3_INSTQUEUE_REG_1__3__SCAN_IN, P3_INSTQUEUE_REG_1__2__SCAN_IN, P3_INSTQUEUE_REG_1__1__SCAN_IN, P3_INSTQUEUE_REG_1__0__SCAN_IN, P3_INSTQUEUE_REG_0__7__SCAN_IN, P3_INSTQUEUE_REG_0__6__SCAN_IN, P3_INSTQUEUE_REG_0__5__SCAN_IN, P3_INSTQUEUE_REG_0__4__SCAN_IN, P3_INSTQUEUE_REG_0__3__SCAN_IN, P3_INSTQUEUE_REG_0__2__SCAN_IN, P3_INSTQUEUE_REG_0__1__SCAN_IN, P3_INSTQUEUE_REG_0__0__SCAN_IN, P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN, P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN, P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN, P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN, P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN, P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN, P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN, P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P3_INSTADDRPOINTER_REG_0__SCAN_IN, P3_INSTADDRPOINTER_REG_1__SCAN_IN, P3_INSTADDRPOINTER_REG_2__SCAN_IN, P3_INSTADDRPOINTER_REG_3__SCAN_IN, P3_INSTADDRPOINTER_REG_4__SCAN_IN, P3_INSTADDRPOINTER_REG_5__SCAN_IN, P3_INSTADDRPOINTER_REG_6__SCAN_IN, P3_INSTADDRPOINTER_REG_7__SCAN_IN, P3_INSTADDRPOINTER_REG_8__SCAN_IN, P3_INSTADDRPOINTER_REG_9__SCAN_IN, P3_INSTADDRPOINTER_REG_10__SCAN_IN, P3_INSTADDRPOINTER_REG_11__SCAN_IN, P3_INSTADDRPOINTER_REG_12__SCAN_IN, P3_INSTADDRPOINTER_REG_13__SCAN_IN, P3_INSTADDRPOINTER_REG_14__SCAN_IN, P3_INSTADDRPOINTER_REG_15__SCAN_IN, P3_INSTADDRPOINTER_REG_16__SCAN_IN, P3_INSTADDRPOINTER_REG_17__SCAN_IN, P3_INSTADDRPOINTER_REG_18__SCAN_IN, P3_INSTADDRPOINTER_REG_19__SCAN_IN, P3_INSTADDRPOINTER_REG_20__SCAN_IN, P3_INSTADDRPOINTER_REG_21__SCAN_IN, P3_INSTADDRPOINTER_REG_22__SCAN_IN, P3_INSTADDRPOINTER_REG_23__SCAN_IN, P3_INSTADDRPOINTER_REG_24__SCAN_IN, P3_INSTADDRPOINTER_REG_25__SCAN_IN, P3_INSTADDRPOINTER_REG_26__SCAN_IN, P3_INSTADDRPOINTER_REG_27__SCAN_IN, P3_INSTADDRPOINTER_REG_28__SCAN_IN, P3_INSTADDRPOINTER_REG_29__SCAN_IN, P3_INSTADDRPOINTER_REG_30__SCAN_IN, P3_INSTADDRPOINTER_REG_31__SCAN_IN, P3_PHYADDRPOINTER_REG_0__SCAN_IN, P3_PHYADDRPOINTER_REG_1__SCAN_IN, P3_PHYADDRPOINTER_REG_2__SCAN_IN, P3_PHYADDRPOINTER_REG_3__SCAN_IN, P3_PHYADDRPOINTER_REG_4__SCAN_IN, P3_PHYADDRPOINTER_REG_5__SCAN_IN, P3_PHYADDRPOINTER_REG_6__SCAN_IN, P3_PHYADDRPOINTER_REG_7__SCAN_IN, P3_PHYADDRPOINTER_REG_8__SCAN_IN, P3_PHYADDRPOINTER_REG_9__SCAN_IN, P3_PHYADDRPOINTER_REG_10__SCAN_IN, P3_PHYADDRPOINTER_REG_11__SCAN_IN, P3_PHYADDRPOINTER_REG_12__SCAN_IN, P3_PHYADDRPOINTER_REG_13__SCAN_IN, P3_PHYADDRPOINTER_REG_14__SCAN_IN, P3_PHYADDRPOINTER_REG_15__SCAN_IN, P3_PHYADDRPOINTER_REG_16__SCAN_IN, P3_PHYADDRPOINTER_REG_17__SCAN_IN, P3_PHYADDRPOINTER_REG_18__SCAN_IN, P3_PHYADDRPOINTER_REG_19__SCAN_IN, P3_PHYADDRPOINTER_REG_20__SCAN_IN, P3_PHYADDRPOINTER_REG_21__SCAN_IN, P3_PHYADDRPOINTER_REG_22__SCAN_IN, P3_PHYADDRPOINTER_REG_23__SCAN_IN, P3_PHYADDRPOINTER_REG_24__SCAN_IN, P3_PHYADDRPOINTER_REG_25__SCAN_IN, P3_PHYADDRPOINTER_REG_26__SCAN_IN, P3_PHYADDRPOINTER_REG_27__SCAN_IN, P3_PHYADDRPOINTER_REG_28__SCAN_IN, P3_PHYADDRPOINTER_REG_29__SCAN_IN, P3_PHYADDRPOINTER_REG_30__SCAN_IN, P3_PHYADDRPOINTER_REG_31__SCAN_IN, P3_LWORD_REG_15__SCAN_IN, P3_LWORD_REG_14__SCAN_IN, P3_LWORD_REG_13__SCAN_IN, P3_LWORD_REG_12__SCAN_IN, P3_LWORD_REG_11__SCAN_IN, P3_LWORD_REG_10__SCAN_IN, P3_LWORD_REG_9__SCAN_IN, P3_LWORD_REG_8__SCAN_IN, P3_LWORD_REG_7__SCAN_IN, P3_LWORD_REG_6__SCAN_IN, P3_LWORD_REG_5__SCAN_IN, P3_LWORD_REG_4__SCAN_IN, P3_LWORD_REG_3__SCAN_IN, P3_LWORD_REG_2__SCAN_IN, P3_LWORD_REG_1__SCAN_IN, P3_LWORD_REG_0__SCAN_IN, P3_UWORD_REG_14__SCAN_IN, P3_UWORD_REG_13__SCAN_IN, P3_UWORD_REG_12__SCAN_IN, P3_UWORD_REG_11__SCAN_IN, P3_UWORD_REG_10__SCAN_IN, P3_UWORD_REG_9__SCAN_IN, P3_UWORD_REG_8__SCAN_IN, P3_UWORD_REG_7__SCAN_IN, P3_UWORD_REG_6__SCAN_IN, P3_UWORD_REG_5__SCAN_IN, P3_UWORD_REG_4__SCAN_IN, P3_UWORD_REG_3__SCAN_IN, P3_UWORD_REG_2__SCAN_IN, P3_UWORD_REG_1__SCAN_IN, P3_UWORD_REG_0__SCAN_IN, P3_DATAO_REG_0__SCAN_IN, P3_DATAO_REG_1__SCAN_IN, P3_DATAO_REG_2__SCAN_IN, P3_DATAO_REG_3__SCAN_IN, P3_DATAO_REG_4__SCAN_IN, P3_DATAO_REG_5__SCAN_IN, P3_DATAO_REG_6__SCAN_IN, P3_DATAO_REG_7__SCAN_IN, P3_DATAO_REG_8__SCAN_IN, P3_DATAO_REG_9__SCAN_IN, P3_DATAO_REG_10__SCAN_IN, P3_DATAO_REG_11__SCAN_IN, P3_DATAO_REG_12__SCAN_IN, P3_DATAO_REG_13__SCAN_IN, P3_DATAO_REG_14__SCAN_IN, P3_DATAO_REG_15__SCAN_IN, P3_DATAO_REG_16__SCAN_IN, P3_DATAO_REG_17__SCAN_IN, P3_DATAO_REG_18__SCAN_IN, P3_DATAO_REG_19__SCAN_IN, P3_DATAO_REG_20__SCAN_IN, P3_DATAO_REG_21__SCAN_IN, P3_DATAO_REG_22__SCAN_IN, P3_DATAO_REG_23__SCAN_IN, P3_DATAO_REG_24__SCAN_IN, P3_DATAO_REG_25__SCAN_IN, P3_DATAO_REG_26__SCAN_IN, P3_DATAO_REG_27__SCAN_IN, P3_DATAO_REG_28__SCAN_IN, P3_DATAO_REG_29__SCAN_IN, P3_DATAO_REG_30__SCAN_IN, P3_DATAO_REG_31__SCAN_IN, P3_EAX_REG_0__SCAN_IN, P3_EAX_REG_1__SCAN_IN, P3_EAX_REG_2__SCAN_IN, P3_EAX_REG_3__SCAN_IN, P3_EAX_REG_4__SCAN_IN, P3_EAX_REG_5__SCAN_IN, P3_EAX_REG_6__SCAN_IN, P3_EAX_REG_7__SCAN_IN, P3_EAX_REG_8__SCAN_IN, P3_EAX_REG_9__SCAN_IN, P3_EAX_REG_10__SCAN_IN, P3_EAX_REG_11__SCAN_IN, P3_EAX_REG_12__SCAN_IN, P3_EAX_REG_13__SCAN_IN, P3_EAX_REG_14__SCAN_IN, P3_EAX_REG_15__SCAN_IN, P3_EAX_REG_16__SCAN_IN, P3_EAX_REG_17__SCAN_IN, P3_EAX_REG_18__SCAN_IN, P3_EAX_REG_19__SCAN_IN, P3_EAX_REG_20__SCAN_IN, P3_EAX_REG_21__SCAN_IN, P3_EAX_REG_22__SCAN_IN, P3_EAX_REG_23__SCAN_IN, P3_EAX_REG_24__SCAN_IN, P3_EAX_REG_25__SCAN_IN, P3_EAX_REG_26__SCAN_IN, P3_EAX_REG_27__SCAN_IN, P3_EAX_REG_28__SCAN_IN, P3_EAX_REG_29__SCAN_IN, P3_EAX_REG_30__SCAN_IN, P3_EAX_REG_31__SCAN_IN, P3_EBX_REG_0__SCAN_IN, P3_EBX_REG_1__SCAN_IN, P3_EBX_REG_2__SCAN_IN, P3_EBX_REG_3__SCAN_IN, P3_EBX_REG_4__SCAN_IN, P3_EBX_REG_5__SCAN_IN, P3_EBX_REG_6__SCAN_IN, P3_EBX_REG_7__SCAN_IN, P3_EBX_REG_8__SCAN_IN, P3_EBX_REG_9__SCAN_IN, P3_EBX_REG_10__SCAN_IN, P3_EBX_REG_11__SCAN_IN, P3_EBX_REG_12__SCAN_IN, P3_EBX_REG_13__SCAN_IN, P3_EBX_REG_14__SCAN_IN, P3_EBX_REG_15__SCAN_IN, P3_EBX_REG_16__SCAN_IN, P3_EBX_REG_17__SCAN_IN, P3_EBX_REG_18__SCAN_IN, P3_EBX_REG_19__SCAN_IN, P3_EBX_REG_20__SCAN_IN, P3_EBX_REG_21__SCAN_IN, P3_EBX_REG_22__SCAN_IN, P3_EBX_REG_23__SCAN_IN, P3_EBX_REG_24__SCAN_IN, P3_EBX_REG_25__SCAN_IN, P3_EBX_REG_26__SCAN_IN, P3_EBX_REG_27__SCAN_IN, P3_EBX_REG_28__SCAN_IN, P3_EBX_REG_29__SCAN_IN, P3_EBX_REG_30__SCAN_IN, P3_EBX_REG_31__SCAN_IN, P3_REIP_REG_0__SCAN_IN, P3_REIP_REG_1__SCAN_IN, P3_REIP_REG_2__SCAN_IN, P3_REIP_REG_3__SCAN_IN, P3_REIP_REG_4__SCAN_IN, P3_REIP_REG_5__SCAN_IN, P3_REIP_REG_6__SCAN_IN, P3_REIP_REG_7__SCAN_IN, P3_REIP_REG_8__SCAN_IN, P3_REIP_REG_9__SCAN_IN, P3_REIP_REG_10__SCAN_IN, P3_REIP_REG_11__SCAN_IN, P3_REIP_REG_12__SCAN_IN, P3_REIP_REG_13__SCAN_IN, P3_REIP_REG_14__SCAN_IN, P3_REIP_REG_15__SCAN_IN, P3_REIP_REG_16__SCAN_IN, P3_REIP_REG_17__SCAN_IN, P3_REIP_REG_18__SCAN_IN, P3_REIP_REG_19__SCAN_IN, P3_REIP_REG_20__SCAN_IN, P3_REIP_REG_21__SCAN_IN, P3_REIP_REG_22__SCAN_IN, P3_REIP_REG_23__SCAN_IN, P3_REIP_REG_24__SCAN_IN, P3_REIP_REG_25__SCAN_IN, P3_REIP_REG_26__SCAN_IN, P3_REIP_REG_27__SCAN_IN, P3_REIP_REG_28__SCAN_IN, P3_REIP_REG_29__SCAN_IN, P3_REIP_REG_30__SCAN_IN, P3_REIP_REG_31__SCAN_IN, P3_BYTEENABLE_REG_3__SCAN_IN, P3_BYTEENABLE_REG_2__SCAN_IN, P3_BYTEENABLE_REG_1__SCAN_IN, P3_BYTEENABLE_REG_0__SCAN_IN, P3_W_R_N_REG_SCAN_IN, P3_FLUSH_REG_SCAN_IN, P3_MORE_REG_SCAN_IN, P3_STATEBS16_REG_SCAN_IN, P3_REQUESTPENDING_REG_SCAN_IN, P3_D_C_N_REG_SCAN_IN, P3_M_IO_N_REG_SCAN_IN, P3_CODEFETCH_REG_SCAN_IN, P3_ADS_N_REG_SCAN_IN, P3_READREQUEST_REG_SCAN_IN, P3_MEMORYFETCH_REG_SCAN_IN, P2_BE_N_REG_3__SCAN_IN, P2_BE_N_REG_2__SCAN_IN, P2_BE_N_REG_1__SCAN_IN, P2_BE_N_REG_0__SCAN_IN, P2_ADDRESS_REG_29__SCAN_IN, P2_ADDRESS_REG_28__SCAN_IN, P2_ADDRESS_REG_27__SCAN_IN, P2_ADDRESS_REG_26__SCAN_IN, P2_ADDRESS_REG_25__SCAN_IN, P2_ADDRESS_REG_24__SCAN_IN, P2_ADDRESS_REG_23__SCAN_IN, P2_ADDRESS_REG_22__SCAN_IN, P2_ADDRESS_REG_21__SCAN_IN, P2_ADDRESS_REG_20__SCAN_IN, P2_ADDRESS_REG_19__SCAN_IN, P2_ADDRESS_REG_18__SCAN_IN, P2_ADDRESS_REG_17__SCAN_IN, P2_ADDRESS_REG_16__SCAN_IN, P2_ADDRESS_REG_15__SCAN_IN, P2_ADDRESS_REG_14__SCAN_IN, P2_ADDRESS_REG_13__SCAN_IN, P2_ADDRESS_REG_12__SCAN_IN, P2_ADDRESS_REG_11__SCAN_IN, P2_ADDRESS_REG_10__SCAN_IN, P2_ADDRESS_REG_9__SCAN_IN, P2_ADDRESS_REG_8__SCAN_IN, P2_ADDRESS_REG_7__SCAN_IN, P2_ADDRESS_REG_6__SCAN_IN, P2_ADDRESS_REG_5__SCAN_IN, P2_ADDRESS_REG_4__SCAN_IN, P2_ADDRESS_REG_3__SCAN_IN, P2_ADDRESS_REG_2__SCAN_IN, P2_ADDRESS_REG_1__SCAN_IN, P2_ADDRESS_REG_0__SCAN_IN, P2_STATE_REG_2__SCAN_IN, P2_STATE_REG_1__SCAN_IN, P2_STATE_REG_0__SCAN_IN, P2_DATAWIDTH_REG_0__SCAN_IN, P2_DATAWIDTH_REG_1__SCAN_IN, P2_DATAWIDTH_REG_2__SCAN_IN, P2_DATAWIDTH_REG_3__SCAN_IN, P2_DATAWIDTH_REG_4__SCAN_IN, P2_DATAWIDTH_REG_5__SCAN_IN, P2_DATAWIDTH_REG_6__SCAN_IN, P2_DATAWIDTH_REG_7__SCAN_IN, P2_DATAWIDTH_REG_8__SCAN_IN, P2_DATAWIDTH_REG_9__SCAN_IN, P2_DATAWIDTH_REG_10__SCAN_IN, P2_DATAWIDTH_REG_11__SCAN_IN, P2_DATAWIDTH_REG_12__SCAN_IN, P2_DATAWIDTH_REG_13__SCAN_IN, P2_DATAWIDTH_REG_14__SCAN_IN, P2_DATAWIDTH_REG_15__SCAN_IN, P2_DATAWIDTH_REG_16__SCAN_IN, P2_DATAWIDTH_REG_17__SCAN_IN, P2_DATAWIDTH_REG_18__SCAN_IN, P2_DATAWIDTH_REG_19__SCAN_IN, P2_DATAWIDTH_REG_20__SCAN_IN, P2_DATAWIDTH_REG_21__SCAN_IN, P2_DATAWIDTH_REG_22__SCAN_IN, P2_DATAWIDTH_REG_23__SCAN_IN, P2_DATAWIDTH_REG_24__SCAN_IN, P2_DATAWIDTH_REG_25__SCAN_IN, P2_DATAWIDTH_REG_26__SCAN_IN, P2_DATAWIDTH_REG_27__SCAN_IN, P2_DATAWIDTH_REG_28__SCAN_IN, P2_DATAWIDTH_REG_29__SCAN_IN, P2_DATAWIDTH_REG_30__SCAN_IN, P2_DATAWIDTH_REG_31__SCAN_IN, P2_STATE2_REG_3__SCAN_IN, P2_STATE2_REG_2__SCAN_IN, P2_STATE2_REG_1__SCAN_IN, P2_STATE2_REG_0__SCAN_IN, P2_INSTQUEUE_REG_15__7__SCAN_IN, P2_INSTQUEUE_REG_15__6__SCAN_IN, P2_INSTQUEUE_REG_15__5__SCAN_IN, P2_INSTQUEUE_REG_15__4__SCAN_IN, P2_INSTQUEUE_REG_15__3__SCAN_IN, P2_INSTQUEUE_REG_15__2__SCAN_IN, P2_INSTQUEUE_REG_15__1__SCAN_IN, P2_INSTQUEUE_REG_15__0__SCAN_IN, P2_INSTQUEUE_REG_14__7__SCAN_IN, P2_INSTQUEUE_REG_14__6__SCAN_IN, P2_INSTQUEUE_REG_14__5__SCAN_IN, P2_INSTQUEUE_REG_14__4__SCAN_IN, P2_INSTQUEUE_REG_14__3__SCAN_IN, P2_INSTQUEUE_REG_14__2__SCAN_IN, P2_INSTQUEUE_REG_14__1__SCAN_IN, P2_INSTQUEUE_REG_14__0__SCAN_IN, P2_INSTQUEUE_REG_13__7__SCAN_IN, P2_INSTQUEUE_REG_13__6__SCAN_IN, P2_INSTQUEUE_REG_13__5__SCAN_IN, P2_INSTQUEUE_REG_13__4__SCAN_IN, P2_INSTQUEUE_REG_13__3__SCAN_IN, P2_INSTQUEUE_REG_13__2__SCAN_IN, P2_INSTQUEUE_REG_13__1__SCAN_IN, P2_INSTQUEUE_REG_13__0__SCAN_IN, P2_INSTQUEUE_REG_12__7__SCAN_IN, P2_INSTQUEUE_REG_12__6__SCAN_IN, P2_INSTQUEUE_REG_12__5__SCAN_IN, P2_INSTQUEUE_REG_12__4__SCAN_IN, P2_INSTQUEUE_REG_12__3__SCAN_IN, P2_INSTQUEUE_REG_12__2__SCAN_IN, P2_INSTQUEUE_REG_12__1__SCAN_IN, P2_INSTQUEUE_REG_12__0__SCAN_IN, P2_INSTQUEUE_REG_11__7__SCAN_IN, P2_INSTQUEUE_REG_11__6__SCAN_IN, P2_INSTQUEUE_REG_11__5__SCAN_IN, P2_INSTQUEUE_REG_11__4__SCAN_IN, P2_INSTQUEUE_REG_11__3__SCAN_IN, P2_INSTQUEUE_REG_11__2__SCAN_IN, P2_INSTQUEUE_REG_11__1__SCAN_IN, P2_INSTQUEUE_REG_11__0__SCAN_IN, P2_INSTQUEUE_REG_10__7__SCAN_IN, P2_INSTQUEUE_REG_10__6__SCAN_IN, P2_INSTQUEUE_REG_10__5__SCAN_IN, P2_INSTQUEUE_REG_10__4__SCAN_IN, P2_INSTQUEUE_REG_10__3__SCAN_IN, P2_INSTQUEUE_REG_10__2__SCAN_IN, P2_INSTQUEUE_REG_10__1__SCAN_IN, P2_INSTQUEUE_REG_10__0__SCAN_IN, P2_INSTQUEUE_REG_9__7__SCAN_IN, P2_INSTQUEUE_REG_9__6__SCAN_IN, P2_INSTQUEUE_REG_9__5__SCAN_IN, P2_INSTQUEUE_REG_9__4__SCAN_IN, P2_INSTQUEUE_REG_9__3__SCAN_IN, P2_INSTQUEUE_REG_9__2__SCAN_IN, P2_INSTQUEUE_REG_9__1__SCAN_IN, P2_INSTQUEUE_REG_9__0__SCAN_IN, P2_INSTQUEUE_REG_8__7__SCAN_IN, P2_INSTQUEUE_REG_8__6__SCAN_IN, P2_INSTQUEUE_REG_8__5__SCAN_IN, P2_INSTQUEUE_REG_8__4__SCAN_IN, P2_INSTQUEUE_REG_8__3__SCAN_IN, P2_INSTQUEUE_REG_8__2__SCAN_IN, P2_INSTQUEUE_REG_8__1__SCAN_IN, P2_INSTQUEUE_REG_8__0__SCAN_IN, P2_INSTQUEUE_REG_7__7__SCAN_IN, P2_INSTQUEUE_REG_7__6__SCAN_IN, P2_INSTQUEUE_REG_7__5__SCAN_IN, P2_INSTQUEUE_REG_7__4__SCAN_IN, P2_INSTQUEUE_REG_7__3__SCAN_IN, P2_INSTQUEUE_REG_7__2__SCAN_IN, P2_INSTQUEUE_REG_7__1__SCAN_IN, P2_INSTQUEUE_REG_7__0__SCAN_IN, P2_INSTQUEUE_REG_6__7__SCAN_IN, P2_INSTQUEUE_REG_6__6__SCAN_IN, P2_INSTQUEUE_REG_6__5__SCAN_IN, P2_INSTQUEUE_REG_6__4__SCAN_IN, P2_INSTQUEUE_REG_6__3__SCAN_IN, P2_INSTQUEUE_REG_6__2__SCAN_IN, P2_INSTQUEUE_REG_6__1__SCAN_IN, P2_INSTQUEUE_REG_6__0__SCAN_IN, P2_INSTQUEUE_REG_5__7__SCAN_IN, P2_INSTQUEUE_REG_5__6__SCAN_IN, P2_INSTQUEUE_REG_5__5__SCAN_IN, P2_INSTQUEUE_REG_5__4__SCAN_IN, P2_INSTQUEUE_REG_5__3__SCAN_IN, P2_INSTQUEUE_REG_5__2__SCAN_IN, P2_INSTQUEUE_REG_5__1__SCAN_IN, P2_INSTQUEUE_REG_5__0__SCAN_IN, P2_INSTQUEUE_REG_4__7__SCAN_IN, P2_INSTQUEUE_REG_4__6__SCAN_IN, P2_INSTQUEUE_REG_4__5__SCAN_IN, P2_INSTQUEUE_REG_4__4__SCAN_IN, P2_INSTQUEUE_REG_4__3__SCAN_IN, P2_INSTQUEUE_REG_4__2__SCAN_IN, P2_INSTQUEUE_REG_4__1__SCAN_IN, P2_INSTQUEUE_REG_4__0__SCAN_IN, P2_INSTQUEUE_REG_3__7__SCAN_IN, P2_INSTQUEUE_REG_3__6__SCAN_IN, P2_INSTQUEUE_REG_3__5__SCAN_IN, P2_INSTQUEUE_REG_3__4__SCAN_IN, P2_INSTQUEUE_REG_3__3__SCAN_IN, P2_INSTQUEUE_REG_3__2__SCAN_IN, P2_INSTQUEUE_REG_3__1__SCAN_IN, P2_INSTQUEUE_REG_3__0__SCAN_IN, P2_INSTQUEUE_REG_2__7__SCAN_IN, P2_INSTQUEUE_REG_2__6__SCAN_IN, P2_INSTQUEUE_REG_2__5__SCAN_IN, P2_INSTQUEUE_REG_2__4__SCAN_IN, P2_INSTQUEUE_REG_2__3__SCAN_IN, P2_INSTQUEUE_REG_2__2__SCAN_IN, P2_INSTQUEUE_REG_2__1__SCAN_IN, P2_INSTQUEUE_REG_2__0__SCAN_IN, P2_INSTQUEUE_REG_1__7__SCAN_IN, P2_INSTQUEUE_REG_1__6__SCAN_IN, P2_INSTQUEUE_REG_1__5__SCAN_IN, P2_INSTQUEUE_REG_1__4__SCAN_IN, P2_INSTQUEUE_REG_1__3__SCAN_IN, P2_INSTQUEUE_REG_1__2__SCAN_IN, P2_INSTQUEUE_REG_1__1__SCAN_IN, P2_INSTQUEUE_REG_1__0__SCAN_IN, P2_INSTQUEUE_REG_0__7__SCAN_IN, P2_INSTQUEUE_REG_0__6__SCAN_IN, P2_INSTQUEUE_REG_0__5__SCAN_IN, P2_INSTQUEUE_REG_0__4__SCAN_IN, P2_INSTQUEUE_REG_0__3__SCAN_IN, P2_INSTQUEUE_REG_0__2__SCAN_IN, P2_INSTQUEUE_REG_0__1__SCAN_IN, P2_INSTQUEUE_REG_0__0__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN, P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN, P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN, P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN, P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN, P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P2_INSTADDRPOINTER_REG_0__SCAN_IN, P2_INSTADDRPOINTER_REG_1__SCAN_IN, P2_INSTADDRPOINTER_REG_2__SCAN_IN, P2_INSTADDRPOINTER_REG_3__SCAN_IN, P2_INSTADDRPOINTER_REG_4__SCAN_IN, P2_INSTADDRPOINTER_REG_5__SCAN_IN, P2_INSTADDRPOINTER_REG_6__SCAN_IN, P2_INSTADDRPOINTER_REG_7__SCAN_IN, P2_INSTADDRPOINTER_REG_8__SCAN_IN, P2_INSTADDRPOINTER_REG_9__SCAN_IN, P2_INSTADDRPOINTER_REG_10__SCAN_IN, P2_INSTADDRPOINTER_REG_11__SCAN_IN, P2_INSTADDRPOINTER_REG_12__SCAN_IN, P2_INSTADDRPOINTER_REG_13__SCAN_IN, P2_INSTADDRPOINTER_REG_14__SCAN_IN, P2_INSTADDRPOINTER_REG_15__SCAN_IN, P2_INSTADDRPOINTER_REG_16__SCAN_IN, P2_INSTADDRPOINTER_REG_17__SCAN_IN, P2_INSTADDRPOINTER_REG_18__SCAN_IN, P2_INSTADDRPOINTER_REG_19__SCAN_IN, P2_INSTADDRPOINTER_REG_20__SCAN_IN, P2_INSTADDRPOINTER_REG_21__SCAN_IN, P2_INSTADDRPOINTER_REG_22__SCAN_IN, P2_INSTADDRPOINTER_REG_23__SCAN_IN, P2_INSTADDRPOINTER_REG_24__SCAN_IN, P2_INSTADDRPOINTER_REG_25__SCAN_IN, P2_INSTADDRPOINTER_REG_26__SCAN_IN, P2_INSTADDRPOINTER_REG_27__SCAN_IN, P2_INSTADDRPOINTER_REG_28__SCAN_IN, P2_INSTADDRPOINTER_REG_29__SCAN_IN, P2_INSTADDRPOINTER_REG_30__SCAN_IN, P2_INSTADDRPOINTER_REG_31__SCAN_IN, P2_PHYADDRPOINTER_REG_0__SCAN_IN, P2_PHYADDRPOINTER_REG_1__SCAN_IN, P2_PHYADDRPOINTER_REG_2__SCAN_IN, P2_PHYADDRPOINTER_REG_3__SCAN_IN, P2_PHYADDRPOINTER_REG_4__SCAN_IN, P2_PHYADDRPOINTER_REG_5__SCAN_IN, P2_PHYADDRPOINTER_REG_6__SCAN_IN, P2_PHYADDRPOINTER_REG_7__SCAN_IN, P2_PHYADDRPOINTER_REG_8__SCAN_IN, P2_PHYADDRPOINTER_REG_9__SCAN_IN, P2_PHYADDRPOINTER_REG_10__SCAN_IN, P2_PHYADDRPOINTER_REG_11__SCAN_IN, P2_PHYADDRPOINTER_REG_12__SCAN_IN, P2_PHYADDRPOINTER_REG_13__SCAN_IN, P2_PHYADDRPOINTER_REG_14__SCAN_IN, P2_PHYADDRPOINTER_REG_15__SCAN_IN, P2_PHYADDRPOINTER_REG_16__SCAN_IN, P2_PHYADDRPOINTER_REG_17__SCAN_IN, P2_PHYADDRPOINTER_REG_18__SCAN_IN, P2_PHYADDRPOINTER_REG_19__SCAN_IN, P2_PHYADDRPOINTER_REG_20__SCAN_IN, P2_PHYADDRPOINTER_REG_21__SCAN_IN, P2_PHYADDRPOINTER_REG_22__SCAN_IN, P2_PHYADDRPOINTER_REG_23__SCAN_IN, P2_PHYADDRPOINTER_REG_24__SCAN_IN, P2_PHYADDRPOINTER_REG_25__SCAN_IN, P2_PHYADDRPOINTER_REG_26__SCAN_IN, P2_PHYADDRPOINTER_REG_27__SCAN_IN, P2_PHYADDRPOINTER_REG_28__SCAN_IN, P2_PHYADDRPOINTER_REG_29__SCAN_IN, P2_PHYADDRPOINTER_REG_30__SCAN_IN, P2_PHYADDRPOINTER_REG_31__SCAN_IN, P2_LWORD_REG_15__SCAN_IN, P2_LWORD_REG_14__SCAN_IN, P2_LWORD_REG_13__SCAN_IN, P2_LWORD_REG_12__SCAN_IN, P2_LWORD_REG_11__SCAN_IN, P2_LWORD_REG_10__SCAN_IN, P2_LWORD_REG_9__SCAN_IN, P2_LWORD_REG_8__SCAN_IN, P2_LWORD_REG_7__SCAN_IN, P2_LWORD_REG_6__SCAN_IN, P2_LWORD_REG_5__SCAN_IN, P2_LWORD_REG_4__SCAN_IN, P2_LWORD_REG_3__SCAN_IN, P2_LWORD_REG_2__SCAN_IN, P2_LWORD_REG_1__SCAN_IN, P2_LWORD_REG_0__SCAN_IN, P2_UWORD_REG_14__SCAN_IN, P2_UWORD_REG_13__SCAN_IN, P2_UWORD_REG_12__SCAN_IN, P2_UWORD_REG_11__SCAN_IN, P2_UWORD_REG_10__SCAN_IN, P2_UWORD_REG_9__SCAN_IN, P2_UWORD_REG_8__SCAN_IN, P2_UWORD_REG_7__SCAN_IN, P2_UWORD_REG_6__SCAN_IN, P2_UWORD_REG_5__SCAN_IN, P2_UWORD_REG_4__SCAN_IN, P2_UWORD_REG_3__SCAN_IN, P2_UWORD_REG_2__SCAN_IN, P2_UWORD_REG_1__SCAN_IN, P2_UWORD_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN, P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN, P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN, P2_DATAO_REG_5__SCAN_IN, P2_DATAO_REG_6__SCAN_IN, P2_DATAO_REG_7__SCAN_IN, P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_9__SCAN_IN, P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_11__SCAN_IN, P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_13__SCAN_IN, P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_15__SCAN_IN, P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_17__SCAN_IN, P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_19__SCAN_IN, P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_21__SCAN_IN, P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_23__SCAN_IN, P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_25__SCAN_IN, P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_27__SCAN_IN, P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_29__SCAN_IN, P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_31__SCAN_IN, P2_EAX_REG_0__SCAN_IN, P2_EAX_REG_1__SCAN_IN, P2_EAX_REG_2__SCAN_IN, P2_EAX_REG_3__SCAN_IN, P2_EAX_REG_4__SCAN_IN, P2_EAX_REG_5__SCAN_IN, P2_EAX_REG_6__SCAN_IN, P2_EAX_REG_7__SCAN_IN, P2_EAX_REG_8__SCAN_IN, P2_EAX_REG_9__SCAN_IN, P2_EAX_REG_10__SCAN_IN, P2_EAX_REG_11__SCAN_IN, P2_EAX_REG_12__SCAN_IN, P2_EAX_REG_13__SCAN_IN, P2_EAX_REG_14__SCAN_IN, P2_EAX_REG_15__SCAN_IN, P2_EAX_REG_16__SCAN_IN, P2_EAX_REG_17__SCAN_IN, P2_EAX_REG_18__SCAN_IN, P2_EAX_REG_19__SCAN_IN, P2_EAX_REG_20__SCAN_IN, P2_EAX_REG_21__SCAN_IN, P2_EAX_REG_22__SCAN_IN, P2_EAX_REG_23__SCAN_IN, P2_EAX_REG_24__SCAN_IN, P2_EAX_REG_25__SCAN_IN, P2_EAX_REG_26__SCAN_IN, P2_EAX_REG_27__SCAN_IN, P2_EAX_REG_28__SCAN_IN, P2_EAX_REG_29__SCAN_IN, P2_EAX_REG_30__SCAN_IN, P2_EAX_REG_31__SCAN_IN, P2_EBX_REG_0__SCAN_IN, P2_EBX_REG_1__SCAN_IN, P2_EBX_REG_2__SCAN_IN, P2_EBX_REG_3__SCAN_IN, P2_EBX_REG_4__SCAN_IN, P2_EBX_REG_5__SCAN_IN, P2_EBX_REG_6__SCAN_IN, P2_EBX_REG_7__SCAN_IN, P2_EBX_REG_8__SCAN_IN, P2_EBX_REG_9__SCAN_IN, P2_EBX_REG_10__SCAN_IN, P2_EBX_REG_11__SCAN_IN, P2_EBX_REG_12__SCAN_IN, P2_EBX_REG_13__SCAN_IN, P2_EBX_REG_14__SCAN_IN, P2_EBX_REG_15__SCAN_IN, P2_EBX_REG_16__SCAN_IN, P2_EBX_REG_17__SCAN_IN, P2_EBX_REG_18__SCAN_IN, P2_EBX_REG_19__SCAN_IN, P2_EBX_REG_20__SCAN_IN, P2_EBX_REG_21__SCAN_IN, P2_EBX_REG_22__SCAN_IN, P2_EBX_REG_23__SCAN_IN, P2_EBX_REG_24__SCAN_IN, P2_EBX_REG_25__SCAN_IN, P2_EBX_REG_26__SCAN_IN, P2_EBX_REG_27__SCAN_IN, P2_EBX_REG_28__SCAN_IN, P2_EBX_REG_29__SCAN_IN, P2_EBX_REG_30__SCAN_IN, P2_EBX_REG_31__SCAN_IN, P2_REIP_REG_0__SCAN_IN, P2_REIP_REG_1__SCAN_IN, P2_REIP_REG_2__SCAN_IN, P2_REIP_REG_3__SCAN_IN, P2_REIP_REG_4__SCAN_IN, P2_REIP_REG_5__SCAN_IN, P2_REIP_REG_6__SCAN_IN, P2_REIP_REG_7__SCAN_IN, P2_REIP_REG_8__SCAN_IN, P2_REIP_REG_9__SCAN_IN, P2_REIP_REG_10__SCAN_IN, P2_REIP_REG_11__SCAN_IN, P2_REIP_REG_12__SCAN_IN, P2_REIP_REG_13__SCAN_IN, P2_REIP_REG_14__SCAN_IN, P2_REIP_REG_15__SCAN_IN, P2_REIP_REG_16__SCAN_IN, P2_REIP_REG_17__SCAN_IN, P2_REIP_REG_18__SCAN_IN, P2_REIP_REG_19__SCAN_IN, P2_REIP_REG_20__SCAN_IN, P2_REIP_REG_21__SCAN_IN, P2_REIP_REG_22__SCAN_IN, P2_REIP_REG_23__SCAN_IN, P2_REIP_REG_24__SCAN_IN, P2_REIP_REG_25__SCAN_IN, P2_REIP_REG_26__SCAN_IN, P2_REIP_REG_27__SCAN_IN, P2_REIP_REG_28__SCAN_IN, P2_REIP_REG_29__SCAN_IN, P2_REIP_REG_30__SCAN_IN, P2_REIP_REG_31__SCAN_IN, P2_BYTEENABLE_REG_3__SCAN_IN, P2_BYTEENABLE_REG_2__SCAN_IN, P2_BYTEENABLE_REG_1__SCAN_IN, P2_BYTEENABLE_REG_0__SCAN_IN, P2_W_R_N_REG_SCAN_IN, P2_FLUSH_REG_SCAN_IN, P2_MORE_REG_SCAN_IN, P2_STATEBS16_REG_SCAN_IN, P2_REQUESTPENDING_REG_SCAN_IN, P2_D_C_N_REG_SCAN_IN, P2_M_IO_N_REG_SCAN_IN, P2_CODEFETCH_REG_SCAN_IN, P2_ADS_N_REG_SCAN_IN, P2_READREQUEST_REG_SCAN_IN, P2_MEMORYFETCH_REG_SCAN_IN, P1_BE_N_REG_3__SCAN_IN, P1_BE_N_REG_2__SCAN_IN, P1_BE_N_REG_1__SCAN_IN, P1_BE_N_REG_0__SCAN_IN, P1_ADDRESS_REG_29__SCAN_IN, P1_ADDRESS_REG_28__SCAN_IN, P1_ADDRESS_REG_27__SCAN_IN, P1_ADDRESS_REG_26__SCAN_IN, P1_ADDRESS_REG_25__SCAN_IN, P1_ADDRESS_REG_24__SCAN_IN, P1_ADDRESS_REG_23__SCAN_IN, P1_ADDRESS_REG_22__SCAN_IN, P1_ADDRESS_REG_21__SCAN_IN, P1_ADDRESS_REG_20__SCAN_IN, P1_ADDRESS_REG_19__SCAN_IN, P1_ADDRESS_REG_18__SCAN_IN, P1_ADDRESS_REG_17__SCAN_IN, P1_ADDRESS_REG_16__SCAN_IN, P1_ADDRESS_REG_15__SCAN_IN, P1_ADDRESS_REG_14__SCAN_IN, P1_ADDRESS_REG_13__SCAN_IN, P1_ADDRESS_REG_12__SCAN_IN, P1_ADDRESS_REG_11__SCAN_IN, P1_ADDRESS_REG_10__SCAN_IN, P1_ADDRESS_REG_9__SCAN_IN, P1_ADDRESS_REG_8__SCAN_IN, P1_ADDRESS_REG_7__SCAN_IN, P1_ADDRESS_REG_6__SCAN_IN, P1_ADDRESS_REG_5__SCAN_IN, P1_ADDRESS_REG_4__SCAN_IN, P1_ADDRESS_REG_3__SCAN_IN, P1_ADDRESS_REG_2__SCAN_IN, P1_ADDRESS_REG_1__SCAN_IN, P1_ADDRESS_REG_0__SCAN_IN, P1_STATE_REG_2__SCAN_IN, P1_STATE_REG_1__SCAN_IN, P1_STATE_REG_0__SCAN_IN, P1_DATAWIDTH_REG_0__SCAN_IN, P1_DATAWIDTH_REG_1__SCAN_IN, P1_DATAWIDTH_REG_2__SCAN_IN, P1_DATAWIDTH_REG_3__SCAN_IN, P1_DATAWIDTH_REG_4__SCAN_IN, P1_DATAWIDTH_REG_5__SCAN_IN, P1_DATAWIDTH_REG_6__SCAN_IN, P1_DATAWIDTH_REG_7__SCAN_IN, P1_DATAWIDTH_REG_8__SCAN_IN, P1_DATAWIDTH_REG_9__SCAN_IN, P1_DATAWIDTH_REG_10__SCAN_IN, P1_DATAWIDTH_REG_11__SCAN_IN, P1_DATAWIDTH_REG_12__SCAN_IN, P1_DATAWIDTH_REG_13__SCAN_IN, P1_DATAWIDTH_REG_14__SCAN_IN, P1_DATAWIDTH_REG_15__SCAN_IN, P1_DATAWIDTH_REG_16__SCAN_IN, P1_DATAWIDTH_REG_17__SCAN_IN, P1_DATAWIDTH_REG_18__SCAN_IN, P1_DATAWIDTH_REG_19__SCAN_IN, P1_DATAWIDTH_REG_20__SCAN_IN, P1_DATAWIDTH_REG_21__SCAN_IN, P1_DATAWIDTH_REG_22__SCAN_IN, P1_DATAWIDTH_REG_23__SCAN_IN, P1_DATAWIDTH_REG_24__SCAN_IN, P1_DATAWIDTH_REG_25__SCAN_IN, P1_DATAWIDTH_REG_26__SCAN_IN, P1_DATAWIDTH_REG_27__SCAN_IN, P1_DATAWIDTH_REG_28__SCAN_IN, P1_DATAWIDTH_REG_29__SCAN_IN, P1_DATAWIDTH_REG_30__SCAN_IN, P1_DATAWIDTH_REG_31__SCAN_IN, P1_STATE2_REG_3__SCAN_IN, P1_STATE2_REG_2__SCAN_IN, P1_STATE2_REG_1__SCAN_IN, P1_STATE2_REG_0__SCAN_IN, P1_INSTQUEUE_REG_15__7__SCAN_IN, P1_INSTQUEUE_REG_15__6__SCAN_IN, P1_INSTQUEUE_REG_15__5__SCAN_IN, P1_INSTQUEUE_REG_15__4__SCAN_IN, P1_INSTQUEUE_REG_15__3__SCAN_IN, P1_INSTQUEUE_REG_15__2__SCAN_IN, P1_INSTQUEUE_REG_15__1__SCAN_IN, P1_INSTQUEUE_REG_15__0__SCAN_IN, P1_INSTQUEUE_REG_14__7__SCAN_IN, P1_INSTQUEUE_REG_14__6__SCAN_IN, P1_INSTQUEUE_REG_14__5__SCAN_IN, P1_INSTQUEUE_REG_14__4__SCAN_IN, P1_INSTQUEUE_REG_14__3__SCAN_IN, P1_INSTQUEUE_REG_14__2__SCAN_IN, P1_INSTQUEUE_REG_14__1__SCAN_IN, P1_INSTQUEUE_REG_14__0__SCAN_IN, P1_INSTQUEUE_REG_13__7__SCAN_IN, P1_INSTQUEUE_REG_13__6__SCAN_IN, P1_INSTQUEUE_REG_13__5__SCAN_IN, P1_INSTQUEUE_REG_13__4__SCAN_IN, P1_INSTQUEUE_REG_13__3__SCAN_IN, P1_INSTQUEUE_REG_13__2__SCAN_IN, P1_INSTQUEUE_REG_13__1__SCAN_IN, P1_INSTQUEUE_REG_13__0__SCAN_IN, P1_INSTQUEUE_REG_12__7__SCAN_IN, P1_INSTQUEUE_REG_12__6__SCAN_IN, P1_INSTQUEUE_REG_12__5__SCAN_IN, P1_INSTQUEUE_REG_12__4__SCAN_IN, P1_INSTQUEUE_REG_12__3__SCAN_IN, P1_INSTQUEUE_REG_12__2__SCAN_IN, P1_INSTQUEUE_REG_12__1__SCAN_IN, P1_INSTQUEUE_REG_12__0__SCAN_IN, P1_INSTQUEUE_REG_11__7__SCAN_IN, P1_INSTQUEUE_REG_11__6__SCAN_IN, P1_INSTQUEUE_REG_11__5__SCAN_IN, P1_INSTQUEUE_REG_11__4__SCAN_IN, P1_INSTQUEUE_REG_11__3__SCAN_IN, P1_INSTQUEUE_REG_11__2__SCAN_IN, P1_INSTQUEUE_REG_11__1__SCAN_IN, P1_INSTQUEUE_REG_11__0__SCAN_IN, P1_INSTQUEUE_REG_10__7__SCAN_IN, P1_INSTQUEUE_REG_10__6__SCAN_IN, P1_INSTQUEUE_REG_10__5__SCAN_IN, P1_INSTQUEUE_REG_10__4__SCAN_IN, P1_INSTQUEUE_REG_10__3__SCAN_IN, P1_INSTQUEUE_REG_10__2__SCAN_IN, P1_INSTQUEUE_REG_10__1__SCAN_IN, P1_INSTQUEUE_REG_10__0__SCAN_IN, P1_INSTQUEUE_REG_9__7__SCAN_IN, P1_INSTQUEUE_REG_9__6__SCAN_IN, P1_INSTQUEUE_REG_9__5__SCAN_IN, P1_INSTQUEUE_REG_9__4__SCAN_IN, P1_INSTQUEUE_REG_9__3__SCAN_IN, P1_INSTQUEUE_REG_9__2__SCAN_IN, P1_INSTQUEUE_REG_9__1__SCAN_IN, P1_INSTQUEUE_REG_9__0__SCAN_IN, P1_INSTQUEUE_REG_8__7__SCAN_IN, P1_INSTQUEUE_REG_8__6__SCAN_IN, P1_INSTQUEUE_REG_8__5__SCAN_IN, P1_INSTQUEUE_REG_8__4__SCAN_IN, P1_INSTQUEUE_REG_8__3__SCAN_IN, P1_INSTQUEUE_REG_8__2__SCAN_IN, P1_INSTQUEUE_REG_8__1__SCAN_IN, P1_INSTQUEUE_REG_8__0__SCAN_IN, P1_INSTQUEUE_REG_7__7__SCAN_IN, P1_INSTQUEUE_REG_7__6__SCAN_IN, P1_INSTQUEUE_REG_7__5__SCAN_IN, P1_INSTQUEUE_REG_7__4__SCAN_IN, P1_INSTQUEUE_REG_7__3__SCAN_IN, P1_INSTQUEUE_REG_7__2__SCAN_IN, P1_INSTQUEUE_REG_7__1__SCAN_IN, P1_INSTQUEUE_REG_7__0__SCAN_IN, P1_INSTQUEUE_REG_6__7__SCAN_IN, P1_INSTQUEUE_REG_6__6__SCAN_IN, P1_INSTQUEUE_REG_6__5__SCAN_IN, P1_INSTQUEUE_REG_6__4__SCAN_IN, P1_INSTQUEUE_REG_6__3__SCAN_IN, P1_INSTQUEUE_REG_6__2__SCAN_IN, P1_INSTQUEUE_REG_6__1__SCAN_IN, P1_INSTQUEUE_REG_6__0__SCAN_IN, P1_INSTQUEUE_REG_5__7__SCAN_IN, P1_INSTQUEUE_REG_5__6__SCAN_IN, P1_INSTQUEUE_REG_5__5__SCAN_IN, P1_INSTQUEUE_REG_5__4__SCAN_IN, P1_INSTQUEUE_REG_5__3__SCAN_IN, P1_INSTQUEUE_REG_5__2__SCAN_IN, P1_INSTQUEUE_REG_5__1__SCAN_IN, P1_INSTQUEUE_REG_5__0__SCAN_IN, P1_INSTQUEUE_REG_4__7__SCAN_IN, P1_INSTQUEUE_REG_4__6__SCAN_IN, P1_INSTQUEUE_REG_4__5__SCAN_IN, P1_INSTQUEUE_REG_4__4__SCAN_IN, P1_INSTQUEUE_REG_4__3__SCAN_IN, P1_INSTQUEUE_REG_4__2__SCAN_IN, P1_INSTQUEUE_REG_4__1__SCAN_IN, keyinput0, keyinput1, keyinput2, keyinput3, keyinput4, keyinput5, keyinput6, keyinput7, keyinput8, keyinput9, keyinput10, keyinput11, keyinput12, keyinput13, keyinput14, keyinput15, keyinput16, keyinput17, keyinput18, keyinput19, keyinput20, keyinput21, keyinput22, keyinput23, keyinput24, keyinput25, keyinput26, keyinput27, keyinput28, keyinput29, keyinput30, keyinput31, keyinput32, keyinput33, keyinput34, keyinput35, keyinput36, keyinput37, keyinput38, keyinput39, keyinput40, keyinput41, keyinput42, keyinput43, keyinput44, keyinput45, keyinput46, keyinput47, keyinput48, keyinput49, keyinput50, keyinput51, keyinput52, keyinput53, keyinput54, keyinput55, keyinput56, keyinput57, keyinput58, keyinput59, keyinput60, keyinput61, keyinput62, keyinput63;
  output P3_DATAO_REG_31__SCAN_IN, P3_DATAO_REG_30__SCAN_IN, P3_DATAO_REG_29__SCAN_IN, P3_DATAO_REG_28__SCAN_IN, P3_DATAO_REG_27__SCAN_IN, P3_DATAO_REG_26__SCAN_IN, P3_DATAO_REG_25__SCAN_IN, P3_DATAO_REG_24__SCAN_IN, P3_DATAO_REG_23__SCAN_IN, P3_DATAO_REG_22__SCAN_IN, P3_DATAO_REG_21__SCAN_IN, P3_DATAO_REG_20__SCAN_IN, P3_DATAO_REG_19__SCAN_IN, P3_DATAO_REG_18__SCAN_IN, P3_DATAO_REG_17__SCAN_IN, P3_DATAO_REG_16__SCAN_IN, P3_DATAO_REG_15__SCAN_IN, P3_DATAO_REG_14__SCAN_IN, P3_DATAO_REG_13__SCAN_IN, P3_DATAO_REG_12__SCAN_IN, P3_DATAO_REG_11__SCAN_IN, P3_DATAO_REG_10__SCAN_IN, P3_DATAO_REG_9__SCAN_IN, P3_DATAO_REG_8__SCAN_IN, P3_DATAO_REG_7__SCAN_IN, P3_DATAO_REG_6__SCAN_IN, P3_DATAO_REG_5__SCAN_IN, P3_DATAO_REG_4__SCAN_IN, P3_DATAO_REG_3__SCAN_IN, P3_DATAO_REG_2__SCAN_IN, P3_DATAO_REG_1__SCAN_IN, P3_DATAO_REG_0__SCAN_IN, P1_ADDRESS_REG_29__SCAN_IN, P1_ADDRESS_REG_28__SCAN_IN, P1_ADDRESS_REG_27__SCAN_IN, P1_ADDRESS_REG_26__SCAN_IN, P1_ADDRESS_REG_25__SCAN_IN, P1_ADDRESS_REG_24__SCAN_IN, P1_ADDRESS_REG_23__SCAN_IN, P1_ADDRESS_REG_22__SCAN_IN, P1_ADDRESS_REG_21__SCAN_IN, P1_ADDRESS_REG_20__SCAN_IN, P1_ADDRESS_REG_19__SCAN_IN, P1_ADDRESS_REG_18__SCAN_IN, P1_ADDRESS_REG_17__SCAN_IN, P1_ADDRESS_REG_16__SCAN_IN, P1_ADDRESS_REG_15__SCAN_IN, P1_ADDRESS_REG_14__SCAN_IN, P1_ADDRESS_REG_13__SCAN_IN, P1_ADDRESS_REG_12__SCAN_IN, P1_ADDRESS_REG_11__SCAN_IN, P1_ADDRESS_REG_10__SCAN_IN, P1_ADDRESS_REG_9__SCAN_IN, P1_ADDRESS_REG_8__SCAN_IN, P1_ADDRESS_REG_7__SCAN_IN, P1_ADDRESS_REG_6__SCAN_IN, P1_ADDRESS_REG_5__SCAN_IN, P1_ADDRESS_REG_4__SCAN_IN, P1_ADDRESS_REG_3__SCAN_IN, P1_ADDRESS_REG_2__SCAN_IN, P1_ADDRESS_REG_1__SCAN_IN, P1_ADDRESS_REG_0__SCAN_IN, U355, U356, U357, U358, U359, U360, U361, U362, U363, U364, U366, U367, U368, U369, U370, U371, U372, U373, U374, U375, U347, U348, U349, U350, U351, U352, U353, U354, U365, U376, P3_W_R_N_REG_SCAN_IN, P3_D_C_N_REG_SCAN_IN, P3_M_IO_N_REG_SCAN_IN, P1_ADS_N_REG_SCAN_IN, P3_ADS_N_REG_SCAN_IN, U247, U246, U245, U244, U243, U242, U241, U240, U239, U238, U237, U236, U235, U234, U233, U232, U231, U230, U229, U228, U227, U226, U225, U224, U223, U222, U221, U220, U219, U218, U217, U216, U251, U252, U253, U254, U255, U256, U257, U258, U259, U260, U261, U262, U263, U264, U265, U266, U267, U268, U269, U270, U271, U272, U273, U274, U275, U276, U277, U278, U279, U280, U281, U282, U212, U215, U213, U214, P3_U3274, P3_U3275, P3_U3276, P3_U3277, P3_U3061, P3_U3060, P3_U3059, P3_U3058, P3_U3057, P3_U3056, P3_U3055, P3_U3054, P3_U3053, P3_U3052, P3_U3051, P3_U3050, P3_U3049, P3_U3048, P3_U3047, P3_U3046, P3_U3045, P3_U3044, P3_U3043, P3_U3042, P3_U3041, P3_U3040, P3_U3039, P3_U3038, P3_U3037, P3_U3036, P3_U3035, P3_U3034, P3_U3033, P3_U3032, P3_U3031, P3_U3030, P3_U3029, P3_U3280, P3_U3281, P3_U3028, P3_U3027, P3_U3026, P3_U3025, P3_U3024, P3_U3023, P3_U3022, P3_U3021, P3_U3020, P3_U3019, P3_U3018, P3_U3017, P3_U3016, P3_U3015, P3_U3014, P3_U3013, P3_U3012, P3_U3011, P3_U3010, P3_U3009, P3_U3008, P3_U3007, P3_U3006, P3_U3005, P3_U3004, P3_U3003, P3_U3002, P3_U3001, P3_U3000, P3_U2999, P3_U3282, P3_U2998, P3_U2997, P3_U2996, P3_U2995, P3_U2994, P3_U2993, P3_U2992, P3_U2991, P3_U2990, P3_U2989, P3_U2988, P3_U2987, P3_U2986, P3_U2985, P3_U2984, P3_U2983, P3_U2982, P3_U2981, P3_U2980, P3_U2979, P3_U2978, P3_U2977, P3_U2976, P3_U2975, P3_U2974, P3_U2973, P3_U2972, P3_U2971, P3_U2970, P3_U2969, P3_U2968, P3_U2967, P3_U2966, P3_U2965, P3_U2964, P3_U2963, P3_U2962, P3_U2961, P3_U2960, P3_U2959, P3_U2958, P3_U2957, P3_U2956, P3_U2955, P3_U2954, P3_U2953, P3_U2952, P3_U2951, P3_U2950, P3_U2949, P3_U2948, P3_U2947, P3_U2946, P3_U2945, P3_U2944, P3_U2943, P3_U2942, P3_U2941, P3_U2940, P3_U2939, P3_U2938, P3_U2937, P3_U2936, P3_U2935, P3_U2934, P3_U2933, P3_U2932, P3_U2931, P3_U2930, P3_U2929, P3_U2928, P3_U2927, P3_U2926, P3_U2925, P3_U2924, P3_U2923, P3_U2922, P3_U2921, P3_U2920, P3_U2919, P3_U2918, P3_U2917, P3_U2916, P3_U2915, P3_U2914, P3_U2913, P3_U2912, P3_U2911, P3_U2910, P3_U2909, P3_U2908, P3_U2907, P3_U2906, P3_U2905, P3_U2904, P3_U2903, P3_U2902, P3_U2901, P3_U2900, P3_U2899, P3_U2898, P3_U2897, P3_U2896, P3_U2895, P3_U2894, P3_U2893, P3_U2892, P3_U2891, P3_U2890, P3_U2889, P3_U2888, P3_U2887, P3_U2886, P3_U2885, P3_U2884, P3_U2883, P3_U2882, P3_U2881, P3_U2880, P3_U2879, P3_U2878, P3_U2877, P3_U2876, P3_U2875, P3_U2874, P3_U2873, P3_U2872, P3_U2871, P3_U2870, P3_U2869, P3_U2868, P3_U3284, P3_U3285, P3_U3288, P3_U3289, P3_U3290, P3_U2867, P3_U2866, P3_U2865, P3_U2864, P3_U2863, P3_U2862, P3_U2861, P3_U2860, P3_U2859, P3_U2858, P3_U2857, P3_U2856, P3_U2855, P3_U2854, P3_U2853, P3_U2852, P3_U2851, P3_U2850, P3_U2849, P3_U2848, P3_U2847, P3_U2846, P3_U2845, P3_U2844, P3_U2843, P3_U2842, P3_U2841, P3_U2840, P3_U2839, P3_U2838, P3_U2837, P3_U2836, P3_U2835, P3_U2834, P3_U2833, P3_U2832, P3_U2831, P3_U2830, P3_U2829, P3_U2828, P3_U2827, P3_U2826, P3_U2825, P3_U2824, P3_U2823, P3_U2822, P3_U2821, P3_U2820, P3_U2819, P3_U2818, P3_U2817, P3_U2816, P3_U2815, P3_U2814, P3_U2813, P3_U2812, P3_U2811, P3_U2810, P3_U2809, P3_U2808, P3_U2807, P3_U2806, P3_U2805, P3_U2804, P3_U2803, P3_U2802, P3_U2801, P3_U2800, P3_U2799, P3_U2798, P3_U2797, P3_U2796, P3_U2795, P3_U2794, P3_U2793, P3_U2792, P3_U2791, P3_U2790, P3_U2789, P3_U2788, P3_U2787, P3_U2786, P3_U2785, P3_U2784, P3_U2783, P3_U2782, P3_U2781, P3_U2780, P3_U2779, P3_U2778, P3_U2777, P3_U2776, P3_U2775, P3_U2774, P3_U2773, P3_U2772, P3_U2771, P3_U2770, P3_U2769, P3_U2768, P3_U2767, P3_U2766, P3_U2765, P3_U2764, P3_U2763, P3_U2762, P3_U2761, P3_U2760, P3_U2759, P3_U2758, P3_U2757, P3_U2756, P3_U2755, P3_U2754, P3_U2753, P3_U2752, P3_U2751, P3_U2750, P3_U2749, P3_U2748, P3_U2747, P3_U2746, P3_U2745, P3_U2744, P3_U2743, P3_U2742, P3_U2741, P3_U2740, P3_U2739, P3_U2738, P3_U2737, P3_U2736, P3_U2735, P3_U2734, P3_U2733, P3_U2732, P3_U2731, P3_U2730, P3_U2729, P3_U2728, P3_U2727, P3_U2726, P3_U2725, P3_U2724, P3_U2723, P3_U2722, P3_U2721, P3_U2720, P3_U2719, P3_U2718, P3_U2717, P3_U2716, P3_U2715, P3_U2714, P3_U2713, P3_U2712, P3_U2711, P3_U2710, P3_U2709, P3_U2708, P3_U2707, P3_U2706, P3_U2705, P3_U2704, P3_U2703, P3_U2702, P3_U2701, P3_U2700, P3_U2699, P3_U2698, P3_U2697, P3_U2696, P3_U2695, P3_U2694, P3_U2693, P3_U2692, P3_U2691, P3_U2690, P3_U2689, P3_U2688, P3_U2687, P3_U2686, P3_U2685, P3_U2684, P3_U2683, P3_U2682, P3_U2681, P3_U2680, P3_U2679, P3_U2678, P3_U2677, P3_U2676, P3_U2675, P3_U2674, P3_U2673, P3_U2672, P3_U2671, P3_U2670, P3_U2669, P3_U2668, P3_U2667, P3_U2666, P3_U2665, P3_U2664, P3_U2663, P3_U2662, P3_U2661, P3_U2660, P3_U2659, P3_U2658, P3_U2657, P3_U2656, P3_U2655, P3_U2654, P3_U2653, P3_U2652, P3_U2651, P3_U2650, P3_U2649, P3_U2648, P3_U2647, P3_U2646, P3_U2645, P3_U2644, P3_U2643, P3_U2642, P3_U2641, P3_U2640, P3_U2639, P3_U3292, P3_U2638, P3_U3293, P3_U3294, P3_U2637, P3_U3295, P3_U2636, P3_U3296, P3_U2635, P3_U3297, P3_U2634, P3_U2633, P3_U3298, P3_U3299, P2_U3585, P2_U3586, P2_U3587, P2_U3588, P2_U3241, P2_U3240, P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234, P2_U3233, P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227, P2_U3226, P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220, P2_U3219, P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3214, P2_U3213, P2_U3212, P2_U3211, P2_U3210, P2_U3209, P2_U3591, P2_U3592, P2_U3208, P2_U3207, P2_U3206, P2_U3205, P2_U3204, P2_U3203, P2_U3202, P2_U3201, P2_U3200, P2_U3199, P2_U3198, P2_U3197, P2_U3196, P2_U3195, P2_U3194, P2_U3193, P2_U3192, P2_U3191, P2_U3190, P2_U3189, P2_U3188, P2_U3187, P2_U3186, P2_U3185, P2_U3184, P2_U3183, P2_U3182, P2_U3181, P2_U3180, P2_U3179, P2_U3593, P2_U3178, P2_U3177, P2_U3176, P2_U3175, P2_U3174, P2_U3173, P2_U3172, P2_U3171, P2_U3170, P2_U3169, P2_U3168, P2_U3167, P2_U3166, P2_U3165, P2_U3164, P2_U3163, P2_U3162, P2_U3161, P2_U3160, P2_U3159, P2_U3158, P2_U3157, P2_U3156, P2_U3155, P2_U3154, P2_U3153, P2_U3152, P2_U3151, P2_U3150, P2_U3149, P2_U3148, P2_U3147, P2_U3146, P2_U3145, P2_U3144, P2_U3143, P2_U3142, P2_U3141, P2_U3140, P2_U3139, P2_U3138, P2_U3137, P2_U3136, P2_U3135, P2_U3134, P2_U3133, P2_U3132, P2_U3131, P2_U3130, P2_U3129, P2_U3128, P2_U3127, P2_U3126, P2_U3125, P2_U3124, P2_U3123, P2_U3122, P2_U3121, P2_U3120, P2_U3119, P2_U3118, P2_U3117, P2_U3116, P2_U3115, P2_U3114, P2_U3113, P2_U3112, P2_U3111, P2_U3110, P2_U3109, P2_U3108, P2_U3107, P2_U3106, P2_U3105, P2_U3104, P2_U3103, P2_U3102, P2_U3101, P2_U3100, P2_U3099, P2_U3098, P2_U3097, P2_U3096, P2_U3095, P2_U3094, P2_U3093, P2_U3092, P2_U3091, P2_U3090, P2_U3089, P2_U3088, P2_U3087, P2_U3086, P2_U3085, P2_U3084, P2_U3083, P2_U3082, P2_U3081, P2_U3080, P2_U3079, P2_U3078, P2_U3077, P2_U3076, P2_U3075, P2_U3074, P2_U3073, P2_U3072, P2_U3071, P2_U3070, P2_U3069, P2_U3068, P2_U3067, P2_U3066, P2_U3065, P2_U3064, P2_U3063, P2_U3062, P2_U3061, P2_U3060, P2_U3059, P2_U3058, P2_U3057, P2_U3056, P2_U3055, P2_U3054, P2_U3053, P2_U3052, P2_U3051, P2_U3050, P2_U3049, P2_U3048, P2_U3595, P2_U3596, P2_U3599, P2_U3600, P2_U3601, P2_U3047, P2_U3602, P2_U3603, P2_U3604, P2_U3605, P2_U3046, P2_U3045, P2_U3044, P2_U3043, P2_U3042, P2_U3041, P2_U3040, P2_U3039, P2_U3038, P2_U3037, P2_U3036, P2_U3035, P2_U3034, P2_U3033, P2_U3032, P2_U3031, P2_U3030, P2_U3029, P2_U3028, P2_U3027, P2_U3026, P2_U3025, P2_U3024, P2_U3023, P2_U3022, P2_U3021, P2_U3020, P2_U3019, P2_U3018, P2_U3017, P2_U3016, P2_U3015, P2_U3014, P2_U3013, P2_U3012, P2_U3011, P2_U3010, P2_U3009, P2_U3008, P2_U3007, P2_U3006, P2_U3005, P2_U3004, P2_U3003, P2_U3002, P2_U3001, P2_U3000, P2_U2999, P2_U2998, P2_U2997, P2_U2996, P2_U2995, P2_U2994, P2_U2993, P2_U2992, P2_U2991, P2_U2990, P2_U2989, P2_U2988, P2_U2987, P2_U2986, P2_U2985, P2_U2984, P2_U2983, P2_U2982, P2_U2981, P2_U2980, P2_U2979, P2_U2978, P2_U2977, P2_U2976, P2_U2975, P2_U2974, P2_U2973, P2_U2972, P2_U2971, P2_U2970, P2_U2969, P2_U2968, P2_U2967, P2_U2966, P2_U2965, P2_U2964, P2_U2963, P2_U2962, P2_U2961, P2_U2960, P2_U2959, P2_U2958, P2_U2957, P2_U2956, P2_U2955, P2_U2954, P2_U2953, P2_U2952, P2_U2951, P2_U2950, P2_U2949, P2_U2948, P2_U2947, P2_U2946, P2_U2945, P2_U2944, P2_U2943, P2_U2942, P2_U2941, P2_U2940, P2_U2939, P2_U2938, P2_U2937, P2_U2936, P2_U2935, P2_U2934, P2_U2933, P2_U2932, P2_U2931, P2_U2930, P2_U2929, P2_U2928, P2_U2927, P2_U2926, P2_U2925, P2_U2924, P2_U2923, P2_U2922, P2_U2921, P2_U2920, P2_U2919, P2_U2918, P2_U2917, P2_U2916, P2_U2915, P2_U2914, P2_U2913, P2_U2912, P2_U2911, P2_U2910, P2_U2909, P2_U2908, P2_U2907, P2_U2906, P2_U2905, P2_U2904, P2_U2903, P2_U2902, P2_U2901, P2_U2900, P2_U2899, P2_U2898, P2_U2897, P2_U2896, P2_U2895, P2_U2894, P2_U2893, P2_U2892, P2_U2891, P2_U2890, P2_U2889, P2_U2888, P2_U2887, P2_U2886, P2_U2885, P2_U2884, P2_U2883, P2_U2882, P2_U2881, P2_U2880, P2_U2879, P2_U2878, P2_U2877, P2_U2876, P2_U2875, P2_U2874, P2_U2873, P2_U2872, P2_U2871, P2_U2870, P2_U2869, P2_U2868, P2_U2867, P2_U2866, P2_U2865, P2_U2864, P2_U2863, P2_U2862, P2_U2861, P2_U2860, P2_U2859, P2_U2858, P2_U2857, P2_U2856, P2_U2855, P2_U2854, P2_U2853, P2_U2852, P2_U2851, P2_U2850, P2_U2849, P2_U2848, P2_U2847, P2_U2846, P2_U2845, P2_U2844, P2_U2843, P2_U2842, P2_U2841, P2_U2840, P2_U2839, P2_U2838, P2_U2837, P2_U2836, P2_U2835, P2_U2834, P2_U2833, P2_U2832, P2_U2831, P2_U2830, P2_U2829, P2_U2828, P2_U2827, P2_U2826, P2_U2825, P2_U2824, P2_U2823, P2_U2822, P2_U2821, P2_U2820, P2_U3608, P2_U2819, P2_U3609, P2_U2818, P2_U3610, P2_U2817, P2_U3611, P2_U2816, P2_U2815, P2_U3612, P2_U2814, P1_U3458, P1_U3459, P1_U3460, P1_U3461, P1_U3226, P1_U3225, P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218, P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3212, P1_U3211, P1_U3210, P1_U3209, P1_U3208, P1_U3207, P1_U3206, P1_U3205, P1_U3204, P1_U3203, P1_U3202, P1_U3201, P1_U3200, P1_U3199, P1_U3198, P1_U3197, P1_U3196, P1_U3195, P1_U3194, P1_U3464, P1_U3465, P1_U3193, P1_U3192, P1_U3191, P1_U3190, P1_U3189, P1_U3188, P1_U3187, P1_U3186, P1_U3185, P1_U3184, P1_U3183, P1_U3182, P1_U3181, P1_U3180, P1_U3179, P1_U3178, P1_U3177, P1_U3176, P1_U3175, P1_U3174, P1_U3173, P1_U3172, P1_U3171, P1_U3170, P1_U3169, P1_U3168, P1_U3167, P1_U3166, P1_U3165, P1_U3164, P1_U3466, P1_U3163, P1_U3162, P1_U3161, P1_U3160, P1_U3159, P1_U3158, P1_U3157, P1_U3156, P1_U3155, P1_U3154, P1_U3153, P1_U3152, P1_U3151, P1_U3150, P1_U3149, P1_U3148, P1_U3147, P1_U3146, P1_U3145, P1_U3144, P1_U3143, P1_U3142, P1_U3141, P1_U3140, P1_U3139, P1_U3138, P1_U3137, P1_U3136, P1_U3135, P1_U3134, P1_U3133, P1_U3132, P1_U3131, P1_U3130, P1_U3129, P1_U3128, P1_U3127, P1_U3126, P1_U3125, P1_U3124, P1_U3123, P1_U3122, P1_U3121, P1_U3120, P1_U3119, P1_U3118, P1_U3117, P1_U3116, P1_U3115, P1_U3114, P1_U3113, P1_U3112, P1_U3111, P1_U3110, P1_U3109, P1_U3108, P1_U3107, P1_U3106, P1_U3105, P1_U3104, P1_U3103, P1_U3102, P1_U3101, P1_U3100, P1_U3099, P1_U3098, P1_U3097, P1_U3096, P1_U3095, P1_U3094, P1_U3093, P1_U3092, P1_U3091, P1_U3090, P1_U3089, P1_U3088, P1_U3087, P1_U3086, P1_U3085, P1_U3084, P1_U3083, P1_U3082, P1_U3081, P1_U3080, P1_U3079, P1_U3078, P1_U3077, P1_U3076, P1_U3075, P1_U3074, P1_U3073, P1_U3072, P1_U3071, P1_U3070, P1_U3069, P1_U3068, P1_U3067, P1_U3066, P1_U3065, P1_U3064, P1_U3063, P1_U3062, P1_U3061, P1_U3060, P1_U3059, P1_U3058, P1_U3057, P1_U3056, P1_U3055, P1_U3054, P1_U3053, P1_U3052, P1_U3051, P1_U3050, P1_U3049, P1_U3048, P1_U3047, P1_U3046, P1_U3045, P1_U3044, P1_U3043, P1_U3042, P1_U3041, P1_U3040, P1_U3039, P1_U3038, P1_U3037, P1_U3036, P1_U3035, P1_U3034, P1_U3033, P1_U3468, P1_U3469, P1_U3472, P1_U3473, P1_U3474, P1_U3032, P1_U3475, P1_U3476, P1_U3477, P1_U3478, P1_U3031, P1_U3030, P1_U3029, P1_U3028, P1_U3027, P1_U3026, P1_U3025, P1_U3024, P1_U3023, P1_U3022, P1_U3021, P1_U3020, P1_U3019, P1_U3018, P1_U3017, P1_U3016, P1_U3015, P1_U3014, P1_U3013, P1_U3012, P1_U3011, P1_U3010, P1_U3009, P1_U3008, P1_U3007, P1_U3006, P1_U3005, P1_U3004, P1_U3003, P1_U3002, P1_U3001, P1_U3000, P1_U2999, P1_U2998, P1_U2997, P1_U2996, P1_U2995, P1_U2994, P1_U2993, P1_U2992, P1_U2991, P1_U2990, P1_U2989, P1_U2988, P1_U2987, P1_U2986, P1_U2985, P1_U2984, P1_U2983, P1_U2982, P1_U2981, P1_U2980, P1_U2979, P1_U2978, P1_U2977, P1_U2976, P1_U2975, P1_U2974, P1_U2973, P1_U2972, P1_U2971, P1_U2970, P1_U2969, P1_U2968, P1_U2967, P1_U2966, P1_U2965, P1_U2964, P1_U2963, P1_U2962, P1_U2961, P1_U2960, P1_U2959, P1_U2958, P1_U2957, P1_U2956, P1_U2955, P1_U2954, P1_U2953, P1_U2952, P1_U2951, P1_U2950, P1_U2949, P1_U2948, P1_U2947, P1_U2946, P1_U2945, P1_U2944, P1_U2943, P1_U2942, P1_U2941, P1_U2940, P1_U2939, P1_U2938, P1_U2937, P1_U2936, P1_U2935, P1_U2934, P1_U2933, P1_U2932, P1_U2931, P1_U2930, P1_U2929, P1_U2928, P1_U2927, P1_U2926, P1_U2925, P1_U2924, P1_U2923, P1_U2922, P1_U2921, P1_U2920, P1_U2919, P1_U2918, P1_U2917, P1_U2916, P1_U2915, P1_U2914, P1_U2913, P1_U2912, P1_U2911, P1_U2910, P1_U2909, P1_U2908, P1_U2907, P1_U2906, P1_U2905, P1_U2904, P1_U2903, P1_U2902, P1_U2901, P1_U2900, P1_U2899, P1_U2898, P1_U2897, P1_U2896, P1_U2895, P1_U2894, P1_U2893, P1_U2892, P1_U2891, P1_U2890, P1_U2889, P1_U2888, P1_U2887, P1_U2886, P1_U2885, P1_U2884, P1_U2883, P1_U2882, P1_U2881, P1_U2880, P1_U2879, P1_U2878, P1_U2877, P1_U2876, P1_U2875, P1_U2874, P1_U2873, P1_U2872, P1_U2871, P1_U2870, P1_U2869, P1_U2868, P1_U2867, P1_U2866, P1_U2865, P1_U2864, P1_U2863, P1_U2862, P1_U2861, P1_U2860, P1_U2859, P1_U2858, P1_U2857, P1_U2856, P1_U2855, P1_U2854, P1_U2853, P1_U2852, P1_U2851, P1_U2850, P1_U2849, P1_U2848, P1_U2847, P1_U2846, P1_U2845, P1_U2844, P1_U2843, P1_U2842, P1_U2841, P1_U2840, P1_U2839, P1_U2838, P1_U2837, P1_U2836, P1_U2835, P1_U2834, P1_U2833, P1_U2832, P1_U2831, P1_U2830, P1_U2829, P1_U2828, P1_U2827, P1_U2826, P1_U2825, P1_U2824, P1_U2823, P1_U2822, P1_U2821, P1_U2820, P1_U2819, P1_U2818, P1_U2817, P1_U2816, P1_U2815, P1_U2814, P1_U2813, P1_U2812, P1_U2811, P1_U2810, P1_U2809, P1_U2808, P1_U3481, P1_U2807, P1_U3482, P1_U3483, P1_U2806, P1_U3484, P1_U2805, P1_U3485, P1_U2804, P1_U3486, P1_U2803, P1_U2802, P1_U3487, P1_U2801;
  wire LT_748_U6, LT_782_119_U6, LT_782_119_U7, LT_782_120_U6, LT_782_120_U7, LT_782_U6, LT_782_U7, P1_ADD_371_U10, P1_ADD_371_U11, P1_ADD_371_U12, P1_ADD_371_U13, P1_ADD_371_U14, P1_ADD_371_U15, P1_ADD_371_U16, P1_ADD_371_U17, P1_ADD_371_U18, P1_ADD_371_U19, P1_ADD_371_U20, P1_ADD_371_U21, P1_ADD_371_U22, P1_ADD_371_U23, P1_ADD_371_U24, P1_ADD_371_U25, P1_ADD_371_U26, P1_ADD_371_U27, P1_ADD_371_U28, P1_ADD_371_U29, P1_ADD_371_U30, P1_ADD_371_U31, P1_ADD_371_U32, P1_ADD_371_U33, P1_ADD_371_U34, P1_ADD_371_U35, P1_ADD_371_U36, P1_ADD_371_U37, P1_ADD_371_U38, P1_ADD_371_U39, P1_ADD_371_U4, P1_ADD_371_U40, P1_ADD_371_U41, P1_ADD_371_U42, P1_ADD_371_U43, P1_ADD_371_U44, P1_ADD_371_U5, P1_ADD_371_U6, P1_ADD_371_U7, P1_ADD_371_U8, P1_ADD_371_U9, P1_ADD_405_U10, P1_ADD_405_U100, P1_ADD_405_U101, P1_ADD_405_U102, P1_ADD_405_U103, P1_ADD_405_U104, P1_ADD_405_U105, P1_ADD_405_U106, P1_ADD_405_U107, P1_ADD_405_U108, P1_ADD_405_U109, P1_ADD_405_U11, P1_ADD_405_U110, P1_ADD_405_U111, P1_ADD_405_U112, P1_ADD_405_U113, P1_ADD_405_U114, P1_ADD_405_U115, P1_ADD_405_U116, P1_ADD_405_U117, P1_ADD_405_U118, P1_ADD_405_U119, P1_ADD_405_U12, P1_ADD_405_U120, P1_ADD_405_U121, P1_ADD_405_U122, P1_ADD_405_U123, P1_ADD_405_U124, P1_ADD_405_U125, P1_ADD_405_U126, P1_ADD_405_U127, P1_ADD_405_U128, P1_ADD_405_U129, P1_ADD_405_U13, P1_ADD_405_U130, P1_ADD_405_U131, P1_ADD_405_U132, P1_ADD_405_U133, P1_ADD_405_U134, P1_ADD_405_U135, P1_ADD_405_U136, P1_ADD_405_U137, P1_ADD_405_U138, P1_ADD_405_U139, P1_ADD_405_U14, P1_ADD_405_U140, P1_ADD_405_U141, P1_ADD_405_U142, P1_ADD_405_U143, P1_ADD_405_U144, P1_ADD_405_U145, P1_ADD_405_U146, P1_ADD_405_U147, P1_ADD_405_U148, P1_ADD_405_U149, P1_ADD_405_U15, P1_ADD_405_U150, P1_ADD_405_U151, P1_ADD_405_U152, P1_ADD_405_U153, P1_ADD_405_U154, P1_ADD_405_U155, P1_ADD_405_U156, P1_ADD_405_U157, P1_ADD_405_U158, P1_ADD_405_U159, P1_ADD_405_U16, P1_ADD_405_U160, P1_ADD_405_U161, P1_ADD_405_U162, P1_ADD_405_U163, P1_ADD_405_U164, P1_ADD_405_U165, P1_ADD_405_U166, P1_ADD_405_U167, P1_ADD_405_U168, P1_ADD_405_U169, P1_ADD_405_U17, P1_ADD_405_U170, P1_ADD_405_U171, P1_ADD_405_U172, P1_ADD_405_U173, P1_ADD_405_U174, P1_ADD_405_U175, P1_ADD_405_U176, P1_ADD_405_U177, P1_ADD_405_U178, P1_ADD_405_U179, P1_ADD_405_U18, P1_ADD_405_U180, P1_ADD_405_U181, P1_ADD_405_U182, P1_ADD_405_U183, P1_ADD_405_U184, P1_ADD_405_U185, P1_ADD_405_U186, P1_ADD_405_U19, P1_ADD_405_U20, P1_ADD_405_U21, P1_ADD_405_U22, P1_ADD_405_U23, P1_ADD_405_U24, P1_ADD_405_U25, P1_ADD_405_U26, P1_ADD_405_U27, P1_ADD_405_U28, P1_ADD_405_U29, P1_ADD_405_U30, P1_ADD_405_U31, P1_ADD_405_U32, P1_ADD_405_U33, P1_ADD_405_U34, P1_ADD_405_U35, P1_ADD_405_U36, P1_ADD_405_U37, P1_ADD_405_U38, P1_ADD_405_U39, P1_ADD_405_U4, P1_ADD_405_U40, P1_ADD_405_U41, P1_ADD_405_U42, P1_ADD_405_U43, P1_ADD_405_U44, P1_ADD_405_U45, P1_ADD_405_U46, P1_ADD_405_U47, P1_ADD_405_U48, P1_ADD_405_U49, P1_ADD_405_U5, P1_ADD_405_U50, P1_ADD_405_U51, P1_ADD_405_U52, P1_ADD_405_U53, P1_ADD_405_U54, P1_ADD_405_U55, P1_ADD_405_U56, P1_ADD_405_U57, P1_ADD_405_U58, P1_ADD_405_U59, P1_ADD_405_U6, P1_ADD_405_U60, P1_ADD_405_U61, P1_ADD_405_U62, P1_ADD_405_U63, P1_ADD_405_U64, P1_ADD_405_U65, P1_ADD_405_U66, P1_ADD_405_U67, P1_ADD_405_U68, P1_ADD_405_U69, P1_ADD_405_U7, P1_ADD_405_U70, P1_ADD_405_U71, P1_ADD_405_U72, P1_ADD_405_U73, P1_ADD_405_U74, P1_ADD_405_U75, P1_ADD_405_U76, P1_ADD_405_U77, P1_ADD_405_U78, P1_ADD_405_U79, P1_ADD_405_U8, P1_ADD_405_U80, P1_ADD_405_U81, P1_ADD_405_U82, P1_ADD_405_U83, P1_ADD_405_U84, P1_ADD_405_U85, P1_ADD_405_U86, P1_ADD_405_U87, P1_ADD_405_U88, P1_ADD_405_U89, P1_ADD_405_U9, P1_ADD_405_U90, P1_ADD_405_U91, P1_ADD_405_U92, P1_ADD_405_U93, P1_ADD_405_U94, P1_ADD_405_U95, P1_ADD_405_U96, P1_ADD_405_U97, P1_ADD_405_U98, P1_ADD_405_U99, P1_ADD_515_U10, P1_ADD_515_U100, P1_ADD_515_U101, P1_ADD_515_U102, P1_ADD_515_U103, P1_ADD_515_U104, P1_ADD_515_U105, P1_ADD_515_U106, P1_ADD_515_U107, P1_ADD_515_U108, P1_ADD_515_U109, P1_ADD_515_U11, P1_ADD_515_U110, P1_ADD_515_U111, P1_ADD_515_U112, P1_ADD_515_U113, P1_ADD_515_U114, P1_ADD_515_U115, P1_ADD_515_U116, P1_ADD_515_U117, P1_ADD_515_U118, P1_ADD_515_U119, P1_ADD_515_U12, P1_ADD_515_U120, P1_ADD_515_U121, P1_ADD_515_U122, P1_ADD_515_U123, P1_ADD_515_U124, P1_ADD_515_U125, P1_ADD_515_U126, P1_ADD_515_U127, P1_ADD_515_U128, P1_ADD_515_U129, P1_ADD_515_U13, P1_ADD_515_U130, P1_ADD_515_U131, P1_ADD_515_U132, P1_ADD_515_U133, P1_ADD_515_U134, P1_ADD_515_U135, P1_ADD_515_U136, P1_ADD_515_U137, P1_ADD_515_U138, P1_ADD_515_U139, P1_ADD_515_U14, P1_ADD_515_U140, P1_ADD_515_U141, P1_ADD_515_U142, P1_ADD_515_U143, P1_ADD_515_U144, P1_ADD_515_U145, P1_ADD_515_U146, P1_ADD_515_U147, P1_ADD_515_U148, P1_ADD_515_U149, P1_ADD_515_U15, P1_ADD_515_U150, P1_ADD_515_U151, P1_ADD_515_U152, P1_ADD_515_U153, P1_ADD_515_U154, P1_ADD_515_U155, P1_ADD_515_U156, P1_ADD_515_U157, P1_ADD_515_U158, P1_ADD_515_U159, P1_ADD_515_U16, P1_ADD_515_U160, P1_ADD_515_U161, P1_ADD_515_U162, P1_ADD_515_U163, P1_ADD_515_U164, P1_ADD_515_U165, P1_ADD_515_U166, P1_ADD_515_U167, P1_ADD_515_U168, P1_ADD_515_U169, P1_ADD_515_U17, P1_ADD_515_U170, P1_ADD_515_U171, P1_ADD_515_U172, P1_ADD_515_U173, P1_ADD_515_U174, P1_ADD_515_U175, P1_ADD_515_U176, P1_ADD_515_U177, P1_ADD_515_U178, P1_ADD_515_U179, P1_ADD_515_U18, P1_ADD_515_U180, P1_ADD_515_U181, P1_ADD_515_U182, P1_ADD_515_U19, P1_ADD_515_U20, P1_ADD_515_U21, P1_ADD_515_U22, P1_ADD_515_U23, P1_ADD_515_U24, P1_ADD_515_U25, P1_ADD_515_U26, P1_ADD_515_U27, P1_ADD_515_U28, P1_ADD_515_U29, P1_ADD_515_U30, P1_ADD_515_U31, P1_ADD_515_U32, P1_ADD_515_U33, P1_ADD_515_U34, P1_ADD_515_U35, P1_ADD_515_U36, P1_ADD_515_U37, P1_ADD_515_U38, P1_ADD_515_U39, P1_ADD_515_U4, P1_ADD_515_U40, P1_ADD_515_U41, P1_ADD_515_U42, P1_ADD_515_U43, P1_ADD_515_U44, P1_ADD_515_U45, P1_ADD_515_U46, P1_ADD_515_U47, P1_ADD_515_U48, P1_ADD_515_U49, P1_ADD_515_U5, P1_ADD_515_U50, P1_ADD_515_U51, P1_ADD_515_U52, P1_ADD_515_U53, P1_ADD_515_U54, P1_ADD_515_U55, P1_ADD_515_U56, P1_ADD_515_U57, P1_ADD_515_U58, P1_ADD_515_U59, P1_ADD_515_U6, P1_ADD_515_U60, P1_ADD_515_U61, P1_ADD_515_U62, P1_ADD_515_U63, P1_ADD_515_U64, P1_ADD_515_U65, P1_ADD_515_U66, P1_ADD_515_U67, P1_ADD_515_U68, P1_ADD_515_U69, P1_ADD_515_U7, P1_ADD_515_U70, P1_ADD_515_U71, P1_ADD_515_U72, P1_ADD_515_U73, P1_ADD_515_U74, P1_ADD_515_U75, P1_ADD_515_U76, P1_ADD_515_U77, P1_ADD_515_U78, P1_ADD_515_U79, P1_ADD_515_U8, P1_ADD_515_U80, P1_ADD_515_U81, P1_ADD_515_U82, P1_ADD_515_U83, P1_ADD_515_U84, P1_ADD_515_U85, P1_ADD_515_U86, P1_ADD_515_U87, P1_ADD_515_U88, P1_ADD_515_U89, P1_ADD_515_U9, P1_ADD_515_U90, P1_ADD_515_U91, P1_ADD_515_U92, P1_ADD_515_U93, P1_ADD_515_U94, P1_ADD_515_U95, P1_ADD_515_U96, P1_ADD_515_U97, P1_ADD_515_U98, P1_ADD_515_U99, P1_GTE_485_U6, P1_GTE_485_U7, P1_LT_563_1260_U6, P1_LT_563_1260_U7, P1_LT_563_1260_U8, P1_LT_563_1260_U9, P1_LT_563_U10, P1_LT_563_U11, P1_LT_563_U12, P1_LT_563_U13, P1_LT_563_U14, P1_LT_563_U15, P1_LT_563_U16, P1_LT_563_U17, P1_LT_563_U18, P1_LT_563_U19, P1_LT_563_U20, P1_LT_563_U21, P1_LT_563_U22, P1_LT_563_U23, P1_LT_563_U24, P1_LT_563_U25, P1_LT_563_U26, P1_LT_563_U27, P1_LT_563_U28, P1_LT_563_U6, P1_LT_563_U7, P1_LT_563_U8, P1_LT_563_U9, P1_LT_589_U6, P1_LT_589_U7, P1_LT_589_U8, P1_R2027_U10, P1_R2027_U100, P1_R2027_U101, P1_R2027_U102, P1_R2027_U103, P1_R2027_U104, P1_R2027_U105, P1_R2027_U106, P1_R2027_U107, P1_R2027_U108, P1_R2027_U109, P1_R2027_U11, P1_R2027_U110, P1_R2027_U111, P1_R2027_U112, P1_R2027_U113, P1_R2027_U114, P1_R2027_U115, P1_R2027_U116, P1_R2027_U117, P1_R2027_U118, P1_R2027_U119, P1_R2027_U12, P1_R2027_U120, P1_R2027_U121, P1_R2027_U122, P1_R2027_U123, P1_R2027_U124, P1_R2027_U125, P1_R2027_U126, P1_R2027_U127, P1_R2027_U128, P1_R2027_U129, P1_R2027_U13, P1_R2027_U130, P1_R2027_U131, P1_R2027_U132, P1_R2027_U133, P1_R2027_U134, P1_R2027_U135, P1_R2027_U136, P1_R2027_U137, P1_R2027_U138, P1_R2027_U139, P1_R2027_U14, P1_R2027_U140, P1_R2027_U141, P1_R2027_U142, P1_R2027_U143, P1_R2027_U144, P1_R2027_U145, P1_R2027_U146, P1_R2027_U147, P1_R2027_U148, P1_R2027_U149, P1_R2027_U15, P1_R2027_U150, P1_R2027_U151, P1_R2027_U152, P1_R2027_U153, P1_R2027_U154, P1_R2027_U155, P1_R2027_U156, P1_R2027_U157, P1_R2027_U158, P1_R2027_U159, P1_R2027_U16, P1_R2027_U160, P1_R2027_U161, P1_R2027_U162, P1_R2027_U163, P1_R2027_U164, P1_R2027_U165, P1_R2027_U166, P1_R2027_U167, P1_R2027_U168, P1_R2027_U169, P1_R2027_U17, P1_R2027_U170, P1_R2027_U171, P1_R2027_U172, P1_R2027_U173, P1_R2027_U174, P1_R2027_U175, P1_R2027_U176, P1_R2027_U177, P1_R2027_U178, P1_R2027_U179, P1_R2027_U18, P1_R2027_U180, P1_R2027_U181, P1_R2027_U182, P1_R2027_U183, P1_R2027_U184, P1_R2027_U185, P1_R2027_U186, P1_R2027_U187, P1_R2027_U188, P1_R2027_U189, P1_R2027_U19, P1_R2027_U190, P1_R2027_U191, P1_R2027_U192, P1_R2027_U193, P1_R2027_U194, P1_R2027_U195, P1_R2027_U196, P1_R2027_U197, P1_R2027_U198, P1_R2027_U199, P1_R2027_U20, P1_R2027_U200, P1_R2027_U201, P1_R2027_U202, P1_R2027_U21, P1_R2027_U22, P1_R2027_U23, P1_R2027_U24, P1_R2027_U25, P1_R2027_U26, P1_R2027_U27, P1_R2027_U28, P1_R2027_U29, P1_R2027_U30, P1_R2027_U31, P1_R2027_U32, P1_R2027_U33, P1_R2027_U34, P1_R2027_U35, P1_R2027_U36, P1_R2027_U37, P1_R2027_U38, P1_R2027_U39, P1_R2027_U40, P1_R2027_U41, P1_R2027_U42, P1_R2027_U43, P1_R2027_U44, P1_R2027_U45, P1_R2027_U46, P1_R2027_U47, P1_R2027_U48, P1_R2027_U49, P1_R2027_U5, P1_R2027_U50, P1_R2027_U51, P1_R2027_U52, P1_R2027_U53, P1_R2027_U54, P1_R2027_U55, P1_R2027_U56, P1_R2027_U57, P1_R2027_U58, P1_R2027_U59, P1_R2027_U6, P1_R2027_U60, P1_R2027_U61, P1_R2027_U62, P1_R2027_U63, P1_R2027_U64, P1_R2027_U65, P1_R2027_U66, P1_R2027_U67, P1_R2027_U68, P1_R2027_U69, P1_R2027_U7, P1_R2027_U70, P1_R2027_U71, P1_R2027_U72, P1_R2027_U73, P1_R2027_U74, P1_R2027_U75, P1_R2027_U76, P1_R2027_U77, P1_R2027_U78, P1_R2027_U79, P1_R2027_U8, P1_R2027_U80, P1_R2027_U81, P1_R2027_U82, P1_R2027_U83, P1_R2027_U84, P1_R2027_U85, P1_R2027_U86, P1_R2027_U87, P1_R2027_U88, P1_R2027_U89, P1_R2027_U9, P1_R2027_U90, P1_R2027_U91, P1_R2027_U92, P1_R2027_U93, P1_R2027_U94, P1_R2027_U95, P1_R2027_U96, P1_R2027_U97, P1_R2027_U98, P1_R2027_U99, P1_R2096_U10, P1_R2096_U100, P1_R2096_U101, P1_R2096_U102, P1_R2096_U103, P1_R2096_U104, P1_R2096_U105, P1_R2096_U106, P1_R2096_U107, P1_R2096_U108, P1_R2096_U109, P1_R2096_U11, P1_R2096_U110, P1_R2096_U111, P1_R2096_U112, P1_R2096_U113, P1_R2096_U114, P1_R2096_U115, P1_R2096_U116, P1_R2096_U117, P1_R2096_U118, P1_R2096_U119, P1_R2096_U12, P1_R2096_U120, P1_R2096_U121, P1_R2096_U122, P1_R2096_U123, P1_R2096_U124, P1_R2096_U125, P1_R2096_U126, P1_R2096_U127, P1_R2096_U128, P1_R2096_U129, P1_R2096_U13, P1_R2096_U130, P1_R2096_U131, P1_R2096_U132, P1_R2096_U133, P1_R2096_U134, P1_R2096_U135, P1_R2096_U136, P1_R2096_U137, P1_R2096_U138, P1_R2096_U139, P1_R2096_U14, P1_R2096_U140, P1_R2096_U141, P1_R2096_U142, P1_R2096_U143, P1_R2096_U144, P1_R2096_U145, P1_R2096_U146, P1_R2096_U147, P1_R2096_U148, P1_R2096_U149, P1_R2096_U15, P1_R2096_U150, P1_R2096_U151, P1_R2096_U152, P1_R2096_U153, P1_R2096_U154, P1_R2096_U155, P1_R2096_U156, P1_R2096_U157, P1_R2096_U158, P1_R2096_U159, P1_R2096_U16, P1_R2096_U160, P1_R2096_U161, P1_R2096_U162, P1_R2096_U163, P1_R2096_U164, P1_R2096_U165, P1_R2096_U166, P1_R2096_U167, P1_R2096_U168, P1_R2096_U169, P1_R2096_U17, P1_R2096_U170, P1_R2096_U171, P1_R2096_U172, P1_R2096_U173, P1_R2096_U174, P1_R2096_U175, P1_R2096_U176, P1_R2096_U177, P1_R2096_U178, P1_R2096_U179, P1_R2096_U18, P1_R2096_U180, P1_R2096_U181, P1_R2096_U182, P1_R2096_U19, P1_R2096_U20, P1_R2096_U21, P1_R2096_U22, P1_R2096_U23, P1_R2096_U24, P1_R2096_U25, P1_R2096_U26, P1_R2096_U27, P1_R2096_U28, P1_R2096_U29, P1_R2096_U30, P1_R2096_U31, P1_R2096_U32, P1_R2096_U33, P1_R2096_U34, P1_R2096_U35, P1_R2096_U36, P1_R2096_U37, P1_R2096_U38, P1_R2096_U39, P1_R2096_U4, P1_R2096_U40, P1_R2096_U41, P1_R2096_U42, P1_R2096_U43, P1_R2096_U44, P1_R2096_U45, P1_R2096_U46, P1_R2096_U47, P1_R2096_U48, P1_R2096_U49, P1_R2096_U5, P1_R2096_U50, P1_R2096_U51, P1_R2096_U52, P1_R2096_U53, P1_R2096_U54, P1_R2096_U55, P1_R2096_U56, P1_R2096_U57, P1_R2096_U58, P1_R2096_U59, P1_R2096_U6, P1_R2096_U60, P1_R2096_U61, P1_R2096_U62, P1_R2096_U63, P1_R2096_U64, P1_R2096_U65, P1_R2096_U66, P1_R2096_U67, P1_R2096_U68, P1_R2096_U69, P1_R2096_U7, P1_R2096_U70, P1_R2096_U71, P1_R2096_U72, P1_R2096_U73, P1_R2096_U74, P1_R2096_U75, P1_R2096_U76, P1_R2096_U77, P1_R2096_U78, P1_R2096_U79, P1_R2096_U8, P1_R2096_U80, P1_R2096_U81, P1_R2096_U82, P1_R2096_U83, P1_R2096_U84, P1_R2096_U85, P1_R2096_U86, P1_R2096_U87, P1_R2096_U88, P1_R2096_U89, P1_R2096_U9, P1_R2096_U90, P1_R2096_U91, P1_R2096_U92, P1_R2096_U93, P1_R2096_U94, P1_R2096_U95, P1_R2096_U96, P1_R2096_U97, P1_R2096_U98, P1_R2096_U99, P1_R2099_U10, P1_R2099_U100, P1_R2099_U101, P1_R2099_U102, P1_R2099_U103, P1_R2099_U104, P1_R2099_U105, P1_R2099_U106, P1_R2099_U107, P1_R2099_U108, P1_R2099_U109, P1_R2099_U11, P1_R2099_U110, P1_R2099_U111, P1_R2099_U112, P1_R2099_U113, P1_R2099_U114, P1_R2099_U115, P1_R2099_U116, P1_R2099_U117, P1_R2099_U118, P1_R2099_U119, P1_R2099_U12, P1_R2099_U120, P1_R2099_U121, P1_R2099_U122, P1_R2099_U123, P1_R2099_U124, P1_R2099_U125, P1_R2099_U126, P1_R2099_U127, P1_R2099_U128, P1_R2099_U129, P1_R2099_U13, P1_R2099_U130, P1_R2099_U131, P1_R2099_U132, P1_R2099_U133, P1_R2099_U134, P1_R2099_U135, P1_R2099_U136, P1_R2099_U137, P1_R2099_U138, P1_R2099_U139, P1_R2099_U14, P1_R2099_U140, P1_R2099_U141, P1_R2099_U142, P1_R2099_U143, P1_R2099_U144, P1_R2099_U145, P1_R2099_U146, P1_R2099_U147, P1_R2099_U148, P1_R2099_U149, P1_R2099_U15, P1_R2099_U150, P1_R2099_U151, P1_R2099_U152, P1_R2099_U153, P1_R2099_U154, P1_R2099_U155, P1_R2099_U156, P1_R2099_U157, P1_R2099_U158, P1_R2099_U159, P1_R2099_U16, P1_R2099_U160, P1_R2099_U161, P1_R2099_U162, P1_R2099_U163, P1_R2099_U164, P1_R2099_U165, P1_R2099_U166, P1_R2099_U167, P1_R2099_U168, P1_R2099_U169, P1_R2099_U17, P1_R2099_U170, P1_R2099_U171, P1_R2099_U172, P1_R2099_U173, P1_R2099_U174, P1_R2099_U175, P1_R2099_U176, P1_R2099_U177, P1_R2099_U178, P1_R2099_U179, P1_R2099_U18, P1_R2099_U180, P1_R2099_U181, P1_R2099_U182, P1_R2099_U183, P1_R2099_U184, P1_R2099_U185, P1_R2099_U186, P1_R2099_U187, P1_R2099_U188, P1_R2099_U189, P1_R2099_U19, P1_R2099_U190, P1_R2099_U191, P1_R2099_U192, P1_R2099_U193, P1_R2099_U194, P1_R2099_U195, P1_R2099_U196, P1_R2099_U197, P1_R2099_U198, P1_R2099_U199, P1_R2099_U20, P1_R2099_U200, P1_R2099_U201, P1_R2099_U202, P1_R2099_U203, P1_R2099_U204, P1_R2099_U205, P1_R2099_U206, P1_R2099_U207, P1_R2099_U208, P1_R2099_U209, P1_R2099_U21, P1_R2099_U210, P1_R2099_U211, P1_R2099_U212, P1_R2099_U213, P1_R2099_U214, P1_R2099_U215, P1_R2099_U216, P1_R2099_U217, P1_R2099_U218, P1_R2099_U219, P1_R2099_U22, P1_R2099_U220, P1_R2099_U221, P1_R2099_U222, P1_R2099_U223, P1_R2099_U224, P1_R2099_U225, P1_R2099_U226, P1_R2099_U227, P1_R2099_U228, P1_R2099_U229, P1_R2099_U23, P1_R2099_U230, P1_R2099_U231, P1_R2099_U232, P1_R2099_U233, P1_R2099_U234, P1_R2099_U235, P1_R2099_U236, P1_R2099_U237, P1_R2099_U238, P1_R2099_U239, P1_R2099_U24, P1_R2099_U240, P1_R2099_U241, P1_R2099_U242, P1_R2099_U243, P1_R2099_U244, P1_R2099_U245, P1_R2099_U246, P1_R2099_U247, P1_R2099_U248, P1_R2099_U249, P1_R2099_U25, P1_R2099_U250, P1_R2099_U251, P1_R2099_U252, P1_R2099_U253, P1_R2099_U254, P1_R2099_U255, P1_R2099_U256, P1_R2099_U257, P1_R2099_U258, P1_R2099_U259, P1_R2099_U26, P1_R2099_U260, P1_R2099_U261, P1_R2099_U262, P1_R2099_U263, P1_R2099_U264, P1_R2099_U265, P1_R2099_U266, P1_R2099_U267, P1_R2099_U268, P1_R2099_U269, P1_R2099_U27, P1_R2099_U270, P1_R2099_U271, P1_R2099_U272, P1_R2099_U273, P1_R2099_U274, P1_R2099_U275, P1_R2099_U276, P1_R2099_U277, P1_R2099_U278, P1_R2099_U279, P1_R2099_U28, P1_R2099_U280, P1_R2099_U281, P1_R2099_U282, P1_R2099_U283, P1_R2099_U284, P1_R2099_U285, P1_R2099_U286, P1_R2099_U287, P1_R2099_U288, P1_R2099_U289, P1_R2099_U29, P1_R2099_U290, P1_R2099_U291, P1_R2099_U292, P1_R2099_U293, P1_R2099_U294, P1_R2099_U295, P1_R2099_U296, P1_R2099_U297, P1_R2099_U298, P1_R2099_U299, P1_R2099_U30, P1_R2099_U300, P1_R2099_U301, P1_R2099_U302, P1_R2099_U303, P1_R2099_U304, P1_R2099_U305, P1_R2099_U306, P1_R2099_U307, P1_R2099_U308, P1_R2099_U309, P1_R2099_U31, P1_R2099_U310, P1_R2099_U311, P1_R2099_U312, P1_R2099_U313, P1_R2099_U314, P1_R2099_U315, P1_R2099_U316, P1_R2099_U317, P1_R2099_U318, P1_R2099_U319, P1_R2099_U32, P1_R2099_U320, P1_R2099_U321, P1_R2099_U322, P1_R2099_U323, P1_R2099_U324, P1_R2099_U325, P1_R2099_U326, P1_R2099_U327, P1_R2099_U328, P1_R2099_U329, P1_R2099_U33, P1_R2099_U330, P1_R2099_U331, P1_R2099_U332, P1_R2099_U333, P1_R2099_U334, P1_R2099_U335, P1_R2099_U336, P1_R2099_U337, P1_R2099_U338, P1_R2099_U339, P1_R2099_U34, P1_R2099_U340, P1_R2099_U341, P1_R2099_U342, P1_R2099_U343, P1_R2099_U344, P1_R2099_U345, P1_R2099_U346, P1_R2099_U347, P1_R2099_U348, P1_R2099_U349, P1_R2099_U35, P1_R2099_U36, P1_R2099_U37, P1_R2099_U38, P1_R2099_U39, P1_R2099_U4, P1_R2099_U40, P1_R2099_U41, P1_R2099_U42, P1_R2099_U43, P1_R2099_U44, P1_R2099_U45, P1_R2099_U46, P1_R2099_U47, P1_R2099_U48, P1_R2099_U49, P1_R2099_U5, P1_R2099_U50, P1_R2099_U51, P1_R2099_U52, P1_R2099_U53, P1_R2099_U54, P1_R2099_U55, P1_R2099_U56, P1_R2099_U57, P1_R2099_U58, P1_R2099_U59, P1_R2099_U6, P1_R2099_U60, P1_R2099_U61, P1_R2099_U62, P1_R2099_U63, P1_R2099_U64, P1_R2099_U65, P1_R2099_U66, P1_R2099_U67, P1_R2099_U68, P1_R2099_U69, P1_R2099_U7, P1_R2099_U70, P1_R2099_U71, P1_R2099_U72, P1_R2099_U73, P1_R2099_U74, P1_R2099_U75, P1_R2099_U76, P1_R2099_U77, P1_R2099_U78, P1_R2099_U79, P1_R2099_U8, P1_R2099_U80, P1_R2099_U81, P1_R2099_U82, P1_R2099_U83, P1_R2099_U84, P1_R2099_U85, P1_R2099_U86, P1_R2099_U87, P1_R2099_U88, P1_R2099_U89, P1_R2099_U9, P1_R2099_U90, P1_R2099_U91, P1_R2099_U92, P1_R2099_U93, P1_R2099_U94, P1_R2099_U95, P1_R2099_U96, P1_R2099_U97, P1_R2099_U98, P1_R2099_U99, P1_R2144_U10, P1_R2144_U100, P1_R2144_U101, P1_R2144_U102, P1_R2144_U103, P1_R2144_U104, P1_R2144_U105, P1_R2144_U106, P1_R2144_U107, P1_R2144_U108, P1_R2144_U109, P1_R2144_U11, P1_R2144_U110, P1_R2144_U111, P1_R2144_U112, P1_R2144_U113, P1_R2144_U114, P1_R2144_U115, P1_R2144_U116, P1_R2144_U117, P1_R2144_U118, P1_R2144_U119, P1_R2144_U12, P1_R2144_U120, P1_R2144_U121, P1_R2144_U122, P1_R2144_U123, P1_R2144_U124, P1_R2144_U125, P1_R2144_U126, P1_R2144_U127, P1_R2144_U128, P1_R2144_U129, P1_R2144_U13, P1_R2144_U130, P1_R2144_U131, P1_R2144_U132, P1_R2144_U133, P1_R2144_U134, P1_R2144_U135, P1_R2144_U136, P1_R2144_U137, P1_R2144_U138, P1_R2144_U139, P1_R2144_U14, P1_R2144_U140, P1_R2144_U141, P1_R2144_U142, P1_R2144_U143, P1_R2144_U144, P1_R2144_U145, P1_R2144_U146, P1_R2144_U147, P1_R2144_U148, P1_R2144_U149, P1_R2144_U15, P1_R2144_U150, P1_R2144_U151, P1_R2144_U152, P1_R2144_U153, P1_R2144_U154, P1_R2144_U155, P1_R2144_U156, P1_R2144_U157, P1_R2144_U158, P1_R2144_U159, P1_R2144_U16, P1_R2144_U160, P1_R2144_U161, P1_R2144_U162, P1_R2144_U163, P1_R2144_U164, P1_R2144_U165, P1_R2144_U166, P1_R2144_U167, P1_R2144_U168, P1_R2144_U169, P1_R2144_U17, P1_R2144_U170, P1_R2144_U171, P1_R2144_U172, P1_R2144_U173, P1_R2144_U174, P1_R2144_U175, P1_R2144_U176, P1_R2144_U177, P1_R2144_U178, P1_R2144_U179, P1_R2144_U18, P1_R2144_U180, P1_R2144_U181, P1_R2144_U182, P1_R2144_U183, P1_R2144_U184, P1_R2144_U185, P1_R2144_U186, P1_R2144_U187, P1_R2144_U188, P1_R2144_U189, P1_R2144_U19, P1_R2144_U190, P1_R2144_U191, P1_R2144_U192, P1_R2144_U193, P1_R2144_U194, P1_R2144_U195, P1_R2144_U196, P1_R2144_U197, P1_R2144_U198, P1_R2144_U199, P1_R2144_U20, P1_R2144_U200, P1_R2144_U201, P1_R2144_U202, P1_R2144_U203, P1_R2144_U204, P1_R2144_U205, P1_R2144_U206, P1_R2144_U207, P1_R2144_U208, P1_R2144_U209, P1_R2144_U21, P1_R2144_U210, P1_R2144_U211, P1_R2144_U212, P1_R2144_U213, P1_R2144_U214, P1_R2144_U215, P1_R2144_U216, P1_R2144_U217, P1_R2144_U218, P1_R2144_U219, P1_R2144_U22, P1_R2144_U220, P1_R2144_U221, P1_R2144_U222, P1_R2144_U223, P1_R2144_U224, P1_R2144_U225, P1_R2144_U226, P1_R2144_U227, P1_R2144_U228, P1_R2144_U229, P1_R2144_U23, P1_R2144_U230, P1_R2144_U231, P1_R2144_U232, P1_R2144_U233, P1_R2144_U234, P1_R2144_U235, P1_R2144_U236, P1_R2144_U237, P1_R2144_U238, P1_R2144_U239, P1_R2144_U24, P1_R2144_U240, P1_R2144_U241, P1_R2144_U242, P1_R2144_U243, P1_R2144_U244, P1_R2144_U245, P1_R2144_U246, P1_R2144_U247, P1_R2144_U248, P1_R2144_U249, P1_R2144_U25, P1_R2144_U250, P1_R2144_U251, P1_R2144_U252, P1_R2144_U253, P1_R2144_U254, P1_R2144_U255, P1_R2144_U256, P1_R2144_U257, P1_R2144_U258, P1_R2144_U259, P1_R2144_U26, P1_R2144_U260, P1_R2144_U27, P1_R2144_U28, P1_R2144_U29, P1_R2144_U30, P1_R2144_U31, P1_R2144_U32, P1_R2144_U33, P1_R2144_U34, P1_R2144_U35, P1_R2144_U36, P1_R2144_U37, P1_R2144_U38, P1_R2144_U39, P1_R2144_U40, P1_R2144_U41, P1_R2144_U42, P1_R2144_U43, P1_R2144_U44, P1_R2144_U45, P1_R2144_U46, P1_R2144_U47, P1_R2144_U48, P1_R2144_U49, P1_R2144_U5, P1_R2144_U50, P1_R2144_U51, P1_R2144_U52, P1_R2144_U53, P1_R2144_U54, P1_R2144_U55, P1_R2144_U56, P1_R2144_U57, P1_R2144_U58, P1_R2144_U59, P1_R2144_U6, P1_R2144_U60, P1_R2144_U61, P1_R2144_U62, P1_R2144_U63, P1_R2144_U64, P1_R2144_U65, P1_R2144_U66, P1_R2144_U67, P1_R2144_U68, P1_R2144_U69, P1_R2144_U7, P1_R2144_U70, P1_R2144_U71, P1_R2144_U72, P1_R2144_U73, P1_R2144_U74, P1_R2144_U75, P1_R2144_U76, P1_R2144_U77, P1_R2144_U78, P1_R2144_U79, P1_R2144_U8, P1_R2144_U80, P1_R2144_U81, P1_R2144_U82, P1_R2144_U83, P1_R2144_U84, P1_R2144_U85, P1_R2144_U86, P1_R2144_U87, P1_R2144_U88, P1_R2144_U89, P1_R2144_U9, P1_R2144_U90, P1_R2144_U91, P1_R2144_U92, P1_R2144_U93, P1_R2144_U94, P1_R2144_U95, P1_R2144_U96, P1_R2144_U97, P1_R2144_U98, P1_R2144_U99, P1_R2167_U10, P1_R2167_U11, P1_R2167_U12, P1_R2167_U13, P1_R2167_U14, P1_R2167_U15, P1_R2167_U16, P1_R2167_U17, P1_R2167_U18, P1_R2167_U19, P1_R2167_U20, P1_R2167_U21, P1_R2167_U22, P1_R2167_U23, P1_R2167_U24, P1_R2167_U25, P1_R2167_U26, P1_R2167_U27, P1_R2167_U28, P1_R2167_U29, P1_R2167_U30, P1_R2167_U31, P1_R2167_U32, P1_R2167_U33, P1_R2167_U34, P1_R2167_U35, P1_R2167_U36, P1_R2167_U37, P1_R2167_U38, P1_R2167_U39, P1_R2167_U40, P1_R2167_U41, P1_R2167_U42, P1_R2167_U43, P1_R2167_U44, P1_R2167_U45, P1_R2167_U46, P1_R2167_U47, P1_R2167_U48, P1_R2167_U49, P1_R2167_U50, P1_R2167_U6, P1_R2167_U7, P1_R2167_U8, P1_R2167_U9, P1_R2182_U10, P1_R2182_U11, P1_R2182_U12, P1_R2182_U13, P1_R2182_U14, P1_R2182_U15, P1_R2182_U16, P1_R2182_U17, P1_R2182_U18, P1_R2182_U19, P1_R2182_U20, P1_R2182_U21, P1_R2182_U22, P1_R2182_U23, P1_R2182_U24, P1_R2182_U25, P1_R2182_U26, P1_R2182_U27, P1_R2182_U28, P1_R2182_U29, P1_R2182_U30, P1_R2182_U31, P1_R2182_U32, P1_R2182_U33, P1_R2182_U34, P1_R2182_U35, P1_R2182_U36, P1_R2182_U37, P1_R2182_U38, P1_R2182_U39, P1_R2182_U40, P1_R2182_U41, P1_R2182_U42, P1_R2182_U43, P1_R2182_U44, P1_R2182_U45, P1_R2182_U46, P1_R2182_U47, P1_R2182_U48, P1_R2182_U49, P1_R2182_U5, P1_R2182_U50, P1_R2182_U51, P1_R2182_U52, P1_R2182_U53, P1_R2182_U54, P1_R2182_U55, P1_R2182_U56, P1_R2182_U57, P1_R2182_U58, P1_R2182_U59, P1_R2182_U6, P1_R2182_U60, P1_R2182_U61, P1_R2182_U62, P1_R2182_U63, P1_R2182_U64, P1_R2182_U65, P1_R2182_U66, P1_R2182_U67, P1_R2182_U68, P1_R2182_U69, P1_R2182_U7, P1_R2182_U70, P1_R2182_U71, P1_R2182_U72, P1_R2182_U73, P1_R2182_U74, P1_R2182_U75, P1_R2182_U76, P1_R2182_U77, P1_R2182_U78, P1_R2182_U79, P1_R2182_U8, P1_R2182_U80, P1_R2182_U81, P1_R2182_U82, P1_R2182_U83, P1_R2182_U84, P1_R2182_U85, P1_R2182_U86, P1_R2182_U9, P1_R2238_U10, P1_R2238_U11, P1_R2238_U12, P1_R2238_U13, P1_R2238_U14, P1_R2238_U15, P1_R2238_U16, P1_R2238_U17, P1_R2238_U18, P1_R2238_U19, P1_R2238_U20, P1_R2238_U21, P1_R2238_U22, P1_R2238_U23, P1_R2238_U24, P1_R2238_U25, P1_R2238_U26, P1_R2238_U27, P1_R2238_U28, P1_R2238_U29, P1_R2238_U30, P1_R2238_U31, P1_R2238_U32, P1_R2238_U33, P1_R2238_U34, P1_R2238_U35, P1_R2238_U36, P1_R2238_U37, P1_R2238_U38, P1_R2238_U39, P1_R2238_U40, P1_R2238_U41, P1_R2238_U42, P1_R2238_U43, P1_R2238_U44, P1_R2238_U45, P1_R2238_U46, P1_R2238_U47, P1_R2238_U48, P1_R2238_U49, P1_R2238_U50, P1_R2238_U51, P1_R2238_U52, P1_R2238_U53, P1_R2238_U54, P1_R2238_U55, P1_R2238_U56, P1_R2238_U57, P1_R2238_U58, P1_R2238_U59, P1_R2238_U6, P1_R2238_U60, P1_R2238_U61, P1_R2238_U62, P1_R2238_U63, P1_R2238_U64, P1_R2238_U65, P1_R2238_U66, P1_R2238_U7, P1_R2238_U8, P1_R2238_U9, P1_R2278_U10, P1_R2278_U100, P1_R2278_U101, P1_R2278_U102, P1_R2278_U103, P1_R2278_U104, P1_R2278_U105, P1_R2278_U106, P1_R2278_U107, P1_R2278_U108, P1_R2278_U109, P1_R2278_U11, P1_R2278_U110, P1_R2278_U111, P1_R2278_U112, P1_R2278_U113, P1_R2278_U114, P1_R2278_U115, P1_R2278_U116, P1_R2278_U117, P1_R2278_U118, P1_R2278_U119, P1_R2278_U12, P1_R2278_U120, P1_R2278_U121, P1_R2278_U122, P1_R2278_U123, P1_R2278_U124, P1_R2278_U125, P1_R2278_U126, P1_R2278_U127, P1_R2278_U128, P1_R2278_U129, P1_R2278_U13, P1_R2278_U130, P1_R2278_U131, P1_R2278_U132, P1_R2278_U133, P1_R2278_U134, P1_R2278_U135, P1_R2278_U136, P1_R2278_U137, P1_R2278_U138, P1_R2278_U139, P1_R2278_U14, P1_R2278_U140, P1_R2278_U141, P1_R2278_U142, P1_R2278_U143, P1_R2278_U144, P1_R2278_U145, P1_R2278_U146, P1_R2278_U147, P1_R2278_U148, P1_R2278_U149, P1_R2278_U15, P1_R2278_U150, P1_R2278_U151, P1_R2278_U152, P1_R2278_U153, P1_R2278_U154, P1_R2278_U155, P1_R2278_U156, P1_R2278_U157, P1_R2278_U158, P1_R2278_U159, P1_R2278_U16, P1_R2278_U160, P1_R2278_U161, P1_R2278_U162, P1_R2278_U163, P1_R2278_U164, P1_R2278_U165, P1_R2278_U166, P1_R2278_U167, P1_R2278_U168, P1_R2278_U169, P1_R2278_U17, P1_R2278_U170, P1_R2278_U171, P1_R2278_U172, P1_R2278_U173, P1_R2278_U174, P1_R2278_U175, P1_R2278_U176, P1_R2278_U177, P1_R2278_U178, P1_R2278_U179, P1_R2278_U18, P1_R2278_U180, P1_R2278_U181, P1_R2278_U182, P1_R2278_U183, P1_R2278_U184, P1_R2278_U185, P1_R2278_U186, P1_R2278_U187, P1_R2278_U188, P1_R2278_U189, P1_R2278_U19, P1_R2278_U190, P1_R2278_U191, P1_R2278_U192, P1_R2278_U193, P1_R2278_U194, P1_R2278_U195, P1_R2278_U196, P1_R2278_U197, P1_R2278_U198, P1_R2278_U199, P1_R2278_U20, P1_R2278_U200, P1_R2278_U201, P1_R2278_U202, P1_R2278_U203, P1_R2278_U204, P1_R2278_U205, P1_R2278_U206, P1_R2278_U207, P1_R2278_U208, P1_R2278_U209, P1_R2278_U21, P1_R2278_U210, P1_R2278_U211, P1_R2278_U212, P1_R2278_U213, P1_R2278_U214, P1_R2278_U215, P1_R2278_U216, P1_R2278_U217, P1_R2278_U218, P1_R2278_U219, P1_R2278_U22, P1_R2278_U220, P1_R2278_U221, P1_R2278_U222, P1_R2278_U223, P1_R2278_U224, P1_R2278_U225, P1_R2278_U226, P1_R2278_U227, P1_R2278_U228, P1_R2278_U229, P1_R2278_U23, P1_R2278_U230, P1_R2278_U231, P1_R2278_U232, P1_R2278_U233, P1_R2278_U234, P1_R2278_U235, P1_R2278_U236, P1_R2278_U237, P1_R2278_U238, P1_R2278_U239, P1_R2278_U24, P1_R2278_U240, P1_R2278_U241, P1_R2278_U242, P1_R2278_U243, P1_R2278_U244, P1_R2278_U245, P1_R2278_U246, P1_R2278_U247, P1_R2278_U248, P1_R2278_U249, P1_R2278_U25, P1_R2278_U250, P1_R2278_U251, P1_R2278_U252, P1_R2278_U253, P1_R2278_U254, P1_R2278_U255, P1_R2278_U256, P1_R2278_U257, P1_R2278_U258, P1_R2278_U259, P1_R2278_U26, P1_R2278_U260, P1_R2278_U261, P1_R2278_U262, P1_R2278_U263, P1_R2278_U264, P1_R2278_U265, P1_R2278_U266, P1_R2278_U267, P1_R2278_U268, P1_R2278_U269, P1_R2278_U27, P1_R2278_U270, P1_R2278_U271, P1_R2278_U272, P1_R2278_U273, P1_R2278_U274, P1_R2278_U275, P1_R2278_U276, P1_R2278_U277, P1_R2278_U278, P1_R2278_U279, P1_R2278_U28, P1_R2278_U280, P1_R2278_U281, P1_R2278_U282, P1_R2278_U283, P1_R2278_U284, P1_R2278_U285, P1_R2278_U286, P1_R2278_U287, P1_R2278_U288, P1_R2278_U289, P1_R2278_U29, P1_R2278_U290, P1_R2278_U291, P1_R2278_U292, P1_R2278_U293, P1_R2278_U294, P1_R2278_U295, P1_R2278_U296, P1_R2278_U297, P1_R2278_U298, P1_R2278_U299, P1_R2278_U30, P1_R2278_U300, P1_R2278_U301, P1_R2278_U302, P1_R2278_U303, P1_R2278_U304, P1_R2278_U305, P1_R2278_U306, P1_R2278_U307, P1_R2278_U308, P1_R2278_U309, P1_R2278_U31, P1_R2278_U310, P1_R2278_U311, P1_R2278_U312, P1_R2278_U313, P1_R2278_U314, P1_R2278_U315, P1_R2278_U316, P1_R2278_U317, P1_R2278_U318, P1_R2278_U319, P1_R2278_U32, P1_R2278_U320, P1_R2278_U321, P1_R2278_U322, P1_R2278_U323, P1_R2278_U324, P1_R2278_U325, P1_R2278_U326, P1_R2278_U327, P1_R2278_U328, P1_R2278_U329, P1_R2278_U33, P1_R2278_U330, P1_R2278_U331, P1_R2278_U332, P1_R2278_U333, P1_R2278_U334, P1_R2278_U335, P1_R2278_U336, P1_R2278_U337, P1_R2278_U338, P1_R2278_U339, P1_R2278_U34, P1_R2278_U340, P1_R2278_U341, P1_R2278_U342, P1_R2278_U343, P1_R2278_U344, P1_R2278_U345, P1_R2278_U346, P1_R2278_U347, P1_R2278_U348, P1_R2278_U349, P1_R2278_U35, P1_R2278_U350, P1_R2278_U351, P1_R2278_U352, P1_R2278_U353, P1_R2278_U354, P1_R2278_U355, P1_R2278_U356, P1_R2278_U357, P1_R2278_U358, P1_R2278_U359, P1_R2278_U36, P1_R2278_U360, P1_R2278_U361, P1_R2278_U362, P1_R2278_U363, P1_R2278_U364, P1_R2278_U365, P1_R2278_U366, P1_R2278_U367, P1_R2278_U368, P1_R2278_U369, P1_R2278_U37, P1_R2278_U370, P1_R2278_U371, P1_R2278_U372, P1_R2278_U373, P1_R2278_U374, P1_R2278_U375, P1_R2278_U376, P1_R2278_U377, P1_R2278_U378, P1_R2278_U379, P1_R2278_U38, P1_R2278_U380, P1_R2278_U381, P1_R2278_U382, P1_R2278_U383, P1_R2278_U384, P1_R2278_U385, P1_R2278_U386, P1_R2278_U387, P1_R2278_U388, P1_R2278_U389, P1_R2278_U39, P1_R2278_U390, P1_R2278_U391, P1_R2278_U392, P1_R2278_U393, P1_R2278_U394, P1_R2278_U395, P1_R2278_U396, P1_R2278_U397, P1_R2278_U398, P1_R2278_U399, P1_R2278_U40, P1_R2278_U400, P1_R2278_U401, P1_R2278_U402, P1_R2278_U403, P1_R2278_U404, P1_R2278_U405, P1_R2278_U406, P1_R2278_U407, P1_R2278_U408, P1_R2278_U409, P1_R2278_U41, P1_R2278_U410, P1_R2278_U411, P1_R2278_U412, P1_R2278_U413, P1_R2278_U414, P1_R2278_U415, P1_R2278_U416, P1_R2278_U417, P1_R2278_U418, P1_R2278_U419, P1_R2278_U42, P1_R2278_U420, P1_R2278_U421, P1_R2278_U422, P1_R2278_U423, P1_R2278_U424, P1_R2278_U425, P1_R2278_U426, P1_R2278_U427, P1_R2278_U428, P1_R2278_U429, P1_R2278_U43, P1_R2278_U430, P1_R2278_U431, P1_R2278_U432, P1_R2278_U433, P1_R2278_U434, P1_R2278_U435, P1_R2278_U436, P1_R2278_U437, P1_R2278_U438, P1_R2278_U439, P1_R2278_U44, P1_R2278_U440, P1_R2278_U441, P1_R2278_U442, P1_R2278_U443, P1_R2278_U444, P1_R2278_U445, P1_R2278_U446, P1_R2278_U447, P1_R2278_U448, P1_R2278_U449, P1_R2278_U45, P1_R2278_U450, P1_R2278_U451, P1_R2278_U452, P1_R2278_U453, P1_R2278_U454, P1_R2278_U455, P1_R2278_U456, P1_R2278_U457, P1_R2278_U458, P1_R2278_U459, P1_R2278_U46, P1_R2278_U460, P1_R2278_U461, P1_R2278_U462, P1_R2278_U463, P1_R2278_U464, P1_R2278_U465, P1_R2278_U466, P1_R2278_U467, P1_R2278_U468, P1_R2278_U469, P1_R2278_U47, P1_R2278_U470, P1_R2278_U471, P1_R2278_U472, P1_R2278_U473, P1_R2278_U474, P1_R2278_U475, P1_R2278_U476, P1_R2278_U477, P1_R2278_U478, P1_R2278_U479, P1_R2278_U48, P1_R2278_U480, P1_R2278_U481, P1_R2278_U482, P1_R2278_U483, P1_R2278_U484, P1_R2278_U485, P1_R2278_U486, P1_R2278_U487, P1_R2278_U488, P1_R2278_U489, P1_R2278_U49, P1_R2278_U490, P1_R2278_U491, P1_R2278_U492, P1_R2278_U493, P1_R2278_U494, P1_R2278_U495, P1_R2278_U496, P1_R2278_U497, P1_R2278_U498, P1_R2278_U499, P1_R2278_U5, P1_R2278_U50, P1_R2278_U500, P1_R2278_U501, P1_R2278_U502, P1_R2278_U503, P1_R2278_U504, P1_R2278_U505, P1_R2278_U506, P1_R2278_U507, P1_R2278_U508, P1_R2278_U509, P1_R2278_U51, P1_R2278_U510, P1_R2278_U511, P1_R2278_U512, P1_R2278_U513, P1_R2278_U514, P1_R2278_U515, P1_R2278_U516, P1_R2278_U517, P1_R2278_U518, P1_R2278_U519, P1_R2278_U52, P1_R2278_U520, P1_R2278_U521, P1_R2278_U522, P1_R2278_U523, P1_R2278_U524, P1_R2278_U525, P1_R2278_U526, P1_R2278_U527, P1_R2278_U528, P1_R2278_U529, P1_R2278_U53, P1_R2278_U530, P1_R2278_U531, P1_R2278_U532, P1_R2278_U533, P1_R2278_U534, P1_R2278_U535, P1_R2278_U536, P1_R2278_U537, P1_R2278_U538, P1_R2278_U539, P1_R2278_U54, P1_R2278_U540, P1_R2278_U541, P1_R2278_U542, P1_R2278_U543, P1_R2278_U544, P1_R2278_U545, P1_R2278_U546, P1_R2278_U547, P1_R2278_U548, P1_R2278_U549, P1_R2278_U55, P1_R2278_U550, P1_R2278_U551, P1_R2278_U552, P1_R2278_U553, P1_R2278_U554, P1_R2278_U555, P1_R2278_U556, P1_R2278_U557, P1_R2278_U558, P1_R2278_U559, P1_R2278_U56, P1_R2278_U560, P1_R2278_U561, P1_R2278_U562, P1_R2278_U563, P1_R2278_U564, P1_R2278_U565, P1_R2278_U566, P1_R2278_U567, P1_R2278_U568, P1_R2278_U569, P1_R2278_U57, P1_R2278_U570, P1_R2278_U571, P1_R2278_U572, P1_R2278_U573, P1_R2278_U574, P1_R2278_U575, P1_R2278_U576, P1_R2278_U577, P1_R2278_U578, P1_R2278_U579, P1_R2278_U58, P1_R2278_U580, P1_R2278_U581, P1_R2278_U582, P1_R2278_U583, P1_R2278_U584, P1_R2278_U585, P1_R2278_U586, P1_R2278_U587, P1_R2278_U588, P1_R2278_U589, P1_R2278_U59, P1_R2278_U590, P1_R2278_U591, P1_R2278_U592, P1_R2278_U593, P1_R2278_U594, P1_R2278_U595, P1_R2278_U596, P1_R2278_U597, P1_R2278_U598, P1_R2278_U599, P1_R2278_U6, P1_R2278_U60, P1_R2278_U600, P1_R2278_U601, P1_R2278_U602, P1_R2278_U603, P1_R2278_U604, P1_R2278_U605, P1_R2278_U606, P1_R2278_U607, P1_R2278_U608, P1_R2278_U609, P1_R2278_U61, P1_R2278_U610, P1_R2278_U62, P1_R2278_U63, P1_R2278_U64, P1_R2278_U65, P1_R2278_U66, P1_R2278_U67, P1_R2278_U68, P1_R2278_U69, P1_R2278_U7, P1_R2278_U70, P1_R2278_U71, P1_R2278_U72, P1_R2278_U73, P1_R2278_U74, P1_R2278_U75, P1_R2278_U76, P1_R2278_U77, P1_R2278_U78, P1_R2278_U79, P1_R2278_U8, P1_R2278_U80, P1_R2278_U81, P1_R2278_U82, P1_R2278_U83, P1_R2278_U84, P1_R2278_U85, P1_R2278_U86, P1_R2278_U87, P1_R2278_U88, P1_R2278_U89, P1_R2278_U9, P1_R2278_U90, P1_R2278_U91, P1_R2278_U92, P1_R2278_U93, P1_R2278_U94, P1_R2278_U95, P1_R2278_U96, P1_R2278_U97, P1_R2278_U98, P1_R2278_U99, P1_R2337_U10, P1_R2337_U100, P1_R2337_U101, P1_R2337_U102, P1_R2337_U103, P1_R2337_U104, P1_R2337_U105, P1_R2337_U106, P1_R2337_U107, P1_R2337_U108, P1_R2337_U109, P1_R2337_U11, P1_R2337_U110, P1_R2337_U111, P1_R2337_U112, P1_R2337_U113, P1_R2337_U114, P1_R2337_U115, P1_R2337_U116, P1_R2337_U117, P1_R2337_U118, P1_R2337_U119, P1_R2337_U12, P1_R2337_U120, P1_R2337_U121, P1_R2337_U122, P1_R2337_U123, P1_R2337_U124, P1_R2337_U125, P1_R2337_U126, P1_R2337_U127, P1_R2337_U128, P1_R2337_U129, P1_R2337_U13, P1_R2337_U130, P1_R2337_U131, P1_R2337_U132, P1_R2337_U133, P1_R2337_U134, P1_R2337_U135, P1_R2337_U136, P1_R2337_U137, P1_R2337_U138, P1_R2337_U139, P1_R2337_U14, P1_R2337_U140, P1_R2337_U141, P1_R2337_U142, P1_R2337_U143, P1_R2337_U144, P1_R2337_U145, P1_R2337_U146, P1_R2337_U147, P1_R2337_U148, P1_R2337_U149, P1_R2337_U15, P1_R2337_U150, P1_R2337_U151, P1_R2337_U152, P1_R2337_U153, P1_R2337_U154, P1_R2337_U155, P1_R2337_U156, P1_R2337_U157, P1_R2337_U158, P1_R2337_U159, P1_R2337_U16, P1_R2337_U160, P1_R2337_U161, P1_R2337_U162, P1_R2337_U163, P1_R2337_U164, P1_R2337_U165, P1_R2337_U166, P1_R2337_U167, P1_R2337_U168, P1_R2337_U169, P1_R2337_U17, P1_R2337_U170, P1_R2337_U171, P1_R2337_U172, P1_R2337_U173, P1_R2337_U174, P1_R2337_U175, P1_R2337_U176, P1_R2337_U177, P1_R2337_U178, P1_R2337_U179, P1_R2337_U18, P1_R2337_U180, P1_R2337_U181, P1_R2337_U182, P1_R2337_U19, P1_R2337_U20, P1_R2337_U21, P1_R2337_U22, P1_R2337_U23, P1_R2337_U24, P1_R2337_U25, P1_R2337_U26, P1_R2337_U27, P1_R2337_U28, P1_R2337_U29, P1_R2337_U30, P1_R2337_U31, P1_R2337_U32, P1_R2337_U33, P1_R2337_U34, P1_R2337_U35, P1_R2337_U36, P1_R2337_U37, P1_R2337_U38, P1_R2337_U39, P1_R2337_U4, P1_R2337_U40, P1_R2337_U41, P1_R2337_U42, P1_R2337_U43, P1_R2337_U44, P1_R2337_U45, P1_R2337_U46, P1_R2337_U47, P1_R2337_U48, P1_R2337_U49, P1_R2337_U5, P1_R2337_U50, P1_R2337_U51, P1_R2337_U52, P1_R2337_U53, P1_R2337_U54, P1_R2337_U55, P1_R2337_U56, P1_R2337_U57, P1_R2337_U58, P1_R2337_U59, P1_R2337_U6, P1_R2337_U60, P1_R2337_U61, P1_R2337_U62, P1_R2337_U63, P1_R2337_U64, P1_R2337_U65, P1_R2337_U66, P1_R2337_U67, P1_R2337_U68, P1_R2337_U69, P1_R2337_U7, P1_R2337_U70, P1_R2337_U71, P1_R2337_U72, P1_R2337_U73, P1_R2337_U74, P1_R2337_U75, P1_R2337_U76, P1_R2337_U77, P1_R2337_U78, P1_R2337_U79, P1_R2337_U8, P1_R2337_U80, P1_R2337_U81, P1_R2337_U82, P1_R2337_U83, P1_R2337_U84, P1_R2337_U85, P1_R2337_U86, P1_R2337_U87, P1_R2337_U88, P1_R2337_U89, P1_R2337_U9, P1_R2337_U90, P1_R2337_U91, P1_R2337_U92, P1_R2337_U93, P1_R2337_U94, P1_R2337_U95, P1_R2337_U96, P1_R2337_U97, P1_R2337_U98, P1_R2337_U99, P1_R2358_U10, P1_R2358_U100, P1_R2358_U101, P1_R2358_U102, P1_R2358_U103, P1_R2358_U104, P1_R2358_U105, P1_R2358_U106, P1_R2358_U107, P1_R2358_U108, P1_R2358_U109, P1_R2358_U11, P1_R2358_U110, P1_R2358_U111, P1_R2358_U112, P1_R2358_U113, P1_R2358_U114, P1_R2358_U115, P1_R2358_U116, P1_R2358_U117, P1_R2358_U118, P1_R2358_U119, P1_R2358_U12, P1_R2358_U120, P1_R2358_U121, P1_R2358_U122, P1_R2358_U123, P1_R2358_U124, P1_R2358_U125, P1_R2358_U126, P1_R2358_U127, P1_R2358_U128, P1_R2358_U129, P1_R2358_U13, P1_R2358_U130, P1_R2358_U131, P1_R2358_U132, P1_R2358_U133, P1_R2358_U134, P1_R2358_U135, P1_R2358_U136, P1_R2358_U137, P1_R2358_U138, P1_R2358_U139, P1_R2358_U14, P1_R2358_U140, P1_R2358_U141, P1_R2358_U142, P1_R2358_U143, P1_R2358_U144, P1_R2358_U145, P1_R2358_U146, P1_R2358_U147, P1_R2358_U148, P1_R2358_U149, P1_R2358_U15, P1_R2358_U150, P1_R2358_U151, P1_R2358_U152, P1_R2358_U153, P1_R2358_U154, P1_R2358_U155, P1_R2358_U156, P1_R2358_U157, P1_R2358_U158, P1_R2358_U159, P1_R2358_U16, P1_R2358_U160, P1_R2358_U161, P1_R2358_U162, P1_R2358_U163, P1_R2358_U164, P1_R2358_U165, P1_R2358_U166, P1_R2358_U167, P1_R2358_U168, P1_R2358_U169, P1_R2358_U17, P1_R2358_U170, P1_R2358_U171, P1_R2358_U172, P1_R2358_U173, P1_R2358_U174, P1_R2358_U175, P1_R2358_U176, P1_R2358_U177, P1_R2358_U178, P1_R2358_U179, P1_R2358_U18, P1_R2358_U180, P1_R2358_U181, P1_R2358_U182, P1_R2358_U183, P1_R2358_U184, P1_R2358_U185, P1_R2358_U186, P1_R2358_U187, P1_R2358_U188, P1_R2358_U189, P1_R2358_U19, P1_R2358_U190, P1_R2358_U191, P1_R2358_U192, P1_R2358_U193, P1_R2358_U194, P1_R2358_U195, P1_R2358_U196, P1_R2358_U197, P1_R2358_U198, P1_R2358_U199, P1_R2358_U20, P1_R2358_U200, P1_R2358_U201, P1_R2358_U202, P1_R2358_U203, P1_R2358_U204, P1_R2358_U205, P1_R2358_U206, P1_R2358_U207, P1_R2358_U208, P1_R2358_U209, P1_R2358_U21, P1_R2358_U210, P1_R2358_U211, P1_R2358_U212, P1_R2358_U213, P1_R2358_U214, P1_R2358_U215, P1_R2358_U216, P1_R2358_U217, P1_R2358_U218, P1_R2358_U219, P1_R2358_U22, P1_R2358_U220, P1_R2358_U221, P1_R2358_U222, P1_R2358_U223, P1_R2358_U224, P1_R2358_U225, P1_R2358_U226, P1_R2358_U227, P1_R2358_U228, P1_R2358_U229, P1_R2358_U23, P1_R2358_U230, P1_R2358_U231, P1_R2358_U232, P1_R2358_U233, P1_R2358_U234, P1_R2358_U235, P1_R2358_U236, P1_R2358_U237, P1_R2358_U238, P1_R2358_U239, P1_R2358_U24, P1_R2358_U240, P1_R2358_U241, P1_R2358_U242, P1_R2358_U243, P1_R2358_U244, P1_R2358_U245, P1_R2358_U246, P1_R2358_U247, P1_R2358_U248, P1_R2358_U249, P1_R2358_U25, P1_R2358_U250, P1_R2358_U251, P1_R2358_U252, P1_R2358_U253, P1_R2358_U254, P1_R2358_U255, P1_R2358_U256, P1_R2358_U257, P1_R2358_U258, P1_R2358_U259, P1_R2358_U26, P1_R2358_U260, P1_R2358_U261, P1_R2358_U262, P1_R2358_U263, P1_R2358_U264, P1_R2358_U265, P1_R2358_U266, P1_R2358_U267, P1_R2358_U268, P1_R2358_U269, P1_R2358_U27, P1_R2358_U270, P1_R2358_U271, P1_R2358_U272, P1_R2358_U273, P1_R2358_U274, P1_R2358_U275, P1_R2358_U276, P1_R2358_U277, P1_R2358_U278, P1_R2358_U279, P1_R2358_U28, P1_R2358_U280, P1_R2358_U281, P1_R2358_U282, P1_R2358_U283, P1_R2358_U284, P1_R2358_U285, P1_R2358_U286, P1_R2358_U287, P1_R2358_U288, P1_R2358_U289, P1_R2358_U29, P1_R2358_U290, P1_R2358_U291, P1_R2358_U292, P1_R2358_U293, P1_R2358_U294, P1_R2358_U295, P1_R2358_U296, P1_R2358_U297, P1_R2358_U298, P1_R2358_U299, P1_R2358_U30, P1_R2358_U300, P1_R2358_U301, P1_R2358_U302, P1_R2358_U303, P1_R2358_U304, P1_R2358_U305, P1_R2358_U306, P1_R2358_U307, P1_R2358_U308, P1_R2358_U309, P1_R2358_U31, P1_R2358_U310, P1_R2358_U311, P1_R2358_U312, P1_R2358_U313, P1_R2358_U314, P1_R2358_U315, P1_R2358_U316, P1_R2358_U317, P1_R2358_U318, P1_R2358_U319, P1_R2358_U32, P1_R2358_U320, P1_R2358_U321, P1_R2358_U322, P1_R2358_U323, P1_R2358_U324, P1_R2358_U325, P1_R2358_U326, P1_R2358_U327, P1_R2358_U328, P1_R2358_U329, P1_R2358_U33, P1_R2358_U330, P1_R2358_U331, P1_R2358_U332, P1_R2358_U333, P1_R2358_U334, P1_R2358_U335, P1_R2358_U336, P1_R2358_U337, P1_R2358_U338, P1_R2358_U339, P1_R2358_U34, P1_R2358_U340, P1_R2358_U341, P1_R2358_U342, P1_R2358_U343, P1_R2358_U344, P1_R2358_U345, P1_R2358_U346, P1_R2358_U347, P1_R2358_U348, P1_R2358_U349, P1_R2358_U35, P1_R2358_U350, P1_R2358_U351, P1_R2358_U352, P1_R2358_U353, P1_R2358_U354, P1_R2358_U355, P1_R2358_U356, P1_R2358_U357, P1_R2358_U358, P1_R2358_U359, P1_R2358_U36, P1_R2358_U360, P1_R2358_U361, P1_R2358_U362, P1_R2358_U363, P1_R2358_U364, P1_R2358_U365, P1_R2358_U366, P1_R2358_U367, P1_R2358_U368, P1_R2358_U369, P1_R2358_U37, P1_R2358_U370, P1_R2358_U371, P1_R2358_U372, P1_R2358_U373, P1_R2358_U374, P1_R2358_U375, P1_R2358_U376, P1_R2358_U377, P1_R2358_U378, P1_R2358_U379, P1_R2358_U38, P1_R2358_U380, P1_R2358_U381, P1_R2358_U382, P1_R2358_U383, P1_R2358_U384, P1_R2358_U385, P1_R2358_U386, P1_R2358_U387, P1_R2358_U388, P1_R2358_U389, P1_R2358_U39, P1_R2358_U390, P1_R2358_U391, P1_R2358_U392, P1_R2358_U393, P1_R2358_U394, P1_R2358_U395, P1_R2358_U396, P1_R2358_U397, P1_R2358_U398, P1_R2358_U399, P1_R2358_U40, P1_R2358_U400, P1_R2358_U401, P1_R2358_U402, P1_R2358_U403, P1_R2358_U404, P1_R2358_U405, P1_R2358_U406, P1_R2358_U407, P1_R2358_U408, P1_R2358_U409, P1_R2358_U41, P1_R2358_U410, P1_R2358_U411, P1_R2358_U412, P1_R2358_U413, P1_R2358_U414, P1_R2358_U415, P1_R2358_U416, P1_R2358_U417, P1_R2358_U418, P1_R2358_U419, P1_R2358_U42, P1_R2358_U420, P1_R2358_U421, P1_R2358_U422, P1_R2358_U423, P1_R2358_U424, P1_R2358_U425, P1_R2358_U426, P1_R2358_U427, P1_R2358_U428, P1_R2358_U429, P1_R2358_U43, P1_R2358_U430, P1_R2358_U431, P1_R2358_U432, P1_R2358_U433, P1_R2358_U434, P1_R2358_U435, P1_R2358_U436, P1_R2358_U437, P1_R2358_U438, P1_R2358_U439, P1_R2358_U44, P1_R2358_U440, P1_R2358_U441, P1_R2358_U442, P1_R2358_U443, P1_R2358_U444, P1_R2358_U445, P1_R2358_U446, P1_R2358_U447, P1_R2358_U448, P1_R2358_U449, P1_R2358_U45, P1_R2358_U450, P1_R2358_U451, P1_R2358_U452, P1_R2358_U453, P1_R2358_U454, P1_R2358_U455, P1_R2358_U456, P1_R2358_U457, P1_R2358_U458, P1_R2358_U459, P1_R2358_U46, P1_R2358_U460, P1_R2358_U461, P1_R2358_U462, P1_R2358_U463, P1_R2358_U464, P1_R2358_U465, P1_R2358_U466, P1_R2358_U467, P1_R2358_U468, P1_R2358_U469, P1_R2358_U47, P1_R2358_U470, P1_R2358_U471, P1_R2358_U472, P1_R2358_U473, P1_R2358_U474, P1_R2358_U475, P1_R2358_U476, P1_R2358_U477, P1_R2358_U478, P1_R2358_U479, P1_R2358_U48, P1_R2358_U480, P1_R2358_U481, P1_R2358_U482, P1_R2358_U483, P1_R2358_U484, P1_R2358_U485, P1_R2358_U486, P1_R2358_U487, P1_R2358_U488, P1_R2358_U489, P1_R2358_U49, P1_R2358_U490, P1_R2358_U491, P1_R2358_U492, P1_R2358_U493, P1_R2358_U494, P1_R2358_U495, P1_R2358_U496, P1_R2358_U497, P1_R2358_U498, P1_R2358_U499, P1_R2358_U5, P1_R2358_U50, P1_R2358_U500, P1_R2358_U501, P1_R2358_U502, P1_R2358_U503, P1_R2358_U504, P1_R2358_U505, P1_R2358_U506, P1_R2358_U507, P1_R2358_U508, P1_R2358_U509, P1_R2358_U51, P1_R2358_U510, P1_R2358_U511, P1_R2358_U512, P1_R2358_U513, P1_R2358_U514, P1_R2358_U515, P1_R2358_U516, P1_R2358_U517, P1_R2358_U518, P1_R2358_U519, P1_R2358_U52, P1_R2358_U520, P1_R2358_U521, P1_R2358_U522, P1_R2358_U523, P1_R2358_U524, P1_R2358_U525, P1_R2358_U526, P1_R2358_U527, P1_R2358_U528, P1_R2358_U529, P1_R2358_U53, P1_R2358_U530, P1_R2358_U531, P1_R2358_U532, P1_R2358_U533, P1_R2358_U534, P1_R2358_U535, P1_R2358_U536, P1_R2358_U537, P1_R2358_U538, P1_R2358_U539, P1_R2358_U54, P1_R2358_U540, P1_R2358_U541, P1_R2358_U542, P1_R2358_U543, P1_R2358_U544, P1_R2358_U545, P1_R2358_U546, P1_R2358_U547, P1_R2358_U548, P1_R2358_U549, P1_R2358_U55, P1_R2358_U550, P1_R2358_U551, P1_R2358_U552, P1_R2358_U553, P1_R2358_U554, P1_R2358_U555, P1_R2358_U556, P1_R2358_U557, P1_R2358_U558, P1_R2358_U559, P1_R2358_U56, P1_R2358_U560, P1_R2358_U561, P1_R2358_U562, P1_R2358_U563, P1_R2358_U564, P1_R2358_U565, P1_R2358_U566, P1_R2358_U567, P1_R2358_U568, P1_R2358_U569, P1_R2358_U57, P1_R2358_U570, P1_R2358_U571, P1_R2358_U572, P1_R2358_U573, P1_R2358_U574, P1_R2358_U575, P1_R2358_U576, P1_R2358_U577, P1_R2358_U578, P1_R2358_U579, P1_R2358_U58, P1_R2358_U580, P1_R2358_U581, P1_R2358_U582, P1_R2358_U583, P1_R2358_U584, P1_R2358_U585, P1_R2358_U586, P1_R2358_U587, P1_R2358_U588, P1_R2358_U589, P1_R2358_U59, P1_R2358_U590, P1_R2358_U591, P1_R2358_U592, P1_R2358_U593, P1_R2358_U594, P1_R2358_U595, P1_R2358_U596, P1_R2358_U597, P1_R2358_U598, P1_R2358_U599, P1_R2358_U6, P1_R2358_U60, P1_R2358_U600, P1_R2358_U601, P1_R2358_U602, P1_R2358_U603, P1_R2358_U604, P1_R2358_U605, P1_R2358_U606, P1_R2358_U607, P1_R2358_U608, P1_R2358_U609, P1_R2358_U61, P1_R2358_U610, P1_R2358_U611, P1_R2358_U62, P1_R2358_U63, P1_R2358_U64, P1_R2358_U65, P1_R2358_U66, P1_R2358_U67, P1_R2358_U68, P1_R2358_U69, P1_R2358_U7, P1_R2358_U70, P1_R2358_U71, P1_R2358_U72, P1_R2358_U73, P1_R2358_U74, P1_R2358_U75, P1_R2358_U76, P1_R2358_U77, P1_R2358_U78, P1_R2358_U79, P1_R2358_U8, P1_R2358_U80, P1_R2358_U81, P1_R2358_U82, P1_R2358_U83, P1_R2358_U84, P1_R2358_U85, P1_R2358_U86, P1_R2358_U87, P1_R2358_U88, P1_R2358_U89, P1_R2358_U9, P1_R2358_U90, P1_R2358_U91, P1_R2358_U92, P1_R2358_U93, P1_R2358_U94, P1_R2358_U95, P1_R2358_U96, P1_R2358_U97, P1_R2358_U98, P1_R2358_U99, P1_R584_U6, P1_R584_U7, P1_R584_U8, P1_R584_U9, P1_SUB_357_U10, P1_SUB_357_U11, P1_SUB_357_U12, P1_SUB_357_U13, P1_SUB_357_U6, P1_SUB_357_U7, P1_SUB_357_U8, P1_SUB_357_U9, P1_SUB_450_U10, P1_SUB_450_U11, P1_SUB_450_U12, P1_SUB_450_U13, P1_SUB_450_U14, P1_SUB_450_U15, P1_SUB_450_U16, P1_SUB_450_U17, P1_SUB_450_U18, P1_SUB_450_U19, P1_SUB_450_U20, P1_SUB_450_U21, P1_SUB_450_U22, P1_SUB_450_U23, P1_SUB_450_U24, P1_SUB_450_U25, P1_SUB_450_U26, P1_SUB_450_U27, P1_SUB_450_U28, P1_SUB_450_U29, P1_SUB_450_U30, P1_SUB_450_U31, P1_SUB_450_U32, P1_SUB_450_U33, P1_SUB_450_U34, P1_SUB_450_U35, P1_SUB_450_U36, P1_SUB_450_U37, P1_SUB_450_U38, P1_SUB_450_U39, P1_SUB_450_U40, P1_SUB_450_U41, P1_SUB_450_U42, P1_SUB_450_U43, P1_SUB_450_U44, P1_SUB_450_U45, P1_SUB_450_U46, P1_SUB_450_U47, P1_SUB_450_U48, P1_SUB_450_U49, P1_SUB_450_U50, P1_SUB_450_U51, P1_SUB_450_U52, P1_SUB_450_U53, P1_SUB_450_U54, P1_SUB_450_U55, P1_SUB_450_U56, P1_SUB_450_U57, P1_SUB_450_U58, P1_SUB_450_U59, P1_SUB_450_U6, P1_SUB_450_U60, P1_SUB_450_U61, P1_SUB_450_U62, P1_SUB_450_U63, P1_SUB_450_U64, P1_SUB_450_U65, P1_SUB_450_U66, P1_SUB_450_U7, P1_SUB_450_U8, P1_SUB_450_U9, P1_SUB_580_U10, P1_SUB_580_U6, P1_SUB_580_U7, P1_SUB_580_U8, P1_SUB_580_U9, P1_U2352, P1_U2353, P1_U2354, P1_U2355, P1_U2356, P1_U2357, P1_U2358, P1_U2359, P1_U2360, P1_U2361, P1_U2362, P1_U2363, P1_U2364, P1_U2365, P1_U2366, P1_U2367, P1_U2368, P1_U2369, P1_U2370, P1_U2371, P1_U2372, P1_U2373, P1_U2374, P1_U2375, P1_U2376, P1_U2377, P1_U2378, P1_U2379, P1_U2380, P1_U2381, P1_U2382, P1_U2383, P1_U2384, P1_U2385, P1_U2386, P1_U2387, P1_U2388, P1_U2389, P1_U2390, P1_U2391, P1_U2392, P1_U2393, P1_U2394, P1_U2395, P1_U2396, P1_U2397, P1_U2398, P1_U2399, P1_U2400, P1_U2401, P1_U2402, P1_U2403, P1_U2404, P1_U2405, P1_U2406, P1_U2407, P1_U2408, P1_U2409, P1_U2410, P1_U2411, P1_U2412, P1_U2413, P1_U2414, P1_U2415, P1_U2416, P1_U2417, P1_U2418, P1_U2419, P1_U2420, P1_U2421, P1_U2422, P1_U2423, P1_U2424, P1_U2425, P1_U2426, P1_U2427, P1_U2428, P1_U2429, P1_U2430, P1_U2431, P1_U2432, P1_U2433, P1_U2434, P1_U2435, P1_U2436, P1_U2437, P1_U2438, P1_U2439, P1_U2440, P1_U2441, P1_U2442, P1_U2443, P1_U2444, P1_U2445, P1_U2446, P1_U2447, P1_U2448, P1_U2449, P1_U2450, P1_U2451, P1_U2452, P1_U2453, P1_U2454, P1_U2455, P1_U2456, P1_U2457, P1_U2458, P1_U2459, P1_U2460, P1_U2461, P1_U2462, P1_U2463, P1_U2464, P1_U2465, P1_U2466, P1_U2467, P1_U2468, P1_U2469, P1_U2470, P1_U2471, P1_U2472, P1_U2473, P1_U2474, P1_U2475, P1_U2476, P1_U2477, P1_U2478, P1_U2479, P1_U2480, P1_U2481, P1_U2482, P1_U2483, P1_U2484, P1_U2485, P1_U2486, P1_U2487, P1_U2488, P1_U2489, P1_U2490, P1_U2491, P1_U2492, P1_U2493, P1_U2494, P1_U2495, P1_U2496, P1_U2497, P1_U2498, P1_U2499, P1_U2500, P1_U2501, P1_U2502, P1_U2503, P1_U2504, P1_U2505, P1_U2506, P1_U2507, P1_U2508, P1_U2509, P1_U2510, P1_U2511, P1_U2512, P1_U2513, P1_U2514, P1_U2515, P1_U2516, P1_U2517, P1_U2518, P1_U2519, P1_U2520, P1_U2521, P1_U2522, P1_U2523, P1_U2524, P1_U2525, P1_U2526, P1_U2527, P1_U2528, P1_U2529, P1_U2530, P1_U2531, P1_U2532, P1_U2533, P1_U2534, P1_U2535, P1_U2536, P1_U2537, P1_U2538, P1_U2539, P1_U2540, P1_U2541, P1_U2542, P1_U2543, P1_U2544, P1_U2545, P1_U2546, P1_U2547, P1_U2548, P1_U2549, P1_U2550, P1_U2551, P1_U2552, P1_U2553, P1_U2554, P1_U2555, P1_U2556, P1_U2557, P1_U2558, P1_U2559, P1_U2560, P1_U2561, P1_U2562, P1_U2563, P1_U2564, P1_U2565, P1_U2566, P1_U2567, P1_U2568, P1_U2569, P1_U2570, P1_U2571, P1_U2572, P1_U2573, P1_U2574, P1_U2575, P1_U2576, P1_U2577, P1_U2578, P1_U2579, P1_U2580, P1_U2581, P1_U2582, P1_U2583, P1_U2584, P1_U2585, P1_U2586, P1_U2587, P1_U2588, P1_U2589, P1_U2590, P1_U2591, P1_U2592, P1_U2593, P1_U2594, P1_U2595, P1_U2596, P1_U2597, P1_U2598, P1_U2599, P1_U2600, P1_U2601, P1_U2602, P1_U2603, P1_U2604, P1_U2605, P1_U2606, P1_U2607, P1_U2608, P1_U2609, P1_U2610, P1_U2611, P1_U2612, P1_U2613, P1_U2614, P1_U2615, P1_U2616, P1_U2617, P1_U2618, P1_U2620, P1_U2621, P1_U2622, P1_U2623, P1_U2624, P1_U2625, P1_U2626, P1_U2627, P1_U2628, P1_U2629, P1_U2630, P1_U2631, P1_U2632, P1_U2633, P1_U2634, P1_U2635, P1_U2636, P1_U2637, P1_U2638, P1_U2639, P1_U2640, P1_U2641, P1_U2642, P1_U2643, P1_U2644, P1_U2645, P1_U2646, P1_U2647, P1_U2648, P1_U2649, P1_U2650, P1_U2651, P1_U2652, P1_U2653, P1_U2654, P1_U2655, P1_U2656, P1_U2657, P1_U2658, P1_U2659, P1_U2660, P1_U2661, P1_U2662, P1_U2663, P1_U2664, P1_U2665, P1_U2666, P1_U2667, P1_U2668, P1_U2669, P1_U2670, P1_U2671, P1_U2672, P1_U2673, P1_U2674, P1_U2675, P1_U2676, P1_U2677, P1_U2678, P1_U2679, P1_U2680, P1_U2681, P1_U2682, P1_U2683, P1_U2684, P1_U2685, P1_U2686, P1_U2687, P1_U2688, P1_U2689, P1_U2690, P1_U2691, P1_U2692, P1_U2693, P1_U2694, P1_U2695, P1_U2696, P1_U2697, P1_U2698, P1_U2699, P1_U2700, P1_U2701, P1_U2702, P1_U2703, P1_U2704, P1_U2705, P1_U2706, P1_U2707, P1_U2708, P1_U2709, P1_U2710, P1_U2711, P1_U2712, P1_U2713, P1_U2714, P1_U2715, P1_U2716, P1_U2717, P1_U2718, P1_U2719, P1_U2720, P1_U2721, P1_U2722, P1_U2723, P1_U2724, P1_U2725, P1_U2726, P1_U2727, P1_U2728, P1_U2729, P1_U2730, P1_U2731, P1_U2732, P1_U2733, P1_U2734, P1_U2735, P1_U2736, P1_U2737, P1_U2738, P1_U2739, P1_U2740, P1_U2741, P1_U2742, P1_U2743, P1_U2744, P1_U2745, P1_U2746, P1_U2747, P1_U2748, P1_U2749, P1_U2750, P1_U2751, P1_U2752, P1_U2753, P1_U2754, P1_U2755, P1_U2756, P1_U2757, P1_U2758, P1_U2759, P1_U2760, P1_U2761, P1_U2762, P1_U2763, P1_U2764, P1_U2765, P1_U2766, P1_U2767, P1_U2768, P1_U2769, P1_U2770, P1_U2771, P1_U2772, P1_U2773, P1_U2774, P1_U2775, P1_U2776, P1_U2777, P1_U2778, P1_U2779, P1_U2780, P1_U2781, P1_U2782, P1_U2783, P1_U2784, P1_U2785, P1_U2786, P1_U2787, P1_U2788, P1_U2789, P1_U2790, P1_U2791, P1_U2792, P1_U2793, P1_U2794, P1_U2795, P1_U2796, P1_U2797, P1_U2798, P1_U2799, P1_U2800, P1_U3227, P1_U3228, P1_U3229, P1_U3230, P1_U3231, P1_U3232, P1_U3233, P1_U3234, P1_U3235, P1_U3236, P1_U3237, P1_U3238, P1_U3239, P1_U3240, P1_U3241, P1_U3242, P1_U3243, P1_U3244, P1_U3245, P1_U3246, P1_U3247, P1_U3248, P1_U3249, P1_U3250, P1_U3251, P1_U3252, P1_U3253, P1_U3254, P1_U3255, P1_U3256, P1_U3257, P1_U3258, P1_U3259, P1_U3260, P1_U3261, P1_U3262, P1_U3263, P1_U3264, P1_U3265, P1_U3266, P1_U3267, P1_U3268, P1_U3269, P1_U3270, P1_U3271, P1_U3272, P1_U3273, P1_U3274, P1_U3275, P1_U3276, P1_U3277, P1_U3278, P1_U3279, P1_U3280, P1_U3281, P1_U3282, P1_U3283, P1_U3284, P1_U3285, P1_U3286, P1_U3287, P1_U3288, P1_U3289, P1_U3290, P1_U3291, P1_U3292, P1_U3293, P1_U3294, P1_U3295, P1_U3296, P1_U3297, P1_U3298, P1_U3299, P1_U3300, P1_U3301, P1_U3302, P1_U3303, P1_U3304, P1_U3305, P1_U3306, P1_U3307, P1_U3308, P1_U3309, P1_U3310, P1_U3311, P1_U3312, P1_U3313, P1_U3314, P1_U3315, P1_U3316, P1_U3317, P1_U3318, P1_U3319, P1_U3320, P1_U3321, P1_U3322, P1_U3323, P1_U3324, P1_U3325, P1_U3326, P1_U3327, P1_U3328, P1_U3329, P1_U3330, P1_U3331, P1_U3332, P1_U3333, P1_U3334, P1_U3335, P1_U3336, P1_U3337, P1_U3338, P1_U3339, P1_U3340, P1_U3341, P1_U3342, P1_U3343, P1_U3344, P1_U3345, P1_U3346, P1_U3347, P1_U3348, P1_U3349, P1_U3350, P1_U3351, P1_U3352, P1_U3353, P1_U3354, P1_U3355, P1_U3356, P1_U3357, P1_U3358, P1_U3359, P1_U3360, P1_U3361, P1_U3362, P1_U3363, P1_U3364, P1_U3365, P1_U3366, P1_U3367, P1_U3368, P1_U3369, P1_U3370, P1_U3371, P1_U3372, P1_U3373, P1_U3374, P1_U3375, P1_U3376, P1_U3377, P1_U3378, P1_U3379, P1_U3380, P1_U3381, P1_U3382, P1_U3383, P1_U3384, P1_U3385, P1_U3386, P1_U3387, P1_U3388, P1_U3389, P1_U3390, P1_U3391, P1_U3392, P1_U3393, P1_U3394, P1_U3395, P1_U3396, P1_U3397, P1_U3398, P1_U3399, P1_U3400, P1_U3401, P1_U3402, P1_U3403, P1_U3404, P1_U3405, P1_U3406, P1_U3407, P1_U3408, P1_U3409, P1_U3410, P1_U3411, P1_U3412, P1_U3413, P1_U3414, P1_U3415, P1_U3416, P1_U3417, P1_U3418, P1_U3419, P1_U3420, P1_U3421, P1_U3422, P1_U3423, P1_U3424, P1_U3425, P1_U3426, P1_U3427, P1_U3428, P1_U3429, P1_U3430, P1_U3431, P1_U3432, P1_U3433, P1_U3434, P1_U3435, P1_U3436, P1_U3437, P1_U3438, P1_U3439, P1_U3440, P1_U3441, P1_U3442, P1_U3443, P1_U3444, P1_U3445, P1_U3446, P1_U3447, P1_U3448, P1_U3449, P1_U3450, P1_U3451, P1_U3452, P1_U3453, P1_U3454, P1_U3455, P1_U3456, P1_U3457, P1_U3462, P1_U3463, P1_U3467, P1_U3470, P1_U3471, P1_U3479, P1_U3480, P1_U3488, P1_U3489, P1_U3490, P1_U3491, P1_U3492, P1_U3493, P1_U3494, P1_U3495, P1_U3496, P1_U3497, P1_U3498, P1_U3499, P1_U3500, P1_U3501, P1_U3502, P1_U3503, P1_U3504, P1_U3505, P1_U3506, P1_U3507, P1_U3508, P1_U3509, P1_U3510, P1_U3511, P1_U3512, P1_U3513, P1_U3514, P1_U3515, P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521, P1_U3522, P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528, P1_U3529, P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535, P1_U3536, P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542, P1_U3543, P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549, P1_U3550, P1_U3551, P1_U3552, P1_U3553, P1_U3554, P1_U3555, P1_U3556, P1_U3557, P1_U3558, P1_U3559, P1_U3560, P1_U3561, P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567, P1_U3568, P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574, P1_U3575, P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581, P1_U3582, P1_U3583, P1_U3584, P1_U3585, P1_U3586, P1_U3587, P1_U3588, P1_U3589, P1_U3590, P1_U3591, P1_U3592, P1_U3593, P1_U3594, P1_U3595, P1_U3596, P1_U3597, P1_U3598, P1_U3599, P1_U3600, P1_U3601, P1_U3602, P1_U3603, P1_U3604, P1_U3605, P1_U3606, P1_U3607, P1_U3608, P1_U3609, P1_U3610, P1_U3611, P1_U3612, P1_U3613, P1_U3614, P1_U3615, P1_U3616, P1_U3617, P1_U3618, P1_U3619, P1_U3620, P1_U3621, P1_U3622, P1_U3623, P1_U3624, P1_U3625, P1_U3626, P1_U3627, P1_U3628, P1_U3629, P1_U3630, P1_U3631, P1_U3632, P1_U3633, P1_U3634, P1_U3635, P1_U3636, P1_U3637, P1_U3638, P1_U3639, P1_U3640, P1_U3641, P1_U3642, P1_U3643, P1_U3644, P1_U3645, P1_U3646, P1_U3647, P1_U3648, P1_U3649, P1_U3650, P1_U3651, P1_U3652, P1_U3653, P1_U3654, P1_U3655, P1_U3656, P1_U3657, P1_U3658, P1_U3659, P1_U3660, P1_U3661, P1_U3662, P1_U3663, P1_U3664, P1_U3665, P1_U3666, P1_U3667, P1_U3668, P1_U3669, P1_U3670, P1_U3671, P1_U3672, P1_U3673, P1_U3674, P1_U3675, P1_U3676, P1_U3677, P1_U3678, P1_U3679, P1_U3680, P1_U3681, P1_U3682, P1_U3683, P1_U3684, P1_U3685, P1_U3686, P1_U3687, P1_U3688, P1_U3689, P1_U3690, P1_U3691, P1_U3692, P1_U3693, P1_U3694, P1_U3695, P1_U3696, P1_U3697, P1_U3698, P1_U3699, P1_U3700, P1_U3701, P1_U3702, P1_U3703, P1_U3704, P1_U3705, P1_U3706, P1_U3707, P1_U3708, P1_U3709, P1_U3710, P1_U3711, P1_U3712, P1_U3713, P1_U3714, P1_U3715, P1_U3716, P1_U3717, P1_U3718, P1_U3719, P1_U3720, P1_U3721, P1_U3722, P1_U3723, P1_U3724, P1_U3725, P1_U3726, P1_U3727, P1_U3728, P1_U3729, P1_U3730, P1_U3731, P1_U3732, P1_U3733, P1_U3734, P1_U3735, P1_U3736, P1_U3737, P1_U3738, P1_U3739, P1_U3740, P1_U3741, P1_U3742, P1_U3743, P1_U3744, P1_U3745, P1_U3746, P1_U3747, P1_U3748, P1_U3749, P1_U3750, P1_U3751, P1_U3752, P1_U3753, P1_U3754, P1_U3755, P1_U3756, P1_U3757, P1_U3758, P1_U3759, P1_U3760, P1_U3761, P1_U3762, P1_U3763, P1_U3764, P1_U3765, P1_U3766, P1_U3767, P1_U3768, P1_U3769, P1_U3770, P1_U3771, P1_U3772, P1_U3773, P1_U3774, P1_U3775, P1_U3776, P1_U3777, P1_U3778, P1_U3779, P1_U3780, P1_U3781, P1_U3782, P1_U3783, P1_U3784, P1_U3785, P1_U3786, P1_U3787, P1_U3788, P1_U3789, P1_U3790, P1_U3791, P1_U3792, P1_U3793, P1_U3794, P1_U3795, P1_U3796, P1_U3797, P1_U3798, P1_U3799, P1_U3800, P1_U3801, P1_U3802, P1_U3803, P1_U3804, P1_U3805, P1_U3806, P1_U3807, P1_U3808, P1_U3809, P1_U3810, P1_U3811, P1_U3812, P1_U3813, P1_U3814, P1_U3815, P1_U3816, P1_U3817, P1_U3818, P1_U3819, P1_U3820, P1_U3821, P1_U3822, P1_U3823, P1_U3824, P1_U3825, P1_U3826, P1_U3827, P1_U3828, P1_U3829, P1_U3830, P1_U3831, P1_U3832, P1_U3833, P1_U3834, P1_U3835, P1_U3836, P1_U3837, P1_U3838, P1_U3839, P1_U3840, P1_U3841, P1_U3842, P1_U3843, P1_U3844, P1_U3845, P1_U3846, P1_U3847, P1_U3848, P1_U3849, P1_U3850, P1_U3851, P1_U3852, P1_U3853, P1_U3854, P1_U3855, P1_U3856, P1_U3857, P1_U3858, P1_U3859, P1_U3860, P1_U3861, P1_U3862, P1_U3863, P1_U3864, P1_U3865, P1_U3866, P1_U3867, P1_U3868, P1_U3869, P1_U3870, P1_U3871, P1_U3872, P1_U3873, P1_U3874, P1_U3875, P1_U3876, P1_U3877, P1_U3878, P1_U3879, P1_U3880, P1_U3881, P1_U3882, P1_U3883, P1_U3884, P1_U3885, P1_U3886, P1_U3887, P1_U3888, P1_U3889, P1_U3890, P1_U3891, P1_U3892, P1_U3893, P1_U3894, P1_U3895, P1_U3896, P1_U3897, P1_U3898, P1_U3899, P1_U3900, P1_U3901, P1_U3902, P1_U3903, P1_U3904, P1_U3905, P1_U3906, P1_U3907, P1_U3908, P1_U3909, P1_U3910, P1_U3911, P1_U3912, P1_U3913, P1_U3914, P1_U3915, P1_U3916, P1_U3917, P1_U3918, P1_U3919, P1_U3920, P1_U3921, P1_U3922, P1_U3923, P1_U3924, P1_U3925, P1_U3926, P1_U3927, P1_U3928, P1_U3929, P1_U3930, P1_U3931, P1_U3932, P1_U3933, P1_U3934, P1_U3935, P1_U3936, P1_U3937, P1_U3938, P1_U3939, P1_U3940, P1_U3941, P1_U3942, P1_U3943, P1_U3944, P1_U3945, P1_U3946, P1_U3947, P1_U3948, P1_U3949, P1_U3950, P1_U3951, P1_U3952, P1_U3953, P1_U3954, P1_U3955, P1_U3956, P1_U3957, P1_U3958, P1_U3959, P1_U3960, P1_U3961, P1_U3962, P1_U3963, P1_U3964, P1_U3965, P1_U3966, P1_U3967, P1_U3968, P1_U3969, P1_U3970, P1_U3971, P1_U3972, P1_U3973, P1_U3974, P1_U3975, P1_U3976, P1_U3977, P1_U3978, P1_U3979, P1_U3980, P1_U3981, P1_U3982, P1_U3983, P1_U3984, P1_U3985, P1_U3986, P1_U3987, P1_U3988, P1_U3989, P1_U3990, P1_U3991, P1_U3992, P1_U3993, P1_U3994, P1_U3995, P1_U3996, P1_U3997, P1_U3998, P1_U3999, P1_U4000, P1_U4001, P1_U4002, P1_U4003, P1_U4004, P1_U4005, P1_U4006, P1_U4007, P1_U4008, P1_U4009, P1_U4010, P1_U4011, P1_U4012, P1_U4013, P1_U4014, P1_U4015, P1_U4016, P1_U4017, P1_U4018, P1_U4019, P1_U4020, P1_U4021, P1_U4022, P1_U4023, P1_U4024, P1_U4025, P1_U4026, P1_U4027, P1_U4028, P1_U4029, P1_U4030, P1_U4031, P1_U4032, P1_U4033, P1_U4034, P1_U4035, P1_U4036, P1_U4037, P1_U4038, P1_U4039, P1_U4040, P1_U4041, P1_U4042, P1_U4043, P1_U4044, P1_U4045, P1_U4046, P1_U4047, P1_U4048, P1_U4049, P1_U4050, P1_U4051, P1_U4052, P1_U4053, P1_U4054, P1_U4055, P1_U4056, P1_U4057, P1_U4058, P1_U4059, P1_U4060, P1_U4061, P1_U4062, P1_U4063, P1_U4064, P1_U4065, P1_U4066, P1_U4067, P1_U4068, P1_U4069, P1_U4070, P1_U4071, P1_U4072, P1_U4073, P1_U4074, P1_U4075, P1_U4076, P1_U4077, P1_U4078, P1_U4079, P1_U4080, P1_U4081, P1_U4082, P1_U4083, P1_U4084, P1_U4085, P1_U4086, P1_U4087, P1_U4088, P1_U4089, P1_U4090, P1_U4091, P1_U4092, P1_U4093, P1_U4094, P1_U4095, P1_U4096, P1_U4097, P1_U4098, P1_U4099, P1_U4100, P1_U4101, P1_U4102, P1_U4103, P1_U4104, P1_U4105, P1_U4106, P1_U4107, P1_U4108, P1_U4109, P1_U4110, P1_U4111, P1_U4112, P1_U4113, P1_U4114, P1_U4115, P1_U4116, P1_U4117, P1_U4118, P1_U4119, P1_U4120, P1_U4121, P1_U4122, P1_U4123, P1_U4124, P1_U4125, P1_U4126, P1_U4127, P1_U4128, P1_U4129, P1_U4130, P1_U4131, P1_U4132, P1_U4133, P1_U4134, P1_U4135, P1_U4136, P1_U4137, P1_U4138, P1_U4139, P1_U4140, P1_U4141, P1_U4142, P1_U4143, P1_U4144, P1_U4145, P1_U4146, P1_U4147, P1_U4148, P1_U4149, P1_U4150, P1_U4151, P1_U4152, P1_U4153, P1_U4154, P1_U4155, P1_U4156, P1_U4157, P1_U4158, P1_U4159, P1_U4160, P1_U4161, P1_U4162, P1_U4163, P1_U4164, P1_U4165, P1_U4166, P1_U4167, P1_U4168, P1_U4169, P1_U4170, P1_U4171, P1_U4172, P1_U4173, P1_U4174, P1_U4175, P1_U4176, P1_U4177, P1_U4178, P1_U4179, P1_U4180, P1_U4181, P1_U4182, P1_U4183, P1_U4184, P1_U4185, P1_U4186, P1_U4187, P1_U4188, P1_U4189, P1_U4190, P1_U4191, P1_U4192, P1_U4193, P1_U4194, P1_U4195, P1_U4196, P1_U4197, P1_U4198, P1_U4199, P1_U4200, P1_U4201, P1_U4202, P1_U4203, P1_U4204, P1_U4205, P1_U4206, P1_U4207, P1_U4208, P1_U4209, P1_U4210, P1_U4211, P1_U4212, P1_U4213, P1_U4214, P1_U4215, P1_U4216, P1_U4217, P1_U4218, P1_U4219, P1_U4220, P1_U4221, P1_U4222, P1_U4223, P1_U4224, P1_U4225, P1_U4226, P1_U4227, P1_U4228, P1_U4229, P1_U4230, P1_U4231, P1_U4232, P1_U4233, P1_U4234, P1_U4235, P1_U4236, P1_U4237, P1_U4238, P1_U4239, P1_U4240, P1_U4241, P1_U4242, P1_U4243, P1_U4244, P1_U4245, P1_U4246, P1_U4247, P1_U4248, P1_U4249, P1_U4250, P1_U4251, P1_U4252, P1_U4253, P1_U4254, P1_U4255, P1_U4256, P1_U4257, P1_U4258, P1_U4259, P1_U4260, P1_U4261, P1_U4262, P1_U4263, P1_U4264, P1_U4265, P1_U4266, P1_U4267, P1_U4268, P1_U4269, P1_U4270, P1_U4271, P1_U4272, P1_U4273, P1_U4274, P1_U4275, P1_U4276, P1_U4277, P1_U4278, P1_U4279, P1_U4280, P1_U4281, P1_U4282, P1_U4283, P1_U4284, P1_U4285, P1_U4286, P1_U4287, P1_U4288, P1_U4289, P1_U4290, P1_U4291, P1_U4292, P1_U4293, P1_U4294, P1_U4295, P1_U4296, P1_U4297, P1_U4298, P1_U4299, P1_U4300, P1_U4301, P1_U4302, P1_U4303, P1_U4304, P1_U4305, P1_U4306, P1_U4307, P1_U4308, P1_U4309, P1_U4310, P1_U4311, P1_U4312, P1_U4313, P1_U4314, P1_U4315, P1_U4316, P1_U4317, P1_U4318, P1_U4319, P1_U4320, P1_U4321, P1_U4322, P1_U4323, P1_U4324, P1_U4325, P1_U4326, P1_U4327, P1_U4328, P1_U4329, P1_U4330, P1_U4331, P1_U4332, P1_U4333, P1_U4334, P1_U4335, P1_U4336, P1_U4337, P1_U4338, P1_U4339, P1_U4340, P1_U4341, P1_U4342, P1_U4343, P1_U4344, P1_U4345, P1_U4346, P1_U4347, P1_U4348, P1_U4349, P1_U4350, P1_U4351, P1_U4352, P1_U4353, P1_U4354, P1_U4355, P1_U4356, P1_U4357, P1_U4358, P1_U4359, P1_U4360, P1_U4361, P1_U4362, P1_U4363, P1_U4364, P1_U4365, P1_U4366, P1_U4367, P1_U4368, P1_U4369, P1_U4370, P1_U4371, P1_U4372, P1_U4373, P1_U4374, P1_U4375, P1_U4376, P1_U4377, P1_U4378, P1_U4379, P1_U4380, P1_U4381, P1_U4382, P1_U4383, P1_U4384, P1_U4385, P1_U4386, P1_U4387, P1_U4388, P1_U4389, P1_U4390, P1_U4391, P1_U4392, P1_U4393, P1_U4394, P1_U4395, P1_U4396, P1_U4397, P1_U4398, P1_U4399, P1_U4400, P1_U4401, P1_U4402, P1_U4403, P1_U4404, P1_U4405, P1_U4406, P1_U4407, P1_U4408, P1_U4409, P1_U4410, P1_U4411, P1_U4412, P1_U4413, P1_U4414, P1_U4415, P1_U4416, P1_U4417, P1_U4418, P1_U4419, P1_U4420, P1_U4421, P1_U4422, P1_U4423, P1_U4424, P1_U4425, P1_U4426, P1_U4427, P1_U4428, P1_U4429, P1_U4430, P1_U4431, P1_U4432, P1_U4433, P1_U4434, P1_U4435, P1_U4436, P1_U4437, P1_U4438, P1_U4439, P1_U4440, P1_U4441, P1_U4442, P1_U4443, P1_U4444, P1_U4445, P1_U4446, P1_U4447, P1_U4448, P1_U4449, P1_U4450, P1_U4451, P1_U4452, P1_U4453, P1_U4454, P1_U4455, P1_U4456, P1_U4457, P1_U4458, P1_U4459, P1_U4460, P1_U4461, P1_U4462, P1_U4463, P1_U4464, P1_U4465, P1_U4466, P1_U4467, P1_U4468, P1_U4469, P1_U4470, P1_U4471, P1_U4472, P1_U4473, P1_U4474, P1_U4475, P1_U4476, P1_U4477, P1_U4478, P1_U4479, P1_U4480, P1_U4481, P1_U4482, P1_U4483, P1_U4484, P1_U4485, P1_U4486, P1_U4487, P1_U4488, P1_U4489, P1_U4490, P1_U4491, P1_U4492, P1_U4493, P1_U4494, P1_U4495, P1_U4496, P1_U4497, P1_U4498, P1_U4499, P1_U4500, P1_U4501, P1_U4502, P1_U4503, P1_U4504, P1_U4505, P1_U4506, P1_U4507, P1_U4508, P1_U4509, P1_U4510, P1_U4511, P1_U4512, P1_U4513, P1_U4514, P1_U4515, P1_U4516, P1_U4517, P1_U4518, P1_U4519, P1_U4520, P1_U4521, P1_U4522, P1_U4523, P1_U4524, P1_U4525, P1_U4526, P1_U4527, P1_U4528, P1_U4529, P1_U4530, P1_U4531, P1_U4532, P1_U4533, P1_U4534, P1_U4535, P1_U4536, P1_U4537, P1_U4538, P1_U4539, P1_U4540, P1_U4541, P1_U4542, P1_U4543, P1_U4544, P1_U4545, P1_U4546, P1_U4547, P1_U4548, P1_U4549, P1_U4550, P1_U4551, P1_U4552, P1_U4553, P1_U4554, P1_U4555, P1_U4556, P1_U4557, P1_U4558, P1_U4559, P1_U4560, P1_U4561, P1_U4562, P1_U4563, P1_U4564, P1_U4565, P1_U4566, P1_U4567, P1_U4568, P1_U4569, P1_U4570, P1_U4571, P1_U4572, P1_U4573, P1_U4574, P1_U4575, P1_U4576, P1_U4577, P1_U4578, P1_U4579, P1_U4580, P1_U4581, P1_U4582, P1_U4583, P1_U4584, P1_U4585, P1_U4586, P1_U4587, P1_U4588, P1_U4589, P1_U4590, P1_U4591, P1_U4592, P1_U4593, P1_U4594, P1_U4595, P1_U4596, P1_U4597, P1_U4598, P1_U4599, P1_U4600, P1_U4601, P1_U4602, P1_U4603, P1_U4604, P1_U4605, P1_U4606, P1_U4607, P1_U4608, P1_U4609, P1_U4610, P1_U4611, P1_U4612, P1_U4613, P1_U4614, P1_U4615, P1_U4616, P1_U4617, P1_U4618, P1_U4619, P1_U4620, P1_U4621, P1_U4622, P1_U4623, P1_U4624, P1_U4625, P1_U4626, P1_U4627, P1_U4628, P1_U4629, P1_U4630, P1_U4631, P1_U4632, P1_U4633, P1_U4634, P1_U4635, P1_U4636, P1_U4637, P1_U4638, P1_U4639, P1_U4640, P1_U4641, P1_U4642, P1_U4643, P1_U4644, P1_U4645, P1_U4646, P1_U4647, P1_U4648, P1_U4649, P1_U4650, P1_U4651, P1_U4652, P1_U4653, P1_U4654, P1_U4655, P1_U4656, P1_U4657, P1_U4658, P1_U4659, P1_U4660, P1_U4661, P1_U4662, P1_U4663, P1_U4664, P1_U4665, P1_U4666, P1_U4667, P1_U4668, P1_U4669, P1_U4670, P1_U4671, P1_U4672, P1_U4673, P1_U4674, P1_U4675, P1_U4676, P1_U4677, P1_U4678, P1_U4679, P1_U4680, P1_U4681, P1_U4682, P1_U4683, P1_U4684, P1_U4685, P1_U4686, P1_U4687, P1_U4688, P1_U4689, P1_U4690, P1_U4691, P1_U4692, P1_U4693, P1_U4694, P1_U4695, P1_U4696, P1_U4697, P1_U4698, P1_U4699, P1_U4700, P1_U4701, P1_U4702, P1_U4703, P1_U4704, P1_U4705, P1_U4706, P1_U4707, P1_U4708, P1_U4709, P1_U4710, P1_U4711, P1_U4712, P1_U4713, P1_U4714, P1_U4715, P1_U4716, P1_U4717, P1_U4718, P1_U4719, P1_U4720, P1_U4721, P1_U4722, P1_U4723, P1_U4724, P1_U4725, P1_U4726, P1_U4727, P1_U4728, P1_U4729, P1_U4730, P1_U4731, P1_U4732, P1_U4733, P1_U4734, P1_U4735, P1_U4736, P1_U4737, P1_U4738, P1_U4739, P1_U4740, P1_U4741, P1_U4742, P1_U4743, P1_U4744, P1_U4745, P1_U4746, P1_U4747, P1_U4748, P1_U4749, P1_U4750, P1_U4751, P1_U4752, P1_U4753, P1_U4754, P1_U4755, P1_U4756, P1_U4757, P1_U4758, P1_U4759, P1_U4760, P1_U4761, P1_U4762, P1_U4763, P1_U4764, P1_U4765, P1_U4766, P1_U4767, P1_U4768, P1_U4769, P1_U4770, P1_U4771, P1_U4772, P1_U4773, P1_U4774, P1_U4775, P1_U4776, P1_U4777, P1_U4778, P1_U4779, P1_U4780, P1_U4781, P1_U4782, P1_U4783, P1_U4784, P1_U4785, P1_U4786, P1_U4787, P1_U4788, P1_U4789, P1_U4790, P1_U4791, P1_U4792, P1_U4793, P1_U4794, P1_U4795, P1_U4796, P1_U4797, P1_U4798, P1_U4799, P1_U4800, P1_U4801, P1_U4802, P1_U4803, P1_U4804, P1_U4805, P1_U4806, P1_U4807, P1_U4808, P1_U4809, P1_U4810, P1_U4811, P1_U4812, P1_U4813, P1_U4814, P1_U4815, P1_U4816, P1_U4817, P1_U4818, P1_U4819, P1_U4820, P1_U4821, P1_U4822, P1_U4823, P1_U4824, P1_U4825, P1_U4826, P1_U4827, P1_U4828, P1_U4829, P1_U4830, P1_U4831, P1_U4832, P1_U4833, P1_U4834, P1_U4835, P1_U4836, P1_U4837, P1_U4838, P1_U4839, P1_U4840, P1_U4841, P1_U4842, P1_U4843, P1_U4844, P1_U4845, P1_U4846, P1_U4847, P1_U4848, P1_U4849, P1_U4850, P1_U4851, P1_U4852, P1_U4853, P1_U4854, P1_U4855, P1_U4856, P1_U4857, P1_U4858, P1_U4859, P1_U4860, P1_U4861, P1_U4862, P1_U4863, P1_U4864, P1_U4865, P1_U4866, P1_U4867, P1_U4868, P1_U4869, P1_U4870, P1_U4871, P1_U4872, P1_U4873, P1_U4874, P1_U4875, P1_U4876, P1_U4877, P1_U4878, P1_U4879, P1_U4880, P1_U4881, P1_U4882, P1_U4883, P1_U4884, P1_U4885, P1_U4886, P1_U4887, P1_U4888, P1_U4889, P1_U4890, P1_U4891, P1_U4892, P1_U4893, P1_U4894, P1_U4895, P1_U4896, P1_U4897, P1_U4898, P1_U4899, P1_U4900, P1_U4901, P1_U4902, P1_U4903, P1_U4904, P1_U4905, P1_U4906, P1_U4907, P1_U4908, P1_U4909, P1_U4910, P1_U4911, P1_U4912, P1_U4913, P1_U4914, P1_U4915, P1_U4916, P1_U4917, P1_U4918, P1_U4919, P1_U4920, P1_U4921, P1_U4922, P1_U4923, P1_U4924, P1_U4925, P1_U4926, P1_U4927, P1_U4928, P1_U4929, P1_U4930, P1_U4931, P1_U4932, P1_U4933, P1_U4934, P1_U4935, P1_U4936, P1_U4937, P1_U4938, P1_U4939, P1_U4940, P1_U4941, P1_U4942, P1_U4943, P1_U4944, P1_U4945, P1_U4946, P1_U4947, P1_U4948, P1_U4949, P1_U4950, P1_U4951, P1_U4952, P1_U4953, P1_U4954, P1_U4955, P1_U4956, P1_U4957, P1_U4958, P1_U4959, P1_U4960, P1_U4961, P1_U4962, P1_U4963, P1_U4964, P1_U4965, P1_U4966, P1_U4967, P1_U4968, P1_U4969, P1_U4970, P1_U4971, P1_U4972, P1_U4973, P1_U4974, P1_U4975, P1_U4976, P1_U4977, P1_U4978, P1_U4979, P1_U4980, P1_U4981, P1_U4982, P1_U4983, P1_U4984, P1_U4985, P1_U4986, P1_U4987, P1_U4988, P1_U4989, P1_U4990, P1_U4991, P1_U4992, P1_U4993, P1_U4994, P1_U4995, P1_U4996, P1_U4997, P1_U4998, P1_U4999, P1_U5000, P1_U5001, P1_U5002, P1_U5003, P1_U5004, P1_U5005, P1_U5006, P1_U5007, P1_U5008, P1_U5009, P1_U5010, P1_U5011, P1_U5012, P1_U5013, P1_U5014, P1_U5015, P1_U5016, P1_U5017, P1_U5018, P1_U5019, P1_U5020, P1_U5021, P1_U5022, P1_U5023, P1_U5024, P1_U5025, P1_U5026, P1_U5027, P1_U5028, P1_U5029, P1_U5030, P1_U5031, P1_U5032, P1_U5033, P1_U5034, P1_U5035, P1_U5036, P1_U5037, P1_U5038, P1_U5039, P1_U5040, P1_U5041, P1_U5042, P1_U5043, P1_U5044, P1_U5045, P1_U5046, P1_U5047, P1_U5048, P1_U5049, P1_U5050, P1_U5051, P1_U5052, P1_U5053, P1_U5054, P1_U5055, P1_U5056, P1_U5057, P1_U5058, P1_U5059, P1_U5060, P1_U5061, P1_U5062, P1_U5063, P1_U5064, P1_U5065, P1_U5066, P1_U5067, P1_U5068, P1_U5069, P1_U5070, P1_U5071, P1_U5072, P1_U5073, P1_U5074, P1_U5075, P1_U5076, P1_U5077, P1_U5078, P1_U5079, P1_U5080, P1_U5081, P1_U5082, P1_U5083, P1_U5084, P1_U5085, P1_U5086, P1_U5087, P1_U5088, P1_U5089, P1_U5090, P1_U5091, P1_U5092, P1_U5093, P1_U5094, P1_U5095, P1_U5096, P1_U5097, P1_U5098, P1_U5099, P1_U5100, P1_U5101, P1_U5102, P1_U5103, P1_U5104, P1_U5105, P1_U5106, P1_U5107, P1_U5108, P1_U5109, P1_U5110, P1_U5111, P1_U5112, P1_U5113, P1_U5114, P1_U5115, P1_U5116, P1_U5117, P1_U5118, P1_U5119, P1_U5120, P1_U5121, P1_U5122, P1_U5123, P1_U5124, P1_U5125, P1_U5126, P1_U5127, P1_U5128, P1_U5129, P1_U5130, P1_U5131, P1_U5132, P1_U5133, P1_U5134, P1_U5135, P1_U5136, P1_U5137, P1_U5138, P1_U5139, P1_U5140, P1_U5141, P1_U5142, P1_U5143, P1_U5144, P1_U5145, P1_U5146, P1_U5147, P1_U5148, P1_U5149, P1_U5150, P1_U5151, P1_U5152, P1_U5153, P1_U5154, P1_U5155, P1_U5156, P1_U5157, P1_U5158, P1_U5159, P1_U5160, P1_U5161, P1_U5162, P1_U5163, P1_U5164, P1_U5165, P1_U5166, P1_U5167, P1_U5168, P1_U5169, P1_U5170, P1_U5171, P1_U5172, P1_U5173, P1_U5174, P1_U5175, P1_U5176, P1_U5177, P1_U5178, P1_U5179, P1_U5180, P1_U5181, P1_U5182, P1_U5183, P1_U5184, P1_U5185, P1_U5186, P1_U5187, P1_U5188, P1_U5189, P1_U5190, P1_U5191, P1_U5192, P1_U5193, P1_U5194, P1_U5195, P1_U5196, P1_U5197, P1_U5198, P1_U5199, P1_U5200, P1_U5201, P1_U5202, P1_U5203, P1_U5204, P1_U5205, P1_U5206, P1_U5207, P1_U5208, P1_U5209, P1_U5210, P1_U5211, P1_U5212, P1_U5213, P1_U5214, P1_U5215, P1_U5216, P1_U5217, P1_U5218, P1_U5219, P1_U5220, P1_U5221, P1_U5222, P1_U5223, P1_U5224, P1_U5225, P1_U5226, P1_U5227, P1_U5228, P1_U5229, P1_U5230, P1_U5231, P1_U5232, P1_U5233, P1_U5234, P1_U5235, P1_U5236, P1_U5237, P1_U5238, P1_U5239, P1_U5240, P1_U5241, P1_U5242, P1_U5243, P1_U5244, P1_U5245, P1_U5246, P1_U5247, P1_U5248, P1_U5249, P1_U5250, P1_U5251, P1_U5252, P1_U5253, P1_U5254, P1_U5255, P1_U5256, P1_U5257, P1_U5258, P1_U5259, P1_U5260, P1_U5261, P1_U5262, P1_U5263, P1_U5264, P1_U5265, P1_U5266, P1_U5267, P1_U5268, P1_U5269, P1_U5270, P1_U5271, P1_U5272, P1_U5273, P1_U5274, P1_U5275, P1_U5276, P1_U5277, P1_U5278, P1_U5279, P1_U5280, P1_U5281, P1_U5282, P1_U5283, P1_U5284, P1_U5285, P1_U5286, P1_U5287, P1_U5288, P1_U5289, P1_U5290, P1_U5291, P1_U5292, P1_U5293, P1_U5294, P1_U5295, P1_U5296, P1_U5297, P1_U5298, P1_U5299, P1_U5300, P1_U5301, P1_U5302, P1_U5303, P1_U5304, P1_U5305, P1_U5306, P1_U5307, P1_U5308, P1_U5309, P1_U5310, P1_U5311, P1_U5312, P1_U5313, P1_U5314, P1_U5315, P1_U5316, P1_U5317, P1_U5318, P1_U5319, P1_U5320, P1_U5321, P1_U5322, P1_U5323, P1_U5324, P1_U5325, P1_U5326, P1_U5327, P1_U5328, P1_U5329, P1_U5330, P1_U5331, P1_U5332, P1_U5333, P1_U5334, P1_U5335, P1_U5336, P1_U5337, P1_U5338, P1_U5339, P1_U5340, P1_U5341, P1_U5342, P1_U5343, P1_U5344, P1_U5345, P1_U5346, P1_U5347, P1_U5348, P1_U5349, P1_U5350, P1_U5351, P1_U5352, P1_U5353, P1_U5354, P1_U5355, P1_U5356, P1_U5357, P1_U5358, P1_U5359, P1_U5360, P1_U5361, P1_U5362, P1_U5363, P1_U5364, P1_U5365, P1_U5366, P1_U5367, P1_U5368, P1_U5369, P1_U5370, P1_U5371, P1_U5372, P1_U5373, P1_U5374, P1_U5375, P1_U5376, P1_U5377, P1_U5378, P1_U5379, P1_U5380, P1_U5381, P1_U5382, P1_U5383, P1_U5384, P1_U5385, P1_U5386, P1_U5387, P1_U5388, P1_U5389, P1_U5390, P1_U5391, P1_U5392, P1_U5393, P1_U5394, P1_U5395, P1_U5396, P1_U5397, P1_U5398, P1_U5399, P1_U5400, P1_U5401, P1_U5402, P1_U5403, P1_U5404, P1_U5405, P1_U5406, P1_U5407, P1_U5408, P1_U5409, P1_U5410, P1_U5411, P1_U5412, P1_U5413, P1_U5414, P1_U5415, P1_U5416, P1_U5417, P1_U5418, P1_U5419, P1_U5420, P1_U5421, P1_U5422, P1_U5423, P1_U5424, P1_U5425, P1_U5426, P1_U5427, P1_U5428, P1_U5429, P1_U5430, P1_U5431, P1_U5432, P1_U5433, P1_U5434, P1_U5435, P1_U5436, P1_U5437, P1_U5438, P1_U5439, P1_U5440, P1_U5441, P1_U5442, P1_U5443, P1_U5444, P1_U5445, P1_U5446, P1_U5447, P1_U5448, P1_U5449, P1_U5450, P1_U5451, P1_U5452, P1_U5453, P1_U5454, P1_U5455, P1_U5456, P1_U5457, P1_U5458, P1_U5459, P1_U5460, P1_U5461, P1_U5462, P1_U5463, P1_U5464, P1_U5465, P1_U5466, P1_U5467, P1_U5468, P1_U5469, P1_U5470, P1_U5471, P1_U5472, P1_U5473, P1_U5474, P1_U5475, P1_U5476, P1_U5477, P1_U5478, P1_U5479, P1_U5480, P1_U5481, P1_U5482, P1_U5483, P1_U5484, P1_U5485, P1_U5486, P1_U5487, P1_U5488, P1_U5489, P1_U5490, P1_U5491, P1_U5492, P1_U5493, P1_U5494, P1_U5495, P1_U5496, P1_U5497, P1_U5498, P1_U5499, P1_U5500, P1_U5501, P1_U5502, P1_U5503, P1_U5504, P1_U5505, P1_U5506, P1_U5507, P1_U5508, P1_U5509, P1_U5510, P1_U5511, P1_U5512, P1_U5513, P1_U5514, P1_U5515, P1_U5516, P1_U5517, P1_U5518, P1_U5519, P1_U5520, P1_U5521, P1_U5522, P1_U5523, P1_U5524, P1_U5525, P1_U5526, P1_U5527, P1_U5528, P1_U5529, P1_U5530, P1_U5531, P1_U5532, P1_U5533, P1_U5534, P1_U5535, P1_U5536, P1_U5537, P1_U5538, P1_U5539, P1_U5540, P1_U5541, P1_U5542, P1_U5543, P1_U5544, P1_U5545, P1_U5546, P1_U5547, P1_U5548, P1_U5549, P1_U5550, P1_U5551, P1_U5552, P1_U5553, P1_U5554, P1_U5555, P1_U5556, P1_U5557, P1_U5558, P1_U5559, P1_U5560, P1_U5561, P1_U5562, P1_U5563, P1_U5564, P1_U5565, P1_U5566, P1_U5567, P1_U5568, P1_U5569, P1_U5570, P1_U5571, P1_U5572, P1_U5573, P1_U5574, P1_U5575, P1_U5576, P1_U5577, P1_U5578, P1_U5579, P1_U5580, P1_U5581, P1_U5582, P1_U5583, P1_U5584, P1_U5585, P1_U5586, P1_U5587, P1_U5588, P1_U5589, P1_U5590, P1_U5591, P1_U5592, P1_U5593, P1_U5594, P1_U5595, P1_U5596, P1_U5597, P1_U5598, P1_U5599, P1_U5600, P1_U5601, P1_U5602, P1_U5603, P1_U5604, P1_U5605, P1_U5606, P1_U5607, P1_U5608, P1_U5609, P1_U5610, P1_U5611, P1_U5612, P1_U5613, P1_U5614, P1_U5615, P1_U5616, P1_U5617, P1_U5618, P1_U5619, P1_U5620, P1_U5621, P1_U5622, P1_U5623, P1_U5624, P1_U5625, P1_U5626, P1_U5627, P1_U5628, P1_U5629, P1_U5630, P1_U5631, P1_U5632, P1_U5633, P1_U5634, P1_U5635, P1_U5636, P1_U5637, P1_U5638, P1_U5639, P1_U5640, P1_U5641, P1_U5642, P1_U5643, P1_U5644, P1_U5645, P1_U5646, P1_U5647, P1_U5648, P1_U5649, P1_U5650, P1_U5651, P1_U5652, P1_U5653, P1_U5654, P1_U5655, P1_U5656, P1_U5657, P1_U5658, P1_U5659, P1_U5660, P1_U5661, P1_U5662, P1_U5663, P1_U5664, P1_U5665, P1_U5666, P1_U5667, P1_U5668, P1_U5669, P1_U5670, P1_U5671, P1_U5672, P1_U5673, P1_U5674, P1_U5675, P1_U5676, P1_U5677, P1_U5678, P1_U5679, P1_U5680, P1_U5681, P1_U5682, P1_U5683, P1_U5684, P1_U5685, P1_U5686, P1_U5687, P1_U5688, P1_U5689, P1_U5690, P1_U5691, P1_U5692, P1_U5693, P1_U5694, P1_U5695, P1_U5696, P1_U5697, P1_U5698, P1_U5699, P1_U5700, P1_U5701, P1_U5702, P1_U5703, P1_U5704, P1_U5705, P1_U5706, P1_U5707, P1_U5708, P1_U5709, P1_U5710, P1_U5711, P1_U5712, P1_U5713, P1_U5714, P1_U5715, P1_U5716, P1_U5717, P1_U5718, P1_U5719, P1_U5720, P1_U5721, P1_U5722, P1_U5723, P1_U5724, P1_U5725, P1_U5726, P1_U5727, P1_U5728, P1_U5729, P1_U5730, P1_U5731, P1_U5732, P1_U5733, P1_U5734, P1_U5735, P1_U5736, P1_U5737, P1_U5738, P1_U5739, P1_U5740, P1_U5741, P1_U5742, P1_U5743, P1_U5744, P1_U5745, P1_U5746, P1_U5747, P1_U5748, P1_U5749, P1_U5750, P1_U5751, P1_U5752, P1_U5753, P1_U5754, P1_U5755, P1_U5756, P1_U5757, P1_U5758, P1_U5759, P1_U5760, P1_U5761, P1_U5762, P1_U5763, P1_U5764, P1_U5765, P1_U5766, P1_U5767, P1_U5768, P1_U5769, P1_U5770, P1_U5771, P1_U5772, P1_U5773, P1_U5774, P1_U5775, P1_U5776, P1_U5777, P1_U5778, P1_U5779, P1_U5780, P1_U5781, P1_U5782, P1_U5783, P1_U5784, P1_U5785, P1_U5786, P1_U5787, P1_U5788, P1_U5789, P1_U5790, P1_U5791, P1_U5792, P1_U5793, P1_U5794, P1_U5795, P1_U5796, P1_U5797, P1_U5798, P1_U5799, P1_U5800, P1_U5801, P1_U5802, P1_U5803, P1_U5804, P1_U5805, P1_U5806, P1_U5807, P1_U5808, P1_U5809, P1_U5810, P1_U5811, P1_U5812, P1_U5813, P1_U5814, P1_U5815, P1_U5816, P1_U5817, P1_U5818, P1_U5819, P1_U5820, P1_U5821, P1_U5822, P1_U5823, P1_U5824, P1_U5825, P1_U5826, P1_U5827, P1_U5828, P1_U5829, P1_U5830, P1_U5831, P1_U5832, P1_U5833, P1_U5834, P1_U5835, P1_U5836, P1_U5837, P1_U5838, P1_U5839, P1_U5840, P1_U5841, P1_U5842, P1_U5843, P1_U5844, P1_U5845, P1_U5846, P1_U5847, P1_U5848, P1_U5849, P1_U5850, P1_U5851, P1_U5852, P1_U5853, P1_U5854, P1_U5855, P1_U5856, P1_U5857, P1_U5858, P1_U5859, P1_U5860, P1_U5861, P1_U5862, P1_U5863, P1_U5864, P1_U5865, P1_U5866, P1_U5867, P1_U5868, P1_U5869, P1_U5870, P1_U5871, P1_U5872, P1_U5873, P1_U5874, P1_U5875, P1_U5876, P1_U5877, P1_U5878, P1_U5879, P1_U5880, P1_U5881, P1_U5882, P1_U5883, P1_U5884, P1_U5885, P1_U5886, P1_U5887, P1_U5888, P1_U5889, P1_U5890, P1_U5891, P1_U5892, P1_U5893, P1_U5894, P1_U5895, P1_U5896, P1_U5897, P1_U5898, P1_U5899, P1_U5900, P1_U5901, P1_U5902, P1_U5903, P1_U5904, P1_U5905, P1_U5906, P1_U5907, P1_U5908, P1_U5909, P1_U5910, P1_U5911, P1_U5912, P1_U5913, P1_U5914, P1_U5915, P1_U5916, P1_U5917, P1_U5918, P1_U5919, P1_U5920, P1_U5921, P1_U5922, P1_U5923, P1_U5924, P1_U5925, P1_U5926, P1_U5927, P1_U5928, P1_U5929, P1_U5930, P1_U5931, P1_U5932, P1_U5933, P1_U5934, P1_U5935, P1_U5936, P1_U5937, P1_U5938, P1_U5939, P1_U5940, P1_U5941, P1_U5942, P1_U5943, P1_U5944, P1_U5945, P1_U5946, P1_U5947, P1_U5948, P1_U5949, P1_U5950, P1_U5951, P1_U5952, P1_U5953, P1_U5954, P1_U5955, P1_U5956, P1_U5957, P1_U5958, P1_U5959, P1_U5960, P1_U5961, P1_U5962, P1_U5963, P1_U5964, P1_U5965, P1_U5966, P1_U5967, P1_U5968, P1_U5969, P1_U5970, P1_U5971, P1_U5972, P1_U5973, P1_U5974, P1_U5975, P1_U5976, P1_U5977, P1_U5978, P1_U5979, P1_U5980, P1_U5981, P1_U5982, P1_U5983, P1_U5984, P1_U5985, P1_U5986, P1_U5987, P1_U5988, P1_U5989, P1_U5990, P1_U5991, P1_U5992, P1_U5993, P1_U5994, P1_U5995, P1_U5996, P1_U5997, P1_U5998, P1_U5999, P1_U6000, P1_U6001, P1_U6002, P1_U6003, P1_U6004, P1_U6005, P1_U6006, P1_U6007, P1_U6008, P1_U6009, P1_U6010, P1_U6011, P1_U6012, P1_U6013, P1_U6014, P1_U6015, P1_U6016, P1_U6017, P1_U6018, P1_U6019, P1_U6020, P1_U6021, P1_U6022, P1_U6023, P1_U6024, P1_U6025, P1_U6026, P1_U6027, P1_U6028, P1_U6029, P1_U6030, P1_U6031, P1_U6032, P1_U6033, P1_U6034, P1_U6035, P1_U6036, P1_U6037, P1_U6038, P1_U6039, P1_U6040, P1_U6041, P1_U6042, P1_U6043, P1_U6044, P1_U6045, P1_U6046, P1_U6047, P1_U6048, P1_U6049, P1_U6050, P1_U6051, P1_U6052, P1_U6053, P1_U6054, P1_U6055, P1_U6056, P1_U6057, P1_U6058, P1_U6059, P1_U6060, P1_U6061, P1_U6062, P1_U6063, P1_U6064, P1_U6065, P1_U6066, P1_U6067, P1_U6068, P1_U6069, P1_U6070, P1_U6071, P1_U6072, P1_U6073, P1_U6074, P1_U6075, P1_U6076, P1_U6077, P1_U6078, P1_U6079, P1_U6080, P1_U6081, P1_U6082, P1_U6083, P1_U6084, P1_U6085, P1_U6086, P1_U6087, P1_U6088, P1_U6089, P1_U6090, P1_U6091, P1_U6092, P1_U6093, P1_U6094, P1_U6095, P1_U6096, P1_U6097, P1_U6098, P1_U6099, P1_U6100, P1_U6101, P1_U6102, P1_U6103, P1_U6104, P1_U6105, P1_U6106, P1_U6107, P1_U6108, P1_U6109, P1_U6110, P1_U6111, P1_U6112, P1_U6113, P1_U6114, P1_U6115, P1_U6116, P1_U6117, P1_U6118, P1_U6119, P1_U6120, P1_U6121, P1_U6122, P1_U6123, P1_U6124, P1_U6125, P1_U6126, P1_U6127, P1_U6128, P1_U6129, P1_U6130, P1_U6131, P1_U6132, P1_U6133, P1_U6134, P1_U6135, P1_U6136, P1_U6137, P1_U6138, P1_U6139, P1_U6140, P1_U6141, P1_U6142, P1_U6143, P1_U6144, P1_U6145, P1_U6146, P1_U6147, P1_U6148, P1_U6149, P1_U6150, P1_U6151, P1_U6152, P1_U6153, P1_U6154, P1_U6155, P1_U6156, P1_U6157, P1_U6158, P1_U6159, P1_U6160, P1_U6161, P1_U6162, P1_U6163, P1_U6164, P1_U6165, P1_U6166, P1_U6167, P1_U6168, P1_U6169, P1_U6170, P1_U6171, P1_U6172, P1_U6173, P1_U6174, P1_U6175, P1_U6176, P1_U6177, P1_U6178, P1_U6179, P1_U6180, P1_U6181, P1_U6182, P1_U6183, P1_U6184, P1_U6185, P1_U6186, P1_U6187, P1_U6188, P1_U6189, P1_U6190, P1_U6191, P1_U6192, P1_U6193, P1_U6194, P1_U6195, P1_U6196, P1_U6197, P1_U6198, P1_U6199, P1_U6200, P1_U6201, P1_U6202, P1_U6203, P1_U6204, P1_U6205, P1_U6206, P1_U6207, P1_U6208, P1_U6209, P1_U6210, P1_U6211, P1_U6212, P1_U6213, P1_U6214, P1_U6215, P1_U6216, P1_U6217, P1_U6218, P1_U6219, P1_U6220, P1_U6221, P1_U6222, P1_U6223, P1_U6224, P1_U6225, P1_U6226, P1_U6227, P1_U6228, P1_U6229, P1_U6230, P1_U6231, P1_U6232, P1_U6233, P1_U6234, P1_U6235, P1_U6236, P1_U6237, P1_U6238, P1_U6239, P1_U6240, P1_U6241, P1_U6242, P1_U6243, P1_U6244, P1_U6245, P1_U6246, P1_U6247, P1_U6248, P1_U6249, P1_U6250, P1_U6251, P1_U6252, P1_U6253, P1_U6254, P1_U6255, P1_U6256, P1_U6257, P1_U6258, P1_U6259, P1_U6260, P1_U6261, P1_U6262, P1_U6263, P1_U6264, P1_U6265, P1_U6266, P1_U6267, P1_U6268, P1_U6269, P1_U6270, P1_U6271, P1_U6272, P1_U6273, P1_U6274, P1_U6275, P1_U6276, P1_U6277, P1_U6278, P1_U6279, P1_U6280, P1_U6281, P1_U6282, P1_U6283, P1_U6284, P1_U6285, P1_U6286, P1_U6287, P1_U6288, P1_U6289, P1_U6290, P1_U6291, P1_U6292, P1_U6293, P1_U6294, P1_U6295, P1_U6296, P1_U6297, P1_U6298, P1_U6299, P1_U6300, P1_U6301, P1_U6302, P1_U6303, P1_U6304, P1_U6305, P1_U6306, P1_U6307, P1_U6308, P1_U6309, P1_U6310, P1_U6311, P1_U6312, P1_U6313, P1_U6314, P1_U6315, P1_U6316, P1_U6317, P1_U6318, P1_U6319, P1_U6320, P1_U6321, P1_U6322, P1_U6323, P1_U6324, P1_U6325, P1_U6326, P1_U6327, P1_U6328, P1_U6329, P1_U6330, P1_U6331, P1_U6332, P1_U6333, P1_U6334, P1_U6335, P1_U6336, P1_U6337, P1_U6338, P1_U6339, P1_U6340, P1_U6341, P1_U6342, P1_U6343, P1_U6344, P1_U6345, P1_U6346, P1_U6347, P1_U6348, P1_U6349, P1_U6350, P1_U6351, P1_U6352, P1_U6353, P1_U6354, P1_U6355, P1_U6356, P1_U6357, P1_U6358, P1_U6359, P1_U6360, P1_U6361, P1_U6362, P1_U6363, P1_U6364, P1_U6365, P1_U6366, P1_U6367, P1_U6368, P1_U6369, P1_U6370, P1_U6371, P1_U6372, P1_U6373, P1_U6374, P1_U6375, P1_U6376, P1_U6377, P1_U6378, P1_U6379, P1_U6380, P1_U6381, P1_U6382, P1_U6383, P1_U6384, P1_U6385, P1_U6386, P1_U6387, P1_U6388, P1_U6389, P1_U6390, P1_U6391, P1_U6392, P1_U6393, P1_U6394, P1_U6395, P1_U6396, P1_U6397, P1_U6398, P1_U6399, P1_U6400, P1_U6401, P1_U6402, P1_U6403, P1_U6404, P1_U6405, P1_U6406, P1_U6407, P1_U6408, P1_U6409, P1_U6410, P1_U6411, P1_U6412, P1_U6413, P1_U6414, P1_U6415, P1_U6416, P1_U6417, P1_U6418, P1_U6419, P1_U6420, P1_U6421, P1_U6422, P1_U6423, P1_U6424, P1_U6425, P1_U6426, P1_U6427, P1_U6428, P1_U6429, P1_U6430, P1_U6431, P1_U6432, P1_U6433, P1_U6434, P1_U6435, P1_U6436, P1_U6437, P1_U6438, P1_U6439, P1_U6440, P1_U6441, P1_U6442, P1_U6443, P1_U6444, P1_U6445, P1_U6446, P1_U6447, P1_U6448, P1_U6449, P1_U6450, P1_U6451, P1_U6452, P1_U6453, P1_U6454, P1_U6455, P1_U6456, P1_U6457, P1_U6458, P1_U6459, P1_U6460, P1_U6461, P1_U6462, P1_U6463, P1_U6464, P1_U6465, P1_U6466, P1_U6467, P1_U6468, P1_U6469, P1_U6470, P1_U6471, P1_U6472, P1_U6473, P1_U6474, P1_U6475, P1_U6476, P1_U6477, P1_U6478, P1_U6479, P1_U6480, P1_U6481, P1_U6482, P1_U6483, P1_U6484, P1_U6485, P1_U6486, P1_U6487, P1_U6488, P1_U6489, P1_U6490, P1_U6491, P1_U6492, P1_U6493, P1_U6494, P1_U6495, P1_U6496, P1_U6497, P1_U6498, P1_U6499, P1_U6500, P1_U6501, P1_U6502, P1_U6503, P1_U6504, P1_U6505, P1_U6506, P1_U6507, P1_U6508, P1_U6509, P1_U6510, P1_U6511, P1_U6512, P1_U6513, P1_U6514, P1_U6515, P1_U6516, P1_U6517, P1_U6518, P1_U6519, P1_U6520, P1_U6521, P1_U6522, P1_U6523, P1_U6524, P1_U6525, P1_U6526, P1_U6527, P1_U6528, P1_U6529, P1_U6530, P1_U6531, P1_U6532, P1_U6533, P1_U6534, P1_U6535, P1_U6536, P1_U6537, P1_U6538, P1_U6539, P1_U6540, P1_U6541, P1_U6542, P1_U6543, P1_U6544, P1_U6545, P1_U6546, P1_U6547, P1_U6548, P1_U6549, P1_U6550, P1_U6551, P1_U6552, P1_U6553, P1_U6554, P1_U6555, P1_U6556, P1_U6557, P1_U6558, P1_U6559, P1_U6560, P1_U6561, P1_U6562, P1_U6563, P1_U6564, P1_U6565, P1_U6566, P1_U6567, P1_U6568, P1_U6569, P1_U6570, P1_U6571, P1_U6572, P1_U6573, P1_U6574, P1_U6575, P1_U6576, P1_U6577, P1_U6578, P1_U6579, P1_U6580, P1_U6581, P1_U6582, P1_U6583, P1_U6584, P1_U6585, P1_U6586, P1_U6587, P1_U6588, P1_U6589, P1_U6590, P1_U6591, P1_U6592, P1_U6593, P1_U6594, P1_U6595, P1_U6596, P1_U6597, P1_U6598, P1_U6599, P1_U6600, P1_U6601, P1_U6602, P1_U6603, P1_U6604, P1_U6605, P1_U6606, P1_U6607, P1_U6608, P1_U6609, P1_U6610, P1_U6611, P1_U6612, P1_U6613, P1_U6614, P1_U6615, P1_U6616, P1_U6617, P1_U6618, P1_U6619, P1_U6620, P1_U6621, P1_U6622, P1_U6623, P1_U6624, P1_U6625, P1_U6626, P1_U6627, P1_U6628, P1_U6629, P1_U6630, P1_U6631, P1_U6632, P1_U6633, P1_U6634, P1_U6635, P1_U6636, P1_U6637, P1_U6638, P1_U6639, P1_U6640, P1_U6641, P1_U6642, P1_U6643, P1_U6644, P1_U6645, P1_U6646, P1_U6647, P1_U6648, P1_U6649, P1_U6650, P1_U6651, P1_U6652, P1_U6653, P1_U6654, P1_U6655, P1_U6656, P1_U6657, P1_U6658, P1_U6659, P1_U6660, P1_U6661, P1_U6662, P1_U6663, P1_U6664, P1_U6665, P1_U6666, P1_U6667, P1_U6668, P1_U6669, P1_U6670, P1_U6671, P1_U6672, P1_U6673, P1_U6674, P1_U6675, P1_U6676, P1_U6677, P1_U6678, P1_U6679, P1_U6680, P1_U6681, P1_U6682, P1_U6683, P1_U6684, P1_U6685, P1_U6686, P1_U6687, P1_U6688, P1_U6689, P1_U6690, P1_U6691, P1_U6692, P1_U6693, P1_U6694, P1_U6695, P1_U6696, P1_U6697, P1_U6698, P1_U6699, P1_U6700, P1_U6701, P1_U6702, P1_U6703, P1_U6704, P1_U6705, P1_U6706, P1_U6707, P1_U6708, P1_U6709, P1_U6710, P1_U6711, P1_U6712, P1_U6713, P1_U6714, P1_U6715, P1_U6716, P1_U6717, P1_U6718, P1_U6719, P1_U6720, P1_U6721, P1_U6722, P1_U6723, P1_U6724, P1_U6725, P1_U6726, P1_U6727, P1_U6728, P1_U6729, P1_U6730, P1_U6731, P1_U6732, P1_U6733, P1_U6734, P1_U6735, P1_U6736, P1_U6737, P1_U6738, P1_U6739, P1_U6740, P1_U6741, P1_U6742, P1_U6743, P1_U6744, P1_U6745, P1_U6746, P1_U6747, P1_U6748, P1_U6749, P1_U6750, P1_U6751, P1_U6752, P1_U6753, P1_U6754, P1_U6755, P1_U6756, P1_U6757, P1_U6758, P1_U6759, P1_U6760, P1_U6761, P1_U6762, P1_U6763, P1_U6764, P1_U6765, P1_U6766, P1_U6767, P1_U6768, P1_U6769, P1_U6770, P1_U6771, P1_U6772, P1_U6773, P1_U6774, P1_U6775, P1_U6776, P1_U6777, P1_U6778, P1_U6779, P1_U6780, P1_U6781, P1_U6782, P1_U6783, P1_U6784, P1_U6785, P1_U6786, P1_U6787, P1_U6788, P1_U6789, P1_U6790, P1_U6791, P1_U6792, P1_U6793, P1_U6794, P1_U6795, P1_U6796, P1_U6797, P1_U6798, P1_U6799, P1_U6800, P1_U6801, P1_U6802, P1_U6803, P1_U6804, P1_U6805, P1_U6806, P1_U6807, P1_U6808, P1_U6809, P1_U6810, P1_U6811, P1_U6812, P1_U6813, P1_U6814, P1_U6815, P1_U6816, P1_U6817, P1_U6818, P1_U6819, P1_U6820, P1_U6821, P1_U6822, P1_U6823, P1_U6824, P1_U6825, P1_U6826, P1_U6827, P1_U6828, P1_U6829, P1_U6830, P1_U6831, P1_U6832, P1_U6833, P1_U6834, P1_U6835, P1_U6836, P1_U6837, P1_U6838, P1_U6839, P1_U6840, P1_U6841, P1_U6842, P1_U6843, P1_U6844, P1_U6845, P1_U6846, P1_U6847, P1_U6848, P1_U6849, P1_U6850, P1_U6851, P1_U6852, P1_U6853, P1_U6854, P1_U6855, P1_U6856, P1_U6857, P1_U6858, P1_U6859, P1_U6860, P1_U6861, P1_U6862, P1_U6863, P1_U6864, P1_U6865, P1_U6866, P1_U6867, P1_U6868, P1_U6869, P1_U6870, P1_U6871, P1_U6872, P1_U6873, P1_U6874, P1_U6875, P1_U6876, P1_U6877, P1_U6878, P1_U6879, P1_U6880, P1_U6881, P1_U6882, P1_U6883, P1_U6884, P1_U6885, P1_U6886, P1_U6887, P1_U6888, P1_U6889, P1_U6890, P1_U6891, P1_U6892, P1_U6893, P1_U6894, P1_U6895, P1_U6896, P1_U6897, P1_U6898, P1_U6899, P1_U6900, P1_U6901, P1_U6902, P1_U6903, P1_U6904, P1_U6905, P1_U6906, P1_U6907, P1_U6908, P1_U6909, P1_U6910, P1_U6911, P1_U6912, P1_U6913, P1_U6914, P1_U6915, P1_U6916, P1_U6917, P1_U6918, P1_U6919, P1_U6920, P1_U6921, P1_U6922, P1_U6923, P1_U6924, P1_U6925, P1_U6926, P1_U6927, P1_U6928, P1_U6929, P1_U6930, P1_U6931, P1_U6932, P1_U6933, P1_U6934, P1_U6935, P1_U6936, P1_U6937, P1_U6938, P1_U6939, P1_U6940, P1_U6941, P1_U6942, P1_U6943, P1_U6944, P1_U6945, P1_U6946, P1_U6947, P1_U6948, P1_U6949, P1_U6950, P1_U6951, P1_U6952, P1_U6953, P1_U6954, P1_U6955, P1_U6956, P1_U6957, P1_U6958, P1_U6959, P1_U6960, P1_U6961, P1_U6962, P1_U6963, P1_U6964, P1_U6965, P1_U6966, P1_U6967, P1_U6968, P1_U6969, P1_U6970, P1_U6971, P1_U6972, P1_U6973, P1_U6974, P1_U6975, P1_U6976, P1_U6977, P1_U6978, P1_U6979, P1_U6980, P1_U6981, P1_U6982, P1_U6983, P1_U6984, P1_U6985, P1_U6986, P1_U6987, P1_U6988, P1_U6989, P1_U6990, P1_U6991, P1_U6992, P1_U6993, P1_U6994, P1_U6995, P1_U6996, P1_U6997, P1_U6998, P1_U6999, P1_U7000, P1_U7001, P1_U7002, P1_U7003, P1_U7004, P1_U7005, P1_U7006, P1_U7007, P1_U7008, P1_U7009, P1_U7010, P1_U7011, P1_U7012, P1_U7013, P1_U7014, P1_U7015, P1_U7016, P1_U7017, P1_U7018, P1_U7019, P1_U7020, P1_U7021, P1_U7022, P1_U7023, P1_U7024, P1_U7025, P1_U7026, P1_U7027, P1_U7028, P1_U7029, P1_U7030, P1_U7031, P1_U7032, P1_U7033, P1_U7034, P1_U7035, P1_U7036, P1_U7037, P1_U7038, P1_U7039, P1_U7040, P1_U7041, P1_U7042, P1_U7043, P1_U7044, P1_U7045, P1_U7046, P1_U7047, P1_U7048, P1_U7049, P1_U7050, P1_U7051, P1_U7052, P1_U7053, P1_U7054, P1_U7055, P1_U7056, P1_U7057, P1_U7058, P1_U7059, P1_U7060, P1_U7061, P1_U7062, P1_U7063, P1_U7064, P1_U7065, P1_U7066, P1_U7067, P1_U7068, P1_U7069, P1_U7070, P1_U7071, P1_U7072, P1_U7073, P1_U7074, P1_U7075, P1_U7076, P1_U7077, P1_U7078, P1_U7079, P1_U7080, P1_U7081, P1_U7082, P1_U7083, P1_U7084, P1_U7085, P1_U7086, P1_U7087, P1_U7088, P1_U7089, P1_U7090, P1_U7091, P1_U7092, P1_U7093, P1_U7094, P1_U7095, P1_U7096, P1_U7097, P1_U7098, P1_U7099, P1_U7100, P1_U7101, P1_U7102, P1_U7103, P1_U7104, P1_U7105, P1_U7106, P1_U7107, P1_U7108, P1_U7109, P1_U7110, P1_U7111, P1_U7112, P1_U7113, P1_U7114, P1_U7115, P1_U7116, P1_U7117, P1_U7118, P1_U7119, P1_U7120, P1_U7121, P1_U7122, P1_U7123, P1_U7124, P1_U7125, P1_U7126, P1_U7127, P1_U7128, P1_U7129, P1_U7130, P1_U7131, P1_U7132, P1_U7133, P1_U7134, P1_U7135, P1_U7136, P1_U7137, P1_U7138, P1_U7139, P1_U7140, P1_U7141, P1_U7142, P1_U7143, P1_U7144, P1_U7145, P1_U7146, P1_U7147, P1_U7148, P1_U7149, P1_U7150, P1_U7151, P1_U7152, P1_U7153, P1_U7154, P1_U7155, P1_U7156, P1_U7157, P1_U7158, P1_U7159, P1_U7160, P1_U7161, P1_U7162, P1_U7163, P1_U7164, P1_U7165, P1_U7166, P1_U7167, P1_U7168, P1_U7169, P1_U7170, P1_U7171, P1_U7172, P1_U7173, P1_U7174, P1_U7175, P1_U7176, P1_U7177, P1_U7178, P1_U7179, P1_U7180, P1_U7181, P1_U7182, P1_U7183, P1_U7184, P1_U7185, P1_U7186, P1_U7187, P1_U7188, P1_U7189, P1_U7190, P1_U7191, P1_U7192, P1_U7193, P1_U7194, P1_U7195, P1_U7196, P1_U7197, P1_U7198, P1_U7199, P1_U7200, P1_U7201, P1_U7202, P1_U7203, P1_U7204, P1_U7205, P1_U7206, P1_U7207, P1_U7208, P1_U7209, P1_U7210, P1_U7211, P1_U7212, P1_U7213, P1_U7214, P1_U7215, P1_U7216, P1_U7217, P1_U7218, P1_U7219, P1_U7220, P1_U7221, P1_U7222, P1_U7223, P1_U7224, P1_U7225, P1_U7226, P1_U7227, P1_U7228, P1_U7229, P1_U7230, P1_U7231, P1_U7232, P1_U7233, P1_U7234, P1_U7235, P1_U7236, P1_U7237, P1_U7238, P1_U7239, P1_U7240, P1_U7241, P1_U7242, P1_U7243, P1_U7244, P1_U7245, P1_U7246, P1_U7247, P1_U7248, P1_U7249, P1_U7250, P1_U7251, P1_U7252, P1_U7253, P1_U7254, P1_U7255, P1_U7256, P1_U7257, P1_U7258, P1_U7259, P1_U7260, P1_U7261, P1_U7262, P1_U7263, P1_U7264, P1_U7265, P1_U7266, P1_U7267, P1_U7268, P1_U7269, P1_U7270, P1_U7271, P1_U7272, P1_U7273, P1_U7274, P1_U7275, P1_U7276, P1_U7277, P1_U7278, P1_U7279, P1_U7280, P1_U7281, P1_U7282, P1_U7283, P1_U7284, P1_U7285, P1_U7286, P1_U7287, P1_U7288, P1_U7289, P1_U7290, P1_U7291, P1_U7292, P1_U7293, P1_U7294, P1_U7295, P1_U7296, P1_U7297, P1_U7298, P1_U7299, P1_U7300, P1_U7301, P1_U7302, P1_U7303, P1_U7304, P1_U7305, P1_U7306, P1_U7307, P1_U7308, P1_U7309, P1_U7310, P1_U7311, P1_U7312, P1_U7313, P1_U7314, P1_U7315, P1_U7316, P1_U7317, P1_U7318, P1_U7319, P1_U7320, P1_U7321, P1_U7322, P1_U7323, P1_U7324, P1_U7325, P1_U7326, P1_U7327, P1_U7328, P1_U7329, P1_U7330, P1_U7331, P1_U7332, P1_U7333, P1_U7334, P1_U7335, P1_U7336, P1_U7337, P1_U7338, P1_U7339, P1_U7340, P1_U7341, P1_U7342, P1_U7343, P1_U7344, P1_U7345, P1_U7346, P1_U7347, P1_U7348, P1_U7349, P1_U7350, P1_U7351, P1_U7352, P1_U7353, P1_U7354, P1_U7355, P1_U7356, P1_U7357, P1_U7358, P1_U7359, P1_U7360, P1_U7361, P1_U7362, P1_U7363, P1_U7364, P1_U7365, P1_U7366, P1_U7367, P1_U7368, P1_U7369, P1_U7370, P1_U7371, P1_U7372, P1_U7373, P1_U7374, P1_U7375, P1_U7376, P1_U7377, P1_U7378, P1_U7379, P1_U7380, P1_U7381, P1_U7382, P1_U7383, P1_U7384, P1_U7385, P1_U7386, P1_U7387, P1_U7388, P1_U7389, P1_U7390, P1_U7391, P1_U7392, P1_U7393, P1_U7394, P1_U7395, P1_U7396, P1_U7397, P1_U7398, P1_U7399, P1_U7400, P1_U7401, P1_U7402, P1_U7403, P1_U7404, P1_U7405, P1_U7406, P1_U7407, P1_U7408, P1_U7409, P1_U7410, P1_U7411, P1_U7412, P1_U7413, P1_U7414, P1_U7415, P1_U7416, P1_U7417, P1_U7418, P1_U7419, P1_U7420, P1_U7421, P1_U7422, P1_U7423, P1_U7424, P1_U7425, P1_U7426, P1_U7427, P1_U7428, P1_U7429, P1_U7430, P1_U7431, P1_U7432, P1_U7433, P1_U7434, P1_U7435, P1_U7436, P1_U7437, P1_U7438, P1_U7439, P1_U7440, P1_U7441, P1_U7442, P1_U7443, P1_U7444, P1_U7445, P1_U7446, P1_U7447, P1_U7448, P1_U7449, P1_U7450, P1_U7451, P1_U7452, P1_U7453, P1_U7454, P1_U7455, P1_U7456, P1_U7457, P1_U7458, P1_U7459, P1_U7460, P1_U7461, P1_U7462, P1_U7463, P1_U7464, P1_U7465, P1_U7466, P1_U7467, P1_U7468, P1_U7469, P1_U7470, P1_U7471, P1_U7472, P1_U7473, P1_U7474, P1_U7475, P1_U7476, P1_U7477, P1_U7478, P1_U7479, P1_U7480, P1_U7481, P1_U7482, P1_U7483, P1_U7484, P1_U7485, P1_U7486, P1_U7487, P1_U7488, P1_U7489, P1_U7490, P1_U7491, P1_U7492, P1_U7493, P1_U7494, P1_U7495, P1_U7496, P1_U7497, P1_U7498, P1_U7499, P1_U7500, P1_U7501, P1_U7502, P1_U7503, P1_U7504, P1_U7505, P1_U7506, P1_U7507, P1_U7508, P1_U7509, P1_U7510, P1_U7511, P1_U7512, P1_U7513, P1_U7514, P1_U7515, P1_U7516, P1_U7517, P1_U7518, P1_U7519, P1_U7520, P1_U7521, P1_U7522, P1_U7523, P1_U7524, P1_U7525, P1_U7526, P1_U7527, P1_U7528, P1_U7529, P1_U7530, P1_U7531, P1_U7532, P1_U7533, P1_U7534, P1_U7535, P1_U7536, P1_U7537, P1_U7538, P1_U7539, P1_U7540, P1_U7541, P1_U7542, P1_U7543, P1_U7544, P1_U7545, P1_U7546, P1_U7547, P1_U7548, P1_U7549, P1_U7550, P1_U7551, P1_U7552, P1_U7553, P1_U7554, P1_U7555, P1_U7556, P1_U7557, P1_U7558, P1_U7559, P1_U7560, P1_U7561, P1_U7562, P1_U7563, P1_U7564, P1_U7565, P1_U7566, P1_U7567, P1_U7568, P1_U7569, P1_U7570, P1_U7571, P1_U7572, P1_U7573, P1_U7574, P1_U7575, P1_U7576, P1_U7577, P1_U7578, P1_U7579, P1_U7580, P1_U7581, P1_U7582, P1_U7583, P1_U7584, P1_U7585, P1_U7586, P1_U7587, P1_U7588, P1_U7589, P1_U7590, P1_U7591, P1_U7592, P1_U7593, P1_U7594, P1_U7595, P1_U7596, P1_U7597, P1_U7598, P1_U7599, P1_U7600, P1_U7601, P1_U7602, P1_U7603, P1_U7604, P1_U7605, P1_U7606, P1_U7607, P1_U7608, P1_U7609, P1_U7610, P1_U7611, P1_U7612, P1_U7613, P1_U7614, P1_U7615, P1_U7616, P1_U7617, P1_U7618, P1_U7619, P1_U7620, P1_U7621, P1_U7622, P1_U7623, P1_U7624, P1_U7625, P1_U7626, P1_U7627, P1_U7628, P1_U7629, P1_U7630, P1_U7631, P1_U7632, P1_U7633, P1_U7634, P1_U7635, P1_U7636, P1_U7637, P1_U7638, P1_U7639, P1_U7640, P1_U7641, P1_U7642, P1_U7643, P1_U7644, P1_U7645, P1_U7646, P1_U7647, P1_U7648, P1_U7649, P1_U7650, P1_U7651, P1_U7652, P1_U7653, P1_U7654, P1_U7655, P1_U7656, P1_U7657, P1_U7658, P1_U7659, P1_U7660, P1_U7661, P1_U7662, P1_U7663, P1_U7664, P1_U7665, P1_U7666, P1_U7667, P1_U7668, P1_U7669, P1_U7670, P1_U7671, P1_U7672, P1_U7673, P1_U7674, P1_U7675, P1_U7676, P1_U7677, P1_U7678, P1_U7679, P1_U7680, P1_U7681, P1_U7682, P1_U7683, P1_U7684, P1_U7685, P1_U7686, P1_U7687, P1_U7688, P1_U7689, P1_U7690, P1_U7691, P1_U7692, P1_U7693, P1_U7694, P1_U7695, P1_U7696, P1_U7697, P1_U7698, P1_U7699, P1_U7700, P1_U7701, P1_U7702, P1_U7703, P1_U7704, P1_U7705, P1_U7706, P1_U7707, P1_U7708, P1_U7709, P1_U7710, P1_U7711, P1_U7712, P1_U7713, P1_U7714, P1_U7715, P1_U7716, P1_U7717, P1_U7718, P1_U7719, P1_U7720, P1_U7721, P1_U7722, P1_U7723, P1_U7724, P1_U7725, P1_U7726, P1_U7727, P1_U7728, P1_U7729, P1_U7730, P1_U7731, P1_U7732, P1_U7733, P1_U7734, P1_U7735, P1_U7736, P1_U7737, P1_U7738, P1_U7739, P1_U7740, P1_U7741, P1_U7742, P1_U7743, P1_U7744, P1_U7745, P1_U7746, P1_U7747, P1_U7748, P1_U7749, P1_U7750, P1_U7751, P1_U7752, P1_U7753, P1_U7754, P1_U7755, P1_U7756, P1_U7757, P1_U7758, P1_U7759, P1_U7760, P1_U7761, P1_U7762, P1_U7763, P1_U7764, P1_U7765, P1_U7766, P1_U7767, P1_U7768, P1_U7769, P1_U7770, P1_U7771, P1_U7772, P1_U7773, P1_U7774, P1_U7775, P1_U7776, P1_U7777, P1_U7778, P1_U7779, P1_U7780, P1_U7781, P1_U7782, P1_U7783, P1_U7784, P1_U7785, P1_U7786, P1_U7787, P1_U7788, P1_U7789, P1_U7790, P1_U7791, P1_U7792, P1_U7793, P1_U7794, P2_ADD_371_1212_U10, P2_ADD_371_1212_U100, P2_ADD_371_1212_U101, P2_ADD_371_1212_U102, P2_ADD_371_1212_U103, P2_ADD_371_1212_U104, P2_ADD_371_1212_U105, P2_ADD_371_1212_U106, P2_ADD_371_1212_U107, P2_ADD_371_1212_U108, P2_ADD_371_1212_U109, P2_ADD_371_1212_U11, P2_ADD_371_1212_U110, P2_ADD_371_1212_U111, P2_ADD_371_1212_U112, P2_ADD_371_1212_U113, P2_ADD_371_1212_U114, P2_ADD_371_1212_U115, P2_ADD_371_1212_U116, P2_ADD_371_1212_U117, P2_ADD_371_1212_U118, P2_ADD_371_1212_U119, P2_ADD_371_1212_U12, P2_ADD_371_1212_U120, P2_ADD_371_1212_U121, P2_ADD_371_1212_U122, P2_ADD_371_1212_U123, P2_ADD_371_1212_U124, P2_ADD_371_1212_U125, P2_ADD_371_1212_U126, P2_ADD_371_1212_U127, P2_ADD_371_1212_U128, P2_ADD_371_1212_U129, P2_ADD_371_1212_U13, P2_ADD_371_1212_U130, P2_ADD_371_1212_U131, P2_ADD_371_1212_U132, P2_ADD_371_1212_U133, P2_ADD_371_1212_U134, P2_ADD_371_1212_U135, P2_ADD_371_1212_U136, P2_ADD_371_1212_U137, P2_ADD_371_1212_U138, P2_ADD_371_1212_U139, P2_ADD_371_1212_U14, P2_ADD_371_1212_U140, P2_ADD_371_1212_U141, P2_ADD_371_1212_U142, P2_ADD_371_1212_U143, P2_ADD_371_1212_U144, P2_ADD_371_1212_U145, P2_ADD_371_1212_U146, P2_ADD_371_1212_U147, P2_ADD_371_1212_U148, P2_ADD_371_1212_U149, P2_ADD_371_1212_U15, P2_ADD_371_1212_U150, P2_ADD_371_1212_U151, P2_ADD_371_1212_U152, P2_ADD_371_1212_U153, P2_ADD_371_1212_U154, P2_ADD_371_1212_U155, P2_ADD_371_1212_U156, P2_ADD_371_1212_U157, P2_ADD_371_1212_U158, P2_ADD_371_1212_U159, P2_ADD_371_1212_U16, P2_ADD_371_1212_U160, P2_ADD_371_1212_U161, P2_ADD_371_1212_U162, P2_ADD_371_1212_U163, P2_ADD_371_1212_U164, P2_ADD_371_1212_U165, P2_ADD_371_1212_U166, P2_ADD_371_1212_U167, P2_ADD_371_1212_U168, P2_ADD_371_1212_U169, P2_ADD_371_1212_U17, P2_ADD_371_1212_U170, P2_ADD_371_1212_U171, P2_ADD_371_1212_U172, P2_ADD_371_1212_U173, P2_ADD_371_1212_U174, P2_ADD_371_1212_U175, P2_ADD_371_1212_U176, P2_ADD_371_1212_U177, P2_ADD_371_1212_U178, P2_ADD_371_1212_U179, P2_ADD_371_1212_U18, P2_ADD_371_1212_U180, P2_ADD_371_1212_U181, P2_ADD_371_1212_U182, P2_ADD_371_1212_U183, P2_ADD_371_1212_U184, P2_ADD_371_1212_U185, P2_ADD_371_1212_U186, P2_ADD_371_1212_U187, P2_ADD_371_1212_U188, P2_ADD_371_1212_U189, P2_ADD_371_1212_U19, P2_ADD_371_1212_U190, P2_ADD_371_1212_U191, P2_ADD_371_1212_U192, P2_ADD_371_1212_U193, P2_ADD_371_1212_U194, P2_ADD_371_1212_U195, P2_ADD_371_1212_U196, P2_ADD_371_1212_U197, P2_ADD_371_1212_U198, P2_ADD_371_1212_U199, P2_ADD_371_1212_U20, P2_ADD_371_1212_U200, P2_ADD_371_1212_U201, P2_ADD_371_1212_U202, P2_ADD_371_1212_U203, P2_ADD_371_1212_U204, P2_ADD_371_1212_U205, P2_ADD_371_1212_U206, P2_ADD_371_1212_U207, P2_ADD_371_1212_U208, P2_ADD_371_1212_U209, P2_ADD_371_1212_U21, P2_ADD_371_1212_U210, P2_ADD_371_1212_U211, P2_ADD_371_1212_U212, P2_ADD_371_1212_U213, P2_ADD_371_1212_U214, P2_ADD_371_1212_U215, P2_ADD_371_1212_U216, P2_ADD_371_1212_U217, P2_ADD_371_1212_U218, P2_ADD_371_1212_U219, P2_ADD_371_1212_U22, P2_ADD_371_1212_U220, P2_ADD_371_1212_U221, P2_ADD_371_1212_U222, P2_ADD_371_1212_U223, P2_ADD_371_1212_U224, P2_ADD_371_1212_U225, P2_ADD_371_1212_U226, P2_ADD_371_1212_U227, P2_ADD_371_1212_U228, P2_ADD_371_1212_U229, P2_ADD_371_1212_U23, P2_ADD_371_1212_U230, P2_ADD_371_1212_U231, P2_ADD_371_1212_U232, P2_ADD_371_1212_U233, P2_ADD_371_1212_U234, P2_ADD_371_1212_U235, P2_ADD_371_1212_U236, P2_ADD_371_1212_U237, P2_ADD_371_1212_U238, P2_ADD_371_1212_U239, P2_ADD_371_1212_U24, P2_ADD_371_1212_U240, P2_ADD_371_1212_U241, P2_ADD_371_1212_U242, P2_ADD_371_1212_U243, P2_ADD_371_1212_U244, P2_ADD_371_1212_U245, P2_ADD_371_1212_U246, P2_ADD_371_1212_U247, P2_ADD_371_1212_U248, P2_ADD_371_1212_U249, P2_ADD_371_1212_U25, P2_ADD_371_1212_U250, P2_ADD_371_1212_U251, P2_ADD_371_1212_U252, P2_ADD_371_1212_U253, P2_ADD_371_1212_U254, P2_ADD_371_1212_U255, P2_ADD_371_1212_U256, P2_ADD_371_1212_U257, P2_ADD_371_1212_U258, P2_ADD_371_1212_U259, P2_ADD_371_1212_U26, P2_ADD_371_1212_U260, P2_ADD_371_1212_U261, P2_ADD_371_1212_U262, P2_ADD_371_1212_U263, P2_ADD_371_1212_U264, P2_ADD_371_1212_U265, P2_ADD_371_1212_U266, P2_ADD_371_1212_U267, P2_ADD_371_1212_U268, P2_ADD_371_1212_U269, P2_ADD_371_1212_U27, P2_ADD_371_1212_U270, P2_ADD_371_1212_U271, P2_ADD_371_1212_U272, P2_ADD_371_1212_U273, P2_ADD_371_1212_U274, P2_ADD_371_1212_U275, P2_ADD_371_1212_U276, P2_ADD_371_1212_U277, P2_ADD_371_1212_U278, P2_ADD_371_1212_U279, P2_ADD_371_1212_U28, P2_ADD_371_1212_U280, P2_ADD_371_1212_U281, P2_ADD_371_1212_U282, P2_ADD_371_1212_U29, P2_ADD_371_1212_U30, P2_ADD_371_1212_U31, P2_ADD_371_1212_U32, P2_ADD_371_1212_U33, P2_ADD_371_1212_U34, P2_ADD_371_1212_U35, P2_ADD_371_1212_U36, P2_ADD_371_1212_U37, P2_ADD_371_1212_U38, P2_ADD_371_1212_U39, P2_ADD_371_1212_U4, P2_ADD_371_1212_U40, P2_ADD_371_1212_U41, P2_ADD_371_1212_U42, P2_ADD_371_1212_U43, P2_ADD_371_1212_U44, P2_ADD_371_1212_U45, P2_ADD_371_1212_U46, P2_ADD_371_1212_U47, P2_ADD_371_1212_U48, P2_ADD_371_1212_U49, P2_ADD_371_1212_U5, P2_ADD_371_1212_U50, P2_ADD_371_1212_U51, P2_ADD_371_1212_U52, P2_ADD_371_1212_U53, P2_ADD_371_1212_U54, P2_ADD_371_1212_U55, P2_ADD_371_1212_U56, P2_ADD_371_1212_U57, P2_ADD_371_1212_U58, P2_ADD_371_1212_U59, P2_ADD_371_1212_U6, P2_ADD_371_1212_U60, P2_ADD_371_1212_U61, P2_ADD_371_1212_U62, P2_ADD_371_1212_U63, P2_ADD_371_1212_U64, P2_ADD_371_1212_U65, P2_ADD_371_1212_U66, P2_ADD_371_1212_U67, P2_ADD_371_1212_U68, P2_ADD_371_1212_U69, P2_ADD_371_1212_U7, P2_ADD_371_1212_U70, P2_ADD_371_1212_U71, P2_ADD_371_1212_U72, P2_ADD_371_1212_U73, P2_ADD_371_1212_U74, P2_ADD_371_1212_U75, P2_ADD_371_1212_U76, P2_ADD_371_1212_U77, P2_ADD_371_1212_U78, P2_ADD_371_1212_U79, P2_ADD_371_1212_U8, P2_ADD_371_1212_U80, P2_ADD_371_1212_U81, P2_ADD_371_1212_U82, P2_ADD_371_1212_U83, P2_ADD_371_1212_U84, P2_ADD_371_1212_U85, P2_ADD_371_1212_U86, P2_ADD_371_1212_U87, P2_ADD_371_1212_U88, P2_ADD_371_1212_U89, P2_ADD_371_1212_U9, P2_ADD_371_1212_U90, P2_ADD_371_1212_U91, P2_ADD_371_1212_U92, P2_ADD_371_1212_U93, P2_ADD_371_1212_U94, P2_ADD_371_1212_U95, P2_ADD_371_1212_U96, P2_ADD_371_1212_U97, P2_ADD_371_1212_U98, P2_ADD_371_1212_U99, P2_ADD_391_1196_U10, P2_ADD_391_1196_U100, P2_ADD_391_1196_U101, P2_ADD_391_1196_U102, P2_ADD_391_1196_U103, P2_ADD_391_1196_U104, P2_ADD_391_1196_U105, P2_ADD_391_1196_U106, P2_ADD_391_1196_U107, P2_ADD_391_1196_U108, P2_ADD_391_1196_U109, P2_ADD_391_1196_U11, P2_ADD_391_1196_U110, P2_ADD_391_1196_U111, P2_ADD_391_1196_U112, P2_ADD_391_1196_U113, P2_ADD_391_1196_U114, P2_ADD_391_1196_U115, P2_ADD_391_1196_U116, P2_ADD_391_1196_U117, P2_ADD_391_1196_U118, P2_ADD_391_1196_U119, P2_ADD_391_1196_U12, P2_ADD_391_1196_U120, P2_ADD_391_1196_U121, P2_ADD_391_1196_U122, P2_ADD_391_1196_U123, P2_ADD_391_1196_U124, P2_ADD_391_1196_U125, P2_ADD_391_1196_U126, P2_ADD_391_1196_U127, P2_ADD_391_1196_U128, P2_ADD_391_1196_U129, P2_ADD_391_1196_U13, P2_ADD_391_1196_U130, P2_ADD_391_1196_U131, P2_ADD_391_1196_U132, P2_ADD_391_1196_U133, P2_ADD_391_1196_U134, P2_ADD_391_1196_U135, P2_ADD_391_1196_U136, P2_ADD_391_1196_U137, P2_ADD_391_1196_U138, P2_ADD_391_1196_U139, P2_ADD_391_1196_U14, P2_ADD_391_1196_U140, P2_ADD_391_1196_U141, P2_ADD_391_1196_U142, P2_ADD_391_1196_U143, P2_ADD_391_1196_U144, P2_ADD_391_1196_U145, P2_ADD_391_1196_U146, P2_ADD_391_1196_U147, P2_ADD_391_1196_U148, P2_ADD_391_1196_U149, P2_ADD_391_1196_U15, P2_ADD_391_1196_U150, P2_ADD_391_1196_U151, P2_ADD_391_1196_U152, P2_ADD_391_1196_U153, P2_ADD_391_1196_U154, P2_ADD_391_1196_U155, P2_ADD_391_1196_U156, P2_ADD_391_1196_U157, P2_ADD_391_1196_U158, P2_ADD_391_1196_U159, P2_ADD_391_1196_U16, P2_ADD_391_1196_U160, P2_ADD_391_1196_U161, P2_ADD_391_1196_U162, P2_ADD_391_1196_U163, P2_ADD_391_1196_U164, P2_ADD_391_1196_U165, P2_ADD_391_1196_U166, P2_ADD_391_1196_U167, P2_ADD_391_1196_U168, P2_ADD_391_1196_U169, P2_ADD_391_1196_U17, P2_ADD_391_1196_U170, P2_ADD_391_1196_U171, P2_ADD_391_1196_U172, P2_ADD_391_1196_U173, P2_ADD_391_1196_U174, P2_ADD_391_1196_U175, P2_ADD_391_1196_U176, P2_ADD_391_1196_U177, P2_ADD_391_1196_U178, P2_ADD_391_1196_U179, P2_ADD_391_1196_U18, P2_ADD_391_1196_U180, P2_ADD_391_1196_U181, P2_ADD_391_1196_U182, P2_ADD_391_1196_U183, P2_ADD_391_1196_U184, P2_ADD_391_1196_U185, P2_ADD_391_1196_U186, P2_ADD_391_1196_U187, P2_ADD_391_1196_U188, P2_ADD_391_1196_U189, P2_ADD_391_1196_U19, P2_ADD_391_1196_U190, P2_ADD_391_1196_U191, P2_ADD_391_1196_U192, P2_ADD_391_1196_U193, P2_ADD_391_1196_U194, P2_ADD_391_1196_U195, P2_ADD_391_1196_U196, P2_ADD_391_1196_U197, P2_ADD_391_1196_U198, P2_ADD_391_1196_U199, P2_ADD_391_1196_U20, P2_ADD_391_1196_U200, P2_ADD_391_1196_U201, P2_ADD_391_1196_U202, P2_ADD_391_1196_U203, P2_ADD_391_1196_U204, P2_ADD_391_1196_U205, P2_ADD_391_1196_U206, P2_ADD_391_1196_U207, P2_ADD_391_1196_U208, P2_ADD_391_1196_U209, P2_ADD_391_1196_U21, P2_ADD_391_1196_U210, P2_ADD_391_1196_U211, P2_ADD_391_1196_U212, P2_ADD_391_1196_U213, P2_ADD_391_1196_U214, P2_ADD_391_1196_U215, P2_ADD_391_1196_U216, P2_ADD_391_1196_U217, P2_ADD_391_1196_U218, P2_ADD_391_1196_U219, P2_ADD_391_1196_U22, P2_ADD_391_1196_U220, P2_ADD_391_1196_U221, P2_ADD_391_1196_U222, P2_ADD_391_1196_U223, P2_ADD_391_1196_U224, P2_ADD_391_1196_U225, P2_ADD_391_1196_U226, P2_ADD_391_1196_U227, P2_ADD_391_1196_U228, P2_ADD_391_1196_U229, P2_ADD_391_1196_U23, P2_ADD_391_1196_U230, P2_ADD_391_1196_U231, P2_ADD_391_1196_U232, P2_ADD_391_1196_U233, P2_ADD_391_1196_U234, P2_ADD_391_1196_U235, P2_ADD_391_1196_U236, P2_ADD_391_1196_U237, P2_ADD_391_1196_U238, P2_ADD_391_1196_U239, P2_ADD_391_1196_U24, P2_ADD_391_1196_U240, P2_ADD_391_1196_U241, P2_ADD_391_1196_U242, P2_ADD_391_1196_U243, P2_ADD_391_1196_U244, P2_ADD_391_1196_U245, P2_ADD_391_1196_U246, P2_ADD_391_1196_U247, P2_ADD_391_1196_U248, P2_ADD_391_1196_U249, P2_ADD_391_1196_U25, P2_ADD_391_1196_U250, P2_ADD_391_1196_U251, P2_ADD_391_1196_U252, P2_ADD_391_1196_U253, P2_ADD_391_1196_U254, P2_ADD_391_1196_U255, P2_ADD_391_1196_U256, P2_ADD_391_1196_U257, P2_ADD_391_1196_U258, P2_ADD_391_1196_U259, P2_ADD_391_1196_U26, P2_ADD_391_1196_U260, P2_ADD_391_1196_U261, P2_ADD_391_1196_U262, P2_ADD_391_1196_U263, P2_ADD_391_1196_U264, P2_ADD_391_1196_U265, P2_ADD_391_1196_U266, P2_ADD_391_1196_U267, P2_ADD_391_1196_U268, P2_ADD_391_1196_U269, P2_ADD_391_1196_U27, P2_ADD_391_1196_U270, P2_ADD_391_1196_U271, P2_ADD_391_1196_U272, P2_ADD_391_1196_U273, P2_ADD_391_1196_U274, P2_ADD_391_1196_U275, P2_ADD_391_1196_U276, P2_ADD_391_1196_U277, P2_ADD_391_1196_U278, P2_ADD_391_1196_U279, P2_ADD_391_1196_U28, P2_ADD_391_1196_U280, P2_ADD_391_1196_U281, P2_ADD_391_1196_U282, P2_ADD_391_1196_U283, P2_ADD_391_1196_U284, P2_ADD_391_1196_U285, P2_ADD_391_1196_U286, P2_ADD_391_1196_U287, P2_ADD_391_1196_U288, P2_ADD_391_1196_U289, P2_ADD_391_1196_U29, P2_ADD_391_1196_U290, P2_ADD_391_1196_U291, P2_ADD_391_1196_U292, P2_ADD_391_1196_U293, P2_ADD_391_1196_U294, P2_ADD_391_1196_U295, P2_ADD_391_1196_U296, P2_ADD_391_1196_U297, P2_ADD_391_1196_U298, P2_ADD_391_1196_U299, P2_ADD_391_1196_U30, P2_ADD_391_1196_U300, P2_ADD_391_1196_U301, P2_ADD_391_1196_U302, P2_ADD_391_1196_U303, P2_ADD_391_1196_U304, P2_ADD_391_1196_U305, P2_ADD_391_1196_U306, P2_ADD_391_1196_U307, P2_ADD_391_1196_U308, P2_ADD_391_1196_U309, P2_ADD_391_1196_U31, P2_ADD_391_1196_U310, P2_ADD_391_1196_U311, P2_ADD_391_1196_U312, P2_ADD_391_1196_U313, P2_ADD_391_1196_U314, P2_ADD_391_1196_U315, P2_ADD_391_1196_U316, P2_ADD_391_1196_U317, P2_ADD_391_1196_U318, P2_ADD_391_1196_U319, P2_ADD_391_1196_U32, P2_ADD_391_1196_U320, P2_ADD_391_1196_U321, P2_ADD_391_1196_U322, P2_ADD_391_1196_U323, P2_ADD_391_1196_U324, P2_ADD_391_1196_U325, P2_ADD_391_1196_U326, P2_ADD_391_1196_U327, P2_ADD_391_1196_U328, P2_ADD_391_1196_U329, P2_ADD_391_1196_U33, P2_ADD_391_1196_U330, P2_ADD_391_1196_U331, P2_ADD_391_1196_U332, P2_ADD_391_1196_U333, P2_ADD_391_1196_U334, P2_ADD_391_1196_U335, P2_ADD_391_1196_U336, P2_ADD_391_1196_U337, P2_ADD_391_1196_U338, P2_ADD_391_1196_U339, P2_ADD_391_1196_U34, P2_ADD_391_1196_U340, P2_ADD_391_1196_U341, P2_ADD_391_1196_U342, P2_ADD_391_1196_U343, P2_ADD_391_1196_U344, P2_ADD_391_1196_U345, P2_ADD_391_1196_U346, P2_ADD_391_1196_U347, P2_ADD_391_1196_U348, P2_ADD_391_1196_U349, P2_ADD_391_1196_U35, P2_ADD_391_1196_U350, P2_ADD_391_1196_U351, P2_ADD_391_1196_U352, P2_ADD_391_1196_U353, P2_ADD_391_1196_U354, P2_ADD_391_1196_U355, P2_ADD_391_1196_U356, P2_ADD_391_1196_U357, P2_ADD_391_1196_U358, P2_ADD_391_1196_U359, P2_ADD_391_1196_U36, P2_ADD_391_1196_U360, P2_ADD_391_1196_U361, P2_ADD_391_1196_U362, P2_ADD_391_1196_U363, P2_ADD_391_1196_U364, P2_ADD_391_1196_U365, P2_ADD_391_1196_U366, P2_ADD_391_1196_U367, P2_ADD_391_1196_U368, P2_ADD_391_1196_U369, P2_ADD_391_1196_U37, P2_ADD_391_1196_U370, P2_ADD_391_1196_U371, P2_ADD_391_1196_U372, P2_ADD_391_1196_U373, P2_ADD_391_1196_U374, P2_ADD_391_1196_U375, P2_ADD_391_1196_U376, P2_ADD_391_1196_U377, P2_ADD_391_1196_U378, P2_ADD_391_1196_U379, P2_ADD_391_1196_U38, P2_ADD_391_1196_U380, P2_ADD_391_1196_U381, P2_ADD_391_1196_U382, P2_ADD_391_1196_U383, P2_ADD_391_1196_U384, P2_ADD_391_1196_U385, P2_ADD_391_1196_U386, P2_ADD_391_1196_U387, P2_ADD_391_1196_U388, P2_ADD_391_1196_U389, P2_ADD_391_1196_U39, P2_ADD_391_1196_U390, P2_ADD_391_1196_U391, P2_ADD_391_1196_U392, P2_ADD_391_1196_U393, P2_ADD_391_1196_U394, P2_ADD_391_1196_U395, P2_ADD_391_1196_U396, P2_ADD_391_1196_U397, P2_ADD_391_1196_U398, P2_ADD_391_1196_U399, P2_ADD_391_1196_U40, P2_ADD_391_1196_U400, P2_ADD_391_1196_U401, P2_ADD_391_1196_U402, P2_ADD_391_1196_U403, P2_ADD_391_1196_U404, P2_ADD_391_1196_U405, P2_ADD_391_1196_U406, P2_ADD_391_1196_U407, P2_ADD_391_1196_U408, P2_ADD_391_1196_U409, P2_ADD_391_1196_U41, P2_ADD_391_1196_U410, P2_ADD_391_1196_U411, P2_ADD_391_1196_U412, P2_ADD_391_1196_U413, P2_ADD_391_1196_U414, P2_ADD_391_1196_U415, P2_ADD_391_1196_U416, P2_ADD_391_1196_U417, P2_ADD_391_1196_U418, P2_ADD_391_1196_U419, P2_ADD_391_1196_U42, P2_ADD_391_1196_U420, P2_ADD_391_1196_U421, P2_ADD_391_1196_U422, P2_ADD_391_1196_U423, P2_ADD_391_1196_U424, P2_ADD_391_1196_U425, P2_ADD_391_1196_U426, P2_ADD_391_1196_U427, P2_ADD_391_1196_U428, P2_ADD_391_1196_U429, P2_ADD_391_1196_U43, P2_ADD_391_1196_U430, P2_ADD_391_1196_U431, P2_ADD_391_1196_U432, P2_ADD_391_1196_U433, P2_ADD_391_1196_U434, P2_ADD_391_1196_U435, P2_ADD_391_1196_U436, P2_ADD_391_1196_U437, P2_ADD_391_1196_U438, P2_ADD_391_1196_U439, P2_ADD_391_1196_U44, P2_ADD_391_1196_U440, P2_ADD_391_1196_U441, P2_ADD_391_1196_U442, P2_ADD_391_1196_U443, P2_ADD_391_1196_U444, P2_ADD_391_1196_U445, P2_ADD_391_1196_U446, P2_ADD_391_1196_U447, P2_ADD_391_1196_U448, P2_ADD_391_1196_U449, P2_ADD_391_1196_U45, P2_ADD_391_1196_U450, P2_ADD_391_1196_U451, P2_ADD_391_1196_U452, P2_ADD_391_1196_U453, P2_ADD_391_1196_U454, P2_ADD_391_1196_U455, P2_ADD_391_1196_U456, P2_ADD_391_1196_U457, P2_ADD_391_1196_U458, P2_ADD_391_1196_U459, P2_ADD_391_1196_U46, P2_ADD_391_1196_U460, P2_ADD_391_1196_U461, P2_ADD_391_1196_U462, P2_ADD_391_1196_U463, P2_ADD_391_1196_U464, P2_ADD_391_1196_U465, P2_ADD_391_1196_U466, P2_ADD_391_1196_U467, P2_ADD_391_1196_U468, P2_ADD_391_1196_U469, P2_ADD_391_1196_U47, P2_ADD_391_1196_U470, P2_ADD_391_1196_U471, P2_ADD_391_1196_U472, P2_ADD_391_1196_U473, P2_ADD_391_1196_U474, P2_ADD_391_1196_U475, P2_ADD_391_1196_U476, P2_ADD_391_1196_U477, P2_ADD_391_1196_U478, P2_ADD_391_1196_U48, P2_ADD_391_1196_U49, P2_ADD_391_1196_U5, P2_ADD_391_1196_U50, P2_ADD_391_1196_U51, P2_ADD_391_1196_U52, P2_ADD_391_1196_U53, P2_ADD_391_1196_U54, P2_ADD_391_1196_U55, P2_ADD_391_1196_U56, P2_ADD_391_1196_U57, P2_ADD_391_1196_U58, P2_ADD_391_1196_U59, P2_ADD_391_1196_U6, P2_ADD_391_1196_U60, P2_ADD_391_1196_U61, P2_ADD_391_1196_U62, P2_ADD_391_1196_U63, P2_ADD_391_1196_U64, P2_ADD_391_1196_U65, P2_ADD_391_1196_U66, P2_ADD_391_1196_U67, P2_ADD_391_1196_U68, P2_ADD_391_1196_U69, P2_ADD_391_1196_U7, P2_ADD_391_1196_U70, P2_ADD_391_1196_U71, P2_ADD_391_1196_U72, P2_ADD_391_1196_U73, P2_ADD_391_1196_U74, P2_ADD_391_1196_U75, P2_ADD_391_1196_U76, P2_ADD_391_1196_U77, P2_ADD_391_1196_U78, P2_ADD_391_1196_U79, P2_ADD_391_1196_U8, P2_ADD_391_1196_U80, P2_ADD_391_1196_U81, P2_ADD_391_1196_U82, P2_ADD_391_1196_U83, P2_ADD_391_1196_U84, P2_ADD_391_1196_U85, P2_ADD_391_1196_U86, P2_ADD_391_1196_U87, P2_ADD_391_1196_U88, P2_ADD_391_1196_U89, P2_ADD_391_1196_U9, P2_ADD_391_1196_U90, P2_ADD_391_1196_U91, P2_ADD_391_1196_U92, P2_ADD_391_1196_U93, P2_ADD_391_1196_U94, P2_ADD_391_1196_U95, P2_ADD_391_1196_U96, P2_ADD_391_1196_U97, P2_ADD_391_1196_U98, P2_ADD_391_1196_U99, P2_ADD_394_U10, P2_ADD_394_U100, P2_ADD_394_U101, P2_ADD_394_U102, P2_ADD_394_U103, P2_ADD_394_U104, P2_ADD_394_U105, P2_ADD_394_U106, P2_ADD_394_U107, P2_ADD_394_U108, P2_ADD_394_U109, P2_ADD_394_U11, P2_ADD_394_U110, P2_ADD_394_U111, P2_ADD_394_U112, P2_ADD_394_U113, P2_ADD_394_U114, P2_ADD_394_U115, P2_ADD_394_U116, P2_ADD_394_U117, P2_ADD_394_U118, P2_ADD_394_U119, P2_ADD_394_U12, P2_ADD_394_U120, P2_ADD_394_U121, P2_ADD_394_U122, P2_ADD_394_U123, P2_ADD_394_U124, P2_ADD_394_U125, P2_ADD_394_U126, P2_ADD_394_U127, P2_ADD_394_U128, P2_ADD_394_U129, P2_ADD_394_U13, P2_ADD_394_U130, P2_ADD_394_U131, P2_ADD_394_U132, P2_ADD_394_U133, P2_ADD_394_U134, P2_ADD_394_U135, P2_ADD_394_U136, P2_ADD_394_U137, P2_ADD_394_U138, P2_ADD_394_U139, P2_ADD_394_U14, P2_ADD_394_U140, P2_ADD_394_U141, P2_ADD_394_U142, P2_ADD_394_U143, P2_ADD_394_U144, P2_ADD_394_U145, P2_ADD_394_U146, P2_ADD_394_U147, P2_ADD_394_U148, P2_ADD_394_U149, P2_ADD_394_U15, P2_ADD_394_U150, P2_ADD_394_U151, P2_ADD_394_U152, P2_ADD_394_U153, P2_ADD_394_U154, P2_ADD_394_U155, P2_ADD_394_U156, P2_ADD_394_U157, P2_ADD_394_U158, P2_ADD_394_U159, P2_ADD_394_U16, P2_ADD_394_U160, P2_ADD_394_U161, P2_ADD_394_U162, P2_ADD_394_U163, P2_ADD_394_U164, P2_ADD_394_U165, P2_ADD_394_U166, P2_ADD_394_U167, P2_ADD_394_U168, P2_ADD_394_U169, P2_ADD_394_U17, P2_ADD_394_U170, P2_ADD_394_U171, P2_ADD_394_U172, P2_ADD_394_U173, P2_ADD_394_U174, P2_ADD_394_U175, P2_ADD_394_U176, P2_ADD_394_U177, P2_ADD_394_U178, P2_ADD_394_U179, P2_ADD_394_U18, P2_ADD_394_U180, P2_ADD_394_U181, P2_ADD_394_U182, P2_ADD_394_U183, P2_ADD_394_U184, P2_ADD_394_U185, P2_ADD_394_U186, P2_ADD_394_U19, P2_ADD_394_U20, P2_ADD_394_U21, P2_ADD_394_U22, P2_ADD_394_U23, P2_ADD_394_U24, P2_ADD_394_U25, P2_ADD_394_U26, P2_ADD_394_U27, P2_ADD_394_U28, P2_ADD_394_U29, P2_ADD_394_U30, P2_ADD_394_U31, P2_ADD_394_U32, P2_ADD_394_U33, P2_ADD_394_U34, P2_ADD_394_U35, P2_ADD_394_U36, P2_ADD_394_U37, P2_ADD_394_U38, P2_ADD_394_U39, P2_ADD_394_U4, P2_ADD_394_U40, P2_ADD_394_U41, P2_ADD_394_U42, P2_ADD_394_U43, P2_ADD_394_U44, P2_ADD_394_U45, P2_ADD_394_U46, P2_ADD_394_U47, P2_ADD_394_U48, P2_ADD_394_U49, P2_ADD_394_U5, P2_ADD_394_U50, P2_ADD_394_U51, P2_ADD_394_U52, P2_ADD_394_U53, P2_ADD_394_U54, P2_ADD_394_U55, P2_ADD_394_U56, P2_ADD_394_U57, P2_ADD_394_U58, P2_ADD_394_U59, P2_ADD_394_U6, P2_ADD_394_U60, P2_ADD_394_U61, P2_ADD_394_U62, P2_ADD_394_U63, P2_ADD_394_U64, P2_ADD_394_U65, P2_ADD_394_U66, P2_ADD_394_U67, P2_ADD_394_U68, P2_ADD_394_U69, P2_ADD_394_U7, P2_ADD_394_U70, P2_ADD_394_U71, P2_ADD_394_U72, P2_ADD_394_U73, P2_ADD_394_U74, P2_ADD_394_U75, P2_ADD_394_U76, P2_ADD_394_U77, P2_ADD_394_U78, P2_ADD_394_U79, P2_ADD_394_U8, P2_ADD_394_U80, P2_ADD_394_U81, P2_ADD_394_U82, P2_ADD_394_U83, P2_ADD_394_U84, P2_ADD_394_U85, P2_ADD_394_U86, P2_ADD_394_U87, P2_ADD_394_U88, P2_ADD_394_U89, P2_ADD_394_U9, P2_ADD_394_U90, P2_ADD_394_U91, P2_ADD_394_U92, P2_ADD_394_U93, P2_ADD_394_U94, P2_ADD_394_U95, P2_ADD_394_U96, P2_ADD_394_U97, P2_ADD_394_U98, P2_ADD_394_U99, P2_ADD_402_1132_U10, P2_ADD_402_1132_U11, P2_ADD_402_1132_U12, P2_ADD_402_1132_U13, P2_ADD_402_1132_U14, P2_ADD_402_1132_U15, P2_ADD_402_1132_U16, P2_ADD_402_1132_U17, P2_ADD_402_1132_U18, P2_ADD_402_1132_U19, P2_ADD_402_1132_U20, P2_ADD_402_1132_U21, P2_ADD_402_1132_U22, P2_ADD_402_1132_U23, P2_ADD_402_1132_U24, P2_ADD_402_1132_U25, P2_ADD_402_1132_U26, P2_ADD_402_1132_U27, P2_ADD_402_1132_U28, P2_ADD_402_1132_U29, P2_ADD_402_1132_U30, P2_ADD_402_1132_U31, P2_ADD_402_1132_U32, P2_ADD_402_1132_U33, P2_ADD_402_1132_U34, P2_ADD_402_1132_U35, P2_ADD_402_1132_U36, P2_ADD_402_1132_U37, P2_ADD_402_1132_U38, P2_ADD_402_1132_U39, P2_ADD_402_1132_U4, P2_ADD_402_1132_U40, P2_ADD_402_1132_U41, P2_ADD_402_1132_U42, P2_ADD_402_1132_U43, P2_ADD_402_1132_U44, P2_ADD_402_1132_U45, P2_ADD_402_1132_U46, P2_ADD_402_1132_U47, P2_ADD_402_1132_U48, P2_ADD_402_1132_U49, P2_ADD_402_1132_U5, P2_ADD_402_1132_U50, P2_ADD_402_1132_U6, P2_ADD_402_1132_U7, P2_ADD_402_1132_U8, P2_ADD_402_1132_U9, P2_GTE_370_U6, P2_GTE_370_U7, P2_GTE_370_U8, P2_GTE_370_U9, P2_LT_563_1260_U6, P2_LT_563_1260_U7, P2_LT_563_U10, P2_LT_563_U11, P2_LT_563_U12, P2_LT_563_U13, P2_LT_563_U14, P2_LT_563_U15, P2_LT_563_U16, P2_LT_563_U17, P2_LT_563_U18, P2_LT_563_U19, P2_LT_563_U20, P2_LT_563_U21, P2_LT_563_U22, P2_LT_563_U23, P2_LT_563_U24, P2_LT_563_U25, P2_LT_563_U26, P2_LT_563_U27, P2_LT_563_U6, P2_LT_563_U7, P2_LT_563_U8, P2_LT_563_U9, P2_R1957_U10, P2_R1957_U100, P2_R1957_U101, P2_R1957_U102, P2_R1957_U103, P2_R1957_U104, P2_R1957_U105, P2_R1957_U106, P2_R1957_U107, P2_R1957_U108, P2_R1957_U109, P2_R1957_U11, P2_R1957_U110, P2_R1957_U111, P2_R1957_U112, P2_R1957_U113, P2_R1957_U114, P2_R1957_U115, P2_R1957_U116, P2_R1957_U117, P2_R1957_U118, P2_R1957_U119, P2_R1957_U12, P2_R1957_U120, P2_R1957_U121, P2_R1957_U122, P2_R1957_U123, P2_R1957_U124, P2_R1957_U125, P2_R1957_U126, P2_R1957_U127, P2_R1957_U128, P2_R1957_U129, P2_R1957_U13, P2_R1957_U130, P2_R1957_U131, P2_R1957_U132, P2_R1957_U133, P2_R1957_U134, P2_R1957_U135, P2_R1957_U136, P2_R1957_U137, P2_R1957_U138, P2_R1957_U139, P2_R1957_U14, P2_R1957_U140, P2_R1957_U141, P2_R1957_U142, P2_R1957_U143, P2_R1957_U144, P2_R1957_U145, P2_R1957_U146, P2_R1957_U147, P2_R1957_U148, P2_R1957_U149, P2_R1957_U15, P2_R1957_U150, P2_R1957_U151, P2_R1957_U152, P2_R1957_U153, P2_R1957_U154, P2_R1957_U155, P2_R1957_U156, P2_R1957_U157, P2_R1957_U158, P2_R1957_U159, P2_R1957_U16, P2_R1957_U17, P2_R1957_U18, P2_R1957_U19, P2_R1957_U20, P2_R1957_U21, P2_R1957_U22, P2_R1957_U23, P2_R1957_U24, P2_R1957_U25, P2_R1957_U26, P2_R1957_U27, P2_R1957_U28, P2_R1957_U29, P2_R1957_U30, P2_R1957_U31, P2_R1957_U32, P2_R1957_U33, P2_R1957_U34, P2_R1957_U35, P2_R1957_U36, P2_R1957_U37, P2_R1957_U38, P2_R1957_U39, P2_R1957_U40, P2_R1957_U41, P2_R1957_U42, P2_R1957_U43, P2_R1957_U44, P2_R1957_U45, P2_R1957_U46, P2_R1957_U47, P2_R1957_U48, P2_R1957_U49, P2_R1957_U50, P2_R1957_U51, P2_R1957_U52, P2_R1957_U53, P2_R1957_U54, P2_R1957_U55, P2_R1957_U56, P2_R1957_U57, P2_R1957_U58, P2_R1957_U59, P2_R1957_U6, P2_R1957_U60, P2_R1957_U61, P2_R1957_U62, P2_R1957_U63, P2_R1957_U64, P2_R1957_U65, P2_R1957_U66, P2_R1957_U67, P2_R1957_U68, P2_R1957_U69, P2_R1957_U7, P2_R1957_U70, P2_R1957_U71, P2_R1957_U72, P2_R1957_U73, P2_R1957_U74, P2_R1957_U75, P2_R1957_U76, P2_R1957_U77, P2_R1957_U78, P2_R1957_U79, P2_R1957_U8, P2_R1957_U80, P2_R1957_U81, P2_R1957_U82, P2_R1957_U83, P2_R1957_U84, P2_R1957_U85, P2_R1957_U86, P2_R1957_U87, P2_R1957_U88, P2_R1957_U89, P2_R1957_U9, P2_R1957_U90, P2_R1957_U91, P2_R1957_U92, P2_R1957_U93, P2_R1957_U94, P2_R1957_U95, P2_R1957_U96, P2_R1957_U97, P2_R1957_U98, P2_R1957_U99, P2_R2027_U10, P2_R2027_U100, P2_R2027_U101, P2_R2027_U102, P2_R2027_U103, P2_R2027_U104, P2_R2027_U105, P2_R2027_U106, P2_R2027_U107, P2_R2027_U108, P2_R2027_U109, P2_R2027_U11, P2_R2027_U110, P2_R2027_U111, P2_R2027_U112, P2_R2027_U113, P2_R2027_U114, P2_R2027_U115, P2_R2027_U116, P2_R2027_U117, P2_R2027_U118, P2_R2027_U119, P2_R2027_U12, P2_R2027_U120, P2_R2027_U121, P2_R2027_U122, P2_R2027_U123, P2_R2027_U124, P2_R2027_U125, P2_R2027_U126, P2_R2027_U127, P2_R2027_U128, P2_R2027_U129, P2_R2027_U13, P2_R2027_U130, P2_R2027_U131, P2_R2027_U132, P2_R2027_U133, P2_R2027_U134, P2_R2027_U135, P2_R2027_U136, P2_R2027_U137, P2_R2027_U138, P2_R2027_U139, P2_R2027_U14, P2_R2027_U140, P2_R2027_U141, P2_R2027_U142, P2_R2027_U143, P2_R2027_U144, P2_R2027_U145, P2_R2027_U146, P2_R2027_U147, P2_R2027_U148, P2_R2027_U149, P2_R2027_U15, P2_R2027_U150, P2_R2027_U151, P2_R2027_U152, P2_R2027_U153, P2_R2027_U154, P2_R2027_U155, P2_R2027_U156, P2_R2027_U157, P2_R2027_U158, P2_R2027_U159, P2_R2027_U16, P2_R2027_U160, P2_R2027_U161, P2_R2027_U162, P2_R2027_U163, P2_R2027_U164, P2_R2027_U165, P2_R2027_U166, P2_R2027_U167, P2_R2027_U168, P2_R2027_U169, P2_R2027_U17, P2_R2027_U170, P2_R2027_U171, P2_R2027_U172, P2_R2027_U173, P2_R2027_U174, P2_R2027_U175, P2_R2027_U176, P2_R2027_U177, P2_R2027_U178, P2_R2027_U179, P2_R2027_U18, P2_R2027_U180, P2_R2027_U181, P2_R2027_U182, P2_R2027_U183, P2_R2027_U184, P2_R2027_U185, P2_R2027_U186, P2_R2027_U187, P2_R2027_U188, P2_R2027_U189, P2_R2027_U19, P2_R2027_U20, P2_R2027_U21, P2_R2027_U22, P2_R2027_U23, P2_R2027_U24, P2_R2027_U25, P2_R2027_U26, P2_R2027_U27, P2_R2027_U28, P2_R2027_U29, P2_R2027_U30, P2_R2027_U31, P2_R2027_U32, P2_R2027_U33, P2_R2027_U34, P2_R2027_U35, P2_R2027_U36, P2_R2027_U37, P2_R2027_U38, P2_R2027_U39, P2_R2027_U40, P2_R2027_U41, P2_R2027_U42, P2_R2027_U43, P2_R2027_U44, P2_R2027_U45, P2_R2027_U46, P2_R2027_U47, P2_R2027_U48, P2_R2027_U49, P2_R2027_U5, P2_R2027_U50, P2_R2027_U51, P2_R2027_U52, P2_R2027_U53, P2_R2027_U54, P2_R2027_U55, P2_R2027_U56, P2_R2027_U57, P2_R2027_U58, P2_R2027_U59, P2_R2027_U6, P2_R2027_U60, P2_R2027_U61, P2_R2027_U62, P2_R2027_U63, P2_R2027_U64, P2_R2027_U65, P2_R2027_U66, P2_R2027_U67, P2_R2027_U68, P2_R2027_U69, P2_R2027_U7, P2_R2027_U70, P2_R2027_U71, P2_R2027_U72, P2_R2027_U73, P2_R2027_U74, P2_R2027_U75, P2_R2027_U76, P2_R2027_U77, P2_R2027_U78, P2_R2027_U79, P2_R2027_U8, P2_R2027_U80, P2_R2027_U81, P2_R2027_U82, P2_R2027_U83, P2_R2027_U84, P2_R2027_U85, P2_R2027_U86, P2_R2027_U87, P2_R2027_U88, P2_R2027_U89, P2_R2027_U9, P2_R2027_U90, P2_R2027_U91, P2_R2027_U92, P2_R2027_U93, P2_R2027_U94, P2_R2027_U95, P2_R2027_U96, P2_R2027_U97, P2_R2027_U98, P2_R2027_U99, P2_R2088_U6, P2_R2088_U7, P2_R2096_U10, P2_R2096_U100, P2_R2096_U101, P2_R2096_U102, P2_R2096_U103, P2_R2096_U104, P2_R2096_U105, P2_R2096_U106, P2_R2096_U107, P2_R2096_U108, P2_R2096_U109, P2_R2096_U11, P2_R2096_U110, P2_R2096_U111, P2_R2096_U112, P2_R2096_U113, P2_R2096_U114, P2_R2096_U115, P2_R2096_U116, P2_R2096_U117, P2_R2096_U118, P2_R2096_U119, P2_R2096_U12, P2_R2096_U120, P2_R2096_U121, P2_R2096_U122, P2_R2096_U123, P2_R2096_U124, P2_R2096_U125, P2_R2096_U126, P2_R2096_U127, P2_R2096_U128, P2_R2096_U129, P2_R2096_U13, P2_R2096_U130, P2_R2096_U131, P2_R2096_U132, P2_R2096_U133, P2_R2096_U134, P2_R2096_U135, P2_R2096_U136, P2_R2096_U137, P2_R2096_U138, P2_R2096_U139, P2_R2096_U14, P2_R2096_U140, P2_R2096_U141, P2_R2096_U142, P2_R2096_U143, P2_R2096_U144, P2_R2096_U145, P2_R2096_U146, P2_R2096_U147, P2_R2096_U148, P2_R2096_U149, P2_R2096_U15, P2_R2096_U150, P2_R2096_U151, P2_R2096_U152, P2_R2096_U153, P2_R2096_U154, P2_R2096_U155, P2_R2096_U156, P2_R2096_U157, P2_R2096_U158, P2_R2096_U159, P2_R2096_U16, P2_R2096_U160, P2_R2096_U161, P2_R2096_U162, P2_R2096_U163, P2_R2096_U164, P2_R2096_U165, P2_R2096_U166, P2_R2096_U167, P2_R2096_U168, P2_R2096_U169, P2_R2096_U17, P2_R2096_U170, P2_R2096_U171, P2_R2096_U172, P2_R2096_U173, P2_R2096_U174, P2_R2096_U175, P2_R2096_U176, P2_R2096_U177, P2_R2096_U178, P2_R2096_U179, P2_R2096_U18, P2_R2096_U180, P2_R2096_U181, P2_R2096_U182, P2_R2096_U183, P2_R2096_U184, P2_R2096_U185, P2_R2096_U186, P2_R2096_U187, P2_R2096_U188, P2_R2096_U189, P2_R2096_U19, P2_R2096_U190, P2_R2096_U191, P2_R2096_U192, P2_R2096_U193, P2_R2096_U194, P2_R2096_U195, P2_R2096_U196, P2_R2096_U197, P2_R2096_U198, P2_R2096_U199, P2_R2096_U20, P2_R2096_U200, P2_R2096_U201, P2_R2096_U202, P2_R2096_U203, P2_R2096_U204, P2_R2096_U205, P2_R2096_U206, P2_R2096_U207, P2_R2096_U208, P2_R2096_U209, P2_R2096_U21, P2_R2096_U210, P2_R2096_U211, P2_R2096_U212, P2_R2096_U213, P2_R2096_U214, P2_R2096_U215, P2_R2096_U216, P2_R2096_U217, P2_R2096_U218, P2_R2096_U219, P2_R2096_U22, P2_R2096_U220, P2_R2096_U221, P2_R2096_U222, P2_R2096_U223, P2_R2096_U224, P2_R2096_U225, P2_R2096_U226, P2_R2096_U227, P2_R2096_U228, P2_R2096_U229, P2_R2096_U23, P2_R2096_U230, P2_R2096_U231, P2_R2096_U232, P2_R2096_U233, P2_R2096_U234, P2_R2096_U235, P2_R2096_U236, P2_R2096_U237, P2_R2096_U238, P2_R2096_U239, P2_R2096_U24, P2_R2096_U240, P2_R2096_U241, P2_R2096_U242, P2_R2096_U243, P2_R2096_U244, P2_R2096_U245, P2_R2096_U246, P2_R2096_U247, P2_R2096_U248, P2_R2096_U249, P2_R2096_U25, P2_R2096_U250, P2_R2096_U251, P2_R2096_U252, P2_R2096_U253, P2_R2096_U254, P2_R2096_U255, P2_R2096_U256, P2_R2096_U257, P2_R2096_U258, P2_R2096_U259, P2_R2096_U26, P2_R2096_U260, P2_R2096_U261, P2_R2096_U262, P2_R2096_U263, P2_R2096_U264, P2_R2096_U265, P2_R2096_U27, P2_R2096_U28, P2_R2096_U29, P2_R2096_U30, P2_R2096_U31, P2_R2096_U32, P2_R2096_U33, P2_R2096_U34, P2_R2096_U35, P2_R2096_U36, P2_R2096_U37, P2_R2096_U38, P2_R2096_U39, P2_R2096_U4, P2_R2096_U40, P2_R2096_U41, P2_R2096_U42, P2_R2096_U43, P2_R2096_U44, P2_R2096_U45, P2_R2096_U46, P2_R2096_U47, P2_R2096_U48, P2_R2096_U49, P2_R2096_U5, P2_R2096_U50, P2_R2096_U51, P2_R2096_U52, P2_R2096_U53, P2_R2096_U54, P2_R2096_U55, P2_R2096_U56, P2_R2096_U57, P2_R2096_U58, P2_R2096_U59, P2_R2096_U6, P2_R2096_U60, P2_R2096_U61, P2_R2096_U62, P2_R2096_U63, P2_R2096_U64, P2_R2096_U65, P2_R2096_U66, P2_R2096_U67, P2_R2096_U68, P2_R2096_U69, P2_R2096_U7, P2_R2096_U70, P2_R2096_U71, P2_R2096_U72, P2_R2096_U73, P2_R2096_U74, P2_R2096_U75, P2_R2096_U76, P2_R2096_U77, P2_R2096_U78, P2_R2096_U79, P2_R2096_U8, P2_R2096_U80, P2_R2096_U81, P2_R2096_U82, P2_R2096_U83, P2_R2096_U84, P2_R2096_U85, P2_R2096_U86, P2_R2096_U87, P2_R2096_U88, P2_R2096_U89, P2_R2096_U9, P2_R2096_U90, P2_R2096_U91, P2_R2096_U92, P2_R2096_U93, P2_R2096_U94, P2_R2096_U95, P2_R2096_U96, P2_R2096_U97, P2_R2096_U98, P2_R2096_U99, P2_R2099_U10, P2_R2099_U100, P2_R2099_U101, P2_R2099_U102, P2_R2099_U103, P2_R2099_U104, P2_R2099_U105, P2_R2099_U106, P2_R2099_U107, P2_R2099_U108, P2_R2099_U109, P2_R2099_U11, P2_R2099_U110, P2_R2099_U111, P2_R2099_U112, P2_R2099_U113, P2_R2099_U114, P2_R2099_U115, P2_R2099_U116, P2_R2099_U117, P2_R2099_U118, P2_R2099_U119, P2_R2099_U12, P2_R2099_U120, P2_R2099_U121, P2_R2099_U122, P2_R2099_U123, P2_R2099_U124, P2_R2099_U125, P2_R2099_U126, P2_R2099_U127, P2_R2099_U128, P2_R2099_U129, P2_R2099_U13, P2_R2099_U130, P2_R2099_U131, P2_R2099_U132, P2_R2099_U133, P2_R2099_U134, P2_R2099_U135, P2_R2099_U136, P2_R2099_U137, P2_R2099_U138, P2_R2099_U139, P2_R2099_U14, P2_R2099_U140, P2_R2099_U141, P2_R2099_U142, P2_R2099_U143, P2_R2099_U144, P2_R2099_U145, P2_R2099_U146, P2_R2099_U147, P2_R2099_U148, P2_R2099_U149, P2_R2099_U15, P2_R2099_U150, P2_R2099_U151, P2_R2099_U152, P2_R2099_U153, P2_R2099_U154, P2_R2099_U155, P2_R2099_U156, P2_R2099_U157, P2_R2099_U158, P2_R2099_U159, P2_R2099_U16, P2_R2099_U160, P2_R2099_U161, P2_R2099_U162, P2_R2099_U163, P2_R2099_U164, P2_R2099_U165, P2_R2099_U166, P2_R2099_U167, P2_R2099_U168, P2_R2099_U169, P2_R2099_U17, P2_R2099_U170, P2_R2099_U171, P2_R2099_U172, P2_R2099_U173, P2_R2099_U174, P2_R2099_U175, P2_R2099_U176, P2_R2099_U177, P2_R2099_U178, P2_R2099_U179, P2_R2099_U18, P2_R2099_U180, P2_R2099_U181, P2_R2099_U182, P2_R2099_U183, P2_R2099_U184, P2_R2099_U185, P2_R2099_U186, P2_R2099_U187, P2_R2099_U188, P2_R2099_U189, P2_R2099_U19, P2_R2099_U190, P2_R2099_U191, P2_R2099_U192, P2_R2099_U193, P2_R2099_U194, P2_R2099_U195, P2_R2099_U196, P2_R2099_U197, P2_R2099_U198, P2_R2099_U199, P2_R2099_U20, P2_R2099_U200, P2_R2099_U201, P2_R2099_U202, P2_R2099_U203, P2_R2099_U204, P2_R2099_U205, P2_R2099_U206, P2_R2099_U207, P2_R2099_U208, P2_R2099_U209, P2_R2099_U21, P2_R2099_U210, P2_R2099_U211, P2_R2099_U212, P2_R2099_U213, P2_R2099_U214, P2_R2099_U215, P2_R2099_U216, P2_R2099_U217, P2_R2099_U218, P2_R2099_U219, P2_R2099_U22, P2_R2099_U220, P2_R2099_U221, P2_R2099_U222, P2_R2099_U223, P2_R2099_U224, P2_R2099_U225, P2_R2099_U23, P2_R2099_U24, P2_R2099_U25, P2_R2099_U26, P2_R2099_U27, P2_R2099_U28, P2_R2099_U29, P2_R2099_U30, P2_R2099_U31, P2_R2099_U32, P2_R2099_U33, P2_R2099_U34, P2_R2099_U35, P2_R2099_U36, P2_R2099_U37, P2_R2099_U38, P2_R2099_U39, P2_R2099_U40, P2_R2099_U41, P2_R2099_U42, P2_R2099_U43, P2_R2099_U44, P2_R2099_U45, P2_R2099_U46, P2_R2099_U47, P2_R2099_U48, P2_R2099_U49, P2_R2099_U5, P2_R2099_U50, P2_R2099_U51, P2_R2099_U52, P2_R2099_U53, P2_R2099_U54, P2_R2099_U55, P2_R2099_U56, P2_R2099_U57, P2_R2099_U58, P2_R2099_U59, P2_R2099_U6, P2_R2099_U60, P2_R2099_U61, P2_R2099_U62, P2_R2099_U63, P2_R2099_U64, P2_R2099_U65, P2_R2099_U66, P2_R2099_U67, P2_R2099_U68, P2_R2099_U69, P2_R2099_U7, P2_R2099_U70, P2_R2099_U71, P2_R2099_U72, P2_R2099_U73, P2_R2099_U74, P2_R2099_U75, P2_R2099_U76, P2_R2099_U77, P2_R2099_U78, P2_R2099_U79, P2_R2099_U8, P2_R2099_U80, P2_R2099_U81, P2_R2099_U82, P2_R2099_U83, P2_R2099_U84, P2_R2099_U85, P2_R2099_U86, P2_R2099_U87, P2_R2099_U88, P2_R2099_U89, P2_R2099_U9, P2_R2099_U90, P2_R2099_U91, P2_R2099_U92, P2_R2099_U93, P2_R2099_U94, P2_R2099_U95, P2_R2099_U96, P2_R2099_U97, P2_R2099_U98, P2_R2099_U99, P2_R2147_U10, P2_R2147_U11, P2_R2147_U12, P2_R2147_U13, P2_R2147_U14, P2_R2147_U15, P2_R2147_U16, P2_R2147_U17, P2_R2147_U18, P2_R2147_U19, P2_R2147_U20, P2_R2147_U4, P2_R2147_U5, P2_R2147_U6, P2_R2147_U7, P2_R2147_U8, P2_R2147_U9, P2_R2167_U10, P2_R2167_U11, P2_R2167_U12, P2_R2167_U13, P2_R2167_U14, P2_R2167_U15, P2_R2167_U16, P2_R2167_U17, P2_R2167_U18, P2_R2167_U19, P2_R2167_U20, P2_R2167_U21, P2_R2167_U22, P2_R2167_U23, P2_R2167_U24, P2_R2167_U25, P2_R2167_U26, P2_R2167_U27, P2_R2167_U28, P2_R2167_U29, P2_R2167_U30, P2_R2167_U31, P2_R2167_U32, P2_R2167_U33, P2_R2167_U34, P2_R2167_U35, P2_R2167_U36, P2_R2167_U37, P2_R2167_U38, P2_R2167_U39, P2_R2167_U40, P2_R2167_U41, P2_R2167_U42, P2_R2167_U6, P2_R2167_U7, P2_R2167_U8, P2_R2167_U9, P2_R2182_U10, P2_R2182_U100, P2_R2182_U101, P2_R2182_U102, P2_R2182_U103, P2_R2182_U104, P2_R2182_U105, P2_R2182_U106, P2_R2182_U107, P2_R2182_U108, P2_R2182_U109, P2_R2182_U11, P2_R2182_U110, P2_R2182_U111, P2_R2182_U112, P2_R2182_U113, P2_R2182_U114, P2_R2182_U115, P2_R2182_U116, P2_R2182_U117, P2_R2182_U118, P2_R2182_U119, P2_R2182_U12, P2_R2182_U120, P2_R2182_U121, P2_R2182_U122, P2_R2182_U123, P2_R2182_U124, P2_R2182_U125, P2_R2182_U126, P2_R2182_U127, P2_R2182_U128, P2_R2182_U129, P2_R2182_U13, P2_R2182_U130, P2_R2182_U131, P2_R2182_U132, P2_R2182_U133, P2_R2182_U134, P2_R2182_U135, P2_R2182_U136, P2_R2182_U137, P2_R2182_U138, P2_R2182_U139, P2_R2182_U14, P2_R2182_U140, P2_R2182_U141, P2_R2182_U142, P2_R2182_U143, P2_R2182_U144, P2_R2182_U145, P2_R2182_U146, P2_R2182_U147, P2_R2182_U148, P2_R2182_U149, P2_R2182_U15, P2_R2182_U150, P2_R2182_U151, P2_R2182_U152, P2_R2182_U153, P2_R2182_U154, P2_R2182_U155, P2_R2182_U156, P2_R2182_U157, P2_R2182_U158, P2_R2182_U159, P2_R2182_U16, P2_R2182_U160, P2_R2182_U161, P2_R2182_U162, P2_R2182_U163, P2_R2182_U164, P2_R2182_U165, P2_R2182_U166, P2_R2182_U167, P2_R2182_U168, P2_R2182_U169, P2_R2182_U17, P2_R2182_U170, P2_R2182_U171, P2_R2182_U172, P2_R2182_U173, P2_R2182_U174, P2_R2182_U175, P2_R2182_U176, P2_R2182_U177, P2_R2182_U178, P2_R2182_U179, P2_R2182_U18, P2_R2182_U180, P2_R2182_U181, P2_R2182_U182, P2_R2182_U183, P2_R2182_U184, P2_R2182_U185, P2_R2182_U186, P2_R2182_U187, P2_R2182_U188, P2_R2182_U189, P2_R2182_U19, P2_R2182_U190, P2_R2182_U191, P2_R2182_U192, P2_R2182_U193, P2_R2182_U194, P2_R2182_U195, P2_R2182_U196, P2_R2182_U197, P2_R2182_U198, P2_R2182_U199, P2_R2182_U20, P2_R2182_U200, P2_R2182_U201, P2_R2182_U202, P2_R2182_U203, P2_R2182_U204, P2_R2182_U205, P2_R2182_U206, P2_R2182_U207, P2_R2182_U208, P2_R2182_U209, P2_R2182_U21, P2_R2182_U210, P2_R2182_U211, P2_R2182_U212, P2_R2182_U213, P2_R2182_U214, P2_R2182_U215, P2_R2182_U216, P2_R2182_U217, P2_R2182_U218, P2_R2182_U219, P2_R2182_U22, P2_R2182_U220, P2_R2182_U221, P2_R2182_U222, P2_R2182_U223, P2_R2182_U224, P2_R2182_U225, P2_R2182_U226, P2_R2182_U227, P2_R2182_U228, P2_R2182_U229, P2_R2182_U23, P2_R2182_U230, P2_R2182_U231, P2_R2182_U232, P2_R2182_U233, P2_R2182_U234, P2_R2182_U235, P2_R2182_U236, P2_R2182_U237, P2_R2182_U238, P2_R2182_U239, P2_R2182_U24, P2_R2182_U240, P2_R2182_U241, P2_R2182_U242, P2_R2182_U243, P2_R2182_U244, P2_R2182_U245, P2_R2182_U246, P2_R2182_U247, P2_R2182_U248, P2_R2182_U249, P2_R2182_U25, P2_R2182_U250, P2_R2182_U251, P2_R2182_U252, P2_R2182_U253, P2_R2182_U254, P2_R2182_U255, P2_R2182_U256, P2_R2182_U257, P2_R2182_U258, P2_R2182_U259, P2_R2182_U26, P2_R2182_U260, P2_R2182_U261, P2_R2182_U262, P2_R2182_U263, P2_R2182_U264, P2_R2182_U265, P2_R2182_U266, P2_R2182_U267, P2_R2182_U268, P2_R2182_U269, P2_R2182_U27, P2_R2182_U270, P2_R2182_U271, P2_R2182_U272, P2_R2182_U273, P2_R2182_U274, P2_R2182_U275, P2_R2182_U276, P2_R2182_U277, P2_R2182_U278, P2_R2182_U279, P2_R2182_U28, P2_R2182_U280, P2_R2182_U281, P2_R2182_U282, P2_R2182_U283, P2_R2182_U284, P2_R2182_U285, P2_R2182_U286, P2_R2182_U287, P2_R2182_U288, P2_R2182_U289, P2_R2182_U29, P2_R2182_U290, P2_R2182_U291, P2_R2182_U292, P2_R2182_U293, P2_R2182_U294, P2_R2182_U295, P2_R2182_U296, P2_R2182_U297, P2_R2182_U298, P2_R2182_U299, P2_R2182_U30, P2_R2182_U300, P2_R2182_U301, P2_R2182_U302, P2_R2182_U303, P2_R2182_U304, P2_R2182_U305, P2_R2182_U31, P2_R2182_U32, P2_R2182_U33, P2_R2182_U34, P2_R2182_U35, P2_R2182_U36, P2_R2182_U37, P2_R2182_U38, P2_R2182_U39, P2_R2182_U4, P2_R2182_U40, P2_R2182_U41, P2_R2182_U42, P2_R2182_U43, P2_R2182_U44, P2_R2182_U45, P2_R2182_U46, P2_R2182_U47, P2_R2182_U48, P2_R2182_U49, P2_R2182_U5, P2_R2182_U50, P2_R2182_U51, P2_R2182_U52, P2_R2182_U53, P2_R2182_U54, P2_R2182_U55, P2_R2182_U56, P2_R2182_U57, P2_R2182_U58, P2_R2182_U59, P2_R2182_U6, P2_R2182_U60, P2_R2182_U61, P2_R2182_U62, P2_R2182_U63, P2_R2182_U64, P2_R2182_U65, P2_R2182_U66, P2_R2182_U67, P2_R2182_U68, P2_R2182_U69, P2_R2182_U7, P2_R2182_U70, P2_R2182_U71, P2_R2182_U72, P2_R2182_U73, P2_R2182_U74, P2_R2182_U75, P2_R2182_U76, P2_R2182_U77, P2_R2182_U78, P2_R2182_U79, P2_R2182_U8, P2_R2182_U80, P2_R2182_U81, P2_R2182_U82, P2_R2182_U83, P2_R2182_U84, P2_R2182_U85, P2_R2182_U86, P2_R2182_U87, P2_R2182_U88, P2_R2182_U89, P2_R2182_U9, P2_R2182_U90, P2_R2182_U91, P2_R2182_U92, P2_R2182_U93, P2_R2182_U94, P2_R2182_U95, P2_R2182_U96, P2_R2182_U97, P2_R2182_U98, P2_R2182_U99, P2_R2219_U10, P2_R2219_U100, P2_R2219_U101, P2_R2219_U102, P2_R2219_U103, P2_R2219_U104, P2_R2219_U105, P2_R2219_U106, P2_R2219_U107, P2_R2219_U108, P2_R2219_U109, P2_R2219_U11, P2_R2219_U110, P2_R2219_U111, P2_R2219_U112, P2_R2219_U113, P2_R2219_U114, P2_R2219_U115, P2_R2219_U116, P2_R2219_U12, P2_R2219_U13, P2_R2219_U14, P2_R2219_U15, P2_R2219_U16, P2_R2219_U17, P2_R2219_U18, P2_R2219_U19, P2_R2219_U20, P2_R2219_U21, P2_R2219_U22, P2_R2219_U23, P2_R2219_U24, P2_R2219_U25, P2_R2219_U26, P2_R2219_U27, P2_R2219_U28, P2_R2219_U29, P2_R2219_U30, P2_R2219_U31, P2_R2219_U32, P2_R2219_U33, P2_R2219_U34, P2_R2219_U35, P2_R2219_U36, P2_R2219_U37, P2_R2219_U38, P2_R2219_U39, P2_R2219_U40, P2_R2219_U41, P2_R2219_U42, P2_R2219_U43, P2_R2219_U44, P2_R2219_U45, P2_R2219_U46, P2_R2219_U47, P2_R2219_U48, P2_R2219_U49, P2_R2219_U50, P2_R2219_U51, P2_R2219_U52, P2_R2219_U53, P2_R2219_U54, P2_R2219_U55, P2_R2219_U56, P2_R2219_U57, P2_R2219_U58, P2_R2219_U59, P2_R2219_U6, P2_R2219_U60, P2_R2219_U61, P2_R2219_U62, P2_R2219_U63, P2_R2219_U64, P2_R2219_U65, P2_R2219_U66, P2_R2219_U67, P2_R2219_U68, P2_R2219_U69, P2_R2219_U7, P2_R2219_U70, P2_R2219_U71, P2_R2219_U72, P2_R2219_U73, P2_R2219_U74, P2_R2219_U75, P2_R2219_U76, P2_R2219_U77, P2_R2219_U78, P2_R2219_U79, P2_R2219_U8, P2_R2219_U80, P2_R2219_U81, P2_R2219_U82, P2_R2219_U83, P2_R2219_U84, P2_R2219_U85, P2_R2219_U86, P2_R2219_U87, P2_R2219_U88, P2_R2219_U89, P2_R2219_U9, P2_R2219_U90, P2_R2219_U91, P2_R2219_U92, P2_R2219_U93, P2_R2219_U94, P2_R2219_U95, P2_R2219_U96, P2_R2219_U97, P2_R2219_U98, P2_R2219_U99, P2_R2238_U10, P2_R2238_U11, P2_R2238_U12, P2_R2238_U13, P2_R2238_U14, P2_R2238_U15, P2_R2238_U16, P2_R2238_U17, P2_R2238_U18, P2_R2238_U19, P2_R2238_U20, P2_R2238_U21, P2_R2238_U22, P2_R2238_U23, P2_R2238_U24, P2_R2238_U25, P2_R2238_U26, P2_R2238_U27, P2_R2238_U28, P2_R2238_U29, P2_R2238_U30, P2_R2238_U31, P2_R2238_U32, P2_R2238_U33, P2_R2238_U34, P2_R2238_U35, P2_R2238_U36, P2_R2238_U37, P2_R2238_U38, P2_R2238_U39, P2_R2238_U40, P2_R2238_U41, P2_R2238_U42, P2_R2238_U43, P2_R2238_U44, P2_R2238_U45, P2_R2238_U46, P2_R2238_U47, P2_R2238_U48, P2_R2238_U49, P2_R2238_U50, P2_R2238_U51, P2_R2238_U52, P2_R2238_U53, P2_R2238_U54, P2_R2238_U55, P2_R2238_U56, P2_R2238_U57, P2_R2238_U58, P2_R2238_U59, P2_R2238_U6, P2_R2238_U60, P2_R2238_U61, P2_R2238_U62, P2_R2238_U63, P2_R2238_U64, P2_R2238_U65, P2_R2238_U66, P2_R2238_U7, P2_R2238_U8, P2_R2238_U9, P2_R2243_U10, P2_R2243_U11, P2_R2243_U6, P2_R2243_U7, P2_R2243_U8, P2_R2243_U9, P2_R2256_U10, P2_R2256_U11, P2_R2256_U12, P2_R2256_U13, P2_R2256_U14, P2_R2256_U15, P2_R2256_U16, P2_R2256_U17, P2_R2256_U18, P2_R2256_U19, P2_R2256_U20, P2_R2256_U21, P2_R2256_U22, P2_R2256_U23, P2_R2256_U24, P2_R2256_U25, P2_R2256_U26, P2_R2256_U27, P2_R2256_U28, P2_R2256_U29, P2_R2256_U30, P2_R2256_U31, P2_R2256_U32, P2_R2256_U33, P2_R2256_U34, P2_R2256_U35, P2_R2256_U36, P2_R2256_U37, P2_R2256_U38, P2_R2256_U39, P2_R2256_U4, P2_R2256_U40, P2_R2256_U41, P2_R2256_U42, P2_R2256_U43, P2_R2256_U44, P2_R2256_U45, P2_R2256_U46, P2_R2256_U47, P2_R2256_U48, P2_R2256_U49, P2_R2256_U5, P2_R2256_U50, P2_R2256_U51, P2_R2256_U52, P2_R2256_U53, P2_R2256_U54, P2_R2256_U55, P2_R2256_U56, P2_R2256_U57, P2_R2256_U58, P2_R2256_U59, P2_R2256_U6, P2_R2256_U60, P2_R2256_U61, P2_R2256_U62, P2_R2256_U63, P2_R2256_U64, P2_R2256_U65, P2_R2256_U66, P2_R2256_U67, P2_R2256_U68, P2_R2256_U69, P2_R2256_U7, P2_R2256_U70, P2_R2256_U8, P2_R2256_U9, P2_R2267_U10, P2_R2267_U100, P2_R2267_U101, P2_R2267_U102, P2_R2267_U103, P2_R2267_U104, P2_R2267_U105, P2_R2267_U106, P2_R2267_U107, P2_R2267_U108, P2_R2267_U109, P2_R2267_U11, P2_R2267_U110, P2_R2267_U111, P2_R2267_U112, P2_R2267_U113, P2_R2267_U114, P2_R2267_U115, P2_R2267_U116, P2_R2267_U117, P2_R2267_U118, P2_R2267_U119, P2_R2267_U12, P2_R2267_U120, P2_R2267_U121, P2_R2267_U122, P2_R2267_U123, P2_R2267_U124, P2_R2267_U125, P2_R2267_U126, P2_R2267_U127, P2_R2267_U128, P2_R2267_U129, P2_R2267_U13, P2_R2267_U130, P2_R2267_U131, P2_R2267_U132, P2_R2267_U133, P2_R2267_U134, P2_R2267_U135, P2_R2267_U136, P2_R2267_U137, P2_R2267_U138, P2_R2267_U139, P2_R2267_U14, P2_R2267_U140, P2_R2267_U141, P2_R2267_U142, P2_R2267_U143, P2_R2267_U144, P2_R2267_U145, P2_R2267_U146, P2_R2267_U147, P2_R2267_U148, P2_R2267_U149, P2_R2267_U15, P2_R2267_U150, P2_R2267_U151, P2_R2267_U152, P2_R2267_U153, P2_R2267_U154, P2_R2267_U155, P2_R2267_U156, P2_R2267_U157, P2_R2267_U158, P2_R2267_U159, P2_R2267_U16, P2_R2267_U160, P2_R2267_U161, P2_R2267_U162, P2_R2267_U163, P2_R2267_U164, P2_R2267_U165, P2_R2267_U166, P2_R2267_U17, P2_R2267_U18, P2_R2267_U19, P2_R2267_U20, P2_R2267_U21, P2_R2267_U22, P2_R2267_U23, P2_R2267_U24, P2_R2267_U25, P2_R2267_U26, P2_R2267_U27, P2_R2267_U28, P2_R2267_U29, P2_R2267_U30, P2_R2267_U31, P2_R2267_U32, P2_R2267_U33, P2_R2267_U34, P2_R2267_U35, P2_R2267_U36, P2_R2267_U37, P2_R2267_U38, P2_R2267_U39, P2_R2267_U40, P2_R2267_U41, P2_R2267_U42, P2_R2267_U43, P2_R2267_U44, P2_R2267_U45, P2_R2267_U46, P2_R2267_U47, P2_R2267_U48, P2_R2267_U49, P2_R2267_U50, P2_R2267_U51, P2_R2267_U52, P2_R2267_U53, P2_R2267_U54, P2_R2267_U55, P2_R2267_U56, P2_R2267_U57, P2_R2267_U58, P2_R2267_U59, P2_R2267_U6, P2_R2267_U60, P2_R2267_U61, P2_R2267_U62, P2_R2267_U63, P2_R2267_U64, P2_R2267_U65, P2_R2267_U66, P2_R2267_U67, P2_R2267_U68, P2_R2267_U69, P2_R2267_U7, P2_R2267_U70, P2_R2267_U71, P2_R2267_U72, P2_R2267_U73, P2_R2267_U74, P2_R2267_U75, P2_R2267_U76, P2_R2267_U77, P2_R2267_U78, P2_R2267_U79, P2_R2267_U8, P2_R2267_U80, P2_R2267_U81, P2_R2267_U82, P2_R2267_U83, P2_R2267_U84, P2_R2267_U85, P2_R2267_U86, P2_R2267_U87, P2_R2267_U88, P2_R2267_U89, P2_R2267_U9, P2_R2267_U90, P2_R2267_U91, P2_R2267_U92, P2_R2267_U93, P2_R2267_U94, P2_R2267_U95, P2_R2267_U96, P2_R2267_U97, P2_R2267_U98, P2_R2267_U99, P2_R2278_U10, P2_R2278_U100, P2_R2278_U101, P2_R2278_U102, P2_R2278_U103, P2_R2278_U104, P2_R2278_U105, P2_R2278_U106, P2_R2278_U107, P2_R2278_U108, P2_R2278_U109, P2_R2278_U11, P2_R2278_U110, P2_R2278_U111, P2_R2278_U112, P2_R2278_U113, P2_R2278_U114, P2_R2278_U115, P2_R2278_U116, P2_R2278_U117, P2_R2278_U118, P2_R2278_U119, P2_R2278_U12, P2_R2278_U120, P2_R2278_U121, P2_R2278_U122, P2_R2278_U123, P2_R2278_U124, P2_R2278_U125, P2_R2278_U126, P2_R2278_U127, P2_R2278_U128, P2_R2278_U129, P2_R2278_U13, P2_R2278_U130, P2_R2278_U131, P2_R2278_U132, P2_R2278_U133, P2_R2278_U134, P2_R2278_U135, P2_R2278_U136, P2_R2278_U137, P2_R2278_U138, P2_R2278_U139, P2_R2278_U14, P2_R2278_U140, P2_R2278_U141, P2_R2278_U142, P2_R2278_U143, P2_R2278_U144, P2_R2278_U145, P2_R2278_U146, P2_R2278_U147, P2_R2278_U148, P2_R2278_U149, P2_R2278_U15, P2_R2278_U150, P2_R2278_U151, P2_R2278_U152, P2_R2278_U153, P2_R2278_U154, P2_R2278_U155, P2_R2278_U156, P2_R2278_U157, P2_R2278_U158, P2_R2278_U159, P2_R2278_U16, P2_R2278_U160, P2_R2278_U161, P2_R2278_U162, P2_R2278_U163, P2_R2278_U164, P2_R2278_U165, P2_R2278_U166, P2_R2278_U167, P2_R2278_U168, P2_R2278_U169, P2_R2278_U17, P2_R2278_U170, P2_R2278_U171, P2_R2278_U172, P2_R2278_U173, P2_R2278_U174, P2_R2278_U175, P2_R2278_U176, P2_R2278_U177, P2_R2278_U178, P2_R2278_U179, P2_R2278_U18, P2_R2278_U180, P2_R2278_U181, P2_R2278_U182, P2_R2278_U183, P2_R2278_U184, P2_R2278_U185, P2_R2278_U186, P2_R2278_U187, P2_R2278_U188, P2_R2278_U189, P2_R2278_U19, P2_R2278_U190, P2_R2278_U191, P2_R2278_U192, P2_R2278_U193, P2_R2278_U194, P2_R2278_U195, P2_R2278_U196, P2_R2278_U197, P2_R2278_U198, P2_R2278_U199, P2_R2278_U20, P2_R2278_U200, P2_R2278_U201, P2_R2278_U202, P2_R2278_U203, P2_R2278_U204, P2_R2278_U205, P2_R2278_U206, P2_R2278_U207, P2_R2278_U208, P2_R2278_U209, P2_R2278_U21, P2_R2278_U210, P2_R2278_U211, P2_R2278_U212, P2_R2278_U213, P2_R2278_U214, P2_R2278_U215, P2_R2278_U216, P2_R2278_U217, P2_R2278_U218, P2_R2278_U219, P2_R2278_U22, P2_R2278_U220, P2_R2278_U221, P2_R2278_U222, P2_R2278_U223, P2_R2278_U224, P2_R2278_U225, P2_R2278_U226, P2_R2278_U227, P2_R2278_U228, P2_R2278_U229, P2_R2278_U23, P2_R2278_U230, P2_R2278_U231, P2_R2278_U232, P2_R2278_U233, P2_R2278_U234, P2_R2278_U235, P2_R2278_U236, P2_R2278_U237, P2_R2278_U238, P2_R2278_U239, P2_R2278_U24, P2_R2278_U240, P2_R2278_U241, P2_R2278_U242, P2_R2278_U243, P2_R2278_U244, P2_R2278_U245, P2_R2278_U246, P2_R2278_U247, P2_R2278_U248, P2_R2278_U249, P2_R2278_U25, P2_R2278_U250, P2_R2278_U251, P2_R2278_U252, P2_R2278_U253, P2_R2278_U254, P2_R2278_U255, P2_R2278_U256, P2_R2278_U257, P2_R2278_U258, P2_R2278_U259, P2_R2278_U26, P2_R2278_U260, P2_R2278_U261, P2_R2278_U262, P2_R2278_U263, P2_R2278_U264, P2_R2278_U265, P2_R2278_U266, P2_R2278_U267, P2_R2278_U268, P2_R2278_U269, P2_R2278_U27, P2_R2278_U270, P2_R2278_U271, P2_R2278_U272, P2_R2278_U273, P2_R2278_U274, P2_R2278_U275, P2_R2278_U276, P2_R2278_U277, P2_R2278_U278, P2_R2278_U279, P2_R2278_U28, P2_R2278_U280, P2_R2278_U281, P2_R2278_U282, P2_R2278_U283, P2_R2278_U284, P2_R2278_U285, P2_R2278_U286, P2_R2278_U287, P2_R2278_U288, P2_R2278_U289, P2_R2278_U29, P2_R2278_U290, P2_R2278_U291, P2_R2278_U292, P2_R2278_U293, P2_R2278_U294, P2_R2278_U295, P2_R2278_U296, P2_R2278_U297, P2_R2278_U298, P2_R2278_U299, P2_R2278_U30, P2_R2278_U300, P2_R2278_U301, P2_R2278_U302, P2_R2278_U303, P2_R2278_U304, P2_R2278_U305, P2_R2278_U306, P2_R2278_U307, P2_R2278_U308, P2_R2278_U309, P2_R2278_U31, P2_R2278_U310, P2_R2278_U311, P2_R2278_U312, P2_R2278_U313, P2_R2278_U314, P2_R2278_U315, P2_R2278_U316, P2_R2278_U317, P2_R2278_U318, P2_R2278_U319, P2_R2278_U32, P2_R2278_U320, P2_R2278_U321, P2_R2278_U322, P2_R2278_U323, P2_R2278_U324, P2_R2278_U325, P2_R2278_U326, P2_R2278_U327, P2_R2278_U328, P2_R2278_U329, P2_R2278_U33, P2_R2278_U330, P2_R2278_U331, P2_R2278_U332, P2_R2278_U333, P2_R2278_U334, P2_R2278_U335, P2_R2278_U336, P2_R2278_U337, P2_R2278_U338, P2_R2278_U339, P2_R2278_U34, P2_R2278_U340, P2_R2278_U341, P2_R2278_U342, P2_R2278_U343, P2_R2278_U344, P2_R2278_U345, P2_R2278_U346, P2_R2278_U347, P2_R2278_U348, P2_R2278_U349, P2_R2278_U35, P2_R2278_U350, P2_R2278_U351, P2_R2278_U352, P2_R2278_U353, P2_R2278_U354, P2_R2278_U355, P2_R2278_U356, P2_R2278_U357, P2_R2278_U358, P2_R2278_U359, P2_R2278_U36, P2_R2278_U360, P2_R2278_U361, P2_R2278_U362, P2_R2278_U363, P2_R2278_U364, P2_R2278_U365, P2_R2278_U366, P2_R2278_U367, P2_R2278_U368, P2_R2278_U369, P2_R2278_U37, P2_R2278_U370, P2_R2278_U371, P2_R2278_U372, P2_R2278_U373, P2_R2278_U374, P2_R2278_U375, P2_R2278_U376, P2_R2278_U377, P2_R2278_U378, P2_R2278_U379, P2_R2278_U38, P2_R2278_U380, P2_R2278_U381, P2_R2278_U382, P2_R2278_U383, P2_R2278_U384, P2_R2278_U385, P2_R2278_U386, P2_R2278_U387, P2_R2278_U388, P2_R2278_U389, P2_R2278_U39, P2_R2278_U390, P2_R2278_U391, P2_R2278_U392, P2_R2278_U393, P2_R2278_U394, P2_R2278_U395, P2_R2278_U396, P2_R2278_U397, P2_R2278_U398, P2_R2278_U399, P2_R2278_U4, P2_R2278_U40, P2_R2278_U400, P2_R2278_U401, P2_R2278_U402, P2_R2278_U403, P2_R2278_U404, P2_R2278_U405, P2_R2278_U406, P2_R2278_U407, P2_R2278_U408, P2_R2278_U409, P2_R2278_U41, P2_R2278_U410, P2_R2278_U411, P2_R2278_U412, P2_R2278_U413, P2_R2278_U414, P2_R2278_U415, P2_R2278_U416, P2_R2278_U417, P2_R2278_U418, P2_R2278_U419, P2_R2278_U42, P2_R2278_U420, P2_R2278_U421, P2_R2278_U422, P2_R2278_U423, P2_R2278_U424, P2_R2278_U425, P2_R2278_U426, P2_R2278_U427, P2_R2278_U428, P2_R2278_U429, P2_R2278_U43, P2_R2278_U430, P2_R2278_U431, P2_R2278_U432, P2_R2278_U433, P2_R2278_U434, P2_R2278_U435, P2_R2278_U436, P2_R2278_U437, P2_R2278_U438, P2_R2278_U439, P2_R2278_U44, P2_R2278_U440, P2_R2278_U441, P2_R2278_U442, P2_R2278_U443, P2_R2278_U444, P2_R2278_U445, P2_R2278_U446, P2_R2278_U447, P2_R2278_U448, P2_R2278_U449, P2_R2278_U45, P2_R2278_U450, P2_R2278_U451, P2_R2278_U452, P2_R2278_U453, P2_R2278_U454, P2_R2278_U455, P2_R2278_U456, P2_R2278_U457, P2_R2278_U458, P2_R2278_U459, P2_R2278_U46, P2_R2278_U460, P2_R2278_U461, P2_R2278_U462, P2_R2278_U463, P2_R2278_U464, P2_R2278_U465, P2_R2278_U466, P2_R2278_U467, P2_R2278_U468, P2_R2278_U469, P2_R2278_U47, P2_R2278_U470, P2_R2278_U471, P2_R2278_U472, P2_R2278_U473, P2_R2278_U474, P2_R2278_U475, P2_R2278_U476, P2_R2278_U477, P2_R2278_U478, P2_R2278_U479, P2_R2278_U48, P2_R2278_U480, P2_R2278_U481, P2_R2278_U482, P2_R2278_U483, P2_R2278_U484, P2_R2278_U485, P2_R2278_U486, P2_R2278_U487, P2_R2278_U488, P2_R2278_U489, P2_R2278_U49, P2_R2278_U490, P2_R2278_U491, P2_R2278_U492, P2_R2278_U493, P2_R2278_U494, P2_R2278_U495, P2_R2278_U496, P2_R2278_U497, P2_R2278_U498, P2_R2278_U499, P2_R2278_U5, P2_R2278_U50, P2_R2278_U500, P2_R2278_U501, P2_R2278_U502, P2_R2278_U503, P2_R2278_U504, P2_R2278_U505, P2_R2278_U506, P2_R2278_U507, P2_R2278_U508, P2_R2278_U509, P2_R2278_U51, P2_R2278_U510, P2_R2278_U511, P2_R2278_U512, P2_R2278_U513, P2_R2278_U514, P2_R2278_U515, P2_R2278_U516, P2_R2278_U517, P2_R2278_U518, P2_R2278_U519, P2_R2278_U52, P2_R2278_U520, P2_R2278_U521, P2_R2278_U522, P2_R2278_U523, P2_R2278_U524, P2_R2278_U525, P2_R2278_U526, P2_R2278_U527, P2_R2278_U528, P2_R2278_U529, P2_R2278_U53, P2_R2278_U530, P2_R2278_U531, P2_R2278_U532, P2_R2278_U533, P2_R2278_U534, P2_R2278_U535, P2_R2278_U536, P2_R2278_U537, P2_R2278_U538, P2_R2278_U539, P2_R2278_U54, P2_R2278_U540, P2_R2278_U541, P2_R2278_U542, P2_R2278_U543, P2_R2278_U544, P2_R2278_U545, P2_R2278_U546, P2_R2278_U547, P2_R2278_U548, P2_R2278_U549, P2_R2278_U55, P2_R2278_U550, P2_R2278_U551, P2_R2278_U552, P2_R2278_U553, P2_R2278_U554, P2_R2278_U555, P2_R2278_U556, P2_R2278_U557, P2_R2278_U558, P2_R2278_U559, P2_R2278_U56, P2_R2278_U560, P2_R2278_U561, P2_R2278_U562, P2_R2278_U57, P2_R2278_U58, P2_R2278_U59, P2_R2278_U6, P2_R2278_U60, P2_R2278_U61, P2_R2278_U62, P2_R2278_U63, P2_R2278_U64, P2_R2278_U65, P2_R2278_U66, P2_R2278_U67, P2_R2278_U68, P2_R2278_U69, P2_R2278_U7, P2_R2278_U70, P2_R2278_U71, P2_R2278_U72, P2_R2278_U73, P2_R2278_U74, P2_R2278_U75, P2_R2278_U76, P2_R2278_U77, P2_R2278_U78, P2_R2278_U79, P2_R2278_U8, P2_R2278_U80, P2_R2278_U81, P2_R2278_U82, P2_R2278_U83, P2_R2278_U84, P2_R2278_U85, P2_R2278_U86, P2_R2278_U87, P2_R2278_U88, P2_R2278_U89, P2_R2278_U9, P2_R2278_U90, P2_R2278_U91, P2_R2278_U92, P2_R2278_U93, P2_R2278_U94, P2_R2278_U95, P2_R2278_U96, P2_R2278_U97, P2_R2278_U98, P2_R2278_U99, P2_R2337_U10, P2_R2337_U100, P2_R2337_U101, P2_R2337_U102, P2_R2337_U103, P2_R2337_U104, P2_R2337_U105, P2_R2337_U106, P2_R2337_U107, P2_R2337_U108, P2_R2337_U109, P2_R2337_U11, P2_R2337_U110, P2_R2337_U111, P2_R2337_U112, P2_R2337_U113, P2_R2337_U114, P2_R2337_U115, P2_R2337_U116, P2_R2337_U117, P2_R2337_U118, P2_R2337_U119, P2_R2337_U12, P2_R2337_U120, P2_R2337_U121, P2_R2337_U122, P2_R2337_U123, P2_R2337_U124, P2_R2337_U125, P2_R2337_U126, P2_R2337_U127, P2_R2337_U128, P2_R2337_U129, P2_R2337_U13, P2_R2337_U130, P2_R2337_U131, P2_R2337_U132, P2_R2337_U133, P2_R2337_U134, P2_R2337_U135, P2_R2337_U136, P2_R2337_U137, P2_R2337_U138, P2_R2337_U139, P2_R2337_U14, P2_R2337_U140, P2_R2337_U141, P2_R2337_U142, P2_R2337_U143, P2_R2337_U144, P2_R2337_U145, P2_R2337_U146, P2_R2337_U147, P2_R2337_U148, P2_R2337_U149, P2_R2337_U15, P2_R2337_U150, P2_R2337_U151, P2_R2337_U152, P2_R2337_U153, P2_R2337_U154, P2_R2337_U155, P2_R2337_U156, P2_R2337_U157, P2_R2337_U158, P2_R2337_U159, P2_R2337_U16, P2_R2337_U160, P2_R2337_U161, P2_R2337_U162, P2_R2337_U163, P2_R2337_U164, P2_R2337_U165, P2_R2337_U166, P2_R2337_U167, P2_R2337_U168, P2_R2337_U169, P2_R2337_U17, P2_R2337_U170, P2_R2337_U171, P2_R2337_U172, P2_R2337_U173, P2_R2337_U174, P2_R2337_U175, P2_R2337_U176, P2_R2337_U177, P2_R2337_U178, P2_R2337_U179, P2_R2337_U18, P2_R2337_U180, P2_R2337_U181, P2_R2337_U182, P2_R2337_U19, P2_R2337_U20, P2_R2337_U21, P2_R2337_U22, P2_R2337_U23, P2_R2337_U24, P2_R2337_U25, P2_R2337_U26, P2_R2337_U27, P2_R2337_U28, P2_R2337_U29, P2_R2337_U30, P2_R2337_U31, P2_R2337_U32, P2_R2337_U33, P2_R2337_U34, P2_R2337_U35, P2_R2337_U36, P2_R2337_U37, P2_R2337_U38, P2_R2337_U39, P2_R2337_U4, P2_R2337_U40, P2_R2337_U41, P2_R2337_U42, P2_R2337_U43, P2_R2337_U44, P2_R2337_U45, P2_R2337_U46, P2_R2337_U47, P2_R2337_U48, P2_R2337_U49, P2_R2337_U5, P2_R2337_U50, P2_R2337_U51, P2_R2337_U52, P2_R2337_U53, P2_R2337_U54, P2_R2337_U55, P2_R2337_U56, P2_R2337_U57, P2_R2337_U58, P2_R2337_U59, P2_R2337_U6, P2_R2337_U60, P2_R2337_U61, P2_R2337_U62, P2_R2337_U63, P2_R2337_U64, P2_R2337_U65, P2_R2337_U66, P2_R2337_U67, P2_R2337_U68, P2_R2337_U69, P2_R2337_U7, P2_R2337_U70, P2_R2337_U71, P2_R2337_U72, P2_R2337_U73, P2_R2337_U74, P2_R2337_U75, P2_R2337_U76, P2_R2337_U77, P2_R2337_U78, P2_R2337_U79, P2_R2337_U8, P2_R2337_U80, P2_R2337_U81, P2_R2337_U82, P2_R2337_U83, P2_R2337_U84, P2_R2337_U85, P2_R2337_U86, P2_R2337_U87, P2_R2337_U88, P2_R2337_U89, P2_R2337_U9, P2_R2337_U90, P2_R2337_U91, P2_R2337_U92, P2_R2337_U93, P2_R2337_U94, P2_R2337_U95, P2_R2337_U96, P2_R2337_U97, P2_R2337_U98, P2_R2337_U99, P2_SUB_450_U10, P2_SUB_450_U11, P2_SUB_450_U12, P2_SUB_450_U13, P2_SUB_450_U14, P2_SUB_450_U15, P2_SUB_450_U16, P2_SUB_450_U17, P2_SUB_450_U18, P2_SUB_450_U19, P2_SUB_450_U20, P2_SUB_450_U21, P2_SUB_450_U22, P2_SUB_450_U23, P2_SUB_450_U24, P2_SUB_450_U25, P2_SUB_450_U26, P2_SUB_450_U27, P2_SUB_450_U28, P2_SUB_450_U29, P2_SUB_450_U30, P2_SUB_450_U31, P2_SUB_450_U32, P2_SUB_450_U33, P2_SUB_450_U34, P2_SUB_450_U35, P2_SUB_450_U36, P2_SUB_450_U37, P2_SUB_450_U38, P2_SUB_450_U39, P2_SUB_450_U40, P2_SUB_450_U41, P2_SUB_450_U42, P2_SUB_450_U43, P2_SUB_450_U44, P2_SUB_450_U45, P2_SUB_450_U46, P2_SUB_450_U47, P2_SUB_450_U48, P2_SUB_450_U49, P2_SUB_450_U50, P2_SUB_450_U51, P2_SUB_450_U52, P2_SUB_450_U53, P2_SUB_450_U54, P2_SUB_450_U55, P2_SUB_450_U56, P2_SUB_450_U57, P2_SUB_450_U58, P2_SUB_450_U59, P2_SUB_450_U6, P2_SUB_450_U60, P2_SUB_450_U61, P2_SUB_450_U62, P2_SUB_450_U63, P2_SUB_450_U7, P2_SUB_450_U8, P2_SUB_450_U9, P2_SUB_563_U6, P2_SUB_563_U7, P2_SUB_589_U6, P2_SUB_589_U7, P2_SUB_589_U8, P2_SUB_589_U9, P2_U2352, P2_U2353, P2_U2354, P2_U2355, P2_U2356, P2_U2357, P2_U2358, P2_U2359, P2_U2360, P2_U2361, P2_U2362, P2_U2363, P2_U2364, P2_U2365, P2_U2366, P2_U2367, P2_U2368, P2_U2369, P2_U2370, P2_U2371, P2_U2372, P2_U2373, P2_U2374, P2_U2375, P2_U2376, P2_U2377, P2_U2378, P2_U2379, P2_U2380, P2_U2381, P2_U2382, P2_U2383, P2_U2384, P2_U2385, P2_U2386, P2_U2387, P2_U2388, P2_U2389, P2_U2390, P2_U2391, P2_U2392, P2_U2393, P2_U2394, P2_U2395, P2_U2396, P2_U2397, P2_U2398, P2_U2399, P2_U2400, P2_U2401, P2_U2402, P2_U2403, P2_U2404, P2_U2405, P2_U2406, P2_U2407, P2_U2408, P2_U2409, P2_U2410, P2_U2411, P2_U2412, P2_U2413, P2_U2414, P2_U2415, P2_U2416, P2_U2417, P2_U2418, P2_U2419, P2_U2420, P2_U2421, P2_U2422, P2_U2423, P2_U2424, P2_U2425, P2_U2426, P2_U2427, P2_U2428, P2_U2429, P2_U2430, P2_U2431, P2_U2432, P2_U2433, P2_U2434, P2_U2435, P2_U2436, P2_U2437, P2_U2438, P2_U2439, P2_U2440, P2_U2441, P2_U2442, P2_U2443, P2_U2444, P2_U2445, P2_U2446, P2_U2447, P2_U2448, P2_U2449, P2_U2450, P2_U2451, P2_U2452, P2_U2453, P2_U2454, P2_U2455, P2_U2456, P2_U2457, P2_U2458, P2_U2459, P2_U2460, P2_U2461, P2_U2462, P2_U2463, P2_U2464, P2_U2465, P2_U2466, P2_U2467, P2_U2468, P2_U2469, P2_U2470, P2_U2471, P2_U2472, P2_U2473, P2_U2474, P2_U2475, P2_U2476, P2_U2477, P2_U2478, P2_U2479, P2_U2480, P2_U2481, P2_U2482, P2_U2483, P2_U2484, P2_U2485, P2_U2486, P2_U2487, P2_U2488, P2_U2489, P2_U2490, P2_U2491, P2_U2492, P2_U2493, P2_U2494, P2_U2495, P2_U2496, P2_U2497, P2_U2498, P2_U2499, P2_U2500, P2_U2501, P2_U2502, P2_U2503, P2_U2504, P2_U2505, P2_U2506, P2_U2507, P2_U2508, P2_U2509, P2_U2510, P2_U2511, P2_U2512, P2_U2513, P2_U2514, P2_U2515, P2_U2516, P2_U2517, P2_U2518, P2_U2519, P2_U2520, P2_U2521, P2_U2522, P2_U2523, P2_U2524, P2_U2525, P2_U2526, P2_U2527, P2_U2528, P2_U2529, P2_U2530, P2_U2531, P2_U2532, P2_U2533, P2_U2534, P2_U2535, P2_U2536, P2_U2537, P2_U2538, P2_U2539, P2_U2540, P2_U2541, P2_U2542, P2_U2543, P2_U2544, P2_U2545, P2_U2546, P2_U2547, P2_U2548, P2_U2549, P2_U2550, P2_U2551, P2_U2552, P2_U2553, P2_U2554, P2_U2555, P2_U2556, P2_U2557, P2_U2558, P2_U2559, P2_U2560, P2_U2561, P2_U2562, P2_U2563, P2_U2564, P2_U2565, P2_U2566, P2_U2567, P2_U2568, P2_U2569, P2_U2570, P2_U2571, P2_U2572, P2_U2573, P2_U2574, P2_U2575, P2_U2576, P2_U2577, P2_U2578, P2_U2579, P2_U2580, P2_U2581, P2_U2582, P2_U2583, P2_U2584, P2_U2585, P2_U2586, P2_U2587, P2_U2588, P2_U2589, P2_U2590, P2_U2591, P2_U2592, P2_U2593, P2_U2594, P2_U2595, P2_U2596, P2_U2597, P2_U2598, P2_U2599, P2_U2600, P2_U2601, P2_U2602, P2_U2603, P2_U2604, P2_U2605, P2_U2606, P2_U2607, P2_U2608, P2_U2609, P2_U2610, P2_U2611, P2_U2612, P2_U2613, P2_U2614, P2_U2615, P2_U2616, P2_U2617, P2_U2618, P2_U2619, P2_U2620, P2_U2621, P2_U2622, P2_U2623, P2_U2624, P2_U2625, P2_U2626, P2_U2627, P2_U2628, P2_U2629, P2_U2630, P2_U2631, P2_U2632, P2_U2633, P2_U2634, P2_U2635, P2_U2636, P2_U2637, P2_U2638, P2_U2639, P2_U2640, P2_U2641, P2_U2642, P2_U2643, P2_U2644, P2_U2645, P2_U2646, P2_U2647, P2_U2648, P2_U2649, P2_U2650, P2_U2651, P2_U2652, P2_U2653, P2_U2654, P2_U2655, P2_U2656, P2_U2657, P2_U2658, P2_U2659, P2_U2660, P2_U2661, P2_U2662, P2_U2663, P2_U2664, P2_U2665, P2_U2666, P2_U2667, P2_U2668, P2_U2669, P2_U2670, P2_U2671, P2_U2672, P2_U2673, P2_U2674, P2_U2675, P2_U2676, P2_U2677, P2_U2678, P2_U2679, P2_U2680, P2_U2681, P2_U2682, P2_U2683, P2_U2684, P2_U2685, P2_U2686, P2_U2687, P2_U2688, P2_U2689, P2_U2690, P2_U2691, P2_U2692, P2_U2693, P2_U2694, P2_U2695, P2_U2696, P2_U2698, P2_U2699, P2_U2700, P2_U2701, P2_U2702, P2_U2703, P2_U2704, P2_U2705, P2_U2706, P2_U2707, P2_U2708, P2_U2709, P2_U2710, P2_U2711, P2_U2712, P2_U2713, P2_U2714, P2_U2715, P2_U2716, P2_U2717, P2_U2718, P2_U2719, P2_U2720, P2_U2721, P2_U2722, P2_U2723, P2_U2724, P2_U2725, P2_U2726, P2_U2727, P2_U2728, P2_U2729, P2_U2730, P2_U2731, P2_U2732, P2_U2733, P2_U2734, P2_U2735, P2_U2736, P2_U2737, P2_U2738, P2_U2739, P2_U2740, P2_U2741, P2_U2742, P2_U2743, P2_U2744, P2_U2745, P2_U2746, P2_U2747, P2_U2748, P2_U2749, P2_U2750, P2_U2751, P2_U2752, P2_U2753, P2_U2754, P2_U2755, P2_U2756, P2_U2757, P2_U2758, P2_U2759, P2_U2760, P2_U2761, P2_U2762, P2_U2763, P2_U2764, P2_U2765, P2_U2766, P2_U2767, P2_U2768, P2_U2769, P2_U2770, P2_U2771, P2_U2772, P2_U2773, P2_U2774, P2_U2775, P2_U2776, P2_U2777, P2_U2778, P2_U2779, P2_U2780, P2_U2781, P2_U2782, P2_U2783, P2_U2784, P2_U2785, P2_U2786, P2_U2787, P2_U2788, P2_U2789, P2_U2790, P2_U2791, P2_U2792, P2_U2793, P2_U2794, P2_U2795, P2_U2796, P2_U2797, P2_U2798, P2_U2799, P2_U2800, P2_U2801, P2_U2802, P2_U2803, P2_U2804, P2_U2805, P2_U2806, P2_U2807, P2_U2808, P2_U2809, P2_U2810, P2_U2811, P2_U2812, P2_U2813, P2_U3242, P2_U3243, P2_U3244, P2_U3245, P2_U3246, P2_U3247, P2_U3248, P2_U3249, P2_U3250, P2_U3251, P2_U3252, P2_U3253, P2_U3254, P2_U3255, P2_U3256, P2_U3257, P2_U3258, P2_U3259, P2_U3260, P2_U3261, P2_U3262, P2_U3263, P2_U3264, P2_U3265, P2_U3266, P2_U3267, P2_U3268, P2_U3269, P2_U3270, P2_U3271, P2_U3272, P2_U3273, P2_U3274, P2_U3275, P2_U3276, P2_U3277, P2_U3278, P2_U3279, P2_U3280, P2_U3281, P2_U3282, P2_U3283, P2_U3284, P2_U3285, P2_U3286, P2_U3287, P2_U3288, P2_U3289, P2_U3290, P2_U3291, P2_U3292, P2_U3293, P2_U3294, P2_U3295, P2_U3296, P2_U3297, P2_U3298, P2_U3299, P2_U3300, P2_U3301, P2_U3302, P2_U3303, P2_U3304, P2_U3305, P2_U3306, P2_U3307, P2_U3308, P2_U3309, P2_U3310, P2_U3311, P2_U3312, P2_U3313, P2_U3314, P2_U3315, P2_U3316, P2_U3317, P2_U3318, P2_U3319, P2_U3320, P2_U3321, P2_U3322, P2_U3323, P2_U3324, P2_U3325, P2_U3326, P2_U3327, P2_U3328, P2_U3329, P2_U3330, P2_U3331, P2_U3332, P2_U3333, P2_U3334, P2_U3335, P2_U3336, P2_U3337, P2_U3338, P2_U3339, P2_U3340, P2_U3341, P2_U3342, P2_U3343, P2_U3344, P2_U3345, P2_U3346, P2_U3347, P2_U3348, P2_U3349, P2_U3350, P2_U3351, P2_U3352, P2_U3353, P2_U3354, P2_U3355, P2_U3356, P2_U3357, P2_U3358, P2_U3359, P2_U3360, P2_U3361, P2_U3362, P2_U3363, P2_U3364, P2_U3365, P2_U3366, P2_U3367, P2_U3368, P2_U3369, P2_U3370, P2_U3371, P2_U3372, P2_U3373, P2_U3374, P2_U3375, P2_U3376, P2_U3377, P2_U3378, P2_U3379, P2_U3380, P2_U3381, P2_U3382, P2_U3383, P2_U3384, P2_U3385, P2_U3386, P2_U3387, P2_U3388, P2_U3389, P2_U3390, P2_U3391, P2_U3392, P2_U3393, P2_U3394, P2_U3395, P2_U3396, P2_U3397, P2_U3398, P2_U3399, P2_U3400, P2_U3401, P2_U3402, P2_U3403, P2_U3404, P2_U3405, P2_U3406, P2_U3407, P2_U3408, P2_U3409, P2_U3410, P2_U3411, P2_U3412, P2_U3413, P2_U3414, P2_U3415, P2_U3416, P2_U3417, P2_U3418, P2_U3419, P2_U3420, P2_U3421, P2_U3422, P2_U3423, P2_U3424, P2_U3425, P2_U3426, P2_U3427, P2_U3428, P2_U3429, P2_U3430, P2_U3431, P2_U3432, P2_U3433, P2_U3434, P2_U3435, P2_U3436, P2_U3437, P2_U3438, P2_U3439, P2_U3440, P2_U3441, P2_U3442, P2_U3443, P2_U3444, P2_U3445, P2_U3446, P2_U3447, P2_U3448, P2_U3449, P2_U3450, P2_U3451, P2_U3452, P2_U3453, P2_U3454, P2_U3455, P2_U3456, P2_U3457, P2_U3458, P2_U3459, P2_U3460, P2_U3461, P2_U3462, P2_U3463, P2_U3464, P2_U3465, P2_U3466, P2_U3467, P2_U3468, P2_U3469, P2_U3470, P2_U3471, P2_U3472, P2_U3473, P2_U3474, P2_U3475, P2_U3476, P2_U3477, P2_U3478, P2_U3479, P2_U3480, P2_U3481, P2_U3482, P2_U3483, P2_U3484, P2_U3485, P2_U3486, P2_U3487, P2_U3488, P2_U3489, P2_U3490, P2_U3491, P2_U3492, P2_U3493, P2_U3494, P2_U3495, P2_U3496, P2_U3497, P2_U3498, P2_U3499, P2_U3500, P2_U3501, P2_U3502, P2_U3503, P2_U3504, P2_U3505, P2_U3506, P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511, P2_U3512, P2_U3513, P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518, P2_U3519, P2_U3520, P2_U3521, P2_U3522, P2_U3523, P2_U3524, P2_U3525, P2_U3526, P2_U3527, P2_U3528, P2_U3529, P2_U3530, P2_U3531, P2_U3532, P2_U3533, P2_U3534, P2_U3535, P2_U3536, P2_U3537, P2_U3538, P2_U3539, P2_U3540, P2_U3541, P2_U3542, P2_U3543, P2_U3544, P2_U3545, P2_U3546, P2_U3547, P2_U3548, P2_U3549, P2_U3550, P2_U3551, P2_U3552, P2_U3553, P2_U3554, P2_U3555, P2_U3556, P2_U3557, P2_U3558, P2_U3559, P2_U3560, P2_U3561, P2_U3562, P2_U3563, P2_U3564, P2_U3565, P2_U3566, P2_U3567, P2_U3568, P2_U3569, P2_U3570, P2_U3571, P2_U3572, P2_U3573, P2_U3574, P2_U3575, P2_U3576, P2_U3577, P2_U3578, P2_U3579, P2_U3580, P2_U3581, P2_U3582, P2_U3583, P2_U3584, P2_U3589, P2_U3590, P2_U3594, P2_U3597, P2_U3598, P2_U3606, P2_U3607, P2_U3613, P2_U3614, P2_U3615, P2_U3616, P2_U3617, P2_U3618, P2_U3619, P2_U3620, P2_U3621, P2_U3622, P2_U3623, P2_U3624, P2_U3625, P2_U3626, P2_U3627, P2_U3628, P2_U3629, P2_U3630, P2_U3631, P2_U3632, P2_U3633, P2_U3634, P2_U3635, P2_U3636, P2_U3637, P2_U3638, P2_U3639, P2_U3640, P2_U3641, P2_U3642, P2_U3643, P2_U3644, P2_U3645, P2_U3646, P2_U3647, P2_U3648, P2_U3649, P2_U3650, P2_U3651, P2_U3652, P2_U3653, P2_U3654, P2_U3655, P2_U3656, P2_U3657, P2_U3658, P2_U3659, P2_U3660, P2_U3661, P2_U3662, P2_U3663, P2_U3664, P2_U3665, P2_U3666, P2_U3667, P2_U3668, P2_U3669, P2_U3670, P2_U3671, P2_U3672, P2_U3673, P2_U3674, P2_U3675, P2_U3676, P2_U3677, P2_U3678, P2_U3679, P2_U3680, P2_U3681, P2_U3682, P2_U3683, P2_U3684, P2_U3685, P2_U3686, P2_U3687, P2_U3688, P2_U3689, P2_U3690, P2_U3691, P2_U3692, P2_U3693, P2_U3694, P2_U3695, P2_U3696, P2_U3697, P2_U3698, P2_U3699, P2_U3700, P2_U3701, P2_U3702, P2_U3703, P2_U3704, P2_U3705, P2_U3706, P2_U3707, P2_U3708, P2_U3709, P2_U3710, P2_U3711, P2_U3712, P2_U3713, P2_U3714, P2_U3715, P2_U3716, P2_U3717, P2_U3718, P2_U3719, P2_U3720, P2_U3721, P2_U3722, P2_U3723, P2_U3724, P2_U3725, P2_U3726, P2_U3727, P2_U3728, P2_U3729, P2_U3730, P2_U3731, P2_U3732, P2_U3733, P2_U3734, P2_U3735, P2_U3736, P2_U3737, P2_U3738, P2_U3739, P2_U3740, P2_U3741, P2_U3742, P2_U3743, P2_U3744, P2_U3745, P2_U3746, P2_U3747, P2_U3748, P2_U3749, P2_U3750, P2_U3751, P2_U3752, P2_U3753, P2_U3754, P2_U3755, P2_U3756, P2_U3757, P2_U3758, P2_U3759, P2_U3760, P2_U3761, P2_U3762, P2_U3763, P2_U3764, P2_U3765, P2_U3766, P2_U3767, P2_U3768, P2_U3769, P2_U3770, P2_U3771, P2_U3772, P2_U3773, P2_U3774, P2_U3775, P2_U3776, P2_U3777, P2_U3778, P2_U3779, P2_U3780, P2_U3781, P2_U3782, P2_U3783, P2_U3784, P2_U3785, P2_U3786, P2_U3787, P2_U3788, P2_U3789, P2_U3790, P2_U3791, P2_U3792, P2_U3793, P2_U3794, P2_U3795, P2_U3796, P2_U3797, P2_U3798, P2_U3799, P2_U3800, P2_U3801, P2_U3802, P2_U3803, P2_U3804, P2_U3805, P2_U3806, P2_U3807, P2_U3808, P2_U3809, P2_U3810, P2_U3811, P2_U3812, P2_U3813, P2_U3814, P2_U3815, P2_U3816, P2_U3817, P2_U3818, P2_U3819, P2_U3820, P2_U3821, P2_U3822, P2_U3823, P2_U3824, P2_U3825, P2_U3826, P2_U3827, P2_U3828, P2_U3829, P2_U3830, P2_U3831, P2_U3832, P2_U3833, P2_U3834, P2_U3835, P2_U3836, P2_U3837, P2_U3838, P2_U3839, P2_U3840, P2_U3841, P2_U3842, P2_U3843, P2_U3844, P2_U3845, P2_U3846, P2_U3847, P2_U3848, P2_U3849, P2_U3850, P2_U3851, P2_U3852, P2_U3853, P2_U3854, P2_U3855, P2_U3856, P2_U3857, P2_U3858, P2_U3859, P2_U3860, P2_U3861, P2_U3862, P2_U3863, P2_U3864, P2_U3865, P2_U3866, P2_U3867, P2_U3868, P2_U3869, P2_U3870, P2_U3871, P2_U3872, P2_U3873, P2_U3874, P2_U3875, P2_U3876, P2_U3877, P2_U3878, P2_U3879, P2_U3880, P2_U3881, P2_U3882, P2_U3883, P2_U3884, P2_U3885, P2_U3886, P2_U3887, P2_U3888, P2_U3889, P2_U3890, P2_U3891, P2_U3892, P2_U3893, P2_U3894, P2_U3895, P2_U3896, P2_U3897, P2_U3898, P2_U3899, P2_U3900, P2_U3901, P2_U3902, P2_U3903, P2_U3904, P2_U3905, P2_U3906, P2_U3907, P2_U3908, P2_U3909, P2_U3910, P2_U3911, P2_U3912, P2_U3913, P2_U3914, P2_U3915, P2_U3916, P2_U3917, P2_U3918, P2_U3919, P2_U3920, P2_U3921, P2_U3922, P2_U3923, P2_U3924, P2_U3925, P2_U3926, P2_U3927, P2_U3928, P2_U3929, P2_U3930, P2_U3931, P2_U3932, P2_U3933, P2_U3934, P2_U3935, P2_U3936, P2_U3937, P2_U3938, P2_U3939, P2_U3940, P2_U3941, P2_U3942, P2_U3943, P2_U3944, P2_U3945, P2_U3946, P2_U3947, P2_U3948, P2_U3949, P2_U3950, P2_U3951, P2_U3952, P2_U3953, P2_U3954, P2_U3955, P2_U3956, P2_U3957, P2_U3958, P2_U3959, P2_U3960, P2_U3961, P2_U3962, P2_U3963, P2_U3964, P2_U3965, P2_U3966, P2_U3967, P2_U3968, P2_U3969, P2_U3970, P2_U3971, P2_U3972, P2_U3973, P2_U3974, P2_U3975, P2_U3976, P2_U3977, P2_U3978, P2_U3979, P2_U3980, P2_U3981, P2_U3982, P2_U3983, P2_U3984, P2_U3985, P2_U3986, P2_U3987, P2_U3988, P2_U3989, P2_U3990, P2_U3991, P2_U3992, P2_U3993, P2_U3994, P2_U3995, P2_U3996, P2_U3997, P2_U3998, P2_U3999, P2_U4000, P2_U4001, P2_U4002, P2_U4003, P2_U4004, P2_U4005, P2_U4006, P2_U4007, P2_U4008, P2_U4009, P2_U4010, P2_U4011, P2_U4012, P2_U4013, P2_U4014, P2_U4015, P2_U4016, P2_U4017, P2_U4018, P2_U4019, P2_U4020, P2_U4021, P2_U4022, P2_U4023, P2_U4024, P2_U4025, P2_U4026, P2_U4027, P2_U4028, P2_U4029, P2_U4030, P2_U4031, P2_U4032, P2_U4033, P2_U4034, P2_U4035, P2_U4036, P2_U4037, P2_U4038, P2_U4039, P2_U4040, P2_U4041, P2_U4042, P2_U4043, P2_U4044, P2_U4045, P2_U4046, P2_U4047, P2_U4048, P2_U4049, P2_U4050, P2_U4051, P2_U4052, P2_U4053, P2_U4054, P2_U4055, P2_U4056, P2_U4057, P2_U4058, P2_U4059, P2_U4060, P2_U4061, P2_U4062, P2_U4063, P2_U4064, P2_U4065, P2_U4066, P2_U4067, P2_U4068, P2_U4069, P2_U4070, P2_U4071, P2_U4072, P2_U4073, P2_U4074, P2_U4075, P2_U4076, P2_U4077, P2_U4078, P2_U4079, P2_U4080, P2_U4081, P2_U4082, P2_U4083, P2_U4084, P2_U4085, P2_U4086, P2_U4087, P2_U4088, P2_U4089, P2_U4090, P2_U4091, P2_U4092, P2_U4093, P2_U4094, P2_U4095, P2_U4096, P2_U4097, P2_U4098, P2_U4099, P2_U4100, P2_U4101, P2_U4102, P2_U4103, P2_U4104, P2_U4105, P2_U4106, P2_U4107, P2_U4108, P2_U4109, P2_U4110, P2_U4111, P2_U4112, P2_U4113, P2_U4114, P2_U4115, P2_U4116, P2_U4117, P2_U4118, P2_U4119, P2_U4120, P2_U4121, P2_U4122, P2_U4123, P2_U4124, P2_U4125, P2_U4126, P2_U4127, P2_U4128, P2_U4129, P2_U4130, P2_U4131, P2_U4132, P2_U4133, P2_U4134, P2_U4135, P2_U4136, P2_U4137, P2_U4138, P2_U4139, P2_U4140, P2_U4141, P2_U4142, P2_U4143, P2_U4144, P2_U4145, P2_U4146, P2_U4147, P2_U4148, P2_U4149, P2_U4150, P2_U4151, P2_U4152, P2_U4153, P2_U4154, P2_U4155, P2_U4156, P2_U4157, P2_U4158, P2_U4159, P2_U4160, P2_U4161, P2_U4162, P2_U4163, P2_U4164, P2_U4165, P2_U4166, P2_U4167, P2_U4168, P2_U4169, P2_U4170, P2_U4171, P2_U4172, P2_U4173, P2_U4174, P2_U4175, P2_U4176, P2_U4177, P2_U4178, P2_U4179, P2_U4180, P2_U4181, P2_U4182, P2_U4183, P2_U4184, P2_U4185, P2_U4186, P2_U4187, P2_U4188, P2_U4189, P2_U4190, P2_U4191, P2_U4192, P2_U4193, P2_U4194, P2_U4195, P2_U4196, P2_U4197, P2_U4198, P2_U4199, P2_U4200, P2_U4201, P2_U4202, P2_U4203, P2_U4204, P2_U4205, P2_U4206, P2_U4207, P2_U4208, P2_U4209, P2_U4210, P2_U4211, P2_U4212, P2_U4213, P2_U4214, P2_U4215, P2_U4216, P2_U4217, P2_U4218, P2_U4219, P2_U4220, P2_U4221, P2_U4222, P2_U4223, P2_U4224, P2_U4225, P2_U4226, P2_U4227, P2_U4228, P2_U4229, P2_U4230, P2_U4231, P2_U4232, P2_U4233, P2_U4234, P2_U4235, P2_U4236, P2_U4237, P2_U4238, P2_U4239, P2_U4240, P2_U4241, P2_U4242, P2_U4243, P2_U4244, P2_U4245, P2_U4246, P2_U4247, P2_U4248, P2_U4249, P2_U4250, P2_U4251, P2_U4252, P2_U4253, P2_U4254, P2_U4255, P2_U4256, P2_U4257, P2_U4258, P2_U4259, P2_U4260, P2_U4261, P2_U4262, P2_U4263, P2_U4264, P2_U4265, P2_U4266, P2_U4267, P2_U4268, P2_U4269, P2_U4270, P2_U4271, P2_U4272, P2_U4273, P2_U4274, P2_U4275, P2_U4276, P2_U4277, P2_U4278, P2_U4279, P2_U4280, P2_U4281, P2_U4282, P2_U4283, P2_U4284, P2_U4285, P2_U4286, P2_U4287, P2_U4288, P2_U4289, P2_U4290, P2_U4291, P2_U4292, P2_U4293, P2_U4294, P2_U4295, P2_U4296, P2_U4297, P2_U4298, P2_U4299, P2_U4300, P2_U4301, P2_U4302, P2_U4303, P2_U4304, P2_U4305, P2_U4306, P2_U4307, P2_U4308, P2_U4309, P2_U4310, P2_U4311, P2_U4312, P2_U4313, P2_U4314, P2_U4315, P2_U4316, P2_U4317, P2_U4318, P2_U4319, P2_U4320, P2_U4321, P2_U4322, P2_U4323, P2_U4324, P2_U4325, P2_U4326, P2_U4327, P2_U4328, P2_U4329, P2_U4330, P2_U4331, P2_U4332, P2_U4333, P2_U4334, P2_U4335, P2_U4336, P2_U4337, P2_U4338, P2_U4339, P2_U4340, P2_U4341, P2_U4342, P2_U4343, P2_U4344, P2_U4345, P2_U4346, P2_U4347, P2_U4348, P2_U4349, P2_U4350, P2_U4351, P2_U4352, P2_U4353, P2_U4354, P2_U4355, P2_U4356, P2_U4357, P2_U4358, P2_U4359, P2_U4360, P2_U4361, P2_U4362, P2_U4363, P2_U4364, P2_U4365, P2_U4366, P2_U4367, P2_U4368, P2_U4369, P2_U4370, P2_U4371, P2_U4372, P2_U4373, P2_U4374, P2_U4375, P2_U4376, P2_U4377, P2_U4378, P2_U4379, P2_U4380, P2_U4381, P2_U4382, P2_U4383, P2_U4384, P2_U4385, P2_U4386, P2_U4387, P2_U4388, P2_U4389, P2_U4390, P2_U4391, P2_U4392, P2_U4393, P2_U4394, P2_U4395, P2_U4396, P2_U4397, P2_U4398, P2_U4399, P2_U4400, P2_U4401, P2_U4402, P2_U4403, P2_U4404, P2_U4405, P2_U4406, P2_U4407, P2_U4408, P2_U4409, P2_U4410, P2_U4411, P2_U4412, P2_U4413, P2_U4414, P2_U4415, P2_U4416, P2_U4417, P2_U4418, P2_U4419, P2_U4420, P2_U4421, P2_U4422, P2_U4423, P2_U4424, P2_U4425, P2_U4426, P2_U4427, P2_U4428, P2_U4429, P2_U4430, P2_U4431, P2_U4432, P2_U4433, P2_U4434, P2_U4435, P2_U4436, P2_U4437, P2_U4438, P2_U4439, P2_U4440, P2_U4441, P2_U4442, P2_U4443, P2_U4444, P2_U4445, P2_U4446, P2_U4447, P2_U4448, P2_U4449, P2_U4450, P2_U4451, P2_U4452, P2_U4453, P2_U4454, P2_U4455, P2_U4456, P2_U4457, P2_U4458, P2_U4459, P2_U4460, P2_U4461, P2_U4462, P2_U4463, P2_U4464, P2_U4465, P2_U4466, P2_U4467, P2_U4468, P2_U4469, P2_U4470, P2_U4471, P2_U4472, P2_U4473, P2_U4474, P2_U4475, P2_U4476, P2_U4477, P2_U4478, P2_U4479, P2_U4480, P2_U4481, P2_U4482, P2_U4483, P2_U4484, P2_U4485, P2_U4486, P2_U4487, P2_U4488, P2_U4489, P2_U4490, P2_U4491, P2_U4492, P2_U4493, P2_U4494, P2_U4495, P2_U4496, P2_U4497, P2_U4498, P2_U4499, P2_U4500, P2_U4501, P2_U4502, P2_U4503, P2_U4504, P2_U4505, P2_U4506, P2_U4507, P2_U4508, P2_U4509, P2_U4510, P2_U4511, P2_U4512, P2_U4513, P2_U4514, P2_U4515, P2_U4516, P2_U4517, P2_U4518, P2_U4519, P2_U4520, P2_U4521, P2_U4522, P2_U4523, P2_U4524, P2_U4525, P2_U4526, P2_U4527, P2_U4528, P2_U4529, P2_U4530, P2_U4531, P2_U4532, P2_U4533, P2_U4534, P2_U4535, P2_U4536, P2_U4537, P2_U4538, P2_U4539, P2_U4540, P2_U4541, P2_U4542, P2_U4543, P2_U4544, P2_U4545, P2_U4546, P2_U4547, P2_U4548, P2_U4549, P2_U4550, P2_U4551, P2_U4552, P2_U4553, P2_U4554, P2_U4555, P2_U4556, P2_U4557, P2_U4558, P2_U4559, P2_U4560, P2_U4561, P2_U4562, P2_U4563, P2_U4564, P2_U4565, P2_U4566, P2_U4567, P2_U4568, P2_U4569, P2_U4570, P2_U4571, P2_U4572, P2_U4573, P2_U4574, P2_U4575, P2_U4576, P2_U4577, P2_U4578, P2_U4579, P2_U4580, P2_U4581, P2_U4582, P2_U4583, P2_U4584, P2_U4585, P2_U4586, P2_U4587, P2_U4588, P2_U4589, P2_U4590, P2_U4591, P2_U4592, P2_U4593, P2_U4594, P2_U4595, P2_U4596, P2_U4597, P2_U4598, P2_U4599, P2_U4600, P2_U4601, P2_U4602, P2_U4603, P2_U4604, P2_U4605, P2_U4606, P2_U4607, P2_U4608, P2_U4609, P2_U4610, P2_U4611, P2_U4612, P2_U4613, P2_U4614, P2_U4615, P2_U4616, P2_U4617, P2_U4618, P2_U4619, P2_U4620, P2_U4621, P2_U4622, P2_U4623, P2_U4624, P2_U4625, P2_U4626, P2_U4627, P2_U4628, P2_U4629, P2_U4630, P2_U4631, P2_U4632, P2_U4633, P2_U4634, P2_U4635, P2_U4636, P2_U4637, P2_U4638, P2_U4639, P2_U4640, P2_U4641, P2_U4642, P2_U4643, P2_U4644, P2_U4645, P2_U4646, P2_U4647, P2_U4648, P2_U4649, P2_U4650, P2_U4651, P2_U4652, P2_U4653, P2_U4654, P2_U4655, P2_U4656, P2_U4657, P2_U4658, P2_U4659, P2_U4660, P2_U4661, P2_U4662, P2_U4663, P2_U4664, P2_U4665, P2_U4666, P2_U4667, P2_U4668, P2_U4669, P2_U4670, P2_U4671, P2_U4672, P2_U4673, P2_U4674, P2_U4675, P2_U4676, P2_U4677, P2_U4678, P2_U4679, P2_U4680, P2_U4681, P2_U4682, P2_U4683, P2_U4684, P2_U4685, P2_U4686, P2_U4687, P2_U4688, P2_U4689, P2_U4690, P2_U4691, P2_U4692, P2_U4693, P2_U4694, P2_U4695, P2_U4696, P2_U4697, P2_U4698, P2_U4699, P2_U4700, P2_U4701, P2_U4702, P2_U4703, P2_U4704, P2_U4705, P2_U4706, P2_U4707, P2_U4708, P2_U4709, P2_U4710, P2_U4711, P2_U4712, P2_U4713, P2_U4714, P2_U4715, P2_U4716, P2_U4717, P2_U4718, P2_U4719, P2_U4720, P2_U4721, P2_U4722, P2_U4723, P2_U4724, P2_U4725, P2_U4726, P2_U4727, P2_U4728, P2_U4729, P2_U4730, P2_U4731, P2_U4732, P2_U4733, P2_U4734, P2_U4735, P2_U4736, P2_U4737, P2_U4738, P2_U4739, P2_U4740, P2_U4741, P2_U4742, P2_U4743, P2_U4744, P2_U4745, P2_U4746, P2_U4747, P2_U4748, P2_U4749, P2_U4750, P2_U4751, P2_U4752, P2_U4753, P2_U4754, P2_U4755, P2_U4756, P2_U4757, P2_U4758, P2_U4759, P2_U4760, P2_U4761, P2_U4762, P2_U4763, P2_U4764, P2_U4765, P2_U4766, P2_U4767, P2_U4768, P2_U4769, P2_U4770, P2_U4771, P2_U4772, P2_U4773, P2_U4774, P2_U4775, P2_U4776, P2_U4777, P2_U4778, P2_U4779, P2_U4780, P2_U4781, P2_U4782, P2_U4783, P2_U4784, P2_U4785, P2_U4786, P2_U4787, P2_U4788, P2_U4789, P2_U4790, P2_U4791, P2_U4792, P2_U4793, P2_U4794, P2_U4795, P2_U4796, P2_U4797, P2_U4798, P2_U4799, P2_U4800, P2_U4801, P2_U4802, P2_U4803, P2_U4804, P2_U4805, P2_U4806, P2_U4807, P2_U4808, P2_U4809, P2_U4810, P2_U4811, P2_U4812, P2_U4813, P2_U4814, P2_U4815, P2_U4816, P2_U4817, P2_U4818, P2_U4819, P2_U4820, P2_U4821, P2_U4822, P2_U4823, P2_U4824, P2_U4825, P2_U4826, P2_U4827, P2_U4828, P2_U4829, P2_U4830, P2_U4831, P2_U4832, P2_U4833, P2_U4834, P2_U4835, P2_U4836, P2_U4837, P2_U4838, P2_U4839, P2_U4840, P2_U4841, P2_U4842, P2_U4843, P2_U4844, P2_U4845, P2_U4846, P2_U4847, P2_U4848, P2_U4849, P2_U4850, P2_U4851, P2_U4852, P2_U4853, P2_U4854, P2_U4855, P2_U4856, P2_U4857, P2_U4858, P2_U4859, P2_U4860, P2_U4861, P2_U4862, P2_U4863, P2_U4864, P2_U4865, P2_U4866, P2_U4867, P2_U4868, P2_U4869, P2_U4870, P2_U4871, P2_U4872, P2_U4873, P2_U4874, P2_U4875, P2_U4876, P2_U4877, P2_U4878, P2_U4879, P2_U4880, P2_U4881, P2_U4882, P2_U4883, P2_U4884, P2_U4885, P2_U4886, P2_U4887, P2_U4888, P2_U4889, P2_U4890, P2_U4891, P2_U4892, P2_U4893, P2_U4894, P2_U4895, P2_U4896, P2_U4897, P2_U4898, P2_U4899, P2_U4900, P2_U4901, P2_U4902, P2_U4903, P2_U4904, P2_U4905, P2_U4906, P2_U4907, P2_U4908, P2_U4909, P2_U4910, P2_U4911, P2_U4912, P2_U4913, P2_U4914, P2_U4915, P2_U4916, P2_U4917, P2_U4918, P2_U4919, P2_U4920, P2_U4921, P2_U4922, P2_U4923, P2_U4924, P2_U4925, P2_U4926, P2_U4927, P2_U4928, P2_U4929, P2_U4930, P2_U4931, P2_U4932, P2_U4933, P2_U4934, P2_U4935, P2_U4936, P2_U4937, P2_U4938, P2_U4939, P2_U4940, P2_U4941, P2_U4942, P2_U4943, P2_U4944, P2_U4945, P2_U4946, P2_U4947, P2_U4948, P2_U4949, P2_U4950, P2_U4951, P2_U4952, P2_U4953, P2_U4954, P2_U4955, P2_U4956, P2_U4957, P2_U4958, P2_U4959, P2_U4960, P2_U4961, P2_U4962, P2_U4963, P2_U4964, P2_U4965, P2_U4966, P2_U4967, P2_U4968, P2_U4969, P2_U4970, P2_U4971, P2_U4972, P2_U4973, P2_U4974, P2_U4975, P2_U4976, P2_U4977, P2_U4978, P2_U4979, P2_U4980, P2_U4981, P2_U4982, P2_U4983, P2_U4984, P2_U4985, P2_U4986, P2_U4987, P2_U4988, P2_U4989, P2_U4990, P2_U4991, P2_U4992, P2_U4993, P2_U4994, P2_U4995, P2_U4996, P2_U4997, P2_U4998, P2_U4999, P2_U5000, P2_U5001, P2_U5002, P2_U5003, P2_U5004, P2_U5005, P2_U5006, P2_U5007, P2_U5008, P2_U5009, P2_U5010, P2_U5011, P2_U5012, P2_U5013, P2_U5014, P2_U5015, P2_U5016, P2_U5017, P2_U5018, P2_U5019, P2_U5020, P2_U5021, P2_U5022, P2_U5023, P2_U5024, P2_U5025, P2_U5026, P2_U5027, P2_U5028, P2_U5029, P2_U5030, P2_U5031, P2_U5032, P2_U5033, P2_U5034, P2_U5035, P2_U5036, P2_U5037, P2_U5038, P2_U5039, P2_U5040, P2_U5041, P2_U5042, P2_U5043, P2_U5044, P2_U5045, P2_U5046, P2_U5047, P2_U5048, P2_U5049, P2_U5050, P2_U5051, P2_U5052, P2_U5053, P2_U5054, P2_U5055, P2_U5056, P2_U5057, P2_U5058, P2_U5059, P2_U5060, P2_U5061, P2_U5062, P2_U5063, P2_U5064, P2_U5065, P2_U5066, P2_U5067, P2_U5068, P2_U5069, P2_U5070, P2_U5071, P2_U5072, P2_U5073, P2_U5074, P2_U5075, P2_U5076, P2_U5077, P2_U5078, P2_U5079, P2_U5080, P2_U5081, P2_U5082, P2_U5083, P2_U5084, P2_U5085, P2_U5086, P2_U5087, P2_U5088, P2_U5089, P2_U5090, P2_U5091, P2_U5092, P2_U5093, P2_U5094, P2_U5095, P2_U5096, P2_U5097, P2_U5098, P2_U5099, P2_U5100, P2_U5101, P2_U5102, P2_U5103, P2_U5104, P2_U5105, P2_U5106, P2_U5107, P2_U5108, P2_U5109, P2_U5110, P2_U5111, P2_U5112, P2_U5113, P2_U5114, P2_U5115, P2_U5116, P2_U5117, P2_U5118, P2_U5119, P2_U5120, P2_U5121, P2_U5122, P2_U5123, P2_U5124, P2_U5125, P2_U5126, P2_U5127, P2_U5128, P2_U5129, P2_U5130, P2_U5131, P2_U5132, P2_U5133, P2_U5134, P2_U5135, P2_U5136, P2_U5137, P2_U5138, P2_U5139, P2_U5140, P2_U5141, P2_U5142, P2_U5143, P2_U5144, P2_U5145, P2_U5146, P2_U5147, P2_U5148, P2_U5149, P2_U5150, P2_U5151, P2_U5152, P2_U5153, P2_U5154, P2_U5155, P2_U5156, P2_U5157, P2_U5158, P2_U5159, P2_U5160, P2_U5161, P2_U5162, P2_U5163, P2_U5164, P2_U5165, P2_U5166, P2_U5167, P2_U5168, P2_U5169, P2_U5170, P2_U5171, P2_U5172, P2_U5173, P2_U5174, P2_U5175, P2_U5176, P2_U5177, P2_U5178, P2_U5179, P2_U5180, P2_U5181, P2_U5182, P2_U5183, P2_U5184, P2_U5185, P2_U5186, P2_U5187, P2_U5188, P2_U5189, P2_U5190, P2_U5191, P2_U5192, P2_U5193, P2_U5194, P2_U5195, P2_U5196, P2_U5197, P2_U5198, P2_U5199, P2_U5200, P2_U5201, P2_U5202, P2_U5203, P2_U5204, P2_U5205, P2_U5206, P2_U5207, P2_U5208, P2_U5209, P2_U5210, P2_U5211, P2_U5212, P2_U5213, P2_U5214, P2_U5215, P2_U5216, P2_U5217, P2_U5218, P2_U5219, P2_U5220, P2_U5221, P2_U5222, P2_U5223, P2_U5224, P2_U5225, P2_U5226, P2_U5227, P2_U5228, P2_U5229, P2_U5230, P2_U5231, P2_U5232, P2_U5233, P2_U5234, P2_U5235, P2_U5236, P2_U5237, P2_U5238, P2_U5239, P2_U5240, P2_U5241, P2_U5242, P2_U5243, P2_U5244, P2_U5245, P2_U5246, P2_U5247, P2_U5248, P2_U5249, P2_U5250, P2_U5251, P2_U5252, P2_U5253, P2_U5254, P2_U5255, P2_U5256, P2_U5257, P2_U5258, P2_U5259, P2_U5260, P2_U5261, P2_U5262, P2_U5263, P2_U5264, P2_U5265, P2_U5266, P2_U5267, P2_U5268, P2_U5269, P2_U5270, P2_U5271, P2_U5272, P2_U5273, P2_U5274, P2_U5275, P2_U5276, P2_U5277, P2_U5278, P2_U5279, P2_U5280, P2_U5281, P2_U5282, P2_U5283, P2_U5284, P2_U5285, P2_U5286, P2_U5287, P2_U5288, P2_U5289, P2_U5290, P2_U5291, P2_U5292, P2_U5293, P2_U5294, P2_U5295, P2_U5296, P2_U5297, P2_U5298, P2_U5299, P2_U5300, P2_U5301, P2_U5302, P2_U5303, P2_U5304, P2_U5305, P2_U5306, P2_U5307, P2_U5308, P2_U5309, P2_U5310, P2_U5311, P2_U5312, P2_U5313, P2_U5314, P2_U5315, P2_U5316, P2_U5317, P2_U5318, P2_U5319, P2_U5320, P2_U5321, P2_U5322, P2_U5323, P2_U5324, P2_U5325, P2_U5326, P2_U5327, P2_U5328, P2_U5329, P2_U5330, P2_U5331, P2_U5332, P2_U5333, P2_U5334, P2_U5335, P2_U5336, P2_U5337, P2_U5338, P2_U5339, P2_U5340, P2_U5341, P2_U5342, P2_U5343, P2_U5344, P2_U5345, P2_U5346, P2_U5347, P2_U5348, P2_U5349, P2_U5350, P2_U5351, P2_U5352, P2_U5353, P2_U5354, P2_U5355, P2_U5356, P2_U5357, P2_U5358, P2_U5359, P2_U5360, P2_U5361, P2_U5362, P2_U5363, P2_U5364, P2_U5365, P2_U5366, P2_U5367, P2_U5368, P2_U5369, P2_U5370, P2_U5371, P2_U5372, P2_U5373, P2_U5374, P2_U5375, P2_U5376, P2_U5377, P2_U5378, P2_U5379, P2_U5380, P2_U5381, P2_U5382, P2_U5383, P2_U5384, P2_U5385, P2_U5386, P2_U5387, P2_U5388, P2_U5389, P2_U5390, P2_U5391, P2_U5392, P2_U5393, P2_U5394, P2_U5395, P2_U5396, P2_U5397, P2_U5398, P2_U5399, P2_U5400, P2_U5401, P2_U5402, P2_U5403, P2_U5404, P2_U5405, P2_U5406, P2_U5407, P2_U5408, P2_U5409, P2_U5410, P2_U5411, P2_U5412, P2_U5413, P2_U5414, P2_U5415, P2_U5416, P2_U5417, P2_U5418, P2_U5419, P2_U5420, P2_U5421, P2_U5422, P2_U5423, P2_U5424, P2_U5425, P2_U5426, P2_U5427, P2_U5428, P2_U5429, P2_U5430, P2_U5431, P2_U5432, P2_U5433, P2_U5434, P2_U5435, P2_U5436, P2_U5437, P2_U5438, P2_U5439, P2_U5440, P2_U5441, P2_U5442, P2_U5443, P2_U5444, P2_U5445, P2_U5446, P2_U5447, P2_U5448, P2_U5449, P2_U5450, P2_U5451, P2_U5452, P2_U5453, P2_U5454, P2_U5455, P2_U5456, P2_U5457, P2_U5458, P2_U5459, P2_U5460, P2_U5461, P2_U5462, P2_U5463, P2_U5464, P2_U5465, P2_U5466, P2_U5467, P2_U5468, P2_U5469, P2_U5470, P2_U5471, P2_U5472, P2_U5473, P2_U5474, P2_U5475, P2_U5476, P2_U5477, P2_U5478, P2_U5479, P2_U5480, P2_U5481, P2_U5482, P2_U5483, P2_U5484, P2_U5485, P2_U5486, P2_U5487, P2_U5488, P2_U5489, P2_U5490, P2_U5491, P2_U5492, P2_U5493, P2_U5494, P2_U5495, P2_U5496, P2_U5497, P2_U5498, P2_U5499, P2_U5500, P2_U5501, P2_U5502, P2_U5503, P2_U5504, P2_U5505, P2_U5506, P2_U5507, P2_U5508, P2_U5509, P2_U5510, P2_U5511, P2_U5512, P2_U5513, P2_U5514, P2_U5515, P2_U5516, P2_U5517, P2_U5518, P2_U5519, P2_U5520, P2_U5521, P2_U5522, P2_U5523, P2_U5524, P2_U5525, P2_U5526, P2_U5527, P2_U5528, P2_U5529, P2_U5530, P2_U5531, P2_U5532, P2_U5533, P2_U5534, P2_U5535, P2_U5536, P2_U5537, P2_U5538, P2_U5539, P2_U5540, P2_U5541, P2_U5542, P2_U5543, P2_U5544, P2_U5545, P2_U5546, P2_U5547, P2_U5548, P2_U5549, P2_U5550, P2_U5551, P2_U5552, P2_U5553, P2_U5554, P2_U5555, P2_U5556, P2_U5557, P2_U5558, P2_U5559, P2_U5560, P2_U5561, P2_U5562, P2_U5563, P2_U5564, P2_U5565, P2_U5566, P2_U5567, P2_U5568, P2_U5569, P2_U5570, P2_U5571, P2_U5572, P2_U5573, P2_U5574, P2_U5575, P2_U5576, P2_U5577, P2_U5578, P2_U5579, P2_U5580, P2_U5581, P2_U5582, P2_U5583, P2_U5584, P2_U5585, P2_U5586, P2_U5587, P2_U5588, P2_U5589, P2_U5590, P2_U5591, P2_U5592, P2_U5593, P2_U5594, P2_U5595, P2_U5596, P2_U5597, P2_U5598, P2_U5599, P2_U5600, P2_U5601, P2_U5602, P2_U5603, P2_U5604, P2_U5605, P2_U5606, P2_U5607, P2_U5608, P2_U5609, P2_U5610, P2_U5611, P2_U5612, P2_U5613, P2_U5614, P2_U5615, P2_U5616, P2_U5617, P2_U5618, P2_U5619, P2_U5620, P2_U5621, P2_U5622, P2_U5623, P2_U5624, P2_U5625, P2_U5626, P2_U5627, P2_U5628, P2_U5629, P2_U5630, P2_U5631, P2_U5632, P2_U5633, P2_U5634, P2_U5635, P2_U5636, P2_U5637, P2_U5638, P2_U5639, P2_U5640, P2_U5641, P2_U5642, P2_U5643, P2_U5644, P2_U5645, P2_U5646, P2_U5647, P2_U5648, P2_U5649, P2_U5650, P2_U5651, P2_U5652, P2_U5653, P2_U5654, P2_U5655, P2_U5656, P2_U5657, P2_U5658, P2_U5659, P2_U5660, P2_U5661, P2_U5662, P2_U5663, P2_U5664, P2_U5665, P2_U5666, P2_U5667, P2_U5668, P2_U5669, P2_U5670, P2_U5671, P2_U5672, P2_U5673, P2_U5674, P2_U5675, P2_U5676, P2_U5677, P2_U5678, P2_U5679, P2_U5680, P2_U5681, P2_U5682, P2_U5683, P2_U5684, P2_U5685, P2_U5686, P2_U5687, P2_U5688, P2_U5689, P2_U5690, P2_U5691, P2_U5692, P2_U5693, P2_U5694, P2_U5695, P2_U5696, P2_U5697, P2_U5698, P2_U5699, P2_U5700, P2_U5701, P2_U5702, P2_U5703, P2_U5704, P2_U5705, P2_U5706, P2_U5707, P2_U5708, P2_U5709, P2_U5710, P2_U5711, P2_U5712, P2_U5713, P2_U5714, P2_U5715, P2_U5716, P2_U5717, P2_U5718, P2_U5719, P2_U5720, P2_U5721, P2_U5722, P2_U5723, P2_U5724, P2_U5725, P2_U5726, P2_U5727, P2_U5728, P2_U5729, P2_U5730, P2_U5731, P2_U5732, P2_U5733, P2_U5734, P2_U5735, P2_U5736, P2_U5737, P2_U5738, P2_U5739, P2_U5740, P2_U5741, P2_U5742, P2_U5743, P2_U5744, P2_U5745, P2_U5746, P2_U5747, P2_U5748, P2_U5749, P2_U5750, P2_U5751, P2_U5752, P2_U5753, P2_U5754, P2_U5755, P2_U5756, P2_U5757, P2_U5758, P2_U5759, P2_U5760, P2_U5761, P2_U5762, P2_U5763, P2_U5764, P2_U5765, P2_U5766, P2_U5767, P2_U5768, P2_U5769, P2_U5770, P2_U5771, P2_U5772, P2_U5773, P2_U5774, P2_U5775, P2_U5776, P2_U5777, P2_U5778, P2_U5779, P2_U5780, P2_U5781, P2_U5782, P2_U5783, P2_U5784, P2_U5785, P2_U5786, P2_U5787, P2_U5788, P2_U5789, P2_U5790, P2_U5791, P2_U5792, P2_U5793, P2_U5794, P2_U5795, P2_U5796, P2_U5797, P2_U5798, P2_U5799, P2_U5800, P2_U5801, P2_U5802, P2_U5803, P2_U5804, P2_U5805, P2_U5806, P2_U5807, P2_U5808, P2_U5809, P2_U5810, P2_U5811, P2_U5812, P2_U5813, P2_U5814, P2_U5815, P2_U5816, P2_U5817, P2_U5818, P2_U5819, P2_U5820, P2_U5821, P2_U5822, P2_U5823, P2_U5824, P2_U5825, P2_U5826, P2_U5827, P2_U5828, P2_U5829, P2_U5830, P2_U5831, P2_U5832, P2_U5833, P2_U5834, P2_U5835, P2_U5836, P2_U5837, P2_U5838, P2_U5839, P2_U5840, P2_U5841, P2_U5842, P2_U5843, P2_U5844, P2_U5845, P2_U5846, P2_U5847, P2_U5848, P2_U5849, P2_U5850, P2_U5851, P2_U5852, P2_U5853, P2_U5854, P2_U5855, P2_U5856, P2_U5857, P2_U5858, P2_U5859, P2_U5860, P2_U5861, P2_U5862, P2_U5863, P2_U5864, P2_U5865, P2_U5866, P2_U5867, P2_U5868, P2_U5869, P2_U5870, P2_U5871, P2_U5872, P2_U5873, P2_U5874, P2_U5875, P2_U5876, P2_U5877, P2_U5878, P2_U5879, P2_U5880, P2_U5881, P2_U5882, P2_U5883, P2_U5884, P2_U5885, P2_U5886, P2_U5887, P2_U5888, P2_U5889, P2_U5890, P2_U5891, P2_U5892, P2_U5893, P2_U5894, P2_U5895, P2_U5896, P2_U5897, P2_U5898, P2_U5899, P2_U5900, P2_U5901, P2_U5902, P2_U5903, P2_U5904, P2_U5905, P2_U5906, P2_U5907, P2_U5908, P2_U5909, P2_U5910, P2_U5911, P2_U5912, P2_U5913, P2_U5914, P2_U5915, P2_U5916, P2_U5917, P2_U5918, P2_U5919, P2_U5920, P2_U5921, P2_U5922, P2_U5923, P2_U5924, P2_U5925, P2_U5926, P2_U5927, P2_U5928, P2_U5929, P2_U5930, P2_U5931, P2_U5932, P2_U5933, P2_U5934, P2_U5935, P2_U5936, P2_U5937, P2_U5938, P2_U5939, P2_U5940, P2_U5941, P2_U5942, P2_U5943, P2_U5944, P2_U5945, P2_U5946, P2_U5947, P2_U5948, P2_U5949, P2_U5950, P2_U5951, P2_U5952, P2_U5953, P2_U5954, P2_U5955, P2_U5956, P2_U5957, P2_U5958, P2_U5959, P2_U5960, P2_U5961, P2_U5962, P2_U5963, P2_U5964, P2_U5965, P2_U5966, P2_U5967, P2_U5968, P2_U5969, P2_U5970, P2_U5971, P2_U5972, P2_U5973, P2_U5974, P2_U5975, P2_U5976, P2_U5977, P2_U5978, P2_U5979, P2_U5980, P2_U5981, P2_U5982, P2_U5983, P2_U5984, P2_U5985, P2_U5986, P2_U5987, P2_U5988, P2_U5989, P2_U5990, P2_U5991, P2_U5992, P2_U5993, P2_U5994, P2_U5995, P2_U5996, P2_U5997, P2_U5998, P2_U5999, P2_U6000, P2_U6001, P2_U6002, P2_U6003, P2_U6004, P2_U6005, P2_U6006, P2_U6007, P2_U6008, P2_U6009, P2_U6010, P2_U6011, P2_U6012, P2_U6013, P2_U6014, P2_U6015, P2_U6016, P2_U6017, P2_U6018, P2_U6019, P2_U6020, P2_U6021, P2_U6022, P2_U6023, P2_U6024, P2_U6025, P2_U6026, P2_U6027, P2_U6028, P2_U6029, P2_U6030, P2_U6031, P2_U6032, P2_U6033, P2_U6034, P2_U6035, P2_U6036, P2_U6037, P2_U6038, P2_U6039, P2_U6040, P2_U6041, P2_U6042, P2_U6043, P2_U6044, P2_U6045, P2_U6046, P2_U6047, P2_U6048, P2_U6049, P2_U6050, P2_U6051, P2_U6052, P2_U6053, P2_U6054, P2_U6055, P2_U6056, P2_U6057, P2_U6058, P2_U6059, P2_U6060, P2_U6061, P2_U6062, P2_U6063, P2_U6064, P2_U6065, P2_U6066, P2_U6067, P2_U6068, P2_U6069, P2_U6070, P2_U6071, P2_U6072, P2_U6073, P2_U6074, P2_U6075, P2_U6076, P2_U6077, P2_U6078, P2_U6079, P2_U6080, P2_U6081, P2_U6082, P2_U6083, P2_U6084, P2_U6085, P2_U6086, P2_U6087, P2_U6088, P2_U6089, P2_U6090, P2_U6091, P2_U6092, P2_U6093, P2_U6094, P2_U6095, P2_U6096, P2_U6097, P2_U6098, P2_U6099, P2_U6100, P2_U6101, P2_U6102, P2_U6103, P2_U6104, P2_U6105, P2_U6106, P2_U6107, P2_U6108, P2_U6109, P2_U6110, P2_U6111, P2_U6112, P2_U6113, P2_U6114, P2_U6115, P2_U6116, P2_U6117, P2_U6118, P2_U6119, P2_U6120, P2_U6121, P2_U6122, P2_U6123, P2_U6124, P2_U6125, P2_U6126, P2_U6127, P2_U6128, P2_U6129, P2_U6130, P2_U6131, P2_U6132, P2_U6133, P2_U6134, P2_U6135, P2_U6136, P2_U6137, P2_U6138, P2_U6139, P2_U6140, P2_U6141, P2_U6142, P2_U6143, P2_U6144, P2_U6145, P2_U6146, P2_U6147, P2_U6148, P2_U6149, P2_U6150, P2_U6151, P2_U6152, P2_U6153, P2_U6154, P2_U6155, P2_U6156, P2_U6157, P2_U6158, P2_U6159, P2_U6160, P2_U6161, P2_U6162, P2_U6163, P2_U6164, P2_U6165, P2_U6166, P2_U6167, P2_U6168, P2_U6169, P2_U6170, P2_U6171, P2_U6172, P2_U6173, P2_U6174, P2_U6175, P2_U6176, P2_U6177, P2_U6178, P2_U6179, P2_U6180, P2_U6181, P2_U6182, P2_U6183, P2_U6184, P2_U6185, P2_U6186, P2_U6187, P2_U6188, P2_U6189, P2_U6190, P2_U6191, P2_U6192, P2_U6193, P2_U6194, P2_U6195, P2_U6196, P2_U6197, P2_U6198, P2_U6199, P2_U6200, P2_U6201, P2_U6202, P2_U6203, P2_U6204, P2_U6205, P2_U6206, P2_U6207, P2_U6208, P2_U6209, P2_U6210, P2_U6211, P2_U6212, P2_U6213, P2_U6214, P2_U6215, P2_U6216, P2_U6217, P2_U6218, P2_U6219, P2_U6220, P2_U6221, P2_U6222, P2_U6223, P2_U6224, P2_U6225, P2_U6226, P2_U6227, P2_U6228, P2_U6229, P2_U6230, P2_U6231, P2_U6232, P2_U6233, P2_U6234, P2_U6235, P2_U6236, P2_U6237, P2_U6238, P2_U6239, P2_U6240, P2_U6241, P2_U6242, P2_U6243, P2_U6244, P2_U6245, P2_U6246, P2_U6247, P2_U6248, P2_U6249, P2_U6250, P2_U6251, P2_U6252, P2_U6253, P2_U6254, P2_U6255, P2_U6256, P2_U6257, P2_U6258, P2_U6259, P2_U6260, P2_U6261, P2_U6262, P2_U6263, P2_U6264, P2_U6265, P2_U6266, P2_U6267, P2_U6268, P2_U6269, P2_U6270, P2_U6271, P2_U6272, P2_U6273, P2_U6274, P2_U6275, P2_U6276, P2_U6277, P2_U6278, P2_U6279, P2_U6280, P2_U6281, P2_U6282, P2_U6283, P2_U6284, P2_U6285, P2_U6286, P2_U6287, P2_U6288, P2_U6289, P2_U6290, P2_U6291, P2_U6292, P2_U6293, P2_U6294, P2_U6295, P2_U6296, P2_U6297, P2_U6298, P2_U6299, P2_U6300, P2_U6301, P2_U6302, P2_U6303, P2_U6304, P2_U6305, P2_U6306, P2_U6307, P2_U6308, P2_U6309, P2_U6310, P2_U6311, P2_U6312, P2_U6313, P2_U6314, P2_U6315, P2_U6316, P2_U6317, P2_U6318, P2_U6319, P2_U6320, P2_U6321, P2_U6322, P2_U6323, P2_U6324, P2_U6325, P2_U6326, P2_U6327, P2_U6328, P2_U6329, P2_U6330, P2_U6331, P2_U6332, P2_U6333, P2_U6334, P2_U6335, P2_U6336, P2_U6337, P2_U6338, P2_U6339, P2_U6340, P2_U6341, P2_U6342, P2_U6343, P2_U6344, P2_U6345, P2_U6346, P2_U6347, P2_U6348, P2_U6349, P2_U6350, P2_U6351, P2_U6352, P2_U6353, P2_U6354, P2_U6355, P2_U6356, P2_U6357, P2_U6358, P2_U6359, P2_U6360, P2_U6361, P2_U6362, P2_U6363, P2_U6364, P2_U6365, P2_U6366, P2_U6367, P2_U6368, P2_U6369, P2_U6370, P2_U6371, P2_U6372, P2_U6373, P2_U6374, P2_U6375, P2_U6376, P2_U6377, P2_U6378, P2_U6379, P2_U6380, P2_U6381, P2_U6382, P2_U6383, P2_U6384, P2_U6385, P2_U6386, P2_U6387, P2_U6388, P2_U6389, P2_U6390, P2_U6391, P2_U6392, P2_U6393, P2_U6394, P2_U6395, P2_U6396, P2_U6397, P2_U6398, P2_U6399, P2_U6400, P2_U6401, P2_U6402, P2_U6403, P2_U6404, P2_U6405, P2_U6406, P2_U6407, P2_U6408, P2_U6409, P2_U6410, P2_U6411, P2_U6412, P2_U6413, P2_U6414, P2_U6415, P2_U6416, P2_U6417, P2_U6418, P2_U6419, P2_U6420, P2_U6421, P2_U6422, P2_U6423, P2_U6424, P2_U6425, P2_U6426, P2_U6427, P2_U6428, P2_U6429, P2_U6430, P2_U6431, P2_U6432, P2_U6433, P2_U6434, P2_U6435, P2_U6436, P2_U6437, P2_U6438, P2_U6439, P2_U6440, P2_U6441, P2_U6442, P2_U6443, P2_U6444, P2_U6445, P2_U6446, P2_U6447, P2_U6448, P2_U6449, P2_U6450, P2_U6451, P2_U6452, P2_U6453, P2_U6454, P2_U6455, P2_U6456, P2_U6457, P2_U6458, P2_U6459, P2_U6460, P2_U6461, P2_U6462, P2_U6463, P2_U6464, P2_U6465, P2_U6466, P2_U6467, P2_U6468, P2_U6469, P2_U6470, P2_U6471, P2_U6472, P2_U6473, P2_U6474, P2_U6475, P2_U6476, P2_U6477, P2_U6478, P2_U6479, P2_U6480, P2_U6481, P2_U6482, P2_U6483, P2_U6484, P2_U6485, P2_U6486, P2_U6487, P2_U6488, P2_U6489, P2_U6490, P2_U6491, P2_U6492, P2_U6493, P2_U6494, P2_U6495, P2_U6496, P2_U6497, P2_U6498, P2_U6499, P2_U6500, P2_U6501, P2_U6502, P2_U6503, P2_U6504, P2_U6505, P2_U6506, P2_U6507, P2_U6508, P2_U6509, P2_U6510, P2_U6511, P2_U6512, P2_U6513, P2_U6514, P2_U6515, P2_U6516, P2_U6517, P2_U6518, P2_U6519, P2_U6520, P2_U6521, P2_U6522, P2_U6523, P2_U6524, P2_U6525, P2_U6526, P2_U6527, P2_U6528, P2_U6529, P2_U6530, P2_U6531, P2_U6532, P2_U6533, P2_U6534, P2_U6535, P2_U6536, P2_U6537, P2_U6538, P2_U6539, P2_U6540, P2_U6541, P2_U6542, P2_U6543, P2_U6544, P2_U6545, P2_U6546, P2_U6547, P2_U6548, P2_U6549, P2_U6550, P2_U6551, P2_U6552, P2_U6553, P2_U6554, P2_U6555, P2_U6556, P2_U6557, P2_U6558, P2_U6559, P2_U6560, P2_U6561, P2_U6562, P2_U6563, P2_U6564, P2_U6565, P2_U6566, P2_U6567, P2_U6568, P2_U6569, P2_U6570, P2_U6571, P2_U6572, P2_U6573, P2_U6574, P2_U6575, P2_U6576, P2_U6577, P2_U6578, P2_U6579, P2_U6580, P2_U6581, P2_U6582, P2_U6583, P2_U6584, P2_U6585, P2_U6586, P2_U6587, P2_U6588, P2_U6589, P2_U6590, P2_U6591, P2_U6592, P2_U6593, P2_U6594, P2_U6595, P2_U6596, P2_U6597, P2_U6598, P2_U6599, P2_U6600, P2_U6601, P2_U6602, P2_U6603, P2_U6604, P2_U6605, P2_U6606, P2_U6607, P2_U6608, P2_U6609, P2_U6610, P2_U6611, P2_U6612, P2_U6613, P2_U6614, P2_U6615, P2_U6616, P2_U6617, P2_U6618, P2_U6619, P2_U6620, P2_U6621, P2_U6622, P2_U6623, P2_U6624, P2_U6625, P2_U6626, P2_U6627, P2_U6628, P2_U6629, P2_U6630, P2_U6631, P2_U6632, P2_U6633, P2_U6634, P2_U6635, P2_U6636, P2_U6637, P2_U6638, P2_U6639, P2_U6640, P2_U6641, P2_U6642, P2_U6643, P2_U6644, P2_U6645, P2_U6646, P2_U6647, P2_U6648, P2_U6649, P2_U6650, P2_U6651, P2_U6652, P2_U6653, P2_U6654, P2_U6655, P2_U6656, P2_U6657, P2_U6658, P2_U6659, P2_U6660, P2_U6661, P2_U6662, P2_U6663, P2_U6664, P2_U6665, P2_U6666, P2_U6667, P2_U6668, P2_U6669, P2_U6670, P2_U6671, P2_U6672, P2_U6673, P2_U6674, P2_U6675, P2_U6676, P2_U6677, P2_U6678, P2_U6679, P2_U6680, P2_U6681, P2_U6682, P2_U6683, P2_U6684, P2_U6685, P2_U6686, P2_U6687, P2_U6688, P2_U6689, P2_U6690, P2_U6691, P2_U6692, P2_U6693, P2_U6694, P2_U6695, P2_U6696, P2_U6697, P2_U6698, P2_U6699, P2_U6700, P2_U6701, P2_U6702, P2_U6703, P2_U6704, P2_U6705, P2_U6706, P2_U6707, P2_U6708, P2_U6709, P2_U6710, P2_U6711, P2_U6712, P2_U6713, P2_U6714, P2_U6715, P2_U6716, P2_U6717, P2_U6718, P2_U6719, P2_U6720, P2_U6721, P2_U6722, P2_U6723, P2_U6724, P2_U6725, P2_U6726, P2_U6727, P2_U6728, P2_U6729, P2_U6730, P2_U6731, P2_U6732, P2_U6733, P2_U6734, P2_U6735, P2_U6736, P2_U6737, P2_U6738, P2_U6739, P2_U6740, P2_U6741, P2_U6742, P2_U6743, P2_U6744, P2_U6745, P2_U6746, P2_U6747, P2_U6748, P2_U6749, P2_U6750, P2_U6751, P2_U6752, P2_U6753, P2_U6754, P2_U6755, P2_U6756, P2_U6757, P2_U6758, P2_U6759, P2_U6760, P2_U6761, P2_U6762, P2_U6763, P2_U6764, P2_U6765, P2_U6766, P2_U6767, P2_U6768, P2_U6769, P2_U6770, P2_U6771, P2_U6772, P2_U6773, P2_U6774, P2_U6775, P2_U6776, P2_U6777, P2_U6778, P2_U6779, P2_U6780, P2_U6781, P2_U6782, P2_U6783, P2_U6784, P2_U6785, P2_U6786, P2_U6787, P2_U6788, P2_U6789, P2_U6790, P2_U6791, P2_U6792, P2_U6793, P2_U6794, P2_U6795, P2_U6796, P2_U6797, P2_U6798, P2_U6799, P2_U6800, P2_U6801, P2_U6802, P2_U6803, P2_U6804, P2_U6805, P2_U6806, P2_U6807, P2_U6808, P2_U6809, P2_U6810, P2_U6811, P2_U6812, P2_U6813, P2_U6814, P2_U6815, P2_U6816, P2_U6817, P2_U6818, P2_U6819, P2_U6820, P2_U6821, P2_U6822, P2_U6823, P2_U6824, P2_U6825, P2_U6826, P2_U6827, P2_U6828, P2_U6829, P2_U6830, P2_U6831, P2_U6832, P2_U6833, P2_U6834, P2_U6835, P2_U6836, P2_U6837, P2_U6838, P2_U6839, P2_U6840, P2_U6841, P2_U6842, P2_U6843, P2_U6844, P2_U6845, P2_U6846, P2_U6847, P2_U6848, P2_U6849, P2_U6850, P2_U6851, P2_U6852, P2_U6853, P2_U6854, P2_U6855, P2_U6856, P2_U6857, P2_U6858, P2_U6859, P2_U6860, P2_U6861, P2_U6862, P2_U6863, P2_U6864, P2_U6865, P2_U6866, P2_U6867, P2_U6868, P2_U6869, P2_U6870, P2_U6871, P2_U6872, P2_U6873, P2_U6874, P2_U6875, P2_U6876, P2_U6877, P2_U6878, P2_U6879, P2_U6880, P2_U6881, P2_U6882, P2_U6883, P2_U6884, P2_U6885, P2_U6886, P2_U6887, P2_U6888, P2_U6889, P2_U6890, P2_U6891, P2_U6892, P2_U6893, P2_U6894, P2_U6895, P2_U6896, P2_U6897, P2_U6898, P2_U6899, P2_U6900, P2_U6901, P2_U6902, P2_U6903, P2_U6904, P2_U6905, P2_U6906, P2_U6907, P2_U6908, P2_U6909, P2_U6910, P2_U6911, P2_U6912, P2_U6913, P2_U6914, P2_U6915, P2_U6916, P2_U6917, P2_U6918, P2_U6919, P2_U6920, P2_U6921, P2_U6922, P2_U6923, P2_U6924, P2_U6925, P2_U6926, P2_U6927, P2_U6928, P2_U6929, P2_U6930, P2_U6931, P2_U6932, P2_U6933, P2_U6934, P2_U6935, P2_U6936, P2_U6937, P2_U6938, P2_U6939, P2_U6940, P2_U6941, P2_U6942, P2_U6943, P2_U6944, P2_U6945, P2_U6946, P2_U6947, P2_U6948, P2_U6949, P2_U6950, P2_U6951, P2_U6952, P2_U6953, P2_U6954, P2_U6955, P2_U6956, P2_U6957, P2_U6958, P2_U6959, P2_U6960, P2_U6961, P2_U6962, P2_U6963, P2_U6964, P2_U6965, P2_U6966, P2_U6967, P2_U6968, P2_U6969, P2_U6970, P2_U6971, P2_U6972, P2_U6973, P2_U6974, P2_U6975, P2_U6976, P2_U6977, P2_U6978, P2_U6979, P2_U6980, P2_U6981, P2_U6982, P2_U6983, P2_U6984, P2_U6985, P2_U6986, P2_U6987, P2_U6988, P2_U6989, P2_U6990, P2_U6991, P2_U6992, P2_U6993, P2_U6994, P2_U6995, P2_U6996, P2_U6997, P2_U6998, P2_U6999, P2_U7000, P2_U7001, P2_U7002, P2_U7003, P2_U7004, P2_U7005, P2_U7006, P2_U7007, P2_U7008, P2_U7009, P2_U7010, P2_U7011, P2_U7012, P2_U7013, P2_U7014, P2_U7015, P2_U7016, P2_U7017, P2_U7018, P2_U7019, P2_U7020, P2_U7021, P2_U7022, P2_U7023, P2_U7024, P2_U7025, P2_U7026, P2_U7027, P2_U7028, P2_U7029, P2_U7030, P2_U7031, P2_U7032, P2_U7033, P2_U7034, P2_U7035, P2_U7036, P2_U7037, P2_U7038, P2_U7039, P2_U7040, P2_U7041, P2_U7042, P2_U7043, P2_U7044, P2_U7045, P2_U7046, P2_U7047, P2_U7048, P2_U7049, P2_U7050, P2_U7051, P2_U7052, P2_U7053, P2_U7054, P2_U7055, P2_U7056, P2_U7057, P2_U7058, P2_U7059, P2_U7060, P2_U7061, P2_U7062, P2_U7063, P2_U7064, P2_U7065, P2_U7066, P2_U7067, P2_U7068, P2_U7069, P2_U7070, P2_U7071, P2_U7072, P2_U7073, P2_U7074, P2_U7075, P2_U7076, P2_U7077, P2_U7078, P2_U7079, P2_U7080, P2_U7081, P2_U7082, P2_U7083, P2_U7084, P2_U7085, P2_U7086, P2_U7087, P2_U7088, P2_U7089, P2_U7090, P2_U7091, P2_U7092, P2_U7093, P2_U7094, P2_U7095, P2_U7096, P2_U7097, P2_U7098, P2_U7099, P2_U7100, P2_U7101, P2_U7102, P2_U7103, P2_U7104, P2_U7105, P2_U7106, P2_U7107, P2_U7108, P2_U7109, P2_U7110, P2_U7111, P2_U7112, P2_U7113, P2_U7114, P2_U7115, P2_U7116, P2_U7117, P2_U7118, P2_U7119, P2_U7120, P2_U7121, P2_U7122, P2_U7123, P2_U7124, P2_U7125, P2_U7126, P2_U7127, P2_U7128, P2_U7129, P2_U7130, P2_U7131, P2_U7132, P2_U7133, P2_U7134, P2_U7135, P2_U7136, P2_U7137, P2_U7138, P2_U7139, P2_U7140, P2_U7141, P2_U7142, P2_U7143, P2_U7144, P2_U7145, P2_U7146, P2_U7147, P2_U7148, P2_U7149, P2_U7150, P2_U7151, P2_U7152, P2_U7153, P2_U7154, P2_U7155, P2_U7156, P2_U7157, P2_U7158, P2_U7159, P2_U7160, P2_U7161, P2_U7162, P2_U7163, P2_U7164, P2_U7165, P2_U7166, P2_U7167, P2_U7168, P2_U7169, P2_U7170, P2_U7171, P2_U7172, P2_U7173, P2_U7174, P2_U7175, P2_U7176, P2_U7177, P2_U7178, P2_U7179, P2_U7180, P2_U7181, P2_U7182, P2_U7183, P2_U7184, P2_U7185, P2_U7186, P2_U7187, P2_U7188, P2_U7189, P2_U7190, P2_U7191, P2_U7192, P2_U7193, P2_U7194, P2_U7195, P2_U7196, P2_U7197, P2_U7198, P2_U7199, P2_U7200, P2_U7201, P2_U7202, P2_U7203, P2_U7204, P2_U7205, P2_U7206, P2_U7207, P2_U7208, P2_U7209, P2_U7210, P2_U7211, P2_U7212, P2_U7213, P2_U7214, P2_U7215, P2_U7216, P2_U7217, P2_U7218, P2_U7219, P2_U7220, P2_U7221, P2_U7222, P2_U7223, P2_U7224, P2_U7225, P2_U7226, P2_U7227, P2_U7228, P2_U7229, P2_U7230, P2_U7231, P2_U7232, P2_U7233, P2_U7234, P2_U7235, P2_U7236, P2_U7237, P2_U7238, P2_U7239, P2_U7240, P2_U7241, P2_U7242, P2_U7243, P2_U7244, P2_U7245, P2_U7246, P2_U7247, P2_U7248, P2_U7249, P2_U7250, P2_U7251, P2_U7252, P2_U7253, P2_U7254, P2_U7255, P2_U7256, P2_U7257, P2_U7258, P2_U7259, P2_U7260, P2_U7261, P2_U7262, P2_U7263, P2_U7264, P2_U7265, P2_U7266, P2_U7267, P2_U7268, P2_U7269, P2_U7270, P2_U7271, P2_U7272, P2_U7273, P2_U7274, P2_U7275, P2_U7276, P2_U7277, P2_U7278, P2_U7279, P2_U7280, P2_U7281, P2_U7282, P2_U7283, P2_U7284, P2_U7285, P2_U7286, P2_U7287, P2_U7288, P2_U7289, P2_U7290, P2_U7291, P2_U7292, P2_U7293, P2_U7294, P2_U7295, P2_U7296, P2_U7297, P2_U7298, P2_U7299, P2_U7300, P2_U7301, P2_U7302, P2_U7303, P2_U7304, P2_U7305, P2_U7306, P2_U7307, P2_U7308, P2_U7309, P2_U7310, P2_U7311, P2_U7312, P2_U7313, P2_U7314, P2_U7315, P2_U7316, P2_U7317, P2_U7318, P2_U7319, P2_U7320, P2_U7321, P2_U7322, P2_U7323, P2_U7324, P2_U7325, P2_U7326, P2_U7327, P2_U7328, P2_U7329, P2_U7330, P2_U7331, P2_U7332, P2_U7333, P2_U7334, P2_U7335, P2_U7336, P2_U7337, P2_U7338, P2_U7339, P2_U7340, P2_U7341, P2_U7342, P2_U7343, P2_U7344, P2_U7345, P2_U7346, P2_U7347, P2_U7348, P2_U7349, P2_U7350, P2_U7351, P2_U7352, P2_U7353, P2_U7354, P2_U7355, P2_U7356, P2_U7357, P2_U7358, P2_U7359, P2_U7360, P2_U7361, P2_U7362, P2_U7363, P2_U7364, P2_U7365, P2_U7366, P2_U7367, P2_U7368, P2_U7369, P2_U7370, P2_U7371, P2_U7372, P2_U7373, P2_U7374, P2_U7375, P2_U7376, P2_U7377, P2_U7378, P2_U7379, P2_U7380, P2_U7381, P2_U7382, P2_U7383, P2_U7384, P2_U7385, P2_U7386, P2_U7387, P2_U7388, P2_U7389, P2_U7390, P2_U7391, P2_U7392, P2_U7393, P2_U7394, P2_U7395, P2_U7396, P2_U7397, P2_U7398, P2_U7399, P2_U7400, P2_U7401, P2_U7402, P2_U7403, P2_U7404, P2_U7405, P2_U7406, P2_U7407, P2_U7408, P2_U7409, P2_U7410, P2_U7411, P2_U7412, P2_U7413, P2_U7414, P2_U7415, P2_U7416, P2_U7417, P2_U7418, P2_U7419, P2_U7420, P2_U7421, P2_U7422, P2_U7423, P2_U7424, P2_U7425, P2_U7426, P2_U7427, P2_U7428, P2_U7429, P2_U7430, P2_U7431, P2_U7432, P2_U7433, P2_U7434, P2_U7435, P2_U7436, P2_U7437, P2_U7438, P2_U7439, P2_U7440, P2_U7441, P2_U7442, P2_U7443, P2_U7444, P2_U7445, P2_U7446, P2_U7447, P2_U7448, P2_U7449, P2_U7450, P2_U7451, P2_U7452, P2_U7453, P2_U7454, P2_U7455, P2_U7456, P2_U7457, P2_U7458, P2_U7459, P2_U7460, P2_U7461, P2_U7462, P2_U7463, P2_U7464, P2_U7465, P2_U7466, P2_U7467, P2_U7468, P2_U7469, P2_U7470, P2_U7471, P2_U7472, P2_U7473, P2_U7474, P2_U7475, P2_U7476, P2_U7477, P2_U7478, P2_U7479, P2_U7480, P2_U7481, P2_U7482, P2_U7483, P2_U7484, P2_U7485, P2_U7486, P2_U7487, P2_U7488, P2_U7489, P2_U7490, P2_U7491, P2_U7492, P2_U7493, P2_U7494, P2_U7495, P2_U7496, P2_U7497, P2_U7498, P2_U7499, P2_U7500, P2_U7501, P2_U7502, P2_U7503, P2_U7504, P2_U7505, P2_U7506, P2_U7507, P2_U7508, P2_U7509, P2_U7510, P2_U7511, P2_U7512, P2_U7513, P2_U7514, P2_U7515, P2_U7516, P2_U7517, P2_U7518, P2_U7519, P2_U7520, P2_U7521, P2_U7522, P2_U7523, P2_U7524, P2_U7525, P2_U7526, P2_U7527, P2_U7528, P2_U7529, P2_U7530, P2_U7531, P2_U7532, P2_U7533, P2_U7534, P2_U7535, P2_U7536, P2_U7537, P2_U7538, P2_U7539, P2_U7540, P2_U7541, P2_U7542, P2_U7543, P2_U7544, P2_U7545, P2_U7546, P2_U7547, P2_U7548, P2_U7549, P2_U7550, P2_U7551, P2_U7552, P2_U7553, P2_U7554, P2_U7555, P2_U7556, P2_U7557, P2_U7558, P2_U7559, P2_U7560, P2_U7561, P2_U7562, P2_U7563, P2_U7564, P2_U7565, P2_U7566, P2_U7567, P2_U7568, P2_U7569, P2_U7570, P2_U7571, P2_U7572, P2_U7573, P2_U7574, P2_U7575, P2_U7576, P2_U7577, P2_U7578, P2_U7579, P2_U7580, P2_U7581, P2_U7582, P2_U7583, P2_U7584, P2_U7585, P2_U7586, P2_U7587, P2_U7588, P2_U7589, P2_U7590, P2_U7591, P2_U7592, P2_U7593, P2_U7594, P2_U7595, P2_U7596, P2_U7597, P2_U7598, P2_U7599, P2_U7600, P2_U7601, P2_U7602, P2_U7603, P2_U7604, P2_U7605, P2_U7606, P2_U7607, P2_U7608, P2_U7609, P2_U7610, P2_U7611, P2_U7612, P2_U7613, P2_U7614, P2_U7615, P2_U7616, P2_U7617, P2_U7618, P2_U7619, P2_U7620, P2_U7621, P2_U7622, P2_U7623, P2_U7624, P2_U7625, P2_U7626, P2_U7627, P2_U7628, P2_U7629, P2_U7630, P2_U7631, P2_U7632, P2_U7633, P2_U7634, P2_U7635, P2_U7636, P2_U7637, P2_U7638, P2_U7639, P2_U7640, P2_U7641, P2_U7642, P2_U7643, P2_U7644, P2_U7645, P2_U7646, P2_U7647, P2_U7648, P2_U7649, P2_U7650, P2_U7651, P2_U7652, P2_U7653, P2_U7654, P2_U7655, P2_U7656, P2_U7657, P2_U7658, P2_U7659, P2_U7660, P2_U7661, P2_U7662, P2_U7663, P2_U7664, P2_U7665, P2_U7666, P2_U7667, P2_U7668, P2_U7669, P2_U7670, P2_U7671, P2_U7672, P2_U7673, P2_U7674, P2_U7675, P2_U7676, P2_U7677, P2_U7678, P2_U7679, P2_U7680, P2_U7681, P2_U7682, P2_U7683, P2_U7684, P2_U7685, P2_U7686, P2_U7687, P2_U7688, P2_U7689, P2_U7690, P2_U7691, P2_U7692, P2_U7693, P2_U7694, P2_U7695, P2_U7696, P2_U7697, P2_U7698, P2_U7699, P2_U7700, P2_U7701, P2_U7702, P2_U7703, P2_U7704, P2_U7705, P2_U7706, P2_U7707, P2_U7708, P2_U7709, P2_U7710, P2_U7711, P2_U7712, P2_U7713, P2_U7714, P2_U7715, P2_U7716, P2_U7717, P2_U7718, P2_U7719, P2_U7720, P2_U7721, P2_U7722, P2_U7723, P2_U7724, P2_U7725, P2_U7726, P2_U7727, P2_U7728, P2_U7729, P2_U7730, P2_U7731, P2_U7732, P2_U7733, P2_U7734, P2_U7735, P2_U7736, P2_U7737, P2_U7738, P2_U7739, P2_U7740, P2_U7741, P2_U7742, P2_U7743, P2_U7744, P2_U7745, P2_U7746, P2_U7747, P2_U7748, P2_U7749, P2_U7750, P2_U7751, P2_U7752, P2_U7753, P2_U7754, P2_U7755, P2_U7756, P2_U7757, P2_U7758, P2_U7759, P2_U7760, P2_U7761, P2_U7762, P2_U7763, P2_U7764, P2_U7765, P2_U7766, P2_U7767, P2_U7768, P2_U7769, P2_U7770, P2_U7771, P2_U7772, P2_U7773, P2_U7774, P2_U7775, P2_U7776, P2_U7777, P2_U7778, P2_U7779, P2_U7780, P2_U7781, P2_U7782, P2_U7783, P2_U7784, P2_U7785, P2_U7786, P2_U7787, P2_U7788, P2_U7789, P2_U7790, P2_U7791, P2_U7792, P2_U7793, P2_U7794, P2_U7795, P2_U7796, P2_U7797, P2_U7798, P2_U7799, P2_U7800, P2_U7801, P2_U7802, P2_U7803, P2_U7804, P2_U7805, P2_U7806, P2_U7807, P2_U7808, P2_U7809, P2_U7810, P2_U7811, P2_U7812, P2_U7813, P2_U7814, P2_U7815, P2_U7816, P2_U7817, P2_U7818, P2_U7819, P2_U7820, P2_U7821, P2_U7822, P2_U7823, P2_U7824, P2_U7825, P2_U7826, P2_U7827, P2_U7828, P2_U7829, P2_U7830, P2_U7831, P2_U7832, P2_U7833, P2_U7834, P2_U7835, P2_U7836, P2_U7837, P2_U7838, P2_U7839, P2_U7840, P2_U7841, P2_U7842, P2_U7843, P2_U7844, P2_U7845, P2_U7846, P2_U7847, P2_U7848, P2_U7849, P2_U7850, P2_U7851, P2_U7852, P2_U7853, P2_U7854, P2_U7855, P2_U7856, P2_U7857, P2_U7858, P2_U7859, P2_U7860, P2_U7861, P2_U7862, P2_U7863, P2_U7864, P2_U7865, P2_U7866, P2_U7867, P2_U7868, P2_U7869, P2_U7870, P2_U7871, P2_U7872, P2_U7873, P2_U7874, P2_U7875, P2_U7876, P2_U7877, P2_U7878, P2_U7879, P2_U7880, P2_U7881, P2_U7882, P2_U7883, P2_U7884, P2_U7885, P2_U7886, P2_U7887, P2_U7888, P2_U7889, P2_U7890, P2_U7891, P2_U7892, P2_U7893, P2_U7894, P2_U7895, P2_U7896, P2_U7897, P2_U7898, P2_U7899, P2_U7900, P2_U7901, P2_U7902, P2_U7903, P2_U7904, P2_U7905, P2_U7906, P2_U7907, P2_U7908, P2_U7909, P2_U7910, P2_U7911, P2_U7912, P2_U7913, P2_U7914, P2_U7915, P2_U7916, P2_U7917, P2_U7918, P2_U7919, P2_U7920, P2_U7921, P2_U7922, P2_U7923, P2_U7924, P2_U7925, P2_U7926, P2_U7927, P2_U7928, P2_U7929, P2_U7930, P2_U7931, P2_U7932, P2_U7933, P2_U7934, P2_U7935, P2_U7936, P2_U7937, P2_U7938, P2_U7939, P2_U7940, P2_U7941, P2_U7942, P2_U7943, P2_U7944, P2_U7945, P2_U7946, P2_U7947, P2_U7948, P2_U7949, P2_U7950, P2_U7951, P2_U7952, P2_U7953, P2_U7954, P2_U7955, P2_U7956, P2_U7957, P2_U7958, P2_U7959, P2_U7960, P2_U7961, P2_U7962, P2_U7963, P2_U7964, P2_U7965, P2_U7966, P2_U7967, P2_U7968, P2_U7969, P2_U7970, P2_U7971, P2_U7972, P2_U7973, P2_U7974, P2_U7975, P2_U7976, P2_U7977, P2_U7978, P2_U7979, P2_U7980, P2_U7981, P2_U7982, P2_U7983, P2_U7984, P2_U7985, P2_U7986, P2_U7987, P2_U7988, P2_U7989, P2_U7990, P2_U7991, P2_U7992, P2_U7993, P2_U7994, P2_U7995, P2_U7996, P2_U7997, P2_U7998, P2_U7999, P2_U8000, P2_U8001, P2_U8002, P2_U8003, P2_U8004, P2_U8005, P2_U8006, P2_U8007, P2_U8008, P2_U8009, P2_U8010, P2_U8011, P2_U8012, P2_U8013, P2_U8014, P2_U8015, P2_U8016, P2_U8017, P2_U8018, P2_U8019, P2_U8020, P2_U8021, P2_U8022, P2_U8023, P2_U8024, P2_U8025, P2_U8026, P2_U8027, P2_U8028, P2_U8029, P2_U8030, P2_U8031, P2_U8032, P2_U8033, P2_U8034, P2_U8035, P2_U8036, P2_U8037, P2_U8038, P2_U8039, P2_U8040, P2_U8041, P2_U8042, P2_U8043, P2_U8044, P2_U8045, P2_U8046, P2_U8047, P2_U8048, P2_U8049, P2_U8050, P2_U8051, P2_U8052, P2_U8053, P2_U8054, P2_U8055, P2_U8056, P2_U8057, P2_U8058, P2_U8059, P2_U8060, P2_U8061, P2_U8062, P2_U8063, P2_U8064, P2_U8065, P2_U8066, P2_U8067, P2_U8068, P2_U8069, P2_U8070, P2_U8071, P2_U8072, P2_U8073, P2_U8074, P2_U8075, P2_U8076, P2_U8077, P2_U8078, P2_U8079, P2_U8080, P2_U8081, P2_U8082, P2_U8083, P2_U8084, P2_U8085, P2_U8086, P2_U8087, P2_U8088, P2_U8089, P2_U8090, P2_U8091, P2_U8092, P2_U8093, P2_U8094, P2_U8095, P2_U8096, P2_U8097, P2_U8098, P2_U8099, P2_U8100, P2_U8101, P2_U8102, P2_U8103, P2_U8104, P2_U8105, P2_U8106, P2_U8107, P2_U8108, P2_U8109, P2_U8110, P2_U8111, P2_U8112, P2_U8113, P2_U8114, P2_U8115, P2_U8116, P2_U8117, P2_U8118, P2_U8119, P2_U8120, P2_U8121, P2_U8122, P2_U8123, P2_U8124, P2_U8125, P2_U8126, P2_U8127, P2_U8128, P2_U8129, P2_U8130, P2_U8131, P2_U8132, P2_U8133, P2_U8134, P2_U8135, P2_U8136, P2_U8137, P2_U8138, P2_U8139, P2_U8140, P2_U8141, P2_U8142, P2_U8143, P2_U8144, P2_U8145, P2_U8146, P2_U8147, P2_U8148, P2_U8149, P2_U8150, P2_U8151, P2_U8152, P2_U8153, P2_U8154, P2_U8155, P2_U8156, P2_U8157, P2_U8158, P2_U8159, P2_U8160, P2_U8161, P2_U8162, P2_U8163, P2_U8164, P2_U8165, P2_U8166, P2_U8167, P2_U8168, P2_U8169, P2_U8170, P2_U8171, P2_U8172, P2_U8173, P2_U8174, P2_U8175, P2_U8176, P2_U8177, P2_U8178, P2_U8179, P2_U8180, P2_U8181, P2_U8182, P2_U8183, P2_U8184, P2_U8185, P2_U8186, P2_U8187, P2_U8188, P2_U8189, P2_U8190, P2_U8191, P2_U8192, P2_U8193, P2_U8194, P2_U8195, P2_U8196, P2_U8197, P2_U8198, P2_U8199, P2_U8200, P2_U8201, P2_U8202, P2_U8203, P2_U8204, P2_U8205, P2_U8206, P2_U8207, P2_U8208, P2_U8209, P2_U8210, P2_U8211, P2_U8212, P2_U8213, P2_U8214, P2_U8215, P2_U8216, P2_U8217, P2_U8218, P2_U8219, P2_U8220, P2_U8221, P2_U8222, P2_U8223, P2_U8224, P2_U8225, P2_U8226, P2_U8227, P2_U8228, P2_U8229, P2_U8230, P2_U8231, P2_U8232, P2_U8233, P2_U8234, P2_U8235, P2_U8236, P2_U8237, P2_U8238, P2_U8239, P2_U8240, P2_U8241, P2_U8242, P2_U8243, P2_U8244, P2_U8245, P2_U8246, P2_U8247, P2_U8248, P2_U8249, P2_U8250, P2_U8251, P2_U8252, P2_U8253, P2_U8254, P2_U8255, P2_U8256, P2_U8257, P2_U8258, P2_U8259, P2_U8260, P2_U8261, P2_U8262, P2_U8263, P2_U8264, P2_U8265, P2_U8266, P2_U8267, P2_U8268, P2_U8269, P2_U8270, P2_U8271, P2_U8272, P2_U8273, P2_U8274, P2_U8275, P2_U8276, P2_U8277, P2_U8278, P2_U8279, P2_U8280, P2_U8281, P2_U8282, P2_U8283, P2_U8284, P2_U8285, P2_U8286, P2_U8287, P2_U8288, P2_U8289, P2_U8290, P2_U8291, P2_U8292, P2_U8293, P2_U8294, P2_U8295, P2_U8296, P2_U8297, P2_U8298, P2_U8299, P2_U8300, P2_U8301, P2_U8302, P2_U8303, P2_U8304, P2_U8305, P2_U8306, P2_U8307, P2_U8308, P2_U8309, P2_U8310, P2_U8311, P2_U8312, P2_U8313, P2_U8314, P2_U8315, P2_U8316, P2_U8317, P2_U8318, P2_U8319, P2_U8320, P2_U8321, P2_U8322, P2_U8323, P2_U8324, P2_U8325, P2_U8326, P2_U8327, P2_U8328, P2_U8329, P2_U8330, P2_U8331, P2_U8332, P2_U8333, P2_U8334, P2_U8335, P2_U8336, P2_U8337, P2_U8338, P2_U8339, P2_U8340, P2_U8341, P2_U8342, P2_U8343, P2_U8344, P2_U8345, P2_U8346, P2_U8347, P2_U8348, P2_U8349, P2_U8350, P2_U8351, P2_U8352, P2_U8353, P2_U8354, P2_U8355, P2_U8356, P2_U8357, P2_U8358, P2_U8359, P2_U8360, P2_U8361, P2_U8362, P2_U8363, P2_U8364, P2_U8365, P2_U8366, P2_U8367, P2_U8368, P2_U8369, P2_U8370, P2_U8371, P2_U8372, P2_U8373, P2_U8374, P2_U8375, P2_U8376, P2_U8377, P2_U8378, P2_U8379, P2_U8380, P2_U8381, P2_U8382, P2_U8383, P2_U8384, P2_U8385, P2_U8386, P2_U8387, P2_U8388, P2_U8389, P2_U8390, P2_U8391, P2_U8392, P2_U8393, P2_U8394, P2_U8395, P2_U8396, P2_U8397, P2_U8398, P2_U8399, P2_U8400, P2_U8401, P2_U8402, P2_U8403, P2_U8404, P2_U8405, P2_U8406, P2_U8407, P2_U8408, P2_U8409, P2_U8410, P2_U8411, P2_U8412, P2_U8413, P2_U8414, P2_U8415, P2_U8416, P2_U8417, P2_U8418, P2_U8419, P2_U8420, P2_U8421, P2_U8422, P2_U8423, P2_U8424, P2_U8425, P2_U8426, P2_U8427, P2_U8428, P2_U8429, P2_U8430, P2_U8431, P2_U8432, P2_U8433, P2_U8434, P3_ADD_315_U10, P3_ADD_315_U100, P3_ADD_315_U101, P3_ADD_315_U102, P3_ADD_315_U103, P3_ADD_315_U104, P3_ADD_315_U105, P3_ADD_315_U106, P3_ADD_315_U107, P3_ADD_315_U108, P3_ADD_315_U109, P3_ADD_315_U11, P3_ADD_315_U110, P3_ADD_315_U111, P3_ADD_315_U112, P3_ADD_315_U113, P3_ADD_315_U114, P3_ADD_315_U115, P3_ADD_315_U116, P3_ADD_315_U117, P3_ADD_315_U118, P3_ADD_315_U119, P3_ADD_315_U12, P3_ADD_315_U120, P3_ADD_315_U121, P3_ADD_315_U122, P3_ADD_315_U123, P3_ADD_315_U124, P3_ADD_315_U125, P3_ADD_315_U126, P3_ADD_315_U127, P3_ADD_315_U128, P3_ADD_315_U129, P3_ADD_315_U13, P3_ADD_315_U130, P3_ADD_315_U131, P3_ADD_315_U132, P3_ADD_315_U133, P3_ADD_315_U134, P3_ADD_315_U135, P3_ADD_315_U136, P3_ADD_315_U137, P3_ADD_315_U138, P3_ADD_315_U139, P3_ADD_315_U14, P3_ADD_315_U140, P3_ADD_315_U141, P3_ADD_315_U142, P3_ADD_315_U143, P3_ADD_315_U144, P3_ADD_315_U145, P3_ADD_315_U146, P3_ADD_315_U147, P3_ADD_315_U148, P3_ADD_315_U149, P3_ADD_315_U15, P3_ADD_315_U150, P3_ADD_315_U151, P3_ADD_315_U152, P3_ADD_315_U153, P3_ADD_315_U154, P3_ADD_315_U155, P3_ADD_315_U156, P3_ADD_315_U157, P3_ADD_315_U158, P3_ADD_315_U159, P3_ADD_315_U16, P3_ADD_315_U160, P3_ADD_315_U161, P3_ADD_315_U162, P3_ADD_315_U163, P3_ADD_315_U164, P3_ADD_315_U165, P3_ADD_315_U166, P3_ADD_315_U167, P3_ADD_315_U168, P3_ADD_315_U169, P3_ADD_315_U17, P3_ADD_315_U170, P3_ADD_315_U171, P3_ADD_315_U172, P3_ADD_315_U173, P3_ADD_315_U174, P3_ADD_315_U175, P3_ADD_315_U176, P3_ADD_315_U18, P3_ADD_315_U19, P3_ADD_315_U20, P3_ADD_315_U21, P3_ADD_315_U22, P3_ADD_315_U23, P3_ADD_315_U24, P3_ADD_315_U25, P3_ADD_315_U26, P3_ADD_315_U27, P3_ADD_315_U28, P3_ADD_315_U29, P3_ADD_315_U30, P3_ADD_315_U31, P3_ADD_315_U32, P3_ADD_315_U33, P3_ADD_315_U34, P3_ADD_315_U35, P3_ADD_315_U36, P3_ADD_315_U37, P3_ADD_315_U38, P3_ADD_315_U39, P3_ADD_315_U4, P3_ADD_315_U40, P3_ADD_315_U41, P3_ADD_315_U42, P3_ADD_315_U43, P3_ADD_315_U44, P3_ADD_315_U45, P3_ADD_315_U46, P3_ADD_315_U47, P3_ADD_315_U48, P3_ADD_315_U49, P3_ADD_315_U5, P3_ADD_315_U50, P3_ADD_315_U51, P3_ADD_315_U52, P3_ADD_315_U53, P3_ADD_315_U54, P3_ADD_315_U55, P3_ADD_315_U56, P3_ADD_315_U57, P3_ADD_315_U58, P3_ADD_315_U59, P3_ADD_315_U6, P3_ADD_315_U60, P3_ADD_315_U61, P3_ADD_315_U62, P3_ADD_315_U63, P3_ADD_315_U64, P3_ADD_315_U65, P3_ADD_315_U66, P3_ADD_315_U67, P3_ADD_315_U68, P3_ADD_315_U69, P3_ADD_315_U7, P3_ADD_315_U70, P3_ADD_315_U71, P3_ADD_315_U72, P3_ADD_315_U73, P3_ADD_315_U74, P3_ADD_315_U75, P3_ADD_315_U76, P3_ADD_315_U77, P3_ADD_315_U78, P3_ADD_315_U79, P3_ADD_315_U8, P3_ADD_315_U80, P3_ADD_315_U81, P3_ADD_315_U82, P3_ADD_315_U83, P3_ADD_315_U84, P3_ADD_315_U85, P3_ADD_315_U86, P3_ADD_315_U87, P3_ADD_315_U88, P3_ADD_315_U89, P3_ADD_315_U9, P3_ADD_315_U90, P3_ADD_315_U91, P3_ADD_315_U92, P3_ADD_315_U93, P3_ADD_315_U94, P3_ADD_315_U95, P3_ADD_315_U96, P3_ADD_315_U97, P3_ADD_315_U98, P3_ADD_315_U99, P3_ADD_318_U10, P3_ADD_318_U100, P3_ADD_318_U101, P3_ADD_318_U102, P3_ADD_318_U103, P3_ADD_318_U104, P3_ADD_318_U105, P3_ADD_318_U106, P3_ADD_318_U107, P3_ADD_318_U108, P3_ADD_318_U109, P3_ADD_318_U11, P3_ADD_318_U110, P3_ADD_318_U111, P3_ADD_318_U112, P3_ADD_318_U113, P3_ADD_318_U114, P3_ADD_318_U115, P3_ADD_318_U116, P3_ADD_318_U117, P3_ADD_318_U118, P3_ADD_318_U119, P3_ADD_318_U12, P3_ADD_318_U120, P3_ADD_318_U121, P3_ADD_318_U122, P3_ADD_318_U123, P3_ADD_318_U124, P3_ADD_318_U125, P3_ADD_318_U126, P3_ADD_318_U127, P3_ADD_318_U128, P3_ADD_318_U129, P3_ADD_318_U13, P3_ADD_318_U130, P3_ADD_318_U131, P3_ADD_318_U132, P3_ADD_318_U133, P3_ADD_318_U134, P3_ADD_318_U135, P3_ADD_318_U136, P3_ADD_318_U137, P3_ADD_318_U138, P3_ADD_318_U139, P3_ADD_318_U14, P3_ADD_318_U140, P3_ADD_318_U141, P3_ADD_318_U142, P3_ADD_318_U143, P3_ADD_318_U144, P3_ADD_318_U145, P3_ADD_318_U146, P3_ADD_318_U147, P3_ADD_318_U148, P3_ADD_318_U149, P3_ADD_318_U15, P3_ADD_318_U150, P3_ADD_318_U151, P3_ADD_318_U152, P3_ADD_318_U153, P3_ADD_318_U154, P3_ADD_318_U155, P3_ADD_318_U156, P3_ADD_318_U157, P3_ADD_318_U158, P3_ADD_318_U159, P3_ADD_318_U16, P3_ADD_318_U160, P3_ADD_318_U161, P3_ADD_318_U162, P3_ADD_318_U163, P3_ADD_318_U164, P3_ADD_318_U165, P3_ADD_318_U166, P3_ADD_318_U167, P3_ADD_318_U168, P3_ADD_318_U169, P3_ADD_318_U17, P3_ADD_318_U170, P3_ADD_318_U171, P3_ADD_318_U172, P3_ADD_318_U173, P3_ADD_318_U174, P3_ADD_318_U175, P3_ADD_318_U176, P3_ADD_318_U177, P3_ADD_318_U178, P3_ADD_318_U179, P3_ADD_318_U18, P3_ADD_318_U180, P3_ADD_318_U181, P3_ADD_318_U182, P3_ADD_318_U19, P3_ADD_318_U20, P3_ADD_318_U21, P3_ADD_318_U22, P3_ADD_318_U23, P3_ADD_318_U24, P3_ADD_318_U25, P3_ADD_318_U26, P3_ADD_318_U27, P3_ADD_318_U28, P3_ADD_318_U29, P3_ADD_318_U30, P3_ADD_318_U31, P3_ADD_318_U32, P3_ADD_318_U33, P3_ADD_318_U34, P3_ADD_318_U35, P3_ADD_318_U36, P3_ADD_318_U37, P3_ADD_318_U38, P3_ADD_318_U39, P3_ADD_318_U4, P3_ADD_318_U40, P3_ADD_318_U41, P3_ADD_318_U42, P3_ADD_318_U43, P3_ADD_318_U44, P3_ADD_318_U45, P3_ADD_318_U46, P3_ADD_318_U47, P3_ADD_318_U48, P3_ADD_318_U49, P3_ADD_318_U5, P3_ADD_318_U50, P3_ADD_318_U51, P3_ADD_318_U52, P3_ADD_318_U53, P3_ADD_318_U54, P3_ADD_318_U55, P3_ADD_318_U56, P3_ADD_318_U57, P3_ADD_318_U58, P3_ADD_318_U59, P3_ADD_318_U6, P3_ADD_318_U60, P3_ADD_318_U61, P3_ADD_318_U62, P3_ADD_318_U63, P3_ADD_318_U64, P3_ADD_318_U65, P3_ADD_318_U66, P3_ADD_318_U67, P3_ADD_318_U68, P3_ADD_318_U69, P3_ADD_318_U7, P3_ADD_318_U70, P3_ADD_318_U71, P3_ADD_318_U72, P3_ADD_318_U73, P3_ADD_318_U74, P3_ADD_318_U75, P3_ADD_318_U76, P3_ADD_318_U77, P3_ADD_318_U78, P3_ADD_318_U79, P3_ADD_318_U8, P3_ADD_318_U80, P3_ADD_318_U81, P3_ADD_318_U82, P3_ADD_318_U83, P3_ADD_318_U84, P3_ADD_318_U85, P3_ADD_318_U86, P3_ADD_318_U87, P3_ADD_318_U88, P3_ADD_318_U89, P3_ADD_318_U9, P3_ADD_318_U90, P3_ADD_318_U91, P3_ADD_318_U92, P3_ADD_318_U93, P3_ADD_318_U94, P3_ADD_318_U95, P3_ADD_318_U96, P3_ADD_318_U97, P3_ADD_318_U98, P3_ADD_318_U99, P3_ADD_339_U10, P3_ADD_339_U100, P3_ADD_339_U101, P3_ADD_339_U102, P3_ADD_339_U103, P3_ADD_339_U104, P3_ADD_339_U105, P3_ADD_339_U106, P3_ADD_339_U107, P3_ADD_339_U108, P3_ADD_339_U109, P3_ADD_339_U11, P3_ADD_339_U110, P3_ADD_339_U111, P3_ADD_339_U112, P3_ADD_339_U113, P3_ADD_339_U114, P3_ADD_339_U115, P3_ADD_339_U116, P3_ADD_339_U117, P3_ADD_339_U118, P3_ADD_339_U119, P3_ADD_339_U12, P3_ADD_339_U120, P3_ADD_339_U121, P3_ADD_339_U122, P3_ADD_339_U123, P3_ADD_339_U124, P3_ADD_339_U125, P3_ADD_339_U126, P3_ADD_339_U127, P3_ADD_339_U128, P3_ADD_339_U129, P3_ADD_339_U13, P3_ADD_339_U130, P3_ADD_339_U131, P3_ADD_339_U132, P3_ADD_339_U133, P3_ADD_339_U134, P3_ADD_339_U135, P3_ADD_339_U136, P3_ADD_339_U137, P3_ADD_339_U138, P3_ADD_339_U139, P3_ADD_339_U14, P3_ADD_339_U140, P3_ADD_339_U141, P3_ADD_339_U142, P3_ADD_339_U143, P3_ADD_339_U144, P3_ADD_339_U145, P3_ADD_339_U146, P3_ADD_339_U147, P3_ADD_339_U148, P3_ADD_339_U149, P3_ADD_339_U15, P3_ADD_339_U150, P3_ADD_339_U151, P3_ADD_339_U152, P3_ADD_339_U153, P3_ADD_339_U154, P3_ADD_339_U155, P3_ADD_339_U156, P3_ADD_339_U157, P3_ADD_339_U158, P3_ADD_339_U159, P3_ADD_339_U16, P3_ADD_339_U160, P3_ADD_339_U161, P3_ADD_339_U162, P3_ADD_339_U163, P3_ADD_339_U164, P3_ADD_339_U165, P3_ADD_339_U166, P3_ADD_339_U167, P3_ADD_339_U168, P3_ADD_339_U169, P3_ADD_339_U17, P3_ADD_339_U170, P3_ADD_339_U171, P3_ADD_339_U172, P3_ADD_339_U173, P3_ADD_339_U174, P3_ADD_339_U175, P3_ADD_339_U176, P3_ADD_339_U177, P3_ADD_339_U178, P3_ADD_339_U179, P3_ADD_339_U18, P3_ADD_339_U180, P3_ADD_339_U181, P3_ADD_339_U182, P3_ADD_339_U19, P3_ADD_339_U20, P3_ADD_339_U21, P3_ADD_339_U22, P3_ADD_339_U23, P3_ADD_339_U24, P3_ADD_339_U25, P3_ADD_339_U26, P3_ADD_339_U27, P3_ADD_339_U28, P3_ADD_339_U29, P3_ADD_339_U30, P3_ADD_339_U31, P3_ADD_339_U32, P3_ADD_339_U33, P3_ADD_339_U34, P3_ADD_339_U35, P3_ADD_339_U36, P3_ADD_339_U37, P3_ADD_339_U38, P3_ADD_339_U39, P3_ADD_339_U4, P3_ADD_339_U40, P3_ADD_339_U41, P3_ADD_339_U42, P3_ADD_339_U43, P3_ADD_339_U44, P3_ADD_339_U45, P3_ADD_339_U46, P3_ADD_339_U47, P3_ADD_339_U48, P3_ADD_339_U49, P3_ADD_339_U5, P3_ADD_339_U50, P3_ADD_339_U51, P3_ADD_339_U52, P3_ADD_339_U53, P3_ADD_339_U54, P3_ADD_339_U55, P3_ADD_339_U56, P3_ADD_339_U57, P3_ADD_339_U58, P3_ADD_339_U59, P3_ADD_339_U6, P3_ADD_339_U60, P3_ADD_339_U61, P3_ADD_339_U62, P3_ADD_339_U63, P3_ADD_339_U64, P3_ADD_339_U65, P3_ADD_339_U66, P3_ADD_339_U67, P3_ADD_339_U68, P3_ADD_339_U69, P3_ADD_339_U7, P3_ADD_339_U70, P3_ADD_339_U71, P3_ADD_339_U72, P3_ADD_339_U73, P3_ADD_339_U74, P3_ADD_339_U75, P3_ADD_339_U76, P3_ADD_339_U77, P3_ADD_339_U78, P3_ADD_339_U79, P3_ADD_339_U8, P3_ADD_339_U80, P3_ADD_339_U81, P3_ADD_339_U82, P3_ADD_339_U83, P3_ADD_339_U84, P3_ADD_339_U85, P3_ADD_339_U86, P3_ADD_339_U87, P3_ADD_339_U88, P3_ADD_339_U89, P3_ADD_339_U9, P3_ADD_339_U90, P3_ADD_339_U91, P3_ADD_339_U92, P3_ADD_339_U93, P3_ADD_339_U94, P3_ADD_339_U95, P3_ADD_339_U96, P3_ADD_339_U97, P3_ADD_339_U98, P3_ADD_339_U99, P3_ADD_344_U10, P3_ADD_344_U100, P3_ADD_344_U101, P3_ADD_344_U102, P3_ADD_344_U103, P3_ADD_344_U104, P3_ADD_344_U105, P3_ADD_344_U106, P3_ADD_344_U107, P3_ADD_344_U108, P3_ADD_344_U109, P3_ADD_344_U11, P3_ADD_344_U110, P3_ADD_344_U111, P3_ADD_344_U112, P3_ADD_344_U113, P3_ADD_344_U114, P3_ADD_344_U115, P3_ADD_344_U116, P3_ADD_344_U117, P3_ADD_344_U118, P3_ADD_344_U119, P3_ADD_344_U12, P3_ADD_344_U120, P3_ADD_344_U121, P3_ADD_344_U122, P3_ADD_344_U123, P3_ADD_344_U124, P3_ADD_344_U125, P3_ADD_344_U126, P3_ADD_344_U127, P3_ADD_344_U128, P3_ADD_344_U129, P3_ADD_344_U13, P3_ADD_344_U130, P3_ADD_344_U131, P3_ADD_344_U132, P3_ADD_344_U133, P3_ADD_344_U134, P3_ADD_344_U135, P3_ADD_344_U136, P3_ADD_344_U137, P3_ADD_344_U138, P3_ADD_344_U139, P3_ADD_344_U14, P3_ADD_344_U140, P3_ADD_344_U141, P3_ADD_344_U142, P3_ADD_344_U143, P3_ADD_344_U144, P3_ADD_344_U145, P3_ADD_344_U146, P3_ADD_344_U147, P3_ADD_344_U148, P3_ADD_344_U149, P3_ADD_344_U15, P3_ADD_344_U150, P3_ADD_344_U151, P3_ADD_344_U152, P3_ADD_344_U153, P3_ADD_344_U154, P3_ADD_344_U155, P3_ADD_344_U156, P3_ADD_344_U157, P3_ADD_344_U158, P3_ADD_344_U159, P3_ADD_344_U16, P3_ADD_344_U160, P3_ADD_344_U161, P3_ADD_344_U162, P3_ADD_344_U163, P3_ADD_344_U164, P3_ADD_344_U165, P3_ADD_344_U166, P3_ADD_344_U167, P3_ADD_344_U168, P3_ADD_344_U169, P3_ADD_344_U17, P3_ADD_344_U170, P3_ADD_344_U171, P3_ADD_344_U172, P3_ADD_344_U173, P3_ADD_344_U174, P3_ADD_344_U175, P3_ADD_344_U176, P3_ADD_344_U177, P3_ADD_344_U178, P3_ADD_344_U179, P3_ADD_344_U18, P3_ADD_344_U180, P3_ADD_344_U181, P3_ADD_344_U182, P3_ADD_344_U183, P3_ADD_344_U184, P3_ADD_344_U185, P3_ADD_344_U186, P3_ADD_344_U187, P3_ADD_344_U188, P3_ADD_344_U189, P3_ADD_344_U19, P3_ADD_344_U20, P3_ADD_344_U21, P3_ADD_344_U22, P3_ADD_344_U23, P3_ADD_344_U24, P3_ADD_344_U25, P3_ADD_344_U26, P3_ADD_344_U27, P3_ADD_344_U28, P3_ADD_344_U29, P3_ADD_344_U30, P3_ADD_344_U31, P3_ADD_344_U32, P3_ADD_344_U33, P3_ADD_344_U34, P3_ADD_344_U35, P3_ADD_344_U36, P3_ADD_344_U37, P3_ADD_344_U38, P3_ADD_344_U39, P3_ADD_344_U40, P3_ADD_344_U41, P3_ADD_344_U42, P3_ADD_344_U43, P3_ADD_344_U44, P3_ADD_344_U45, P3_ADD_344_U46, P3_ADD_344_U47, P3_ADD_344_U48, P3_ADD_344_U49, P3_ADD_344_U5, P3_ADD_344_U50, P3_ADD_344_U51, P3_ADD_344_U52, P3_ADD_344_U53, P3_ADD_344_U54, P3_ADD_344_U55, P3_ADD_344_U56, P3_ADD_344_U57, P3_ADD_344_U58, P3_ADD_344_U59, P3_ADD_344_U6, P3_ADD_344_U60, P3_ADD_344_U61, P3_ADD_344_U62, P3_ADD_344_U63, P3_ADD_344_U64, P3_ADD_344_U65, P3_ADD_344_U66, P3_ADD_344_U67, P3_ADD_344_U68, P3_ADD_344_U69, P3_ADD_344_U7, P3_ADD_344_U70, P3_ADD_344_U71, P3_ADD_344_U72, P3_ADD_344_U73, P3_ADD_344_U74, P3_ADD_344_U75, P3_ADD_344_U76, P3_ADD_344_U77, P3_ADD_344_U78, P3_ADD_344_U79, P3_ADD_344_U8, P3_ADD_344_U80, P3_ADD_344_U81, P3_ADD_344_U82, P3_ADD_344_U83, P3_ADD_344_U84, P3_ADD_344_U85, P3_ADD_344_U86, P3_ADD_344_U87, P3_ADD_344_U88, P3_ADD_344_U89, P3_ADD_344_U9, P3_ADD_344_U90, P3_ADD_344_U91, P3_ADD_344_U92, P3_ADD_344_U93, P3_ADD_344_U94, P3_ADD_344_U95, P3_ADD_344_U96, P3_ADD_344_U97, P3_ADD_344_U98, P3_ADD_344_U99, P3_ADD_349_U10, P3_ADD_349_U100, P3_ADD_349_U101, P3_ADD_349_U102, P3_ADD_349_U103, P3_ADD_349_U104, P3_ADD_349_U105, P3_ADD_349_U106, P3_ADD_349_U107, P3_ADD_349_U108, P3_ADD_349_U109, P3_ADD_349_U11, P3_ADD_349_U110, P3_ADD_349_U111, P3_ADD_349_U112, P3_ADD_349_U113, P3_ADD_349_U114, P3_ADD_349_U115, P3_ADD_349_U116, P3_ADD_349_U117, P3_ADD_349_U118, P3_ADD_349_U119, P3_ADD_349_U12, P3_ADD_349_U120, P3_ADD_349_U121, P3_ADD_349_U122, P3_ADD_349_U123, P3_ADD_349_U124, P3_ADD_349_U125, P3_ADD_349_U126, P3_ADD_349_U127, P3_ADD_349_U128, P3_ADD_349_U129, P3_ADD_349_U13, P3_ADD_349_U130, P3_ADD_349_U131, P3_ADD_349_U132, P3_ADD_349_U133, P3_ADD_349_U134, P3_ADD_349_U135, P3_ADD_349_U136, P3_ADD_349_U137, P3_ADD_349_U138, P3_ADD_349_U139, P3_ADD_349_U14, P3_ADD_349_U140, P3_ADD_349_U141, P3_ADD_349_U142, P3_ADD_349_U143, P3_ADD_349_U144, P3_ADD_349_U145, P3_ADD_349_U146, P3_ADD_349_U147, P3_ADD_349_U148, P3_ADD_349_U149, P3_ADD_349_U15, P3_ADD_349_U150, P3_ADD_349_U151, P3_ADD_349_U152, P3_ADD_349_U153, P3_ADD_349_U154, P3_ADD_349_U155, P3_ADD_349_U156, P3_ADD_349_U157, P3_ADD_349_U158, P3_ADD_349_U159, P3_ADD_349_U16, P3_ADD_349_U160, P3_ADD_349_U161, P3_ADD_349_U162, P3_ADD_349_U163, P3_ADD_349_U164, P3_ADD_349_U165, P3_ADD_349_U166, P3_ADD_349_U167, P3_ADD_349_U168, P3_ADD_349_U169, P3_ADD_349_U17, P3_ADD_349_U170, P3_ADD_349_U171, P3_ADD_349_U172, P3_ADD_349_U173, P3_ADD_349_U174, P3_ADD_349_U175, P3_ADD_349_U176, P3_ADD_349_U177, P3_ADD_349_U178, P3_ADD_349_U179, P3_ADD_349_U18, P3_ADD_349_U180, P3_ADD_349_U181, P3_ADD_349_U182, P3_ADD_349_U183, P3_ADD_349_U184, P3_ADD_349_U185, P3_ADD_349_U186, P3_ADD_349_U187, P3_ADD_349_U188, P3_ADD_349_U189, P3_ADD_349_U19, P3_ADD_349_U20, P3_ADD_349_U21, P3_ADD_349_U22, P3_ADD_349_U23, P3_ADD_349_U24, P3_ADD_349_U25, P3_ADD_349_U26, P3_ADD_349_U27, P3_ADD_349_U28, P3_ADD_349_U29, P3_ADD_349_U30, P3_ADD_349_U31, P3_ADD_349_U32, P3_ADD_349_U33, P3_ADD_349_U34, P3_ADD_349_U35, P3_ADD_349_U36, P3_ADD_349_U37, P3_ADD_349_U38, P3_ADD_349_U39, P3_ADD_349_U40, P3_ADD_349_U41, P3_ADD_349_U42, P3_ADD_349_U43, P3_ADD_349_U44, P3_ADD_349_U45, P3_ADD_349_U46, P3_ADD_349_U47, P3_ADD_349_U48, P3_ADD_349_U49, P3_ADD_349_U5, P3_ADD_349_U50, P3_ADD_349_U51, P3_ADD_349_U52, P3_ADD_349_U53, P3_ADD_349_U54, P3_ADD_349_U55, P3_ADD_349_U56, P3_ADD_349_U57, P3_ADD_349_U58, P3_ADD_349_U59, P3_ADD_349_U6, P3_ADD_349_U60, P3_ADD_349_U61, P3_ADD_349_U62, P3_ADD_349_U63, P3_ADD_349_U64, P3_ADD_349_U65, P3_ADD_349_U66, P3_ADD_349_U67, P3_ADD_349_U68, P3_ADD_349_U69, P3_ADD_349_U7, P3_ADD_349_U70, P3_ADD_349_U71, P3_ADD_349_U72, P3_ADD_349_U73, P3_ADD_349_U74, P3_ADD_349_U75, P3_ADD_349_U76, P3_ADD_349_U77, P3_ADD_349_U78, P3_ADD_349_U79, P3_ADD_349_U8, P3_ADD_349_U80, P3_ADD_349_U81, P3_ADD_349_U82, P3_ADD_349_U83, P3_ADD_349_U84, P3_ADD_349_U85, P3_ADD_349_U86, P3_ADD_349_U87, P3_ADD_349_U88, P3_ADD_349_U89, P3_ADD_349_U9, P3_ADD_349_U90, P3_ADD_349_U91, P3_ADD_349_U92, P3_ADD_349_U93, P3_ADD_349_U94, P3_ADD_349_U95, P3_ADD_349_U96, P3_ADD_349_U97, P3_ADD_349_U98, P3_ADD_349_U99, P3_ADD_357_U10, P3_ADD_357_U11, P3_ADD_357_U12, P3_ADD_357_U13, P3_ADD_357_U14, P3_ADD_357_U15, P3_ADD_357_U16, P3_ADD_357_U17, P3_ADD_357_U18, P3_ADD_357_U19, P3_ADD_357_U20, P3_ADD_357_U21, P3_ADD_357_U22, P3_ADD_357_U23, P3_ADD_357_U24, P3_ADD_357_U25, P3_ADD_357_U26, P3_ADD_357_U27, P3_ADD_357_U28, P3_ADD_357_U29, P3_ADD_357_U30, P3_ADD_357_U31, P3_ADD_357_U32, P3_ADD_357_U33, P3_ADD_357_U34, P3_ADD_357_U35, P3_ADD_357_U6, P3_ADD_357_U7, P3_ADD_357_U8, P3_ADD_357_U9, P3_ADD_360_1242_U10, P3_ADD_360_1242_U100, P3_ADD_360_1242_U101, P3_ADD_360_1242_U102, P3_ADD_360_1242_U103, P3_ADD_360_1242_U104, P3_ADD_360_1242_U105, P3_ADD_360_1242_U106, P3_ADD_360_1242_U107, P3_ADD_360_1242_U108, P3_ADD_360_1242_U109, P3_ADD_360_1242_U11, P3_ADD_360_1242_U110, P3_ADD_360_1242_U111, P3_ADD_360_1242_U112, P3_ADD_360_1242_U113, P3_ADD_360_1242_U114, P3_ADD_360_1242_U115, P3_ADD_360_1242_U116, P3_ADD_360_1242_U117, P3_ADD_360_1242_U118, P3_ADD_360_1242_U119, P3_ADD_360_1242_U12, P3_ADD_360_1242_U120, P3_ADD_360_1242_U121, P3_ADD_360_1242_U122, P3_ADD_360_1242_U123, P3_ADD_360_1242_U124, P3_ADD_360_1242_U125, P3_ADD_360_1242_U126, P3_ADD_360_1242_U127, P3_ADD_360_1242_U128, P3_ADD_360_1242_U129, P3_ADD_360_1242_U13, P3_ADD_360_1242_U130, P3_ADD_360_1242_U131, P3_ADD_360_1242_U132, P3_ADD_360_1242_U133, P3_ADD_360_1242_U134, P3_ADD_360_1242_U135, P3_ADD_360_1242_U136, P3_ADD_360_1242_U137, P3_ADD_360_1242_U138, P3_ADD_360_1242_U139, P3_ADD_360_1242_U14, P3_ADD_360_1242_U140, P3_ADD_360_1242_U141, P3_ADD_360_1242_U142, P3_ADD_360_1242_U143, P3_ADD_360_1242_U144, P3_ADD_360_1242_U145, P3_ADD_360_1242_U146, P3_ADD_360_1242_U147, P3_ADD_360_1242_U148, P3_ADD_360_1242_U149, P3_ADD_360_1242_U15, P3_ADD_360_1242_U150, P3_ADD_360_1242_U151, P3_ADD_360_1242_U152, P3_ADD_360_1242_U153, P3_ADD_360_1242_U154, P3_ADD_360_1242_U155, P3_ADD_360_1242_U156, P3_ADD_360_1242_U157, P3_ADD_360_1242_U158, P3_ADD_360_1242_U159, P3_ADD_360_1242_U16, P3_ADD_360_1242_U160, P3_ADD_360_1242_U161, P3_ADD_360_1242_U162, P3_ADD_360_1242_U163, P3_ADD_360_1242_U164, P3_ADD_360_1242_U165, P3_ADD_360_1242_U166, P3_ADD_360_1242_U167, P3_ADD_360_1242_U168, P3_ADD_360_1242_U169, P3_ADD_360_1242_U17, P3_ADD_360_1242_U170, P3_ADD_360_1242_U171, P3_ADD_360_1242_U172, P3_ADD_360_1242_U173, P3_ADD_360_1242_U174, P3_ADD_360_1242_U175, P3_ADD_360_1242_U176, P3_ADD_360_1242_U177, P3_ADD_360_1242_U178, P3_ADD_360_1242_U179, P3_ADD_360_1242_U18, P3_ADD_360_1242_U180, P3_ADD_360_1242_U181, P3_ADD_360_1242_U182, P3_ADD_360_1242_U183, P3_ADD_360_1242_U184, P3_ADD_360_1242_U185, P3_ADD_360_1242_U186, P3_ADD_360_1242_U187, P3_ADD_360_1242_U188, P3_ADD_360_1242_U189, P3_ADD_360_1242_U19, P3_ADD_360_1242_U190, P3_ADD_360_1242_U191, P3_ADD_360_1242_U192, P3_ADD_360_1242_U193, P3_ADD_360_1242_U194, P3_ADD_360_1242_U195, P3_ADD_360_1242_U196, P3_ADD_360_1242_U197, P3_ADD_360_1242_U198, P3_ADD_360_1242_U199, P3_ADD_360_1242_U20, P3_ADD_360_1242_U200, P3_ADD_360_1242_U201, P3_ADD_360_1242_U202, P3_ADD_360_1242_U203, P3_ADD_360_1242_U204, P3_ADD_360_1242_U205, P3_ADD_360_1242_U206, P3_ADD_360_1242_U207, P3_ADD_360_1242_U208, P3_ADD_360_1242_U209, P3_ADD_360_1242_U21, P3_ADD_360_1242_U210, P3_ADD_360_1242_U211, P3_ADD_360_1242_U212, P3_ADD_360_1242_U213, P3_ADD_360_1242_U214, P3_ADD_360_1242_U215, P3_ADD_360_1242_U216, P3_ADD_360_1242_U217, P3_ADD_360_1242_U218, P3_ADD_360_1242_U219, P3_ADD_360_1242_U22, P3_ADD_360_1242_U220, P3_ADD_360_1242_U221, P3_ADD_360_1242_U222, P3_ADD_360_1242_U223, P3_ADD_360_1242_U224, P3_ADD_360_1242_U225, P3_ADD_360_1242_U226, P3_ADD_360_1242_U227, P3_ADD_360_1242_U228, P3_ADD_360_1242_U229, P3_ADD_360_1242_U23, P3_ADD_360_1242_U230, P3_ADD_360_1242_U231, P3_ADD_360_1242_U232, P3_ADD_360_1242_U233, P3_ADD_360_1242_U234, P3_ADD_360_1242_U235, P3_ADD_360_1242_U236, P3_ADD_360_1242_U237, P3_ADD_360_1242_U238, P3_ADD_360_1242_U239, P3_ADD_360_1242_U24, P3_ADD_360_1242_U240, P3_ADD_360_1242_U241, P3_ADD_360_1242_U242, P3_ADD_360_1242_U243, P3_ADD_360_1242_U244, P3_ADD_360_1242_U245, P3_ADD_360_1242_U246, P3_ADD_360_1242_U247, P3_ADD_360_1242_U248, P3_ADD_360_1242_U249, P3_ADD_360_1242_U25, P3_ADD_360_1242_U250, P3_ADD_360_1242_U251, P3_ADD_360_1242_U252, P3_ADD_360_1242_U253, P3_ADD_360_1242_U254, P3_ADD_360_1242_U255, P3_ADD_360_1242_U256, P3_ADD_360_1242_U257, P3_ADD_360_1242_U258, P3_ADD_360_1242_U26, P3_ADD_360_1242_U27, P3_ADD_360_1242_U28, P3_ADD_360_1242_U29, P3_ADD_360_1242_U30, P3_ADD_360_1242_U31, P3_ADD_360_1242_U32, P3_ADD_360_1242_U33, P3_ADD_360_1242_U34, P3_ADD_360_1242_U35, P3_ADD_360_1242_U36, P3_ADD_360_1242_U37, P3_ADD_360_1242_U38, P3_ADD_360_1242_U39, P3_ADD_360_1242_U4, P3_ADD_360_1242_U40, P3_ADD_360_1242_U41, P3_ADD_360_1242_U42, P3_ADD_360_1242_U43, P3_ADD_360_1242_U44, P3_ADD_360_1242_U45, P3_ADD_360_1242_U46, P3_ADD_360_1242_U47, P3_ADD_360_1242_U48, P3_ADD_360_1242_U49, P3_ADD_360_1242_U5, P3_ADD_360_1242_U50, P3_ADD_360_1242_U51, P3_ADD_360_1242_U52, P3_ADD_360_1242_U53, P3_ADD_360_1242_U54, P3_ADD_360_1242_U55, P3_ADD_360_1242_U56, P3_ADD_360_1242_U57, P3_ADD_360_1242_U58, P3_ADD_360_1242_U59, P3_ADD_360_1242_U6, P3_ADD_360_1242_U60, P3_ADD_360_1242_U61, P3_ADD_360_1242_U62, P3_ADD_360_1242_U63, P3_ADD_360_1242_U64, P3_ADD_360_1242_U65, P3_ADD_360_1242_U66, P3_ADD_360_1242_U67, P3_ADD_360_1242_U68, P3_ADD_360_1242_U69, P3_ADD_360_1242_U7, P3_ADD_360_1242_U70, P3_ADD_360_1242_U71, P3_ADD_360_1242_U72, P3_ADD_360_1242_U73, P3_ADD_360_1242_U74, P3_ADD_360_1242_U75, P3_ADD_360_1242_U76, P3_ADD_360_1242_U77, P3_ADD_360_1242_U78, P3_ADD_360_1242_U79, P3_ADD_360_1242_U8, P3_ADD_360_1242_U80, P3_ADD_360_1242_U81, P3_ADD_360_1242_U82, P3_ADD_360_1242_U83, P3_ADD_360_1242_U84, P3_ADD_360_1242_U85, P3_ADD_360_1242_U86, P3_ADD_360_1242_U87, P3_ADD_360_1242_U88, P3_ADD_360_1242_U89, P3_ADD_360_1242_U9, P3_ADD_360_1242_U90, P3_ADD_360_1242_U91, P3_ADD_360_1242_U92, P3_ADD_360_1242_U93, P3_ADD_360_1242_U94, P3_ADD_360_1242_U95, P3_ADD_360_1242_U96, P3_ADD_360_1242_U97, P3_ADD_360_1242_U98, P3_ADD_360_1242_U99, P3_ADD_360_U10, P3_ADD_360_U11, P3_ADD_360_U12, P3_ADD_360_U13, P3_ADD_360_U14, P3_ADD_360_U15, P3_ADD_360_U16, P3_ADD_360_U17, P3_ADD_360_U18, P3_ADD_360_U19, P3_ADD_360_U20, P3_ADD_360_U21, P3_ADD_360_U22, P3_ADD_360_U23, P3_ADD_360_U24, P3_ADD_360_U25, P3_ADD_360_U26, P3_ADD_360_U27, P3_ADD_360_U28, P3_ADD_360_U29, P3_ADD_360_U30, P3_ADD_360_U31, P3_ADD_360_U32, P3_ADD_360_U33, P3_ADD_360_U34, P3_ADD_360_U35, P3_ADD_360_U36, P3_ADD_360_U37, P3_ADD_360_U38, P3_ADD_360_U39, P3_ADD_360_U4, P3_ADD_360_U40, P3_ADD_360_U5, P3_ADD_360_U6, P3_ADD_360_U7, P3_ADD_360_U8, P3_ADD_360_U9, P3_ADD_371_1212_U10, P3_ADD_371_1212_U100, P3_ADD_371_1212_U101, P3_ADD_371_1212_U102, P3_ADD_371_1212_U103, P3_ADD_371_1212_U104, P3_ADD_371_1212_U105, P3_ADD_371_1212_U106, P3_ADD_371_1212_U107, P3_ADD_371_1212_U108, P3_ADD_371_1212_U109, P3_ADD_371_1212_U11, P3_ADD_371_1212_U110, P3_ADD_371_1212_U111, P3_ADD_371_1212_U112, P3_ADD_371_1212_U113, P3_ADD_371_1212_U114, P3_ADD_371_1212_U115, P3_ADD_371_1212_U116, P3_ADD_371_1212_U117, P3_ADD_371_1212_U118, P3_ADD_371_1212_U119, P3_ADD_371_1212_U12, P3_ADD_371_1212_U120, P3_ADD_371_1212_U121, P3_ADD_371_1212_U122, P3_ADD_371_1212_U123, P3_ADD_371_1212_U124, P3_ADD_371_1212_U125, P3_ADD_371_1212_U126, P3_ADD_371_1212_U127, P3_ADD_371_1212_U128, P3_ADD_371_1212_U129, P3_ADD_371_1212_U13, P3_ADD_371_1212_U130, P3_ADD_371_1212_U131, P3_ADD_371_1212_U132, P3_ADD_371_1212_U133, P3_ADD_371_1212_U134, P3_ADD_371_1212_U135, P3_ADD_371_1212_U136, P3_ADD_371_1212_U137, P3_ADD_371_1212_U138, P3_ADD_371_1212_U139, P3_ADD_371_1212_U14, P3_ADD_371_1212_U140, P3_ADD_371_1212_U141, P3_ADD_371_1212_U142, P3_ADD_371_1212_U143, P3_ADD_371_1212_U144, P3_ADD_371_1212_U145, P3_ADD_371_1212_U146, P3_ADD_371_1212_U147, P3_ADD_371_1212_U148, P3_ADD_371_1212_U149, P3_ADD_371_1212_U15, P3_ADD_371_1212_U150, P3_ADD_371_1212_U151, P3_ADD_371_1212_U152, P3_ADD_371_1212_U153, P3_ADD_371_1212_U154, P3_ADD_371_1212_U155, P3_ADD_371_1212_U156, P3_ADD_371_1212_U157, P3_ADD_371_1212_U158, P3_ADD_371_1212_U159, P3_ADD_371_1212_U16, P3_ADD_371_1212_U160, P3_ADD_371_1212_U161, P3_ADD_371_1212_U162, P3_ADD_371_1212_U163, P3_ADD_371_1212_U164, P3_ADD_371_1212_U165, P3_ADD_371_1212_U166, P3_ADD_371_1212_U167, P3_ADD_371_1212_U168, P3_ADD_371_1212_U169, P3_ADD_371_1212_U17, P3_ADD_371_1212_U170, P3_ADD_371_1212_U171, P3_ADD_371_1212_U172, P3_ADD_371_1212_U173, P3_ADD_371_1212_U174, P3_ADD_371_1212_U175, P3_ADD_371_1212_U176, P3_ADD_371_1212_U177, P3_ADD_371_1212_U178, P3_ADD_371_1212_U179, P3_ADD_371_1212_U18, P3_ADD_371_1212_U180, P3_ADD_371_1212_U181, P3_ADD_371_1212_U182, P3_ADD_371_1212_U183, P3_ADD_371_1212_U184, P3_ADD_371_1212_U185, P3_ADD_371_1212_U186, P3_ADD_371_1212_U187, P3_ADD_371_1212_U188, P3_ADD_371_1212_U189, P3_ADD_371_1212_U19, P3_ADD_371_1212_U190, P3_ADD_371_1212_U191, P3_ADD_371_1212_U192, P3_ADD_371_1212_U193, P3_ADD_371_1212_U194, P3_ADD_371_1212_U195, P3_ADD_371_1212_U196, P3_ADD_371_1212_U197, P3_ADD_371_1212_U198, P3_ADD_371_1212_U199, P3_ADD_371_1212_U20, P3_ADD_371_1212_U200, P3_ADD_371_1212_U201, P3_ADD_371_1212_U202, P3_ADD_371_1212_U203, P3_ADD_371_1212_U204, P3_ADD_371_1212_U205, P3_ADD_371_1212_U206, P3_ADD_371_1212_U207, P3_ADD_371_1212_U208, P3_ADD_371_1212_U209, P3_ADD_371_1212_U21, P3_ADD_371_1212_U210, P3_ADD_371_1212_U211, P3_ADD_371_1212_U212, P3_ADD_371_1212_U213, P3_ADD_371_1212_U214, P3_ADD_371_1212_U215, P3_ADD_371_1212_U216, P3_ADD_371_1212_U217, P3_ADD_371_1212_U218, P3_ADD_371_1212_U219, P3_ADD_371_1212_U22, P3_ADD_371_1212_U220, P3_ADD_371_1212_U221, P3_ADD_371_1212_U222, P3_ADD_371_1212_U223, P3_ADD_371_1212_U224, P3_ADD_371_1212_U225, P3_ADD_371_1212_U226, P3_ADD_371_1212_U227, P3_ADD_371_1212_U228, P3_ADD_371_1212_U229, P3_ADD_371_1212_U23, P3_ADD_371_1212_U230, P3_ADD_371_1212_U231, P3_ADD_371_1212_U232, P3_ADD_371_1212_U233, P3_ADD_371_1212_U234, P3_ADD_371_1212_U235, P3_ADD_371_1212_U236, P3_ADD_371_1212_U237, P3_ADD_371_1212_U238, P3_ADD_371_1212_U239, P3_ADD_371_1212_U24, P3_ADD_371_1212_U240, P3_ADD_371_1212_U241, P3_ADD_371_1212_U242, P3_ADD_371_1212_U243, P3_ADD_371_1212_U244, P3_ADD_371_1212_U245, P3_ADD_371_1212_U246, P3_ADD_371_1212_U247, P3_ADD_371_1212_U248, P3_ADD_371_1212_U249, P3_ADD_371_1212_U25, P3_ADD_371_1212_U250, P3_ADD_371_1212_U251, P3_ADD_371_1212_U252, P3_ADD_371_1212_U253, P3_ADD_371_1212_U254, P3_ADD_371_1212_U255, P3_ADD_371_1212_U256, P3_ADD_371_1212_U257, P3_ADD_371_1212_U258, P3_ADD_371_1212_U259, P3_ADD_371_1212_U26, P3_ADD_371_1212_U260, P3_ADD_371_1212_U261, P3_ADD_371_1212_U262, P3_ADD_371_1212_U263, P3_ADD_371_1212_U264, P3_ADD_371_1212_U265, P3_ADD_371_1212_U27, P3_ADD_371_1212_U28, P3_ADD_371_1212_U29, P3_ADD_371_1212_U30, P3_ADD_371_1212_U31, P3_ADD_371_1212_U32, P3_ADD_371_1212_U33, P3_ADD_371_1212_U34, P3_ADD_371_1212_U35, P3_ADD_371_1212_U36, P3_ADD_371_1212_U37, P3_ADD_371_1212_U38, P3_ADD_371_1212_U39, P3_ADD_371_1212_U4, P3_ADD_371_1212_U40, P3_ADD_371_1212_U41, P3_ADD_371_1212_U42, P3_ADD_371_1212_U43, P3_ADD_371_1212_U44, P3_ADD_371_1212_U45, P3_ADD_371_1212_U46, P3_ADD_371_1212_U47, P3_ADD_371_1212_U48, P3_ADD_371_1212_U49, P3_ADD_371_1212_U5, P3_ADD_371_1212_U50, P3_ADD_371_1212_U51, P3_ADD_371_1212_U52, P3_ADD_371_1212_U53, P3_ADD_371_1212_U54, P3_ADD_371_1212_U55, P3_ADD_371_1212_U56, P3_ADD_371_1212_U57, P3_ADD_371_1212_U58, P3_ADD_371_1212_U59, P3_ADD_371_1212_U6, P3_ADD_371_1212_U60, P3_ADD_371_1212_U61, P3_ADD_371_1212_U62, P3_ADD_371_1212_U63, P3_ADD_371_1212_U64, P3_ADD_371_1212_U65, P3_ADD_371_1212_U66, P3_ADD_371_1212_U67, P3_ADD_371_1212_U68, P3_ADD_371_1212_U69, P3_ADD_371_1212_U7, P3_ADD_371_1212_U70, P3_ADD_371_1212_U71, P3_ADD_371_1212_U72, P3_ADD_371_1212_U73, P3_ADD_371_1212_U74, P3_ADD_371_1212_U75, P3_ADD_371_1212_U76, P3_ADD_371_1212_U77, P3_ADD_371_1212_U78, P3_ADD_371_1212_U79, P3_ADD_371_1212_U8, P3_ADD_371_1212_U80, P3_ADD_371_1212_U81, P3_ADD_371_1212_U82, P3_ADD_371_1212_U83, P3_ADD_371_1212_U84, P3_ADD_371_1212_U85, P3_ADD_371_1212_U86, P3_ADD_371_1212_U87, P3_ADD_371_1212_U88, P3_ADD_371_1212_U89, P3_ADD_371_1212_U9, P3_ADD_371_1212_U90, P3_ADD_371_1212_U91, P3_ADD_371_1212_U92, P3_ADD_371_1212_U93, P3_ADD_371_1212_U94, P3_ADD_371_1212_U95, P3_ADD_371_1212_U96, P3_ADD_371_1212_U97, P3_ADD_371_1212_U98, P3_ADD_371_1212_U99, P3_ADD_371_U10, P3_ADD_371_U11, P3_ADD_371_U12, P3_ADD_371_U13, P3_ADD_371_U14, P3_ADD_371_U15, P3_ADD_371_U16, P3_ADD_371_U17, P3_ADD_371_U18, P3_ADD_371_U19, P3_ADD_371_U20, P3_ADD_371_U21, P3_ADD_371_U22, P3_ADD_371_U23, P3_ADD_371_U24, P3_ADD_371_U25, P3_ADD_371_U26, P3_ADD_371_U27, P3_ADD_371_U28, P3_ADD_371_U29, P3_ADD_371_U30, P3_ADD_371_U31, P3_ADD_371_U32, P3_ADD_371_U33, P3_ADD_371_U34, P3_ADD_371_U35, P3_ADD_371_U36, P3_ADD_371_U37, P3_ADD_371_U38, P3_ADD_371_U39, P3_ADD_371_U4, P3_ADD_371_U40, P3_ADD_371_U41, P3_ADD_371_U42, P3_ADD_371_U43, P3_ADD_371_U44, P3_ADD_371_U5, P3_ADD_371_U6, P3_ADD_371_U7, P3_ADD_371_U8, P3_ADD_371_U9, P3_ADD_380_U10, P3_ADD_380_U100, P3_ADD_380_U101, P3_ADD_380_U102, P3_ADD_380_U103, P3_ADD_380_U104, P3_ADD_380_U105, P3_ADD_380_U106, P3_ADD_380_U107, P3_ADD_380_U108, P3_ADD_380_U109, P3_ADD_380_U11, P3_ADD_380_U110, P3_ADD_380_U111, P3_ADD_380_U112, P3_ADD_380_U113, P3_ADD_380_U114, P3_ADD_380_U115, P3_ADD_380_U116, P3_ADD_380_U117, P3_ADD_380_U118, P3_ADD_380_U119, P3_ADD_380_U12, P3_ADD_380_U120, P3_ADD_380_U121, P3_ADD_380_U122, P3_ADD_380_U123, P3_ADD_380_U124, P3_ADD_380_U125, P3_ADD_380_U126, P3_ADD_380_U127, P3_ADD_380_U128, P3_ADD_380_U129, P3_ADD_380_U13, P3_ADD_380_U130, P3_ADD_380_U131, P3_ADD_380_U132, P3_ADD_380_U133, P3_ADD_380_U134, P3_ADD_380_U135, P3_ADD_380_U136, P3_ADD_380_U137, P3_ADD_380_U138, P3_ADD_380_U139, P3_ADD_380_U14, P3_ADD_380_U140, P3_ADD_380_U141, P3_ADD_380_U142, P3_ADD_380_U143, P3_ADD_380_U144, P3_ADD_380_U145, P3_ADD_380_U146, P3_ADD_380_U147, P3_ADD_380_U148, P3_ADD_380_U149, P3_ADD_380_U15, P3_ADD_380_U150, P3_ADD_380_U151, P3_ADD_380_U152, P3_ADD_380_U153, P3_ADD_380_U154, P3_ADD_380_U155, P3_ADD_380_U156, P3_ADD_380_U157, P3_ADD_380_U158, P3_ADD_380_U159, P3_ADD_380_U16, P3_ADD_380_U160, P3_ADD_380_U161, P3_ADD_380_U162, P3_ADD_380_U163, P3_ADD_380_U164, P3_ADD_380_U165, P3_ADD_380_U166, P3_ADD_380_U167, P3_ADD_380_U168, P3_ADD_380_U169, P3_ADD_380_U17, P3_ADD_380_U170, P3_ADD_380_U171, P3_ADD_380_U172, P3_ADD_380_U173, P3_ADD_380_U174, P3_ADD_380_U175, P3_ADD_380_U176, P3_ADD_380_U177, P3_ADD_380_U178, P3_ADD_380_U179, P3_ADD_380_U18, P3_ADD_380_U180, P3_ADD_380_U181, P3_ADD_380_U182, P3_ADD_380_U183, P3_ADD_380_U184, P3_ADD_380_U185, P3_ADD_380_U186, P3_ADD_380_U187, P3_ADD_380_U188, P3_ADD_380_U189, P3_ADD_380_U19, P3_ADD_380_U20, P3_ADD_380_U21, P3_ADD_380_U22, P3_ADD_380_U23, P3_ADD_380_U24, P3_ADD_380_U25, P3_ADD_380_U26, P3_ADD_380_U27, P3_ADD_380_U28, P3_ADD_380_U29, P3_ADD_380_U30, P3_ADD_380_U31, P3_ADD_380_U32, P3_ADD_380_U33, P3_ADD_380_U34, P3_ADD_380_U35, P3_ADD_380_U36, P3_ADD_380_U37, P3_ADD_380_U38, P3_ADD_380_U39, P3_ADD_380_U40, P3_ADD_380_U41, P3_ADD_380_U42, P3_ADD_380_U43, P3_ADD_380_U44, P3_ADD_380_U45, P3_ADD_380_U46, P3_ADD_380_U47, P3_ADD_380_U48, P3_ADD_380_U49, P3_ADD_380_U5, P3_ADD_380_U50, P3_ADD_380_U51, P3_ADD_380_U52, P3_ADD_380_U53, P3_ADD_380_U54, P3_ADD_380_U55, P3_ADD_380_U56, P3_ADD_380_U57, P3_ADD_380_U58, P3_ADD_380_U59, P3_ADD_380_U6, P3_ADD_380_U60, P3_ADD_380_U61, P3_ADD_380_U62, P3_ADD_380_U63, P3_ADD_380_U64, P3_ADD_380_U65, P3_ADD_380_U66, P3_ADD_380_U67, P3_ADD_380_U68, P3_ADD_380_U69, P3_ADD_380_U7, P3_ADD_380_U70, P3_ADD_380_U71, P3_ADD_380_U72, P3_ADD_380_U73, P3_ADD_380_U74, P3_ADD_380_U75, P3_ADD_380_U76, P3_ADD_380_U77, P3_ADD_380_U78, P3_ADD_380_U79, P3_ADD_380_U8, P3_ADD_380_U80, P3_ADD_380_U81, P3_ADD_380_U82, P3_ADD_380_U83, P3_ADD_380_U84, P3_ADD_380_U85, P3_ADD_380_U86, P3_ADD_380_U87, P3_ADD_380_U88, P3_ADD_380_U89, P3_ADD_380_U9, P3_ADD_380_U90, P3_ADD_380_U91, P3_ADD_380_U92, P3_ADD_380_U93, P3_ADD_380_U94, P3_ADD_380_U95, P3_ADD_380_U96, P3_ADD_380_U97, P3_ADD_380_U98, P3_ADD_380_U99, P3_ADD_385_U10, P3_ADD_385_U100, P3_ADD_385_U101, P3_ADD_385_U102, P3_ADD_385_U103, P3_ADD_385_U104, P3_ADD_385_U105, P3_ADD_385_U106, P3_ADD_385_U107, P3_ADD_385_U108, P3_ADD_385_U109, P3_ADD_385_U11, P3_ADD_385_U110, P3_ADD_385_U111, P3_ADD_385_U112, P3_ADD_385_U113, P3_ADD_385_U114, P3_ADD_385_U115, P3_ADD_385_U116, P3_ADD_385_U117, P3_ADD_385_U118, P3_ADD_385_U119, P3_ADD_385_U12, P3_ADD_385_U120, P3_ADD_385_U121, P3_ADD_385_U122, P3_ADD_385_U123, P3_ADD_385_U124, P3_ADD_385_U125, P3_ADD_385_U126, P3_ADD_385_U127, P3_ADD_385_U128, P3_ADD_385_U129, P3_ADD_385_U13, P3_ADD_385_U130, P3_ADD_385_U131, P3_ADD_385_U132, P3_ADD_385_U133, P3_ADD_385_U134, P3_ADD_385_U135, P3_ADD_385_U136, P3_ADD_385_U137, P3_ADD_385_U138, P3_ADD_385_U139, P3_ADD_385_U14, P3_ADD_385_U140, P3_ADD_385_U141, P3_ADD_385_U142, P3_ADD_385_U143, P3_ADD_385_U144, P3_ADD_385_U145, P3_ADD_385_U146, P3_ADD_385_U147, P3_ADD_385_U148, P3_ADD_385_U149, P3_ADD_385_U15, P3_ADD_385_U150, P3_ADD_385_U151, P3_ADD_385_U152, P3_ADD_385_U153, P3_ADD_385_U154, P3_ADD_385_U155, P3_ADD_385_U156, P3_ADD_385_U157, P3_ADD_385_U158, P3_ADD_385_U159, P3_ADD_385_U16, P3_ADD_385_U160, P3_ADD_385_U161, P3_ADD_385_U162, P3_ADD_385_U163, P3_ADD_385_U164, P3_ADD_385_U165, P3_ADD_385_U166, P3_ADD_385_U167, P3_ADD_385_U168, P3_ADD_385_U169, P3_ADD_385_U17, P3_ADD_385_U170, P3_ADD_385_U171, P3_ADD_385_U172, P3_ADD_385_U173, P3_ADD_385_U174, P3_ADD_385_U175, P3_ADD_385_U176, P3_ADD_385_U177, P3_ADD_385_U178, P3_ADD_385_U179, P3_ADD_385_U18, P3_ADD_385_U180, P3_ADD_385_U181, P3_ADD_385_U182, P3_ADD_385_U183, P3_ADD_385_U184, P3_ADD_385_U185, P3_ADD_385_U186, P3_ADD_385_U187, P3_ADD_385_U188, P3_ADD_385_U189, P3_ADD_385_U19, P3_ADD_385_U20, P3_ADD_385_U21, P3_ADD_385_U22, P3_ADD_385_U23, P3_ADD_385_U24, P3_ADD_385_U25, P3_ADD_385_U26, P3_ADD_385_U27, P3_ADD_385_U28, P3_ADD_385_U29, P3_ADD_385_U30, P3_ADD_385_U31, P3_ADD_385_U32, P3_ADD_385_U33, P3_ADD_385_U34, P3_ADD_385_U35, P3_ADD_385_U36, P3_ADD_385_U37, P3_ADD_385_U38, P3_ADD_385_U39, P3_ADD_385_U40, P3_ADD_385_U41, P3_ADD_385_U42, P3_ADD_385_U43, P3_ADD_385_U44, P3_ADD_385_U45, P3_ADD_385_U46, P3_ADD_385_U47, P3_ADD_385_U48, P3_ADD_385_U49, P3_ADD_385_U5, P3_ADD_385_U50, P3_ADD_385_U51, P3_ADD_385_U52, P3_ADD_385_U53, P3_ADD_385_U54, P3_ADD_385_U55, P3_ADD_385_U56, P3_ADD_385_U57, P3_ADD_385_U58, P3_ADD_385_U59, P3_ADD_385_U6, P3_ADD_385_U60, P3_ADD_385_U61, P3_ADD_385_U62, P3_ADD_385_U63, P3_ADD_385_U64, P3_ADD_385_U65, P3_ADD_385_U66, P3_ADD_385_U67, P3_ADD_385_U68, P3_ADD_385_U69, P3_ADD_385_U7, P3_ADD_385_U70, P3_ADD_385_U71, P3_ADD_385_U72, P3_ADD_385_U73, P3_ADD_385_U74, P3_ADD_385_U75, P3_ADD_385_U76, P3_ADD_385_U77, P3_ADD_385_U78, P3_ADD_385_U79, P3_ADD_385_U8, P3_ADD_385_U80, P3_ADD_385_U81, P3_ADD_385_U82, P3_ADD_385_U83, P3_ADD_385_U84, P3_ADD_385_U85, P3_ADD_385_U86, P3_ADD_385_U87, P3_ADD_385_U88, P3_ADD_385_U89, P3_ADD_385_U9, P3_ADD_385_U90, P3_ADD_385_U91, P3_ADD_385_U92, P3_ADD_385_U93, P3_ADD_385_U94, P3_ADD_385_U95, P3_ADD_385_U96, P3_ADD_385_U97, P3_ADD_385_U98, P3_ADD_385_U99, P3_ADD_391_1180_U10, P3_ADD_391_1180_U11, P3_ADD_391_1180_U12, P3_ADD_391_1180_U13, P3_ADD_391_1180_U14, P3_ADD_391_1180_U15, P3_ADD_391_1180_U16, P3_ADD_391_1180_U17, P3_ADD_391_1180_U18, P3_ADD_391_1180_U19, P3_ADD_391_1180_U20, P3_ADD_391_1180_U21, P3_ADD_391_1180_U22, P3_ADD_391_1180_U23, P3_ADD_391_1180_U24, P3_ADD_391_1180_U25, P3_ADD_391_1180_U26, P3_ADD_391_1180_U27, P3_ADD_391_1180_U28, P3_ADD_391_1180_U29, P3_ADD_391_1180_U30, P3_ADD_391_1180_U31, P3_ADD_391_1180_U32, P3_ADD_391_1180_U33, P3_ADD_391_1180_U34, P3_ADD_391_1180_U35, P3_ADD_391_1180_U36, P3_ADD_391_1180_U37, P3_ADD_391_1180_U38, P3_ADD_391_1180_U39, P3_ADD_391_1180_U4, P3_ADD_391_1180_U40, P3_ADD_391_1180_U41, P3_ADD_391_1180_U42, P3_ADD_391_1180_U43, P3_ADD_391_1180_U44, P3_ADD_391_1180_U45, P3_ADD_391_1180_U46, P3_ADD_391_1180_U47, P3_ADD_391_1180_U48, P3_ADD_391_1180_U49, P3_ADD_391_1180_U5, P3_ADD_391_1180_U50, P3_ADD_391_1180_U6, P3_ADD_391_1180_U7, P3_ADD_391_1180_U8, P3_ADD_391_1180_U9, P3_ADD_394_U10, P3_ADD_394_U100, P3_ADD_394_U101, P3_ADD_394_U102, P3_ADD_394_U103, P3_ADD_394_U104, P3_ADD_394_U105, P3_ADD_394_U106, P3_ADD_394_U107, P3_ADD_394_U108, P3_ADD_394_U109, P3_ADD_394_U11, P3_ADD_394_U110, P3_ADD_394_U111, P3_ADD_394_U112, P3_ADD_394_U113, P3_ADD_394_U114, P3_ADD_394_U115, P3_ADD_394_U116, P3_ADD_394_U117, P3_ADD_394_U118, P3_ADD_394_U119, P3_ADD_394_U12, P3_ADD_394_U120, P3_ADD_394_U121, P3_ADD_394_U122, P3_ADD_394_U123, P3_ADD_394_U124, P3_ADD_394_U125, P3_ADD_394_U126, P3_ADD_394_U127, P3_ADD_394_U128, P3_ADD_394_U129, P3_ADD_394_U13, P3_ADD_394_U130, P3_ADD_394_U131, P3_ADD_394_U132, P3_ADD_394_U133, P3_ADD_394_U134, P3_ADD_394_U135, P3_ADD_394_U136, P3_ADD_394_U137, P3_ADD_394_U138, P3_ADD_394_U139, P3_ADD_394_U14, P3_ADD_394_U140, P3_ADD_394_U141, P3_ADD_394_U142, P3_ADD_394_U143, P3_ADD_394_U144, P3_ADD_394_U145, P3_ADD_394_U146, P3_ADD_394_U147, P3_ADD_394_U148, P3_ADD_394_U149, P3_ADD_394_U15, P3_ADD_394_U150, P3_ADD_394_U151, P3_ADD_394_U152, P3_ADD_394_U153, P3_ADD_394_U154, P3_ADD_394_U155, P3_ADD_394_U156, P3_ADD_394_U157, P3_ADD_394_U158, P3_ADD_394_U159, P3_ADD_394_U16, P3_ADD_394_U160, P3_ADD_394_U161, P3_ADD_394_U162, P3_ADD_394_U163, P3_ADD_394_U164, P3_ADD_394_U165, P3_ADD_394_U166, P3_ADD_394_U167, P3_ADD_394_U168, P3_ADD_394_U169, P3_ADD_394_U17, P3_ADD_394_U170, P3_ADD_394_U171, P3_ADD_394_U172, P3_ADD_394_U173, P3_ADD_394_U174, P3_ADD_394_U175, P3_ADD_394_U176, P3_ADD_394_U177, P3_ADD_394_U178, P3_ADD_394_U179, P3_ADD_394_U18, P3_ADD_394_U180, P3_ADD_394_U181, P3_ADD_394_U182, P3_ADD_394_U183, P3_ADD_394_U184, P3_ADD_394_U185, P3_ADD_394_U186, P3_ADD_394_U19, P3_ADD_394_U20, P3_ADD_394_U21, P3_ADD_394_U22, P3_ADD_394_U23, P3_ADD_394_U24, P3_ADD_394_U25, P3_ADD_394_U26, P3_ADD_394_U27, P3_ADD_394_U28, P3_ADD_394_U29, P3_ADD_394_U30, P3_ADD_394_U31, P3_ADD_394_U32, P3_ADD_394_U33, P3_ADD_394_U34, P3_ADD_394_U35, P3_ADD_394_U36, P3_ADD_394_U37, P3_ADD_394_U38, P3_ADD_394_U39, P3_ADD_394_U4, P3_ADD_394_U40, P3_ADD_394_U41, P3_ADD_394_U42, P3_ADD_394_U43, P3_ADD_394_U44, P3_ADD_394_U45, P3_ADD_394_U46, P3_ADD_394_U47, P3_ADD_394_U48, P3_ADD_394_U49, P3_ADD_394_U5, P3_ADD_394_U50, P3_ADD_394_U51, P3_ADD_394_U52, P3_ADD_394_U53, P3_ADD_394_U54, P3_ADD_394_U55, P3_ADD_394_U56, P3_ADD_394_U57, P3_ADD_394_U58, P3_ADD_394_U59, P3_ADD_394_U6, P3_ADD_394_U60, P3_ADD_394_U61, P3_ADD_394_U62, P3_ADD_394_U63, P3_ADD_394_U64, P3_ADD_394_U65, P3_ADD_394_U66, P3_ADD_394_U67, P3_ADD_394_U68, P3_ADD_394_U69, P3_ADD_394_U7, P3_ADD_394_U70, P3_ADD_394_U71, P3_ADD_394_U72, P3_ADD_394_U73, P3_ADD_394_U74, P3_ADD_394_U75, P3_ADD_394_U76, P3_ADD_394_U77, P3_ADD_394_U78, P3_ADD_394_U79, P3_ADD_394_U8, P3_ADD_394_U80, P3_ADD_394_U81, P3_ADD_394_U82, P3_ADD_394_U83, P3_ADD_394_U84, P3_ADD_394_U85, P3_ADD_394_U86, P3_ADD_394_U87, P3_ADD_394_U88, P3_ADD_394_U89, P3_ADD_394_U9, P3_ADD_394_U90, P3_ADD_394_U91, P3_ADD_394_U92, P3_ADD_394_U93, P3_ADD_394_U94, P3_ADD_394_U95, P3_ADD_394_U96, P3_ADD_394_U97, P3_ADD_394_U98, P3_ADD_394_U99, P3_ADD_402_1132_U10, P3_ADD_402_1132_U11, P3_ADD_402_1132_U12, P3_ADD_402_1132_U13, P3_ADD_402_1132_U14, P3_ADD_402_1132_U15, P3_ADD_402_1132_U16, P3_ADD_402_1132_U17, P3_ADD_402_1132_U18, P3_ADD_402_1132_U19, P3_ADD_402_1132_U20, P3_ADD_402_1132_U21, P3_ADD_402_1132_U22, P3_ADD_402_1132_U23, P3_ADD_402_1132_U24, P3_ADD_402_1132_U25, P3_ADD_402_1132_U26, P3_ADD_402_1132_U27, P3_ADD_402_1132_U28, P3_ADD_402_1132_U29, P3_ADD_402_1132_U30, P3_ADD_402_1132_U31, P3_ADD_402_1132_U32, P3_ADD_402_1132_U33, P3_ADD_402_1132_U34, P3_ADD_402_1132_U35, P3_ADD_402_1132_U36, P3_ADD_402_1132_U37, P3_ADD_402_1132_U38, P3_ADD_402_1132_U39, P3_ADD_402_1132_U4, P3_ADD_402_1132_U40, P3_ADD_402_1132_U41, P3_ADD_402_1132_U42, P3_ADD_402_1132_U43, P3_ADD_402_1132_U44, P3_ADD_402_1132_U45, P3_ADD_402_1132_U46, P3_ADD_402_1132_U47, P3_ADD_402_1132_U48, P3_ADD_402_1132_U49, P3_ADD_402_1132_U5, P3_ADD_402_1132_U50, P3_ADD_402_1132_U6, P3_ADD_402_1132_U7, P3_ADD_402_1132_U8, P3_ADD_402_1132_U9, P3_ADD_405_U10, P3_ADD_405_U100, P3_ADD_405_U101, P3_ADD_405_U102, P3_ADD_405_U103, P3_ADD_405_U104, P3_ADD_405_U105, P3_ADD_405_U106, P3_ADD_405_U107, P3_ADD_405_U108, P3_ADD_405_U109, P3_ADD_405_U11, P3_ADD_405_U110, P3_ADD_405_U111, P3_ADD_405_U112, P3_ADD_405_U113, P3_ADD_405_U114, P3_ADD_405_U115, P3_ADD_405_U116, P3_ADD_405_U117, P3_ADD_405_U118, P3_ADD_405_U119, P3_ADD_405_U12, P3_ADD_405_U120, P3_ADD_405_U121, P3_ADD_405_U122, P3_ADD_405_U123, P3_ADD_405_U124, P3_ADD_405_U125, P3_ADD_405_U126, P3_ADD_405_U127, P3_ADD_405_U128, P3_ADD_405_U129, P3_ADD_405_U13, P3_ADD_405_U130, P3_ADD_405_U131, P3_ADD_405_U132, P3_ADD_405_U133, P3_ADD_405_U134, P3_ADD_405_U135, P3_ADD_405_U136, P3_ADD_405_U137, P3_ADD_405_U138, P3_ADD_405_U139, P3_ADD_405_U14, P3_ADD_405_U140, P3_ADD_405_U141, P3_ADD_405_U142, P3_ADD_405_U143, P3_ADD_405_U144, P3_ADD_405_U145, P3_ADD_405_U146, P3_ADD_405_U147, P3_ADD_405_U148, P3_ADD_405_U149, P3_ADD_405_U15, P3_ADD_405_U150, P3_ADD_405_U151, P3_ADD_405_U152, P3_ADD_405_U153, P3_ADD_405_U154, P3_ADD_405_U155, P3_ADD_405_U156, P3_ADD_405_U157, P3_ADD_405_U158, P3_ADD_405_U159, P3_ADD_405_U16, P3_ADD_405_U160, P3_ADD_405_U161, P3_ADD_405_U162, P3_ADD_405_U163, P3_ADD_405_U164, P3_ADD_405_U165, P3_ADD_405_U166, P3_ADD_405_U167, P3_ADD_405_U168, P3_ADD_405_U169, P3_ADD_405_U17, P3_ADD_405_U170, P3_ADD_405_U171, P3_ADD_405_U172, P3_ADD_405_U173, P3_ADD_405_U174, P3_ADD_405_U175, P3_ADD_405_U176, P3_ADD_405_U177, P3_ADD_405_U178, P3_ADD_405_U179, P3_ADD_405_U18, P3_ADD_405_U180, P3_ADD_405_U181, P3_ADD_405_U182, P3_ADD_405_U183, P3_ADD_405_U184, P3_ADD_405_U185, P3_ADD_405_U186, P3_ADD_405_U19, P3_ADD_405_U20, P3_ADD_405_U21, P3_ADD_405_U22, P3_ADD_405_U23, P3_ADD_405_U24, P3_ADD_405_U25, P3_ADD_405_U26, P3_ADD_405_U27, P3_ADD_405_U28, P3_ADD_405_U29, P3_ADD_405_U30, P3_ADD_405_U31, P3_ADD_405_U32, P3_ADD_405_U33, P3_ADD_405_U34, P3_ADD_405_U35, P3_ADD_405_U36, P3_ADD_405_U37, P3_ADD_405_U38, P3_ADD_405_U39, P3_ADD_405_U4, P3_ADD_405_U40, P3_ADD_405_U41, P3_ADD_405_U42, P3_ADD_405_U43, P3_ADD_405_U44, P3_ADD_405_U45, P3_ADD_405_U46, P3_ADD_405_U47, P3_ADD_405_U48, P3_ADD_405_U49, P3_ADD_405_U5, P3_ADD_405_U50, P3_ADD_405_U51, P3_ADD_405_U52, P3_ADD_405_U53, P3_ADD_405_U54, P3_ADD_405_U55, P3_ADD_405_U56, P3_ADD_405_U57, P3_ADD_405_U58, P3_ADD_405_U59, P3_ADD_405_U6, P3_ADD_405_U60, P3_ADD_405_U61, P3_ADD_405_U62, P3_ADD_405_U63, P3_ADD_405_U64, P3_ADD_405_U65, P3_ADD_405_U66, P3_ADD_405_U67, P3_ADD_405_U68, P3_ADD_405_U69, P3_ADD_405_U7, P3_ADD_405_U70, P3_ADD_405_U71, P3_ADD_405_U72, P3_ADD_405_U73, P3_ADD_405_U74, P3_ADD_405_U75, P3_ADD_405_U76, P3_ADD_405_U77, P3_ADD_405_U78, P3_ADD_405_U79, P3_ADD_405_U8, P3_ADD_405_U80, P3_ADD_405_U81, P3_ADD_405_U82, P3_ADD_405_U83, P3_ADD_405_U84, P3_ADD_405_U85, P3_ADD_405_U86, P3_ADD_405_U87, P3_ADD_405_U88, P3_ADD_405_U89, P3_ADD_405_U9, P3_ADD_405_U90, P3_ADD_405_U91, P3_ADD_405_U92, P3_ADD_405_U93, P3_ADD_405_U94, P3_ADD_405_U95, P3_ADD_405_U96, P3_ADD_405_U97, P3_ADD_405_U98, P3_ADD_405_U99, P3_ADD_430_U10, P3_ADD_430_U100, P3_ADD_430_U101, P3_ADD_430_U102, P3_ADD_430_U103, P3_ADD_430_U104, P3_ADD_430_U105, P3_ADD_430_U106, P3_ADD_430_U107, P3_ADD_430_U108, P3_ADD_430_U109, P3_ADD_430_U11, P3_ADD_430_U110, P3_ADD_430_U111, P3_ADD_430_U112, P3_ADD_430_U113, P3_ADD_430_U114, P3_ADD_430_U115, P3_ADD_430_U116, P3_ADD_430_U117, P3_ADD_430_U118, P3_ADD_430_U119, P3_ADD_430_U12, P3_ADD_430_U120, P3_ADD_430_U121, P3_ADD_430_U122, P3_ADD_430_U123, P3_ADD_430_U124, P3_ADD_430_U125, P3_ADD_430_U126, P3_ADD_430_U127, P3_ADD_430_U128, P3_ADD_430_U129, P3_ADD_430_U13, P3_ADD_430_U130, P3_ADD_430_U131, P3_ADD_430_U132, P3_ADD_430_U133, P3_ADD_430_U134, P3_ADD_430_U135, P3_ADD_430_U136, P3_ADD_430_U137, P3_ADD_430_U138, P3_ADD_430_U139, P3_ADD_430_U14, P3_ADD_430_U140, P3_ADD_430_U141, P3_ADD_430_U142, P3_ADD_430_U143, P3_ADD_430_U144, P3_ADD_430_U145, P3_ADD_430_U146, P3_ADD_430_U147, P3_ADD_430_U148, P3_ADD_430_U149, P3_ADD_430_U15, P3_ADD_430_U150, P3_ADD_430_U151, P3_ADD_430_U152, P3_ADD_430_U153, P3_ADD_430_U154, P3_ADD_430_U155, P3_ADD_430_U156, P3_ADD_430_U157, P3_ADD_430_U158, P3_ADD_430_U159, P3_ADD_430_U16, P3_ADD_430_U160, P3_ADD_430_U161, P3_ADD_430_U162, P3_ADD_430_U163, P3_ADD_430_U164, P3_ADD_430_U165, P3_ADD_430_U166, P3_ADD_430_U167, P3_ADD_430_U168, P3_ADD_430_U169, P3_ADD_430_U17, P3_ADD_430_U170, P3_ADD_430_U171, P3_ADD_430_U172, P3_ADD_430_U173, P3_ADD_430_U174, P3_ADD_430_U175, P3_ADD_430_U176, P3_ADD_430_U177, P3_ADD_430_U178, P3_ADD_430_U179, P3_ADD_430_U18, P3_ADD_430_U180, P3_ADD_430_U181, P3_ADD_430_U182, P3_ADD_430_U19, P3_ADD_430_U20, P3_ADD_430_U21, P3_ADD_430_U22, P3_ADD_430_U23, P3_ADD_430_U24, P3_ADD_430_U25, P3_ADD_430_U26, P3_ADD_430_U27, P3_ADD_430_U28, P3_ADD_430_U29, P3_ADD_430_U30, P3_ADD_430_U31, P3_ADD_430_U32, P3_ADD_430_U33, P3_ADD_430_U34, P3_ADD_430_U35, P3_ADD_430_U36, P3_ADD_430_U37, P3_ADD_430_U38, P3_ADD_430_U39, P3_ADD_430_U4, P3_ADD_430_U40, P3_ADD_430_U41, P3_ADD_430_U42, P3_ADD_430_U43, P3_ADD_430_U44, P3_ADD_430_U45, P3_ADD_430_U46, P3_ADD_430_U47, P3_ADD_430_U48, P3_ADD_430_U49, P3_ADD_430_U5, P3_ADD_430_U50, P3_ADD_430_U51, P3_ADD_430_U52, P3_ADD_430_U53, P3_ADD_430_U54, P3_ADD_430_U55, P3_ADD_430_U56, P3_ADD_430_U57, P3_ADD_430_U58, P3_ADD_430_U59, P3_ADD_430_U6, P3_ADD_430_U60, P3_ADD_430_U61, P3_ADD_430_U62, P3_ADD_430_U63, P3_ADD_430_U64, P3_ADD_430_U65, P3_ADD_430_U66, P3_ADD_430_U67, P3_ADD_430_U68, P3_ADD_430_U69, P3_ADD_430_U7, P3_ADD_430_U70, P3_ADD_430_U71, P3_ADD_430_U72, P3_ADD_430_U73, P3_ADD_430_U74, P3_ADD_430_U75, P3_ADD_430_U76, P3_ADD_430_U77, P3_ADD_430_U78, P3_ADD_430_U79, P3_ADD_430_U8, P3_ADD_430_U80, P3_ADD_430_U81, P3_ADD_430_U82, P3_ADD_430_U83, P3_ADD_430_U84, P3_ADD_430_U85, P3_ADD_430_U86, P3_ADD_430_U87, P3_ADD_430_U88, P3_ADD_430_U89, P3_ADD_430_U9, P3_ADD_430_U90, P3_ADD_430_U91, P3_ADD_430_U92, P3_ADD_430_U93, P3_ADD_430_U94, P3_ADD_430_U95, P3_ADD_430_U96, P3_ADD_430_U97, P3_ADD_430_U98, P3_ADD_430_U99, P3_ADD_441_U10, P3_ADD_441_U100, P3_ADD_441_U101, P3_ADD_441_U102, P3_ADD_441_U103, P3_ADD_441_U104, P3_ADD_441_U105, P3_ADD_441_U106, P3_ADD_441_U107, P3_ADD_441_U108, P3_ADD_441_U109, P3_ADD_441_U11, P3_ADD_441_U110, P3_ADD_441_U111, P3_ADD_441_U112, P3_ADD_441_U113, P3_ADD_441_U114, P3_ADD_441_U115, P3_ADD_441_U116, P3_ADD_441_U117, P3_ADD_441_U118, P3_ADD_441_U119, P3_ADD_441_U12, P3_ADD_441_U120, P3_ADD_441_U121, P3_ADD_441_U122, P3_ADD_441_U123, P3_ADD_441_U124, P3_ADD_441_U125, P3_ADD_441_U126, P3_ADD_441_U127, P3_ADD_441_U128, P3_ADD_441_U129, P3_ADD_441_U13, P3_ADD_441_U130, P3_ADD_441_U131, P3_ADD_441_U132, P3_ADD_441_U133, P3_ADD_441_U134, P3_ADD_441_U135, P3_ADD_441_U136, P3_ADD_441_U137, P3_ADD_441_U138, P3_ADD_441_U139, P3_ADD_441_U14, P3_ADD_441_U140, P3_ADD_441_U141, P3_ADD_441_U142, P3_ADD_441_U143, P3_ADD_441_U144, P3_ADD_441_U145, P3_ADD_441_U146, P3_ADD_441_U147, P3_ADD_441_U148, P3_ADD_441_U149, P3_ADD_441_U15, P3_ADD_441_U150, P3_ADD_441_U151, P3_ADD_441_U152, P3_ADD_441_U153, P3_ADD_441_U154, P3_ADD_441_U155, P3_ADD_441_U156, P3_ADD_441_U157, P3_ADD_441_U158, P3_ADD_441_U159, P3_ADD_441_U16, P3_ADD_441_U160, P3_ADD_441_U161, P3_ADD_441_U162, P3_ADD_441_U163, P3_ADD_441_U164, P3_ADD_441_U165, P3_ADD_441_U166, P3_ADD_441_U167, P3_ADD_441_U168, P3_ADD_441_U169, P3_ADD_441_U17, P3_ADD_441_U170, P3_ADD_441_U171, P3_ADD_441_U172, P3_ADD_441_U173, P3_ADD_441_U174, P3_ADD_441_U175, P3_ADD_441_U176, P3_ADD_441_U177, P3_ADD_441_U178, P3_ADD_441_U179, P3_ADD_441_U18, P3_ADD_441_U180, P3_ADD_441_U181, P3_ADD_441_U182, P3_ADD_441_U19, P3_ADD_441_U20, P3_ADD_441_U21, P3_ADD_441_U22, P3_ADD_441_U23, P3_ADD_441_U24, P3_ADD_441_U25, P3_ADD_441_U26, P3_ADD_441_U27, P3_ADD_441_U28, P3_ADD_441_U29, P3_ADD_441_U30, P3_ADD_441_U31, P3_ADD_441_U32, P3_ADD_441_U33, P3_ADD_441_U34, P3_ADD_441_U35, P3_ADD_441_U36, P3_ADD_441_U37, P3_ADD_441_U38, P3_ADD_441_U39, P3_ADD_441_U4, P3_ADD_441_U40, P3_ADD_441_U41, P3_ADD_441_U42, P3_ADD_441_U43, P3_ADD_441_U44, P3_ADD_441_U45, P3_ADD_441_U46, P3_ADD_441_U47, P3_ADD_441_U48, P3_ADD_441_U49, P3_ADD_441_U5, P3_ADD_441_U50, P3_ADD_441_U51, P3_ADD_441_U52, P3_ADD_441_U53, P3_ADD_441_U54, P3_ADD_441_U55, P3_ADD_441_U56, P3_ADD_441_U57, P3_ADD_441_U58, P3_ADD_441_U59, P3_ADD_441_U6, P3_ADD_441_U60, P3_ADD_441_U61, P3_ADD_441_U62, P3_ADD_441_U63, P3_ADD_441_U64, P3_ADD_441_U65, P3_ADD_441_U66, P3_ADD_441_U67, P3_ADD_441_U68, P3_ADD_441_U69, P3_ADD_441_U7, P3_ADD_441_U70, P3_ADD_441_U71, P3_ADD_441_U72, P3_ADD_441_U73, P3_ADD_441_U74, P3_ADD_441_U75, P3_ADD_441_U76, P3_ADD_441_U77, P3_ADD_441_U78, P3_ADD_441_U79, P3_ADD_441_U8, P3_ADD_441_U80, P3_ADD_441_U81, P3_ADD_441_U82, P3_ADD_441_U83, P3_ADD_441_U84, P3_ADD_441_U85, P3_ADD_441_U86, P3_ADD_441_U87, P3_ADD_441_U88, P3_ADD_441_U89, P3_ADD_441_U9, P3_ADD_441_U90, P3_ADD_441_U91, P3_ADD_441_U92, P3_ADD_441_U93, P3_ADD_441_U94, P3_ADD_441_U95, P3_ADD_441_U96, P3_ADD_441_U97, P3_ADD_441_U98, P3_ADD_441_U99, P3_ADD_467_U10, P3_ADD_467_U100, P3_ADD_467_U101, P3_ADD_467_U102, P3_ADD_467_U103, P3_ADD_467_U104, P3_ADD_467_U105, P3_ADD_467_U106, P3_ADD_467_U107, P3_ADD_467_U108, P3_ADD_467_U109, P3_ADD_467_U11, P3_ADD_467_U110, P3_ADD_467_U111, P3_ADD_467_U112, P3_ADD_467_U113, P3_ADD_467_U114, P3_ADD_467_U115, P3_ADD_467_U116, P3_ADD_467_U117, P3_ADD_467_U118, P3_ADD_467_U119, P3_ADD_467_U12, P3_ADD_467_U120, P3_ADD_467_U121, P3_ADD_467_U122, P3_ADD_467_U123, P3_ADD_467_U124, P3_ADD_467_U125, P3_ADD_467_U126, P3_ADD_467_U127, P3_ADD_467_U128, P3_ADD_467_U129, P3_ADD_467_U13, P3_ADD_467_U130, P3_ADD_467_U131, P3_ADD_467_U132, P3_ADD_467_U133, P3_ADD_467_U134, P3_ADD_467_U135, P3_ADD_467_U136, P3_ADD_467_U137, P3_ADD_467_U138, P3_ADD_467_U139, P3_ADD_467_U14, P3_ADD_467_U140, P3_ADD_467_U141, P3_ADD_467_U142, P3_ADD_467_U143, P3_ADD_467_U144, P3_ADD_467_U145, P3_ADD_467_U146, P3_ADD_467_U147, P3_ADD_467_U148, P3_ADD_467_U149, P3_ADD_467_U15, P3_ADD_467_U150, P3_ADD_467_U151, P3_ADD_467_U152, P3_ADD_467_U153, P3_ADD_467_U154, P3_ADD_467_U155, P3_ADD_467_U156, P3_ADD_467_U157, P3_ADD_467_U158, P3_ADD_467_U159, P3_ADD_467_U16, P3_ADD_467_U160, P3_ADD_467_U161, P3_ADD_467_U162, P3_ADD_467_U163, P3_ADD_467_U164, P3_ADD_467_U165, P3_ADD_467_U166, P3_ADD_467_U167, P3_ADD_467_U168, P3_ADD_467_U169, P3_ADD_467_U17, P3_ADD_467_U170, P3_ADD_467_U171, P3_ADD_467_U172, P3_ADD_467_U173, P3_ADD_467_U174, P3_ADD_467_U175, P3_ADD_467_U176, P3_ADD_467_U177, P3_ADD_467_U178, P3_ADD_467_U179, P3_ADD_467_U18, P3_ADD_467_U180, P3_ADD_467_U181, P3_ADD_467_U182, P3_ADD_467_U19, P3_ADD_467_U20, P3_ADD_467_U21, P3_ADD_467_U22, P3_ADD_467_U23, P3_ADD_467_U24, P3_ADD_467_U25, P3_ADD_467_U26, P3_ADD_467_U27, P3_ADD_467_U28, P3_ADD_467_U29, P3_ADD_467_U30, P3_ADD_467_U31, P3_ADD_467_U32, P3_ADD_467_U33, P3_ADD_467_U34, P3_ADD_467_U35, P3_ADD_467_U36, P3_ADD_467_U37, P3_ADD_467_U38, P3_ADD_467_U39, P3_ADD_467_U4, P3_ADD_467_U40, P3_ADD_467_U41, P3_ADD_467_U42, P3_ADD_467_U43, P3_ADD_467_U44, P3_ADD_467_U45, P3_ADD_467_U46, P3_ADD_467_U47, P3_ADD_467_U48, P3_ADD_467_U49, P3_ADD_467_U5, P3_ADD_467_U50, P3_ADD_467_U51, P3_ADD_467_U52, P3_ADD_467_U53, P3_ADD_467_U54, P3_ADD_467_U55, P3_ADD_467_U56, P3_ADD_467_U57, P3_ADD_467_U58, P3_ADD_467_U59, P3_ADD_467_U6, P3_ADD_467_U60, P3_ADD_467_U61, P3_ADD_467_U62, P3_ADD_467_U63, P3_ADD_467_U64, P3_ADD_467_U65, P3_ADD_467_U66, P3_ADD_467_U67, P3_ADD_467_U68, P3_ADD_467_U69, P3_ADD_467_U7, P3_ADD_467_U70, P3_ADD_467_U71, P3_ADD_467_U72, P3_ADD_467_U73, P3_ADD_467_U74, P3_ADD_467_U75, P3_ADD_467_U76, P3_ADD_467_U77, P3_ADD_467_U78, P3_ADD_467_U79, P3_ADD_467_U8, P3_ADD_467_U80, P3_ADD_467_U81, P3_ADD_467_U82, P3_ADD_467_U83, P3_ADD_467_U84, P3_ADD_467_U85, P3_ADD_467_U86, P3_ADD_467_U87, P3_ADD_467_U88, P3_ADD_467_U89, P3_ADD_467_U9, P3_ADD_467_U90, P3_ADD_467_U91, P3_ADD_467_U92, P3_ADD_467_U93, P3_ADD_467_U94, P3_ADD_467_U95, P3_ADD_467_U96, P3_ADD_467_U97, P3_ADD_467_U98, P3_ADD_467_U99, P3_ADD_476_U10, P3_ADD_476_U100, P3_ADD_476_U101, P3_ADD_476_U102, P3_ADD_476_U103, P3_ADD_476_U104, P3_ADD_476_U105, P3_ADD_476_U106, P3_ADD_476_U107, P3_ADD_476_U108, P3_ADD_476_U109, P3_ADD_476_U11, P3_ADD_476_U110, P3_ADD_476_U111, P3_ADD_476_U112, P3_ADD_476_U113, P3_ADD_476_U114, P3_ADD_476_U115, P3_ADD_476_U116, P3_ADD_476_U117, P3_ADD_476_U118, P3_ADD_476_U119, P3_ADD_476_U12, P3_ADD_476_U120, P3_ADD_476_U121, P3_ADD_476_U122, P3_ADD_476_U123, P3_ADD_476_U124, P3_ADD_476_U125, P3_ADD_476_U126, P3_ADD_476_U127, P3_ADD_476_U128, P3_ADD_476_U129, P3_ADD_476_U13, P3_ADD_476_U130, P3_ADD_476_U131, P3_ADD_476_U132, P3_ADD_476_U133, P3_ADD_476_U134, P3_ADD_476_U135, P3_ADD_476_U136, P3_ADD_476_U137, P3_ADD_476_U138, P3_ADD_476_U139, P3_ADD_476_U14, P3_ADD_476_U140, P3_ADD_476_U141, P3_ADD_476_U142, P3_ADD_476_U143, P3_ADD_476_U144, P3_ADD_476_U145, P3_ADD_476_U146, P3_ADD_476_U147, P3_ADD_476_U148, P3_ADD_476_U149, P3_ADD_476_U15, P3_ADD_476_U150, P3_ADD_476_U151, P3_ADD_476_U152, P3_ADD_476_U153, P3_ADD_476_U154, P3_ADD_476_U155, P3_ADD_476_U156, P3_ADD_476_U157, P3_ADD_476_U158, P3_ADD_476_U159, P3_ADD_476_U16, P3_ADD_476_U160, P3_ADD_476_U161, P3_ADD_476_U162, P3_ADD_476_U163, P3_ADD_476_U164, P3_ADD_476_U165, P3_ADD_476_U166, P3_ADD_476_U167, P3_ADD_476_U168, P3_ADD_476_U169, P3_ADD_476_U17, P3_ADD_476_U170, P3_ADD_476_U171, P3_ADD_476_U172, P3_ADD_476_U173, P3_ADD_476_U174, P3_ADD_476_U175, P3_ADD_476_U176, P3_ADD_476_U177, P3_ADD_476_U178, P3_ADD_476_U179, P3_ADD_476_U18, P3_ADD_476_U180, P3_ADD_476_U181, P3_ADD_476_U182, P3_ADD_476_U19, P3_ADD_476_U20, P3_ADD_476_U21, P3_ADD_476_U22, P3_ADD_476_U23, P3_ADD_476_U24, P3_ADD_476_U25, P3_ADD_476_U26, P3_ADD_476_U27, P3_ADD_476_U28, P3_ADD_476_U29, P3_ADD_476_U30, P3_ADD_476_U31, P3_ADD_476_U32, P3_ADD_476_U33, P3_ADD_476_U34, P3_ADD_476_U35, P3_ADD_476_U36, P3_ADD_476_U37, P3_ADD_476_U38, P3_ADD_476_U39, P3_ADD_476_U4, P3_ADD_476_U40, P3_ADD_476_U41, P3_ADD_476_U42, P3_ADD_476_U43, P3_ADD_476_U44, P3_ADD_476_U45, P3_ADD_476_U46, P3_ADD_476_U47, P3_ADD_476_U48, P3_ADD_476_U49, P3_ADD_476_U5, P3_ADD_476_U50, P3_ADD_476_U51, P3_ADD_476_U52, P3_ADD_476_U53, P3_ADD_476_U54, P3_ADD_476_U55, P3_ADD_476_U56, P3_ADD_476_U57, P3_ADD_476_U58, P3_ADD_476_U59, P3_ADD_476_U6, P3_ADD_476_U60, P3_ADD_476_U61, P3_ADD_476_U62, P3_ADD_476_U63, P3_ADD_476_U64, P3_ADD_476_U65, P3_ADD_476_U66, P3_ADD_476_U67, P3_ADD_476_U68, P3_ADD_476_U69, P3_ADD_476_U7, P3_ADD_476_U70, P3_ADD_476_U71, P3_ADD_476_U72, P3_ADD_476_U73, P3_ADD_476_U74, P3_ADD_476_U75, P3_ADD_476_U76, P3_ADD_476_U77, P3_ADD_476_U78, P3_ADD_476_U79, P3_ADD_476_U8, P3_ADD_476_U80, P3_ADD_476_U81, P3_ADD_476_U82, P3_ADD_476_U83, P3_ADD_476_U84, P3_ADD_476_U85, P3_ADD_476_U86, P3_ADD_476_U87, P3_ADD_476_U88, P3_ADD_476_U89, P3_ADD_476_U9, P3_ADD_476_U90, P3_ADD_476_U91, P3_ADD_476_U92, P3_ADD_476_U93, P3_ADD_476_U94, P3_ADD_476_U95, P3_ADD_476_U96, P3_ADD_476_U97, P3_ADD_476_U98, P3_ADD_476_U99, P3_ADD_486_U10, P3_ADD_486_U11, P3_ADD_486_U12, P3_ADD_486_U13, P3_ADD_486_U14, P3_ADD_486_U15, P3_ADD_486_U16, P3_ADD_486_U17, P3_ADD_486_U18, P3_ADD_486_U19, P3_ADD_486_U20, P3_ADD_486_U21, P3_ADD_486_U22, P3_ADD_486_U23, P3_ADD_486_U24, P3_ADD_486_U25, P3_ADD_486_U26, P3_ADD_486_U27, P3_ADD_486_U28, P3_ADD_486_U5, P3_ADD_486_U6, P3_ADD_486_U7, P3_ADD_486_U8, P3_ADD_486_U9, P3_ADD_494_U10, P3_ADD_494_U100, P3_ADD_494_U101, P3_ADD_494_U102, P3_ADD_494_U103, P3_ADD_494_U104, P3_ADD_494_U105, P3_ADD_494_U106, P3_ADD_494_U107, P3_ADD_494_U108, P3_ADD_494_U109, P3_ADD_494_U11, P3_ADD_494_U110, P3_ADD_494_U111, P3_ADD_494_U112, P3_ADD_494_U113, P3_ADD_494_U114, P3_ADD_494_U115, P3_ADD_494_U116, P3_ADD_494_U117, P3_ADD_494_U118, P3_ADD_494_U119, P3_ADD_494_U12, P3_ADD_494_U120, P3_ADD_494_U121, P3_ADD_494_U122, P3_ADD_494_U123, P3_ADD_494_U124, P3_ADD_494_U125, P3_ADD_494_U126, P3_ADD_494_U127, P3_ADD_494_U128, P3_ADD_494_U129, P3_ADD_494_U13, P3_ADD_494_U130, P3_ADD_494_U131, P3_ADD_494_U132, P3_ADD_494_U133, P3_ADD_494_U134, P3_ADD_494_U135, P3_ADD_494_U136, P3_ADD_494_U137, P3_ADD_494_U138, P3_ADD_494_U139, P3_ADD_494_U14, P3_ADD_494_U140, P3_ADD_494_U141, P3_ADD_494_U142, P3_ADD_494_U143, P3_ADD_494_U144, P3_ADD_494_U145, P3_ADD_494_U146, P3_ADD_494_U147, P3_ADD_494_U148, P3_ADD_494_U149, P3_ADD_494_U15, P3_ADD_494_U150, P3_ADD_494_U151, P3_ADD_494_U152, P3_ADD_494_U153, P3_ADD_494_U154, P3_ADD_494_U155, P3_ADD_494_U156, P3_ADD_494_U157, P3_ADD_494_U158, P3_ADD_494_U159, P3_ADD_494_U16, P3_ADD_494_U160, P3_ADD_494_U161, P3_ADD_494_U162, P3_ADD_494_U163, P3_ADD_494_U164, P3_ADD_494_U165, P3_ADD_494_U166, P3_ADD_494_U167, P3_ADD_494_U168, P3_ADD_494_U169, P3_ADD_494_U17, P3_ADD_494_U170, P3_ADD_494_U171, P3_ADD_494_U172, P3_ADD_494_U173, P3_ADD_494_U174, P3_ADD_494_U175, P3_ADD_494_U176, P3_ADD_494_U177, P3_ADD_494_U178, P3_ADD_494_U179, P3_ADD_494_U18, P3_ADD_494_U180, P3_ADD_494_U181, P3_ADD_494_U182, P3_ADD_494_U19, P3_ADD_494_U20, P3_ADD_494_U21, P3_ADD_494_U22, P3_ADD_494_U23, P3_ADD_494_U24, P3_ADD_494_U25, P3_ADD_494_U26, P3_ADD_494_U27, P3_ADD_494_U28, P3_ADD_494_U29, P3_ADD_494_U30, P3_ADD_494_U31, P3_ADD_494_U32, P3_ADD_494_U33, P3_ADD_494_U34, P3_ADD_494_U35, P3_ADD_494_U36, P3_ADD_494_U37, P3_ADD_494_U38, P3_ADD_494_U39, P3_ADD_494_U4, P3_ADD_494_U40, P3_ADD_494_U41, P3_ADD_494_U42, P3_ADD_494_U43, P3_ADD_494_U44, P3_ADD_494_U45, P3_ADD_494_U46, P3_ADD_494_U47, P3_ADD_494_U48, P3_ADD_494_U49, P3_ADD_494_U5, P3_ADD_494_U50, P3_ADD_494_U51, P3_ADD_494_U52, P3_ADD_494_U53, P3_ADD_494_U54, P3_ADD_494_U55, P3_ADD_494_U56, P3_ADD_494_U57, P3_ADD_494_U58, P3_ADD_494_U59, P3_ADD_494_U6, P3_ADD_494_U60, P3_ADD_494_U61, P3_ADD_494_U62, P3_ADD_494_U63, P3_ADD_494_U64, P3_ADD_494_U65, P3_ADD_494_U66, P3_ADD_494_U67, P3_ADD_494_U68, P3_ADD_494_U69, P3_ADD_494_U7, P3_ADD_494_U70, P3_ADD_494_U71, P3_ADD_494_U72, P3_ADD_494_U73, P3_ADD_494_U74, P3_ADD_494_U75, P3_ADD_494_U76, P3_ADD_494_U77, P3_ADD_494_U78, P3_ADD_494_U79, P3_ADD_494_U8, P3_ADD_494_U80, P3_ADD_494_U81, P3_ADD_494_U82, P3_ADD_494_U83, P3_ADD_494_U84, P3_ADD_494_U85, P3_ADD_494_U86, P3_ADD_494_U87, P3_ADD_494_U88, P3_ADD_494_U89, P3_ADD_494_U9, P3_ADD_494_U90, P3_ADD_494_U91, P3_ADD_494_U92, P3_ADD_494_U93, P3_ADD_494_U94, P3_ADD_494_U95, P3_ADD_494_U96, P3_ADD_494_U97, P3_ADD_494_U98, P3_ADD_494_U99, P3_ADD_495_U10, P3_ADD_495_U11, P3_ADD_495_U12, P3_ADD_495_U13, P3_ADD_495_U14, P3_ADD_495_U15, P3_ADD_495_U16, P3_ADD_495_U17, P3_ADD_495_U18, P3_ADD_495_U19, P3_ADD_495_U20, P3_ADD_495_U4, P3_ADD_495_U5, P3_ADD_495_U6, P3_ADD_495_U7, P3_ADD_495_U8, P3_ADD_495_U9, P3_ADD_505_U10, P3_ADD_505_U11, P3_ADD_505_U12, P3_ADD_505_U13, P3_ADD_505_U14, P3_ADD_505_U15, P3_ADD_505_U16, P3_ADD_505_U17, P3_ADD_505_U18, P3_ADD_505_U19, P3_ADD_505_U20, P3_ADD_505_U21, P3_ADD_505_U22, P3_ADD_505_U23, P3_ADD_505_U24, P3_ADD_505_U25, P3_ADD_505_U26, P3_ADD_505_U27, P3_ADD_505_U28, P3_ADD_505_U5, P3_ADD_505_U6, P3_ADD_505_U7, P3_ADD_505_U8, P3_ADD_505_U9, P3_ADD_515_U10, P3_ADD_515_U100, P3_ADD_515_U101, P3_ADD_515_U102, P3_ADD_515_U103, P3_ADD_515_U104, P3_ADD_515_U105, P3_ADD_515_U106, P3_ADD_515_U107, P3_ADD_515_U108, P3_ADD_515_U109, P3_ADD_515_U11, P3_ADD_515_U110, P3_ADD_515_U111, P3_ADD_515_U112, P3_ADD_515_U113, P3_ADD_515_U114, P3_ADD_515_U115, P3_ADD_515_U116, P3_ADD_515_U117, P3_ADD_515_U118, P3_ADD_515_U119, P3_ADD_515_U12, P3_ADD_515_U120, P3_ADD_515_U121, P3_ADD_515_U122, P3_ADD_515_U123, P3_ADD_515_U124, P3_ADD_515_U125, P3_ADD_515_U126, P3_ADD_515_U127, P3_ADD_515_U128, P3_ADD_515_U129, P3_ADD_515_U13, P3_ADD_515_U130, P3_ADD_515_U131, P3_ADD_515_U132, P3_ADD_515_U133, P3_ADD_515_U134, P3_ADD_515_U135, P3_ADD_515_U136, P3_ADD_515_U137, P3_ADD_515_U138, P3_ADD_515_U139, P3_ADD_515_U14, P3_ADD_515_U140, P3_ADD_515_U141, P3_ADD_515_U142, P3_ADD_515_U143, P3_ADD_515_U144, P3_ADD_515_U145, P3_ADD_515_U146, P3_ADD_515_U147, P3_ADD_515_U148, P3_ADD_515_U149, P3_ADD_515_U15, P3_ADD_515_U150, P3_ADD_515_U151, P3_ADD_515_U152, P3_ADD_515_U153, P3_ADD_515_U154, P3_ADD_515_U155, P3_ADD_515_U156, P3_ADD_515_U157, P3_ADD_515_U158, P3_ADD_515_U159, P3_ADD_515_U16, P3_ADD_515_U160, P3_ADD_515_U161, P3_ADD_515_U162, P3_ADD_515_U163, P3_ADD_515_U164, P3_ADD_515_U165, P3_ADD_515_U166, P3_ADD_515_U167, P3_ADD_515_U168, P3_ADD_515_U169, P3_ADD_515_U17, P3_ADD_515_U170, P3_ADD_515_U171, P3_ADD_515_U172, P3_ADD_515_U173, P3_ADD_515_U174, P3_ADD_515_U175, P3_ADD_515_U176, P3_ADD_515_U177, P3_ADD_515_U178, P3_ADD_515_U179, P3_ADD_515_U18, P3_ADD_515_U180, P3_ADD_515_U181, P3_ADD_515_U182, P3_ADD_515_U19, P3_ADD_515_U20, P3_ADD_515_U21, P3_ADD_515_U22, P3_ADD_515_U23, P3_ADD_515_U24, P3_ADD_515_U25, P3_ADD_515_U26, P3_ADD_515_U27, P3_ADD_515_U28, P3_ADD_515_U29, P3_ADD_515_U30, P3_ADD_515_U31, P3_ADD_515_U32, P3_ADD_515_U33, P3_ADD_515_U34, P3_ADD_515_U35, P3_ADD_515_U36, P3_ADD_515_U37, P3_ADD_515_U38, P3_ADD_515_U39, P3_ADD_515_U4, P3_ADD_515_U40, P3_ADD_515_U41, P3_ADD_515_U42, P3_ADD_515_U43, P3_ADD_515_U44, P3_ADD_515_U45, P3_ADD_515_U46, P3_ADD_515_U47, P3_ADD_515_U48, P3_ADD_515_U49, P3_ADD_515_U5, P3_ADD_515_U50, P3_ADD_515_U51, P3_ADD_515_U52, P3_ADD_515_U53, P3_ADD_515_U54, P3_ADD_515_U55, P3_ADD_515_U56, P3_ADD_515_U57, P3_ADD_515_U58, P3_ADD_515_U59, P3_ADD_515_U6, P3_ADD_515_U60, P3_ADD_515_U61, P3_ADD_515_U62, P3_ADD_515_U63, P3_ADD_515_U64, P3_ADD_515_U65, P3_ADD_515_U66, P3_ADD_515_U67, P3_ADD_515_U68, P3_ADD_515_U69, P3_ADD_515_U7, P3_ADD_515_U70, P3_ADD_515_U71, P3_ADD_515_U72, P3_ADD_515_U73, P3_ADD_515_U74, P3_ADD_515_U75, P3_ADD_515_U76, P3_ADD_515_U77, P3_ADD_515_U78, P3_ADD_515_U79, P3_ADD_515_U8, P3_ADD_515_U80, P3_ADD_515_U81, P3_ADD_515_U82, P3_ADD_515_U83, P3_ADD_515_U84, P3_ADD_515_U85, P3_ADD_515_U86, P3_ADD_515_U87, P3_ADD_515_U88, P3_ADD_515_U89, P3_ADD_515_U9, P3_ADD_515_U90, P3_ADD_515_U91, P3_ADD_515_U92, P3_ADD_515_U93, P3_ADD_515_U94, P3_ADD_515_U95, P3_ADD_515_U96, P3_ADD_515_U97, P3_ADD_515_U98, P3_ADD_515_U99, P3_ADD_526_U10, P3_ADD_526_U100, P3_ADD_526_U101, P3_ADD_526_U102, P3_ADD_526_U103, P3_ADD_526_U104, P3_ADD_526_U105, P3_ADD_526_U106, P3_ADD_526_U107, P3_ADD_526_U108, P3_ADD_526_U109, P3_ADD_526_U11, P3_ADD_526_U110, P3_ADD_526_U111, P3_ADD_526_U112, P3_ADD_526_U113, P3_ADD_526_U114, P3_ADD_526_U115, P3_ADD_526_U116, P3_ADD_526_U117, P3_ADD_526_U118, P3_ADD_526_U119, P3_ADD_526_U12, P3_ADD_526_U120, P3_ADD_526_U121, P3_ADD_526_U122, P3_ADD_526_U123, P3_ADD_526_U124, P3_ADD_526_U125, P3_ADD_526_U126, P3_ADD_526_U127, P3_ADD_526_U128, P3_ADD_526_U129, P3_ADD_526_U13, P3_ADD_526_U130, P3_ADD_526_U131, P3_ADD_526_U132, P3_ADD_526_U133, P3_ADD_526_U134, P3_ADD_526_U135, P3_ADD_526_U136, P3_ADD_526_U137, P3_ADD_526_U138, P3_ADD_526_U139, P3_ADD_526_U14, P3_ADD_526_U140, P3_ADD_526_U141, P3_ADD_526_U142, P3_ADD_526_U143, P3_ADD_526_U144, P3_ADD_526_U145, P3_ADD_526_U146, P3_ADD_526_U147, P3_ADD_526_U148, P3_ADD_526_U149, P3_ADD_526_U15, P3_ADD_526_U150, P3_ADD_526_U151, P3_ADD_526_U152, P3_ADD_526_U153, P3_ADD_526_U154, P3_ADD_526_U155, P3_ADD_526_U156, P3_ADD_526_U157, P3_ADD_526_U158, P3_ADD_526_U159, P3_ADD_526_U16, P3_ADD_526_U160, P3_ADD_526_U161, P3_ADD_526_U162, P3_ADD_526_U163, P3_ADD_526_U164, P3_ADD_526_U165, P3_ADD_526_U166, P3_ADD_526_U167, P3_ADD_526_U168, P3_ADD_526_U169, P3_ADD_526_U17, P3_ADD_526_U170, P3_ADD_526_U171, P3_ADD_526_U172, P3_ADD_526_U173, P3_ADD_526_U174, P3_ADD_526_U175, P3_ADD_526_U176, P3_ADD_526_U177, P3_ADD_526_U178, P3_ADD_526_U179, P3_ADD_526_U18, P3_ADD_526_U180, P3_ADD_526_U181, P3_ADD_526_U182, P3_ADD_526_U183, P3_ADD_526_U184, P3_ADD_526_U185, P3_ADD_526_U186, P3_ADD_526_U187, P3_ADD_526_U188, P3_ADD_526_U189, P3_ADD_526_U19, P3_ADD_526_U190, P3_ADD_526_U191, P3_ADD_526_U192, P3_ADD_526_U193, P3_ADD_526_U194, P3_ADD_526_U195, P3_ADD_526_U196, P3_ADD_526_U197, P3_ADD_526_U198, P3_ADD_526_U199, P3_ADD_526_U20, P3_ADD_526_U200, P3_ADD_526_U201, P3_ADD_526_U202, P3_ADD_526_U21, P3_ADD_526_U22, P3_ADD_526_U23, P3_ADD_526_U24, P3_ADD_526_U25, P3_ADD_526_U26, P3_ADD_526_U27, P3_ADD_526_U28, P3_ADD_526_U29, P3_ADD_526_U30, P3_ADD_526_U31, P3_ADD_526_U32, P3_ADD_526_U33, P3_ADD_526_U34, P3_ADD_526_U35, P3_ADD_526_U36, P3_ADD_526_U37, P3_ADD_526_U38, P3_ADD_526_U39, P3_ADD_526_U40, P3_ADD_526_U41, P3_ADD_526_U42, P3_ADD_526_U43, P3_ADD_526_U44, P3_ADD_526_U45, P3_ADD_526_U46, P3_ADD_526_U47, P3_ADD_526_U48, P3_ADD_526_U49, P3_ADD_526_U5, P3_ADD_526_U50, P3_ADD_526_U51, P3_ADD_526_U52, P3_ADD_526_U53, P3_ADD_526_U54, P3_ADD_526_U55, P3_ADD_526_U56, P3_ADD_526_U57, P3_ADD_526_U58, P3_ADD_526_U59, P3_ADD_526_U6, P3_ADD_526_U60, P3_ADD_526_U61, P3_ADD_526_U62, P3_ADD_526_U63, P3_ADD_526_U64, P3_ADD_526_U65, P3_ADD_526_U66, P3_ADD_526_U67, P3_ADD_526_U68, P3_ADD_526_U69, P3_ADD_526_U7, P3_ADD_526_U70, P3_ADD_526_U71, P3_ADD_526_U72, P3_ADD_526_U73, P3_ADD_526_U74, P3_ADD_526_U75, P3_ADD_526_U76, P3_ADD_526_U77, P3_ADD_526_U78, P3_ADD_526_U79, P3_ADD_526_U8, P3_ADD_526_U80, P3_ADD_526_U81, P3_ADD_526_U82, P3_ADD_526_U83, P3_ADD_526_U84, P3_ADD_526_U85, P3_ADD_526_U86, P3_ADD_526_U87, P3_ADD_526_U88, P3_ADD_526_U89, P3_ADD_526_U9, P3_ADD_526_U90, P3_ADD_526_U91, P3_ADD_526_U92, P3_ADD_526_U93, P3_ADD_526_U94, P3_ADD_526_U95, P3_ADD_526_U96, P3_ADD_526_U97, P3_ADD_526_U98, P3_ADD_526_U99, P3_ADD_531_U10, P3_ADD_531_U100, P3_ADD_531_U101, P3_ADD_531_U102, P3_ADD_531_U103, P3_ADD_531_U104, P3_ADD_531_U105, P3_ADD_531_U106, P3_ADD_531_U107, P3_ADD_531_U108, P3_ADD_531_U109, P3_ADD_531_U11, P3_ADD_531_U110, P3_ADD_531_U111, P3_ADD_531_U112, P3_ADD_531_U113, P3_ADD_531_U114, P3_ADD_531_U115, P3_ADD_531_U116, P3_ADD_531_U117, P3_ADD_531_U118, P3_ADD_531_U119, P3_ADD_531_U12, P3_ADD_531_U120, P3_ADD_531_U121, P3_ADD_531_U122, P3_ADD_531_U123, P3_ADD_531_U124, P3_ADD_531_U125, P3_ADD_531_U126, P3_ADD_531_U127, P3_ADD_531_U128, P3_ADD_531_U129, P3_ADD_531_U13, P3_ADD_531_U130, P3_ADD_531_U131, P3_ADD_531_U132, P3_ADD_531_U133, P3_ADD_531_U134, P3_ADD_531_U135, P3_ADD_531_U136, P3_ADD_531_U137, P3_ADD_531_U138, P3_ADD_531_U139, P3_ADD_531_U14, P3_ADD_531_U140, P3_ADD_531_U141, P3_ADD_531_U142, P3_ADD_531_U143, P3_ADD_531_U144, P3_ADD_531_U145, P3_ADD_531_U146, P3_ADD_531_U147, P3_ADD_531_U148, P3_ADD_531_U149, P3_ADD_531_U15, P3_ADD_531_U150, P3_ADD_531_U151, P3_ADD_531_U152, P3_ADD_531_U153, P3_ADD_531_U154, P3_ADD_531_U155, P3_ADD_531_U156, P3_ADD_531_U157, P3_ADD_531_U158, P3_ADD_531_U159, P3_ADD_531_U16, P3_ADD_531_U160, P3_ADD_531_U161, P3_ADD_531_U162, P3_ADD_531_U163, P3_ADD_531_U164, P3_ADD_531_U165, P3_ADD_531_U166, P3_ADD_531_U167, P3_ADD_531_U168, P3_ADD_531_U169, P3_ADD_531_U17, P3_ADD_531_U170, P3_ADD_531_U171, P3_ADD_531_U172, P3_ADD_531_U173, P3_ADD_531_U174, P3_ADD_531_U175, P3_ADD_531_U176, P3_ADD_531_U177, P3_ADD_531_U178, P3_ADD_531_U179, P3_ADD_531_U18, P3_ADD_531_U180, P3_ADD_531_U181, P3_ADD_531_U182, P3_ADD_531_U183, P3_ADD_531_U184, P3_ADD_531_U185, P3_ADD_531_U186, P3_ADD_531_U187, P3_ADD_531_U188, P3_ADD_531_U189, P3_ADD_531_U19, P3_ADD_531_U20, P3_ADD_531_U21, P3_ADD_531_U22, P3_ADD_531_U23, P3_ADD_531_U24, P3_ADD_531_U25, P3_ADD_531_U26, P3_ADD_531_U27, P3_ADD_531_U28, P3_ADD_531_U29, P3_ADD_531_U30, P3_ADD_531_U31, P3_ADD_531_U32, P3_ADD_531_U33, P3_ADD_531_U34, P3_ADD_531_U35, P3_ADD_531_U36, P3_ADD_531_U37, P3_ADD_531_U38, P3_ADD_531_U39, P3_ADD_531_U40, P3_ADD_531_U41, P3_ADD_531_U42, P3_ADD_531_U43, P3_ADD_531_U44, P3_ADD_531_U45, P3_ADD_531_U46, P3_ADD_531_U47, P3_ADD_531_U48, P3_ADD_531_U49, P3_ADD_531_U5, P3_ADD_531_U50, P3_ADD_531_U51, P3_ADD_531_U52, P3_ADD_531_U53, P3_ADD_531_U54, P3_ADD_531_U55, P3_ADD_531_U56, P3_ADD_531_U57, P3_ADD_531_U58, P3_ADD_531_U59, P3_ADD_531_U6, P3_ADD_531_U60, P3_ADD_531_U61, P3_ADD_531_U62, P3_ADD_531_U63, P3_ADD_531_U64, P3_ADD_531_U65, P3_ADD_531_U66, P3_ADD_531_U67, P3_ADD_531_U68, P3_ADD_531_U69, P3_ADD_531_U7, P3_ADD_531_U70, P3_ADD_531_U71, P3_ADD_531_U72, P3_ADD_531_U73, P3_ADD_531_U74, P3_ADD_531_U75, P3_ADD_531_U76, P3_ADD_531_U77, P3_ADD_531_U78, P3_ADD_531_U79, P3_ADD_531_U8, P3_ADD_531_U80, P3_ADD_531_U81, P3_ADD_531_U82, P3_ADD_531_U83, P3_ADD_531_U84, P3_ADD_531_U85, P3_ADD_531_U86, P3_ADD_531_U87, P3_ADD_531_U88, P3_ADD_531_U89, P3_ADD_531_U9, P3_ADD_531_U90, P3_ADD_531_U91, P3_ADD_531_U92, P3_ADD_531_U93, P3_ADD_531_U94, P3_ADD_531_U95, P3_ADD_531_U96, P3_ADD_531_U97, P3_ADD_531_U98, P3_ADD_531_U99, P3_ADD_536_U10, P3_ADD_536_U100, P3_ADD_536_U101, P3_ADD_536_U102, P3_ADD_536_U103, P3_ADD_536_U104, P3_ADD_536_U105, P3_ADD_536_U106, P3_ADD_536_U107, P3_ADD_536_U108, P3_ADD_536_U109, P3_ADD_536_U11, P3_ADD_536_U110, P3_ADD_536_U111, P3_ADD_536_U112, P3_ADD_536_U113, P3_ADD_536_U114, P3_ADD_536_U115, P3_ADD_536_U116, P3_ADD_536_U117, P3_ADD_536_U118, P3_ADD_536_U119, P3_ADD_536_U12, P3_ADD_536_U120, P3_ADD_536_U121, P3_ADD_536_U122, P3_ADD_536_U123, P3_ADD_536_U124, P3_ADD_536_U125, P3_ADD_536_U126, P3_ADD_536_U127, P3_ADD_536_U128, P3_ADD_536_U129, P3_ADD_536_U13, P3_ADD_536_U130, P3_ADD_536_U131, P3_ADD_536_U132, P3_ADD_536_U133, P3_ADD_536_U134, P3_ADD_536_U135, P3_ADD_536_U136, P3_ADD_536_U137, P3_ADD_536_U138, P3_ADD_536_U139, P3_ADD_536_U14, P3_ADD_536_U140, P3_ADD_536_U141, P3_ADD_536_U142, P3_ADD_536_U143, P3_ADD_536_U144, P3_ADD_536_U145, P3_ADD_536_U146, P3_ADD_536_U147, P3_ADD_536_U148, P3_ADD_536_U149, P3_ADD_536_U15, P3_ADD_536_U150, P3_ADD_536_U151, P3_ADD_536_U152, P3_ADD_536_U153, P3_ADD_536_U154, P3_ADD_536_U155, P3_ADD_536_U156, P3_ADD_536_U157, P3_ADD_536_U158, P3_ADD_536_U159, P3_ADD_536_U16, P3_ADD_536_U160, P3_ADD_536_U161, P3_ADD_536_U162, P3_ADD_536_U163, P3_ADD_536_U164, P3_ADD_536_U165, P3_ADD_536_U166, P3_ADD_536_U167, P3_ADD_536_U168, P3_ADD_536_U169, P3_ADD_536_U17, P3_ADD_536_U170, P3_ADD_536_U171, P3_ADD_536_U172, P3_ADD_536_U173, P3_ADD_536_U174, P3_ADD_536_U175, P3_ADD_536_U176, P3_ADD_536_U177, P3_ADD_536_U178, P3_ADD_536_U179, P3_ADD_536_U18, P3_ADD_536_U180, P3_ADD_536_U181, P3_ADD_536_U182, P3_ADD_536_U19, P3_ADD_536_U20, P3_ADD_536_U21, P3_ADD_536_U22, P3_ADD_536_U23, P3_ADD_536_U24, P3_ADD_536_U25, P3_ADD_536_U26, P3_ADD_536_U27, P3_ADD_536_U28, P3_ADD_536_U29, P3_ADD_536_U30, P3_ADD_536_U31, P3_ADD_536_U32, P3_ADD_536_U33, P3_ADD_536_U34, P3_ADD_536_U35, P3_ADD_536_U36, P3_ADD_536_U37, P3_ADD_536_U38, P3_ADD_536_U39, P3_ADD_536_U4, P3_ADD_536_U40, P3_ADD_536_U41, P3_ADD_536_U42, P3_ADD_536_U43, P3_ADD_536_U44, P3_ADD_536_U45, P3_ADD_536_U46, P3_ADD_536_U47, P3_ADD_536_U48, P3_ADD_536_U49, P3_ADD_536_U5, P3_ADD_536_U50, P3_ADD_536_U51, P3_ADD_536_U52, P3_ADD_536_U53, P3_ADD_536_U54, P3_ADD_536_U55, P3_ADD_536_U56, P3_ADD_536_U57, P3_ADD_536_U58, P3_ADD_536_U59, P3_ADD_536_U6, P3_ADD_536_U60, P3_ADD_536_U61, P3_ADD_536_U62, P3_ADD_536_U63, P3_ADD_536_U64, P3_ADD_536_U65, P3_ADD_536_U66, P3_ADD_536_U67, P3_ADD_536_U68, P3_ADD_536_U69, P3_ADD_536_U7, P3_ADD_536_U70, P3_ADD_536_U71, P3_ADD_536_U72, P3_ADD_536_U73, P3_ADD_536_U74, P3_ADD_536_U75, P3_ADD_536_U76, P3_ADD_536_U77, P3_ADD_536_U78, P3_ADD_536_U79, P3_ADD_536_U8, P3_ADD_536_U80, P3_ADD_536_U81, P3_ADD_536_U82, P3_ADD_536_U83, P3_ADD_536_U84, P3_ADD_536_U85, P3_ADD_536_U86, P3_ADD_536_U87, P3_ADD_536_U88, P3_ADD_536_U89, P3_ADD_536_U9, P3_ADD_536_U90, P3_ADD_536_U91, P3_ADD_536_U92, P3_ADD_536_U93, P3_ADD_536_U94, P3_ADD_536_U95, P3_ADD_536_U96, P3_ADD_536_U97, P3_ADD_536_U98, P3_ADD_536_U99, P3_ADD_541_U10, P3_ADD_541_U100, P3_ADD_541_U101, P3_ADD_541_U102, P3_ADD_541_U103, P3_ADD_541_U104, P3_ADD_541_U105, P3_ADD_541_U106, P3_ADD_541_U107, P3_ADD_541_U108, P3_ADD_541_U109, P3_ADD_541_U11, P3_ADD_541_U110, P3_ADD_541_U111, P3_ADD_541_U112, P3_ADD_541_U113, P3_ADD_541_U114, P3_ADD_541_U115, P3_ADD_541_U116, P3_ADD_541_U117, P3_ADD_541_U118, P3_ADD_541_U119, P3_ADD_541_U12, P3_ADD_541_U120, P3_ADD_541_U121, P3_ADD_541_U122, P3_ADD_541_U123, P3_ADD_541_U124, P3_ADD_541_U125, P3_ADD_541_U126, P3_ADD_541_U127, P3_ADD_541_U128, P3_ADD_541_U129, P3_ADD_541_U13, P3_ADD_541_U130, P3_ADD_541_U131, P3_ADD_541_U132, P3_ADD_541_U133, P3_ADD_541_U134, P3_ADD_541_U135, P3_ADD_541_U136, P3_ADD_541_U137, P3_ADD_541_U138, P3_ADD_541_U139, P3_ADD_541_U14, P3_ADD_541_U140, P3_ADD_541_U141, P3_ADD_541_U142, P3_ADD_541_U143, P3_ADD_541_U144, P3_ADD_541_U145, P3_ADD_541_U146, P3_ADD_541_U147, P3_ADD_541_U148, P3_ADD_541_U149, P3_ADD_541_U15, P3_ADD_541_U150, P3_ADD_541_U151, P3_ADD_541_U152, P3_ADD_541_U153, P3_ADD_541_U154, P3_ADD_541_U155, P3_ADD_541_U156, P3_ADD_541_U157, P3_ADD_541_U158, P3_ADD_541_U159, P3_ADD_541_U16, P3_ADD_541_U160, P3_ADD_541_U161, P3_ADD_541_U162, P3_ADD_541_U163, P3_ADD_541_U164, P3_ADD_541_U165, P3_ADD_541_U166, P3_ADD_541_U167, P3_ADD_541_U168, P3_ADD_541_U169, P3_ADD_541_U17, P3_ADD_541_U170, P3_ADD_541_U171, P3_ADD_541_U172, P3_ADD_541_U173, P3_ADD_541_U174, P3_ADD_541_U175, P3_ADD_541_U176, P3_ADD_541_U177, P3_ADD_541_U178, P3_ADD_541_U179, P3_ADD_541_U18, P3_ADD_541_U180, P3_ADD_541_U181, P3_ADD_541_U182, P3_ADD_541_U19, P3_ADD_541_U20, P3_ADD_541_U21, P3_ADD_541_U22, P3_ADD_541_U23, P3_ADD_541_U24, P3_ADD_541_U25, P3_ADD_541_U26, P3_ADD_541_U27, P3_ADD_541_U28, P3_ADD_541_U29, P3_ADD_541_U30, P3_ADD_541_U31, P3_ADD_541_U32, P3_ADD_541_U33, P3_ADD_541_U34, P3_ADD_541_U35, P3_ADD_541_U36, P3_ADD_541_U37, P3_ADD_541_U38, P3_ADD_541_U39, P3_ADD_541_U4, P3_ADD_541_U40, P3_ADD_541_U41, P3_ADD_541_U42, P3_ADD_541_U43, P3_ADD_541_U44, P3_ADD_541_U45, P3_ADD_541_U46, P3_ADD_541_U47, P3_ADD_541_U48, P3_ADD_541_U49, P3_ADD_541_U5, P3_ADD_541_U50, P3_ADD_541_U51, P3_ADD_541_U52, P3_ADD_541_U53, P3_ADD_541_U54, P3_ADD_541_U55, P3_ADD_541_U56, P3_ADD_541_U57, P3_ADD_541_U58, P3_ADD_541_U59, P3_ADD_541_U6, P3_ADD_541_U60, P3_ADD_541_U61, P3_ADD_541_U62, P3_ADD_541_U63, P3_ADD_541_U64, P3_ADD_541_U65, P3_ADD_541_U66, P3_ADD_541_U67, P3_ADD_541_U68, P3_ADD_541_U69, P3_ADD_541_U7, P3_ADD_541_U70, P3_ADD_541_U71, P3_ADD_541_U72, P3_ADD_541_U73, P3_ADD_541_U74, P3_ADD_541_U75, P3_ADD_541_U76, P3_ADD_541_U77, P3_ADD_541_U78, P3_ADD_541_U79, P3_ADD_541_U8, P3_ADD_541_U80, P3_ADD_541_U81, P3_ADD_541_U82, P3_ADD_541_U83, P3_ADD_541_U84, P3_ADD_541_U85, P3_ADD_541_U86, P3_ADD_541_U87, P3_ADD_541_U88, P3_ADD_541_U89, P3_ADD_541_U9, P3_ADD_541_U90, P3_ADD_541_U91, P3_ADD_541_U92, P3_ADD_541_U93, P3_ADD_541_U94, P3_ADD_541_U95, P3_ADD_541_U96, P3_ADD_541_U97, P3_ADD_541_U98, P3_ADD_541_U99, P3_ADD_546_U10, P3_ADD_546_U100, P3_ADD_546_U101, P3_ADD_546_U102, P3_ADD_546_U103, P3_ADD_546_U104, P3_ADD_546_U105, P3_ADD_546_U106, P3_ADD_546_U107, P3_ADD_546_U108, P3_ADD_546_U109, P3_ADD_546_U11, P3_ADD_546_U110, P3_ADD_546_U111, P3_ADD_546_U112, P3_ADD_546_U113, P3_ADD_546_U114, P3_ADD_546_U115, P3_ADD_546_U116, P3_ADD_546_U117, P3_ADD_546_U118, P3_ADD_546_U119, P3_ADD_546_U12, P3_ADD_546_U120, P3_ADD_546_U121, P3_ADD_546_U122, P3_ADD_546_U123, P3_ADD_546_U124, P3_ADD_546_U125, P3_ADD_546_U126, P3_ADD_546_U127, P3_ADD_546_U128, P3_ADD_546_U129, P3_ADD_546_U13, P3_ADD_546_U130, P3_ADD_546_U131, P3_ADD_546_U132, P3_ADD_546_U133, P3_ADD_546_U134, P3_ADD_546_U135, P3_ADD_546_U136, P3_ADD_546_U137, P3_ADD_546_U138, P3_ADD_546_U139, P3_ADD_546_U14, P3_ADD_546_U140, P3_ADD_546_U141, P3_ADD_546_U142, P3_ADD_546_U143, P3_ADD_546_U144, P3_ADD_546_U145, P3_ADD_546_U146, P3_ADD_546_U147, P3_ADD_546_U148, P3_ADD_546_U149, P3_ADD_546_U15, P3_ADD_546_U150, P3_ADD_546_U151, P3_ADD_546_U152, P3_ADD_546_U153, P3_ADD_546_U154, P3_ADD_546_U155, P3_ADD_546_U156, P3_ADD_546_U157, P3_ADD_546_U158, P3_ADD_546_U159, P3_ADD_546_U16, P3_ADD_546_U160, P3_ADD_546_U161, P3_ADD_546_U162, P3_ADD_546_U163, P3_ADD_546_U164, P3_ADD_546_U165, P3_ADD_546_U166, P3_ADD_546_U167, P3_ADD_546_U168, P3_ADD_546_U169, P3_ADD_546_U17, P3_ADD_546_U170, P3_ADD_546_U171, P3_ADD_546_U172, P3_ADD_546_U173, P3_ADD_546_U174, P3_ADD_546_U175, P3_ADD_546_U176, P3_ADD_546_U177, P3_ADD_546_U178, P3_ADD_546_U179, P3_ADD_546_U18, P3_ADD_546_U180, P3_ADD_546_U181, P3_ADD_546_U182, P3_ADD_546_U183, P3_ADD_546_U184, P3_ADD_546_U185, P3_ADD_546_U186, P3_ADD_546_U187, P3_ADD_546_U188, P3_ADD_546_U189, P3_ADD_546_U19, P3_ADD_546_U190, P3_ADD_546_U191, P3_ADD_546_U192, P3_ADD_546_U193, P3_ADD_546_U194, P3_ADD_546_U195, P3_ADD_546_U196, P3_ADD_546_U197, P3_ADD_546_U198, P3_ADD_546_U199, P3_ADD_546_U20, P3_ADD_546_U200, P3_ADD_546_U201, P3_ADD_546_U202, P3_ADD_546_U21, P3_ADD_546_U22, P3_ADD_546_U23, P3_ADD_546_U24, P3_ADD_546_U25, P3_ADD_546_U26, P3_ADD_546_U27, P3_ADD_546_U28, P3_ADD_546_U29, P3_ADD_546_U30, P3_ADD_546_U31, P3_ADD_546_U32, P3_ADD_546_U33, P3_ADD_546_U34, P3_ADD_546_U35, P3_ADD_546_U36, P3_ADD_546_U37, P3_ADD_546_U38, P3_ADD_546_U39, P3_ADD_546_U40, P3_ADD_546_U41, P3_ADD_546_U42, P3_ADD_546_U43, P3_ADD_546_U44, P3_ADD_546_U45, P3_ADD_546_U46, P3_ADD_546_U47, P3_ADD_546_U48, P3_ADD_546_U49, P3_ADD_546_U5, P3_ADD_546_U50, P3_ADD_546_U51, P3_ADD_546_U52, P3_ADD_546_U53, P3_ADD_546_U54, P3_ADD_546_U55, P3_ADD_546_U56, P3_ADD_546_U57, P3_ADD_546_U58, P3_ADD_546_U59, P3_ADD_546_U6, P3_ADD_546_U60, P3_ADD_546_U61, P3_ADD_546_U62, P3_ADD_546_U63, P3_ADD_546_U64, P3_ADD_546_U65, P3_ADD_546_U66, P3_ADD_546_U67, P3_ADD_546_U68, P3_ADD_546_U69, P3_ADD_546_U7, P3_ADD_546_U70, P3_ADD_546_U71, P3_ADD_546_U72, P3_ADD_546_U73, P3_ADD_546_U74, P3_ADD_546_U75, P3_ADD_546_U76, P3_ADD_546_U77, P3_ADD_546_U78, P3_ADD_546_U79, P3_ADD_546_U8, P3_ADD_546_U80, P3_ADD_546_U81, P3_ADD_546_U82, P3_ADD_546_U83, P3_ADD_546_U84, P3_ADD_546_U85, P3_ADD_546_U86, P3_ADD_546_U87, P3_ADD_546_U88, P3_ADD_546_U89, P3_ADD_546_U9, P3_ADD_546_U90, P3_ADD_546_U91, P3_ADD_546_U92, P3_ADD_546_U93, P3_ADD_546_U94, P3_ADD_546_U95, P3_ADD_546_U96, P3_ADD_546_U97, P3_ADD_546_U98, P3_ADD_546_U99, P3_ADD_547_U10, P3_ADD_547_U100, P3_ADD_547_U101, P3_ADD_547_U102, P3_ADD_547_U103, P3_ADD_547_U104, P3_ADD_547_U105, P3_ADD_547_U106, P3_ADD_547_U107, P3_ADD_547_U108, P3_ADD_547_U109, P3_ADD_547_U11, P3_ADD_547_U110, P3_ADD_547_U111, P3_ADD_547_U112, P3_ADD_547_U113, P3_ADD_547_U114, P3_ADD_547_U115, P3_ADD_547_U116, P3_ADD_547_U117, P3_ADD_547_U118, P3_ADD_547_U119, P3_ADD_547_U12, P3_ADD_547_U120, P3_ADD_547_U121, P3_ADD_547_U122, P3_ADD_547_U123, P3_ADD_547_U124, P3_ADD_547_U125, P3_ADD_547_U126, P3_ADD_547_U127, P3_ADD_547_U128, P3_ADD_547_U129, P3_ADD_547_U13, P3_ADD_547_U130, P3_ADD_547_U131, P3_ADD_547_U132, P3_ADD_547_U133, P3_ADD_547_U134, P3_ADD_547_U135, P3_ADD_547_U136, P3_ADD_547_U137, P3_ADD_547_U138, P3_ADD_547_U139, P3_ADD_547_U14, P3_ADD_547_U140, P3_ADD_547_U141, P3_ADD_547_U142, P3_ADD_547_U143, P3_ADD_547_U144, P3_ADD_547_U145, P3_ADD_547_U146, P3_ADD_547_U147, P3_ADD_547_U148, P3_ADD_547_U149, P3_ADD_547_U15, P3_ADD_547_U150, P3_ADD_547_U151, P3_ADD_547_U152, P3_ADD_547_U153, P3_ADD_547_U154, P3_ADD_547_U155, P3_ADD_547_U156, P3_ADD_547_U157, P3_ADD_547_U158, P3_ADD_547_U159, P3_ADD_547_U16, P3_ADD_547_U160, P3_ADD_547_U161, P3_ADD_547_U162, P3_ADD_547_U163, P3_ADD_547_U164, P3_ADD_547_U165, P3_ADD_547_U166, P3_ADD_547_U167, P3_ADD_547_U168, P3_ADD_547_U169, P3_ADD_547_U17, P3_ADD_547_U170, P3_ADD_547_U171, P3_ADD_547_U172, P3_ADD_547_U173, P3_ADD_547_U174, P3_ADD_547_U175, P3_ADD_547_U176, P3_ADD_547_U177, P3_ADD_547_U178, P3_ADD_547_U179, P3_ADD_547_U18, P3_ADD_547_U180, P3_ADD_547_U181, P3_ADD_547_U182, P3_ADD_547_U183, P3_ADD_547_U184, P3_ADD_547_U185, P3_ADD_547_U186, P3_ADD_547_U187, P3_ADD_547_U188, P3_ADD_547_U189, P3_ADD_547_U19, P3_ADD_547_U20, P3_ADD_547_U21, P3_ADD_547_U22, P3_ADD_547_U23, P3_ADD_547_U24, P3_ADD_547_U25, P3_ADD_547_U26, P3_ADD_547_U27, P3_ADD_547_U28, P3_ADD_547_U29, P3_ADD_547_U30, P3_ADD_547_U31, P3_ADD_547_U32, P3_ADD_547_U33, P3_ADD_547_U34, P3_ADD_547_U35, P3_ADD_547_U36, P3_ADD_547_U37, P3_ADD_547_U38, P3_ADD_547_U39, P3_ADD_547_U40, P3_ADD_547_U41, P3_ADD_547_U42, P3_ADD_547_U43, P3_ADD_547_U44, P3_ADD_547_U45, P3_ADD_547_U46, P3_ADD_547_U47, P3_ADD_547_U48, P3_ADD_547_U49, P3_ADD_547_U5, P3_ADD_547_U50, P3_ADD_547_U51, P3_ADD_547_U52, P3_ADD_547_U53, P3_ADD_547_U54, P3_ADD_547_U55, P3_ADD_547_U56, P3_ADD_547_U57, P3_ADD_547_U58, P3_ADD_547_U59, P3_ADD_547_U6, P3_ADD_547_U60, P3_ADD_547_U61, P3_ADD_547_U62, P3_ADD_547_U63, P3_ADD_547_U64, P3_ADD_547_U65, P3_ADD_547_U66, P3_ADD_547_U67, P3_ADD_547_U68, P3_ADD_547_U69, P3_ADD_547_U7, P3_ADD_547_U70, P3_ADD_547_U71, P3_ADD_547_U72, P3_ADD_547_U73, P3_ADD_547_U74, P3_ADD_547_U75, P3_ADD_547_U76, P3_ADD_547_U77, P3_ADD_547_U78, P3_ADD_547_U79, P3_ADD_547_U8, P3_ADD_547_U80, P3_ADD_547_U81, P3_ADD_547_U82, P3_ADD_547_U83, P3_ADD_547_U84, P3_ADD_547_U85, P3_ADD_547_U86, P3_ADD_547_U87, P3_ADD_547_U88, P3_ADD_547_U89, P3_ADD_547_U9, P3_ADD_547_U90, P3_ADD_547_U91, P3_ADD_547_U92, P3_ADD_547_U93, P3_ADD_547_U94, P3_ADD_547_U95, P3_ADD_547_U96, P3_ADD_547_U97, P3_ADD_547_U98, P3_ADD_547_U99, P3_ADD_552_U10, P3_ADD_552_U100, P3_ADD_552_U101, P3_ADD_552_U102, P3_ADD_552_U103, P3_ADD_552_U104, P3_ADD_552_U105, P3_ADD_552_U106, P3_ADD_552_U107, P3_ADD_552_U108, P3_ADD_552_U109, P3_ADD_552_U11, P3_ADD_552_U110, P3_ADD_552_U111, P3_ADD_552_U112, P3_ADD_552_U113, P3_ADD_552_U114, P3_ADD_552_U115, P3_ADD_552_U116, P3_ADD_552_U117, P3_ADD_552_U118, P3_ADD_552_U119, P3_ADD_552_U12, P3_ADD_552_U120, P3_ADD_552_U121, P3_ADD_552_U122, P3_ADD_552_U123, P3_ADD_552_U124, P3_ADD_552_U125, P3_ADD_552_U126, P3_ADD_552_U127, P3_ADD_552_U128, P3_ADD_552_U129, P3_ADD_552_U13, P3_ADD_552_U130, P3_ADD_552_U131, P3_ADD_552_U132, P3_ADD_552_U133, P3_ADD_552_U134, P3_ADD_552_U135, P3_ADD_552_U136, P3_ADD_552_U137, P3_ADD_552_U138, P3_ADD_552_U139, P3_ADD_552_U14, P3_ADD_552_U140, P3_ADD_552_U141, P3_ADD_552_U142, P3_ADD_552_U143, P3_ADD_552_U144, P3_ADD_552_U145, P3_ADD_552_U146, P3_ADD_552_U147, P3_ADD_552_U148, P3_ADD_552_U149, P3_ADD_552_U15, P3_ADD_552_U150, P3_ADD_552_U151, P3_ADD_552_U152, P3_ADD_552_U153, P3_ADD_552_U154, P3_ADD_552_U155, P3_ADD_552_U156, P3_ADD_552_U157, P3_ADD_552_U158, P3_ADD_552_U159, P3_ADD_552_U16, P3_ADD_552_U160, P3_ADD_552_U161, P3_ADD_552_U162, P3_ADD_552_U163, P3_ADD_552_U164, P3_ADD_552_U165, P3_ADD_552_U166, P3_ADD_552_U167, P3_ADD_552_U168, P3_ADD_552_U169, P3_ADD_552_U17, P3_ADD_552_U170, P3_ADD_552_U171, P3_ADD_552_U172, P3_ADD_552_U173, P3_ADD_552_U174, P3_ADD_552_U175, P3_ADD_552_U176, P3_ADD_552_U177, P3_ADD_552_U178, P3_ADD_552_U179, P3_ADD_552_U18, P3_ADD_552_U180, P3_ADD_552_U181, P3_ADD_552_U182, P3_ADD_552_U183, P3_ADD_552_U184, P3_ADD_552_U185, P3_ADD_552_U186, P3_ADD_552_U187, P3_ADD_552_U188, P3_ADD_552_U189, P3_ADD_552_U19, P3_ADD_552_U190, P3_ADD_552_U191, P3_ADD_552_U192, P3_ADD_552_U193, P3_ADD_552_U194, P3_ADD_552_U195, P3_ADD_552_U196, P3_ADD_552_U197, P3_ADD_552_U198, P3_ADD_552_U199, P3_ADD_552_U20, P3_ADD_552_U200, P3_ADD_552_U201, P3_ADD_552_U202, P3_ADD_552_U21, P3_ADD_552_U22, P3_ADD_552_U23, P3_ADD_552_U24, P3_ADD_552_U25, P3_ADD_552_U26, P3_ADD_552_U27, P3_ADD_552_U28, P3_ADD_552_U29, P3_ADD_552_U30, P3_ADD_552_U31, P3_ADD_552_U32, P3_ADD_552_U33, P3_ADD_552_U34, P3_ADD_552_U35, P3_ADD_552_U36, P3_ADD_552_U37, P3_ADD_552_U38, P3_ADD_552_U39, P3_ADD_552_U40, P3_ADD_552_U41, P3_ADD_552_U42, P3_ADD_552_U43, P3_ADD_552_U44, P3_ADD_552_U45, P3_ADD_552_U46, P3_ADD_552_U47, P3_ADD_552_U48, P3_ADD_552_U49, P3_ADD_552_U5, P3_ADD_552_U50, P3_ADD_552_U51, P3_ADD_552_U52, P3_ADD_552_U53, P3_ADD_552_U54, P3_ADD_552_U55, P3_ADD_552_U56, P3_ADD_552_U57, P3_ADD_552_U58, P3_ADD_552_U59, P3_ADD_552_U6, P3_ADD_552_U60, P3_ADD_552_U61, P3_ADD_552_U62, P3_ADD_552_U63, P3_ADD_552_U64, P3_ADD_552_U65, P3_ADD_552_U66, P3_ADD_552_U67, P3_ADD_552_U68, P3_ADD_552_U69, P3_ADD_552_U7, P3_ADD_552_U70, P3_ADD_552_U71, P3_ADD_552_U72, P3_ADD_552_U73, P3_ADD_552_U74, P3_ADD_552_U75, P3_ADD_552_U76, P3_ADD_552_U77, P3_ADD_552_U78, P3_ADD_552_U79, P3_ADD_552_U8, P3_ADD_552_U80, P3_ADD_552_U81, P3_ADD_552_U82, P3_ADD_552_U83, P3_ADD_552_U84, P3_ADD_552_U85, P3_ADD_552_U86, P3_ADD_552_U87, P3_ADD_552_U88, P3_ADD_552_U89, P3_ADD_552_U9, P3_ADD_552_U90, P3_ADD_552_U91, P3_ADD_552_U92, P3_ADD_552_U93, P3_ADD_552_U94, P3_ADD_552_U95, P3_ADD_552_U96, P3_ADD_552_U97, P3_ADD_552_U98, P3_ADD_552_U99, P3_ADD_553_U10, P3_ADD_553_U100, P3_ADD_553_U101, P3_ADD_553_U102, P3_ADD_553_U103, P3_ADD_553_U104, P3_ADD_553_U105, P3_ADD_553_U106, P3_ADD_553_U107, P3_ADD_553_U108, P3_ADD_553_U109, P3_ADD_553_U11, P3_ADD_553_U110, P3_ADD_553_U111, P3_ADD_553_U112, P3_ADD_553_U113, P3_ADD_553_U114, P3_ADD_553_U115, P3_ADD_553_U116, P3_ADD_553_U117, P3_ADD_553_U118, P3_ADD_553_U119, P3_ADD_553_U12, P3_ADD_553_U120, P3_ADD_553_U121, P3_ADD_553_U122, P3_ADD_553_U123, P3_ADD_553_U124, P3_ADD_553_U125, P3_ADD_553_U126, P3_ADD_553_U127, P3_ADD_553_U128, P3_ADD_553_U129, P3_ADD_553_U13, P3_ADD_553_U130, P3_ADD_553_U131, P3_ADD_553_U132, P3_ADD_553_U133, P3_ADD_553_U134, P3_ADD_553_U135, P3_ADD_553_U136, P3_ADD_553_U137, P3_ADD_553_U138, P3_ADD_553_U139, P3_ADD_553_U14, P3_ADD_553_U140, P3_ADD_553_U141, P3_ADD_553_U142, P3_ADD_553_U143, P3_ADD_553_U144, P3_ADD_553_U145, P3_ADD_553_U146, P3_ADD_553_U147, P3_ADD_553_U148, P3_ADD_553_U149, P3_ADD_553_U15, P3_ADD_553_U150, P3_ADD_553_U151, P3_ADD_553_U152, P3_ADD_553_U153, P3_ADD_553_U154, P3_ADD_553_U155, P3_ADD_553_U156, P3_ADD_553_U157, P3_ADD_553_U158, P3_ADD_553_U159, P3_ADD_553_U16, P3_ADD_553_U160, P3_ADD_553_U161, P3_ADD_553_U162, P3_ADD_553_U163, P3_ADD_553_U164, P3_ADD_553_U165, P3_ADD_553_U166, P3_ADD_553_U167, P3_ADD_553_U168, P3_ADD_553_U169, P3_ADD_553_U17, P3_ADD_553_U170, P3_ADD_553_U171, P3_ADD_553_U172, P3_ADD_553_U173, P3_ADD_553_U174, P3_ADD_553_U175, P3_ADD_553_U176, P3_ADD_553_U177, P3_ADD_553_U178, P3_ADD_553_U179, P3_ADD_553_U18, P3_ADD_553_U180, P3_ADD_553_U181, P3_ADD_553_U182, P3_ADD_553_U183, P3_ADD_553_U184, P3_ADD_553_U185, P3_ADD_553_U186, P3_ADD_553_U187, P3_ADD_553_U188, P3_ADD_553_U189, P3_ADD_553_U19, P3_ADD_553_U20, P3_ADD_553_U21, P3_ADD_553_U22, P3_ADD_553_U23, P3_ADD_553_U24, P3_ADD_553_U25, P3_ADD_553_U26, P3_ADD_553_U27, P3_ADD_553_U28, P3_ADD_553_U29, P3_ADD_553_U30, P3_ADD_553_U31, P3_ADD_553_U32, P3_ADD_553_U33, P3_ADD_553_U34, P3_ADD_553_U35, P3_ADD_553_U36, P3_ADD_553_U37, P3_ADD_553_U38, P3_ADD_553_U39, P3_ADD_553_U40, P3_ADD_553_U41, P3_ADD_553_U42, P3_ADD_553_U43, P3_ADD_553_U44, P3_ADD_553_U45, P3_ADD_553_U46, P3_ADD_553_U47, P3_ADD_553_U48, P3_ADD_553_U49, P3_ADD_553_U5, P3_ADD_553_U50, P3_ADD_553_U51, P3_ADD_553_U52, P3_ADD_553_U53, P3_ADD_553_U54, P3_ADD_553_U55, P3_ADD_553_U56, P3_ADD_553_U57, P3_ADD_553_U58, P3_ADD_553_U59, P3_ADD_553_U6, P3_ADD_553_U60, P3_ADD_553_U61, P3_ADD_553_U62, P3_ADD_553_U63, P3_ADD_553_U64, P3_ADD_553_U65, P3_ADD_553_U66, P3_ADD_553_U67, P3_ADD_553_U68, P3_ADD_553_U69, P3_ADD_553_U7, P3_ADD_553_U70, P3_ADD_553_U71, P3_ADD_553_U72, P3_ADD_553_U73, P3_ADD_553_U74, P3_ADD_553_U75, P3_ADD_553_U76, P3_ADD_553_U77, P3_ADD_553_U78, P3_ADD_553_U79, P3_ADD_553_U8, P3_ADD_553_U80, P3_ADD_553_U81, P3_ADD_553_U82, P3_ADD_553_U83, P3_ADD_553_U84, P3_ADD_553_U85, P3_ADD_553_U86, P3_ADD_553_U87, P3_ADD_553_U88, P3_ADD_553_U89, P3_ADD_553_U9, P3_ADD_553_U90, P3_ADD_553_U91, P3_ADD_553_U92, P3_ADD_553_U93, P3_ADD_553_U94, P3_ADD_553_U95, P3_ADD_553_U96, P3_ADD_553_U97, P3_ADD_553_U98, P3_ADD_553_U99, P3_ADD_558_U10, P3_ADD_558_U100, P3_ADD_558_U101, P3_ADD_558_U102, P3_ADD_558_U103, P3_ADD_558_U104, P3_ADD_558_U105, P3_ADD_558_U106, P3_ADD_558_U107, P3_ADD_558_U108, P3_ADD_558_U109, P3_ADD_558_U11, P3_ADD_558_U110, P3_ADD_558_U111, P3_ADD_558_U112, P3_ADD_558_U113, P3_ADD_558_U114, P3_ADD_558_U115, P3_ADD_558_U116, P3_ADD_558_U117, P3_ADD_558_U118, P3_ADD_558_U119, P3_ADD_558_U12, P3_ADD_558_U120, P3_ADD_558_U121, P3_ADD_558_U122, P3_ADD_558_U123, P3_ADD_558_U124, P3_ADD_558_U125, P3_ADD_558_U126, P3_ADD_558_U127, P3_ADD_558_U128, P3_ADD_558_U129, P3_ADD_558_U13, P3_ADD_558_U130, P3_ADD_558_U131, P3_ADD_558_U132, P3_ADD_558_U133, P3_ADD_558_U134, P3_ADD_558_U135, P3_ADD_558_U136, P3_ADD_558_U137, P3_ADD_558_U138, P3_ADD_558_U139, P3_ADD_558_U14, P3_ADD_558_U140, P3_ADD_558_U141, P3_ADD_558_U142, P3_ADD_558_U143, P3_ADD_558_U144, P3_ADD_558_U145, P3_ADD_558_U146, P3_ADD_558_U147, P3_ADD_558_U148, P3_ADD_558_U149, P3_ADD_558_U15, P3_ADD_558_U150, P3_ADD_558_U151, P3_ADD_558_U152, P3_ADD_558_U153, P3_ADD_558_U154, P3_ADD_558_U155, P3_ADD_558_U156, P3_ADD_558_U157, P3_ADD_558_U158, P3_ADD_558_U159, P3_ADD_558_U16, P3_ADD_558_U160, P3_ADD_558_U161, P3_ADD_558_U162, P3_ADD_558_U163, P3_ADD_558_U164, P3_ADD_558_U165, P3_ADD_558_U166, P3_ADD_558_U167, P3_ADD_558_U168, P3_ADD_558_U169, P3_ADD_558_U17, P3_ADD_558_U170, P3_ADD_558_U171, P3_ADD_558_U172, P3_ADD_558_U173, P3_ADD_558_U174, P3_ADD_558_U175, P3_ADD_558_U176, P3_ADD_558_U177, P3_ADD_558_U178, P3_ADD_558_U179, P3_ADD_558_U18, P3_ADD_558_U180, P3_ADD_558_U181, P3_ADD_558_U182, P3_ADD_558_U183, P3_ADD_558_U184, P3_ADD_558_U185, P3_ADD_558_U186, P3_ADD_558_U187, P3_ADD_558_U188, P3_ADD_558_U189, P3_ADD_558_U19, P3_ADD_558_U20, P3_ADD_558_U21, P3_ADD_558_U22, P3_ADD_558_U23, P3_ADD_558_U24, P3_ADD_558_U25, P3_ADD_558_U26, P3_ADD_558_U27, P3_ADD_558_U28, P3_ADD_558_U29, P3_ADD_558_U30, P3_ADD_558_U31, P3_ADD_558_U32, P3_ADD_558_U33, P3_ADD_558_U34, P3_ADD_558_U35, P3_ADD_558_U36, P3_ADD_558_U37, P3_ADD_558_U38, P3_ADD_558_U39, P3_ADD_558_U40, P3_ADD_558_U41, P3_ADD_558_U42, P3_ADD_558_U43, P3_ADD_558_U44, P3_ADD_558_U45, P3_ADD_558_U46, P3_ADD_558_U47, P3_ADD_558_U48, P3_ADD_558_U49, P3_ADD_558_U5, P3_ADD_558_U50, P3_ADD_558_U51, P3_ADD_558_U52, P3_ADD_558_U53, P3_ADD_558_U54, P3_ADD_558_U55, P3_ADD_558_U56, P3_ADD_558_U57, P3_ADD_558_U58, P3_ADD_558_U59, P3_ADD_558_U6, P3_ADD_558_U60, P3_ADD_558_U61, P3_ADD_558_U62, P3_ADD_558_U63, P3_ADD_558_U64, P3_ADD_558_U65, P3_ADD_558_U66, P3_ADD_558_U67, P3_ADD_558_U68, P3_ADD_558_U69, P3_ADD_558_U7, P3_ADD_558_U70, P3_ADD_558_U71, P3_ADD_558_U72, P3_ADD_558_U73, P3_ADD_558_U74, P3_ADD_558_U75, P3_ADD_558_U76, P3_ADD_558_U77, P3_ADD_558_U78, P3_ADD_558_U79, P3_ADD_558_U8, P3_ADD_558_U80, P3_ADD_558_U81, P3_ADD_558_U82, P3_ADD_558_U83, P3_ADD_558_U84, P3_ADD_558_U85, P3_ADD_558_U86, P3_ADD_558_U87, P3_ADD_558_U88, P3_ADD_558_U89, P3_ADD_558_U9, P3_ADD_558_U90, P3_ADD_558_U91, P3_ADD_558_U92, P3_ADD_558_U93, P3_ADD_558_U94, P3_ADD_558_U95, P3_ADD_558_U96, P3_ADD_558_U97, P3_ADD_558_U98, P3_ADD_558_U99, P3_GTE_355_U6, P3_GTE_355_U7, P3_GTE_355_U8, P3_GTE_370_U6, P3_GTE_370_U7, P3_GTE_370_U8, P3_GTE_370_U9, P3_GTE_390_U6, P3_GTE_390_U7, P3_GTE_390_U8, P3_GTE_390_U9, P3_GTE_401_U6, P3_GTE_401_U7, P3_GTE_401_U8, P3_GTE_401_U9, P3_GTE_412_U6, P3_GTE_412_U7, P3_GTE_450_U6, P3_GTE_450_U7, P3_GTE_485_U6, P3_GTE_485_U7, P3_GTE_504_U6, P3_GTE_504_U7, P3_LTE_597_U6, P3_LT_563_1260_U6, P3_LT_563_1260_U7, P3_LT_563_U10, P3_LT_563_U11, P3_LT_563_U12, P3_LT_563_U13, P3_LT_563_U14, P3_LT_563_U15, P3_LT_563_U16, P3_LT_563_U17, P3_LT_563_U18, P3_LT_563_U19, P3_LT_563_U20, P3_LT_563_U21, P3_LT_563_U22, P3_LT_563_U23, P3_LT_563_U24, P3_LT_563_U25, P3_LT_563_U26, P3_LT_563_U27, P3_LT_563_U28, P3_LT_563_U6, P3_LT_563_U7, P3_LT_563_U8, P3_LT_563_U9, P3_LT_589_U6, P3_LT_589_U7, P3_LT_589_U8, P3_SUB_320_U10, P3_SUB_320_U100, P3_SUB_320_U101, P3_SUB_320_U102, P3_SUB_320_U103, P3_SUB_320_U104, P3_SUB_320_U105, P3_SUB_320_U106, P3_SUB_320_U107, P3_SUB_320_U108, P3_SUB_320_U109, P3_SUB_320_U11, P3_SUB_320_U110, P3_SUB_320_U111, P3_SUB_320_U112, P3_SUB_320_U113, P3_SUB_320_U114, P3_SUB_320_U115, P3_SUB_320_U116, P3_SUB_320_U117, P3_SUB_320_U118, P3_SUB_320_U119, P3_SUB_320_U12, P3_SUB_320_U120, P3_SUB_320_U121, P3_SUB_320_U122, P3_SUB_320_U123, P3_SUB_320_U124, P3_SUB_320_U125, P3_SUB_320_U126, P3_SUB_320_U127, P3_SUB_320_U128, P3_SUB_320_U129, P3_SUB_320_U13, P3_SUB_320_U130, P3_SUB_320_U131, P3_SUB_320_U132, P3_SUB_320_U133, P3_SUB_320_U134, P3_SUB_320_U135, P3_SUB_320_U136, P3_SUB_320_U137, P3_SUB_320_U138, P3_SUB_320_U139, P3_SUB_320_U14, P3_SUB_320_U140, P3_SUB_320_U141, P3_SUB_320_U142, P3_SUB_320_U143, P3_SUB_320_U144, P3_SUB_320_U145, P3_SUB_320_U146, P3_SUB_320_U147, P3_SUB_320_U148, P3_SUB_320_U149, P3_SUB_320_U15, P3_SUB_320_U150, P3_SUB_320_U151, P3_SUB_320_U152, P3_SUB_320_U153, P3_SUB_320_U154, P3_SUB_320_U155, P3_SUB_320_U156, P3_SUB_320_U157, P3_SUB_320_U158, P3_SUB_320_U159, P3_SUB_320_U16, P3_SUB_320_U17, P3_SUB_320_U18, P3_SUB_320_U19, P3_SUB_320_U20, P3_SUB_320_U21, P3_SUB_320_U22, P3_SUB_320_U23, P3_SUB_320_U24, P3_SUB_320_U25, P3_SUB_320_U26, P3_SUB_320_U27, P3_SUB_320_U28, P3_SUB_320_U29, P3_SUB_320_U30, P3_SUB_320_U31, P3_SUB_320_U32, P3_SUB_320_U33, P3_SUB_320_U34, P3_SUB_320_U35, P3_SUB_320_U36, P3_SUB_320_U37, P3_SUB_320_U38, P3_SUB_320_U39, P3_SUB_320_U40, P3_SUB_320_U41, P3_SUB_320_U42, P3_SUB_320_U43, P3_SUB_320_U44, P3_SUB_320_U45, P3_SUB_320_U46, P3_SUB_320_U47, P3_SUB_320_U48, P3_SUB_320_U49, P3_SUB_320_U50, P3_SUB_320_U51, P3_SUB_320_U52, P3_SUB_320_U53, P3_SUB_320_U54, P3_SUB_320_U55, P3_SUB_320_U56, P3_SUB_320_U57, P3_SUB_320_U58, P3_SUB_320_U59, P3_SUB_320_U6, P3_SUB_320_U60, P3_SUB_320_U61, P3_SUB_320_U62, P3_SUB_320_U63, P3_SUB_320_U64, P3_SUB_320_U65, P3_SUB_320_U66, P3_SUB_320_U67, P3_SUB_320_U68, P3_SUB_320_U69, P3_SUB_320_U7, P3_SUB_320_U70, P3_SUB_320_U71, P3_SUB_320_U72, P3_SUB_320_U73, P3_SUB_320_U74, P3_SUB_320_U75, P3_SUB_320_U76, P3_SUB_320_U77, P3_SUB_320_U78, P3_SUB_320_U79, P3_SUB_320_U8, P3_SUB_320_U80, P3_SUB_320_U81, P3_SUB_320_U82, P3_SUB_320_U83, P3_SUB_320_U84, P3_SUB_320_U85, P3_SUB_320_U86, P3_SUB_320_U87, P3_SUB_320_U88, P3_SUB_320_U89, P3_SUB_320_U9, P3_SUB_320_U90, P3_SUB_320_U91, P3_SUB_320_U92, P3_SUB_320_U93, P3_SUB_320_U94, P3_SUB_320_U95, P3_SUB_320_U96, P3_SUB_320_U97, P3_SUB_320_U98, P3_SUB_320_U99, P3_SUB_355_U10, P3_SUB_355_U11, P3_SUB_355_U12, P3_SUB_355_U13, P3_SUB_355_U14, P3_SUB_355_U15, P3_SUB_355_U16, P3_SUB_355_U17, P3_SUB_355_U18, P3_SUB_355_U19, P3_SUB_355_U20, P3_SUB_355_U21, P3_SUB_355_U22, P3_SUB_355_U23, P3_SUB_355_U24, P3_SUB_355_U25, P3_SUB_355_U26, P3_SUB_355_U27, P3_SUB_355_U28, P3_SUB_355_U29, P3_SUB_355_U30, P3_SUB_355_U31, P3_SUB_355_U32, P3_SUB_355_U33, P3_SUB_355_U34, P3_SUB_355_U35, P3_SUB_355_U36, P3_SUB_355_U37, P3_SUB_355_U38, P3_SUB_355_U39, P3_SUB_355_U40, P3_SUB_355_U41, P3_SUB_355_U42, P3_SUB_355_U43, P3_SUB_355_U44, P3_SUB_355_U45, P3_SUB_355_U46, P3_SUB_355_U47, P3_SUB_355_U48, P3_SUB_355_U49, P3_SUB_355_U50, P3_SUB_355_U51, P3_SUB_355_U52, P3_SUB_355_U53, P3_SUB_355_U54, P3_SUB_355_U55, P3_SUB_355_U56, P3_SUB_355_U57, P3_SUB_355_U58, P3_SUB_355_U59, P3_SUB_355_U6, P3_SUB_355_U60, P3_SUB_355_U61, P3_SUB_355_U62, P3_SUB_355_U63, P3_SUB_355_U64, P3_SUB_355_U65, P3_SUB_355_U66, P3_SUB_355_U7, P3_SUB_355_U8, P3_SUB_355_U9, P3_SUB_357_1258_U10, P3_SUB_357_1258_U100, P3_SUB_357_1258_U101, P3_SUB_357_1258_U102, P3_SUB_357_1258_U103, P3_SUB_357_1258_U104, P3_SUB_357_1258_U105, P3_SUB_357_1258_U106, P3_SUB_357_1258_U107, P3_SUB_357_1258_U108, P3_SUB_357_1258_U109, P3_SUB_357_1258_U11, P3_SUB_357_1258_U110, P3_SUB_357_1258_U111, P3_SUB_357_1258_U112, P3_SUB_357_1258_U113, P3_SUB_357_1258_U114, P3_SUB_357_1258_U115, P3_SUB_357_1258_U116, P3_SUB_357_1258_U117, P3_SUB_357_1258_U118, P3_SUB_357_1258_U119, P3_SUB_357_1258_U12, P3_SUB_357_1258_U120, P3_SUB_357_1258_U121, P3_SUB_357_1258_U122, P3_SUB_357_1258_U123, P3_SUB_357_1258_U124, P3_SUB_357_1258_U125, P3_SUB_357_1258_U126, P3_SUB_357_1258_U127, P3_SUB_357_1258_U128, P3_SUB_357_1258_U129, P3_SUB_357_1258_U13, P3_SUB_357_1258_U130, P3_SUB_357_1258_U131, P3_SUB_357_1258_U132, P3_SUB_357_1258_U133, P3_SUB_357_1258_U134, P3_SUB_357_1258_U135, P3_SUB_357_1258_U136, P3_SUB_357_1258_U137, P3_SUB_357_1258_U138, P3_SUB_357_1258_U139, P3_SUB_357_1258_U14, P3_SUB_357_1258_U140, P3_SUB_357_1258_U141, P3_SUB_357_1258_U142, P3_SUB_357_1258_U143, P3_SUB_357_1258_U144, P3_SUB_357_1258_U145, P3_SUB_357_1258_U146, P3_SUB_357_1258_U147, P3_SUB_357_1258_U148, P3_SUB_357_1258_U149, P3_SUB_357_1258_U15, P3_SUB_357_1258_U150, P3_SUB_357_1258_U151, P3_SUB_357_1258_U152, P3_SUB_357_1258_U153, P3_SUB_357_1258_U154, P3_SUB_357_1258_U155, P3_SUB_357_1258_U156, P3_SUB_357_1258_U157, P3_SUB_357_1258_U158, P3_SUB_357_1258_U159, P3_SUB_357_1258_U16, P3_SUB_357_1258_U160, P3_SUB_357_1258_U161, P3_SUB_357_1258_U162, P3_SUB_357_1258_U163, P3_SUB_357_1258_U164, P3_SUB_357_1258_U165, P3_SUB_357_1258_U166, P3_SUB_357_1258_U167, P3_SUB_357_1258_U168, P3_SUB_357_1258_U169, P3_SUB_357_1258_U17, P3_SUB_357_1258_U170, P3_SUB_357_1258_U171, P3_SUB_357_1258_U172, P3_SUB_357_1258_U173, P3_SUB_357_1258_U174, P3_SUB_357_1258_U175, P3_SUB_357_1258_U176, P3_SUB_357_1258_U177, P3_SUB_357_1258_U178, P3_SUB_357_1258_U179, P3_SUB_357_1258_U18, P3_SUB_357_1258_U180, P3_SUB_357_1258_U181, P3_SUB_357_1258_U182, P3_SUB_357_1258_U183, P3_SUB_357_1258_U184, P3_SUB_357_1258_U185, P3_SUB_357_1258_U186, P3_SUB_357_1258_U187, P3_SUB_357_1258_U188, P3_SUB_357_1258_U189, P3_SUB_357_1258_U19, P3_SUB_357_1258_U190, P3_SUB_357_1258_U191, P3_SUB_357_1258_U192, P3_SUB_357_1258_U193, P3_SUB_357_1258_U194, P3_SUB_357_1258_U195, P3_SUB_357_1258_U196, P3_SUB_357_1258_U197, P3_SUB_357_1258_U198, P3_SUB_357_1258_U199, P3_SUB_357_1258_U20, P3_SUB_357_1258_U200, P3_SUB_357_1258_U201, P3_SUB_357_1258_U202, P3_SUB_357_1258_U203, P3_SUB_357_1258_U204, P3_SUB_357_1258_U205, P3_SUB_357_1258_U206, P3_SUB_357_1258_U207, P3_SUB_357_1258_U208, P3_SUB_357_1258_U209, P3_SUB_357_1258_U21, P3_SUB_357_1258_U210, P3_SUB_357_1258_U211, P3_SUB_357_1258_U212, P3_SUB_357_1258_U213, P3_SUB_357_1258_U214, P3_SUB_357_1258_U215, P3_SUB_357_1258_U216, P3_SUB_357_1258_U217, P3_SUB_357_1258_U218, P3_SUB_357_1258_U219, P3_SUB_357_1258_U22, P3_SUB_357_1258_U220, P3_SUB_357_1258_U221, P3_SUB_357_1258_U222, P3_SUB_357_1258_U223, P3_SUB_357_1258_U224, P3_SUB_357_1258_U225, P3_SUB_357_1258_U226, P3_SUB_357_1258_U227, P3_SUB_357_1258_U228, P3_SUB_357_1258_U229, P3_SUB_357_1258_U23, P3_SUB_357_1258_U230, P3_SUB_357_1258_U231, P3_SUB_357_1258_U232, P3_SUB_357_1258_U233, P3_SUB_357_1258_U234, P3_SUB_357_1258_U235, P3_SUB_357_1258_U236, P3_SUB_357_1258_U237, P3_SUB_357_1258_U238, P3_SUB_357_1258_U239, P3_SUB_357_1258_U24, P3_SUB_357_1258_U240, P3_SUB_357_1258_U241, P3_SUB_357_1258_U242, P3_SUB_357_1258_U243, P3_SUB_357_1258_U244, P3_SUB_357_1258_U245, P3_SUB_357_1258_U246, P3_SUB_357_1258_U247, P3_SUB_357_1258_U248, P3_SUB_357_1258_U249, P3_SUB_357_1258_U25, P3_SUB_357_1258_U250, P3_SUB_357_1258_U251, P3_SUB_357_1258_U252, P3_SUB_357_1258_U253, P3_SUB_357_1258_U254, P3_SUB_357_1258_U255, P3_SUB_357_1258_U256, P3_SUB_357_1258_U257, P3_SUB_357_1258_U258, P3_SUB_357_1258_U259, P3_SUB_357_1258_U26, P3_SUB_357_1258_U260, P3_SUB_357_1258_U261, P3_SUB_357_1258_U262, P3_SUB_357_1258_U263, P3_SUB_357_1258_U264, P3_SUB_357_1258_U265, P3_SUB_357_1258_U266, P3_SUB_357_1258_U267, P3_SUB_357_1258_U268, P3_SUB_357_1258_U269, P3_SUB_357_1258_U27, P3_SUB_357_1258_U270, P3_SUB_357_1258_U271, P3_SUB_357_1258_U272, P3_SUB_357_1258_U273, P3_SUB_357_1258_U274, P3_SUB_357_1258_U275, P3_SUB_357_1258_U276, P3_SUB_357_1258_U277, P3_SUB_357_1258_U278, P3_SUB_357_1258_U279, P3_SUB_357_1258_U28, P3_SUB_357_1258_U280, P3_SUB_357_1258_U281, P3_SUB_357_1258_U282, P3_SUB_357_1258_U283, P3_SUB_357_1258_U284, P3_SUB_357_1258_U285, P3_SUB_357_1258_U286, P3_SUB_357_1258_U287, P3_SUB_357_1258_U288, P3_SUB_357_1258_U289, P3_SUB_357_1258_U29, P3_SUB_357_1258_U290, P3_SUB_357_1258_U291, P3_SUB_357_1258_U292, P3_SUB_357_1258_U293, P3_SUB_357_1258_U294, P3_SUB_357_1258_U295, P3_SUB_357_1258_U296, P3_SUB_357_1258_U297, P3_SUB_357_1258_U298, P3_SUB_357_1258_U299, P3_SUB_357_1258_U30, P3_SUB_357_1258_U300, P3_SUB_357_1258_U301, P3_SUB_357_1258_U302, P3_SUB_357_1258_U303, P3_SUB_357_1258_U304, P3_SUB_357_1258_U305, P3_SUB_357_1258_U306, P3_SUB_357_1258_U307, P3_SUB_357_1258_U308, P3_SUB_357_1258_U309, P3_SUB_357_1258_U31, P3_SUB_357_1258_U310, P3_SUB_357_1258_U311, P3_SUB_357_1258_U312, P3_SUB_357_1258_U313, P3_SUB_357_1258_U314, P3_SUB_357_1258_U315, P3_SUB_357_1258_U316, P3_SUB_357_1258_U317, P3_SUB_357_1258_U318, P3_SUB_357_1258_U319, P3_SUB_357_1258_U32, P3_SUB_357_1258_U320, P3_SUB_357_1258_U321, P3_SUB_357_1258_U322, P3_SUB_357_1258_U323, P3_SUB_357_1258_U324, P3_SUB_357_1258_U325, P3_SUB_357_1258_U326, P3_SUB_357_1258_U327, P3_SUB_357_1258_U328, P3_SUB_357_1258_U329, P3_SUB_357_1258_U33, P3_SUB_357_1258_U330, P3_SUB_357_1258_U331, P3_SUB_357_1258_U332, P3_SUB_357_1258_U333, P3_SUB_357_1258_U334, P3_SUB_357_1258_U335, P3_SUB_357_1258_U336, P3_SUB_357_1258_U337, P3_SUB_357_1258_U338, P3_SUB_357_1258_U339, P3_SUB_357_1258_U34, P3_SUB_357_1258_U340, P3_SUB_357_1258_U341, P3_SUB_357_1258_U342, P3_SUB_357_1258_U343, P3_SUB_357_1258_U344, P3_SUB_357_1258_U345, P3_SUB_357_1258_U346, P3_SUB_357_1258_U347, P3_SUB_357_1258_U348, P3_SUB_357_1258_U349, P3_SUB_357_1258_U35, P3_SUB_357_1258_U350, P3_SUB_357_1258_U351, P3_SUB_357_1258_U352, P3_SUB_357_1258_U353, P3_SUB_357_1258_U354, P3_SUB_357_1258_U355, P3_SUB_357_1258_U356, P3_SUB_357_1258_U357, P3_SUB_357_1258_U358, P3_SUB_357_1258_U359, P3_SUB_357_1258_U36, P3_SUB_357_1258_U360, P3_SUB_357_1258_U361, P3_SUB_357_1258_U362, P3_SUB_357_1258_U363, P3_SUB_357_1258_U364, P3_SUB_357_1258_U365, P3_SUB_357_1258_U366, P3_SUB_357_1258_U367, P3_SUB_357_1258_U368, P3_SUB_357_1258_U369, P3_SUB_357_1258_U37, P3_SUB_357_1258_U370, P3_SUB_357_1258_U371, P3_SUB_357_1258_U372, P3_SUB_357_1258_U373, P3_SUB_357_1258_U374, P3_SUB_357_1258_U375, P3_SUB_357_1258_U376, P3_SUB_357_1258_U377, P3_SUB_357_1258_U378, P3_SUB_357_1258_U379, P3_SUB_357_1258_U38, P3_SUB_357_1258_U380, P3_SUB_357_1258_U381, P3_SUB_357_1258_U382, P3_SUB_357_1258_U383, P3_SUB_357_1258_U384, P3_SUB_357_1258_U385, P3_SUB_357_1258_U386, P3_SUB_357_1258_U387, P3_SUB_357_1258_U388, P3_SUB_357_1258_U389, P3_SUB_357_1258_U39, P3_SUB_357_1258_U390, P3_SUB_357_1258_U391, P3_SUB_357_1258_U392, P3_SUB_357_1258_U393, P3_SUB_357_1258_U394, P3_SUB_357_1258_U395, P3_SUB_357_1258_U396, P3_SUB_357_1258_U397, P3_SUB_357_1258_U398, P3_SUB_357_1258_U399, P3_SUB_357_1258_U4, P3_SUB_357_1258_U40, P3_SUB_357_1258_U400, P3_SUB_357_1258_U401, P3_SUB_357_1258_U402, P3_SUB_357_1258_U403, P3_SUB_357_1258_U404, P3_SUB_357_1258_U405, P3_SUB_357_1258_U406, P3_SUB_357_1258_U407, P3_SUB_357_1258_U408, P3_SUB_357_1258_U409, P3_SUB_357_1258_U41, P3_SUB_357_1258_U410, P3_SUB_357_1258_U411, P3_SUB_357_1258_U412, P3_SUB_357_1258_U413, P3_SUB_357_1258_U414, P3_SUB_357_1258_U415, P3_SUB_357_1258_U416, P3_SUB_357_1258_U417, P3_SUB_357_1258_U418, P3_SUB_357_1258_U419, P3_SUB_357_1258_U42, P3_SUB_357_1258_U420, P3_SUB_357_1258_U421, P3_SUB_357_1258_U422, P3_SUB_357_1258_U423, P3_SUB_357_1258_U424, P3_SUB_357_1258_U425, P3_SUB_357_1258_U426, P3_SUB_357_1258_U427, P3_SUB_357_1258_U428, P3_SUB_357_1258_U429, P3_SUB_357_1258_U43, P3_SUB_357_1258_U430, P3_SUB_357_1258_U431, P3_SUB_357_1258_U432, P3_SUB_357_1258_U433, P3_SUB_357_1258_U434, P3_SUB_357_1258_U435, P3_SUB_357_1258_U436, P3_SUB_357_1258_U437, P3_SUB_357_1258_U438, P3_SUB_357_1258_U439, P3_SUB_357_1258_U44, P3_SUB_357_1258_U440, P3_SUB_357_1258_U441, P3_SUB_357_1258_U442, P3_SUB_357_1258_U443, P3_SUB_357_1258_U444, P3_SUB_357_1258_U445, P3_SUB_357_1258_U446, P3_SUB_357_1258_U447, P3_SUB_357_1258_U448, P3_SUB_357_1258_U449, P3_SUB_357_1258_U45, P3_SUB_357_1258_U450, P3_SUB_357_1258_U451, P3_SUB_357_1258_U452, P3_SUB_357_1258_U453, P3_SUB_357_1258_U454, P3_SUB_357_1258_U455, P3_SUB_357_1258_U456, P3_SUB_357_1258_U457, P3_SUB_357_1258_U458, P3_SUB_357_1258_U459, P3_SUB_357_1258_U46, P3_SUB_357_1258_U460, P3_SUB_357_1258_U461, P3_SUB_357_1258_U462, P3_SUB_357_1258_U463, P3_SUB_357_1258_U464, P3_SUB_357_1258_U465, P3_SUB_357_1258_U466, P3_SUB_357_1258_U467, P3_SUB_357_1258_U468, P3_SUB_357_1258_U469, P3_SUB_357_1258_U47, P3_SUB_357_1258_U470, P3_SUB_357_1258_U471, P3_SUB_357_1258_U472, P3_SUB_357_1258_U473, P3_SUB_357_1258_U474, P3_SUB_357_1258_U475, P3_SUB_357_1258_U476, P3_SUB_357_1258_U477, P3_SUB_357_1258_U478, P3_SUB_357_1258_U479, P3_SUB_357_1258_U48, P3_SUB_357_1258_U480, P3_SUB_357_1258_U481, P3_SUB_357_1258_U482, P3_SUB_357_1258_U483, P3_SUB_357_1258_U484, P3_SUB_357_1258_U49, P3_SUB_357_1258_U5, P3_SUB_357_1258_U50, P3_SUB_357_1258_U51, P3_SUB_357_1258_U52, P3_SUB_357_1258_U53, P3_SUB_357_1258_U54, P3_SUB_357_1258_U55, P3_SUB_357_1258_U56, P3_SUB_357_1258_U57, P3_SUB_357_1258_U58, P3_SUB_357_1258_U59, P3_SUB_357_1258_U6, P3_SUB_357_1258_U60, P3_SUB_357_1258_U61, P3_SUB_357_1258_U62, P3_SUB_357_1258_U63, P3_SUB_357_1258_U64, P3_SUB_357_1258_U65, P3_SUB_357_1258_U66, P3_SUB_357_1258_U67, P3_SUB_357_1258_U68, P3_SUB_357_1258_U69, P3_SUB_357_1258_U7, P3_SUB_357_1258_U70, P3_SUB_357_1258_U71, P3_SUB_357_1258_U72, P3_SUB_357_1258_U73, P3_SUB_357_1258_U74, P3_SUB_357_1258_U75, P3_SUB_357_1258_U76, P3_SUB_357_1258_U77, P3_SUB_357_1258_U78, P3_SUB_357_1258_U79, P3_SUB_357_1258_U8, P3_SUB_357_1258_U80, P3_SUB_357_1258_U81, P3_SUB_357_1258_U82, P3_SUB_357_1258_U83, P3_SUB_357_1258_U84, P3_SUB_357_1258_U85, P3_SUB_357_1258_U86, P3_SUB_357_1258_U87, P3_SUB_357_1258_U88, P3_SUB_357_1258_U89, P3_SUB_357_1258_U9, P3_SUB_357_1258_U90, P3_SUB_357_1258_U91, P3_SUB_357_1258_U92, P3_SUB_357_1258_U93, P3_SUB_357_1258_U94, P3_SUB_357_1258_U95, P3_SUB_357_1258_U96, P3_SUB_357_1258_U97, P3_SUB_357_1258_U98, P3_SUB_357_1258_U99, P3_SUB_357_U10, P3_SUB_357_U11, P3_SUB_357_U12, P3_SUB_357_U13, P3_SUB_357_U6, P3_SUB_357_U7, P3_SUB_357_U8, P3_SUB_357_U9, P3_SUB_370_U10, P3_SUB_370_U11, P3_SUB_370_U12, P3_SUB_370_U13, P3_SUB_370_U14, P3_SUB_370_U15, P3_SUB_370_U16, P3_SUB_370_U17, P3_SUB_370_U18, P3_SUB_370_U19, P3_SUB_370_U20, P3_SUB_370_U21, P3_SUB_370_U22, P3_SUB_370_U23, P3_SUB_370_U24, P3_SUB_370_U25, P3_SUB_370_U26, P3_SUB_370_U27, P3_SUB_370_U28, P3_SUB_370_U29, P3_SUB_370_U30, P3_SUB_370_U31, P3_SUB_370_U32, P3_SUB_370_U33, P3_SUB_370_U34, P3_SUB_370_U35, P3_SUB_370_U36, P3_SUB_370_U37, P3_SUB_370_U38, P3_SUB_370_U39, P3_SUB_370_U40, P3_SUB_370_U41, P3_SUB_370_U42, P3_SUB_370_U43, P3_SUB_370_U44, P3_SUB_370_U45, P3_SUB_370_U46, P3_SUB_370_U47, P3_SUB_370_U48, P3_SUB_370_U49, P3_SUB_370_U50, P3_SUB_370_U51, P3_SUB_370_U52, P3_SUB_370_U53, P3_SUB_370_U54, P3_SUB_370_U55, P3_SUB_370_U56, P3_SUB_370_U57, P3_SUB_370_U58, P3_SUB_370_U59, P3_SUB_370_U6, P3_SUB_370_U60, P3_SUB_370_U61, P3_SUB_370_U62, P3_SUB_370_U63, P3_SUB_370_U64, P3_SUB_370_U65, P3_SUB_370_U66, P3_SUB_370_U7, P3_SUB_370_U8, P3_SUB_370_U9, P3_SUB_390_U10, P3_SUB_390_U11, P3_SUB_390_U12, P3_SUB_390_U13, P3_SUB_390_U14, P3_SUB_390_U15, P3_SUB_390_U16, P3_SUB_390_U17, P3_SUB_390_U18, P3_SUB_390_U19, P3_SUB_390_U20, P3_SUB_390_U21, P3_SUB_390_U22, P3_SUB_390_U23, P3_SUB_390_U24, P3_SUB_390_U25, P3_SUB_390_U26, P3_SUB_390_U27, P3_SUB_390_U28, P3_SUB_390_U29, P3_SUB_390_U30, P3_SUB_390_U31, P3_SUB_390_U32, P3_SUB_390_U33, P3_SUB_390_U34, P3_SUB_390_U35, P3_SUB_390_U36, P3_SUB_390_U37, P3_SUB_390_U38, P3_SUB_390_U39, P3_SUB_390_U40, P3_SUB_390_U41, P3_SUB_390_U42, P3_SUB_390_U43, P3_SUB_390_U44, P3_SUB_390_U45, P3_SUB_390_U46, P3_SUB_390_U47, P3_SUB_390_U48, P3_SUB_390_U49, P3_SUB_390_U50, P3_SUB_390_U51, P3_SUB_390_U52, P3_SUB_390_U53, P3_SUB_390_U54, P3_SUB_390_U55, P3_SUB_390_U56, P3_SUB_390_U57, P3_SUB_390_U58, P3_SUB_390_U59, P3_SUB_390_U6, P3_SUB_390_U60, P3_SUB_390_U61, P3_SUB_390_U62, P3_SUB_390_U63, P3_SUB_390_U64, P3_SUB_390_U65, P3_SUB_390_U66, P3_SUB_390_U7, P3_SUB_390_U8, P3_SUB_390_U9, P3_SUB_401_U10, P3_SUB_401_U11, P3_SUB_401_U12, P3_SUB_401_U13, P3_SUB_401_U14, P3_SUB_401_U15, P3_SUB_401_U16, P3_SUB_401_U17, P3_SUB_401_U18, P3_SUB_401_U19, P3_SUB_401_U20, P3_SUB_401_U21, P3_SUB_401_U22, P3_SUB_401_U23, P3_SUB_401_U24, P3_SUB_401_U25, P3_SUB_401_U26, P3_SUB_401_U27, P3_SUB_401_U28, P3_SUB_401_U29, P3_SUB_401_U30, P3_SUB_401_U31, P3_SUB_401_U32, P3_SUB_401_U33, P3_SUB_401_U34, P3_SUB_401_U35, P3_SUB_401_U36, P3_SUB_401_U37, P3_SUB_401_U38, P3_SUB_401_U39, P3_SUB_401_U40, P3_SUB_401_U41, P3_SUB_401_U42, P3_SUB_401_U43, P3_SUB_401_U44, P3_SUB_401_U45, P3_SUB_401_U46, P3_SUB_401_U47, P3_SUB_401_U48, P3_SUB_401_U49, P3_SUB_401_U50, P3_SUB_401_U51, P3_SUB_401_U52, P3_SUB_401_U53, P3_SUB_401_U54, P3_SUB_401_U55, P3_SUB_401_U56, P3_SUB_401_U57, P3_SUB_401_U58, P3_SUB_401_U59, P3_SUB_401_U6, P3_SUB_401_U60, P3_SUB_401_U61, P3_SUB_401_U62, P3_SUB_401_U63, P3_SUB_401_U64, P3_SUB_401_U65, P3_SUB_401_U66, P3_SUB_401_U7, P3_SUB_401_U8, P3_SUB_401_U9, P3_SUB_412_U10, P3_SUB_412_U11, P3_SUB_412_U12, P3_SUB_412_U13, P3_SUB_412_U14, P3_SUB_412_U15, P3_SUB_412_U16, P3_SUB_412_U17, P3_SUB_412_U18, P3_SUB_412_U19, P3_SUB_412_U20, P3_SUB_412_U21, P3_SUB_412_U22, P3_SUB_412_U23, P3_SUB_412_U24, P3_SUB_412_U25, P3_SUB_412_U26, P3_SUB_412_U27, P3_SUB_412_U28, P3_SUB_412_U29, P3_SUB_412_U30, P3_SUB_412_U31, P3_SUB_412_U32, P3_SUB_412_U33, P3_SUB_412_U34, P3_SUB_412_U35, P3_SUB_412_U36, P3_SUB_412_U37, P3_SUB_412_U38, P3_SUB_412_U39, P3_SUB_412_U40, P3_SUB_412_U41, P3_SUB_412_U42, P3_SUB_412_U43, P3_SUB_412_U44, P3_SUB_412_U45, P3_SUB_412_U46, P3_SUB_412_U47, P3_SUB_412_U48, P3_SUB_412_U49, P3_SUB_412_U50, P3_SUB_412_U51, P3_SUB_412_U52, P3_SUB_412_U53, P3_SUB_412_U54, P3_SUB_412_U55, P3_SUB_412_U56, P3_SUB_412_U57, P3_SUB_412_U58, P3_SUB_412_U59, P3_SUB_412_U6, P3_SUB_412_U60, P3_SUB_412_U61, P3_SUB_412_U62, P3_SUB_412_U63, P3_SUB_412_U7, P3_SUB_412_U8, P3_SUB_412_U9, P3_SUB_414_U10, P3_SUB_414_U100, P3_SUB_414_U101, P3_SUB_414_U102, P3_SUB_414_U103, P3_SUB_414_U104, P3_SUB_414_U105, P3_SUB_414_U106, P3_SUB_414_U107, P3_SUB_414_U108, P3_SUB_414_U109, P3_SUB_414_U11, P3_SUB_414_U110, P3_SUB_414_U111, P3_SUB_414_U112, P3_SUB_414_U113, P3_SUB_414_U114, P3_SUB_414_U115, P3_SUB_414_U116, P3_SUB_414_U117, P3_SUB_414_U118, P3_SUB_414_U119, P3_SUB_414_U12, P3_SUB_414_U120, P3_SUB_414_U121, P3_SUB_414_U122, P3_SUB_414_U123, P3_SUB_414_U124, P3_SUB_414_U125, P3_SUB_414_U126, P3_SUB_414_U127, P3_SUB_414_U128, P3_SUB_414_U129, P3_SUB_414_U13, P3_SUB_414_U130, P3_SUB_414_U131, P3_SUB_414_U132, P3_SUB_414_U133, P3_SUB_414_U134, P3_SUB_414_U135, P3_SUB_414_U136, P3_SUB_414_U137, P3_SUB_414_U138, P3_SUB_414_U139, P3_SUB_414_U14, P3_SUB_414_U140, P3_SUB_414_U141, P3_SUB_414_U142, P3_SUB_414_U143, P3_SUB_414_U144, P3_SUB_414_U145, P3_SUB_414_U146, P3_SUB_414_U147, P3_SUB_414_U148, P3_SUB_414_U149, P3_SUB_414_U15, P3_SUB_414_U150, P3_SUB_414_U151, P3_SUB_414_U152, P3_SUB_414_U153, P3_SUB_414_U154, P3_SUB_414_U155, P3_SUB_414_U156, P3_SUB_414_U157, P3_SUB_414_U158, P3_SUB_414_U159, P3_SUB_414_U16, P3_SUB_414_U17, P3_SUB_414_U18, P3_SUB_414_U19, P3_SUB_414_U20, P3_SUB_414_U21, P3_SUB_414_U22, P3_SUB_414_U23, P3_SUB_414_U24, P3_SUB_414_U25, P3_SUB_414_U26, P3_SUB_414_U27, P3_SUB_414_U28, P3_SUB_414_U29, P3_SUB_414_U30, P3_SUB_414_U31, P3_SUB_414_U32, P3_SUB_414_U33, P3_SUB_414_U34, P3_SUB_414_U35, P3_SUB_414_U36, P3_SUB_414_U37, P3_SUB_414_U38, P3_SUB_414_U39, P3_SUB_414_U40, P3_SUB_414_U41, P3_SUB_414_U42, P3_SUB_414_U43, P3_SUB_414_U44, P3_SUB_414_U45, P3_SUB_414_U46, P3_SUB_414_U47, P3_SUB_414_U48, P3_SUB_414_U49, P3_SUB_414_U50, P3_SUB_414_U51, P3_SUB_414_U52, P3_SUB_414_U53, P3_SUB_414_U54, P3_SUB_414_U55, P3_SUB_414_U56, P3_SUB_414_U57, P3_SUB_414_U58, P3_SUB_414_U59, P3_SUB_414_U6, P3_SUB_414_U60, P3_SUB_414_U61, P3_SUB_414_U62, P3_SUB_414_U63, P3_SUB_414_U64, P3_SUB_414_U65, P3_SUB_414_U66, P3_SUB_414_U67, P3_SUB_414_U68, P3_SUB_414_U69, P3_SUB_414_U7, P3_SUB_414_U70, P3_SUB_414_U71, P3_SUB_414_U72, P3_SUB_414_U73, P3_SUB_414_U74, P3_SUB_414_U75, P3_SUB_414_U76, P3_SUB_414_U77, P3_SUB_414_U78, P3_SUB_414_U79, P3_SUB_414_U8, P3_SUB_414_U80, P3_SUB_414_U81, P3_SUB_414_U82, P3_SUB_414_U83, P3_SUB_414_U84, P3_SUB_414_U85, P3_SUB_414_U86, P3_SUB_414_U87, P3_SUB_414_U88, P3_SUB_414_U89, P3_SUB_414_U9, P3_SUB_414_U90, P3_SUB_414_U91, P3_SUB_414_U92, P3_SUB_414_U93, P3_SUB_414_U94, P3_SUB_414_U95, P3_SUB_414_U96, P3_SUB_414_U97, P3_SUB_414_U98, P3_SUB_414_U99, P3_SUB_450_U10, P3_SUB_450_U11, P3_SUB_450_U12, P3_SUB_450_U13, P3_SUB_450_U14, P3_SUB_450_U15, P3_SUB_450_U16, P3_SUB_450_U17, P3_SUB_450_U18, P3_SUB_450_U19, P3_SUB_450_U20, P3_SUB_450_U21, P3_SUB_450_U22, P3_SUB_450_U23, P3_SUB_450_U24, P3_SUB_450_U25, P3_SUB_450_U26, P3_SUB_450_U27, P3_SUB_450_U28, P3_SUB_450_U29, P3_SUB_450_U30, P3_SUB_450_U31, P3_SUB_450_U32, P3_SUB_450_U33, P3_SUB_450_U34, P3_SUB_450_U35, P3_SUB_450_U36, P3_SUB_450_U37, P3_SUB_450_U38, P3_SUB_450_U39, P3_SUB_450_U40, P3_SUB_450_U41, P3_SUB_450_U42, P3_SUB_450_U43, P3_SUB_450_U44, P3_SUB_450_U45, P3_SUB_450_U46, P3_SUB_450_U47, P3_SUB_450_U48, P3_SUB_450_U49, P3_SUB_450_U50, P3_SUB_450_U51, P3_SUB_450_U52, P3_SUB_450_U53, P3_SUB_450_U54, P3_SUB_450_U55, P3_SUB_450_U56, P3_SUB_450_U57, P3_SUB_450_U58, P3_SUB_450_U59, P3_SUB_450_U6, P3_SUB_450_U60, P3_SUB_450_U61, P3_SUB_450_U62, P3_SUB_450_U63, P3_SUB_450_U7, P3_SUB_450_U8, P3_SUB_450_U9, P3_SUB_485_U10, P3_SUB_485_U11, P3_SUB_485_U12, P3_SUB_485_U13, P3_SUB_485_U14, P3_SUB_485_U15, P3_SUB_485_U16, P3_SUB_485_U17, P3_SUB_485_U18, P3_SUB_485_U19, P3_SUB_485_U20, P3_SUB_485_U21, P3_SUB_485_U22, P3_SUB_485_U23, P3_SUB_485_U24, P3_SUB_485_U25, P3_SUB_485_U26, P3_SUB_485_U27, P3_SUB_485_U28, P3_SUB_485_U29, P3_SUB_485_U30, P3_SUB_485_U31, P3_SUB_485_U32, P3_SUB_485_U33, P3_SUB_485_U34, P3_SUB_485_U35, P3_SUB_485_U36, P3_SUB_485_U37, P3_SUB_485_U38, P3_SUB_485_U39, P3_SUB_485_U40, P3_SUB_485_U41, P3_SUB_485_U42, P3_SUB_485_U43, P3_SUB_485_U44, P3_SUB_485_U45, P3_SUB_485_U46, P3_SUB_485_U47, P3_SUB_485_U48, P3_SUB_485_U49, P3_SUB_485_U50, P3_SUB_485_U51, P3_SUB_485_U52, P3_SUB_485_U53, P3_SUB_485_U54, P3_SUB_485_U55, P3_SUB_485_U56, P3_SUB_485_U57, P3_SUB_485_U58, P3_SUB_485_U59, P3_SUB_485_U6, P3_SUB_485_U60, P3_SUB_485_U61, P3_SUB_485_U62, P3_SUB_485_U63, P3_SUB_485_U7, P3_SUB_485_U8, P3_SUB_485_U9, P3_SUB_504_U10, P3_SUB_504_U11, P3_SUB_504_U12, P3_SUB_504_U13, P3_SUB_504_U14, P3_SUB_504_U15, P3_SUB_504_U16, P3_SUB_504_U17, P3_SUB_504_U18, P3_SUB_504_U19, P3_SUB_504_U20, P3_SUB_504_U21, P3_SUB_504_U22, P3_SUB_504_U23, P3_SUB_504_U24, P3_SUB_504_U25, P3_SUB_504_U26, P3_SUB_504_U27, P3_SUB_504_U28, P3_SUB_504_U29, P3_SUB_504_U30, P3_SUB_504_U31, P3_SUB_504_U32, P3_SUB_504_U33, P3_SUB_504_U34, P3_SUB_504_U35, P3_SUB_504_U36, P3_SUB_504_U37, P3_SUB_504_U38, P3_SUB_504_U39, P3_SUB_504_U40, P3_SUB_504_U41, P3_SUB_504_U42, P3_SUB_504_U43, P3_SUB_504_U44, P3_SUB_504_U45, P3_SUB_504_U46, P3_SUB_504_U47, P3_SUB_504_U48, P3_SUB_504_U49, P3_SUB_504_U50, P3_SUB_504_U51, P3_SUB_504_U52, P3_SUB_504_U53, P3_SUB_504_U54, P3_SUB_504_U55, P3_SUB_504_U56, P3_SUB_504_U57, P3_SUB_504_U58, P3_SUB_504_U59, P3_SUB_504_U6, P3_SUB_504_U60, P3_SUB_504_U61, P3_SUB_504_U62, P3_SUB_504_U63, P3_SUB_504_U7, P3_SUB_504_U8, P3_SUB_504_U9, P3_SUB_563_U6, P3_SUB_563_U7, P3_SUB_580_U10, P3_SUB_580_U6, P3_SUB_580_U7, P3_SUB_580_U8, P3_SUB_580_U9, P3_SUB_589_U6, P3_SUB_589_U7, P3_SUB_589_U8, P3_SUB_589_U9, P3_U2352, P3_U2353, P3_U2354, P3_U2355, P3_U2356, P3_U2357, P3_U2358, P3_U2359, P3_U2360, P3_U2361, P3_U2362, P3_U2363, P3_U2364, P3_U2365, P3_U2366, P3_U2367, P3_U2368, P3_U2369, P3_U2370, P3_U2371, P3_U2372, P3_U2373, P3_U2374, P3_U2375, P3_U2376, P3_U2377, P3_U2378, P3_U2379, P3_U2380, P3_U2381, P3_U2382, P3_U2383, P3_U2384, P3_U2385, P3_U2386, P3_U2387, P3_U2388, P3_U2389, P3_U2390, P3_U2391, P3_U2392, P3_U2393, P3_U2394, P3_U2395, P3_U2396, P3_U2397, P3_U2398, P3_U2399, P3_U2400, P3_U2401, P3_U2402, P3_U2403, P3_U2404, P3_U2405, P3_U2406, P3_U2407, P3_U2408, P3_U2409, P3_U2410, P3_U2411, P3_U2412, P3_U2413, P3_U2414, P3_U2415, P3_U2416, P3_U2417, P3_U2418, P3_U2419, P3_U2420, P3_U2421, P3_U2422, P3_U2423, P3_U2424, P3_U2425, P3_U2426, P3_U2427, P3_U2428, P3_U2429, P3_U2430, P3_U2431, P3_U2432, P3_U2433, P3_U2434, P3_U2435, P3_U2436, P3_U2437, P3_U2438, P3_U2439, P3_U2440, P3_U2441, P3_U2442, P3_U2443, P3_U2444, P3_U2445, P3_U2446, P3_U2447, P3_U2448, P3_U2449, P3_U2450, P3_U2451, P3_U2452, P3_U2453, P3_U2454, P3_U2455, P3_U2456, P3_U2457, P3_U2458, P3_U2459, P3_U2460, P3_U2461, P3_U2462, P3_U2463, P3_U2464, P3_U2465, P3_U2466, P3_U2467, P3_U2468, P3_U2469, P3_U2470, P3_U2471, P3_U2472, P3_U2473, P3_U2474, P3_U2475, P3_U2476, P3_U2477, P3_U2478, P3_U2479, P3_U2480, P3_U2481, P3_U2482, P3_U2483, P3_U2484, P3_U2485, P3_U2486, P3_U2487, P3_U2488, P3_U2489, P3_U2490, P3_U2491, P3_U2492, P3_U2493, P3_U2494, P3_U2495, P3_U2496, P3_U2497, P3_U2498, P3_U2499, P3_U2500, P3_U2501, P3_U2502, P3_U2503, P3_U2504, P3_U2505, P3_U2506, P3_U2507, P3_U2508, P3_U2509, P3_U2510, P3_U2511, P3_U2512, P3_U2513, P3_U2514, P3_U2515, P3_U2516, P3_U2517, P3_U2518, P3_U2519, P3_U2520, P3_U2521, P3_U2522, P3_U2523, P3_U2524, P3_U2525, P3_U2526, P3_U2527, P3_U2528, P3_U2529, P3_U2530, P3_U2531, P3_U2532, P3_U2533, P3_U2534, P3_U2535, P3_U2536, P3_U2537, P3_U2538, P3_U2539, P3_U2540, P3_U2541, P3_U2542, P3_U2543, P3_U2544, P3_U2545, P3_U2546, P3_U2547, P3_U2548, P3_U2549, P3_U2550, P3_U2551, P3_U2552, P3_U2553, P3_U2554, P3_U2555, P3_U2556, P3_U2557, P3_U2558, P3_U2559, P3_U2560, P3_U2561, P3_U2562, P3_U2563, P3_U2564, P3_U2565, P3_U2566, P3_U2567, P3_U2568, P3_U2569, P3_U2570, P3_U2571, P3_U2572, P3_U2573, P3_U2574, P3_U2575, P3_U2576, P3_U2577, P3_U2578, P3_U2579, P3_U2580, P3_U2581, P3_U2582, P3_U2583, P3_U2584, P3_U2585, P3_U2586, P3_U2587, P3_U2588, P3_U2589, P3_U2590, P3_U2591, P3_U2592, P3_U2593, P3_U2594, P3_U2595, P3_U2596, P3_U2597, P3_U2598, P3_U2599, P3_U2600, P3_U2601, P3_U2602, P3_U2603, P3_U2604, P3_U2605, P3_U2606, P3_U2607, P3_U2608, P3_U2609, P3_U2610, P3_U2611, P3_U2612, P3_U2613, P3_U2614, P3_U2615, P3_U2616, P3_U2617, P3_U2618, P3_U2619, P3_U2620, P3_U2621, P3_U2622, P3_U2623, P3_U2624, P3_U2625, P3_U2626, P3_U2627, P3_U2628, P3_U2629, P3_U2630, P3_U2631, P3_U2632, P3_U3062, P3_U3063, P3_U3064, P3_U3065, P3_U3066, P3_U3067, P3_U3068, P3_U3069, P3_U3070, P3_U3071, P3_U3072, P3_U3073, P3_U3074, P3_U3075, P3_U3076, P3_U3077, P3_U3078, P3_U3079, P3_U3080, P3_U3081, P3_U3082, P3_U3083, P3_U3084, P3_U3085, P3_U3086, P3_U3087, P3_U3088, P3_U3089, P3_U3090, P3_U3091, P3_U3092, P3_U3093, P3_U3094, P3_U3095, P3_U3096, P3_U3097, P3_U3098, P3_U3099, P3_U3100, P3_U3101, P3_U3102, P3_U3103, P3_U3104, P3_U3105, P3_U3106, P3_U3107, P3_U3108, P3_U3109, P3_U3110, P3_U3111, P3_U3112, P3_U3113, P3_U3114, P3_U3115, P3_U3116, P3_U3117, P3_U3118, P3_U3119, P3_U3120, P3_U3121, P3_U3122, P3_U3123, P3_U3124, P3_U3125, P3_U3126, P3_U3127, P3_U3128, P3_U3129, P3_U3130, P3_U3131, P3_U3132, P3_U3133, P3_U3134, P3_U3135, P3_U3136, P3_U3137, P3_U3138, P3_U3139, P3_U3140, P3_U3141, P3_U3142, P3_U3143, P3_U3144, P3_U3145, P3_U3146, P3_U3147, P3_U3148, P3_U3149, P3_U3150, P3_U3151, P3_U3152, P3_U3153, P3_U3154, P3_U3155, P3_U3156, P3_U3157, P3_U3158, P3_U3159, P3_U3160, P3_U3161, P3_U3162, P3_U3163, P3_U3164, P3_U3165, P3_U3166, P3_U3167, P3_U3168, P3_U3169, P3_U3170, P3_U3171, P3_U3172, P3_U3173, P3_U3174, P3_U3175, P3_U3176, P3_U3177, P3_U3178, P3_U3179, P3_U3180, P3_U3181, P3_U3182, P3_U3183, P3_U3184, P3_U3185, P3_U3186, P3_U3187, P3_U3188, P3_U3189, P3_U3190, P3_U3191, P3_U3192, P3_U3193, P3_U3194, P3_U3195, P3_U3196, P3_U3197, P3_U3198, P3_U3199, P3_U3200, P3_U3201, P3_U3202, P3_U3203, P3_U3204, P3_U3205, P3_U3206, P3_U3207, P3_U3208, P3_U3209, P3_U3210, P3_U3211, P3_U3212, P3_U3213, P3_U3214, P3_U3215, P3_U3216, P3_U3217, P3_U3218, P3_U3219, P3_U3220, P3_U3221, P3_U3222, P3_U3223, P3_U3224, P3_U3225, P3_U3226, P3_U3227, P3_U3228, P3_U3229, P3_U3230, P3_U3231, P3_U3232, P3_U3233, P3_U3234, P3_U3235, P3_U3236, P3_U3237, P3_U3238, P3_U3239, P3_U3240, P3_U3241, P3_U3242, P3_U3243, P3_U3244, P3_U3245, P3_U3246, P3_U3247, P3_U3248, P3_U3249, P3_U3250, P3_U3251, P3_U3252, P3_U3253, P3_U3254, P3_U3255, P3_U3256, P3_U3257, P3_U3258, P3_U3259, P3_U3260, P3_U3261, P3_U3262, P3_U3263, P3_U3264, P3_U3265, P3_U3266, P3_U3267, P3_U3268, P3_U3269, P3_U3270, P3_U3271, P3_U3272, P3_U3273, P3_U3278, P3_U3279, P3_U3283, P3_U3286, P3_U3287, P3_U3291, P3_U3300, P3_U3301, P3_U3302, P3_U3303, P3_U3304, P3_U3305, P3_U3306, P3_U3307, P3_U3308, P3_U3309, P3_U3310, P3_U3311, P3_U3312, P3_U3313, P3_U3314, P3_U3315, P3_U3316, P3_U3317, P3_U3318, P3_U3319, P3_U3320, P3_U3321, P3_U3322, P3_U3323, P3_U3324, P3_U3325, P3_U3326, P3_U3327, P3_U3328, P3_U3329, P3_U3330, P3_U3331, P3_U3332, P3_U3333, P3_U3334, P3_U3335, P3_U3336, P3_U3337, P3_U3338, P3_U3339, P3_U3340, P3_U3341, P3_U3342, P3_U3343, P3_U3344, P3_U3345, P3_U3346, P3_U3347, P3_U3348, P3_U3349, P3_U3350, P3_U3351, P3_U3352, P3_U3353, P3_U3354, P3_U3355, P3_U3356, P3_U3357, P3_U3358, P3_U3359, P3_U3360, P3_U3361, P3_U3362, P3_U3363, P3_U3364, P3_U3365, P3_U3366, P3_U3367, P3_U3368, P3_U3369, P3_U3370, P3_U3371, P3_U3372, P3_U3373, P3_U3374, P3_U3375, P3_U3376, P3_U3377, P3_U3378, P3_U3379, P3_U3380, P3_U3381, P3_U3382, P3_U3383, P3_U3384, P3_U3385, P3_U3386, P3_U3387, P3_U3388, P3_U3389, P3_U3390, P3_U3391, P3_U3392, P3_U3393, P3_U3394, P3_U3395, P3_U3396, P3_U3397, P3_U3398, P3_U3399, P3_U3400, P3_U3401, P3_U3402, P3_U3403, P3_U3404, P3_U3405, P3_U3406, P3_U3407, P3_U3408, P3_U3409, P3_U3410, P3_U3411, P3_U3412, P3_U3413, P3_U3414, P3_U3415, P3_U3416, P3_U3417, P3_U3418, P3_U3419, P3_U3420, P3_U3421, P3_U3422, P3_U3423, P3_U3424, P3_U3425, P3_U3426, P3_U3427, P3_U3428, P3_U3429, P3_U3430, P3_U3431, P3_U3432, P3_U3433, P3_U3434, P3_U3435, P3_U3436, P3_U3437, P3_U3438, P3_U3439, P3_U3440, P3_U3441, P3_U3442, P3_U3443, P3_U3444, P3_U3445, P3_U3446, P3_U3447, P3_U3448, P3_U3449, P3_U3450, P3_U3451, P3_U3452, P3_U3453, P3_U3454, P3_U3455, P3_U3456, P3_U3457, P3_U3458, P3_U3459, P3_U3460, P3_U3461, P3_U3462, P3_U3463, P3_U3464, P3_U3465, P3_U3466, P3_U3467, P3_U3468, P3_U3469, P3_U3470, P3_U3471, P3_U3472, P3_U3473, P3_U3474, P3_U3475, P3_U3476, P3_U3477, P3_U3478, P3_U3479, P3_U3480, P3_U3481, P3_U3482, P3_U3483, P3_U3484, P3_U3485, P3_U3486, P3_U3487, P3_U3488, P3_U3489, P3_U3490, P3_U3491, P3_U3492, P3_U3493, P3_U3494, P3_U3495, P3_U3496, P3_U3497, P3_U3498, P3_U3499, P3_U3500, P3_U3501, P3_U3502, P3_U3503, P3_U3504, P3_U3505, P3_U3506, P3_U3507, P3_U3508, P3_U3509, P3_U3510, P3_U3511, P3_U3512, P3_U3513, P3_U3514, P3_U3515, P3_U3516, P3_U3517, P3_U3518, P3_U3519, P3_U3520, P3_U3521, P3_U3522, P3_U3523, P3_U3524, P3_U3525, P3_U3526, P3_U3527, P3_U3528, P3_U3529, P3_U3530, P3_U3531, P3_U3532, P3_U3533, P3_U3534, P3_U3535, P3_U3536, P3_U3537, P3_U3538, P3_U3539, P3_U3540, P3_U3541, P3_U3542, P3_U3543, P3_U3544, P3_U3545, P3_U3546, P3_U3547, P3_U3548, P3_U3549, P3_U3550, P3_U3551, P3_U3552, P3_U3553, P3_U3554, P3_U3555, P3_U3556, P3_U3557, P3_U3558, P3_U3559, P3_U3560, P3_U3561, P3_U3562, P3_U3563, P3_U3564, P3_U3565, P3_U3566, P3_U3567, P3_U3568, P3_U3569, P3_U3570, P3_U3571, P3_U3572, P3_U3573, P3_U3574, P3_U3575, P3_U3576, P3_U3577, P3_U3578, P3_U3579, P3_U3580, P3_U3581, P3_U3582, P3_U3583, P3_U3584, P3_U3585, P3_U3586, P3_U3587, P3_U3588, P3_U3589, P3_U3590, P3_U3591, P3_U3592, P3_U3593, P3_U3594, P3_U3595, P3_U3596, P3_U3597, P3_U3598, P3_U3599, P3_U3600, P3_U3601, P3_U3602, P3_U3603, P3_U3604, P3_U3605, P3_U3606, P3_U3607, P3_U3608, P3_U3609, P3_U3610, P3_U3611, P3_U3612, P3_U3613, P3_U3614, P3_U3615, P3_U3616, P3_U3617, P3_U3618, P3_U3619, P3_U3620, P3_U3621, P3_U3622, P3_U3623, P3_U3624, P3_U3625, P3_U3626, P3_U3627, P3_U3628, P3_U3629, P3_U3630, P3_U3631, P3_U3632, P3_U3633, P3_U3634, P3_U3635, P3_U3636, P3_U3637, P3_U3638, P3_U3639, P3_U3640, P3_U3641, P3_U3642, P3_U3643, P3_U3644, P3_U3645, P3_U3646, P3_U3647, P3_U3648, P3_U3649, P3_U3650, P3_U3651, P3_U3652, P3_U3653, P3_U3654, P3_U3655, P3_U3656, P3_U3657, P3_U3658, P3_U3659, P3_U3660, P3_U3661, P3_U3662, P3_U3663, P3_U3664, P3_U3665, P3_U3666, P3_U3667, P3_U3668, P3_U3669, P3_U3670, P3_U3671, P3_U3672, P3_U3673, P3_U3674, P3_U3675, P3_U3676, P3_U3677, P3_U3678, P3_U3679, P3_U3680, P3_U3681, P3_U3682, P3_U3683, P3_U3684, P3_U3685, P3_U3686, P3_U3687, P3_U3688, P3_U3689, P3_U3690, P3_U3691, P3_U3692, P3_U3693, P3_U3694, P3_U3695, P3_U3696, P3_U3697, P3_U3698, P3_U3699, P3_U3700, P3_U3701, P3_U3702, P3_U3703, P3_U3704, P3_U3705, P3_U3706, P3_U3707, P3_U3708, P3_U3709, P3_U3710, P3_U3711, P3_U3712, P3_U3713, P3_U3714, P3_U3715, P3_U3716, P3_U3717, P3_U3718, P3_U3719, P3_U3720, P3_U3721, P3_U3722, P3_U3723, P3_U3724, P3_U3725, P3_U3726, P3_U3727, P3_U3728, P3_U3729, P3_U3730, P3_U3731, P3_U3732, P3_U3733, P3_U3734, P3_U3735, P3_U3736, P3_U3737, P3_U3738, P3_U3739, P3_U3740, P3_U3741, P3_U3742, P3_U3743, P3_U3744, P3_U3745, P3_U3746, P3_U3747, P3_U3748, P3_U3749, P3_U3750, P3_U3751, P3_U3752, P3_U3753, P3_U3754, P3_U3755, P3_U3756, P3_U3757, P3_U3758, P3_U3759, P3_U3760, P3_U3761, P3_U3762, P3_U3763, P3_U3764, P3_U3765, P3_U3766, P3_U3767, P3_U3768, P3_U3769, P3_U3770, P3_U3771, P3_U3772, P3_U3773, P3_U3774, P3_U3775, P3_U3776, P3_U3777, P3_U3778, P3_U3779, P3_U3780, P3_U3781, P3_U3782, P3_U3783, P3_U3784, P3_U3785, P3_U3786, P3_U3787, P3_U3788, P3_U3789, P3_U3790, P3_U3791, P3_U3792, P3_U3793, P3_U3794, P3_U3795, P3_U3796, P3_U3797, P3_U3798, P3_U3799, P3_U3800, P3_U3801, P3_U3802, P3_U3803, P3_U3804, P3_U3805, P3_U3806, P3_U3807, P3_U3808, P3_U3809, P3_U3810, P3_U3811, P3_U3812, P3_U3813, P3_U3814, P3_U3815, P3_U3816, P3_U3817, P3_U3818, P3_U3819, P3_U3820, P3_U3821, P3_U3822, P3_U3823, P3_U3824, P3_U3825, P3_U3826, P3_U3827, P3_U3828, P3_U3829, P3_U3830, P3_U3831, P3_U3832, P3_U3833, P3_U3834, P3_U3835, P3_U3836, P3_U3837, P3_U3838, P3_U3839, P3_U3840, P3_U3841, P3_U3842, P3_U3843, P3_U3844, P3_U3845, P3_U3846, P3_U3847, P3_U3848, P3_U3849, P3_U3850, P3_U3851, P3_U3852, P3_U3853, P3_U3854, P3_U3855, P3_U3856, P3_U3857, P3_U3858, P3_U3859, P3_U3860, P3_U3861, P3_U3862, P3_U3863, P3_U3864, P3_U3865, P3_U3866, P3_U3867, P3_U3868, P3_U3869, P3_U3870, P3_U3871, P3_U3872, P3_U3873, P3_U3874, P3_U3875, P3_U3876, P3_U3877, P3_U3878, P3_U3879, P3_U3880, P3_U3881, P3_U3882, P3_U3883, P3_U3884, P3_U3885, P3_U3886, P3_U3887, P3_U3888, P3_U3889, P3_U3890, P3_U3891, P3_U3892, P3_U3893, P3_U3894, P3_U3895, P3_U3896, P3_U3897, P3_U3898, P3_U3899, P3_U3900, P3_U3901, P3_U3902, P3_U3903, P3_U3904, P3_U3905, P3_U3906, P3_U3907, P3_U3908, P3_U3909, P3_U3910, P3_U3911, P3_U3912, P3_U3913, P3_U3914, P3_U3915, P3_U3916, P3_U3917, P3_U3918, P3_U3919, P3_U3920, P3_U3921, P3_U3922, P3_U3923, P3_U3924, P3_U3925, P3_U3926, P3_U3927, P3_U3928, P3_U3929, P3_U3930, P3_U3931, P3_U3932, P3_U3933, P3_U3934, P3_U3935, P3_U3936, P3_U3937, P3_U3938, P3_U3939, P3_U3940, P3_U3941, P3_U3942, P3_U3943, P3_U3944, P3_U3945, P3_U3946, P3_U3947, P3_U3948, P3_U3949, P3_U3950, P3_U3951, P3_U3952, P3_U3953, P3_U3954, P3_U3955, P3_U3956, P3_U3957, P3_U3958, P3_U3959, P3_U3960, P3_U3961, P3_U3962, P3_U3963, P3_U3964, P3_U3965, P3_U3966, P3_U3967, P3_U3968, P3_U3969, P3_U3970, P3_U3971, P3_U3972, P3_U3973, P3_U3974, P3_U3975, P3_U3976, P3_U3977, P3_U3978, P3_U3979, P3_U3980, P3_U3981, P3_U3982, P3_U3983, P3_U3984, P3_U3985, P3_U3986, P3_U3987, P3_U3988, P3_U3989, P3_U3990, P3_U3991, P3_U3992, P3_U3993, P3_U3994, P3_U3995, P3_U3996, P3_U3997, P3_U3998, P3_U3999, P3_U4000, P3_U4001, P3_U4002, P3_U4003, P3_U4004, P3_U4005, P3_U4006, P3_U4007, P3_U4008, P3_U4009, P3_U4010, P3_U4011, P3_U4012, P3_U4013, P3_U4014, P3_U4015, P3_U4016, P3_U4017, P3_U4018, P3_U4019, P3_U4020, P3_U4021, P3_U4022, P3_U4023, P3_U4024, P3_U4025, P3_U4026, P3_U4027, P3_U4028, P3_U4029, P3_U4030, P3_U4031, P3_U4032, P3_U4033, P3_U4034, P3_U4035, P3_U4036, P3_U4037, P3_U4038, P3_U4039, P3_U4040, P3_U4041, P3_U4042, P3_U4043, P3_U4044, P3_U4045, P3_U4046, P3_U4047, P3_U4048, P3_U4049, P3_U4050, P3_U4051, P3_U4052, P3_U4053, P3_U4054, P3_U4055, P3_U4056, P3_U4057, P3_U4058, P3_U4059, P3_U4060, P3_U4061, P3_U4062, P3_U4063, P3_U4064, P3_U4065, P3_U4066, P3_U4067, P3_U4068, P3_U4069, P3_U4070, P3_U4071, P3_U4072, P3_U4073, P3_U4074, P3_U4075, P3_U4076, P3_U4077, P3_U4078, P3_U4079, P3_U4080, P3_U4081, P3_U4082, P3_U4083, P3_U4084, P3_U4085, P3_U4086, P3_U4087, P3_U4088, P3_U4089, P3_U4090, P3_U4091, P3_U4092, P3_U4093, P3_U4094, P3_U4095, P3_U4096, P3_U4097, P3_U4098, P3_U4099, P3_U4100, P3_U4101, P3_U4102, P3_U4103, P3_U4104, P3_U4105, P3_U4106, P3_U4107, P3_U4108, P3_U4109, P3_U4110, P3_U4111, P3_U4112, P3_U4113, P3_U4114, P3_U4115, P3_U4116, P3_U4117, P3_U4118, P3_U4119, P3_U4120, P3_U4121, P3_U4122, P3_U4123, P3_U4124, P3_U4125, P3_U4126, P3_U4127, P3_U4128, P3_U4129, P3_U4130, P3_U4131, P3_U4132, P3_U4133, P3_U4134, P3_U4135, P3_U4136, P3_U4137, P3_U4138, P3_U4139, P3_U4140, P3_U4141, P3_U4142, P3_U4143, P3_U4144, P3_U4145, P3_U4146, P3_U4147, P3_U4148, P3_U4149, P3_U4150, P3_U4151, P3_U4152, P3_U4153, P3_U4154, P3_U4155, P3_U4156, P3_U4157, P3_U4158, P3_U4159, P3_U4160, P3_U4161, P3_U4162, P3_U4163, P3_U4164, P3_U4165, P3_U4166, P3_U4167, P3_U4168, P3_U4169, P3_U4170, P3_U4171, P3_U4172, P3_U4173, P3_U4174, P3_U4175, P3_U4176, P3_U4177, P3_U4178, P3_U4179, P3_U4180, P3_U4181, P3_U4182, P3_U4183, P3_U4184, P3_U4185, P3_U4186, P3_U4187, P3_U4188, P3_U4189, P3_U4190, P3_U4191, P3_U4192, P3_U4193, P3_U4194, P3_U4195, P3_U4196, P3_U4197, P3_U4198, P3_U4199, P3_U4200, P3_U4201, P3_U4202, P3_U4203, P3_U4204, P3_U4205, P3_U4206, P3_U4207, P3_U4208, P3_U4209, P3_U4210, P3_U4211, P3_U4212, P3_U4213, P3_U4214, P3_U4215, P3_U4216, P3_U4217, P3_U4218, P3_U4219, P3_U4220, P3_U4221, P3_U4222, P3_U4223, P3_U4224, P3_U4225, P3_U4226, P3_U4227, P3_U4228, P3_U4229, P3_U4230, P3_U4231, P3_U4232, P3_U4233, P3_U4234, P3_U4235, P3_U4236, P3_U4237, P3_U4238, P3_U4239, P3_U4240, P3_U4241, P3_U4242, P3_U4243, P3_U4244, P3_U4245, P3_U4246, P3_U4247, P3_U4248, P3_U4249, P3_U4250, P3_U4251, P3_U4252, P3_U4253, P3_U4254, P3_U4255, P3_U4256, P3_U4257, P3_U4258, P3_U4259, P3_U4260, P3_U4261, P3_U4262, P3_U4263, P3_U4264, P3_U4265, P3_U4266, P3_U4267, P3_U4268, P3_U4269, P3_U4270, P3_U4271, P3_U4272, P3_U4273, P3_U4274, P3_U4275, P3_U4276, P3_U4277, P3_U4278, P3_U4279, P3_U4280, P3_U4281, P3_U4282, P3_U4283, P3_U4284, P3_U4285, P3_U4286, P3_U4287, P3_U4288, P3_U4289, P3_U4290, P3_U4291, P3_U4292, P3_U4293, P3_U4294, P3_U4295, P3_U4296, P3_U4297, P3_U4298, P3_U4299, P3_U4300, P3_U4301, P3_U4302, P3_U4303, P3_U4304, P3_U4305, P3_U4306, P3_U4307, P3_U4308, P3_U4309, P3_U4310, P3_U4311, P3_U4312, P3_U4313, P3_U4314, P3_U4315, P3_U4316, P3_U4317, P3_U4318, P3_U4319, P3_U4320, P3_U4321, P3_U4322, P3_U4323, P3_U4324, P3_U4325, P3_U4326, P3_U4327, P3_U4328, P3_U4329, P3_U4330, P3_U4331, P3_U4332, P3_U4333, P3_U4334, P3_U4335, P3_U4336, P3_U4337, P3_U4338, P3_U4339, P3_U4340, P3_U4341, P3_U4342, P3_U4343, P3_U4344, P3_U4345, P3_U4346, P3_U4347, P3_U4348, P3_U4349, P3_U4350, P3_U4351, P3_U4352, P3_U4353, P3_U4354, P3_U4355, P3_U4356, P3_U4357, P3_U4358, P3_U4359, P3_U4360, P3_U4361, P3_U4362, P3_U4363, P3_U4364, P3_U4365, P3_U4366, P3_U4367, P3_U4368, P3_U4369, P3_U4370, P3_U4371, P3_U4372, P3_U4373, P3_U4374, P3_U4375, P3_U4376, P3_U4377, P3_U4378, P3_U4379, P3_U4380, P3_U4381, P3_U4382, P3_U4383, P3_U4384, P3_U4385, P3_U4386, P3_U4387, P3_U4388, P3_U4389, P3_U4390, P3_U4391, P3_U4392, P3_U4393, P3_U4394, P3_U4395, P3_U4396, P3_U4397, P3_U4398, P3_U4399, P3_U4400, P3_U4401, P3_U4402, P3_U4403, P3_U4404, P3_U4405, P3_U4406, P3_U4407, P3_U4408, P3_U4409, P3_U4410, P3_U4411, P3_U4412, P3_U4413, P3_U4414, P3_U4415, P3_U4416, P3_U4417, P3_U4418, P3_U4419, P3_U4420, P3_U4421, P3_U4422, P3_U4423, P3_U4424, P3_U4425, P3_U4426, P3_U4427, P3_U4428, P3_U4429, P3_U4430, P3_U4431, P3_U4432, P3_U4433, P3_U4434, P3_U4435, P3_U4436, P3_U4437, P3_U4438, P3_U4439, P3_U4440, P3_U4441, P3_U4442, P3_U4443, P3_U4444, P3_U4445, P3_U4446, P3_U4447, P3_U4448, P3_U4449, P3_U4450, P3_U4451, P3_U4452, P3_U4453, P3_U4454, P3_U4455, P3_U4456, P3_U4457, P3_U4458, P3_U4459, P3_U4460, P3_U4461, P3_U4462, P3_U4463, P3_U4464, P3_U4465, P3_U4466, P3_U4467, P3_U4468, P3_U4469, P3_U4470, P3_U4471, P3_U4472, P3_U4473, P3_U4474, P3_U4475, P3_U4476, P3_U4477, P3_U4478, P3_U4479, P3_U4480, P3_U4481, P3_U4482, P3_U4483, P3_U4484, P3_U4485, P3_U4486, P3_U4487, P3_U4488, P3_U4489, P3_U4490, P3_U4491, P3_U4492, P3_U4493, P3_U4494, P3_U4495, P3_U4496, P3_U4497, P3_U4498, P3_U4499, P3_U4500, P3_U4501, P3_U4502, P3_U4503, P3_U4504, P3_U4505, P3_U4506, P3_U4507, P3_U4508, P3_U4509, P3_U4510, P3_U4511, P3_U4512, P3_U4513, P3_U4514, P3_U4515, P3_U4516, P3_U4517, P3_U4518, P3_U4519, P3_U4520, P3_U4521, P3_U4522, P3_U4523, P3_U4524, P3_U4525, P3_U4526, P3_U4527, P3_U4528, P3_U4529, P3_U4530, P3_U4531, P3_U4532, P3_U4533, P3_U4534, P3_U4535, P3_U4536, P3_U4537, P3_U4538, P3_U4539, P3_U4540, P3_U4541, P3_U4542, P3_U4543, P3_U4544, P3_U4545, P3_U4546, P3_U4547, P3_U4548, P3_U4549, P3_U4550, P3_U4551, P3_U4552, P3_U4553, P3_U4554, P3_U4555, P3_U4556, P3_U4557, P3_U4558, P3_U4559, P3_U4560, P3_U4561, P3_U4562, P3_U4563, P3_U4564, P3_U4565, P3_U4566, P3_U4567, P3_U4568, P3_U4569, P3_U4570, P3_U4571, P3_U4572, P3_U4573, P3_U4574, P3_U4575, P3_U4576, P3_U4577, P3_U4578, P3_U4579, P3_U4580, P3_U4581, P3_U4582, P3_U4583, P3_U4584, P3_U4585, P3_U4586, P3_U4587, P3_U4588, P3_U4589, P3_U4590, P3_U4591, P3_U4592, P3_U4593, P3_U4594, P3_U4595, P3_U4596, P3_U4597, P3_U4598, P3_U4599, P3_U4600, P3_U4601, P3_U4602, P3_U4603, P3_U4604, P3_U4605, P3_U4606, P3_U4607, P3_U4608, P3_U4609, P3_U4610, P3_U4611, P3_U4612, P3_U4613, P3_U4614, P3_U4615, P3_U4616, P3_U4617, P3_U4618, P3_U4619, P3_U4620, P3_U4621, P3_U4622, P3_U4623, P3_U4624, P3_U4625, P3_U4626, P3_U4627, P3_U4628, P3_U4629, P3_U4630, P3_U4631, P3_U4632, P3_U4633, P3_U4634, P3_U4635, P3_U4636, P3_U4637, P3_U4638, P3_U4639, P3_U4640, P3_U4641, P3_U4642, P3_U4643, P3_U4644, P3_U4645, P3_U4646, P3_U4647, P3_U4648, P3_U4649, P3_U4650, P3_U4651, P3_U4652, P3_U4653, P3_U4654, P3_U4655, P3_U4656, P3_U4657, P3_U4658, P3_U4659, P3_U4660, P3_U4661, P3_U4662, P3_U4663, P3_U4664, P3_U4665, P3_U4666, P3_U4667, P3_U4668, P3_U4669, P3_U4670, P3_U4671, P3_U4672, P3_U4673, P3_U4674, P3_U4675, P3_U4676, P3_U4677, P3_U4678, P3_U4679, P3_U4680, P3_U4681, P3_U4682, P3_U4683, P3_U4684, P3_U4685, P3_U4686, P3_U4687, P3_U4688, P3_U4689, P3_U4690, P3_U4691, P3_U4692, P3_U4693, P3_U4694, P3_U4695, P3_U4696, P3_U4697, P3_U4698, P3_U4699, P3_U4700, P3_U4701, P3_U4702, P3_U4703, P3_U4704, P3_U4705, P3_U4706, P3_U4707, P3_U4708, P3_U4709, P3_U4710, P3_U4711, P3_U4712, P3_U4713, P3_U4714, P3_U4715, P3_U4716, P3_U4717, P3_U4718, P3_U4719, P3_U4720, P3_U4721, P3_U4722, P3_U4723, P3_U4724, P3_U4725, P3_U4726, P3_U4727, P3_U4728, P3_U4729, P3_U4730, P3_U4731, P3_U4732, P3_U4733, P3_U4734, P3_U4735, P3_U4736, P3_U4737, P3_U4738, P3_U4739, P3_U4740, P3_U4741, P3_U4742, P3_U4743, P3_U4744, P3_U4745, P3_U4746, P3_U4747, P3_U4748, P3_U4749, P3_U4750, P3_U4751, P3_U4752, P3_U4753, P3_U4754, P3_U4755, P3_U4756, P3_U4757, P3_U4758, P3_U4759, P3_U4760, P3_U4761, P3_U4762, P3_U4763, P3_U4764, P3_U4765, P3_U4766, P3_U4767, P3_U4768, P3_U4769, P3_U4770, P3_U4771, P3_U4772, P3_U4773, P3_U4774, P3_U4775, P3_U4776, P3_U4777, P3_U4778, P3_U4779, P3_U4780, P3_U4781, P3_U4782, P3_U4783, P3_U4784, P3_U4785, P3_U4786, P3_U4787, P3_U4788, P3_U4789, P3_U4790, P3_U4791, P3_U4792, P3_U4793, P3_U4794, P3_U4795, P3_U4796, P3_U4797, P3_U4798, P3_U4799, P3_U4800, P3_U4801, P3_U4802, P3_U4803, P3_U4804, P3_U4805, P3_U4806, P3_U4807, P3_U4808, P3_U4809, P3_U4810, P3_U4811, P3_U4812, P3_U4813, P3_U4814, P3_U4815, P3_U4816, P3_U4817, P3_U4818, P3_U4819, P3_U4820, P3_U4821, P3_U4822, P3_U4823, P3_U4824, P3_U4825, P3_U4826, P3_U4827, P3_U4828, P3_U4829, P3_U4830, P3_U4831, P3_U4832, P3_U4833, P3_U4834, P3_U4835, P3_U4836, P3_U4837, P3_U4838, P3_U4839, P3_U4840, P3_U4841, P3_U4842, P3_U4843, P3_U4844, P3_U4845, P3_U4846, P3_U4847, P3_U4848, P3_U4849, P3_U4850, P3_U4851, P3_U4852, P3_U4853, P3_U4854, P3_U4855, P3_U4856, P3_U4857, P3_U4858, P3_U4859, P3_U4860, P3_U4861, P3_U4862, P3_U4863, P3_U4864, P3_U4865, P3_U4866, P3_U4867, P3_U4868, P3_U4869, P3_U4870, P3_U4871, P3_U4872, P3_U4873, P3_U4874, P3_U4875, P3_U4876, P3_U4877, P3_U4878, P3_U4879, P3_U4880, P3_U4881, P3_U4882, P3_U4883, P3_U4884, P3_U4885, P3_U4886, P3_U4887, P3_U4888, P3_U4889, P3_U4890, P3_U4891, P3_U4892, P3_U4893, P3_U4894, P3_U4895, P3_U4896, P3_U4897, P3_U4898, P3_U4899, P3_U4900, P3_U4901, P3_U4902, P3_U4903, P3_U4904, P3_U4905, P3_U4906, P3_U4907, P3_U4908, P3_U4909, P3_U4910, P3_U4911, P3_U4912, P3_U4913, P3_U4914, P3_U4915, P3_U4916, P3_U4917, P3_U4918, P3_U4919, P3_U4920, P3_U4921, P3_U4922, P3_U4923, P3_U4924, P3_U4925, P3_U4926, P3_U4927, P3_U4928, P3_U4929, P3_U4930, P3_U4931, P3_U4932, P3_U4933, P3_U4934, P3_U4935, P3_U4936, P3_U4937, P3_U4938, P3_U4939, P3_U4940, P3_U4941, P3_U4942, P3_U4943, P3_U4944, P3_U4945, P3_U4946, P3_U4947, P3_U4948, P3_U4949, P3_U4950, P3_U4951, P3_U4952, P3_U4953, P3_U4954, P3_U4955, P3_U4956, P3_U4957, P3_U4958, P3_U4959, P3_U4960, P3_U4961, P3_U4962, P3_U4963, P3_U4964, P3_U4965, P3_U4966, P3_U4967, P3_U4968, P3_U4969, P3_U4970, P3_U4971, P3_U4972, P3_U4973, P3_U4974, P3_U4975, P3_U4976, P3_U4977, P3_U4978, P3_U4979, P3_U4980, P3_U4981, P3_U4982, P3_U4983, P3_U4984, P3_U4985, P3_U4986, P3_U4987, P3_U4988, P3_U4989, P3_U4990, P3_U4991, P3_U4992, P3_U4993, P3_U4994, P3_U4995, P3_U4996, P3_U4997, P3_U4998, P3_U4999, P3_U5000, P3_U5001, P3_U5002, P3_U5003, P3_U5004, P3_U5005, P3_U5006, P3_U5007, P3_U5008, P3_U5009, P3_U5010, P3_U5011, P3_U5012, P3_U5013, P3_U5014, P3_U5015, P3_U5016, P3_U5017, P3_U5018, P3_U5019, P3_U5020, P3_U5021, P3_U5022, P3_U5023, P3_U5024, P3_U5025, P3_U5026, P3_U5027, P3_U5028, P3_U5029, P3_U5030, P3_U5031, P3_U5032, P3_U5033, P3_U5034, P3_U5035, P3_U5036, P3_U5037, P3_U5038, P3_U5039, P3_U5040, P3_U5041, P3_U5042, P3_U5043, P3_U5044, P3_U5045, P3_U5046, P3_U5047, P3_U5048, P3_U5049, P3_U5050, P3_U5051, P3_U5052, P3_U5053, P3_U5054, P3_U5055, P3_U5056, P3_U5057, P3_U5058, P3_U5059, P3_U5060, P3_U5061, P3_U5062, P3_U5063, P3_U5064, P3_U5065, P3_U5066, P3_U5067, P3_U5068, P3_U5069, P3_U5070, P3_U5071, P3_U5072, P3_U5073, P3_U5074, P3_U5075, P3_U5076, P3_U5077, P3_U5078, P3_U5079, P3_U5080, P3_U5081, P3_U5082, P3_U5083, P3_U5084, P3_U5085, P3_U5086, P3_U5087, P3_U5088, P3_U5089, P3_U5090, P3_U5091, P3_U5092, P3_U5093, P3_U5094, P3_U5095, P3_U5096, P3_U5097, P3_U5098, P3_U5099, P3_U5100, P3_U5101, P3_U5102, P3_U5103, P3_U5104, P3_U5105, P3_U5106, P3_U5107, P3_U5108, P3_U5109, P3_U5110, P3_U5111, P3_U5112, P3_U5113, P3_U5114, P3_U5115, P3_U5116, P3_U5117, P3_U5118, P3_U5119, P3_U5120, P3_U5121, P3_U5122, P3_U5123, P3_U5124, P3_U5125, P3_U5126, P3_U5127, P3_U5128, P3_U5129, P3_U5130, P3_U5131, P3_U5132, P3_U5133, P3_U5134, P3_U5135, P3_U5136, P3_U5137, P3_U5138, P3_U5139, P3_U5140, P3_U5141, P3_U5142, P3_U5143, P3_U5144, P3_U5145, P3_U5146, P3_U5147, P3_U5148, P3_U5149, P3_U5150, P3_U5151, P3_U5152, P3_U5153, P3_U5154, P3_U5155, P3_U5156, P3_U5157, P3_U5158, P3_U5159, P3_U5160, P3_U5161, P3_U5162, P3_U5163, P3_U5164, P3_U5165, P3_U5166, P3_U5167, P3_U5168, P3_U5169, P3_U5170, P3_U5171, P3_U5172, P3_U5173, P3_U5174, P3_U5175, P3_U5176, P3_U5177, P3_U5178, P3_U5179, P3_U5180, P3_U5181, P3_U5182, P3_U5183, P3_U5184, P3_U5185, P3_U5186, P3_U5187, P3_U5188, P3_U5189, P3_U5190, P3_U5191, P3_U5192, P3_U5193, P3_U5194, P3_U5195, P3_U5196, P3_U5197, P3_U5198, P3_U5199, P3_U5200, P3_U5201, P3_U5202, P3_U5203, P3_U5204, P3_U5205, P3_U5206, P3_U5207, P3_U5208, P3_U5209, P3_U5210, P3_U5211, P3_U5212, P3_U5213, P3_U5214, P3_U5215, P3_U5216, P3_U5217, P3_U5218, P3_U5219, P3_U5220, P3_U5221, P3_U5222, P3_U5223, P3_U5224, P3_U5225, P3_U5226, P3_U5227, P3_U5228, P3_U5229, P3_U5230, P3_U5231, P3_U5232, P3_U5233, P3_U5234, P3_U5235, P3_U5236, P3_U5237, P3_U5238, P3_U5239, P3_U5240, P3_U5241, P3_U5242, P3_U5243, P3_U5244, P3_U5245, P3_U5246, P3_U5247, P3_U5248, P3_U5249, P3_U5250, P3_U5251, P3_U5252, P3_U5253, P3_U5254, P3_U5255, P3_U5256, P3_U5257, P3_U5258, P3_U5259, P3_U5260, P3_U5261, P3_U5262, P3_U5263, P3_U5264, P3_U5265, P3_U5266, P3_U5267, P3_U5268, P3_U5269, P3_U5270, P3_U5271, P3_U5272, P3_U5273, P3_U5274, P3_U5275, P3_U5276, P3_U5277, P3_U5278, P3_U5279, P3_U5280, P3_U5281, P3_U5282, P3_U5283, P3_U5284, P3_U5285, P3_U5286, P3_U5287, P3_U5288, P3_U5289, P3_U5290, P3_U5291, P3_U5292, P3_U5293, P3_U5294, P3_U5295, P3_U5296, P3_U5297, P3_U5298, P3_U5299, P3_U5300, P3_U5301, P3_U5302, P3_U5303, P3_U5304, P3_U5305, P3_U5306, P3_U5307, P3_U5308, P3_U5309, P3_U5310, P3_U5311, P3_U5312, P3_U5313, P3_U5314, P3_U5315, P3_U5316, P3_U5317, P3_U5318, P3_U5319, P3_U5320, P3_U5321, P3_U5322, P3_U5323, P3_U5324, P3_U5325, P3_U5326, P3_U5327, P3_U5328, P3_U5329, P3_U5330, P3_U5331, P3_U5332, P3_U5333, P3_U5334, P3_U5335, P3_U5336, P3_U5337, P3_U5338, P3_U5339, P3_U5340, P3_U5341, P3_U5342, P3_U5343, P3_U5344, P3_U5345, P3_U5346, P3_U5347, P3_U5348, P3_U5349, P3_U5350, P3_U5351, P3_U5352, P3_U5353, P3_U5354, P3_U5355, P3_U5356, P3_U5357, P3_U5358, P3_U5359, P3_U5360, P3_U5361, P3_U5362, P3_U5363, P3_U5364, P3_U5365, P3_U5366, P3_U5367, P3_U5368, P3_U5369, P3_U5370, P3_U5371, P3_U5372, P3_U5373, P3_U5374, P3_U5375, P3_U5376, P3_U5377, P3_U5378, P3_U5379, P3_U5380, P3_U5381, P3_U5382, P3_U5383, P3_U5384, P3_U5385, P3_U5386, P3_U5387, P3_U5388, P3_U5389, P3_U5390, P3_U5391, P3_U5392, P3_U5393, P3_U5394, P3_U5395, P3_U5396, P3_U5397, P3_U5398, P3_U5399, P3_U5400, P3_U5401, P3_U5402, P3_U5403, P3_U5404, P3_U5405, P3_U5406, P3_U5407, P3_U5408, P3_U5409, P3_U5410, P3_U5411, P3_U5412, P3_U5413, P3_U5414, P3_U5415, P3_U5416, P3_U5417, P3_U5418, P3_U5419, P3_U5420, P3_U5421, P3_U5422, P3_U5423, P3_U5424, P3_U5425, P3_U5426, P3_U5427, P3_U5428, P3_U5429, P3_U5430, P3_U5431, P3_U5432, P3_U5433, P3_U5434, P3_U5435, P3_U5436, P3_U5437, P3_U5438, P3_U5439, P3_U5440, P3_U5441, P3_U5442, P3_U5443, P3_U5444, P3_U5445, P3_U5446, P3_U5447, P3_U5448, P3_U5449, P3_U5450, P3_U5451, P3_U5452, P3_U5453, P3_U5454, P3_U5455, P3_U5456, P3_U5457, P3_U5458, P3_U5459, P3_U5460, P3_U5461, P3_U5462, P3_U5463, P3_U5464, P3_U5465, P3_U5466, P3_U5467, P3_U5468, P3_U5469, P3_U5470, P3_U5471, P3_U5472, P3_U5473, P3_U5474, P3_U5475, P3_U5476, P3_U5477, P3_U5478, P3_U5479, P3_U5480, P3_U5481, P3_U5482, P3_U5483, P3_U5484, P3_U5485, P3_U5486, P3_U5487, P3_U5488, P3_U5489, P3_U5490, P3_U5491, P3_U5492, P3_U5493, P3_U5494, P3_U5495, P3_U5496, P3_U5497, P3_U5498, P3_U5499, P3_U5500, P3_U5501, P3_U5502, P3_U5503, P3_U5504, P3_U5505, P3_U5506, P3_U5507, P3_U5508, P3_U5509, P3_U5510, P3_U5511, P3_U5512, P3_U5513, P3_U5514, P3_U5515, P3_U5516, P3_U5517, P3_U5518, P3_U5519, P3_U5520, P3_U5521, P3_U5522, P3_U5523, P3_U5524, P3_U5525, P3_U5526, P3_U5527, P3_U5528, P3_U5529, P3_U5530, P3_U5531, P3_U5532, P3_U5533, P3_U5534, P3_U5535, P3_U5536, P3_U5537, P3_U5538, P3_U5539, P3_U5540, P3_U5541, P3_U5542, P3_U5543, P3_U5544, P3_U5545, P3_U5546, P3_U5547, P3_U5548, P3_U5549, P3_U5550, P3_U5551, P3_U5552, P3_U5553, P3_U5554, P3_U5555, P3_U5556, P3_U5557, P3_U5558, P3_U5559, P3_U5560, P3_U5561, P3_U5562, P3_U5563, P3_U5564, P3_U5565, P3_U5566, P3_U5567, P3_U5568, P3_U5569, P3_U5570, P3_U5571, P3_U5572, P3_U5573, P3_U5574, P3_U5575, P3_U5576, P3_U5577, P3_U5578, P3_U5579, P3_U5580, P3_U5581, P3_U5582, P3_U5583, P3_U5584, P3_U5585, P3_U5586, P3_U5587, P3_U5588, P3_U5589, P3_U5590, P3_U5591, P3_U5592, P3_U5593, P3_U5594, P3_U5595, P3_U5596, P3_U5597, P3_U5598, P3_U5599, P3_U5600, P3_U5601, P3_U5602, P3_U5603, P3_U5604, P3_U5605, P3_U5606, P3_U5607, P3_U5608, P3_U5609, P3_U5610, P3_U5611, P3_U5612, P3_U5613, P3_U5614, P3_U5615, P3_U5616, P3_U5617, P3_U5618, P3_U5619, P3_U5620, P3_U5621, P3_U5622, P3_U5623, P3_U5624, P3_U5625, P3_U5626, P3_U5627, P3_U5628, P3_U5629, P3_U5630, P3_U5631, P3_U5632, P3_U5633, P3_U5634, P3_U5635, P3_U5636, P3_U5637, P3_U5638, P3_U5639, P3_U5640, P3_U5641, P3_U5642, P3_U5643, P3_U5644, P3_U5645, P3_U5646, P3_U5647, P3_U5648, P3_U5649, P3_U5650, P3_U5651, P3_U5652, P3_U5653, P3_U5654, P3_U5655, P3_U5656, P3_U5657, P3_U5658, P3_U5659, P3_U5660, P3_U5661, P3_U5662, P3_U5663, P3_U5664, P3_U5665, P3_U5666, P3_U5667, P3_U5668, P3_U5669, P3_U5670, P3_U5671, P3_U5672, P3_U5673, P3_U5674, P3_U5675, P3_U5676, P3_U5677, P3_U5678, P3_U5679, P3_U5680, P3_U5681, P3_U5682, P3_U5683, P3_U5684, P3_U5685, P3_U5686, P3_U5687, P3_U5688, P3_U5689, P3_U5690, P3_U5691, P3_U5692, P3_U5693, P3_U5694, P3_U5695, P3_U5696, P3_U5697, P3_U5698, P3_U5699, P3_U5700, P3_U5701, P3_U5702, P3_U5703, P3_U5704, P3_U5705, P3_U5706, P3_U5707, P3_U5708, P3_U5709, P3_U5710, P3_U5711, P3_U5712, P3_U5713, P3_U5714, P3_U5715, P3_U5716, P3_U5717, P3_U5718, P3_U5719, P3_U5720, P3_U5721, P3_U5722, P3_U5723, P3_U5724, P3_U5725, P3_U5726, P3_U5727, P3_U5728, P3_U5729, P3_U5730, P3_U5731, P3_U5732, P3_U5733, P3_U5734, P3_U5735, P3_U5736, P3_U5737, P3_U5738, P3_U5739, P3_U5740, P3_U5741, P3_U5742, P3_U5743, P3_U5744, P3_U5745, P3_U5746, P3_U5747, P3_U5748, P3_U5749, P3_U5750, P3_U5751, P3_U5752, P3_U5753, P3_U5754, P3_U5755, P3_U5756, P3_U5757, P3_U5758, P3_U5759, P3_U5760, P3_U5761, P3_U5762, P3_U5763, P3_U5764, P3_U5765, P3_U5766, P3_U5767, P3_U5768, P3_U5769, P3_U5770, P3_U5771, P3_U5772, P3_U5773, P3_U5774, P3_U5775, P3_U5776, P3_U5777, P3_U5778, P3_U5779, P3_U5780, P3_U5781, P3_U5782, P3_U5783, P3_U5784, P3_U5785, P3_U5786, P3_U5787, P3_U5788, P3_U5789, P3_U5790, P3_U5791, P3_U5792, P3_U5793, P3_U5794, P3_U5795, P3_U5796, P3_U5797, P3_U5798, P3_U5799, P3_U5800, P3_U5801, P3_U5802, P3_U5803, P3_U5804, P3_U5805, P3_U5806, P3_U5807, P3_U5808, P3_U5809, P3_U5810, P3_U5811, P3_U5812, P3_U5813, P3_U5814, P3_U5815, P3_U5816, P3_U5817, P3_U5818, P3_U5819, P3_U5820, P3_U5821, P3_U5822, P3_U5823, P3_U5824, P3_U5825, P3_U5826, P3_U5827, P3_U5828, P3_U5829, P3_U5830, P3_U5831, P3_U5832, P3_U5833, P3_U5834, P3_U5835, P3_U5836, P3_U5837, P3_U5838, P3_U5839, P3_U5840, P3_U5841, P3_U5842, P3_U5843, P3_U5844, P3_U5845, P3_U5846, P3_U5847, P3_U5848, P3_U5849, P3_U5850, P3_U5851, P3_U5852, P3_U5853, P3_U5854, P3_U5855, P3_U5856, P3_U5857, P3_U5858, P3_U5859, P3_U5860, P3_U5861, P3_U5862, P3_U5863, P3_U5864, P3_U5865, P3_U5866, P3_U5867, P3_U5868, P3_U5869, P3_U5870, P3_U5871, P3_U5872, P3_U5873, P3_U5874, P3_U5875, P3_U5876, P3_U5877, P3_U5878, P3_U5879, P3_U5880, P3_U5881, P3_U5882, P3_U5883, P3_U5884, P3_U5885, P3_U5886, P3_U5887, P3_U5888, P3_U5889, P3_U5890, P3_U5891, P3_U5892, P3_U5893, P3_U5894, P3_U5895, P3_U5896, P3_U5897, P3_U5898, P3_U5899, P3_U5900, P3_U5901, P3_U5902, P3_U5903, P3_U5904, P3_U5905, P3_U5906, P3_U5907, P3_U5908, P3_U5909, P3_U5910, P3_U5911, P3_U5912, P3_U5913, P3_U5914, P3_U5915, P3_U5916, P3_U5917, P3_U5918, P3_U5919, P3_U5920, P3_U5921, P3_U5922, P3_U5923, P3_U5924, P3_U5925, P3_U5926, P3_U5927, P3_U5928, P3_U5929, P3_U5930, P3_U5931, P3_U5932, P3_U5933, P3_U5934, P3_U5935, P3_U5936, P3_U5937, P3_U5938, P3_U5939, P3_U5940, P3_U5941, P3_U5942, P3_U5943, P3_U5944, P3_U5945, P3_U5946, P3_U5947, P3_U5948, P3_U5949, P3_U5950, P3_U5951, P3_U5952, P3_U5953, P3_U5954, P3_U5955, P3_U5956, P3_U5957, P3_U5958, P3_U5959, P3_U5960, P3_U5961, P3_U5962, P3_U5963, P3_U5964, P3_U5965, P3_U5966, P3_U5967, P3_U5968, P3_U5969, P3_U5970, P3_U5971, P3_U5972, P3_U5973, P3_U5974, P3_U5975, P3_U5976, P3_U5977, P3_U5978, P3_U5979, P3_U5980, P3_U5981, P3_U5982, P3_U5983, P3_U5984, P3_U5985, P3_U5986, P3_U5987, P3_U5988, P3_U5989, P3_U5990, P3_U5991, P3_U5992, P3_U5993, P3_U5994, P3_U5995, P3_U5996, P3_U5997, P3_U5998, P3_U5999, P3_U6000, P3_U6001, P3_U6002, P3_U6003, P3_U6004, P3_U6005, P3_U6006, P3_U6007, P3_U6008, P3_U6009, P3_U6010, P3_U6011, P3_U6012, P3_U6013, P3_U6014, P3_U6015, P3_U6016, P3_U6017, P3_U6018, P3_U6019, P3_U6020, P3_U6021, P3_U6022, P3_U6023, P3_U6024, P3_U6025, P3_U6026, P3_U6027, P3_U6028, P3_U6029, P3_U6030, P3_U6031, P3_U6032, P3_U6033, P3_U6034, P3_U6035, P3_U6036, P3_U6037, P3_U6038, P3_U6039, P3_U6040, P3_U6041, P3_U6042, P3_U6043, P3_U6044, P3_U6045, P3_U6046, P3_U6047, P3_U6048, P3_U6049, P3_U6050, P3_U6051, P3_U6052, P3_U6053, P3_U6054, P3_U6055, P3_U6056, P3_U6057, P3_U6058, P3_U6059, P3_U6060, P3_U6061, P3_U6062, P3_U6063, P3_U6064, P3_U6065, P3_U6066, P3_U6067, P3_U6068, P3_U6069, P3_U6070, P3_U6071, P3_U6072, P3_U6073, P3_U6074, P3_U6075, P3_U6076, P3_U6077, P3_U6078, P3_U6079, P3_U6080, P3_U6081, P3_U6082, P3_U6083, P3_U6084, P3_U6085, P3_U6086, P3_U6087, P3_U6088, P3_U6089, P3_U6090, P3_U6091, P3_U6092, P3_U6093, P3_U6094, P3_U6095, P3_U6096, P3_U6097, P3_U6098, P3_U6099, P3_U6100, P3_U6101, P3_U6102, P3_U6103, P3_U6104, P3_U6105, P3_U6106, P3_U6107, P3_U6108, P3_U6109, P3_U6110, P3_U6111, P3_U6112, P3_U6113, P3_U6114, P3_U6115, P3_U6116, P3_U6117, P3_U6118, P3_U6119, P3_U6120, P3_U6121, P3_U6122, P3_U6123, P3_U6124, P3_U6125, P3_U6126, P3_U6127, P3_U6128, P3_U6129, P3_U6130, P3_U6131, P3_U6132, P3_U6133, P3_U6134, P3_U6135, P3_U6136, P3_U6137, P3_U6138, P3_U6139, P3_U6140, P3_U6141, P3_U6142, P3_U6143, P3_U6144, P3_U6145, P3_U6146, P3_U6147, P3_U6148, P3_U6149, P3_U6150, P3_U6151, P3_U6152, P3_U6153, P3_U6154, P3_U6155, P3_U6156, P3_U6157, P3_U6158, P3_U6159, P3_U6160, P3_U6161, P3_U6162, P3_U6163, P3_U6164, P3_U6165, P3_U6166, P3_U6167, P3_U6168, P3_U6169, P3_U6170, P3_U6171, P3_U6172, P3_U6173, P3_U6174, P3_U6175, P3_U6176, P3_U6177, P3_U6178, P3_U6179, P3_U6180, P3_U6181, P3_U6182, P3_U6183, P3_U6184, P3_U6185, P3_U6186, P3_U6187, P3_U6188, P3_U6189, P3_U6190, P3_U6191, P3_U6192, P3_U6193, P3_U6194, P3_U6195, P3_U6196, P3_U6197, P3_U6198, P3_U6199, P3_U6200, P3_U6201, P3_U6202, P3_U6203, P3_U6204, P3_U6205, P3_U6206, P3_U6207, P3_U6208, P3_U6209, P3_U6210, P3_U6211, P3_U6212, P3_U6213, P3_U6214, P3_U6215, P3_U6216, P3_U6217, P3_U6218, P3_U6219, P3_U6220, P3_U6221, P3_U6222, P3_U6223, P3_U6224, P3_U6225, P3_U6226, P3_U6227, P3_U6228, P3_U6229, P3_U6230, P3_U6231, P3_U6232, P3_U6233, P3_U6234, P3_U6235, P3_U6236, P3_U6237, P3_U6238, P3_U6239, P3_U6240, P3_U6241, P3_U6242, P3_U6243, P3_U6244, P3_U6245, P3_U6246, P3_U6247, P3_U6248, P3_U6249, P3_U6250, P3_U6251, P3_U6252, P3_U6253, P3_U6254, P3_U6255, P3_U6256, P3_U6257, P3_U6258, P3_U6259, P3_U6260, P3_U6261, P3_U6262, P3_U6263, P3_U6264, P3_U6265, P3_U6266, P3_U6267, P3_U6268, P3_U6269, P3_U6270, P3_U6271, P3_U6272, P3_U6273, P3_U6274, P3_U6275, P3_U6276, P3_U6277, P3_U6278, P3_U6279, P3_U6280, P3_U6281, P3_U6282, P3_U6283, P3_U6284, P3_U6285, P3_U6286, P3_U6287, P3_U6288, P3_U6289, P3_U6290, P3_U6291, P3_U6292, P3_U6293, P3_U6294, P3_U6295, P3_U6296, P3_U6297, P3_U6298, P3_U6299, P3_U6300, P3_U6301, P3_U6302, P3_U6303, P3_U6304, P3_U6305, P3_U6306, P3_U6307, P3_U6308, P3_U6309, P3_U6310, P3_U6311, P3_U6312, P3_U6313, P3_U6314, P3_U6315, P3_U6316, P3_U6317, P3_U6318, P3_U6319, P3_U6320, P3_U6321, P3_U6322, P3_U6323, P3_U6324, P3_U6325, P3_U6326, P3_U6327, P3_U6328, P3_U6329, P3_U6330, P3_U6331, P3_U6332, P3_U6333, P3_U6334, P3_U6335, P3_U6336, P3_U6337, P3_U6338, P3_U6339, P3_U6340, P3_U6341, P3_U6342, P3_U6343, P3_U6344, P3_U6345, P3_U6346, P3_U6347, P3_U6348, P3_U6349, P3_U6350, P3_U6351, P3_U6352, P3_U6353, P3_U6354, P3_U6355, P3_U6356, P3_U6357, P3_U6358, P3_U6359, P3_U6360, P3_U6361, P3_U6362, P3_U6363, P3_U6364, P3_U6365, P3_U6366, P3_U6367, P3_U6368, P3_U6369, P3_U6370, P3_U6371, P3_U6372, P3_U6373, P3_U6374, P3_U6375, P3_U6376, P3_U6377, P3_U6378, P3_U6379, P3_U6380, P3_U6381, P3_U6382, P3_U6383, P3_U6384, P3_U6385, P3_U6386, P3_U6387, P3_U6388, P3_U6389, P3_U6390, P3_U6391, P3_U6392, P3_U6393, P3_U6394, P3_U6395, P3_U6396, P3_U6397, P3_U6398, P3_U6399, P3_U6400, P3_U6401, P3_U6402, P3_U6403, P3_U6404, P3_U6405, P3_U6406, P3_U6407, P3_U6408, P3_U6409, P3_U6410, P3_U6411, P3_U6412, P3_U6413, P3_U6414, P3_U6415, P3_U6416, P3_U6417, P3_U6418, P3_U6419, P3_U6420, P3_U6421, P3_U6422, P3_U6423, P3_U6424, P3_U6425, P3_U6426, P3_U6427, P3_U6428, P3_U6429, P3_U6430, P3_U6431, P3_U6432, P3_U6433, P3_U6434, P3_U6435, P3_U6436, P3_U6437, P3_U6438, P3_U6439, P3_U6440, P3_U6441, P3_U6442, P3_U6443, P3_U6444, P3_U6445, P3_U6446, P3_U6447, P3_U6448, P3_U6449, P3_U6450, P3_U6451, P3_U6452, P3_U6453, P3_U6454, P3_U6455, P3_U6456, P3_U6457, P3_U6458, P3_U6459, P3_U6460, P3_U6461, P3_U6462, P3_U6463, P3_U6464, P3_U6465, P3_U6466, P3_U6467, P3_U6468, P3_U6469, P3_U6470, P3_U6471, P3_U6472, P3_U6473, P3_U6474, P3_U6475, P3_U6476, P3_U6477, P3_U6478, P3_U6479, P3_U6480, P3_U6481, P3_U6482, P3_U6483, P3_U6484, P3_U6485, P3_U6486, P3_U6487, P3_U6488, P3_U6489, P3_U6490, P3_U6491, P3_U6492, P3_U6493, P3_U6494, P3_U6495, P3_U6496, P3_U6497, P3_U6498, P3_U6499, P3_U6500, P3_U6501, P3_U6502, P3_U6503, P3_U6504, P3_U6505, P3_U6506, P3_U6507, P3_U6508, P3_U6509, P3_U6510, P3_U6511, P3_U6512, P3_U6513, P3_U6514, P3_U6515, P3_U6516, P3_U6517, P3_U6518, P3_U6519, P3_U6520, P3_U6521, P3_U6522, P3_U6523, P3_U6524, P3_U6525, P3_U6526, P3_U6527, P3_U6528, P3_U6529, P3_U6530, P3_U6531, P3_U6532, P3_U6533, P3_U6534, P3_U6535, P3_U6536, P3_U6537, P3_U6538, P3_U6539, P3_U6540, P3_U6541, P3_U6542, P3_U6543, P3_U6544, P3_U6545, P3_U6546, P3_U6547, P3_U6548, P3_U6549, P3_U6550, P3_U6551, P3_U6552, P3_U6553, P3_U6554, P3_U6555, P3_U6556, P3_U6557, P3_U6558, P3_U6559, P3_U6560, P3_U6561, P3_U6562, P3_U6563, P3_U6564, P3_U6565, P3_U6566, P3_U6567, P3_U6568, P3_U6569, P3_U6570, P3_U6571, P3_U6572, P3_U6573, P3_U6574, P3_U6575, P3_U6576, P3_U6577, P3_U6578, P3_U6579, P3_U6580, P3_U6581, P3_U6582, P3_U6583, P3_U6584, P3_U6585, P3_U6586, P3_U6587, P3_U6588, P3_U6589, P3_U6590, P3_U6591, P3_U6592, P3_U6593, P3_U6594, P3_U6595, P3_U6596, P3_U6597, P3_U6598, P3_U6599, P3_U6600, P3_U6601, P3_U6602, P3_U6603, P3_U6604, P3_U6605, P3_U6606, P3_U6607, P3_U6608, P3_U6609, P3_U6610, P3_U6611, P3_U6612, P3_U6613, P3_U6614, P3_U6615, P3_U6616, P3_U6617, P3_U6618, P3_U6619, P3_U6620, P3_U6621, P3_U6622, P3_U6623, P3_U6624, P3_U6625, P3_U6626, P3_U6627, P3_U6628, P3_U6629, P3_U6630, P3_U6631, P3_U6632, P3_U6633, P3_U6634, P3_U6635, P3_U6636, P3_U6637, P3_U6638, P3_U6639, P3_U6640, P3_U6641, P3_U6642, P3_U6643, P3_U6644, P3_U6645, P3_U6646, P3_U6647, P3_U6648, P3_U6649, P3_U6650, P3_U6651, P3_U6652, P3_U6653, P3_U6654, P3_U6655, P3_U6656, P3_U6657, P3_U6658, P3_U6659, P3_U6660, P3_U6661, P3_U6662, P3_U6663, P3_U6664, P3_U6665, P3_U6666, P3_U6667, P3_U6668, P3_U6669, P3_U6670, P3_U6671, P3_U6672, P3_U6673, P3_U6674, P3_U6675, P3_U6676, P3_U6677, P3_U6678, P3_U6679, P3_U6680, P3_U6681, P3_U6682, P3_U6683, P3_U6684, P3_U6685, P3_U6686, P3_U6687, P3_U6688, P3_U6689, P3_U6690, P3_U6691, P3_U6692, P3_U6693, P3_U6694, P3_U6695, P3_U6696, P3_U6697, P3_U6698, P3_U6699, P3_U6700, P3_U6701, P3_U6702, P3_U6703, P3_U6704, P3_U6705, P3_U6706, P3_U6707, P3_U6708, P3_U6709, P3_U6710, P3_U6711, P3_U6712, P3_U6713, P3_U6714, P3_U6715, P3_U6716, P3_U6717, P3_U6718, P3_U6719, P3_U6720, P3_U6721, P3_U6722, P3_U6723, P3_U6724, P3_U6725, P3_U6726, P3_U6727, P3_U6728, P3_U6729, P3_U6730, P3_U6731, P3_U6732, P3_U6733, P3_U6734, P3_U6735, P3_U6736, P3_U6737, P3_U6738, P3_U6739, P3_U6740, P3_U6741, P3_U6742, P3_U6743, P3_U6744, P3_U6745, P3_U6746, P3_U6747, P3_U6748, P3_U6749, P3_U6750, P3_U6751, P3_U6752, P3_U6753, P3_U6754, P3_U6755, P3_U6756, P3_U6757, P3_U6758, P3_U6759, P3_U6760, P3_U6761, P3_U6762, P3_U6763, P3_U6764, P3_U6765, P3_U6766, P3_U6767, P3_U6768, P3_U6769, P3_U6770, P3_U6771, P3_U6772, P3_U6773, P3_U6774, P3_U6775, P3_U6776, P3_U6777, P3_U6778, P3_U6779, P3_U6780, P3_U6781, P3_U6782, P3_U6783, P3_U6784, P3_U6785, P3_U6786, P3_U6787, P3_U6788, P3_U6789, P3_U6790, P3_U6791, P3_U6792, P3_U6793, P3_U6794, P3_U6795, P3_U6796, P3_U6797, P3_U6798, P3_U6799, P3_U6800, P3_U6801, P3_U6802, P3_U6803, P3_U6804, P3_U6805, P3_U6806, P3_U6807, P3_U6808, P3_U6809, P3_U6810, P3_U6811, P3_U6812, P3_U6813, P3_U6814, P3_U6815, P3_U6816, P3_U6817, P3_U6818, P3_U6819, P3_U6820, P3_U6821, P3_U6822, P3_U6823, P3_U6824, P3_U6825, P3_U6826, P3_U6827, P3_U6828, P3_U6829, P3_U6830, P3_U6831, P3_U6832, P3_U6833, P3_U6834, P3_U6835, P3_U6836, P3_U6837, P3_U6838, P3_U6839, P3_U6840, P3_U6841, P3_U6842, P3_U6843, P3_U6844, P3_U6845, P3_U6846, P3_U6847, P3_U6848, P3_U6849, P3_U6850, P3_U6851, P3_U6852, P3_U6853, P3_U6854, P3_U6855, P3_U6856, P3_U6857, P3_U6858, P3_U6859, P3_U6860, P3_U6861, P3_U6862, P3_U6863, P3_U6864, P3_U6865, P3_U6866, P3_U6867, P3_U6868, P3_U6869, P3_U6870, P3_U6871, P3_U6872, P3_U6873, P3_U6874, P3_U6875, P3_U6876, P3_U6877, P3_U6878, P3_U6879, P3_U6880, P3_U6881, P3_U6882, P3_U6883, P3_U6884, P3_U6885, P3_U6886, P3_U6887, P3_U6888, P3_U6889, P3_U6890, P3_U6891, P3_U6892, P3_U6893, P3_U6894, P3_U6895, P3_U6896, P3_U6897, P3_U6898, P3_U6899, P3_U6900, P3_U6901, P3_U6902, P3_U6903, P3_U6904, P3_U6905, P3_U6906, P3_U6907, P3_U6908, P3_U6909, P3_U6910, P3_U6911, P3_U6912, P3_U6913, P3_U6914, P3_U6915, P3_U6916, P3_U6917, P3_U6918, P3_U6919, P3_U6920, P3_U6921, P3_U6922, P3_U6923, P3_U6924, P3_U6925, P3_U6926, P3_U6927, P3_U6928, P3_U6929, P3_U6930, P3_U6931, P3_U6932, P3_U6933, P3_U6934, P3_U6935, P3_U6936, P3_U6937, P3_U6938, P3_U6939, P3_U6940, P3_U6941, P3_U6942, P3_U6943, P3_U6944, P3_U6945, P3_U6946, P3_U6947, P3_U6948, P3_U6949, P3_U6950, P3_U6951, P3_U6952, P3_U6953, P3_U6954, P3_U6955, P3_U6956, P3_U6957, P3_U6958, P3_U6959, P3_U6960, P3_U6961, P3_U6962, P3_U6963, P3_U6964, P3_U6965, P3_U6966, P3_U6967, P3_U6968, P3_U6969, P3_U6970, P3_U6971, P3_U6972, P3_U6973, P3_U6974, P3_U6975, P3_U6976, P3_U6977, P3_U6978, P3_U6979, P3_U6980, P3_U6981, P3_U6982, P3_U6983, P3_U6984, P3_U6985, P3_U6986, P3_U6987, P3_U6988, P3_U6989, P3_U6990, P3_U6991, P3_U6992, P3_U6993, P3_U6994, P3_U6995, P3_U6996, P3_U6997, P3_U6998, P3_U6999, P3_U7000, P3_U7001, P3_U7002, P3_U7003, P3_U7004, P3_U7005, P3_U7006, P3_U7007, P3_U7008, P3_U7009, P3_U7010, P3_U7011, P3_U7012, P3_U7013, P3_U7014, P3_U7015, P3_U7016, P3_U7017, P3_U7018, P3_U7019, P3_U7020, P3_U7021, P3_U7022, P3_U7023, P3_U7024, P3_U7025, P3_U7026, P3_U7027, P3_U7028, P3_U7029, P3_U7030, P3_U7031, P3_U7032, P3_U7033, P3_U7034, P3_U7035, P3_U7036, P3_U7037, P3_U7038, P3_U7039, P3_U7040, P3_U7041, P3_U7042, P3_U7043, P3_U7044, P3_U7045, P3_U7046, P3_U7047, P3_U7048, P3_U7049, P3_U7050, P3_U7051, P3_U7052, P3_U7053, P3_U7054, P3_U7055, P3_U7056, P3_U7057, P3_U7058, P3_U7059, P3_U7060, P3_U7061, P3_U7062, P3_U7063, P3_U7064, P3_U7065, P3_U7066, P3_U7067, P3_U7068, P3_U7069, P3_U7070, P3_U7071, P3_U7072, P3_U7073, P3_U7074, P3_U7075, P3_U7076, P3_U7077, P3_U7078, P3_U7079, P3_U7080, P3_U7081, P3_U7082, P3_U7083, P3_U7084, P3_U7085, P3_U7086, P3_U7087, P3_U7088, P3_U7089, P3_U7090, P3_U7091, P3_U7092, P3_U7093, P3_U7094, P3_U7095, P3_U7096, P3_U7097, P3_U7098, P3_U7099, P3_U7100, P3_U7101, P3_U7102, P3_U7103, P3_U7104, P3_U7105, P3_U7106, P3_U7107, P3_U7108, P3_U7109, P3_U7110, P3_U7111, P3_U7112, P3_U7113, P3_U7114, P3_U7115, P3_U7116, P3_U7117, P3_U7118, P3_U7119, P3_U7120, P3_U7121, P3_U7122, P3_U7123, P3_U7124, P3_U7125, P3_U7126, P3_U7127, P3_U7128, P3_U7129, P3_U7130, P3_U7131, P3_U7132, P3_U7133, P3_U7134, P3_U7135, P3_U7136, P3_U7137, P3_U7138, P3_U7139, P3_U7140, P3_U7141, P3_U7142, P3_U7143, P3_U7144, P3_U7145, P3_U7146, P3_U7147, P3_U7148, P3_U7149, P3_U7150, P3_U7151, P3_U7152, P3_U7153, P3_U7154, P3_U7155, P3_U7156, P3_U7157, P3_U7158, P3_U7159, P3_U7160, P3_U7161, P3_U7162, P3_U7163, P3_U7164, P3_U7165, P3_U7166, P3_U7167, P3_U7168, P3_U7169, P3_U7170, P3_U7171, P3_U7172, P3_U7173, P3_U7174, P3_U7175, P3_U7176, P3_U7177, P3_U7178, P3_U7179, P3_U7180, P3_U7181, P3_U7182, P3_U7183, P3_U7184, P3_U7185, P3_U7186, P3_U7187, P3_U7188, P3_U7189, P3_U7190, P3_U7191, P3_U7192, P3_U7193, P3_U7194, P3_U7195, P3_U7196, P3_U7197, P3_U7198, P3_U7199, P3_U7200, P3_U7201, P3_U7202, P3_U7203, P3_U7204, P3_U7205, P3_U7206, P3_U7207, P3_U7208, P3_U7209, P3_U7210, P3_U7211, P3_U7212, P3_U7213, P3_U7214, P3_U7215, P3_U7216, P3_U7217, P3_U7218, P3_U7219, P3_U7220, P3_U7221, P3_U7222, P3_U7223, P3_U7224, P3_U7225, P3_U7226, P3_U7227, P3_U7228, P3_U7229, P3_U7230, P3_U7231, P3_U7232, P3_U7233, P3_U7234, P3_U7235, P3_U7236, P3_U7237, P3_U7238, P3_U7239, P3_U7240, P3_U7241, P3_U7242, P3_U7243, P3_U7244, P3_U7245, P3_U7246, P3_U7247, P3_U7248, P3_U7249, P3_U7250, P3_U7251, P3_U7252, P3_U7253, P3_U7254, P3_U7255, P3_U7256, P3_U7257, P3_U7258, P3_U7259, P3_U7260, P3_U7261, P3_U7262, P3_U7263, P3_U7264, P3_U7265, P3_U7266, P3_U7267, P3_U7268, P3_U7269, P3_U7270, P3_U7271, P3_U7272, P3_U7273, P3_U7274, P3_U7275, P3_U7276, P3_U7277, P3_U7278, P3_U7279, P3_U7280, P3_U7281, P3_U7282, P3_U7283, P3_U7284, P3_U7285, P3_U7286, P3_U7287, P3_U7288, P3_U7289, P3_U7290, P3_U7291, P3_U7292, P3_U7293, P3_U7294, P3_U7295, P3_U7296, P3_U7297, P3_U7298, P3_U7299, P3_U7300, P3_U7301, P3_U7302, P3_U7303, P3_U7304, P3_U7305, P3_U7306, P3_U7307, P3_U7308, P3_U7309, P3_U7310, P3_U7311, P3_U7312, P3_U7313, P3_U7314, P3_U7315, P3_U7316, P3_U7317, P3_U7318, P3_U7319, P3_U7320, P3_U7321, P3_U7322, P3_U7323, P3_U7324, P3_U7325, P3_U7326, P3_U7327, P3_U7328, P3_U7329, P3_U7330, P3_U7331, P3_U7332, P3_U7333, P3_U7334, P3_U7335, P3_U7336, P3_U7337, P3_U7338, P3_U7339, P3_U7340, P3_U7341, P3_U7342, P3_U7343, P3_U7344, P3_U7345, P3_U7346, P3_U7347, P3_U7348, P3_U7349, P3_U7350, P3_U7351, P3_U7352, P3_U7353, P3_U7354, P3_U7355, P3_U7356, P3_U7357, P3_U7358, P3_U7359, P3_U7360, P3_U7361, P3_U7362, P3_U7363, P3_U7364, P3_U7365, P3_U7366, P3_U7367, P3_U7368, P3_U7369, P3_U7370, P3_U7371, P3_U7372, P3_U7373, P3_U7374, P3_U7375, P3_U7376, P3_U7377, P3_U7378, P3_U7379, P3_U7380, P3_U7381, P3_U7382, P3_U7383, P3_U7384, P3_U7385, P3_U7386, P3_U7387, P3_U7388, P3_U7389, P3_U7390, P3_U7391, P3_U7392, P3_U7393, P3_U7394, P3_U7395, P3_U7396, P3_U7397, P3_U7398, P3_U7399, P3_U7400, P3_U7401, P3_U7402, P3_U7403, P3_U7404, P3_U7405, P3_U7406, P3_U7407, P3_U7408, P3_U7409, P3_U7410, P3_U7411, P3_U7412, P3_U7413, P3_U7414, P3_U7415, P3_U7416, P3_U7417, P3_U7418, P3_U7419, P3_U7420, P3_U7421, P3_U7422, P3_U7423, P3_U7424, P3_U7425, P3_U7426, P3_U7427, P3_U7428, P3_U7429, P3_U7430, P3_U7431, P3_U7432, P3_U7433, P3_U7434, P3_U7435, P3_U7436, P3_U7437, P3_U7438, P3_U7439, P3_U7440, P3_U7441, P3_U7442, P3_U7443, P3_U7444, P3_U7445, P3_U7446, P3_U7447, P3_U7448, P3_U7449, P3_U7450, P3_U7451, P3_U7452, P3_U7453, P3_U7454, P3_U7455, P3_U7456, P3_U7457, P3_U7458, P3_U7459, P3_U7460, P3_U7461, P3_U7462, P3_U7463, P3_U7464, P3_U7465, P3_U7466, P3_U7467, P3_U7468, P3_U7469, P3_U7470, P3_U7471, P3_U7472, P3_U7473, P3_U7474, P3_U7475, P3_U7476, P3_U7477, P3_U7478, P3_U7479, P3_U7480, P3_U7481, P3_U7482, P3_U7483, P3_U7484, P3_U7485, P3_U7486, P3_U7487, P3_U7488, P3_U7489, P3_U7490, P3_U7491, P3_U7492, P3_U7493, P3_U7494, P3_U7495, P3_U7496, P3_U7497, P3_U7498, P3_U7499, P3_U7500, P3_U7501, P3_U7502, P3_U7503, P3_U7504, P3_U7505, P3_U7506, P3_U7507, P3_U7508, P3_U7509, P3_U7510, P3_U7511, P3_U7512, P3_U7513, P3_U7514, P3_U7515, P3_U7516, P3_U7517, P3_U7518, P3_U7519, P3_U7520, P3_U7521, P3_U7522, P3_U7523, P3_U7524, P3_U7525, P3_U7526, P3_U7527, P3_U7528, P3_U7529, P3_U7530, P3_U7531, P3_U7532, P3_U7533, P3_U7534, P3_U7535, P3_U7536, P3_U7537, P3_U7538, P3_U7539, P3_U7540, P3_U7541, P3_U7542, P3_U7543, P3_U7544, P3_U7545, P3_U7546, P3_U7547, P3_U7548, P3_U7549, P3_U7550, P3_U7551, P3_U7552, P3_U7553, P3_U7554, P3_U7555, P3_U7556, P3_U7557, P3_U7558, P3_U7559, P3_U7560, P3_U7561, P3_U7562, P3_U7563, P3_U7564, P3_U7565, P3_U7566, P3_U7567, P3_U7568, P3_U7569, P3_U7570, P3_U7571, P3_U7572, P3_U7573, P3_U7574, P3_U7575, P3_U7576, P3_U7577, P3_U7578, P3_U7579, P3_U7580, P3_U7581, P3_U7582, P3_U7583, P3_U7584, P3_U7585, P3_U7586, P3_U7587, P3_U7588, P3_U7589, P3_U7590, P3_U7591, P3_U7592, P3_U7593, P3_U7594, P3_U7595, P3_U7596, P3_U7597, P3_U7598, P3_U7599, P3_U7600, P3_U7601, P3_U7602, P3_U7603, P3_U7604, P3_U7605, P3_U7606, P3_U7607, P3_U7608, P3_U7609, P3_U7610, P3_U7611, P3_U7612, P3_U7613, P3_U7614, P3_U7615, P3_U7616, P3_U7617, P3_U7618, P3_U7619, P3_U7620, P3_U7621, P3_U7622, P3_U7623, P3_U7624, P3_U7625, P3_U7626, P3_U7627, P3_U7628, P3_U7629, P3_U7630, P3_U7631, P3_U7632, P3_U7633, P3_U7634, P3_U7635, P3_U7636, P3_U7637, P3_U7638, P3_U7639, P3_U7640, P3_U7641, P3_U7642, P3_U7643, P3_U7644, P3_U7645, P3_U7646, P3_U7647, P3_U7648, P3_U7649, P3_U7650, P3_U7651, P3_U7652, P3_U7653, P3_U7654, P3_U7655, P3_U7656, P3_U7657, P3_U7658, P3_U7659, P3_U7660, P3_U7661, P3_U7662, P3_U7663, P3_U7664, P3_U7665, P3_U7666, P3_U7667, P3_U7668, P3_U7669, P3_U7670, P3_U7671, P3_U7672, P3_U7673, P3_U7674, P3_U7675, P3_U7676, P3_U7677, P3_U7678, P3_U7679, P3_U7680, P3_U7681, P3_U7682, P3_U7683, P3_U7684, P3_U7685, P3_U7686, P3_U7687, P3_U7688, P3_U7689, P3_U7690, P3_U7691, P3_U7692, P3_U7693, P3_U7694, P3_U7695, P3_U7696, P3_U7697, P3_U7698, P3_U7699, P3_U7700, P3_U7701, P3_U7702, P3_U7703, P3_U7704, P3_U7705, P3_U7706, P3_U7707, P3_U7708, P3_U7709, P3_U7710, P3_U7711, P3_U7712, P3_U7713, P3_U7714, P3_U7715, P3_U7716, P3_U7717, P3_U7718, P3_U7719, P3_U7720, P3_U7721, P3_U7722, P3_U7723, P3_U7724, P3_U7725, P3_U7726, P3_U7727, P3_U7728, P3_U7729, P3_U7730, P3_U7731, P3_U7732, P3_U7733, P3_U7734, P3_U7735, P3_U7736, P3_U7737, P3_U7738, P3_U7739, P3_U7740, P3_U7741, P3_U7742, P3_U7743, P3_U7744, P3_U7745, P3_U7746, P3_U7747, P3_U7748, P3_U7749, P3_U7750, P3_U7751, P3_U7752, P3_U7753, P3_U7754, P3_U7755, P3_U7756, P3_U7757, P3_U7758, P3_U7759, P3_U7760, P3_U7761, P3_U7762, P3_U7763, P3_U7764, P3_U7765, P3_U7766, P3_U7767, P3_U7768, P3_U7769, P3_U7770, P3_U7771, P3_U7772, P3_U7773, P3_U7774, P3_U7775, P3_U7776, P3_U7777, P3_U7778, P3_U7779, P3_U7780, P3_U7781, P3_U7782, P3_U7783, P3_U7784, P3_U7785, P3_U7786, P3_U7787, P3_U7788, P3_U7789, P3_U7790, P3_U7791, P3_U7792, P3_U7793, P3_U7794, P3_U7795, P3_U7796, P3_U7797, P3_U7798, P3_U7799, P3_U7800, P3_U7801, P3_U7802, P3_U7803, P3_U7804, P3_U7805, P3_U7806, P3_U7807, P3_U7808, P3_U7809, P3_U7810, P3_U7811, P3_U7812, P3_U7813, P3_U7814, P3_U7815, P3_U7816, P3_U7817, P3_U7818, P3_U7819, P3_U7820, P3_U7821, P3_U7822, P3_U7823, P3_U7824, P3_U7825, P3_U7826, P3_U7827, P3_U7828, P3_U7829, P3_U7830, P3_U7831, P3_U7832, P3_U7833, P3_U7834, P3_U7835, P3_U7836, P3_U7837, P3_U7838, P3_U7839, P3_U7840, P3_U7841, P3_U7842, P3_U7843, P3_U7844, P3_U7845, P3_U7846, P3_U7847, P3_U7848, P3_U7849, P3_U7850, P3_U7851, P3_U7852, P3_U7853, P3_U7854, P3_U7855, P3_U7856, P3_U7857, P3_U7858, P3_U7859, P3_U7860, P3_U7861, P3_U7862, P3_U7863, P3_U7864, P3_U7865, P3_U7866, P3_U7867, P3_U7868, P3_U7869, P3_U7870, P3_U7871, P3_U7872, P3_U7873, P3_U7874, P3_U7875, P3_U7876, P3_U7877, P3_U7878, P3_U7879, P3_U7880, P3_U7881, P3_U7882, P3_U7883, P3_U7884, P3_U7885, P3_U7886, P3_U7887, P3_U7888, P3_U7889, P3_U7890, P3_U7891, P3_U7892, P3_U7893, P3_U7894, P3_U7895, P3_U7896, P3_U7897, P3_U7898, P3_U7899, P3_U7900, P3_U7901, P3_U7902, P3_U7903, P3_U7904, P3_U7905, P3_U7906, P3_U7907, P3_U7908, P3_U7909, P3_U7910, P3_U7911, P3_U7912, P3_U7913, P3_U7914, P3_U7915, P3_U7916, P3_U7917, P3_U7918, P3_U7919, P3_U7920, P3_U7921, P3_U7922, P3_U7923, P3_U7924, P3_U7925, P3_U7926, P3_U7927, P3_U7928, P3_U7929, P3_U7930, P3_U7931, P3_U7932, P3_U7933, P3_U7934, P3_U7935, P3_U7936, P3_U7937, P3_U7938, P3_U7939, P3_U7940, P3_U7941, P3_U7942, P3_U7943, P3_U7944, P3_U7945, P3_U7946, P3_U7947, P3_U7948, P3_U7949, P3_U7950, P3_U7951, P3_U7952, P3_U7953, P3_U7954, P3_U7955, P3_U7956, P3_U7957, P3_U7958, P3_U7959, P3_U7960, P3_U7961, P3_U7962, P3_U7963, P3_U7964, P3_U7965, P3_U7966, P3_U7967, P3_U7968, P3_U7969, P3_U7970, P3_U7971, P3_U7972, P3_U7973, P3_U7974, P3_U7975, P3_U7976, P3_U7977, P3_U7978, P3_U7979, P3_U7980, P3_U7981, P3_U7982, P3_U7983, P3_U7984, P3_U7985, P3_U7986, P3_U7987, P3_U7988, P3_U7989, P3_U7990, P3_U7991, P3_U7992, P3_U7993, P3_U7994, P3_U7995, P3_U7996, P3_U7997, P3_U7998, P3_U7999, P3_U8000, P3_U8001, P3_U8002, P3_U8003, P3_U8004, P3_U8005, P3_U8006, P3_U8007, P3_U8008, P3_U8009, P3_U8010, P3_U8011, P3_U8012, P3_U8013, P3_U8014, P3_U8015, P3_U8016, P3_U8017, P3_U8018, P3_U8019, P3_U8020, P3_U8021, P3_U8022, P3_U8023, P3_U8024, P3_U8025, P3_U8026, P3_U8027, P3_U8028, P3_U8029, P3_U8030, P3_U8031, P3_U8032, P3_U8033, P3_U8034, P3_U8035, P3_U8036, P3_U8037, P3_U8038, P3_U8039, P3_U8040, P3_U8041, P3_U8042, P3_U8043, P3_U8044, P3_U8045, P3_U8046, P3_U8047, P3_U8048, P3_U8049, P3_U8050, P3_U8051, P3_U8052, P3_U8053, R165_U10, R165_U11, R165_U12, R165_U13, R165_U14, R165_U15, R165_U6, R165_U7, R165_U8, R165_U9, R170_U10, R170_U11, R170_U12, R170_U13, R170_U14, R170_U15, R170_U6, R170_U7, R170_U8, R170_U9, U207, U208, U209, U210, U211, U248, U249, U250, U283, U284, U285, U286, U287, U288, U289, U290, U291, U292, U293, U294, U295, U296, U297, U298, U299, U300, U301, U302, U303, U304, U305, U306, U307, U308, U309, U310, U311, U312, U313, U314, U315, U316, U317, U318, U319, U320, U321, U322, U323, U324, U325, U326, U327, U328, U329, U330, U331, U332, U333, U334, U335, U336, U337, U338, U339, U340, U341, U342, U343, U344, U345, U346, U377, U378, U379, U380, U381, U382, U383, U384, U385, U386, U387, U388, U389, U390, U391, U392, U393, U394, U395, U396, U397, U398, U399, U400, U401, U402, U403, U404, U405, U406, U407, U408, U409, U410, U411, U412, U413, U414, U415, U416, U417, U418, U419, U420, U421, U422, U423, U424, U425, U426, U427, U428, U429, U430, U431, U432, U433, U434, U435, U436, U437, U438, U439, U440, U441, U442, U443, U444, U445, U446, U447, U448, U449, U450, U451, U452, U453, U454, U455, U456, U457, U458, U459, U460, U461, U462, U463, U464, U465, U466, U467, U468, U469, U470, U471, U472, U473, U474, U475, U476, U477, U478, U479, U480, U481, U482, U483, U484, U485, U486, U487, U488, U489, U490, U491, U492, U493, U494, U495, U496, U497, U498, U499, U500, U501, U502, U503, U504, U505, U506, U507, U508, U509, U510, U511, U512, U513, U514, U515, U516, U517, U518, U519, U520, U521, U522, U523, U524, U525, U526, U527, U528, U529, U530, U531, U532, U533, U534, U535, U536, U537, U538, U539, U540, U541, U542, U543, U544, U545, U546, U547, U548, U549, U550, U551, U552, U553, U554, U555, U556, U557, U558, U559, U560, U561, U562, U563, U564, U565, U566, U567, U568, U569, U570, U571, U572, U573, U574, U575, U576, U577, U578, U579, U580, U581, U582, U583, U584, U585, U586, U587, U588, U589, U590, U591, U592, U593, U594, U595, U596, U597, U598, U599, U600, U601, U602, U603, U604, U605, U606, U607, U608, U609, U610, U611, U612, U613, U614, U615, U616, U617, U618, U619, U620, U621, U622, U623, U624, U625, U626, U627, U628, U629, U630, U631, U632, U633, U634, U635, U636, U637, U638, U639, U640, U641, U642, U643, U644, U645, U646, U647, U648, U649, U650, U651, U652, U653, U654, U655, U656, U657, U658, U659, U660, U661, U662, U663, U664, U665, U666, U667, U668, U669, U670, U671, U672, U673, U674, U675, U676, U677, U678, U679, U680, U681, U682, U683, U684, U685, U686, U687, U688, U689, U690, U691, U692, U693, U694, U695, U696, U697, U698, U699, U700, U701, U702, U703, U704, U705, U706, U707, U708, U709, U710, U711, U712, U713, U714, U715, U716, U717, U718, U719, U720, U721, U722, U723, U724, U725, U726, U727, U728, U729, U730, U731, U732, U733, U734, U735, U736, P1_U3149_in, flip_signal;

  not ginst1 (LT_748_U6, P2_ADDRESS_REG_29__SCAN_IN);
  nand ginst2 (LT_782_119_U6, P2_DATAO_REG_30__SCAN_IN, LT_782_119_U7);
  not ginst3 (LT_782_119_U7, P2_DATAO_REG_31__SCAN_IN);
  nand ginst4 (LT_782_120_U6, P3_DATAO_REG_30__SCAN_IN, LT_782_120_U7);
  not ginst5 (LT_782_120_U7, P3_DATAO_REG_31__SCAN_IN);
  nand ginst6 (LT_782_U6, P1_DATAO_REG_30__SCAN_IN, LT_782_U7);
  not ginst7 (LT_782_U7, P1_DATAO_REG_31__SCAN_IN);
  not ginst8 (P1_ADD_371_U10, P1_U3231);
  nand ginst9 (P1_ADD_371_U11, P1_ADD_371_U28, P1_U3231);
  not ginst10 (P1_ADD_371_U12, P1_U3232);
  not ginst11 (P1_ADD_371_U13, P1_U3233);
  nand ginst12 (P1_ADD_371_U14, P1_ADD_371_U29, P1_U3232);
  not ginst13 (P1_ADD_371_U15, P1_U3229);
  not ginst14 (P1_ADD_371_U16, P1_U3234);
  nand ginst15 (P1_ADD_371_U17, P1_ADD_371_U33, P1_ADD_371_U34);
  nand ginst16 (P1_ADD_371_U18, P1_ADD_371_U35, P1_ADD_371_U36);
  nand ginst17 (P1_ADD_371_U19, P1_ADD_371_U37, P1_ADD_371_U38);
  nand ginst18 (P1_ADD_371_U20, P1_ADD_371_U41, P1_ADD_371_U42);
  nand ginst19 (P1_ADD_371_U21, P1_ADD_371_U43, P1_ADD_371_U44);
  and ginst20 (P1_ADD_371_U22, P1_U3233, P1_U3234);
  nand ginst21 (P1_ADD_371_U23, P1_ADD_371_U15, P1_ADD_371_U26);
  and ginst22 (P1_ADD_371_U24, P1_ADD_371_U39, P1_ADD_371_U40);
  nand ginst23 (P1_ADD_371_U25, P1_ADD_371_U30, P1_U3233);
  nand ginst24 (P1_ADD_371_U26, P1_U3227, P1_U3228);
  not ginst25 (P1_ADD_371_U27, P1_ADD_371_U23);
  not ginst26 (P1_ADD_371_U28, P1_ADD_371_U9);
  not ginst27 (P1_ADD_371_U29, P1_ADD_371_U11);
  not ginst28 (P1_ADD_371_U30, P1_ADD_371_U14);
  nand ginst29 (P1_ADD_371_U31, P1_U3227, P1_U3228, P1_U3229);
  not ginst30 (P1_ADD_371_U32, P1_ADD_371_U25);
  nand ginst31 (P1_ADD_371_U33, P1_ADD_371_U14, P1_U3233);
  nand ginst32 (P1_ADD_371_U34, P1_ADD_371_U13, P1_ADD_371_U30);
  nand ginst33 (P1_ADD_371_U35, P1_ADD_371_U9, P1_U3231);
  nand ginst34 (P1_ADD_371_U36, P1_ADD_371_U10, P1_ADD_371_U28);
  nand ginst35 (P1_ADD_371_U37, P1_ADD_371_U11, P1_U3232);
  nand ginst36 (P1_ADD_371_U38, P1_ADD_371_U12, P1_ADD_371_U29);
  nand ginst37 (P1_ADD_371_U39, P1_ADD_371_U23, P1_U3230);
  not ginst38 (P1_ADD_371_U4, P1_U3227);
  nand ginst39 (P1_ADD_371_U40, P1_ADD_371_U27, P1_ADD_371_U8);
  nand ginst40 (P1_ADD_371_U41, P1_ADD_371_U4, P1_U3228);
  nand ginst41 (P1_ADD_371_U42, P1_ADD_371_U7, P1_U3227);
  nand ginst42 (P1_ADD_371_U43, P1_ADD_371_U25, P1_U3234);
  nand ginst43 (P1_ADD_371_U44, P1_ADD_371_U16, P1_ADD_371_U32);
  nand ginst44 (P1_ADD_371_U5, P1_ADD_371_U23, P1_ADD_371_U31);
  and ginst45 (P1_ADD_371_U6, P1_ADD_371_U22, P1_ADD_371_U30);
  not ginst46 (P1_ADD_371_U7, P1_U3228);
  not ginst47 (P1_ADD_371_U8, P1_U3230);
  nand ginst48 (P1_ADD_371_U9, P1_ADD_371_U23, P1_U3230);
  nand ginst49 (P1_ADD_405_U10, P1_INSTADDRPOINTER_REG_4__SCAN_IN, P1_ADD_405_U98);
  not ginst50 (P1_ADD_405_U100, P1_ADD_405_U13);
  not ginst51 (P1_ADD_405_U101, P1_ADD_405_U14);
  not ginst52 (P1_ADD_405_U102, P1_ADD_405_U16);
  not ginst53 (P1_ADD_405_U103, P1_ADD_405_U18);
  not ginst54 (P1_ADD_405_U104, P1_ADD_405_U20);
  not ginst55 (P1_ADD_405_U105, P1_ADD_405_U22);
  not ginst56 (P1_ADD_405_U106, P1_ADD_405_U24);
  not ginst57 (P1_ADD_405_U107, P1_ADD_405_U26);
  not ginst58 (P1_ADD_405_U108, P1_ADD_405_U28);
  not ginst59 (P1_ADD_405_U109, P1_ADD_405_U30);
  not ginst60 (P1_ADD_405_U11, P1_INSTADDRPOINTER_REG_5__SCAN_IN);
  not ginst61 (P1_ADD_405_U110, P1_ADD_405_U32);
  not ginst62 (P1_ADD_405_U111, P1_ADD_405_U34);
  not ginst63 (P1_ADD_405_U112, P1_ADD_405_U36);
  not ginst64 (P1_ADD_405_U113, P1_ADD_405_U38);
  not ginst65 (P1_ADD_405_U114, P1_ADD_405_U40);
  not ginst66 (P1_ADD_405_U115, P1_ADD_405_U42);
  not ginst67 (P1_ADD_405_U116, P1_ADD_405_U44);
  not ginst68 (P1_ADD_405_U117, P1_ADD_405_U46);
  not ginst69 (P1_ADD_405_U118, P1_ADD_405_U48);
  not ginst70 (P1_ADD_405_U119, P1_ADD_405_U50);
  not ginst71 (P1_ADD_405_U12, P1_INSTADDRPOINTER_REG_6__SCAN_IN);
  not ginst72 (P1_ADD_405_U120, P1_ADD_405_U52);
  not ginst73 (P1_ADD_405_U121, P1_ADD_405_U54);
  not ginst74 (P1_ADD_405_U122, P1_ADD_405_U56);
  not ginst75 (P1_ADD_405_U123, P1_ADD_405_U58);
  not ginst76 (P1_ADD_405_U124, P1_ADD_405_U61);
  nand ginst77 (P1_ADD_405_U125, P1_INSTADDRPOINTER_REG_2__SCAN_IN, P1_INSTADDRPOINTER_REG_1__SCAN_IN, P1_INSTADDRPOINTER_REG_0__SCAN_IN);
  not ginst78 (P1_ADD_405_U126, P1_ADD_405_U93);
  nand ginst79 (P1_ADD_405_U127, P1_INSTADDRPOINTER_REG_6__SCAN_IN, P1_ADD_405_U13);
  nand ginst80 (P1_ADD_405_U128, P1_ADD_405_U100, P1_ADD_405_U12);
  nand ginst81 (P1_ADD_405_U129, P1_INSTADDRPOINTER_REG_30__SCAN_IN, P1_ADD_405_U61);
  nand ginst82 (P1_ADD_405_U13, P1_INSTADDRPOINTER_REG_5__SCAN_IN, P1_ADD_405_U99);
  nand ginst83 (P1_ADD_405_U130, P1_ADD_405_U124, P1_ADD_405_U60);
  nand ginst84 (P1_ADD_405_U131, P1_INSTADDRPOINTER_REG_29__SCAN_IN, P1_ADD_405_U58);
  nand ginst85 (P1_ADD_405_U132, P1_ADD_405_U123, P1_ADD_405_U59);
  nand ginst86 (P1_ADD_405_U133, P1_INSTADDRPOINTER_REG_24__SCAN_IN, P1_ADD_405_U48);
  nand ginst87 (P1_ADD_405_U134, P1_ADD_405_U118, P1_ADD_405_U49);
  nand ginst88 (P1_ADD_405_U135, P1_INSTADDRPOINTER_REG_17__SCAN_IN, P1_ADD_405_U34);
  nand ginst89 (P1_ADD_405_U136, P1_ADD_405_U111, P1_ADD_405_U35);
  nand ginst90 (P1_ADD_405_U137, P1_INSTADDRPOINTER_REG_20__SCAN_IN, P1_ADD_405_U40);
  nand ginst91 (P1_ADD_405_U138, P1_ADD_405_U114, P1_ADD_405_U41);
  nand ginst92 (P1_ADD_405_U139, P1_INSTADDRPOINTER_REG_13__SCAN_IN, P1_ADD_405_U26);
  nand ginst93 (P1_ADD_405_U14, P1_INSTADDRPOINTER_REG_6__SCAN_IN, P1_ADD_405_U100);
  nand ginst94 (P1_ADD_405_U140, P1_ADD_405_U107, P1_ADD_405_U27);
  nand ginst95 (P1_ADD_405_U141, P1_INSTADDRPOINTER_REG_9__SCAN_IN, P1_ADD_405_U18);
  nand ginst96 (P1_ADD_405_U142, P1_ADD_405_U103, P1_ADD_405_U19);
  nand ginst97 (P1_ADD_405_U143, P1_INSTADDRPOINTER_REG_22__SCAN_IN, P1_ADD_405_U44);
  nand ginst98 (P1_ADD_405_U144, P1_ADD_405_U116, P1_ADD_405_U45);
  nand ginst99 (P1_ADD_405_U145, P1_INSTADDRPOINTER_REG_18__SCAN_IN, P1_ADD_405_U36);
  nand ginst100 (P1_ADD_405_U146, P1_ADD_405_U112, P1_ADD_405_U37);
  nand ginst101 (P1_ADD_405_U147, P1_INSTADDRPOINTER_REG_11__SCAN_IN, P1_ADD_405_U22);
  nand ginst102 (P1_ADD_405_U148, P1_ADD_405_U105, P1_ADD_405_U23);
  nand ginst103 (P1_ADD_405_U149, P1_INSTADDRPOINTER_REG_26__SCAN_IN, P1_ADD_405_U52);
  not ginst104 (P1_ADD_405_U15, P1_INSTADDRPOINTER_REG_7__SCAN_IN);
  nand ginst105 (P1_ADD_405_U150, P1_ADD_405_U120, P1_ADD_405_U53);
  nand ginst106 (P1_ADD_405_U151, P1_INSTADDRPOINTER_REG_15__SCAN_IN, P1_ADD_405_U30);
  nand ginst107 (P1_ADD_405_U152, P1_ADD_405_U109, P1_ADD_405_U31);
  nand ginst108 (P1_ADD_405_U153, P1_INSTADDRPOINTER_REG_4__SCAN_IN, P1_ADD_405_U8);
  nand ginst109 (P1_ADD_405_U154, P1_ADD_405_U9, P1_ADD_405_U98);
  nand ginst110 (P1_ADD_405_U155, P1_INSTADDRPOINTER_REG_27__SCAN_IN, P1_ADD_405_U54);
  nand ginst111 (P1_ADD_405_U156, P1_ADD_405_U121, P1_ADD_405_U55);
  nand ginst112 (P1_ADD_405_U157, P1_INSTADDRPOINTER_REG_14__SCAN_IN, P1_ADD_405_U28);
  nand ginst113 (P1_ADD_405_U158, P1_ADD_405_U108, P1_ADD_405_U29);
  nand ginst114 (P1_ADD_405_U159, P1_INSTADDRPOINTER_REG_5__SCAN_IN, P1_ADD_405_U10);
  nand ginst115 (P1_ADD_405_U16, P1_INSTADDRPOINTER_REG_7__SCAN_IN, P1_ADD_405_U101);
  nand ginst116 (P1_ADD_405_U160, P1_ADD_405_U11, P1_ADD_405_U99);
  nand ginst117 (P1_ADD_405_U161, P1_INSTADDRPOINTER_REG_8__SCAN_IN, P1_ADD_405_U16);
  nand ginst118 (P1_ADD_405_U162, P1_ADD_405_U102, P1_ADD_405_U17);
  nand ginst119 (P1_ADD_405_U163, P1_INSTADDRPOINTER_REG_23__SCAN_IN, P1_ADD_405_U46);
  nand ginst120 (P1_ADD_405_U164, P1_ADD_405_U117, P1_ADD_405_U47);
  nand ginst121 (P1_ADD_405_U165, P1_INSTADDRPOINTER_REG_19__SCAN_IN, P1_ADD_405_U38);
  nand ginst122 (P1_ADD_405_U166, P1_ADD_405_U113, P1_ADD_405_U39);
  nand ginst123 (P1_ADD_405_U167, P1_INSTADDRPOINTER_REG_10__SCAN_IN, P1_ADD_405_U20);
  nand ginst124 (P1_ADD_405_U168, P1_ADD_405_U104, P1_ADD_405_U21);
  nand ginst125 (P1_ADD_405_U169, P1_INSTADDRPOINTER_REG_31__SCAN_IN, P1_ADD_405_U93);
  not ginst126 (P1_ADD_405_U17, P1_INSTADDRPOINTER_REG_8__SCAN_IN);
  nand ginst127 (P1_ADD_405_U170, P1_ADD_405_U126, P1_ADD_405_U92);
  nand ginst128 (P1_ADD_405_U171, P1_INSTADDRPOINTER_REG_3__SCAN_IN, P1_ADD_405_U94);
  nand ginst129 (P1_ADD_405_U172, P1_ADD_405_U7, P1_ADD_405_U97);
  nand ginst130 (P1_ADD_405_U173, P1_INSTADDRPOINTER_REG_1__SCAN_IN, P1_ADD_405_U4);
  nand ginst131 (P1_ADD_405_U174, P1_INSTADDRPOINTER_REG_0__SCAN_IN, P1_ADD_405_U6);
  nand ginst132 (P1_ADD_405_U175, P1_INSTADDRPOINTER_REG_28__SCAN_IN, P1_ADD_405_U56);
  nand ginst133 (P1_ADD_405_U176, P1_ADD_405_U122, P1_ADD_405_U57);
  nand ginst134 (P1_ADD_405_U177, P1_INSTADDRPOINTER_REG_21__SCAN_IN, P1_ADD_405_U42);
  nand ginst135 (P1_ADD_405_U178, P1_ADD_405_U115, P1_ADD_405_U43);
  nand ginst136 (P1_ADD_405_U179, P1_INSTADDRPOINTER_REG_12__SCAN_IN, P1_ADD_405_U24);
  nand ginst137 (P1_ADD_405_U18, P1_INSTADDRPOINTER_REG_8__SCAN_IN, P1_ADD_405_U102);
  nand ginst138 (P1_ADD_405_U180, P1_ADD_405_U106, P1_ADD_405_U25);
  nand ginst139 (P1_ADD_405_U181, P1_INSTADDRPOINTER_REG_7__SCAN_IN, P1_ADD_405_U14);
  nand ginst140 (P1_ADD_405_U182, P1_ADD_405_U101, P1_ADD_405_U15);
  nand ginst141 (P1_ADD_405_U183, P1_INSTADDRPOINTER_REG_25__SCAN_IN, P1_ADD_405_U50);
  nand ginst142 (P1_ADD_405_U184, P1_ADD_405_U119, P1_ADD_405_U51);
  nand ginst143 (P1_ADD_405_U185, P1_INSTADDRPOINTER_REG_16__SCAN_IN, P1_ADD_405_U32);
  nand ginst144 (P1_ADD_405_U186, P1_ADD_405_U110, P1_ADD_405_U33);
  not ginst145 (P1_ADD_405_U19, P1_INSTADDRPOINTER_REG_9__SCAN_IN);
  nand ginst146 (P1_ADD_405_U20, P1_INSTADDRPOINTER_REG_9__SCAN_IN, P1_ADD_405_U103);
  not ginst147 (P1_ADD_405_U21, P1_INSTADDRPOINTER_REG_10__SCAN_IN);
  nand ginst148 (P1_ADD_405_U22, P1_INSTADDRPOINTER_REG_10__SCAN_IN, P1_ADD_405_U104);
  not ginst149 (P1_ADD_405_U23, P1_INSTADDRPOINTER_REG_11__SCAN_IN);
  nand ginst150 (P1_ADD_405_U24, P1_INSTADDRPOINTER_REG_11__SCAN_IN, P1_ADD_405_U105);
  not ginst151 (P1_ADD_405_U25, P1_INSTADDRPOINTER_REG_12__SCAN_IN);
  nand ginst152 (P1_ADD_405_U26, P1_INSTADDRPOINTER_REG_12__SCAN_IN, P1_ADD_405_U106);
  not ginst153 (P1_ADD_405_U27, P1_INSTADDRPOINTER_REG_13__SCAN_IN);
  nand ginst154 (P1_ADD_405_U28, P1_INSTADDRPOINTER_REG_13__SCAN_IN, P1_ADD_405_U107);
  not ginst155 (P1_ADD_405_U29, P1_INSTADDRPOINTER_REG_14__SCAN_IN);
  nand ginst156 (P1_ADD_405_U30, P1_INSTADDRPOINTER_REG_14__SCAN_IN, P1_ADD_405_U108);
  not ginst157 (P1_ADD_405_U31, P1_INSTADDRPOINTER_REG_15__SCAN_IN);
  nand ginst158 (P1_ADD_405_U32, P1_INSTADDRPOINTER_REG_15__SCAN_IN, P1_ADD_405_U109);
  not ginst159 (P1_ADD_405_U33, P1_INSTADDRPOINTER_REG_16__SCAN_IN);
  nand ginst160 (P1_ADD_405_U34, P1_INSTADDRPOINTER_REG_16__SCAN_IN, P1_ADD_405_U110);
  not ginst161 (P1_ADD_405_U35, P1_INSTADDRPOINTER_REG_17__SCAN_IN);
  nand ginst162 (P1_ADD_405_U36, P1_INSTADDRPOINTER_REG_17__SCAN_IN, P1_ADD_405_U111);
  not ginst163 (P1_ADD_405_U37, P1_INSTADDRPOINTER_REG_18__SCAN_IN);
  nand ginst164 (P1_ADD_405_U38, P1_INSTADDRPOINTER_REG_18__SCAN_IN, P1_ADD_405_U112);
  not ginst165 (P1_ADD_405_U39, P1_INSTADDRPOINTER_REG_19__SCAN_IN);
  not ginst166 (P1_ADD_405_U4, P1_INSTADDRPOINTER_REG_0__SCAN_IN);
  nand ginst167 (P1_ADD_405_U40, P1_INSTADDRPOINTER_REG_19__SCAN_IN, P1_ADD_405_U113);
  not ginst168 (P1_ADD_405_U41, P1_INSTADDRPOINTER_REG_20__SCAN_IN);
  nand ginst169 (P1_ADD_405_U42, P1_INSTADDRPOINTER_REG_20__SCAN_IN, P1_ADD_405_U114);
  not ginst170 (P1_ADD_405_U43, P1_INSTADDRPOINTER_REG_21__SCAN_IN);
  nand ginst171 (P1_ADD_405_U44, P1_INSTADDRPOINTER_REG_21__SCAN_IN, P1_ADD_405_U115);
  not ginst172 (P1_ADD_405_U45, P1_INSTADDRPOINTER_REG_22__SCAN_IN);
  nand ginst173 (P1_ADD_405_U46, P1_INSTADDRPOINTER_REG_22__SCAN_IN, P1_ADD_405_U116);
  not ginst174 (P1_ADD_405_U47, P1_INSTADDRPOINTER_REG_23__SCAN_IN);
  nand ginst175 (P1_ADD_405_U48, P1_INSTADDRPOINTER_REG_23__SCAN_IN, P1_ADD_405_U117);
  not ginst176 (P1_ADD_405_U49, P1_INSTADDRPOINTER_REG_24__SCAN_IN);
  nand ginst177 (P1_ADD_405_U5, P1_ADD_405_U125, P1_ADD_405_U94);
  nand ginst178 (P1_ADD_405_U50, P1_INSTADDRPOINTER_REG_24__SCAN_IN, P1_ADD_405_U118);
  not ginst179 (P1_ADD_405_U51, P1_INSTADDRPOINTER_REG_25__SCAN_IN);
  nand ginst180 (P1_ADD_405_U52, P1_INSTADDRPOINTER_REG_25__SCAN_IN, P1_ADD_405_U119);
  not ginst181 (P1_ADD_405_U53, P1_INSTADDRPOINTER_REG_26__SCAN_IN);
  nand ginst182 (P1_ADD_405_U54, P1_INSTADDRPOINTER_REG_26__SCAN_IN, P1_ADD_405_U120);
  not ginst183 (P1_ADD_405_U55, P1_INSTADDRPOINTER_REG_27__SCAN_IN);
  nand ginst184 (P1_ADD_405_U56, P1_INSTADDRPOINTER_REG_27__SCAN_IN, P1_ADD_405_U121);
  not ginst185 (P1_ADD_405_U57, P1_INSTADDRPOINTER_REG_28__SCAN_IN);
  nand ginst186 (P1_ADD_405_U58, P1_INSTADDRPOINTER_REG_28__SCAN_IN, P1_ADD_405_U122);
  not ginst187 (P1_ADD_405_U59, P1_INSTADDRPOINTER_REG_29__SCAN_IN);
  not ginst188 (P1_ADD_405_U6, P1_INSTADDRPOINTER_REG_1__SCAN_IN);
  not ginst189 (P1_ADD_405_U60, P1_INSTADDRPOINTER_REG_30__SCAN_IN);
  nand ginst190 (P1_ADD_405_U61, P1_INSTADDRPOINTER_REG_29__SCAN_IN, P1_ADD_405_U123);
  not ginst191 (P1_ADD_405_U62, P1_INSTADDRPOINTER_REG_2__SCAN_IN);
  nand ginst192 (P1_ADD_405_U63, P1_ADD_405_U127, P1_ADD_405_U128);
  nand ginst193 (P1_ADD_405_U64, P1_ADD_405_U129, P1_ADD_405_U130);
  nand ginst194 (P1_ADD_405_U65, P1_ADD_405_U131, P1_ADD_405_U132);
  nand ginst195 (P1_ADD_405_U66, P1_ADD_405_U133, P1_ADD_405_U134);
  nand ginst196 (P1_ADD_405_U67, P1_ADD_405_U135, P1_ADD_405_U136);
  nand ginst197 (P1_ADD_405_U68, P1_ADD_405_U137, P1_ADD_405_U138);
  nand ginst198 (P1_ADD_405_U69, P1_ADD_405_U139, P1_ADD_405_U140);
  not ginst199 (P1_ADD_405_U7, P1_INSTADDRPOINTER_REG_3__SCAN_IN);
  nand ginst200 (P1_ADD_405_U70, P1_ADD_405_U141, P1_ADD_405_U142);
  nand ginst201 (P1_ADD_405_U71, P1_ADD_405_U143, P1_ADD_405_U144);
  nand ginst202 (P1_ADD_405_U72, P1_ADD_405_U145, P1_ADD_405_U146);
  nand ginst203 (P1_ADD_405_U73, P1_ADD_405_U147, P1_ADD_405_U148);
  nand ginst204 (P1_ADD_405_U74, P1_ADD_405_U149, P1_ADD_405_U150);
  nand ginst205 (P1_ADD_405_U75, P1_ADD_405_U151, P1_ADD_405_U152);
  nand ginst206 (P1_ADD_405_U76, P1_ADD_405_U153, P1_ADD_405_U154);
  nand ginst207 (P1_ADD_405_U77, P1_ADD_405_U155, P1_ADD_405_U156);
  nand ginst208 (P1_ADD_405_U78, P1_ADD_405_U157, P1_ADD_405_U158);
  nand ginst209 (P1_ADD_405_U79, P1_ADD_405_U159, P1_ADD_405_U160);
  nand ginst210 (P1_ADD_405_U8, P1_INSTADDRPOINTER_REG_3__SCAN_IN, P1_ADD_405_U94);
  nand ginst211 (P1_ADD_405_U80, P1_ADD_405_U161, P1_ADD_405_U162);
  nand ginst212 (P1_ADD_405_U81, P1_ADD_405_U163, P1_ADD_405_U164);
  nand ginst213 (P1_ADD_405_U82, P1_ADD_405_U165, P1_ADD_405_U166);
  nand ginst214 (P1_ADD_405_U83, P1_ADD_405_U167, P1_ADD_405_U168);
  nand ginst215 (P1_ADD_405_U84, P1_ADD_405_U169, P1_ADD_405_U170);
  nand ginst216 (P1_ADD_405_U85, P1_ADD_405_U173, P1_ADD_405_U174);
  nand ginst217 (P1_ADD_405_U86, P1_ADD_405_U175, P1_ADD_405_U176);
  nand ginst218 (P1_ADD_405_U87, P1_ADD_405_U177, P1_ADD_405_U178);
  nand ginst219 (P1_ADD_405_U88, P1_ADD_405_U179, P1_ADD_405_U180);
  nand ginst220 (P1_ADD_405_U89, P1_ADD_405_U181, P1_ADD_405_U182);
  not ginst221 (P1_ADD_405_U9, P1_INSTADDRPOINTER_REG_4__SCAN_IN);
  nand ginst222 (P1_ADD_405_U90, P1_ADD_405_U183, P1_ADD_405_U184);
  nand ginst223 (P1_ADD_405_U91, P1_ADD_405_U185, P1_ADD_405_U186);
  not ginst224 (P1_ADD_405_U92, P1_INSTADDRPOINTER_REG_31__SCAN_IN);
  nand ginst225 (P1_ADD_405_U93, P1_INSTADDRPOINTER_REG_30__SCAN_IN, P1_ADD_405_U124);
  nand ginst226 (P1_ADD_405_U94, P1_ADD_405_U62, P1_ADD_405_U96);
  and ginst227 (P1_ADD_405_U95, P1_ADD_405_U171, P1_ADD_405_U172);
  nand ginst228 (P1_ADD_405_U96, P1_INSTADDRPOINTER_REG_1__SCAN_IN, P1_INSTADDRPOINTER_REG_0__SCAN_IN);
  not ginst229 (P1_ADD_405_U97, P1_ADD_405_U94);
  not ginst230 (P1_ADD_405_U98, P1_ADD_405_U8);
  not ginst231 (P1_ADD_405_U99, P1_ADD_405_U10);
  nand ginst232 (P1_ADD_515_U10, P1_INSTADDRPOINTER_REG_4__SCAN_IN, P1_ADD_515_U95);
  not ginst233 (P1_ADD_515_U100, P1_ADD_515_U18);
  not ginst234 (P1_ADD_515_U101, P1_ADD_515_U20);
  not ginst235 (P1_ADD_515_U102, P1_ADD_515_U22);
  not ginst236 (P1_ADD_515_U103, P1_ADD_515_U24);
  not ginst237 (P1_ADD_515_U104, P1_ADD_515_U26);
  not ginst238 (P1_ADD_515_U105, P1_ADD_515_U28);
  not ginst239 (P1_ADD_515_U106, P1_ADD_515_U30);
  not ginst240 (P1_ADD_515_U107, P1_ADD_515_U32);
  not ginst241 (P1_ADD_515_U108, P1_ADD_515_U34);
  not ginst242 (P1_ADD_515_U109, P1_ADD_515_U36);
  not ginst243 (P1_ADD_515_U11, P1_INSTADDRPOINTER_REG_5__SCAN_IN);
  not ginst244 (P1_ADD_515_U110, P1_ADD_515_U38);
  not ginst245 (P1_ADD_515_U111, P1_ADD_515_U40);
  not ginst246 (P1_ADD_515_U112, P1_ADD_515_U42);
  not ginst247 (P1_ADD_515_U113, P1_ADD_515_U44);
  not ginst248 (P1_ADD_515_U114, P1_ADD_515_U46);
  not ginst249 (P1_ADD_515_U115, P1_ADD_515_U48);
  not ginst250 (P1_ADD_515_U116, P1_ADD_515_U50);
  not ginst251 (P1_ADD_515_U117, P1_ADD_515_U52);
  not ginst252 (P1_ADD_515_U118, P1_ADD_515_U54);
  not ginst253 (P1_ADD_515_U119, P1_ADD_515_U56);
  not ginst254 (P1_ADD_515_U12, P1_INSTADDRPOINTER_REG_6__SCAN_IN);
  not ginst255 (P1_ADD_515_U120, P1_ADD_515_U58);
  not ginst256 (P1_ADD_515_U121, P1_ADD_515_U61);
  not ginst257 (P1_ADD_515_U122, P1_ADD_515_U93);
  nand ginst258 (P1_ADD_515_U123, P1_INSTADDRPOINTER_REG_6__SCAN_IN, P1_ADD_515_U13);
  nand ginst259 (P1_ADD_515_U124, P1_ADD_515_U12, P1_ADD_515_U97);
  nand ginst260 (P1_ADD_515_U125, P1_INSTADDRPOINTER_REG_30__SCAN_IN, P1_ADD_515_U61);
  nand ginst261 (P1_ADD_515_U126, P1_ADD_515_U121, P1_ADD_515_U60);
  nand ginst262 (P1_ADD_515_U127, P1_INSTADDRPOINTER_REG_29__SCAN_IN, P1_ADD_515_U58);
  nand ginst263 (P1_ADD_515_U128, P1_ADD_515_U120, P1_ADD_515_U59);
  nand ginst264 (P1_ADD_515_U129, P1_INSTADDRPOINTER_REG_24__SCAN_IN, P1_ADD_515_U48);
  nand ginst265 (P1_ADD_515_U13, P1_INSTADDRPOINTER_REG_5__SCAN_IN, P1_ADD_515_U96);
  nand ginst266 (P1_ADD_515_U130, P1_ADD_515_U115, P1_ADD_515_U49);
  nand ginst267 (P1_ADD_515_U131, P1_INSTADDRPOINTER_REG_17__SCAN_IN, P1_ADD_515_U34);
  nand ginst268 (P1_ADD_515_U132, P1_ADD_515_U108, P1_ADD_515_U35);
  nand ginst269 (P1_ADD_515_U133, P1_INSTADDRPOINTER_REG_2__SCAN_IN, P1_ADD_515_U4);
  nand ginst270 (P1_ADD_515_U134, P1_INSTADDRPOINTER_REG_1__SCAN_IN, P1_ADD_515_U5);
  nand ginst271 (P1_ADD_515_U135, P1_INSTADDRPOINTER_REG_20__SCAN_IN, P1_ADD_515_U40);
  nand ginst272 (P1_ADD_515_U136, P1_ADD_515_U111, P1_ADD_515_U41);
  nand ginst273 (P1_ADD_515_U137, P1_INSTADDRPOINTER_REG_13__SCAN_IN, P1_ADD_515_U26);
  nand ginst274 (P1_ADD_515_U138, P1_ADD_515_U104, P1_ADD_515_U27);
  nand ginst275 (P1_ADD_515_U139, P1_INSTADDRPOINTER_REG_9__SCAN_IN, P1_ADD_515_U18);
  nand ginst276 (P1_ADD_515_U14, P1_INSTADDRPOINTER_REG_6__SCAN_IN, P1_ADD_515_U97);
  nand ginst277 (P1_ADD_515_U140, P1_ADD_515_U100, P1_ADD_515_U19);
  nand ginst278 (P1_ADD_515_U141, P1_INSTADDRPOINTER_REG_22__SCAN_IN, P1_ADD_515_U44);
  nand ginst279 (P1_ADD_515_U142, P1_ADD_515_U113, P1_ADD_515_U45);
  nand ginst280 (P1_ADD_515_U143, P1_INSTADDRPOINTER_REG_18__SCAN_IN, P1_ADD_515_U36);
  nand ginst281 (P1_ADD_515_U144, P1_ADD_515_U109, P1_ADD_515_U37);
  nand ginst282 (P1_ADD_515_U145, P1_INSTADDRPOINTER_REG_11__SCAN_IN, P1_ADD_515_U22);
  nand ginst283 (P1_ADD_515_U146, P1_ADD_515_U102, P1_ADD_515_U23);
  nand ginst284 (P1_ADD_515_U147, P1_INSTADDRPOINTER_REG_26__SCAN_IN, P1_ADD_515_U52);
  nand ginst285 (P1_ADD_515_U148, P1_ADD_515_U117, P1_ADD_515_U53);
  nand ginst286 (P1_ADD_515_U149, P1_INSTADDRPOINTER_REG_15__SCAN_IN, P1_ADD_515_U30);
  not ginst287 (P1_ADD_515_U15, P1_INSTADDRPOINTER_REG_7__SCAN_IN);
  nand ginst288 (P1_ADD_515_U150, P1_ADD_515_U106, P1_ADD_515_U31);
  nand ginst289 (P1_ADD_515_U151, P1_INSTADDRPOINTER_REG_4__SCAN_IN, P1_ADD_515_U8);
  nand ginst290 (P1_ADD_515_U152, P1_ADD_515_U9, P1_ADD_515_U95);
  nand ginst291 (P1_ADD_515_U153, P1_INSTADDRPOINTER_REG_27__SCAN_IN, P1_ADD_515_U54);
  nand ginst292 (P1_ADD_515_U154, P1_ADD_515_U118, P1_ADD_515_U55);
  nand ginst293 (P1_ADD_515_U155, P1_INSTADDRPOINTER_REG_14__SCAN_IN, P1_ADD_515_U28);
  nand ginst294 (P1_ADD_515_U156, P1_ADD_515_U105, P1_ADD_515_U29);
  nand ginst295 (P1_ADD_515_U157, P1_INSTADDRPOINTER_REG_5__SCAN_IN, P1_ADD_515_U10);
  nand ginst296 (P1_ADD_515_U158, P1_ADD_515_U11, P1_ADD_515_U96);
  nand ginst297 (P1_ADD_515_U159, P1_INSTADDRPOINTER_REG_8__SCAN_IN, P1_ADD_515_U16);
  nand ginst298 (P1_ADD_515_U16, P1_INSTADDRPOINTER_REG_7__SCAN_IN, P1_ADD_515_U98);
  nand ginst299 (P1_ADD_515_U160, P1_ADD_515_U17, P1_ADD_515_U99);
  nand ginst300 (P1_ADD_515_U161, P1_INSTADDRPOINTER_REG_23__SCAN_IN, P1_ADD_515_U46);
  nand ginst301 (P1_ADD_515_U162, P1_ADD_515_U114, P1_ADD_515_U47);
  nand ginst302 (P1_ADD_515_U163, P1_INSTADDRPOINTER_REG_19__SCAN_IN, P1_ADD_515_U38);
  nand ginst303 (P1_ADD_515_U164, P1_ADD_515_U110, P1_ADD_515_U39);
  nand ginst304 (P1_ADD_515_U165, P1_INSTADDRPOINTER_REG_10__SCAN_IN, P1_ADD_515_U20);
  nand ginst305 (P1_ADD_515_U166, P1_ADD_515_U101, P1_ADD_515_U21);
  nand ginst306 (P1_ADD_515_U167, P1_INSTADDRPOINTER_REG_31__SCAN_IN, P1_ADD_515_U93);
  nand ginst307 (P1_ADD_515_U168, P1_ADD_515_U122, P1_ADD_515_U92);
  nand ginst308 (P1_ADD_515_U169, P1_INSTADDRPOINTER_REG_3__SCAN_IN, P1_ADD_515_U6);
  not ginst309 (P1_ADD_515_U17, P1_INSTADDRPOINTER_REG_8__SCAN_IN);
  nand ginst310 (P1_ADD_515_U170, P1_ADD_515_U7, P1_ADD_515_U94);
  nand ginst311 (P1_ADD_515_U171, P1_INSTADDRPOINTER_REG_28__SCAN_IN, P1_ADD_515_U56);
  nand ginst312 (P1_ADD_515_U172, P1_ADD_515_U119, P1_ADD_515_U57);
  nand ginst313 (P1_ADD_515_U173, P1_INSTADDRPOINTER_REG_21__SCAN_IN, P1_ADD_515_U42);
  nand ginst314 (P1_ADD_515_U174, P1_ADD_515_U112, P1_ADD_515_U43);
  nand ginst315 (P1_ADD_515_U175, P1_INSTADDRPOINTER_REG_12__SCAN_IN, P1_ADD_515_U24);
  nand ginst316 (P1_ADD_515_U176, P1_ADD_515_U103, P1_ADD_515_U25);
  nand ginst317 (P1_ADD_515_U177, P1_INSTADDRPOINTER_REG_7__SCAN_IN, P1_ADD_515_U14);
  nand ginst318 (P1_ADD_515_U178, P1_ADD_515_U15, P1_ADD_515_U98);
  nand ginst319 (P1_ADD_515_U179, P1_INSTADDRPOINTER_REG_25__SCAN_IN, P1_ADD_515_U50);
  nand ginst320 (P1_ADD_515_U18, P1_INSTADDRPOINTER_REG_8__SCAN_IN, P1_ADD_515_U99);
  nand ginst321 (P1_ADD_515_U180, P1_ADD_515_U116, P1_ADD_515_U51);
  nand ginst322 (P1_ADD_515_U181, P1_INSTADDRPOINTER_REG_16__SCAN_IN, P1_ADD_515_U32);
  nand ginst323 (P1_ADD_515_U182, P1_ADD_515_U107, P1_ADD_515_U33);
  not ginst324 (P1_ADD_515_U19, P1_INSTADDRPOINTER_REG_9__SCAN_IN);
  nand ginst325 (P1_ADD_515_U20, P1_INSTADDRPOINTER_REG_9__SCAN_IN, P1_ADD_515_U100);
  not ginst326 (P1_ADD_515_U21, P1_INSTADDRPOINTER_REG_10__SCAN_IN);
  nand ginst327 (P1_ADD_515_U22, P1_INSTADDRPOINTER_REG_10__SCAN_IN, P1_ADD_515_U101);
  not ginst328 (P1_ADD_515_U23, P1_INSTADDRPOINTER_REG_11__SCAN_IN);
  nand ginst329 (P1_ADD_515_U24, P1_INSTADDRPOINTER_REG_11__SCAN_IN, P1_ADD_515_U102);
  not ginst330 (P1_ADD_515_U25, P1_INSTADDRPOINTER_REG_12__SCAN_IN);
  nand ginst331 (P1_ADD_515_U26, P1_INSTADDRPOINTER_REG_12__SCAN_IN, P1_ADD_515_U103);
  not ginst332 (P1_ADD_515_U27, P1_INSTADDRPOINTER_REG_13__SCAN_IN);
  nand ginst333 (P1_ADD_515_U28, P1_INSTADDRPOINTER_REG_13__SCAN_IN, P1_ADD_515_U104);
  not ginst334 (P1_ADD_515_U29, P1_INSTADDRPOINTER_REG_14__SCAN_IN);
  nand ginst335 (P1_ADD_515_U30, P1_INSTADDRPOINTER_REG_14__SCAN_IN, P1_ADD_515_U105);
  not ginst336 (P1_ADD_515_U31, P1_INSTADDRPOINTER_REG_15__SCAN_IN);
  nand ginst337 (P1_ADD_515_U32, P1_INSTADDRPOINTER_REG_15__SCAN_IN, P1_ADD_515_U106);
  not ginst338 (P1_ADD_515_U33, P1_INSTADDRPOINTER_REG_16__SCAN_IN);
  nand ginst339 (P1_ADD_515_U34, P1_INSTADDRPOINTER_REG_16__SCAN_IN, P1_ADD_515_U107);
  not ginst340 (P1_ADD_515_U35, P1_INSTADDRPOINTER_REG_17__SCAN_IN);
  nand ginst341 (P1_ADD_515_U36, P1_INSTADDRPOINTER_REG_17__SCAN_IN, P1_ADD_515_U108);
  not ginst342 (P1_ADD_515_U37, P1_INSTADDRPOINTER_REG_18__SCAN_IN);
  nand ginst343 (P1_ADD_515_U38, P1_INSTADDRPOINTER_REG_18__SCAN_IN, P1_ADD_515_U109);
  not ginst344 (P1_ADD_515_U39, P1_INSTADDRPOINTER_REG_19__SCAN_IN);
  not ginst345 (P1_ADD_515_U4, P1_INSTADDRPOINTER_REG_1__SCAN_IN);
  nand ginst346 (P1_ADD_515_U40, P1_INSTADDRPOINTER_REG_19__SCAN_IN, P1_ADD_515_U110);
  not ginst347 (P1_ADD_515_U41, P1_INSTADDRPOINTER_REG_20__SCAN_IN);
  nand ginst348 (P1_ADD_515_U42, P1_INSTADDRPOINTER_REG_20__SCAN_IN, P1_ADD_515_U111);
  not ginst349 (P1_ADD_515_U43, P1_INSTADDRPOINTER_REG_21__SCAN_IN);
  nand ginst350 (P1_ADD_515_U44, P1_INSTADDRPOINTER_REG_21__SCAN_IN, P1_ADD_515_U112);
  not ginst351 (P1_ADD_515_U45, P1_INSTADDRPOINTER_REG_22__SCAN_IN);
  nand ginst352 (P1_ADD_515_U46, P1_INSTADDRPOINTER_REG_22__SCAN_IN, P1_ADD_515_U113);
  not ginst353 (P1_ADD_515_U47, P1_INSTADDRPOINTER_REG_23__SCAN_IN);
  nand ginst354 (P1_ADD_515_U48, P1_INSTADDRPOINTER_REG_23__SCAN_IN, P1_ADD_515_U114);
  not ginst355 (P1_ADD_515_U49, P1_INSTADDRPOINTER_REG_24__SCAN_IN);
  not ginst356 (P1_ADD_515_U5, P1_INSTADDRPOINTER_REG_2__SCAN_IN);
  nand ginst357 (P1_ADD_515_U50, P1_INSTADDRPOINTER_REG_24__SCAN_IN, P1_ADD_515_U115);
  not ginst358 (P1_ADD_515_U51, P1_INSTADDRPOINTER_REG_25__SCAN_IN);
  nand ginst359 (P1_ADD_515_U52, P1_INSTADDRPOINTER_REG_25__SCAN_IN, P1_ADD_515_U116);
  not ginst360 (P1_ADD_515_U53, P1_INSTADDRPOINTER_REG_26__SCAN_IN);
  nand ginst361 (P1_ADD_515_U54, P1_INSTADDRPOINTER_REG_26__SCAN_IN, P1_ADD_515_U117);
  not ginst362 (P1_ADD_515_U55, P1_INSTADDRPOINTER_REG_27__SCAN_IN);
  nand ginst363 (P1_ADD_515_U56, P1_INSTADDRPOINTER_REG_27__SCAN_IN, P1_ADD_515_U118);
  not ginst364 (P1_ADD_515_U57, P1_INSTADDRPOINTER_REG_28__SCAN_IN);
  nand ginst365 (P1_ADD_515_U58, P1_INSTADDRPOINTER_REG_28__SCAN_IN, P1_ADD_515_U119);
  not ginst366 (P1_ADD_515_U59, P1_INSTADDRPOINTER_REG_29__SCAN_IN);
  nand ginst367 (P1_ADD_515_U6, P1_INSTADDRPOINTER_REG_2__SCAN_IN, P1_INSTADDRPOINTER_REG_1__SCAN_IN);
  not ginst368 (P1_ADD_515_U60, P1_INSTADDRPOINTER_REG_30__SCAN_IN);
  nand ginst369 (P1_ADD_515_U61, P1_INSTADDRPOINTER_REG_29__SCAN_IN, P1_ADD_515_U120);
  nand ginst370 (P1_ADD_515_U62, P1_ADD_515_U123, P1_ADD_515_U124);
  nand ginst371 (P1_ADD_515_U63, P1_ADD_515_U125, P1_ADD_515_U126);
  nand ginst372 (P1_ADD_515_U64, P1_ADD_515_U127, P1_ADD_515_U128);
  nand ginst373 (P1_ADD_515_U65, P1_ADD_515_U129, P1_ADD_515_U130);
  nand ginst374 (P1_ADD_515_U66, P1_ADD_515_U131, P1_ADD_515_U132);
  nand ginst375 (P1_ADD_515_U67, P1_ADD_515_U133, P1_ADD_515_U134);
  nand ginst376 (P1_ADD_515_U68, P1_ADD_515_U135, P1_ADD_515_U136);
  nand ginst377 (P1_ADD_515_U69, P1_ADD_515_U137, P1_ADD_515_U138);
  not ginst378 (P1_ADD_515_U7, P1_INSTADDRPOINTER_REG_3__SCAN_IN);
  nand ginst379 (P1_ADD_515_U70, P1_ADD_515_U139, P1_ADD_515_U140);
  nand ginst380 (P1_ADD_515_U71, P1_ADD_515_U141, P1_ADD_515_U142);
  nand ginst381 (P1_ADD_515_U72, P1_ADD_515_U143, P1_ADD_515_U144);
  nand ginst382 (P1_ADD_515_U73, P1_ADD_515_U145, P1_ADD_515_U146);
  nand ginst383 (P1_ADD_515_U74, P1_ADD_515_U147, P1_ADD_515_U148);
  nand ginst384 (P1_ADD_515_U75, P1_ADD_515_U149, P1_ADD_515_U150);
  nand ginst385 (P1_ADD_515_U76, P1_ADD_515_U151, P1_ADD_515_U152);
  nand ginst386 (P1_ADD_515_U77, P1_ADD_515_U153, P1_ADD_515_U154);
  nand ginst387 (P1_ADD_515_U78, P1_ADD_515_U155, P1_ADD_515_U156);
  nand ginst388 (P1_ADD_515_U79, P1_ADD_515_U157, P1_ADD_515_U158);
  nand ginst389 (P1_ADD_515_U8, P1_INSTADDRPOINTER_REG_3__SCAN_IN, P1_ADD_515_U94);
  nand ginst390 (P1_ADD_515_U80, P1_ADD_515_U159, P1_ADD_515_U160);
  nand ginst391 (P1_ADD_515_U81, P1_ADD_515_U161, P1_ADD_515_U162);
  nand ginst392 (P1_ADD_515_U82, P1_ADD_515_U163, P1_ADD_515_U164);
  nand ginst393 (P1_ADD_515_U83, P1_ADD_515_U165, P1_ADD_515_U166);
  nand ginst394 (P1_ADD_515_U84, P1_ADD_515_U167, P1_ADD_515_U168);
  nand ginst395 (P1_ADD_515_U85, P1_ADD_515_U169, P1_ADD_515_U170);
  nand ginst396 (P1_ADD_515_U86, P1_ADD_515_U171, P1_ADD_515_U172);
  nand ginst397 (P1_ADD_515_U87, P1_ADD_515_U173, P1_ADD_515_U174);
  nand ginst398 (P1_ADD_515_U88, P1_ADD_515_U175, P1_ADD_515_U176);
  nand ginst399 (P1_ADD_515_U89, P1_ADD_515_U177, P1_ADD_515_U178);
  not ginst400 (P1_ADD_515_U9, P1_INSTADDRPOINTER_REG_4__SCAN_IN);
  nand ginst401 (P1_ADD_515_U90, P1_ADD_515_U179, P1_ADD_515_U180);
  nand ginst402 (P1_ADD_515_U91, P1_ADD_515_U181, P1_ADD_515_U182);
  not ginst403 (P1_ADD_515_U92, P1_INSTADDRPOINTER_REG_31__SCAN_IN);
  nand ginst404 (P1_ADD_515_U93, P1_INSTADDRPOINTER_REG_30__SCAN_IN, P1_ADD_515_U121);
  not ginst405 (P1_ADD_515_U94, P1_ADD_515_U6);
  not ginst406 (P1_ADD_515_U95, P1_ADD_515_U8);
  not ginst407 (P1_ADD_515_U96, P1_ADD_515_U10);
  not ginst408 (P1_ADD_515_U97, P1_ADD_515_U13);
  not ginst409 (P1_ADD_515_U98, P1_ADD_515_U14);
  not ginst410 (P1_ADD_515_U99, P1_ADD_515_U16);
  nor ginst411 (P1_GTE_485_U6, P1_GTE_485_U7, P1_R2238_U6);
  nor ginst412 (P1_GTE_485_U7, P1_R2238_U19, P1_R2238_U20, P1_R2238_U21, P1_R2238_U22);
  and ginst413 (P1_LT_563_1260_U6, P1_LT_563_1260_U8, P1_LT_563_1260_U9);
  not ginst414 (P1_LT_563_1260_U7, P1_U2673);
  nand ginst415 (P1_LT_563_1260_U8, P1_LT_563_1260_U7, P1_R584_U8);
  nand ginst416 (P1_LT_563_1260_U9, P1_LT_563_1260_U7, P1_R584_U9);
  not ginst417 (P1_LT_563_U10, P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN);
  not ginst418 (P1_LT_563_U11, P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN);
  not ginst419 (P1_LT_563_U12, P1_U3489);
  and ginst420 (P1_LT_563_U13, P1_LT_563_U21, P1_LT_563_U22);
  and ginst421 (P1_LT_563_U14, P1_LT_563_U24, P1_LT_563_U25);
  not ginst422 (P1_LT_563_U15, P1_U3492);
  not ginst423 (P1_LT_563_U16, P1_U3493);
  nand ginst424 (P1_LT_563_U17, P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P1_LT_563_U15, P1_LT_563_U16);
  nand ginst425 (P1_LT_563_U18, P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN, P1_LT_563_U15);
  nand ginst426 (P1_LT_563_U19, P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN, P1_LT_563_U8);
  nand ginst427 (P1_LT_563_U20, P1_LT_563_U17, P1_LT_563_U18, P1_LT_563_U19, P1_LT_563_U28);
  nand ginst428 (P1_LT_563_U21, P1_LT_563_U7, P1_U3491);
  nand ginst429 (P1_LT_563_U22, P1_LT_563_U10, P1_U3490);
  nand ginst430 (P1_LT_563_U23, P1_LT_563_U13, P1_LT_563_U20);
  nand ginst431 (P1_LT_563_U24, P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN, P1_LT_563_U9);
  nand ginst432 (P1_LT_563_U25, P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN, P1_LT_563_U12);
  nand ginst433 (P1_LT_563_U26, P1_LT_563_U14, P1_LT_563_U23);
  nand ginst434 (P1_LT_563_U27, P1_LT_563_U11, P1_U3489);
  nand ginst435 (P1_LT_563_U28, P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN, P1_LT_563_U16);
  and ginst436 (P1_LT_563_U6, P1_LT_563_U26, P1_LT_563_U27);
  not ginst437 (P1_LT_563_U7, P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN);
  not ginst438 (P1_LT_563_U8, P1_U3491);
  not ginst439 (P1_LT_563_U9, P1_U3490);
  or ginst440 (P1_LT_589_U6, P1_LT_589_U8, P1_U2673);
  and ginst441 (P1_LT_589_U7, P1_R584_U6, P1_R584_U7);
  nor ginst442 (P1_LT_589_U8, P1_LT_589_U7, P1_R584_U8, P1_R584_U9);
  nand ginst443 (P1_R2027_U10, P1_INSTADDRPOINTER_REG_2__SCAN_IN, P1_INSTADDRPOINTER_REG_1__SCAN_IN, P1_INSTADDRPOINTER_REG_0__SCAN_IN);
  nand ginst444 (P1_R2027_U100, P1_INSTADDRPOINTER_REG_1__SCAN_IN, P1_INSTADDRPOINTER_REG_0__SCAN_IN);
  nand ginst445 (P1_R2027_U101, P1_INSTADDRPOINTER_REG_27__SCAN_IN, P1_R2027_U122);
  nand ginst446 (P1_R2027_U102, P1_INSTADDRPOINTER_REG_25__SCAN_IN, P1_R2027_U116);
  nand ginst447 (P1_R2027_U103, P1_INSTADDRPOINTER_REG_23__SCAN_IN, P1_R2027_U115);
  nand ginst448 (P1_R2027_U104, P1_INSTADDRPOINTER_REG_21__SCAN_IN, P1_R2027_U121);
  nand ginst449 (P1_R2027_U105, P1_INSTADDRPOINTER_REG_19__SCAN_IN, P1_R2027_U114);
  nand ginst450 (P1_R2027_U106, P1_INSTADDRPOINTER_REG_17__SCAN_IN, P1_R2027_U117);
  nand ginst451 (P1_R2027_U107, P1_INSTADDRPOINTER_REG_15__SCAN_IN, P1_R2027_U124);
  nand ginst452 (P1_R2027_U108, P1_INSTADDRPOINTER_REG_13__SCAN_IN, P1_R2027_U119);
  nand ginst453 (P1_R2027_U109, P1_INSTADDRPOINTER_REG_11__SCAN_IN, P1_R2027_U113);
  not ginst454 (P1_R2027_U11, P1_INSTADDRPOINTER_REG_6__SCAN_IN);
  nand ginst455 (P1_R2027_U110, P1_INSTADDRPOINTER_REG_9__SCAN_IN, P1_R2027_U120);
  not ginst456 (P1_R2027_U111, P1_R2027_U10);
  not ginst457 (P1_R2027_U112, P1_R2027_U13);
  not ginst458 (P1_R2027_U113, P1_R2027_U22);
  not ginst459 (P1_R2027_U114, P1_R2027_U34);
  not ginst460 (P1_R2027_U115, P1_R2027_U40);
  not ginst461 (P1_R2027_U116, P1_R2027_U43);
  not ginst462 (P1_R2027_U117, P1_R2027_U31);
  not ginst463 (P1_R2027_U118, P1_R2027_U16);
  not ginst464 (P1_R2027_U119, P1_R2027_U25);
  not ginst465 (P1_R2027_U12, P1_INSTADDRPOINTER_REG_5__SCAN_IN);
  not ginst466 (P1_R2027_U120, P1_R2027_U17);
  not ginst467 (P1_R2027_U121, P1_R2027_U36);
  not ginst468 (P1_R2027_U122, P1_R2027_U46);
  not ginst469 (P1_R2027_U123, P1_R2027_U48);
  not ginst470 (P1_R2027_U124, P1_R2027_U27);
  not ginst471 (P1_R2027_U125, P1_R2027_U95);
  not ginst472 (P1_R2027_U126, P1_R2027_U96);
  not ginst473 (P1_R2027_U127, P1_R2027_U97);
  not ginst474 (P1_R2027_U128, P1_R2027_U49);
  not ginst475 (P1_R2027_U129, P1_R2027_U99);
  nand ginst476 (P1_R2027_U13, P1_R2027_U111, P1_R2027_U82);
  not ginst477 (P1_R2027_U130, P1_R2027_U100);
  not ginst478 (P1_R2027_U131, P1_R2027_U101);
  not ginst479 (P1_R2027_U132, P1_R2027_U102);
  not ginst480 (P1_R2027_U133, P1_R2027_U103);
  not ginst481 (P1_R2027_U134, P1_R2027_U104);
  not ginst482 (P1_R2027_U135, P1_R2027_U105);
  not ginst483 (P1_R2027_U136, P1_R2027_U106);
  not ginst484 (P1_R2027_U137, P1_R2027_U107);
  not ginst485 (P1_R2027_U138, P1_R2027_U108);
  not ginst486 (P1_R2027_U139, P1_R2027_U109);
  not ginst487 (P1_R2027_U14, P1_INSTADDRPOINTER_REG_8__SCAN_IN);
  not ginst488 (P1_R2027_U140, P1_R2027_U110);
  nand ginst489 (P1_R2027_U141, P1_R2027_U120, P1_R2027_U18);
  nand ginst490 (P1_R2027_U142, P1_INSTADDRPOINTER_REG_9__SCAN_IN, P1_R2027_U17);
  nand ginst491 (P1_R2027_U143, P1_INSTADDRPOINTER_REG_8__SCAN_IN, P1_R2027_U95);
  nand ginst492 (P1_R2027_U144, P1_R2027_U125, P1_R2027_U14);
  nand ginst493 (P1_R2027_U145, P1_R2027_U118, P1_R2027_U15);
  nand ginst494 (P1_R2027_U146, P1_INSTADDRPOINTER_REG_7__SCAN_IN, P1_R2027_U16);
  nand ginst495 (P1_R2027_U147, P1_INSTADDRPOINTER_REG_6__SCAN_IN, P1_R2027_U96);
  nand ginst496 (P1_R2027_U148, P1_R2027_U11, P1_R2027_U126);
  nand ginst497 (P1_R2027_U149, P1_R2027_U112, P1_R2027_U12);
  not ginst498 (P1_R2027_U15, P1_INSTADDRPOINTER_REG_7__SCAN_IN);
  nand ginst499 (P1_R2027_U150, P1_INSTADDRPOINTER_REG_5__SCAN_IN, P1_R2027_U13);
  nand ginst500 (P1_R2027_U151, P1_INSTADDRPOINTER_REG_4__SCAN_IN, P1_R2027_U97);
  nand ginst501 (P1_R2027_U152, P1_R2027_U127, P1_R2027_U8);
  nand ginst502 (P1_R2027_U153, P1_R2027_U111, P1_R2027_U9);
  nand ginst503 (P1_R2027_U154, P1_INSTADDRPOINTER_REG_3__SCAN_IN, P1_R2027_U10);
  nand ginst504 (P1_R2027_U155, P1_INSTADDRPOINTER_REG_31__SCAN_IN, P1_R2027_U99);
  nand ginst505 (P1_R2027_U156, P1_R2027_U129, P1_R2027_U98);
  nand ginst506 (P1_R2027_U157, P1_INSTADDRPOINTER_REG_30__SCAN_IN, P1_R2027_U49);
  nand ginst507 (P1_R2027_U158, P1_R2027_U128, P1_R2027_U50);
  nand ginst508 (P1_R2027_U159, P1_INSTADDRPOINTER_REG_2__SCAN_IN, P1_R2027_U100);
  nand ginst509 (P1_R2027_U16, P1_R2027_U112, P1_R2027_U83);
  nand ginst510 (P1_R2027_U160, P1_R2027_U130, P1_R2027_U6);
  nand ginst511 (P1_R2027_U161, P1_R2027_U123, P1_R2027_U47);
  nand ginst512 (P1_R2027_U162, P1_INSTADDRPOINTER_REG_29__SCAN_IN, P1_R2027_U48);
  nand ginst513 (P1_R2027_U163, P1_INSTADDRPOINTER_REG_28__SCAN_IN, P1_R2027_U101);
  nand ginst514 (P1_R2027_U164, P1_R2027_U131, P1_R2027_U45);
  nand ginst515 (P1_R2027_U165, P1_R2027_U122, P1_R2027_U44);
  nand ginst516 (P1_R2027_U166, P1_INSTADDRPOINTER_REG_27__SCAN_IN, P1_R2027_U46);
  nand ginst517 (P1_R2027_U167, P1_INSTADDRPOINTER_REG_26__SCAN_IN, P1_R2027_U102);
  nand ginst518 (P1_R2027_U168, P1_R2027_U132, P1_R2027_U41);
  nand ginst519 (P1_R2027_U169, P1_R2027_U116, P1_R2027_U42);
  nand ginst520 (P1_R2027_U17, P1_R2027_U118, P1_R2027_U84);
  nand ginst521 (P1_R2027_U170, P1_INSTADDRPOINTER_REG_25__SCAN_IN, P1_R2027_U43);
  nand ginst522 (P1_R2027_U171, P1_INSTADDRPOINTER_REG_24__SCAN_IN, P1_R2027_U103);
  nand ginst523 (P1_R2027_U172, P1_R2027_U133, P1_R2027_U38);
  nand ginst524 (P1_R2027_U173, P1_R2027_U115, P1_R2027_U39);
  nand ginst525 (P1_R2027_U174, P1_INSTADDRPOINTER_REG_23__SCAN_IN, P1_R2027_U40);
  nand ginst526 (P1_R2027_U175, P1_INSTADDRPOINTER_REG_22__SCAN_IN, P1_R2027_U104);
  nand ginst527 (P1_R2027_U176, P1_R2027_U134, P1_R2027_U37);
  nand ginst528 (P1_R2027_U177, P1_R2027_U121, P1_R2027_U35);
  nand ginst529 (P1_R2027_U178, P1_INSTADDRPOINTER_REG_21__SCAN_IN, P1_R2027_U36);
  nand ginst530 (P1_R2027_U179, P1_INSTADDRPOINTER_REG_20__SCAN_IN, P1_R2027_U105);
  not ginst531 (P1_R2027_U18, P1_INSTADDRPOINTER_REG_9__SCAN_IN);
  nand ginst532 (P1_R2027_U180, P1_R2027_U135, P1_R2027_U32);
  nand ginst533 (P1_R2027_U181, P1_INSTADDRPOINTER_REG_0__SCAN_IN, P1_R2027_U7);
  nand ginst534 (P1_R2027_U182, P1_INSTADDRPOINTER_REG_1__SCAN_IN, P1_R2027_U5);
  nand ginst535 (P1_R2027_U183, P1_R2027_U114, P1_R2027_U33);
  nand ginst536 (P1_R2027_U184, P1_INSTADDRPOINTER_REG_19__SCAN_IN, P1_R2027_U34);
  nand ginst537 (P1_R2027_U185, P1_INSTADDRPOINTER_REG_18__SCAN_IN, P1_R2027_U106);
  nand ginst538 (P1_R2027_U186, P1_R2027_U136, P1_R2027_U29);
  nand ginst539 (P1_R2027_U187, P1_R2027_U117, P1_R2027_U30);
  nand ginst540 (P1_R2027_U188, P1_INSTADDRPOINTER_REG_17__SCAN_IN, P1_R2027_U31);
  nand ginst541 (P1_R2027_U189, P1_INSTADDRPOINTER_REG_16__SCAN_IN, P1_R2027_U107);
  not ginst542 (P1_R2027_U19, P1_INSTADDRPOINTER_REG_10__SCAN_IN);
  nand ginst543 (P1_R2027_U190, P1_R2027_U137, P1_R2027_U28);
  nand ginst544 (P1_R2027_U191, P1_R2027_U124, P1_R2027_U26);
  nand ginst545 (P1_R2027_U192, P1_INSTADDRPOINTER_REG_15__SCAN_IN, P1_R2027_U27);
  nand ginst546 (P1_R2027_U193, P1_INSTADDRPOINTER_REG_14__SCAN_IN, P1_R2027_U108);
  nand ginst547 (P1_R2027_U194, P1_R2027_U138, P1_R2027_U23);
  nand ginst548 (P1_R2027_U195, P1_R2027_U119, P1_R2027_U24);
  nand ginst549 (P1_R2027_U196, P1_INSTADDRPOINTER_REG_13__SCAN_IN, P1_R2027_U25);
  nand ginst550 (P1_R2027_U197, P1_INSTADDRPOINTER_REG_12__SCAN_IN, P1_R2027_U109);
  nand ginst551 (P1_R2027_U198, P1_R2027_U139, P1_R2027_U20);
  nand ginst552 (P1_R2027_U199, P1_R2027_U113, P1_R2027_U21);
  not ginst553 (P1_R2027_U20, P1_INSTADDRPOINTER_REG_12__SCAN_IN);
  nand ginst554 (P1_R2027_U200, P1_INSTADDRPOINTER_REG_11__SCAN_IN, P1_R2027_U22);
  nand ginst555 (P1_R2027_U201, P1_INSTADDRPOINTER_REG_10__SCAN_IN, P1_R2027_U110);
  nand ginst556 (P1_R2027_U202, P1_R2027_U140, P1_R2027_U19);
  not ginst557 (P1_R2027_U21, P1_INSTADDRPOINTER_REG_11__SCAN_IN);
  nand ginst558 (P1_R2027_U22, P1_R2027_U120, P1_R2027_U85);
  not ginst559 (P1_R2027_U23, P1_INSTADDRPOINTER_REG_14__SCAN_IN);
  not ginst560 (P1_R2027_U24, P1_INSTADDRPOINTER_REG_13__SCAN_IN);
  nand ginst561 (P1_R2027_U25, P1_R2027_U113, P1_R2027_U86);
  not ginst562 (P1_R2027_U26, P1_INSTADDRPOINTER_REG_15__SCAN_IN);
  nand ginst563 (P1_R2027_U27, P1_R2027_U119, P1_R2027_U87);
  not ginst564 (P1_R2027_U28, P1_INSTADDRPOINTER_REG_16__SCAN_IN);
  not ginst565 (P1_R2027_U29, P1_INSTADDRPOINTER_REG_18__SCAN_IN);
  not ginst566 (P1_R2027_U30, P1_INSTADDRPOINTER_REG_17__SCAN_IN);
  nand ginst567 (P1_R2027_U31, P1_R2027_U124, P1_R2027_U88);
  not ginst568 (P1_R2027_U32, P1_INSTADDRPOINTER_REG_20__SCAN_IN);
  not ginst569 (P1_R2027_U33, P1_INSTADDRPOINTER_REG_19__SCAN_IN);
  nand ginst570 (P1_R2027_U34, P1_R2027_U117, P1_R2027_U89);
  not ginst571 (P1_R2027_U35, P1_INSTADDRPOINTER_REG_21__SCAN_IN);
  nand ginst572 (P1_R2027_U36, P1_R2027_U114, P1_R2027_U90);
  not ginst573 (P1_R2027_U37, P1_INSTADDRPOINTER_REG_22__SCAN_IN);
  not ginst574 (P1_R2027_U38, P1_INSTADDRPOINTER_REG_24__SCAN_IN);
  not ginst575 (P1_R2027_U39, P1_INSTADDRPOINTER_REG_23__SCAN_IN);
  nand ginst576 (P1_R2027_U40, P1_R2027_U121, P1_R2027_U91);
  not ginst577 (P1_R2027_U41, P1_INSTADDRPOINTER_REG_26__SCAN_IN);
  not ginst578 (P1_R2027_U42, P1_INSTADDRPOINTER_REG_25__SCAN_IN);
  nand ginst579 (P1_R2027_U43, P1_R2027_U115, P1_R2027_U92);
  not ginst580 (P1_R2027_U44, P1_INSTADDRPOINTER_REG_27__SCAN_IN);
  not ginst581 (P1_R2027_U45, P1_INSTADDRPOINTER_REG_28__SCAN_IN);
  nand ginst582 (P1_R2027_U46, P1_R2027_U116, P1_R2027_U93);
  not ginst583 (P1_R2027_U47, P1_INSTADDRPOINTER_REG_29__SCAN_IN);
  nand ginst584 (P1_R2027_U48, P1_R2027_U122, P1_R2027_U94);
  nand ginst585 (P1_R2027_U49, P1_INSTADDRPOINTER_REG_29__SCAN_IN, P1_R2027_U123);
  not ginst586 (P1_R2027_U5, P1_INSTADDRPOINTER_REG_0__SCAN_IN);
  not ginst587 (P1_R2027_U50, P1_INSTADDRPOINTER_REG_30__SCAN_IN);
  nand ginst588 (P1_R2027_U51, P1_R2027_U141, P1_R2027_U142);
  nand ginst589 (P1_R2027_U52, P1_R2027_U143, P1_R2027_U144);
  nand ginst590 (P1_R2027_U53, P1_R2027_U145, P1_R2027_U146);
  nand ginst591 (P1_R2027_U54, P1_R2027_U147, P1_R2027_U148);
  nand ginst592 (P1_R2027_U55, P1_R2027_U149, P1_R2027_U150);
  nand ginst593 (P1_R2027_U56, P1_R2027_U151, P1_R2027_U152);
  nand ginst594 (P1_R2027_U57, P1_R2027_U153, P1_R2027_U154);
  nand ginst595 (P1_R2027_U58, P1_R2027_U155, P1_R2027_U156);
  nand ginst596 (P1_R2027_U59, P1_R2027_U157, P1_R2027_U158);
  not ginst597 (P1_R2027_U6, P1_INSTADDRPOINTER_REG_2__SCAN_IN);
  nand ginst598 (P1_R2027_U60, P1_R2027_U159, P1_R2027_U160);
  nand ginst599 (P1_R2027_U61, P1_R2027_U161, P1_R2027_U162);
  nand ginst600 (P1_R2027_U62, P1_R2027_U163, P1_R2027_U164);
  nand ginst601 (P1_R2027_U63, P1_R2027_U165, P1_R2027_U166);
  nand ginst602 (P1_R2027_U64, P1_R2027_U167, P1_R2027_U168);
  nand ginst603 (P1_R2027_U65, P1_R2027_U169, P1_R2027_U170);
  nand ginst604 (P1_R2027_U66, P1_R2027_U171, P1_R2027_U172);
  nand ginst605 (P1_R2027_U67, P1_R2027_U173, P1_R2027_U174);
  nand ginst606 (P1_R2027_U68, P1_R2027_U175, P1_R2027_U176);
  nand ginst607 (P1_R2027_U69, P1_R2027_U177, P1_R2027_U178);
  not ginst608 (P1_R2027_U7, P1_INSTADDRPOINTER_REG_1__SCAN_IN);
  nand ginst609 (P1_R2027_U70, P1_R2027_U179, P1_R2027_U180);
  nand ginst610 (P1_R2027_U71, P1_R2027_U181, P1_R2027_U182);
  nand ginst611 (P1_R2027_U72, P1_R2027_U183, P1_R2027_U184);
  nand ginst612 (P1_R2027_U73, P1_R2027_U185, P1_R2027_U186);
  nand ginst613 (P1_R2027_U74, P1_R2027_U187, P1_R2027_U188);
  nand ginst614 (P1_R2027_U75, P1_R2027_U189, P1_R2027_U190);
  nand ginst615 (P1_R2027_U76, P1_R2027_U191, P1_R2027_U192);
  nand ginst616 (P1_R2027_U77, P1_R2027_U193, P1_R2027_U194);
  nand ginst617 (P1_R2027_U78, P1_R2027_U195, P1_R2027_U196);
  nand ginst618 (P1_R2027_U79, P1_R2027_U197, P1_R2027_U198);
  not ginst619 (P1_R2027_U8, P1_INSTADDRPOINTER_REG_4__SCAN_IN);
  nand ginst620 (P1_R2027_U80, P1_R2027_U199, P1_R2027_U200);
  nand ginst621 (P1_R2027_U81, P1_R2027_U201, P1_R2027_U202);
  and ginst622 (P1_R2027_U82, P1_INSTADDRPOINTER_REG_4__SCAN_IN, P1_INSTADDRPOINTER_REG_3__SCAN_IN);
  and ginst623 (P1_R2027_U83, P1_INSTADDRPOINTER_REG_6__SCAN_IN, P1_INSTADDRPOINTER_REG_5__SCAN_IN);
  and ginst624 (P1_R2027_U84, P1_INSTADDRPOINTER_REG_8__SCAN_IN, P1_INSTADDRPOINTER_REG_7__SCAN_IN);
  and ginst625 (P1_R2027_U85, P1_INSTADDRPOINTER_REG_10__SCAN_IN, P1_INSTADDRPOINTER_REG_9__SCAN_IN);
  and ginst626 (P1_R2027_U86, P1_INSTADDRPOINTER_REG_12__SCAN_IN, P1_INSTADDRPOINTER_REG_11__SCAN_IN);
  and ginst627 (P1_R2027_U87, P1_INSTADDRPOINTER_REG_14__SCAN_IN, P1_INSTADDRPOINTER_REG_13__SCAN_IN);
  and ginst628 (P1_R2027_U88, P1_INSTADDRPOINTER_REG_16__SCAN_IN, P1_INSTADDRPOINTER_REG_15__SCAN_IN);
  and ginst629 (P1_R2027_U89, P1_INSTADDRPOINTER_REG_18__SCAN_IN, P1_INSTADDRPOINTER_REG_17__SCAN_IN);
  not ginst630 (P1_R2027_U9, P1_INSTADDRPOINTER_REG_3__SCAN_IN);
  and ginst631 (P1_R2027_U90, P1_INSTADDRPOINTER_REG_20__SCAN_IN, P1_INSTADDRPOINTER_REG_19__SCAN_IN);
  and ginst632 (P1_R2027_U91, P1_INSTADDRPOINTER_REG_22__SCAN_IN, P1_INSTADDRPOINTER_REG_21__SCAN_IN);
  and ginst633 (P1_R2027_U92, P1_INSTADDRPOINTER_REG_24__SCAN_IN, P1_INSTADDRPOINTER_REG_23__SCAN_IN);
  and ginst634 (P1_R2027_U93, P1_INSTADDRPOINTER_REG_26__SCAN_IN, P1_INSTADDRPOINTER_REG_25__SCAN_IN);
  and ginst635 (P1_R2027_U94, P1_INSTADDRPOINTER_REG_28__SCAN_IN, P1_INSTADDRPOINTER_REG_27__SCAN_IN);
  nand ginst636 (P1_R2027_U95, P1_INSTADDRPOINTER_REG_7__SCAN_IN, P1_R2027_U118);
  nand ginst637 (P1_R2027_U96, P1_INSTADDRPOINTER_REG_5__SCAN_IN, P1_R2027_U112);
  nand ginst638 (P1_R2027_U97, P1_INSTADDRPOINTER_REG_3__SCAN_IN, P1_R2027_U111);
  not ginst639 (P1_R2027_U98, P1_INSTADDRPOINTER_REG_31__SCAN_IN);
  nand ginst640 (P1_R2027_U99, P1_INSTADDRPOINTER_REG_30__SCAN_IN, P1_R2027_U128);
  nand ginst641 (P1_R2096_U10, P1_REIP_REG_4__SCAN_IN, P1_R2096_U95);
  not ginst642 (P1_R2096_U100, P1_R2096_U19);
  not ginst643 (P1_R2096_U101, P1_R2096_U20);
  not ginst644 (P1_R2096_U102, P1_R2096_U22);
  not ginst645 (P1_R2096_U103, P1_R2096_U24);
  not ginst646 (P1_R2096_U104, P1_R2096_U26);
  not ginst647 (P1_R2096_U105, P1_R2096_U28);
  not ginst648 (P1_R2096_U106, P1_R2096_U30);
  not ginst649 (P1_R2096_U107, P1_R2096_U32);
  not ginst650 (P1_R2096_U108, P1_R2096_U34);
  not ginst651 (P1_R2096_U109, P1_R2096_U36);
  not ginst652 (P1_R2096_U11, P1_REIP_REG_5__SCAN_IN);
  not ginst653 (P1_R2096_U110, P1_R2096_U38);
  not ginst654 (P1_R2096_U111, P1_R2096_U40);
  not ginst655 (P1_R2096_U112, P1_R2096_U42);
  not ginst656 (P1_R2096_U113, P1_R2096_U44);
  not ginst657 (P1_R2096_U114, P1_R2096_U46);
  not ginst658 (P1_R2096_U115, P1_R2096_U48);
  not ginst659 (P1_R2096_U116, P1_R2096_U50);
  not ginst660 (P1_R2096_U117, P1_R2096_U52);
  not ginst661 (P1_R2096_U118, P1_R2096_U54);
  not ginst662 (P1_R2096_U119, P1_R2096_U56);
  nand ginst663 (P1_R2096_U12, P1_REIP_REG_5__SCAN_IN, P1_R2096_U96);
  not ginst664 (P1_R2096_U120, P1_R2096_U58);
  not ginst665 (P1_R2096_U121, P1_R2096_U60);
  not ginst666 (P1_R2096_U122, P1_R2096_U93);
  nand ginst667 (P1_R2096_U123, P1_REIP_REG_9__SCAN_IN, P1_R2096_U19);
  nand ginst668 (P1_R2096_U124, P1_R2096_U100, P1_R2096_U18);
  nand ginst669 (P1_R2096_U125, P1_REIP_REG_8__SCAN_IN, P1_R2096_U16);
  nand ginst670 (P1_R2096_U126, P1_R2096_U17, P1_R2096_U99);
  nand ginst671 (P1_R2096_U127, P1_REIP_REG_7__SCAN_IN, P1_R2096_U14);
  nand ginst672 (P1_R2096_U128, P1_R2096_U15, P1_R2096_U98);
  nand ginst673 (P1_R2096_U129, P1_REIP_REG_6__SCAN_IN, P1_R2096_U12);
  not ginst674 (P1_R2096_U13, P1_REIP_REG_6__SCAN_IN);
  nand ginst675 (P1_R2096_U130, P1_R2096_U13, P1_R2096_U97);
  nand ginst676 (P1_R2096_U131, P1_REIP_REG_5__SCAN_IN, P1_R2096_U10);
  nand ginst677 (P1_R2096_U132, P1_R2096_U11, P1_R2096_U96);
  nand ginst678 (P1_R2096_U133, P1_REIP_REG_4__SCAN_IN, P1_R2096_U8);
  nand ginst679 (P1_R2096_U134, P1_R2096_U9, P1_R2096_U95);
  nand ginst680 (P1_R2096_U135, P1_REIP_REG_3__SCAN_IN, P1_R2096_U6);
  nand ginst681 (P1_R2096_U136, P1_R2096_U7, P1_R2096_U94);
  nand ginst682 (P1_R2096_U137, P1_REIP_REG_31__SCAN_IN, P1_R2096_U93);
  nand ginst683 (P1_R2096_U138, P1_R2096_U122, P1_R2096_U92);
  nand ginst684 (P1_R2096_U139, P1_REIP_REG_30__SCAN_IN, P1_R2096_U60);
  nand ginst685 (P1_R2096_U14, P1_REIP_REG_6__SCAN_IN, P1_R2096_U97);
  nand ginst686 (P1_R2096_U140, P1_R2096_U121, P1_R2096_U61);
  nand ginst687 (P1_R2096_U141, P1_REIP_REG_2__SCAN_IN, P1_R2096_U4);
  nand ginst688 (P1_R2096_U142, P1_REIP_REG_1__SCAN_IN, P1_R2096_U5);
  nand ginst689 (P1_R2096_U143, P1_REIP_REG_29__SCAN_IN, P1_R2096_U58);
  nand ginst690 (P1_R2096_U144, P1_R2096_U120, P1_R2096_U59);
  nand ginst691 (P1_R2096_U145, P1_REIP_REG_28__SCAN_IN, P1_R2096_U56);
  nand ginst692 (P1_R2096_U146, P1_R2096_U119, P1_R2096_U57);
  nand ginst693 (P1_R2096_U147, P1_REIP_REG_27__SCAN_IN, P1_R2096_U54);
  nand ginst694 (P1_R2096_U148, P1_R2096_U118, P1_R2096_U55);
  nand ginst695 (P1_R2096_U149, P1_REIP_REG_26__SCAN_IN, P1_R2096_U52);
  not ginst696 (P1_R2096_U15, P1_REIP_REG_7__SCAN_IN);
  nand ginst697 (P1_R2096_U150, P1_R2096_U117, P1_R2096_U53);
  nand ginst698 (P1_R2096_U151, P1_REIP_REG_25__SCAN_IN, P1_R2096_U50);
  nand ginst699 (P1_R2096_U152, P1_R2096_U116, P1_R2096_U51);
  nand ginst700 (P1_R2096_U153, P1_REIP_REG_24__SCAN_IN, P1_R2096_U48);
  nand ginst701 (P1_R2096_U154, P1_R2096_U115, P1_R2096_U49);
  nand ginst702 (P1_R2096_U155, P1_REIP_REG_23__SCAN_IN, P1_R2096_U46);
  nand ginst703 (P1_R2096_U156, P1_R2096_U114, P1_R2096_U47);
  nand ginst704 (P1_R2096_U157, P1_REIP_REG_22__SCAN_IN, P1_R2096_U44);
  nand ginst705 (P1_R2096_U158, P1_R2096_U113, P1_R2096_U45);
  nand ginst706 (P1_R2096_U159, P1_REIP_REG_21__SCAN_IN, P1_R2096_U42);
  nand ginst707 (P1_R2096_U16, P1_REIP_REG_7__SCAN_IN, P1_R2096_U98);
  nand ginst708 (P1_R2096_U160, P1_R2096_U112, P1_R2096_U43);
  nand ginst709 (P1_R2096_U161, P1_REIP_REG_20__SCAN_IN, P1_R2096_U40);
  nand ginst710 (P1_R2096_U162, P1_R2096_U111, P1_R2096_U41);
  nand ginst711 (P1_R2096_U163, P1_REIP_REG_19__SCAN_IN, P1_R2096_U38);
  nand ginst712 (P1_R2096_U164, P1_R2096_U110, P1_R2096_U39);
  nand ginst713 (P1_R2096_U165, P1_REIP_REG_18__SCAN_IN, P1_R2096_U36);
  nand ginst714 (P1_R2096_U166, P1_R2096_U109, P1_R2096_U37);
  nand ginst715 (P1_R2096_U167, P1_REIP_REG_17__SCAN_IN, P1_R2096_U34);
  nand ginst716 (P1_R2096_U168, P1_R2096_U108, P1_R2096_U35);
  nand ginst717 (P1_R2096_U169, P1_REIP_REG_16__SCAN_IN, P1_R2096_U32);
  not ginst718 (P1_R2096_U17, P1_REIP_REG_8__SCAN_IN);
  nand ginst719 (P1_R2096_U170, P1_R2096_U107, P1_R2096_U33);
  nand ginst720 (P1_R2096_U171, P1_REIP_REG_15__SCAN_IN, P1_R2096_U30);
  nand ginst721 (P1_R2096_U172, P1_R2096_U106, P1_R2096_U31);
  nand ginst722 (P1_R2096_U173, P1_REIP_REG_14__SCAN_IN, P1_R2096_U28);
  nand ginst723 (P1_R2096_U174, P1_R2096_U105, P1_R2096_U29);
  nand ginst724 (P1_R2096_U175, P1_REIP_REG_13__SCAN_IN, P1_R2096_U26);
  nand ginst725 (P1_R2096_U176, P1_R2096_U104, P1_R2096_U27);
  nand ginst726 (P1_R2096_U177, P1_REIP_REG_12__SCAN_IN, P1_R2096_U24);
  nand ginst727 (P1_R2096_U178, P1_R2096_U103, P1_R2096_U25);
  nand ginst728 (P1_R2096_U179, P1_REIP_REG_11__SCAN_IN, P1_R2096_U22);
  not ginst729 (P1_R2096_U18, P1_REIP_REG_9__SCAN_IN);
  nand ginst730 (P1_R2096_U180, P1_R2096_U102, P1_R2096_U23);
  nand ginst731 (P1_R2096_U181, P1_REIP_REG_10__SCAN_IN, P1_R2096_U20);
  nand ginst732 (P1_R2096_U182, P1_R2096_U101, P1_R2096_U21);
  nand ginst733 (P1_R2096_U19, P1_REIP_REG_8__SCAN_IN, P1_R2096_U99);
  nand ginst734 (P1_R2096_U20, P1_REIP_REG_9__SCAN_IN, P1_R2096_U100);
  not ginst735 (P1_R2096_U21, P1_REIP_REG_10__SCAN_IN);
  nand ginst736 (P1_R2096_U22, P1_REIP_REG_10__SCAN_IN, P1_R2096_U101);
  not ginst737 (P1_R2096_U23, P1_REIP_REG_11__SCAN_IN);
  nand ginst738 (P1_R2096_U24, P1_REIP_REG_11__SCAN_IN, P1_R2096_U102);
  not ginst739 (P1_R2096_U25, P1_REIP_REG_12__SCAN_IN);
  nand ginst740 (P1_R2096_U26, P1_REIP_REG_12__SCAN_IN, P1_R2096_U103);
  not ginst741 (P1_R2096_U27, P1_REIP_REG_13__SCAN_IN);
  nand ginst742 (P1_R2096_U28, P1_REIP_REG_13__SCAN_IN, P1_R2096_U104);
  not ginst743 (P1_R2096_U29, P1_REIP_REG_14__SCAN_IN);
  nand ginst744 (P1_R2096_U30, P1_REIP_REG_14__SCAN_IN, P1_R2096_U105);
  not ginst745 (P1_R2096_U31, P1_REIP_REG_15__SCAN_IN);
  nand ginst746 (P1_R2096_U32, P1_REIP_REG_15__SCAN_IN, P1_R2096_U106);
  not ginst747 (P1_R2096_U33, P1_REIP_REG_16__SCAN_IN);
  nand ginst748 (P1_R2096_U34, P1_REIP_REG_16__SCAN_IN, P1_R2096_U107);
  not ginst749 (P1_R2096_U35, P1_REIP_REG_17__SCAN_IN);
  nand ginst750 (P1_R2096_U36, P1_REIP_REG_17__SCAN_IN, P1_R2096_U108);
  not ginst751 (P1_R2096_U37, P1_REIP_REG_18__SCAN_IN);
  nand ginst752 (P1_R2096_U38, P1_REIP_REG_18__SCAN_IN, P1_R2096_U109);
  not ginst753 (P1_R2096_U39, P1_REIP_REG_19__SCAN_IN);
  not ginst754 (P1_R2096_U4, P1_REIP_REG_1__SCAN_IN);
  nand ginst755 (P1_R2096_U40, P1_REIP_REG_19__SCAN_IN, P1_R2096_U110);
  not ginst756 (P1_R2096_U41, P1_REIP_REG_20__SCAN_IN);
  nand ginst757 (P1_R2096_U42, P1_REIP_REG_20__SCAN_IN, P1_R2096_U111);
  not ginst758 (P1_R2096_U43, P1_REIP_REG_21__SCAN_IN);
  nand ginst759 (P1_R2096_U44, P1_REIP_REG_21__SCAN_IN, P1_R2096_U112);
  not ginst760 (P1_R2096_U45, P1_REIP_REG_22__SCAN_IN);
  nand ginst761 (P1_R2096_U46, P1_REIP_REG_22__SCAN_IN, P1_R2096_U113);
  not ginst762 (P1_R2096_U47, P1_REIP_REG_23__SCAN_IN);
  nand ginst763 (P1_R2096_U48, P1_REIP_REG_23__SCAN_IN, P1_R2096_U114);
  not ginst764 (P1_R2096_U49, P1_REIP_REG_24__SCAN_IN);
  not ginst765 (P1_R2096_U5, P1_REIP_REG_2__SCAN_IN);
  nand ginst766 (P1_R2096_U50, P1_REIP_REG_24__SCAN_IN, P1_R2096_U115);
  not ginst767 (P1_R2096_U51, P1_REIP_REG_25__SCAN_IN);
  nand ginst768 (P1_R2096_U52, P1_REIP_REG_25__SCAN_IN, P1_R2096_U116);
  not ginst769 (P1_R2096_U53, P1_REIP_REG_26__SCAN_IN);
  nand ginst770 (P1_R2096_U54, P1_REIP_REG_26__SCAN_IN, P1_R2096_U117);
  not ginst771 (P1_R2096_U55, P1_REIP_REG_27__SCAN_IN);
  nand ginst772 (P1_R2096_U56, P1_REIP_REG_27__SCAN_IN, P1_R2096_U118);
  not ginst773 (P1_R2096_U57, P1_REIP_REG_28__SCAN_IN);
  nand ginst774 (P1_R2096_U58, P1_REIP_REG_28__SCAN_IN, P1_R2096_U119);
  not ginst775 (P1_R2096_U59, P1_REIP_REG_29__SCAN_IN);
  nand ginst776 (P1_R2096_U6, P1_REIP_REG_2__SCAN_IN, P1_REIP_REG_1__SCAN_IN);
  nand ginst777 (P1_R2096_U60, P1_REIP_REG_29__SCAN_IN, P1_R2096_U120);
  not ginst778 (P1_R2096_U61, P1_REIP_REG_30__SCAN_IN);
  nand ginst779 (P1_R2096_U62, P1_R2096_U123, P1_R2096_U124);
  nand ginst780 (P1_R2096_U63, P1_R2096_U125, P1_R2096_U126);
  nand ginst781 (P1_R2096_U64, P1_R2096_U127, P1_R2096_U128);
  nand ginst782 (P1_R2096_U65, P1_R2096_U129, P1_R2096_U130);
  nand ginst783 (P1_R2096_U66, P1_R2096_U131, P1_R2096_U132);
  nand ginst784 (P1_R2096_U67, P1_R2096_U133, P1_R2096_U134);
  nand ginst785 (P1_R2096_U68, P1_R2096_U135, P1_R2096_U136);
  nand ginst786 (P1_R2096_U69, P1_R2096_U137, P1_R2096_U138);
  not ginst787 (P1_R2096_U7, P1_REIP_REG_3__SCAN_IN);
  nand ginst788 (P1_R2096_U70, P1_R2096_U139, P1_R2096_U140);
  nand ginst789 (P1_R2096_U71, P1_R2096_U141, P1_R2096_U142);
  nand ginst790 (P1_R2096_U72, P1_R2096_U143, P1_R2096_U144);
  nand ginst791 (P1_R2096_U73, P1_R2096_U145, P1_R2096_U146);
  nand ginst792 (P1_R2096_U74, P1_R2096_U147, P1_R2096_U148);
  nand ginst793 (P1_R2096_U75, P1_R2096_U149, P1_R2096_U150);
  nand ginst794 (P1_R2096_U76, P1_R2096_U151, P1_R2096_U152);
  nand ginst795 (P1_R2096_U77, P1_R2096_U153, P1_R2096_U154);
  nand ginst796 (P1_R2096_U78, P1_R2096_U155, P1_R2096_U156);
  nand ginst797 (P1_R2096_U79, P1_R2096_U157, P1_R2096_U158);
  nand ginst798 (P1_R2096_U8, P1_REIP_REG_3__SCAN_IN, P1_R2096_U94);
  nand ginst799 (P1_R2096_U80, P1_R2096_U159, P1_R2096_U160);
  nand ginst800 (P1_R2096_U81, P1_R2096_U161, P1_R2096_U162);
  nand ginst801 (P1_R2096_U82, P1_R2096_U163, P1_R2096_U164);
  nand ginst802 (P1_R2096_U83, P1_R2096_U165, P1_R2096_U166);
  nand ginst803 (P1_R2096_U84, P1_R2096_U167, P1_R2096_U168);
  nand ginst804 (P1_R2096_U85, P1_R2096_U169, P1_R2096_U170);
  nand ginst805 (P1_R2096_U86, P1_R2096_U171, P1_R2096_U172);
  nand ginst806 (P1_R2096_U87, P1_R2096_U173, P1_R2096_U174);
  nand ginst807 (P1_R2096_U88, P1_R2096_U175, P1_R2096_U176);
  nand ginst808 (P1_R2096_U89, P1_R2096_U177, P1_R2096_U178);
  not ginst809 (P1_R2096_U9, P1_REIP_REG_4__SCAN_IN);
  nand ginst810 (P1_R2096_U90, P1_R2096_U179, P1_R2096_U180);
  nand ginst811 (P1_R2096_U91, P1_R2096_U181, P1_R2096_U182);
  not ginst812 (P1_R2096_U92, P1_REIP_REG_31__SCAN_IN);
  nand ginst813 (P1_R2096_U93, P1_REIP_REG_30__SCAN_IN, P1_R2096_U121);
  not ginst814 (P1_R2096_U94, P1_R2096_U6);
  not ginst815 (P1_R2096_U95, P1_R2096_U8);
  not ginst816 (P1_R2096_U96, P1_R2096_U10);
  not ginst817 (P1_R2096_U97, P1_R2096_U12);
  not ginst818 (P1_R2096_U98, P1_R2096_U14);
  not ginst819 (P1_R2096_U99, P1_R2096_U16);
  nand ginst820 (P1_R2099_U10, P1_R2099_U159, P1_R2099_U91);
  not ginst821 (P1_R2099_U100, P1_U2710);
  not ginst822 (P1_R2099_U101, P1_U2709);
  not ginst823 (P1_R2099_U102, P1_U2708);
  not ginst824 (P1_R2099_U103, P1_U2707);
  not ginst825 (P1_R2099_U104, P1_U2706);
  not ginst826 (P1_R2099_U105, P1_U2705);
  not ginst827 (P1_R2099_U106, P1_U2704);
  not ginst828 (P1_R2099_U107, P1_U2703);
  not ginst829 (P1_R2099_U108, P1_U2701);
  nand ginst830 (P1_R2099_U109, P1_R2099_U159, P1_R2099_U27);
  nand ginst831 (P1_R2099_U11, P1_R2099_U161, P1_R2099_U92);
  nand ginst832 (P1_R2099_U110, P1_R2099_U157, P1_R2099_U28);
  nand ginst833 (P1_R2099_U111, P1_R2099_U155, P1_R2099_U30);
  nand ginst834 (P1_R2099_U112, P1_R2099_U137, P1_R2099_U35);
  not ginst835 (P1_R2099_U113, P1_U2682);
  not ginst836 (P1_R2099_U114, P1_U2683);
  not ginst837 (P1_R2099_U115, P1_U2684);
  not ginst838 (P1_R2099_U116, P1_U2685);
  not ginst839 (P1_R2099_U117, P1_U2686);
  not ginst840 (P1_R2099_U118, P1_U2687);
  not ginst841 (P1_R2099_U119, P1_U2688);
  nand ginst842 (P1_R2099_U12, P1_R2099_U163, P1_R2099_U93);
  not ginst843 (P1_R2099_U120, P1_U2689);
  not ginst844 (P1_R2099_U121, P1_U2690);
  not ginst845 (P1_R2099_U122, P1_U2691);
  not ginst846 (P1_R2099_U123, P1_U2692);
  not ginst847 (P1_R2099_U124, P1_U2700);
  not ginst848 (P1_R2099_U125, P1_U2699);
  not ginst849 (P1_R2099_U126, P1_U2698);
  not ginst850 (P1_R2099_U127, P1_U2697);
  not ginst851 (P1_R2099_U128, P1_U2696);
  not ginst852 (P1_R2099_U129, P1_U2695);
  nand ginst853 (P1_R2099_U13, P1_R2099_U165, P1_R2099_U94);
  not ginst854 (P1_R2099_U130, P1_U2694);
  not ginst855 (P1_R2099_U131, P1_U2693);
  not ginst856 (P1_R2099_U132, P1_U2680);
  not ginst857 (P1_R2099_U133, P1_U2681);
  not ginst858 (P1_R2099_U134, P1_U2679);
  nand ginst859 (P1_R2099_U135, P1_R2099_U180, P1_R2099_U96);
  nand ginst860 (P1_R2099_U136, P1_R2099_U180, P1_R2099_U44);
  nand ginst861 (P1_R2099_U137, P1_R2099_U151, P1_R2099_U152);
  and ginst862 (P1_R2099_U138, P1_R2099_U296, P1_R2099_U297);
  and ginst863 (P1_R2099_U139, P1_R2099_U318, P1_R2099_U319);
  nand ginst864 (P1_R2099_U14, P1_R2099_U167, P1_R2099_U95);
  nand ginst865 (P1_R2099_U140, P1_R2099_U147, P1_R2099_U148);
  nand ginst866 (P1_R2099_U141, P1_R2099_U167, P1_R2099_U56);
  nand ginst867 (P1_R2099_U142, P1_R2099_U165, P1_R2099_U58);
  nand ginst868 (P1_R2099_U143, P1_R2099_U163, P1_R2099_U60);
  nand ginst869 (P1_R2099_U144, P1_R2099_U161, P1_R2099_U62);
  not ginst870 (P1_R2099_U145, P1_R2099_U135);
  or ginst871 (P1_R2099_U146, P1_U4189, P1_U4190);
  nand ginst872 (P1_R2099_U147, P1_R2099_U146, P1_R2099_U32);
  nand ginst873 (P1_R2099_U148, P1_U4189, P1_U4190);
  not ginst874 (P1_R2099_U149, P1_R2099_U140);
  nand ginst875 (P1_R2099_U15, P1_R2099_U169, P1_R2099_U55);
  nand ginst876 (P1_R2099_U150, P1_R2099_U190, P1_R2099_U6);
  nand ginst877 (P1_R2099_U151, P1_R2099_U140, P1_R2099_U150);
  nand ginst878 (P1_R2099_U152, P1_R2099_U33, P1_U2678);
  not ginst879 (P1_R2099_U153, P1_R2099_U137);
  not ginst880 (P1_R2099_U154, P1_R2099_U112);
  not ginst881 (P1_R2099_U155, P1_R2099_U7);
  not ginst882 (P1_R2099_U156, P1_R2099_U111);
  not ginst883 (P1_R2099_U157, P1_R2099_U8);
  not ginst884 (P1_R2099_U158, P1_R2099_U110);
  not ginst885 (P1_R2099_U159, P1_R2099_U9);
  nand ginst886 (P1_R2099_U16, P1_R2099_U170, P1_R2099_U54);
  not ginst887 (P1_R2099_U160, P1_R2099_U109);
  not ginst888 (P1_R2099_U161, P1_R2099_U10);
  not ginst889 (P1_R2099_U162, P1_R2099_U144);
  not ginst890 (P1_R2099_U163, P1_R2099_U11);
  not ginst891 (P1_R2099_U164, P1_R2099_U143);
  not ginst892 (P1_R2099_U165, P1_R2099_U12);
  not ginst893 (P1_R2099_U166, P1_R2099_U142);
  not ginst894 (P1_R2099_U167, P1_R2099_U13);
  not ginst895 (P1_R2099_U168, P1_R2099_U141);
  not ginst896 (P1_R2099_U169, P1_R2099_U14);
  nand ginst897 (P1_R2099_U17, P1_R2099_U171, P1_R2099_U53);
  not ginst898 (P1_R2099_U170, P1_R2099_U15);
  not ginst899 (P1_R2099_U171, P1_R2099_U16);
  not ginst900 (P1_R2099_U172, P1_R2099_U17);
  not ginst901 (P1_R2099_U173, P1_R2099_U18);
  not ginst902 (P1_R2099_U174, P1_R2099_U19);
  not ginst903 (P1_R2099_U175, P1_R2099_U20);
  not ginst904 (P1_R2099_U176, P1_R2099_U21);
  not ginst905 (P1_R2099_U177, P1_R2099_U22);
  not ginst906 (P1_R2099_U178, P1_R2099_U23);
  not ginst907 (P1_R2099_U179, P1_R2099_U24);
  nand ginst908 (P1_R2099_U18, P1_R2099_U172, P1_R2099_U52);
  not ginst909 (P1_R2099_U180, P1_R2099_U25);
  not ginst910 (P1_R2099_U181, P1_R2099_U136);
  nand ginst911 (P1_R2099_U182, P1_R2099_U99, P1_U4190);
  nand ginst912 (P1_R2099_U183, P1_R2099_U4, P1_U2702);
  not ginst913 (P1_R2099_U184, P1_R2099_U27);
  nand ginst914 (P1_R2099_U185, P1_R2099_U100, P1_U4190);
  nand ginst915 (P1_R2099_U186, P1_R2099_U4, P1_U2710);
  not ginst916 (P1_R2099_U187, P1_R2099_U32);
  nand ginst917 (P1_R2099_U188, P1_R2099_U101, P1_U4190);
  nand ginst918 (P1_R2099_U189, P1_R2099_U4, P1_U2709);
  nand ginst919 (P1_R2099_U19, P1_R2099_U173, P1_R2099_U51);
  not ginst920 (P1_R2099_U190, P1_R2099_U33);
  nand ginst921 (P1_R2099_U191, P1_R2099_U102, P1_U4190);
  nand ginst922 (P1_R2099_U192, P1_R2099_U4, P1_U2708);
  not ginst923 (P1_R2099_U193, P1_R2099_U35);
  nand ginst924 (P1_R2099_U194, P1_R2099_U103, P1_U4190);
  nand ginst925 (P1_R2099_U195, P1_R2099_U4, P1_U2707);
  not ginst926 (P1_R2099_U196, P1_R2099_U34);
  nand ginst927 (P1_R2099_U197, P1_R2099_U104, P1_U4190);
  nand ginst928 (P1_R2099_U198, P1_R2099_U4, P1_U2706);
  not ginst929 (P1_R2099_U199, P1_R2099_U30);
  nand ginst930 (P1_R2099_U20, P1_R2099_U174, P1_R2099_U50);
  nand ginst931 (P1_R2099_U200, P1_R2099_U105, P1_U4190);
  nand ginst932 (P1_R2099_U201, P1_R2099_U4, P1_U2705);
  not ginst933 (P1_R2099_U202, P1_R2099_U31);
  nand ginst934 (P1_R2099_U203, P1_R2099_U106, P1_U4190);
  nand ginst935 (P1_R2099_U204, P1_R2099_U4, P1_U2704);
  not ginst936 (P1_R2099_U205, P1_R2099_U28);
  nand ginst937 (P1_R2099_U206, P1_R2099_U107, P1_U4190);
  nand ginst938 (P1_R2099_U207, P1_R2099_U4, P1_U2703);
  not ginst939 (P1_R2099_U208, P1_R2099_U29);
  nand ginst940 (P1_R2099_U209, P1_R2099_U108, P1_U4190);
  nand ginst941 (P1_R2099_U21, P1_R2099_U175, P1_R2099_U49);
  nand ginst942 (P1_R2099_U210, P1_R2099_U4, P1_U2701);
  not ginst943 (P1_R2099_U211, P1_R2099_U26);
  nand ginst944 (P1_R2099_U212, P1_R2099_U160, P1_R2099_U211);
  nand ginst945 (P1_R2099_U213, P1_R2099_U109, P1_R2099_U26);
  nand ginst946 (P1_R2099_U214, P1_R2099_U159, P1_R2099_U184);
  nand ginst947 (P1_R2099_U215, P1_R2099_U27, P1_R2099_U9);
  nand ginst948 (P1_R2099_U216, P1_R2099_U158, P1_R2099_U208);
  nand ginst949 (P1_R2099_U217, P1_R2099_U110, P1_R2099_U29);
  nand ginst950 (P1_R2099_U218, P1_R2099_U157, P1_R2099_U205);
  nand ginst951 (P1_R2099_U219, P1_R2099_U28, P1_R2099_U8);
  nand ginst952 (P1_R2099_U22, P1_R2099_U176, P1_R2099_U48);
  nand ginst953 (P1_R2099_U220, P1_R2099_U156, P1_R2099_U202);
  nand ginst954 (P1_R2099_U221, P1_R2099_U111, P1_R2099_U31);
  nand ginst955 (P1_R2099_U222, P1_R2099_U155, P1_R2099_U199);
  nand ginst956 (P1_R2099_U223, P1_R2099_U30, P1_R2099_U7);
  nand ginst957 (P1_R2099_U224, P1_R2099_U154, P1_R2099_U196);
  nand ginst958 (P1_R2099_U225, P1_R2099_U112, P1_R2099_U34);
  nand ginst959 (P1_R2099_U226, P1_R2099_U113, P1_U4190);
  nand ginst960 (P1_R2099_U227, P1_R2099_U4, P1_U2682);
  not ginst961 (P1_R2099_U228, P1_R2099_U45);
  nand ginst962 (P1_R2099_U229, P1_R2099_U114, P1_U4190);
  nand ginst963 (P1_R2099_U23, P1_R2099_U177, P1_R2099_U47);
  nand ginst964 (P1_R2099_U230, P1_R2099_U4, P1_U2683);
  not ginst965 (P1_R2099_U231, P1_R2099_U46);
  nand ginst966 (P1_R2099_U232, P1_R2099_U115, P1_U4190);
  nand ginst967 (P1_R2099_U233, P1_R2099_U4, P1_U2684);
  not ginst968 (P1_R2099_U234, P1_R2099_U47);
  nand ginst969 (P1_R2099_U235, P1_R2099_U116, P1_U4190);
  nand ginst970 (P1_R2099_U236, P1_R2099_U4, P1_U2685);
  not ginst971 (P1_R2099_U237, P1_R2099_U48);
  nand ginst972 (P1_R2099_U238, P1_R2099_U117, P1_U4190);
  nand ginst973 (P1_R2099_U239, P1_R2099_U4, P1_U2686);
  nand ginst974 (P1_R2099_U24, P1_R2099_U178, P1_R2099_U46);
  not ginst975 (P1_R2099_U240, P1_R2099_U49);
  nand ginst976 (P1_R2099_U241, P1_R2099_U118, P1_U4190);
  nand ginst977 (P1_R2099_U242, P1_R2099_U4, P1_U2687);
  not ginst978 (P1_R2099_U243, P1_R2099_U50);
  nand ginst979 (P1_R2099_U244, P1_R2099_U119, P1_U4190);
  nand ginst980 (P1_R2099_U245, P1_R2099_U4, P1_U2688);
  not ginst981 (P1_R2099_U246, P1_R2099_U51);
  nand ginst982 (P1_R2099_U247, P1_R2099_U120, P1_U4190);
  nand ginst983 (P1_R2099_U248, P1_R2099_U4, P1_U2689);
  not ginst984 (P1_R2099_U249, P1_R2099_U52);
  nand ginst985 (P1_R2099_U25, P1_R2099_U179, P1_R2099_U45);
  nand ginst986 (P1_R2099_U250, P1_R2099_U121, P1_U4190);
  nand ginst987 (P1_R2099_U251, P1_R2099_U4, P1_U2690);
  not ginst988 (P1_R2099_U252, P1_R2099_U53);
  nand ginst989 (P1_R2099_U253, P1_R2099_U122, P1_U4190);
  nand ginst990 (P1_R2099_U254, P1_R2099_U4, P1_U2691);
  not ginst991 (P1_R2099_U255, P1_R2099_U54);
  nand ginst992 (P1_R2099_U256, P1_R2099_U123, P1_U4190);
  nand ginst993 (P1_R2099_U257, P1_R2099_U4, P1_U2692);
  not ginst994 (P1_R2099_U258, P1_R2099_U55);
  nand ginst995 (P1_R2099_U259, P1_R2099_U124, P1_U4190);
  nand ginst996 (P1_R2099_U26, P1_R2099_U209, P1_R2099_U210);
  nand ginst997 (P1_R2099_U260, P1_R2099_U4, P1_U2700);
  not ginst998 (P1_R2099_U261, P1_R2099_U62);
  nand ginst999 (P1_R2099_U262, P1_R2099_U125, P1_U4190);
  nand ginst1000 (P1_R2099_U263, P1_R2099_U4, P1_U2699);
  not ginst1001 (P1_R2099_U264, P1_R2099_U63);
  nand ginst1002 (P1_R2099_U265, P1_R2099_U126, P1_U4190);
  nand ginst1003 (P1_R2099_U266, P1_R2099_U4, P1_U2698);
  not ginst1004 (P1_R2099_U267, P1_R2099_U60);
  nand ginst1005 (P1_R2099_U268, P1_R2099_U127, P1_U4190);
  nand ginst1006 (P1_R2099_U269, P1_R2099_U4, P1_U2697);
  nand ginst1007 (P1_R2099_U27, P1_R2099_U182, P1_R2099_U183);
  not ginst1008 (P1_R2099_U270, P1_R2099_U61);
  nand ginst1009 (P1_R2099_U271, P1_R2099_U128, P1_U4190);
  nand ginst1010 (P1_R2099_U272, P1_R2099_U4, P1_U2696);
  not ginst1011 (P1_R2099_U273, P1_R2099_U58);
  nand ginst1012 (P1_R2099_U274, P1_R2099_U129, P1_U4190);
  nand ginst1013 (P1_R2099_U275, P1_R2099_U4, P1_U2695);
  not ginst1014 (P1_R2099_U276, P1_R2099_U59);
  nand ginst1015 (P1_R2099_U277, P1_R2099_U130, P1_U4190);
  nand ginst1016 (P1_R2099_U278, P1_R2099_U4, P1_U2694);
  not ginst1017 (P1_R2099_U279, P1_R2099_U56);
  nand ginst1018 (P1_R2099_U28, P1_R2099_U203, P1_R2099_U204);
  nand ginst1019 (P1_R2099_U280, P1_R2099_U131, P1_U4190);
  nand ginst1020 (P1_R2099_U281, P1_R2099_U4, P1_U2693);
  not ginst1021 (P1_R2099_U282, P1_R2099_U57);
  nand ginst1022 (P1_R2099_U283, P1_R2099_U132, P1_U4190);
  nand ginst1023 (P1_R2099_U284, P1_R2099_U4, P1_U2680);
  not ginst1024 (P1_R2099_U285, P1_R2099_U43);
  nand ginst1025 (P1_R2099_U286, P1_R2099_U133, P1_U4190);
  nand ginst1026 (P1_R2099_U287, P1_R2099_U4, P1_U2681);
  not ginst1027 (P1_R2099_U288, P1_R2099_U44);
  nand ginst1028 (P1_R2099_U289, P1_R2099_U134, P1_U4190);
  nand ginst1029 (P1_R2099_U29, P1_R2099_U206, P1_R2099_U207);
  nand ginst1030 (P1_R2099_U290, P1_R2099_U4, P1_U2679);
  not ginst1031 (P1_R2099_U291, P1_R2099_U97);
  nand ginst1032 (P1_R2099_U292, P1_R2099_U145, P1_R2099_U291);
  nand ginst1033 (P1_R2099_U293, P1_R2099_U135, P1_R2099_U97);
  nand ginst1034 (P1_R2099_U294, P1_R2099_U181, P1_R2099_U285);
  nand ginst1035 (P1_R2099_U295, P1_R2099_U136, P1_R2099_U43);
  nand ginst1036 (P1_R2099_U296, P1_R2099_U153, P1_R2099_U193);
  nand ginst1037 (P1_R2099_U297, P1_R2099_U137, P1_R2099_U35);
  nand ginst1038 (P1_R2099_U298, P1_R2099_U180, P1_R2099_U288);
  nand ginst1039 (P1_R2099_U299, P1_R2099_U25, P1_R2099_U44);
  nand ginst1040 (P1_R2099_U30, P1_R2099_U197, P1_R2099_U198);
  nand ginst1041 (P1_R2099_U300, P1_R2099_U179, P1_R2099_U228);
  nand ginst1042 (P1_R2099_U301, P1_R2099_U24, P1_R2099_U45);
  nand ginst1043 (P1_R2099_U302, P1_R2099_U178, P1_R2099_U231);
  nand ginst1044 (P1_R2099_U303, P1_R2099_U23, P1_R2099_U46);
  nand ginst1045 (P1_R2099_U304, P1_R2099_U177, P1_R2099_U234);
  nand ginst1046 (P1_R2099_U305, P1_R2099_U22, P1_R2099_U47);
  nand ginst1047 (P1_R2099_U306, P1_R2099_U176, P1_R2099_U237);
  nand ginst1048 (P1_R2099_U307, P1_R2099_U21, P1_R2099_U48);
  nand ginst1049 (P1_R2099_U308, P1_R2099_U175, P1_R2099_U240);
  nand ginst1050 (P1_R2099_U309, P1_R2099_U20, P1_R2099_U49);
  nand ginst1051 (P1_R2099_U31, P1_R2099_U200, P1_R2099_U201);
  nand ginst1052 (P1_R2099_U310, P1_R2099_U174, P1_R2099_U243);
  nand ginst1053 (P1_R2099_U311, P1_R2099_U19, P1_R2099_U50);
  nand ginst1054 (P1_R2099_U312, P1_R2099_U173, P1_R2099_U246);
  nand ginst1055 (P1_R2099_U313, P1_R2099_U18, P1_R2099_U51);
  nand ginst1056 (P1_R2099_U314, P1_R2099_U172, P1_R2099_U249);
  nand ginst1057 (P1_R2099_U315, P1_R2099_U17, P1_R2099_U52);
  nand ginst1058 (P1_R2099_U316, P1_R2099_U171, P1_R2099_U252);
  nand ginst1059 (P1_R2099_U317, P1_R2099_U16, P1_R2099_U53);
  nand ginst1060 (P1_R2099_U318, P1_R2099_U190, P1_U2678);
  nand ginst1061 (P1_R2099_U319, P1_R2099_U33, P1_R2099_U6);
  nand ginst1062 (P1_R2099_U32, P1_R2099_U185, P1_R2099_U186);
  nand ginst1063 (P1_R2099_U320, P1_R2099_U190, P1_U2678);
  nand ginst1064 (P1_R2099_U321, P1_R2099_U33, P1_R2099_U6);
  nand ginst1065 (P1_R2099_U322, P1_R2099_U320, P1_R2099_U321);
  nand ginst1066 (P1_R2099_U323, P1_R2099_U139, P1_R2099_U140);
  nand ginst1067 (P1_R2099_U324, P1_R2099_U149, P1_R2099_U322);
  nand ginst1068 (P1_R2099_U325, P1_R2099_U170, P1_R2099_U255);
  nand ginst1069 (P1_R2099_U326, P1_R2099_U15, P1_R2099_U54);
  nand ginst1070 (P1_R2099_U327, P1_R2099_U169, P1_R2099_U258);
  nand ginst1071 (P1_R2099_U328, P1_R2099_U14, P1_R2099_U55);
  nand ginst1072 (P1_R2099_U329, P1_R2099_U168, P1_R2099_U282);
  nand ginst1073 (P1_R2099_U33, P1_R2099_U188, P1_R2099_U189);
  nand ginst1074 (P1_R2099_U330, P1_R2099_U141, P1_R2099_U57);
  nand ginst1075 (P1_R2099_U331, P1_R2099_U167, P1_R2099_U279);
  nand ginst1076 (P1_R2099_U332, P1_R2099_U13, P1_R2099_U56);
  nand ginst1077 (P1_R2099_U333, P1_R2099_U166, P1_R2099_U276);
  nand ginst1078 (P1_R2099_U334, P1_R2099_U142, P1_R2099_U59);
  nand ginst1079 (P1_R2099_U335, P1_R2099_U165, P1_R2099_U273);
  nand ginst1080 (P1_R2099_U336, P1_R2099_U12, P1_R2099_U58);
  nand ginst1081 (P1_R2099_U337, P1_R2099_U164, P1_R2099_U270);
  nand ginst1082 (P1_R2099_U338, P1_R2099_U143, P1_R2099_U61);
  nand ginst1083 (P1_R2099_U339, P1_R2099_U163, P1_R2099_U267);
  nand ginst1084 (P1_R2099_U34, P1_R2099_U194, P1_R2099_U195);
  nand ginst1085 (P1_R2099_U340, P1_R2099_U11, P1_R2099_U60);
  nand ginst1086 (P1_R2099_U341, P1_R2099_U162, P1_R2099_U264);
  nand ginst1087 (P1_R2099_U342, P1_R2099_U144, P1_R2099_U63);
  nand ginst1088 (P1_R2099_U343, P1_R2099_U161, P1_R2099_U261);
  nand ginst1089 (P1_R2099_U344, P1_R2099_U10, P1_R2099_U62);
  nand ginst1090 (P1_R2099_U345, P1_R2099_U4, P1_U4189);
  nand ginst1091 (P1_R2099_U346, P1_R2099_U5, P1_U4190);
  not ginst1092 (P1_R2099_U347, P1_R2099_U98);
  nand ginst1093 (P1_R2099_U348, P1_R2099_U32, P1_R2099_U347);
  nand ginst1094 (P1_R2099_U349, P1_R2099_U187, P1_R2099_U98);
  nand ginst1095 (P1_R2099_U35, P1_R2099_U191, P1_R2099_U192);
  nand ginst1096 (P1_R2099_U36, P1_R2099_U212, P1_R2099_U213);
  nand ginst1097 (P1_R2099_U37, P1_R2099_U214, P1_R2099_U215);
  nand ginst1098 (P1_R2099_U38, P1_R2099_U216, P1_R2099_U217);
  nand ginst1099 (P1_R2099_U39, P1_R2099_U218, P1_R2099_U219);
  not ginst1100 (P1_R2099_U4, P1_U4190);
  nand ginst1101 (P1_R2099_U40, P1_R2099_U220, P1_R2099_U221);
  nand ginst1102 (P1_R2099_U41, P1_R2099_U222, P1_R2099_U223);
  nand ginst1103 (P1_R2099_U42, P1_R2099_U224, P1_R2099_U225);
  nand ginst1104 (P1_R2099_U43, P1_R2099_U283, P1_R2099_U284);
  nand ginst1105 (P1_R2099_U44, P1_R2099_U286, P1_R2099_U287);
  nand ginst1106 (P1_R2099_U45, P1_R2099_U226, P1_R2099_U227);
  nand ginst1107 (P1_R2099_U46, P1_R2099_U229, P1_R2099_U230);
  nand ginst1108 (P1_R2099_U47, P1_R2099_U232, P1_R2099_U233);
  nand ginst1109 (P1_R2099_U48, P1_R2099_U235, P1_R2099_U236);
  nand ginst1110 (P1_R2099_U49, P1_R2099_U238, P1_R2099_U239);
  not ginst1111 (P1_R2099_U5, P1_U4189);
  nand ginst1112 (P1_R2099_U50, P1_R2099_U241, P1_R2099_U242);
  nand ginst1113 (P1_R2099_U51, P1_R2099_U244, P1_R2099_U245);
  nand ginst1114 (P1_R2099_U52, P1_R2099_U247, P1_R2099_U248);
  nand ginst1115 (P1_R2099_U53, P1_R2099_U250, P1_R2099_U251);
  nand ginst1116 (P1_R2099_U54, P1_R2099_U253, P1_R2099_U254);
  nand ginst1117 (P1_R2099_U55, P1_R2099_U256, P1_R2099_U257);
  nand ginst1118 (P1_R2099_U56, P1_R2099_U277, P1_R2099_U278);
  nand ginst1119 (P1_R2099_U57, P1_R2099_U280, P1_R2099_U281);
  nand ginst1120 (P1_R2099_U58, P1_R2099_U271, P1_R2099_U272);
  nand ginst1121 (P1_R2099_U59, P1_R2099_U274, P1_R2099_U275);
  not ginst1122 (P1_R2099_U6, P1_U2678);
  nand ginst1123 (P1_R2099_U60, P1_R2099_U265, P1_R2099_U266);
  nand ginst1124 (P1_R2099_U61, P1_R2099_U268, P1_R2099_U269);
  nand ginst1125 (P1_R2099_U62, P1_R2099_U259, P1_R2099_U260);
  nand ginst1126 (P1_R2099_U63, P1_R2099_U262, P1_R2099_U263);
  nand ginst1127 (P1_R2099_U64, P1_R2099_U292, P1_R2099_U293);
  nand ginst1128 (P1_R2099_U65, P1_R2099_U294, P1_R2099_U295);
  nand ginst1129 (P1_R2099_U66, P1_R2099_U298, P1_R2099_U299);
  nand ginst1130 (P1_R2099_U67, P1_R2099_U300, P1_R2099_U301);
  nand ginst1131 (P1_R2099_U68, P1_R2099_U302, P1_R2099_U303);
  nand ginst1132 (P1_R2099_U69, P1_R2099_U304, P1_R2099_U305);
  nand ginst1133 (P1_R2099_U7, P1_R2099_U137, P1_R2099_U88);
  nand ginst1134 (P1_R2099_U70, P1_R2099_U306, P1_R2099_U307);
  nand ginst1135 (P1_R2099_U71, P1_R2099_U308, P1_R2099_U309);
  nand ginst1136 (P1_R2099_U72, P1_R2099_U310, P1_R2099_U311);
  nand ginst1137 (P1_R2099_U73, P1_R2099_U312, P1_R2099_U313);
  nand ginst1138 (P1_R2099_U74, P1_R2099_U314, P1_R2099_U315);
  nand ginst1139 (P1_R2099_U75, P1_R2099_U316, P1_R2099_U317);
  nand ginst1140 (P1_R2099_U76, P1_R2099_U325, P1_R2099_U326);
  nand ginst1141 (P1_R2099_U77, P1_R2099_U327, P1_R2099_U328);
  nand ginst1142 (P1_R2099_U78, P1_R2099_U329, P1_R2099_U330);
  nand ginst1143 (P1_R2099_U79, P1_R2099_U331, P1_R2099_U332);
  nand ginst1144 (P1_R2099_U8, P1_R2099_U155, P1_R2099_U89);
  nand ginst1145 (P1_R2099_U80, P1_R2099_U333, P1_R2099_U334);
  nand ginst1146 (P1_R2099_U81, P1_R2099_U335, P1_R2099_U336);
  nand ginst1147 (P1_R2099_U82, P1_R2099_U337, P1_R2099_U338);
  nand ginst1148 (P1_R2099_U83, P1_R2099_U339, P1_R2099_U340);
  nand ginst1149 (P1_R2099_U84, P1_R2099_U341, P1_R2099_U342);
  nand ginst1150 (P1_R2099_U85, P1_R2099_U343, P1_R2099_U344);
  nand ginst1151 (P1_R2099_U86, P1_R2099_U348, P1_R2099_U349);
  nand ginst1152 (P1_R2099_U87, P1_R2099_U323, P1_R2099_U324);
  and ginst1153 (P1_R2099_U88, P1_R2099_U34, P1_R2099_U35);
  and ginst1154 (P1_R2099_U89, P1_R2099_U30, P1_R2099_U31);
  nand ginst1155 (P1_R2099_U9, P1_R2099_U157, P1_R2099_U90);
  and ginst1156 (P1_R2099_U90, P1_R2099_U28, P1_R2099_U29);
  and ginst1157 (P1_R2099_U91, P1_R2099_U26, P1_R2099_U27);
  and ginst1158 (P1_R2099_U92, P1_R2099_U62, P1_R2099_U63);
  and ginst1159 (P1_R2099_U93, P1_R2099_U60, P1_R2099_U61);
  and ginst1160 (P1_R2099_U94, P1_R2099_U58, P1_R2099_U59);
  and ginst1161 (P1_R2099_U95, P1_R2099_U56, P1_R2099_U57);
  and ginst1162 (P1_R2099_U96, P1_R2099_U43, P1_R2099_U44);
  nand ginst1163 (P1_R2099_U97, P1_R2099_U289, P1_R2099_U290);
  nand ginst1164 (P1_R2099_U98, P1_R2099_U345, P1_R2099_U346);
  not ginst1165 (P1_R2099_U99, P1_U2702);
  and ginst1166 (P1_R2144_U10, P1_R2144_U212, P1_R2144_U213, P1_R2144_U82);
  nand ginst1167 (P1_R2144_U100, P1_R2144_U28, P1_U2751);
  not ginst1168 (P1_R2144_U101, P1_R2144_U24);
  not ginst1169 (P1_R2144_U102, P1_R2144_U81);
  nand ginst1170 (P1_R2144_U103, P1_R2144_U181, P1_U2745);
  nand ginst1171 (P1_R2144_U104, P1_R2144_U166, P1_R2144_U167, P1_R2144_U17);
  nand ginst1172 (P1_R2144_U105, P1_R2144_U174, P1_R2144_U175, P1_R2144_U20);
  nand ginst1173 (P1_R2144_U106, P1_R2144_U18, P1_R2144_U200, P1_R2144_U201);
  not ginst1174 (P1_R2144_U107, P1_R2144_U21);
  not ginst1175 (P1_R2144_U108, P1_R2144_U23);
  nand ginst1176 (P1_R2144_U109, P1_R2144_U13, P1_R2144_U193, P1_R2144_U194);
  nand ginst1177 (P1_R2144_U11, P1_R2144_U144, P1_R2144_U146);
  nand ginst1178 (P1_R2144_U110, P1_R2144_U16, P1_R2144_U195, P1_R2144_U196);
  nand ginst1179 (P1_R2144_U111, P1_R2144_U199, P1_U2749);
  nand ginst1180 (P1_R2144_U112, P1_R2144_U15, P1_R2144_U188, P1_R2144_U189);
  nand ginst1181 (P1_R2144_U113, P1_R2144_U192, P1_U2752);
  nand ginst1182 (P1_R2144_U114, P1_R2144_U14, P1_R2144_U187);
  nand ginst1183 (P1_R2144_U115, P1_R2144_U112, P1_U2355);
  nand ginst1184 (P1_R2144_U116, P1_R2144_U184, P1_U2750);
  nand ginst1185 (P1_R2144_U117, P1_R2144_U155, P1_R2144_U157);
  nand ginst1186 (P1_R2144_U118, P1_R2144_U117, P1_R2144_U51);
  not ginst1187 (P1_R2144_U119, P1_R2144_U84);
  not ginst1188 (P1_R2144_U12, P1_U2355);
  not ginst1189 (P1_R2144_U120, P1_R2144_U19);
  not ginst1190 (P1_R2144_U121, P1_R2144_U79);
  not ginst1191 (P1_R2144_U122, P1_R2144_U78);
  not ginst1192 (P1_R2144_U123, P1_R2144_U83);
  nand ginst1193 (P1_R2144_U124, P1_R2144_U105, P1_R2144_U83);
  nand ginst1194 (P1_R2144_U125, P1_R2144_U124, P1_R2144_U21);
  nand ginst1195 (P1_R2144_U126, P1_R2144_U23, P1_R2144_U81);
  nand ginst1196 (P1_R2144_U127, P1_R2144_U124, P1_R2144_U60);
  nand ginst1197 (P1_R2144_U128, P1_R2144_U125, P1_R2144_U61);
  nand ginst1198 (P1_R2144_U129, P1_R2144_U112, P1_U2355);
  not ginst1199 (P1_R2144_U13, P1_U2750);
  not ginst1200 (P1_R2144_U130, P1_R2144_U93);
  nand ginst1201 (P1_R2144_U131, P1_R2144_U14, P1_R2144_U187);
  nand ginst1202 (P1_R2144_U132, P1_R2144_U131, P1_R2144_U93);
  not ginst1203 (P1_R2144_U133, P1_R2144_U91);
  nand ginst1204 (P1_R2144_U134, P1_R2144_U109, P1_R2144_U91);
  nand ginst1205 (P1_R2144_U135, P1_R2144_U116, P1_R2144_U134);
  nand ginst1206 (P1_R2144_U136, P1_R2144_U135, P1_R2144_U62);
  nand ginst1207 (P1_R2144_U137, P1_R2144_U110, P1_R2144_U161);
  nand ginst1208 (P1_R2144_U138, P1_R2144_U116, P1_R2144_U134, P1_R2144_U137);
  not ginst1209 (P1_R2144_U139, P1_R2144_U97);
  not ginst1210 (P1_R2144_U14, P1_U2751);
  not ginst1211 (P1_R2144_U140, P1_R2144_U96);
  not ginst1212 (P1_R2144_U141, P1_R2144_U25);
  not ginst1213 (P1_R2144_U142, P1_R2144_U95);
  not ginst1214 (P1_R2144_U143, P1_R2144_U26);
  nand ginst1215 (P1_R2144_U144, P1_R2144_U24, P1_U2355);
  not ginst1216 (P1_R2144_U145, P1_R2144_U144);
  nand ginst1217 (P1_R2144_U146, P1_R2144_U101, P1_R2144_U12);
  not ginst1218 (P1_R2144_U147, P1_R2144_U94);
  not ginst1219 (P1_R2144_U148, P1_R2144_U98);
  nand ginst1220 (P1_R2144_U149, P1_R2144_U105, P1_R2144_U21);
  not ginst1221 (P1_R2144_U15, P1_U2752);
  nand ginst1222 (P1_R2144_U150, P1_R2144_U106, P1_R2144_U19);
  nand ginst1223 (P1_R2144_U151, P1_R2144_U105, P1_R2144_U120, P1_R2144_U7);
  nand ginst1224 (P1_R2144_U152, P1_R2144_U107, P1_R2144_U7);
  nand ginst1225 (P1_R2144_U153, P1_R2144_U108, P1_R2144_U7);
  nand ginst1226 (P1_R2144_U154, P1_R2144_U100, P1_R2144_U113, P1_R2144_U115);
  nand ginst1227 (P1_R2144_U155, P1_R2144_U114, P1_R2144_U154);
  nand ginst1228 (P1_R2144_U156, P1_R2144_U103, P1_R2144_U104);
  nand ginst1229 (P1_R2144_U157, P1_R2144_U184, P1_U2750);
  nand ginst1230 (P1_R2144_U158, P1_R2144_U110, P1_R2144_U117, P1_R2144_U55);
  nand ginst1231 (P1_R2144_U159, P1_R2144_U106, P1_R2144_U199, P1_U2749);
  not ginst1232 (P1_R2144_U16, P1_U2749);
  nand ginst1233 (P1_R2144_U160, P1_R2144_U158, P1_R2144_U58);
  nand ginst1234 (P1_R2144_U161, P1_R2144_U199, P1_U2749);
  nand ginst1235 (P1_R2144_U162, P1_R2144_U184, P1_U2750);
  nand ginst1236 (P1_R2144_U163, P1_R2144_U109, P1_R2144_U116);
  nand ginst1237 (P1_R2144_U164, P1_R2144_U68, P1_U2355);
  nand ginst1238 (P1_R2144_U165, P1_R2144_U12, P1_U2762);
  nand ginst1239 (P1_R2144_U166, P1_R2144_U69, P1_U2355);
  nand ginst1240 (P1_R2144_U167, P1_R2144_U12, P1_U2761);
  nand ginst1241 (P1_R2144_U168, P1_R2144_U70, P1_U2355);
  nand ginst1242 (P1_R2144_U169, P1_R2144_U12, P1_U2763);
  not ginst1243 (P1_R2144_U17, P1_U2745);
  nand ginst1244 (P1_R2144_U170, P1_R2144_U168, P1_R2144_U169);
  nand ginst1245 (P1_R2144_U171, P1_R2144_U68, P1_U2355);
  nand ginst1246 (P1_R2144_U172, P1_R2144_U12, P1_U2762);
  nand ginst1247 (P1_R2144_U173, P1_R2144_U171, P1_R2144_U172);
  nand ginst1248 (P1_R2144_U174, P1_R2144_U70, P1_U2355);
  nand ginst1249 (P1_R2144_U175, P1_R2144_U12, P1_U2763);
  nand ginst1250 (P1_R2144_U176, P1_R2144_U71, P1_U2355);
  nand ginst1251 (P1_R2144_U177, P1_R2144_U12, P1_U2764);
  nand ginst1252 (P1_R2144_U178, P1_R2144_U176, P1_R2144_U177);
  nand ginst1253 (P1_R2144_U179, P1_R2144_U69, P1_U2355);
  not ginst1254 (P1_R2144_U18, P1_U2748);
  nand ginst1255 (P1_R2144_U180, P1_R2144_U12, P1_U2761);
  nand ginst1256 (P1_R2144_U181, P1_R2144_U179, P1_R2144_U180);
  nand ginst1257 (P1_R2144_U182, P1_R2144_U72, P1_U2355);
  nand ginst1258 (P1_R2144_U183, P1_R2144_U12, P1_U2766);
  nand ginst1259 (P1_R2144_U184, P1_R2144_U182, P1_R2144_U183);
  nand ginst1260 (P1_R2144_U185, P1_R2144_U73, P1_U2355);
  nand ginst1261 (P1_R2144_U186, P1_R2144_U12, P1_U2767);
  not ginst1262 (P1_R2144_U187, P1_R2144_U28);
  nand ginst1263 (P1_R2144_U188, P1_R2144_U74, P1_U2355);
  nand ginst1264 (P1_R2144_U189, P1_R2144_U12, P1_U2768);
  nand ginst1265 (P1_R2144_U19, P1_R2144_U178, P1_U2748);
  nand ginst1266 (P1_R2144_U190, P1_R2144_U74, P1_U2355);
  nand ginst1267 (P1_R2144_U191, P1_R2144_U12, P1_U2768);
  nand ginst1268 (P1_R2144_U192, P1_R2144_U190, P1_R2144_U191);
  nand ginst1269 (P1_R2144_U193, P1_R2144_U72, P1_U2355);
  nand ginst1270 (P1_R2144_U194, P1_R2144_U12, P1_U2766);
  nand ginst1271 (P1_R2144_U195, P1_R2144_U75, P1_U2355);
  nand ginst1272 (P1_R2144_U196, P1_R2144_U12, P1_U2765);
  nand ginst1273 (P1_R2144_U197, P1_R2144_U75, P1_U2355);
  nand ginst1274 (P1_R2144_U198, P1_R2144_U12, P1_U2765);
  nand ginst1275 (P1_R2144_U199, P1_R2144_U197, P1_R2144_U198);
  not ginst1276 (P1_R2144_U20, P1_U2747);
  nand ginst1277 (P1_R2144_U200, P1_R2144_U71, P1_U2355);
  nand ginst1278 (P1_R2144_U201, P1_R2144_U12, P1_U2764);
  nand ginst1279 (P1_R2144_U202, P1_R2144_U76, P1_U2355);
  nand ginst1280 (P1_R2144_U203, P1_R2144_U12, P1_U2760);
  not ginst1281 (P1_R2144_U204, P1_R2144_U29);
  nand ginst1282 (P1_R2144_U205, P1_R2144_U77, P1_U2355);
  nand ginst1283 (P1_R2144_U206, P1_R2144_U12, P1_U2759);
  not ginst1284 (P1_R2144_U207, P1_R2144_U27);
  nand ginst1285 (P1_R2144_U208, P1_R2144_U122, P1_R2144_U207);
  nand ginst1286 (P1_R2144_U209, P1_R2144_U27, P1_R2144_U78);
  nand ginst1287 (P1_R2144_U21, P1_R2144_U170, P1_U2747);
  nand ginst1288 (P1_R2144_U210, P1_R2144_U121, P1_R2144_U204);
  nand ginst1289 (P1_R2144_U211, P1_R2144_U29, P1_R2144_U79);
  nand ginst1290 (P1_R2144_U212, P1_R2144_U124, P1_R2144_U23, P1_R2144_U57);
  nand ginst1291 (P1_R2144_U213, P1_R2144_U108, P1_R2144_U5);
  nand ginst1292 (P1_R2144_U214, P1_R2144_U102, P1_R2144_U156);
  nand ginst1293 (P1_R2144_U215, P1_R2144_U160, P1_R2144_U59, P1_R2144_U81);
  nand ginst1294 (P1_R2144_U216, P1_R2144_U149, P1_R2144_U83);
  nand ginst1295 (P1_R2144_U217, P1_R2144_U123, P1_R2144_U44);
  nand ginst1296 (P1_R2144_U218, P1_R2144_U150, P1_R2144_U84);
  nand ginst1297 (P1_R2144_U219, P1_R2144_U119, P1_R2144_U46);
  not ginst1298 (P1_R2144_U22, P1_U2746);
  nand ginst1299 (P1_R2144_U220, P1_R2144_U85, P1_U2355);
  nand ginst1300 (P1_R2144_U221, P1_R2144_U12, P1_U2754);
  not ginst1301 (P1_R2144_U222, P1_R2144_U32);
  nand ginst1302 (P1_R2144_U223, P1_R2144_U86, P1_U2355);
  nand ginst1303 (P1_R2144_U224, P1_R2144_U12, P1_U2753);
  not ginst1304 (P1_R2144_U225, P1_R2144_U31);
  nand ginst1305 (P1_R2144_U226, P1_R2144_U87, P1_U2355);
  nand ginst1306 (P1_R2144_U227, P1_R2144_U12, P1_U2755);
  not ginst1307 (P1_R2144_U228, P1_R2144_U33);
  nand ginst1308 (P1_R2144_U229, P1_R2144_U88, P1_U2355);
  nand ginst1309 (P1_R2144_U23, P1_R2144_U173, P1_U2746);
  nand ginst1310 (P1_R2144_U230, P1_R2144_U12, P1_U2756);
  not ginst1311 (P1_R2144_U231, P1_R2144_U34);
  nand ginst1312 (P1_R2144_U232, P1_R2144_U89, P1_U2355);
  nand ginst1313 (P1_R2144_U233, P1_R2144_U12, P1_U2757);
  not ginst1314 (P1_R2144_U234, P1_R2144_U35);
  nand ginst1315 (P1_R2144_U235, P1_R2144_U90, P1_U2355);
  nand ginst1316 (P1_R2144_U236, P1_R2144_U12, P1_U2758);
  not ginst1317 (P1_R2144_U237, P1_R2144_U36);
  nand ginst1318 (P1_R2144_U238, P1_R2144_U163, P1_R2144_U91);
  nand ginst1319 (P1_R2144_U239, P1_R2144_U133, P1_R2144_U48);
  nand ginst1320 (P1_R2144_U24, P1_R2144_U63, P1_R2144_U79);
  nand ginst1321 (P1_R2144_U240, P1_R2144_U187, P1_U2751);
  nand ginst1322 (P1_R2144_U241, P1_R2144_U14, P1_R2144_U28);
  nand ginst1323 (P1_R2144_U242, P1_R2144_U187, P1_U2751);
  nand ginst1324 (P1_R2144_U243, P1_R2144_U14, P1_R2144_U28);
  nand ginst1325 (P1_R2144_U244, P1_R2144_U242, P1_R2144_U243);
  nand ginst1326 (P1_R2144_U245, P1_R2144_U92, P1_R2144_U93);
  nand ginst1327 (P1_R2144_U246, P1_R2144_U130, P1_R2144_U244);
  nand ginst1328 (P1_R2144_U247, P1_R2144_U147, P1_R2144_U225);
  nand ginst1329 (P1_R2144_U248, P1_R2144_U31, P1_R2144_U94);
  nand ginst1330 (P1_R2144_U249, P1_R2144_U143, P1_R2144_U222);
  nand ginst1331 (P1_R2144_U25, P1_R2144_U6, P1_R2144_U79);
  nand ginst1332 (P1_R2144_U250, P1_R2144_U26, P1_R2144_U32);
  nand ginst1333 (P1_R2144_U251, P1_R2144_U142, P1_R2144_U228);
  nand ginst1334 (P1_R2144_U252, P1_R2144_U33, P1_R2144_U95);
  nand ginst1335 (P1_R2144_U253, P1_R2144_U141, P1_R2144_U231);
  nand ginst1336 (P1_R2144_U254, P1_R2144_U25, P1_R2144_U34);
  nand ginst1337 (P1_R2144_U255, P1_R2144_U140, P1_R2144_U234);
  nand ginst1338 (P1_R2144_U256, P1_R2144_U35, P1_R2144_U96);
  nand ginst1339 (P1_R2144_U257, P1_R2144_U139, P1_R2144_U237);
  nand ginst1340 (P1_R2144_U258, P1_R2144_U36, P1_R2144_U97);
  nand ginst1341 (P1_R2144_U259, P1_R2144_U98, P1_U2355);
  nand ginst1342 (P1_R2144_U26, P1_R2144_U141, P1_R2144_U65);
  nand ginst1343 (P1_R2144_U260, P1_R2144_U12, P1_R2144_U148);
  nand ginst1344 (P1_R2144_U27, P1_R2144_U205, P1_R2144_U206);
  nand ginst1345 (P1_R2144_U28, P1_R2144_U185, P1_R2144_U186);
  nand ginst1346 (P1_R2144_U29, P1_R2144_U202, P1_R2144_U203);
  nand ginst1347 (P1_R2144_U30, P1_R2144_U208, P1_R2144_U209);
  nand ginst1348 (P1_R2144_U31, P1_R2144_U223, P1_R2144_U224);
  nand ginst1349 (P1_R2144_U32, P1_R2144_U220, P1_R2144_U221);
  nand ginst1350 (P1_R2144_U33, P1_R2144_U226, P1_R2144_U227);
  nand ginst1351 (P1_R2144_U34, P1_R2144_U229, P1_R2144_U230);
  nand ginst1352 (P1_R2144_U35, P1_R2144_U232, P1_R2144_U233);
  nand ginst1353 (P1_R2144_U36, P1_R2144_U235, P1_R2144_U236);
  nand ginst1354 (P1_R2144_U37, P1_R2144_U247, P1_R2144_U248);
  nand ginst1355 (P1_R2144_U38, P1_R2144_U249, P1_R2144_U250);
  nand ginst1356 (P1_R2144_U39, P1_R2144_U251, P1_R2144_U252);
  nand ginst1357 (P1_R2144_U40, P1_R2144_U253, P1_R2144_U254);
  nand ginst1358 (P1_R2144_U41, P1_R2144_U255, P1_R2144_U256);
  nand ginst1359 (P1_R2144_U42, P1_R2144_U257, P1_R2144_U258);
  nand ginst1360 (P1_R2144_U43, P1_R2144_U259, P1_R2144_U260);
  and ginst1361 (P1_R2144_U44, P1_R2144_U105, P1_R2144_U21);
  nand ginst1362 (P1_R2144_U45, P1_R2144_U216, P1_R2144_U217);
  and ginst1363 (P1_R2144_U46, P1_R2144_U106, P1_R2144_U19);
  nand ginst1364 (P1_R2144_U47, P1_R2144_U218, P1_R2144_U219);
  and ginst1365 (P1_R2144_U48, P1_R2144_U109, P1_R2144_U162);
  nand ginst1366 (P1_R2144_U49, P1_R2144_U238, P1_R2144_U239);
  and ginst1367 (P1_R2144_U5, P1_R2144_U103, P1_R2144_U104);
  nand ginst1368 (P1_R2144_U50, P1_R2144_U245, P1_R2144_U246);
  and ginst1369 (P1_R2144_U51, P1_R2144_U109, P1_R2144_U110);
  and ginst1370 (P1_R2144_U52, P1_R2144_U105, P1_R2144_U106);
  and ginst1371 (P1_R2144_U53, P1_R2144_U52, P1_R2144_U7);
  and ginst1372 (P1_R2144_U54, P1_R2144_U103, P1_R2144_U151, P1_R2144_U152, P1_R2144_U153);
  and ginst1373 (P1_R2144_U55, P1_R2144_U106, P1_R2144_U109);
  and ginst1374 (P1_R2144_U56, P1_R2144_U159, P1_R2144_U19);
  and ginst1375 (P1_R2144_U57, P1_R2144_U156, P1_R2144_U21);
  and ginst1376 (P1_R2144_U58, P1_R2144_U159, P1_R2144_U19, P1_R2144_U21);
  and ginst1377 (P1_R2144_U59, P1_R2144_U105, P1_R2144_U5);
  and ginst1378 (P1_R2144_U6, P1_R2144_U27, P1_R2144_U29, P1_R2144_U35, P1_R2144_U36);
  and ginst1379 (P1_R2144_U60, P1_R2144_U126, P1_R2144_U21);
  and ginst1380 (P1_R2144_U61, P1_R2144_U23, P1_R2144_U81);
  and ginst1381 (P1_R2144_U62, P1_R2144_U110, P1_R2144_U111);
  and ginst1382 (P1_R2144_U63, P1_R2144_U6, P1_R2144_U64);
  and ginst1383 (P1_R2144_U64, P1_R2144_U31, P1_R2144_U32, P1_R2144_U33, P1_R2144_U34);
  and ginst1384 (P1_R2144_U65, P1_R2144_U33, P1_R2144_U34);
  and ginst1385 (P1_R2144_U66, P1_R2144_U27, P1_R2144_U29, P1_R2144_U36);
  and ginst1386 (P1_R2144_U67, P1_R2144_U27, P1_R2144_U29);
  not ginst1387 (P1_R2144_U68, P1_U2762);
  not ginst1388 (P1_R2144_U69, P1_U2761);
  and ginst1389 (P1_R2144_U7, P1_R2144_U104, P1_R2144_U81);
  not ginst1390 (P1_R2144_U70, P1_U2763);
  not ginst1391 (P1_R2144_U71, P1_U2764);
  not ginst1392 (P1_R2144_U72, P1_U2766);
  not ginst1393 (P1_R2144_U73, P1_U2767);
  not ginst1394 (P1_R2144_U74, P1_U2768);
  not ginst1395 (P1_R2144_U75, P1_U2765);
  not ginst1396 (P1_R2144_U76, P1_U2760);
  not ginst1397 (P1_R2144_U77, P1_U2759);
  nand ginst1398 (P1_R2144_U78, P1_R2144_U29, P1_R2144_U79);
  nand ginst1399 (P1_R2144_U79, P1_R2144_U54, P1_R2144_U99);
  and ginst1400 (P1_R2144_U8, P1_R2144_U136, P1_R2144_U138);
  and ginst1401 (P1_R2144_U80, P1_R2144_U210, P1_R2144_U211);
  nand ginst1402 (P1_R2144_U81, P1_R2144_U164, P1_R2144_U165, P1_R2144_U22);
  and ginst1403 (P1_R2144_U82, P1_R2144_U214, P1_R2144_U215);
  nand ginst1404 (P1_R2144_U83, P1_R2144_U158, P1_R2144_U56);
  nand ginst1405 (P1_R2144_U84, P1_R2144_U111, P1_R2144_U118);
  not ginst1406 (P1_R2144_U85, P1_U2754);
  not ginst1407 (P1_R2144_U86, P1_U2753);
  not ginst1408 (P1_R2144_U87, P1_U2755);
  not ginst1409 (P1_R2144_U88, P1_U2756);
  not ginst1410 (P1_R2144_U89, P1_U2757);
  and ginst1411 (P1_R2144_U9, P1_R2144_U127, P1_R2144_U128);
  not ginst1412 (P1_R2144_U90, P1_U2758);
  nand ginst1413 (P1_R2144_U91, P1_R2144_U100, P1_R2144_U132);
  and ginst1414 (P1_R2144_U92, P1_R2144_U240, P1_R2144_U241);
  nand ginst1415 (P1_R2144_U93, P1_R2144_U113, P1_R2144_U129);
  nand ginst1416 (P1_R2144_U94, P1_R2144_U143, P1_R2144_U32);
  nand ginst1417 (P1_R2144_U95, P1_R2144_U141, P1_R2144_U34);
  nand ginst1418 (P1_R2144_U96, P1_R2144_U66, P1_R2144_U79);
  nand ginst1419 (P1_R2144_U97, P1_R2144_U67, P1_R2144_U79);
  nand ginst1420 (P1_R2144_U98, P1_R2144_U112, P1_R2144_U113);
  nand ginst1421 (P1_R2144_U99, P1_R2144_U53, P1_R2144_U84);
  not ginst1422 (P1_R2167_U10, P1_U2713);
  not ginst1423 (P1_R2167_U11, P1_U2712);
  not ginst1424 (P1_R2167_U12, P1_U2718);
  not ginst1425 (P1_R2167_U13, P1_U2717);
  not ginst1426 (P1_R2167_U14, P1_U2711);
  not ginst1427 (P1_R2167_U15, P1_U2356);
  not ginst1428 (P1_R2167_U16, P1_STATE2_REG_0__SCAN_IN);
  nand ginst1429 (P1_R2167_U17, P1_R2167_U49, P1_R2167_U50);
  and ginst1430 (P1_R2167_U18, P1_R2167_U29, P1_R2167_U30);
  and ginst1431 (P1_R2167_U19, P1_R2167_U32, P1_R2167_U33);
  and ginst1432 (P1_R2167_U20, P1_R2167_U35, P1_R2167_U36);
  and ginst1433 (P1_R2167_U21, P1_R2167_U38, P1_R2167_U39);
  not ginst1434 (P1_R2167_U22, P1_U2721);
  not ginst1435 (P1_R2167_U23, P1_U2722);
  nand ginst1436 (P1_R2167_U24, P1_R2167_U23, P1_U2715);
  nand ginst1437 (P1_R2167_U25, P1_R2167_U22, P1_U2715);
  or ginst1438 (P1_R2167_U26, P1_U2721, P1_U2722);
  nand ginst1439 (P1_R2167_U27, P1_R2167_U8, P1_U2714);
  nand ginst1440 (P1_R2167_U28, P1_R2167_U24, P1_R2167_U25, P1_R2167_U26, P1_R2167_U27);
  nand ginst1441 (P1_R2167_U29, P1_R2167_U7, P1_U2720);
  nand ginst1442 (P1_R2167_U30, P1_R2167_U10, P1_U2719);
  nand ginst1443 (P1_R2167_U31, P1_R2167_U18, P1_R2167_U28);
  nand ginst1444 (P1_R2167_U32, P1_R2167_U9, P1_U2713);
  nand ginst1445 (P1_R2167_U33, P1_R2167_U12, P1_U2712);
  nand ginst1446 (P1_R2167_U34, P1_R2167_U19, P1_R2167_U31);
  nand ginst1447 (P1_R2167_U35, P1_R2167_U11, P1_U2718);
  nand ginst1448 (P1_R2167_U36, P1_R2167_U14, P1_U2717);
  nand ginst1449 (P1_R2167_U37, P1_R2167_U20, P1_R2167_U34);
  nand ginst1450 (P1_R2167_U38, P1_R2167_U13, P1_U2711);
  nand ginst1451 (P1_R2167_U39, P1_R2167_U6, P1_U2356);
  nand ginst1452 (P1_R2167_U40, P1_R2167_U21, P1_R2167_U37);
  nand ginst1453 (P1_R2167_U41, P1_R2167_U15, P1_U2716);
  nand ginst1454 (P1_R2167_U42, P1_R2167_U40, P1_R2167_U41);
  nand ginst1455 (P1_R2167_U43, P1_R2167_U16, P1_U2716);
  nand ginst1456 (P1_R2167_U44, P1_R2167_U42, P1_R2167_U6);
  nand ginst1457 (P1_R2167_U45, P1_R2167_U43, P1_R2167_U44);
  nand ginst1458 (P1_R2167_U46, P1_STATE2_REG_0__SCAN_IN, P1_R2167_U6);
  nand ginst1459 (P1_R2167_U47, P1_R2167_U42, P1_U2716);
  nand ginst1460 (P1_R2167_U48, P1_R2167_U46, P1_R2167_U47);
  nand ginst1461 (P1_R2167_U49, P1_R2167_U15, P1_R2167_U45);
  nand ginst1462 (P1_R2167_U50, P1_R2167_U48, P1_U2356);
  not ginst1463 (P1_R2167_U6, P1_U2716);
  not ginst1464 (P1_R2167_U7, P1_U2714);
  not ginst1465 (P1_R2167_U8, P1_U2720);
  not ginst1466 (P1_R2167_U9, P1_U2719);
  not ginst1467 (P1_R2182_U10, P1_U2742);
  not ginst1468 (P1_R2182_U11, P1_U2741);
  not ginst1469 (P1_R2182_U12, P1_U2740);
  nand ginst1470 (P1_R2182_U13, P1_R2182_U35, P1_R2182_U41);
  not ginst1471 (P1_R2182_U14, P1_U2737);
  not ginst1472 (P1_R2182_U15, P1_U2738);
  nand ginst1473 (P1_R2182_U16, P1_U2723, P1_U2739);
  not ginst1474 (P1_R2182_U17, P1_U2736);
  not ginst1475 (P1_R2182_U18, P1_U2735);
  nand ginst1476 (P1_R2182_U19, P1_R2182_U36, P1_R2182_U49);
  not ginst1477 (P1_R2182_U20, P1_U2734);
  nand ginst1478 (P1_R2182_U21, P1_R2182_U37, P1_R2182_U46);
  nand ginst1479 (P1_R2182_U22, P1_R2182_U48, P1_U2734);
  not ginst1480 (P1_R2182_U23, P1_U2733);
  nand ginst1481 (P1_R2182_U24, P1_R2182_U63, P1_R2182_U64);
  nand ginst1482 (P1_R2182_U25, P1_R2182_U65, P1_R2182_U66);
  nand ginst1483 (P1_R2182_U26, P1_R2182_U67, P1_R2182_U68);
  nand ginst1484 (P1_R2182_U27, P1_R2182_U71, P1_R2182_U72);
  nand ginst1485 (P1_R2182_U28, P1_R2182_U73, P1_R2182_U74);
  nand ginst1486 (P1_R2182_U29, P1_R2182_U75, P1_R2182_U76);
  nand ginst1487 (P1_R2182_U30, P1_R2182_U77, P1_R2182_U78);
  nand ginst1488 (P1_R2182_U31, P1_R2182_U79, P1_R2182_U80);
  nand ginst1489 (P1_R2182_U32, P1_R2182_U81, P1_R2182_U82);
  nand ginst1490 (P1_R2182_U33, P1_R2182_U83, P1_R2182_U84);
  nand ginst1491 (P1_R2182_U34, P1_R2182_U85, P1_R2182_U86);
  and ginst1492 (P1_R2182_U35, P1_U2741, P1_U2742);
  and ginst1493 (P1_R2182_U36, P1_U2737, P1_U2738);
  and ginst1494 (P1_R2182_U37, P1_U2735, P1_U2736);
  nand ginst1495 (P1_R2182_U38, P1_R2182_U41, P1_U2742);
  not ginst1496 (P1_R2182_U39, P1_U2732);
  nand ginst1497 (P1_R2182_U40, P1_R2182_U56, P1_U2733);
  nand ginst1498 (P1_R2182_U41, P1_R2182_U52, P1_R2182_U53);
  and ginst1499 (P1_R2182_U42, P1_R2182_U69, P1_R2182_U70);
  nand ginst1500 (P1_R2182_U43, P1_R2182_U46, P1_U2736);
  nand ginst1501 (P1_R2182_U44, P1_R2182_U49, P1_U2738);
  nand ginst1502 (P1_R2182_U45, P1_R2182_U51, P1_R2182_U62);
  not ginst1503 (P1_R2182_U46, P1_R2182_U19);
  not ginst1504 (P1_R2182_U47, P1_R2182_U13);
  not ginst1505 (P1_R2182_U48, P1_R2182_U21);
  not ginst1506 (P1_R2182_U49, P1_R2182_U16);
  and ginst1507 (P1_R2182_U5, P1_R2182_U47, P1_U2740);
  not ginst1508 (P1_R2182_U50, P1_R2182_U9);
  or ginst1509 (P1_R2182_U51, P1_U2731, P1_U2743);
  nand ginst1510 (P1_R2182_U52, P1_U2731, P1_U2743);
  nand ginst1511 (P1_R2182_U53, P1_R2182_U50, P1_R2182_U51);
  not ginst1512 (P1_R2182_U54, P1_R2182_U41);
  not ginst1513 (P1_R2182_U55, P1_R2182_U38);
  not ginst1514 (P1_R2182_U56, P1_R2182_U22);
  not ginst1515 (P1_R2182_U57, P1_R2182_U40);
  not ginst1516 (P1_R2182_U58, P1_R2182_U43);
  not ginst1517 (P1_R2182_U59, P1_R2182_U44);
  and ginst1518 (P1_R2182_U6, P1_R2182_U16, P1_R2182_U60);
  or ginst1519 (P1_R2182_U60, P1_U2723, P1_U2739);
  not ginst1520 (P1_R2182_U61, P1_R2182_U45);
  nand ginst1521 (P1_R2182_U62, P1_U2731, P1_U2743);
  nand ginst1522 (P1_R2182_U63, P1_R2182_U12, P1_R2182_U47);
  nand ginst1523 (P1_R2182_U64, P1_R2182_U13, P1_U2740);
  nand ginst1524 (P1_R2182_U65, P1_R2182_U38, P1_U2741);
  nand ginst1525 (P1_R2182_U66, P1_R2182_U11, P1_R2182_U55);
  nand ginst1526 (P1_R2182_U67, P1_R2182_U40, P1_U2732);
  nand ginst1527 (P1_R2182_U68, P1_R2182_U39, P1_R2182_U57);
  nand ginst1528 (P1_R2182_U69, P1_R2182_U41, P1_U2742);
  not ginst1529 (P1_R2182_U7, P1_U2744);
  nand ginst1530 (P1_R2182_U70, P1_R2182_U10, P1_R2182_U54);
  nand ginst1531 (P1_R2182_U71, P1_R2182_U22, P1_U2733);
  nand ginst1532 (P1_R2182_U72, P1_R2182_U23, P1_R2182_U56);
  nand ginst1533 (P1_R2182_U73, P1_R2182_U20, P1_R2182_U48);
  nand ginst1534 (P1_R2182_U74, P1_R2182_U21, P1_U2734);
  nand ginst1535 (P1_R2182_U75, P1_R2182_U43, P1_U2735);
  nand ginst1536 (P1_R2182_U76, P1_R2182_U18, P1_R2182_U58);
  nand ginst1537 (P1_R2182_U77, P1_R2182_U17, P1_R2182_U46);
  nand ginst1538 (P1_R2182_U78, P1_R2182_U19, P1_U2736);
  nand ginst1539 (P1_R2182_U79, P1_R2182_U44, P1_U2737);
  not ginst1540 (P1_R2182_U8, P1_U3246);
  nand ginst1541 (P1_R2182_U80, P1_R2182_U14, P1_R2182_U59);
  nand ginst1542 (P1_R2182_U81, P1_R2182_U15, P1_R2182_U49);
  nand ginst1543 (P1_R2182_U82, P1_R2182_U16, P1_U2738);
  nand ginst1544 (P1_R2182_U83, P1_R2182_U45, P1_R2182_U50);
  nand ginst1545 (P1_R2182_U84, P1_R2182_U61, P1_R2182_U9);
  nand ginst1546 (P1_R2182_U85, P1_R2182_U7, P1_U3246);
  nand ginst1547 (P1_R2182_U86, P1_R2182_U8, P1_U2744);
  nand ginst1548 (P1_R2182_U9, P1_U2744, P1_U3246);
  not ginst1549 (P1_R2238_U10, P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN);
  not ginst1550 (P1_R2238_U11, P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN);
  not ginst1551 (P1_R2238_U12, P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN);
  not ginst1552 (P1_R2238_U13, P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN);
  not ginst1553 (P1_R2238_U14, P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN);
  not ginst1554 (P1_R2238_U15, P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN);
  nand ginst1555 (P1_R2238_U16, P1_R2238_U40, P1_R2238_U41);
  not ginst1556 (P1_R2238_U17, P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN);
  not ginst1557 (P1_R2238_U18, P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN);
  nand ginst1558 (P1_R2238_U19, P1_R2238_U50, P1_R2238_U51);
  nand ginst1559 (P1_R2238_U20, P1_R2238_U55, P1_R2238_U56);
  nand ginst1560 (P1_R2238_U21, P1_R2238_U60, P1_R2238_U61);
  nand ginst1561 (P1_R2238_U22, P1_R2238_U65, P1_R2238_U66);
  nand ginst1562 (P1_R2238_U23, P1_R2238_U47, P1_R2238_U48);
  nand ginst1563 (P1_R2238_U24, P1_R2238_U52, P1_R2238_U53);
  nand ginst1564 (P1_R2238_U25, P1_R2238_U57, P1_R2238_U58);
  nand ginst1565 (P1_R2238_U26, P1_R2238_U62, P1_R2238_U63);
  nand ginst1566 (P1_R2238_U27, P1_R2238_U36, P1_R2238_U37);
  nand ginst1567 (P1_R2238_U28, P1_R2238_U32, P1_R2238_U33);
  not ginst1568 (P1_R2238_U29, P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN);
  not ginst1569 (P1_R2238_U30, P1_R2238_U9);
  nand ginst1570 (P1_R2238_U31, P1_R2238_U10, P1_R2238_U30);
  nand ginst1571 (P1_R2238_U32, P1_R2238_U29, P1_R2238_U31);
  nand ginst1572 (P1_R2238_U33, P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN, P1_R2238_U9);
  not ginst1573 (P1_R2238_U34, P1_R2238_U28);
  nand ginst1574 (P1_R2238_U35, P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN, P1_R2238_U12);
  nand ginst1575 (P1_R2238_U36, P1_R2238_U28, P1_R2238_U35);
  nand ginst1576 (P1_R2238_U37, P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN, P1_R2238_U11);
  not ginst1577 (P1_R2238_U38, P1_R2238_U27);
  nand ginst1578 (P1_R2238_U39, P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P1_R2238_U14);
  nand ginst1579 (P1_R2238_U40, P1_R2238_U27, P1_R2238_U39);
  nand ginst1580 (P1_R2238_U41, P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN, P1_R2238_U13);
  not ginst1581 (P1_R2238_U42, P1_R2238_U16);
  nand ginst1582 (P1_R2238_U43, P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN, P1_R2238_U17);
  nand ginst1583 (P1_R2238_U44, P1_R2238_U42, P1_R2238_U43);
  nand ginst1584 (P1_R2238_U45, P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN, P1_R2238_U15);
  nand ginst1585 (P1_R2238_U46, P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P1_R2238_U8);
  nand ginst1586 (P1_R2238_U47, P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN, P1_R2238_U15);
  nand ginst1587 (P1_R2238_U48, P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN, P1_R2238_U17);
  not ginst1588 (P1_R2238_U49, P1_R2238_U23);
  nand ginst1589 (P1_R2238_U50, P1_R2238_U42, P1_R2238_U49);
  nand ginst1590 (P1_R2238_U51, P1_R2238_U16, P1_R2238_U23);
  nand ginst1591 (P1_R2238_U52, P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P1_R2238_U14);
  nand ginst1592 (P1_R2238_U53, P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN, P1_R2238_U13);
  not ginst1593 (P1_R2238_U54, P1_R2238_U24);
  nand ginst1594 (P1_R2238_U55, P1_R2238_U38, P1_R2238_U54);
  nand ginst1595 (P1_R2238_U56, P1_R2238_U24, P1_R2238_U27);
  nand ginst1596 (P1_R2238_U57, P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN, P1_R2238_U12);
  nand ginst1597 (P1_R2238_U58, P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN, P1_R2238_U11);
  not ginst1598 (P1_R2238_U59, P1_R2238_U25);
  nand ginst1599 (P1_R2238_U6, P1_R2238_U44, P1_R2238_U45);
  nand ginst1600 (P1_R2238_U60, P1_R2238_U34, P1_R2238_U59);
  nand ginst1601 (P1_R2238_U61, P1_R2238_U25, P1_R2238_U28);
  nand ginst1602 (P1_R2238_U62, P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P1_R2238_U10);
  nand ginst1603 (P1_R2238_U63, P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN, P1_R2238_U29);
  not ginst1604 (P1_R2238_U64, P1_R2238_U26);
  nand ginst1605 (P1_R2238_U65, P1_R2238_U30, P1_R2238_U64);
  nand ginst1606 (P1_R2238_U66, P1_R2238_U26, P1_R2238_U9);
  nand ginst1607 (P1_R2238_U7, P1_R2238_U46, P1_R2238_U9);
  not ginst1608 (P1_R2238_U8, P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN);
  nand ginst1609 (P1_R2238_U9, P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN, P1_R2238_U18);
  and ginst1610 (P1_R2278_U10, P1_R2278_U311, P1_R2278_U313, P1_R2278_U315);
  and ginst1611 (P1_R2278_U100, P1_R2278_U261, P1_R2278_U262);
  nand ginst1612 (P1_R2278_U101, P1_R2278_U430, P1_R2278_U431);
  nand ginst1613 (P1_R2278_U102, P1_R2278_U437, P1_R2278_U438);
  nand ginst1614 (P1_R2278_U103, P1_R2278_U444, P1_R2278_U445);
  nand ginst1615 (P1_R2278_U104, P1_R2278_U453, P1_R2278_U454);
  nand ginst1616 (P1_R2278_U105, P1_R2278_U460, P1_R2278_U461);
  nand ginst1617 (P1_R2278_U106, P1_R2278_U476, P1_R2278_U477);
  nand ginst1618 (P1_R2278_U107, P1_R2278_U483, P1_R2278_U484);
  nand ginst1619 (P1_R2278_U108, P1_R2278_U490, P1_R2278_U491);
  nand ginst1620 (P1_R2278_U109, P1_R2278_U497, P1_R2278_U498);
  and ginst1621 (P1_R2278_U11, P1_R2278_U10, P1_R2278_U134);
  nand ginst1622 (P1_R2278_U110, P1_R2278_U504, P1_R2278_U505);
  nand ginst1623 (P1_R2278_U111, P1_R2278_U511, P1_R2278_U512);
  nand ginst1624 (P1_R2278_U112, P1_R2278_U518, P1_R2278_U519);
  nand ginst1625 (P1_R2278_U113, P1_R2278_U525, P1_R2278_U526);
  nand ginst1626 (P1_R2278_U114, P1_R2278_U532, P1_R2278_U533);
  nand ginst1627 (P1_R2278_U115, P1_R2278_U539, P1_R2278_U540);
  nand ginst1628 (P1_R2278_U116, P1_R2278_U546, P1_R2278_U547);
  nand ginst1629 (P1_R2278_U117, P1_R2278_U553, P1_R2278_U554);
  nand ginst1630 (P1_R2278_U118, P1_R2278_U565, P1_R2278_U566);
  nand ginst1631 (P1_R2278_U119, P1_R2278_U572, P1_R2278_U573);
  and ginst1632 (P1_R2278_U12, P1_R2278_U292, P1_R2278_U295);
  nand ginst1633 (P1_R2278_U120, P1_R2278_U579, P1_R2278_U580);
  nand ginst1634 (P1_R2278_U121, P1_R2278_U586, P1_R2278_U587);
  nand ginst1635 (P1_R2278_U122, P1_R2278_U593, P1_R2278_U594);
  nand ginst1636 (P1_R2278_U123, P1_R2278_U598, P1_R2278_U599);
  and ginst1637 (P1_R2278_U124, P1_R2278_U281, P1_R2278_U68);
  nand ginst1638 (P1_R2278_U125, P1_R2278_U600, P1_R2278_U601);
  nand ginst1639 (P1_R2278_U126, P1_R2278_U607, P1_R2278_U608);
  and ginst1640 (P1_R2278_U127, P1_INSTADDRPOINTER_REG_7__SCAN_IN, P1_U2793);
  and ginst1641 (P1_R2278_U128, P1_R2278_U254, P1_R2278_U258);
  and ginst1642 (P1_R2278_U129, P1_R2278_U259, P1_R2278_U352);
  and ginst1643 (P1_R2278_U13, P1_R2278_U321, P1_R2278_U9);
  and ginst1644 (P1_R2278_U130, P1_INSTADDRPOINTER_REG_23__SCAN_IN, P1_U2777);
  and ginst1645 (P1_R2278_U131, P1_R2278_U316, P1_R2278_U318);
  and ginst1646 (P1_R2278_U132, P1_R2278_U317, P1_R2278_U319, P1_R2278_U321);
  and ginst1647 (P1_R2278_U133, P1_INSTADDRPOINTER_REG_19__SCAN_IN, P1_U2781);
  and ginst1648 (P1_R2278_U134, P1_R2278_U317, P1_R2278_U319);
  and ginst1649 (P1_R2278_U135, P1_R2278_U308, P1_R2278_U321);
  and ginst1650 (P1_R2278_U136, P1_R2278_U11, P1_R2278_U135);
  and ginst1651 (P1_R2278_U137, P1_R2278_U228, P1_R2278_U259, P1_R2278_U273);
  and ginst1652 (P1_R2278_U138, P1_R2278_U276, P1_R2278_U389);
  and ginst1653 (P1_R2278_U139, P1_R2278_U140, P1_R2278_U357);
  and ginst1654 (P1_R2278_U14, P1_R2278_U462, P1_R2278_U463);
  and ginst1655 (P1_R2278_U140, P1_R2278_U281, P1_R2278_U283, P1_R2278_U284);
  and ginst1656 (P1_R2278_U141, P1_R2278_U286, P1_R2278_U410);
  and ginst1657 (P1_R2278_U142, P1_R2278_U13, P1_R2278_U7);
  and ginst1658 (P1_R2278_U143, P1_R2278_U309, P1_R2278_U321);
  and ginst1659 (P1_R2278_U144, P1_R2278_U296, P1_R2278_U308);
  and ginst1660 (P1_R2278_U145, P1_R2278_U94, P1_R2278_U95);
  and ginst1661 (P1_R2278_U146, P1_R2278_U401, P1_R2278_U96);
  and ginst1662 (P1_R2278_U147, P1_R2278_U324, P1_R2278_U5);
  and ginst1663 (P1_R2278_U148, P1_R2278_U317, P1_R2278_U319, P1_R2278_U321, P1_R2278_U324);
  and ginst1664 (P1_R2278_U149, P1_R2278_U308, P1_R2278_U321, P1_R2278_U324);
  and ginst1665 (P1_R2278_U15, P1_R2278_U342, P1_R2278_U344);
  and ginst1666 (P1_R2278_U150, P1_R2278_U11, P1_R2278_U149);
  and ginst1667 (P1_R2278_U151, P1_R2278_U286, P1_R2278_U412);
  and ginst1668 (P1_R2278_U152, P1_R2278_U11, P1_R2278_U324);
  and ginst1669 (P1_R2278_U153, P1_R2278_U13, P1_R2278_U7);
  and ginst1670 (P1_R2278_U154, P1_R2278_U321, P1_R2278_U324);
  and ginst1671 (P1_R2278_U155, P1_R2278_U156, P1_R2278_U393, P1_R2278_U394, P1_R2278_U395, P1_R2278_U398);
  and ginst1672 (P1_R2278_U156, P1_R2278_U14, P1_R2278_U399, P1_R2278_U400);
  and ginst1673 (P1_R2278_U157, P1_R2278_U11, P1_R2278_U324);
  and ginst1674 (P1_R2278_U158, P1_R2278_U13, P1_R2278_U7);
  and ginst1675 (P1_R2278_U159, P1_R2278_U187, P1_R2278_U403, P1_R2278_U404);
  and ginst1676 (P1_R2278_U16, P1_R2278_U188, P1_R2278_U375, P1_R2278_U467, P1_R2278_U468);
  and ginst1677 (P1_R2278_U160, P1_R2278_U286, P1_R2278_U417);
  and ginst1678 (P1_R2278_U161, P1_R2278_U7, P1_R2278_U9);
  and ginst1679 (P1_R2278_U162, P1_R2278_U369, P1_R2278_U76);
  and ginst1680 (P1_R2278_U163, P1_R2278_U73, P1_R2278_U80);
  and ginst1681 (P1_R2278_U164, P1_R2278_U10, P1_R2278_U317);
  and ginst1682 (P1_R2278_U165, P1_R2278_U316, P1_R2278_U371);
  and ginst1683 (P1_R2278_U166, P1_R2278_U311, P1_R2278_U313);
  and ginst1684 (P1_R2278_U167, P1_R2278_U314, P1_R2278_U370);
  and ginst1685 (P1_R2278_U168, P1_R2278_U286, P1_R2278_U415);
  and ginst1686 (P1_R2278_U169, P1_R2278_U362, P1_R2278_U79);
  and ginst1687 (P1_R2278_U17, P1_R2278_U270, P1_R2278_U272);
  and ginst1688 (P1_R2278_U170, P1_R2278_U306, P1_R2278_U367);
  and ginst1689 (P1_R2278_U171, P1_R2278_U298, P1_R2278_U302);
  and ginst1690 (P1_R2278_U172, P1_R2278_U303, P1_R2278_U364);
  and ginst1691 (P1_R2278_U173, P1_R2278_U285, P1_R2278_U588, P1_R2278_U589);
  and ginst1692 (P1_R2278_U174, P1_R2278_U227, P1_R2278_U337);
  and ginst1693 (P1_R2278_U175, P1_R2278_U228, P1_R2278_U602, P1_R2278_U603);
  nand ginst1694 (P1_R2278_U176, P1_R2278_U129, P1_R2278_U353);
  and ginst1695 (P1_R2278_U177, P1_R2278_U432, P1_R2278_U433);
  nand ginst1696 (P1_R2278_U178, P1_R2278_U256, P1_R2278_U41);
  and ginst1697 (P1_R2278_U179, P1_R2278_U439, P1_R2278_U440);
  and ginst1698 (P1_R2278_U18, P1_R2278_U266, P1_R2278_U268);
  and ginst1699 (P1_R2278_U180, P1_R2278_U446, P1_R2278_U447);
  and ginst1700 (P1_R2278_U181, P1_R2278_U448, P1_R2278_U449);
  nand ginst1701 (P1_R2278_U182, P1_R2278_U241, P1_R2278_U242);
  and ginst1702 (P1_R2278_U183, P1_R2278_U455, P1_R2278_U456);
  nand ginst1703 (P1_R2278_U184, P1_R2278_U237, P1_R2278_U238);
  not ginst1704 (P1_R2278_U185, P1_INSTADDRPOINTER_REG_31__SCAN_IN);
  not ginst1705 (P1_R2278_U186, P1_U2769);
  nand ginst1706 (P1_R2278_U187, P1_INSTADDRPOINTER_REG_29__SCAN_IN, P1_U2771);
  and ginst1707 (P1_R2278_U188, P1_R2278_U469, P1_R2278_U470);
  and ginst1708 (P1_R2278_U189, P1_R2278_U471, P1_R2278_U472);
  nand ginst1709 (P1_R2278_U19, P1_R2278_U214, P1_R2278_U429);
  nand ginst1710 (P1_R2278_U190, P1_R2278_U159, P1_R2278_U405, P1_R2278_U406, P1_R2278_U407);
  and ginst1711 (P1_R2278_U191, P1_R2278_U478, P1_R2278_U479);
  nand ginst1712 (P1_R2278_U192, P1_R2278_U213, P1_R2278_U234);
  and ginst1713 (P1_R2278_U193, P1_R2278_U485, P1_R2278_U486);
  nand ginst1714 (P1_R2278_U194, P1_R2278_U145, P1_R2278_U146, P1_R2278_U385);
  and ginst1715 (P1_R2278_U195, P1_R2278_U492, P1_R2278_U493);
  nand ginst1716 (P1_R2278_U196, P1_R2278_U409, P1_R2278_U419);
  and ginst1717 (P1_R2278_U197, P1_R2278_U499, P1_R2278_U500);
  nand ginst1718 (P1_R2278_U198, P1_R2278_U373, P1_R2278_U425);
  and ginst1719 (P1_R2278_U199, P1_R2278_U506, P1_R2278_U507);
  and ginst1720 (P1_R2278_U20, P1_R2278_U335, P1_R2278_U414);
  nand ginst1721 (P1_R2278_U200, P1_R2278_U165, P1_R2278_U423);
  and ginst1722 (P1_R2278_U201, P1_R2278_U513, P1_R2278_U514);
  nand ginst1723 (P1_R2278_U202, P1_R2278_U167, P1_R2278_U427);
  and ginst1724 (P1_R2278_U203, P1_R2278_U520, P1_R2278_U521);
  nand ginst1725 (P1_R2278_U204, P1_R2278_U312, P1_R2278_U421);
  and ginst1726 (P1_R2278_U205, P1_R2278_U527, P1_R2278_U528);
  nand ginst1727 (P1_R2278_U206, P1_R2278_U162, P1_R2278_U163, P1_R2278_U376);
  and ginst1728 (P1_R2278_U207, P1_R2278_U534, P1_R2278_U535);
  nand ginst1729 (P1_R2278_U208, P1_R2278_U170, P1_R2278_U365);
  and ginst1730 (P1_R2278_U209, P1_R2278_U541, P1_R2278_U542);
  not ginst1731 (P1_R2278_U21, P1_INSTADDRPOINTER_REG_8__SCAN_IN);
  nand ginst1732 (P1_R2278_U210, P1_R2278_U172, P1_R2278_U363);
  and ginst1733 (P1_R2278_U211, P1_R2278_U548, P1_R2278_U549);
  nand ginst1734 (P1_R2278_U212, P1_R2278_U299, P1_R2278_U300);
  nand ginst1735 (P1_R2278_U213, P1_R2278_U232, P1_U2799);
  and ginst1736 (P1_R2278_U214, P1_R2278_U558, P1_R2278_U559);
  and ginst1737 (P1_R2278_U215, P1_R2278_U560, P1_R2278_U561);
  nand ginst1738 (P1_R2278_U216, P1_R2278_U169, P1_R2278_U361);
  and ginst1739 (P1_R2278_U217, P1_R2278_U567, P1_R2278_U568);
  nand ginst1740 (P1_R2278_U218, P1_R2278_U358, P1_R2278_U360);
  and ginst1741 (P1_R2278_U219, P1_R2278_U574, P1_R2278_U575);
  not ginst1742 (P1_R2278_U22, P1_U2792);
  nand ginst1743 (P1_R2278_U220, P1_R2278_U289, P1_R2278_U290);
  and ginst1744 (P1_R2278_U221, P1_R2278_U581, P1_R2278_U582);
  nand ginst1745 (P1_R2278_U222, P1_R2278_U168, P1_R2278_U226);
  nand ginst1746 (P1_R2278_U223, P1_R2278_U328, P1_R2278_U68);
  nand ginst1747 (P1_R2278_U224, P1_R2278_U279, P1_R2278_U98);
  nand ginst1748 (P1_R2278_U225, P1_R2278_U273, P1_R2278_U274);
  nand ginst1749 (P1_R2278_U226, P1_R2278_U139, P1_R2278_U224);
  nand ginst1750 (P1_R2278_U227, P1_R2278_U355, P1_R2278_U356);
  nand ginst1751 (P1_R2278_U228, P1_INSTADDRPOINTER_REG_10__SCAN_IN, P1_U2790);
  nand ginst1752 (P1_R2278_U229, P1_INSTADDRPOINTER_REG_13__SCAN_IN, P1_U2787);
  not ginst1753 (P1_R2278_U23, P1_INSTADDRPOINTER_REG_7__SCAN_IN);
  not ginst1754 (P1_R2278_U230, P1_R2278_U213);
  nand ginst1755 (P1_R2278_U231, P1_INSTADDRPOINTER_REG_6__SCAN_IN, P1_U2794);
  not ginst1756 (P1_R2278_U232, P1_R2278_U32);
  nand ginst1757 (P1_R2278_U233, P1_R2278_U32, P1_R2278_U33);
  nand ginst1758 (P1_R2278_U234, P1_INSTADDRPOINTER_REG_1__SCAN_IN, P1_R2278_U233);
  not ginst1759 (P1_R2278_U235, P1_R2278_U192);
  or ginst1760 (P1_R2278_U236, P1_INSTADDRPOINTER_REG_2__SCAN_IN, P1_U2798);
  nand ginst1761 (P1_R2278_U237, P1_R2278_U192, P1_R2278_U236);
  nand ginst1762 (P1_R2278_U238, P1_INSTADDRPOINTER_REG_2__SCAN_IN, P1_U2798);
  not ginst1763 (P1_R2278_U239, P1_R2278_U184);
  not ginst1764 (P1_R2278_U24, P1_U2793);
  or ginst1765 (P1_R2278_U240, P1_INSTADDRPOINTER_REG_3__SCAN_IN, P1_U2797);
  nand ginst1766 (P1_R2278_U241, P1_R2278_U184, P1_R2278_U240);
  nand ginst1767 (P1_R2278_U242, P1_INSTADDRPOINTER_REG_3__SCAN_IN, P1_U2797);
  not ginst1768 (P1_R2278_U243, P1_R2278_U182);
  or ginst1769 (P1_R2278_U244, P1_INSTADDRPOINTER_REG_4__SCAN_IN, P1_U2796);
  nand ginst1770 (P1_R2278_U245, P1_R2278_U182, P1_R2278_U244);
  nand ginst1771 (P1_R2278_U246, P1_INSTADDRPOINTER_REG_4__SCAN_IN, P1_U2796);
  not ginst1772 (P1_R2278_U247, P1_R2278_U42);
  or ginst1773 (P1_R2278_U248, P1_INSTADDRPOINTER_REG_5__SCAN_IN, P1_U2795);
  not ginst1774 (P1_R2278_U249, P1_R2278_U43);
  not ginst1775 (P1_R2278_U25, P1_INSTADDRPOINTER_REG_6__SCAN_IN);
  nand ginst1776 (P1_R2278_U250, P1_INSTADDRPOINTER_REG_5__SCAN_IN, P1_U2795);
  not ginst1777 (P1_R2278_U251, P1_R2278_U40);
  nand ginst1778 (P1_R2278_U252, P1_R2278_U231, P1_R2278_U251);
  or ginst1779 (P1_R2278_U253, P1_INSTADDRPOINTER_REG_7__SCAN_IN, P1_U2793);
  or ginst1780 (P1_R2278_U254, P1_INSTADDRPOINTER_REG_6__SCAN_IN, P1_U2794);
  not ginst1781 (P1_R2278_U255, P1_R2278_U41);
  nand ginst1782 (P1_R2278_U256, P1_INSTADDRPOINTER_REG_7__SCAN_IN, P1_U2793);
  not ginst1783 (P1_R2278_U257, P1_R2278_U178);
  or ginst1784 (P1_R2278_U258, P1_INSTADDRPOINTER_REG_8__SCAN_IN, P1_U2792);
  nand ginst1785 (P1_R2278_U259, P1_INSTADDRPOINTER_REG_8__SCAN_IN, P1_U2792);
  not ginst1786 (P1_R2278_U26, P1_U2794);
  not ginst1787 (P1_R2278_U260, P1_R2278_U176);
  or ginst1788 (P1_R2278_U261, P1_INSTADDRPOINTER_REG_9__SCAN_IN, P1_U2791);
  nand ginst1789 (P1_R2278_U262, P1_INSTADDRPOINTER_REG_9__SCAN_IN, P1_U2791);
  nand ginst1790 (P1_R2278_U263, P1_INSTADDRPOINTER_REG_9__SCAN_IN, P1_U2791);
  or ginst1791 (P1_R2278_U264, P1_INSTADDRPOINTER_REG_6__SCAN_IN, P1_U2794);
  nand ginst1792 (P1_R2278_U265, P1_R2278_U264, P1_R2278_U40);
  nand ginst1793 (P1_R2278_U266, P1_R2278_U179, P1_R2278_U231, P1_R2278_U265);
  nand ginst1794 (P1_R2278_U267, P1_INSTADDRPOINTER_REG_7__SCAN_IN, P1_U2793);
  nand ginst1795 (P1_R2278_U268, P1_R2278_U255, P1_R2278_U267);
  or ginst1796 (P1_R2278_U269, P1_INSTADDRPOINTER_REG_6__SCAN_IN, P1_U2794);
  not ginst1797 (P1_R2278_U27, P1_INSTADDRPOINTER_REG_5__SCAN_IN);
  nand ginst1798 (P1_R2278_U270, P1_R2278_U180, P1_R2278_U247);
  nand ginst1799 (P1_R2278_U271, P1_INSTADDRPOINTER_REG_5__SCAN_IN, P1_U2795);
  nand ginst1800 (P1_R2278_U272, P1_R2278_U249, P1_R2278_U271);
  nand ginst1801 (P1_R2278_U273, P1_INSTADDRPOINTER_REG_9__SCAN_IN, P1_U2791);
  nand ginst1802 (P1_R2278_U274, P1_R2278_U176, P1_R2278_U261);
  not ginst1803 (P1_R2278_U275, P1_R2278_U225);
  or ginst1804 (P1_R2278_U276, P1_INSTADDRPOINTER_REG_11__SCAN_IN, P1_U2789);
  or ginst1805 (P1_R2278_U277, P1_INSTADDRPOINTER_REG_10__SCAN_IN, P1_U2790);
  not ginst1806 (P1_R2278_U278, P1_R2278_U98);
  nand ginst1807 (P1_R2278_U279, P1_INSTADDRPOINTER_REG_11__SCAN_IN, P1_U2789);
  not ginst1808 (P1_R2278_U28, P1_U2795);
  not ginst1809 (P1_R2278_U280, P1_R2278_U224);
  or ginst1810 (P1_R2278_U281, P1_INSTADDRPOINTER_REG_12__SCAN_IN, P1_U2788);
  not ginst1811 (P1_R2278_U282, P1_R2278_U68);
  or ginst1812 (P1_R2278_U283, P1_INSTADDRPOINTER_REG_13__SCAN_IN, P1_U2787);
  or ginst1813 (P1_R2278_U284, P1_INSTADDRPOINTER_REG_14__SCAN_IN, P1_U2786);
  nand ginst1814 (P1_R2278_U285, P1_INSTADDRPOINTER_REG_14__SCAN_IN, P1_U2786);
  nand ginst1815 (P1_R2278_U286, P1_INSTADDRPOINTER_REG_15__SCAN_IN, P1_U2785);
  nand ginst1816 (P1_R2278_U287, P1_R2278_U229, P1_R2278_U285, P1_R2278_U391);
  or ginst1817 (P1_R2278_U288, P1_INSTADDRPOINTER_REG_16__SCAN_IN, P1_U2784);
  nand ginst1818 (P1_R2278_U289, P1_R2278_U222, P1_R2278_U288);
  not ginst1819 (P1_R2278_U29, P1_U2800);
  nand ginst1820 (P1_R2278_U290, P1_INSTADDRPOINTER_REG_16__SCAN_IN, P1_U2784);
  not ginst1821 (P1_R2278_U291, P1_R2278_U220);
  or ginst1822 (P1_R2278_U292, P1_INSTADDRPOINTER_REG_17__SCAN_IN, P1_U2783);
  nand ginst1823 (P1_R2278_U293, P1_INSTADDRPOINTER_REG_17__SCAN_IN, P1_U2783);
  not ginst1824 (P1_R2278_U294, P1_R2278_U218);
  or ginst1825 (P1_R2278_U295, P1_INSTADDRPOINTER_REG_18__SCAN_IN, P1_U2782);
  not ginst1826 (P1_R2278_U296, P1_R2278_U79);
  not ginst1827 (P1_R2278_U297, P1_R2278_U216);
  or ginst1828 (P1_R2278_U298, P1_INSTADDRPOINTER_REG_19__SCAN_IN, P1_U2781);
  nand ginst1829 (P1_R2278_U299, P1_R2278_U216, P1_R2278_U298);
  not ginst1830 (P1_R2278_U30, P1_INSTADDRPOINTER_REG_0__SCAN_IN);
  nand ginst1831 (P1_R2278_U300, P1_INSTADDRPOINTER_REG_19__SCAN_IN, P1_U2781);
  not ginst1832 (P1_R2278_U301, P1_R2278_U212);
  or ginst1833 (P1_R2278_U302, P1_INSTADDRPOINTER_REG_20__SCAN_IN, P1_U2780);
  nand ginst1834 (P1_R2278_U303, P1_INSTADDRPOINTER_REG_20__SCAN_IN, P1_U2780);
  not ginst1835 (P1_R2278_U304, P1_R2278_U210);
  or ginst1836 (P1_R2278_U305, P1_INSTADDRPOINTER_REG_21__SCAN_IN, P1_U2779);
  nand ginst1837 (P1_R2278_U306, P1_INSTADDRPOINTER_REG_21__SCAN_IN, P1_U2779);
  not ginst1838 (P1_R2278_U307, P1_R2278_U208);
  or ginst1839 (P1_R2278_U308, P1_INSTADDRPOINTER_REG_22__SCAN_IN, P1_U2778);
  not ginst1840 (P1_R2278_U309, P1_R2278_U76);
  not ginst1841 (P1_R2278_U31, P1_INSTADDRPOINTER_REG_1__SCAN_IN);
  not ginst1842 (P1_R2278_U310, P1_R2278_U206);
  or ginst1843 (P1_R2278_U311, P1_INSTADDRPOINTER_REG_23__SCAN_IN, P1_U2777);
  nand ginst1844 (P1_R2278_U312, P1_INSTADDRPOINTER_REG_23__SCAN_IN, P1_U2777);
  or ginst1845 (P1_R2278_U313, P1_INSTADDRPOINTER_REG_24__SCAN_IN, P1_U2776);
  nand ginst1846 (P1_R2278_U314, P1_INSTADDRPOINTER_REG_24__SCAN_IN, P1_U2776);
  or ginst1847 (P1_R2278_U315, P1_INSTADDRPOINTER_REG_25__SCAN_IN, P1_U2775);
  nand ginst1848 (P1_R2278_U316, P1_INSTADDRPOINTER_REG_25__SCAN_IN, P1_U2775);
  or ginst1849 (P1_R2278_U317, P1_INSTADDRPOINTER_REG_26__SCAN_IN, P1_U2774);
  nand ginst1850 (P1_R2278_U318, P1_INSTADDRPOINTER_REG_26__SCAN_IN, P1_U2774);
  or ginst1851 (P1_R2278_U319, P1_INSTADDRPOINTER_REG_27__SCAN_IN, P1_U2773);
  nand ginst1852 (P1_R2278_U32, P1_INSTADDRPOINTER_REG_0__SCAN_IN, P1_U2800);
  not ginst1853 (P1_R2278_U320, P1_R2278_U85);
  or ginst1854 (P1_R2278_U321, P1_INSTADDRPOINTER_REG_28__SCAN_IN, P1_U2772);
  nand ginst1855 (P1_R2278_U322, P1_INSTADDRPOINTER_REG_28__SCAN_IN, P1_U2772);
  not ginst1856 (P1_R2278_U323, P1_R2278_U194);
  or ginst1857 (P1_R2278_U324, P1_INSTADDRPOINTER_REG_29__SCAN_IN, P1_U2771);
  not ginst1858 (P1_R2278_U325, P1_R2278_U187);
  not ginst1859 (P1_R2278_U326, P1_R2278_U190);
  or ginst1860 (P1_R2278_U327, P1_INSTADDRPOINTER_REG_30__SCAN_IN, P1_U2770);
  nand ginst1861 (P1_R2278_U328, P1_R2278_U224, P1_R2278_U281);
  not ginst1862 (P1_R2278_U329, P1_R2278_U223);
  not ginst1863 (P1_R2278_U33, P1_U2799);
  or ginst1864 (P1_R2278_U330, P1_INSTADDRPOINTER_REG_13__SCAN_IN, P1_U2787);
  nand ginst1865 (P1_R2278_U331, P1_R2278_U223, P1_R2278_U330);
  not ginst1866 (P1_R2278_U332, P1_R2278_U97);
  or ginst1867 (P1_R2278_U333, P1_INSTADDRPOINTER_REG_14__SCAN_IN, P1_U2786);
  nand ginst1868 (P1_R2278_U334, P1_R2278_U333, P1_R2278_U97);
  nand ginst1869 (P1_R2278_U335, P1_R2278_U173, P1_R2278_U334);
  nand ginst1870 (P1_R2278_U336, P1_R2278_U285, P1_R2278_U332);
  nand ginst1871 (P1_R2278_U337, P1_INSTADDRPOINTER_REG_15__SCAN_IN, P1_U2785);
  or ginst1872 (P1_R2278_U338, P1_INSTADDRPOINTER_REG_14__SCAN_IN, P1_U2786);
  or ginst1873 (P1_R2278_U339, P1_INSTADDRPOINTER_REG_13__SCAN_IN, P1_U2787);
  not ginst1874 (P1_R2278_U34, P1_INSTADDRPOINTER_REG_2__SCAN_IN);
  or ginst1875 (P1_R2278_U340, P1_INSTADDRPOINTER_REG_10__SCAN_IN, P1_U2790);
  nand ginst1876 (P1_R2278_U341, P1_R2278_U225, P1_R2278_U340);
  nand ginst1877 (P1_R2278_U342, P1_R2278_U175, P1_R2278_U341);
  nand ginst1878 (P1_R2278_U343, P1_INSTADDRPOINTER_REG_11__SCAN_IN, P1_U2789);
  nand ginst1879 (P1_R2278_U344, P1_R2278_U278, P1_R2278_U343);
  or ginst1880 (P1_R2278_U345, P1_INSTADDRPOINTER_REG_10__SCAN_IN, P1_U2790);
  nand ginst1881 (P1_R2278_U346, P1_R2278_U261, P1_R2278_U263);
  nand ginst1882 (P1_R2278_U347, P1_R2278_U231, P1_R2278_U269);
  nand ginst1883 (P1_R2278_U348, P1_R2278_U285, P1_R2278_U338);
  nand ginst1884 (P1_R2278_U349, P1_R2278_U229, P1_R2278_U339);
  not ginst1885 (P1_R2278_U35, P1_U2798);
  nand ginst1886 (P1_R2278_U350, P1_R2278_U281, P1_R2278_U68);
  nand ginst1887 (P1_R2278_U351, P1_R2278_U228, P1_R2278_U345);
  nand ginst1888 (P1_R2278_U352, P1_R2278_U127, P1_R2278_U258);
  nand ginst1889 (P1_R2278_U353, P1_R2278_U128, P1_R2278_U252, P1_R2278_U253);
  nand ginst1890 (P1_R2278_U354, P1_R2278_U137, P1_R2278_U352, P1_R2278_U353);
  nand ginst1891 (P1_R2278_U355, P1_R2278_U284, P1_U2785);
  nand ginst1892 (P1_R2278_U356, P1_INSTADDRPOINTER_REG_15__SCAN_IN, P1_R2278_U284);
  nand ginst1893 (P1_R2278_U357, P1_R2278_U356, P1_R2278_U63);
  nand ginst1894 (P1_R2278_U358, P1_R2278_U222, P1_R2278_U6);
  nand ginst1895 (P1_R2278_U359, P1_R2278_U290, P1_R2278_U293);
  not ginst1896 (P1_R2278_U36, P1_INSTADDRPOINTER_REG_3__SCAN_IN);
  nand ginst1897 (P1_R2278_U360, P1_R2278_U292, P1_R2278_U359);
  nand ginst1898 (P1_R2278_U361, P1_R2278_U222, P1_R2278_U7);
  nand ginst1899 (P1_R2278_U362, P1_R2278_U12, P1_R2278_U359);
  nand ginst1900 (P1_R2278_U363, P1_R2278_U171, P1_R2278_U216);
  nand ginst1901 (P1_R2278_U364, P1_R2278_U133, P1_R2278_U302);
  nand ginst1902 (P1_R2278_U365, P1_R2278_U216, P1_R2278_U8);
  nand ginst1903 (P1_R2278_U366, P1_R2278_U303, P1_R2278_U364);
  nand ginst1904 (P1_R2278_U367, P1_R2278_U305, P1_R2278_U366);
  nand ginst1905 (P1_R2278_U368, P1_R2278_U306, P1_R2278_U367);
  nand ginst1906 (P1_R2278_U369, P1_R2278_U308, P1_R2278_U368);
  not ginst1907 (P1_R2278_U37, P1_U2797);
  nand ginst1908 (P1_R2278_U370, P1_R2278_U130, P1_R2278_U313);
  nand ginst1909 (P1_R2278_U371, P1_R2278_U315, P1_R2278_U381);
  nand ginst1910 (P1_R2278_U372, P1_R2278_U131, P1_R2278_U371);
  nand ginst1911 (P1_R2278_U373, P1_R2278_U317, P1_R2278_U372);
  nand ginst1912 (P1_R2278_U374, P1_R2278_U317, P1_R2278_U372);
  nand ginst1913 (P1_R2278_U375, P1_R2278_U147, P1_R2278_U194);
  nand ginst1914 (P1_R2278_U376, P1_R2278_U161, P1_R2278_U418);
  not ginst1915 (P1_R2278_U377, P1_R2278_U80);
  not ginst1916 (P1_R2278_U378, P1_R2278_U73);
  nand ginst1917 (P1_R2278_U379, P1_R2278_U320, P1_R2278_U321);
  not ginst1918 (P1_R2278_U38, P1_INSTADDRPOINTER_REG_4__SCAN_IN);
  not ginst1919 (P1_R2278_U380, P1_R2278_U94);
  nand ginst1920 (P1_R2278_U381, P1_R2278_U314, P1_R2278_U370);
  nand ginst1921 (P1_R2278_U382, P1_R2278_U229, P1_R2278_U285, P1_R2278_U391);
  not ginst1922 (P1_R2278_U383, P1_R2278_U92);
  not ginst1923 (P1_R2278_U384, P1_R2278_U95);
  nand ginst1924 (P1_R2278_U385, P1_R2278_U11, P1_R2278_U142, P1_R2278_U411);
  not ginst1925 (P1_R2278_U386, P1_R2278_U93);
  not ginst1926 (P1_R2278_U387, P1_R2278_U96);
  nand ginst1927 (P1_R2278_U388, P1_R2278_U261, P1_R2278_U277);
  nand ginst1928 (P1_R2278_U389, P1_R2278_U228, P1_R2278_U388);
  not ginst1929 (P1_R2278_U39, P1_U2796);
  nand ginst1930 (P1_R2278_U390, P1_R2278_U229, P1_R2278_U285, P1_R2278_U391);
  nand ginst1931 (P1_R2278_U391, P1_R2278_U282, P1_R2278_U283);
  not ginst1932 (P1_R2278_U392, P1_R2278_U86);
  nand ginst1933 (P1_R2278_U393, P1_INSTADDRPOINTER_REG_30__SCAN_IN, P1_U2770);
  nand ginst1934 (P1_R2278_U394, P1_R2278_U148, P1_R2278_U372);
  nand ginst1935 (P1_R2278_U395, P1_R2278_U324, P1_R2278_U383);
  nand ginst1936 (P1_R2278_U396, P1_R2278_U150, P1_R2278_U368);
  nand ginst1937 (P1_R2278_U397, P1_R2278_U152, P1_R2278_U153, P1_R2278_U413);
  nand ginst1938 (P1_R2278_U398, P1_R2278_U324, P1_R2278_U386);
  nand ginst1939 (P1_R2278_U399, P1_R2278_U11, P1_R2278_U154, P1_R2278_U378);
  nand ginst1940 (P1_R2278_U40, P1_R2278_U250, P1_R2278_U43);
  nand ginst1941 (P1_R2278_U400, P1_R2278_U324, P1_R2278_U86);
  not ginst1942 (P1_R2278_U401, P1_R2278_U87);
  nand ginst1943 (P1_R2278_U402, P1_R2278_U229, P1_R2278_U285, P1_R2278_U391);
  nand ginst1944 (P1_R2278_U403, P1_R2278_U324, P1_R2278_U380);
  nand ginst1945 (P1_R2278_U404, P1_R2278_U324, P1_R2278_U384);
  nand ginst1946 (P1_R2278_U405, P1_R2278_U157, P1_R2278_U158, P1_R2278_U411);
  nand ginst1947 (P1_R2278_U406, P1_R2278_U324, P1_R2278_U387);
  nand ginst1948 (P1_R2278_U407, P1_R2278_U324, P1_R2278_U87);
  nand ginst1949 (P1_R2278_U408, P1_R2278_U374, P1_R2278_U85);
  nand ginst1950 (P1_R2278_U409, P1_R2278_U319, P1_R2278_U408);
  nand ginst1951 (P1_R2278_U41, P1_R2278_U252, P1_R2278_U253, P1_R2278_U254);
  nand ginst1952 (P1_R2278_U410, P1_R2278_U227, P1_R2278_U402);
  nand ginst1953 (P1_R2278_U411, P1_R2278_U141, P1_R2278_U226);
  nand ginst1954 (P1_R2278_U412, P1_R2278_U227, P1_R2278_U390);
  nand ginst1955 (P1_R2278_U413, P1_R2278_U151, P1_R2278_U226);
  nand ginst1956 (P1_R2278_U414, P1_R2278_U174, P1_R2278_U336);
  nand ginst1957 (P1_R2278_U415, P1_R2278_U227, P1_R2278_U287);
  not ginst1958 (P1_R2278_U416, P1_R2278_U222);
  nand ginst1959 (P1_R2278_U417, P1_R2278_U227, P1_R2278_U382);
  nand ginst1960 (P1_R2278_U418, P1_R2278_U160, P1_R2278_U226);
  nand ginst1961 (P1_R2278_U419, P1_R2278_U11, P1_R2278_U206);
  nand ginst1962 (P1_R2278_U42, P1_R2278_U245, P1_R2278_U246);
  not ginst1963 (P1_R2278_U420, P1_R2278_U196);
  nand ginst1964 (P1_R2278_U421, P1_R2278_U206, P1_R2278_U311);
  not ginst1965 (P1_R2278_U422, P1_R2278_U204);
  nand ginst1966 (P1_R2278_U423, P1_R2278_U10, P1_R2278_U206);
  not ginst1967 (P1_R2278_U424, P1_R2278_U200);
  nand ginst1968 (P1_R2278_U425, P1_R2278_U164, P1_R2278_U206);
  not ginst1969 (P1_R2278_U426, P1_R2278_U198);
  nand ginst1970 (P1_R2278_U427, P1_R2278_U166, P1_R2278_U206);
  not ginst1971 (P1_R2278_U428, P1_R2278_U202);
  nand ginst1972 (P1_R2278_U429, P1_R2278_U33, P1_R2278_U557);
  nand ginst1973 (P1_R2278_U43, P1_R2278_U248, P1_R2278_U42);
  nand ginst1974 (P1_R2278_U430, P1_R2278_U176, P1_R2278_U346);
  nand ginst1975 (P1_R2278_U431, P1_R2278_U100, P1_R2278_U260);
  nand ginst1976 (P1_R2278_U432, P1_R2278_U21, P1_U2792);
  nand ginst1977 (P1_R2278_U433, P1_INSTADDRPOINTER_REG_8__SCAN_IN, P1_R2278_U22);
  nand ginst1978 (P1_R2278_U434, P1_R2278_U21, P1_U2792);
  nand ginst1979 (P1_R2278_U435, P1_INSTADDRPOINTER_REG_8__SCAN_IN, P1_R2278_U22);
  nand ginst1980 (P1_R2278_U436, P1_R2278_U434, P1_R2278_U435);
  nand ginst1981 (P1_R2278_U437, P1_R2278_U177, P1_R2278_U178);
  nand ginst1982 (P1_R2278_U438, P1_R2278_U257, P1_R2278_U436);
  nand ginst1983 (P1_R2278_U439, P1_R2278_U23, P1_U2793);
  not ginst1984 (P1_R2278_U44, P1_INSTADDRPOINTER_REG_25__SCAN_IN);
  nand ginst1985 (P1_R2278_U440, P1_INSTADDRPOINTER_REG_7__SCAN_IN, P1_R2278_U24);
  nand ginst1986 (P1_R2278_U441, P1_R2278_U25, P1_U2794);
  nand ginst1987 (P1_R2278_U442, P1_INSTADDRPOINTER_REG_6__SCAN_IN, P1_R2278_U26);
  nand ginst1988 (P1_R2278_U443, P1_R2278_U441, P1_R2278_U442);
  nand ginst1989 (P1_R2278_U444, P1_R2278_U347, P1_R2278_U40);
  nand ginst1990 (P1_R2278_U445, P1_R2278_U251, P1_R2278_U443);
  nand ginst1991 (P1_R2278_U446, P1_R2278_U27, P1_U2795);
  nand ginst1992 (P1_R2278_U447, P1_INSTADDRPOINTER_REG_5__SCAN_IN, P1_R2278_U28);
  nand ginst1993 (P1_R2278_U448, P1_R2278_U38, P1_U2796);
  nand ginst1994 (P1_R2278_U449, P1_INSTADDRPOINTER_REG_4__SCAN_IN, P1_R2278_U39);
  not ginst1995 (P1_R2278_U45, P1_U2775);
  nand ginst1996 (P1_R2278_U450, P1_R2278_U38, P1_U2796);
  nand ginst1997 (P1_R2278_U451, P1_INSTADDRPOINTER_REG_4__SCAN_IN, P1_R2278_U39);
  nand ginst1998 (P1_R2278_U452, P1_R2278_U450, P1_R2278_U451);
  nand ginst1999 (P1_R2278_U453, P1_R2278_U181, P1_R2278_U182);
  nand ginst2000 (P1_R2278_U454, P1_R2278_U243, P1_R2278_U452);
  nand ginst2001 (P1_R2278_U455, P1_R2278_U36, P1_U2797);
  nand ginst2002 (P1_R2278_U456, P1_INSTADDRPOINTER_REG_3__SCAN_IN, P1_R2278_U37);
  nand ginst2003 (P1_R2278_U457, P1_R2278_U36, P1_U2797);
  nand ginst2004 (P1_R2278_U458, P1_INSTADDRPOINTER_REG_3__SCAN_IN, P1_R2278_U37);
  nand ginst2005 (P1_R2278_U459, P1_R2278_U457, P1_R2278_U458);
  not ginst2006 (P1_R2278_U46, P1_INSTADDRPOINTER_REG_26__SCAN_IN);
  nand ginst2007 (P1_R2278_U460, P1_R2278_U183, P1_R2278_U184);
  nand ginst2008 (P1_R2278_U461, P1_R2278_U239, P1_R2278_U459);
  nand ginst2009 (P1_R2278_U462, P1_INSTADDRPOINTER_REG_31__SCAN_IN, P1_R2278_U186);
  nand ginst2010 (P1_R2278_U463, P1_R2278_U185, P1_U2769);
  nand ginst2011 (P1_R2278_U464, P1_INSTADDRPOINTER_REG_31__SCAN_IN, P1_R2278_U186);
  nand ginst2012 (P1_R2278_U465, P1_R2278_U185, P1_U2769);
  nand ginst2013 (P1_R2278_U466, P1_R2278_U464, P1_R2278_U465);
  nand ginst2014 (P1_R2278_U467, P1_R2278_U155, P1_R2278_U187, P1_R2278_U396, P1_R2278_U397);
  nand ginst2015 (P1_R2278_U468, P1_R2278_U325, P1_R2278_U5);
  nand ginst2016 (P1_R2278_U469, P1_R2278_U14, P1_R2278_U88, P1_R2278_U89);
  not ginst2017 (P1_R2278_U47, P1_U2774);
  nand ginst2018 (P1_R2278_U470, P1_INSTADDRPOINTER_REG_30__SCAN_IN, P1_R2278_U466, P1_U2770);
  nand ginst2019 (P1_R2278_U471, P1_INSTADDRPOINTER_REG_30__SCAN_IN, P1_R2278_U88);
  nand ginst2020 (P1_R2278_U472, P1_R2278_U89, P1_U2770);
  nand ginst2021 (P1_R2278_U473, P1_INSTADDRPOINTER_REG_30__SCAN_IN, P1_R2278_U88);
  nand ginst2022 (P1_R2278_U474, P1_R2278_U89, P1_U2770);
  nand ginst2023 (P1_R2278_U475, P1_R2278_U473, P1_R2278_U474);
  nand ginst2024 (P1_R2278_U476, P1_R2278_U189, P1_R2278_U190);
  nand ginst2025 (P1_R2278_U477, P1_R2278_U326, P1_R2278_U475);
  nand ginst2026 (P1_R2278_U478, P1_R2278_U34, P1_U2798);
  nand ginst2027 (P1_R2278_U479, P1_INSTADDRPOINTER_REG_2__SCAN_IN, P1_R2278_U35);
  not ginst2028 (P1_R2278_U48, P1_INSTADDRPOINTER_REG_24__SCAN_IN);
  nand ginst2029 (P1_R2278_U480, P1_R2278_U34, P1_U2798);
  nand ginst2030 (P1_R2278_U481, P1_INSTADDRPOINTER_REG_2__SCAN_IN, P1_R2278_U35);
  nand ginst2031 (P1_R2278_U482, P1_R2278_U480, P1_R2278_U481);
  nand ginst2032 (P1_R2278_U483, P1_R2278_U191, P1_R2278_U192);
  nand ginst2033 (P1_R2278_U484, P1_R2278_U235, P1_R2278_U482);
  nand ginst2034 (P1_R2278_U485, P1_INSTADDRPOINTER_REG_29__SCAN_IN, P1_R2278_U90);
  nand ginst2035 (P1_R2278_U486, P1_R2278_U91, P1_U2771);
  nand ginst2036 (P1_R2278_U487, P1_INSTADDRPOINTER_REG_29__SCAN_IN, P1_R2278_U90);
  nand ginst2037 (P1_R2278_U488, P1_R2278_U91, P1_U2771);
  nand ginst2038 (P1_R2278_U489, P1_R2278_U487, P1_R2278_U488);
  not ginst2039 (P1_R2278_U49, P1_U2776);
  nand ginst2040 (P1_R2278_U490, P1_R2278_U193, P1_R2278_U194);
  nand ginst2041 (P1_R2278_U491, P1_R2278_U323, P1_R2278_U489);
  nand ginst2042 (P1_R2278_U492, P1_INSTADDRPOINTER_REG_28__SCAN_IN, P1_R2278_U81);
  nand ginst2043 (P1_R2278_U493, P1_R2278_U82, P1_U2772);
  nand ginst2044 (P1_R2278_U494, P1_INSTADDRPOINTER_REG_28__SCAN_IN, P1_R2278_U81);
  nand ginst2045 (P1_R2278_U495, P1_R2278_U82, P1_U2772);
  nand ginst2046 (P1_R2278_U496, P1_R2278_U494, P1_R2278_U495);
  nand ginst2047 (P1_R2278_U497, P1_R2278_U195, P1_R2278_U196);
  nand ginst2048 (P1_R2278_U498, P1_R2278_U420, P1_R2278_U496);
  nand ginst2049 (P1_R2278_U499, P1_R2278_U83, P1_U2773);
  and ginst2050 (P1_R2278_U5, P1_R2278_U327, P1_R2278_U466);
  not ginst2051 (P1_R2278_U50, P1_INSTADDRPOINTER_REG_23__SCAN_IN);
  nand ginst2052 (P1_R2278_U500, P1_INSTADDRPOINTER_REG_27__SCAN_IN, P1_R2278_U84);
  nand ginst2053 (P1_R2278_U501, P1_R2278_U83, P1_U2773);
  nand ginst2054 (P1_R2278_U502, P1_INSTADDRPOINTER_REG_27__SCAN_IN, P1_R2278_U84);
  nand ginst2055 (P1_R2278_U503, P1_R2278_U501, P1_R2278_U502);
  nand ginst2056 (P1_R2278_U504, P1_R2278_U197, P1_R2278_U198);
  nand ginst2057 (P1_R2278_U505, P1_R2278_U426, P1_R2278_U503);
  nand ginst2058 (P1_R2278_U506, P1_R2278_U46, P1_U2774);
  nand ginst2059 (P1_R2278_U507, P1_INSTADDRPOINTER_REG_26__SCAN_IN, P1_R2278_U47);
  nand ginst2060 (P1_R2278_U508, P1_R2278_U46, P1_U2774);
  nand ginst2061 (P1_R2278_U509, P1_INSTADDRPOINTER_REG_26__SCAN_IN, P1_R2278_U47);
  not ginst2062 (P1_R2278_U51, P1_U2777);
  nand ginst2063 (P1_R2278_U510, P1_R2278_U508, P1_R2278_U509);
  nand ginst2064 (P1_R2278_U511, P1_R2278_U199, P1_R2278_U200);
  nand ginst2065 (P1_R2278_U512, P1_R2278_U424, P1_R2278_U510);
  nand ginst2066 (P1_R2278_U513, P1_R2278_U44, P1_U2775);
  nand ginst2067 (P1_R2278_U514, P1_INSTADDRPOINTER_REG_25__SCAN_IN, P1_R2278_U45);
  nand ginst2068 (P1_R2278_U515, P1_R2278_U44, P1_U2775);
  nand ginst2069 (P1_R2278_U516, P1_INSTADDRPOINTER_REG_25__SCAN_IN, P1_R2278_U45);
  nand ginst2070 (P1_R2278_U517, P1_R2278_U515, P1_R2278_U516);
  nand ginst2071 (P1_R2278_U518, P1_R2278_U201, P1_R2278_U202);
  nand ginst2072 (P1_R2278_U519, P1_R2278_U428, P1_R2278_U517);
  not ginst2073 (P1_R2278_U52, P1_INSTADDRPOINTER_REG_21__SCAN_IN);
  nand ginst2074 (P1_R2278_U520, P1_R2278_U48, P1_U2776);
  nand ginst2075 (P1_R2278_U521, P1_INSTADDRPOINTER_REG_24__SCAN_IN, P1_R2278_U49);
  nand ginst2076 (P1_R2278_U522, P1_R2278_U48, P1_U2776);
  nand ginst2077 (P1_R2278_U523, P1_INSTADDRPOINTER_REG_24__SCAN_IN, P1_R2278_U49);
  nand ginst2078 (P1_R2278_U524, P1_R2278_U522, P1_R2278_U523);
  nand ginst2079 (P1_R2278_U525, P1_R2278_U203, P1_R2278_U204);
  nand ginst2080 (P1_R2278_U526, P1_R2278_U422, P1_R2278_U524);
  nand ginst2081 (P1_R2278_U527, P1_R2278_U50, P1_U2777);
  nand ginst2082 (P1_R2278_U528, P1_INSTADDRPOINTER_REG_23__SCAN_IN, P1_R2278_U51);
  nand ginst2083 (P1_R2278_U529, P1_R2278_U50, P1_U2777);
  not ginst2084 (P1_R2278_U53, P1_U2779);
  nand ginst2085 (P1_R2278_U530, P1_INSTADDRPOINTER_REG_23__SCAN_IN, P1_R2278_U51);
  nand ginst2086 (P1_R2278_U531, P1_R2278_U529, P1_R2278_U530);
  nand ginst2087 (P1_R2278_U532, P1_R2278_U205, P1_R2278_U206);
  nand ginst2088 (P1_R2278_U533, P1_R2278_U310, P1_R2278_U531);
  nand ginst2089 (P1_R2278_U534, P1_R2278_U74, P1_U2778);
  nand ginst2090 (P1_R2278_U535, P1_INSTADDRPOINTER_REG_22__SCAN_IN, P1_R2278_U75);
  nand ginst2091 (P1_R2278_U536, P1_R2278_U74, P1_U2778);
  nand ginst2092 (P1_R2278_U537, P1_INSTADDRPOINTER_REG_22__SCAN_IN, P1_R2278_U75);
  nand ginst2093 (P1_R2278_U538, P1_R2278_U536, P1_R2278_U537);
  nand ginst2094 (P1_R2278_U539, P1_R2278_U207, P1_R2278_U208);
  not ginst2095 (P1_R2278_U54, P1_INSTADDRPOINTER_REG_20__SCAN_IN);
  nand ginst2096 (P1_R2278_U540, P1_R2278_U307, P1_R2278_U538);
  nand ginst2097 (P1_R2278_U541, P1_R2278_U52, P1_U2779);
  nand ginst2098 (P1_R2278_U542, P1_INSTADDRPOINTER_REG_21__SCAN_IN, P1_R2278_U53);
  nand ginst2099 (P1_R2278_U543, P1_R2278_U52, P1_U2779);
  nand ginst2100 (P1_R2278_U544, P1_INSTADDRPOINTER_REG_21__SCAN_IN, P1_R2278_U53);
  nand ginst2101 (P1_R2278_U545, P1_R2278_U543, P1_R2278_U544);
  nand ginst2102 (P1_R2278_U546, P1_R2278_U209, P1_R2278_U210);
  nand ginst2103 (P1_R2278_U547, P1_R2278_U304, P1_R2278_U545);
  nand ginst2104 (P1_R2278_U548, P1_R2278_U54, P1_U2780);
  nand ginst2105 (P1_R2278_U549, P1_INSTADDRPOINTER_REG_20__SCAN_IN, P1_R2278_U55);
  not ginst2106 (P1_R2278_U55, P1_U2780);
  nand ginst2107 (P1_R2278_U550, P1_R2278_U54, P1_U2780);
  nand ginst2108 (P1_R2278_U551, P1_INSTADDRPOINTER_REG_20__SCAN_IN, P1_R2278_U55);
  nand ginst2109 (P1_R2278_U552, P1_R2278_U550, P1_R2278_U551);
  nand ginst2110 (P1_R2278_U553, P1_R2278_U211, P1_R2278_U212);
  nand ginst2111 (P1_R2278_U554, P1_R2278_U301, P1_R2278_U552);
  nand ginst2112 (P1_R2278_U555, P1_INSTADDRPOINTER_REG_1__SCAN_IN, P1_R2278_U32);
  nand ginst2113 (P1_R2278_U556, P1_R2278_U232, P1_R2278_U31);
  nand ginst2114 (P1_R2278_U557, P1_R2278_U555, P1_R2278_U556);
  nand ginst2115 (P1_R2278_U558, P1_R2278_U31, P1_R2278_U32, P1_U2799);
  nand ginst2116 (P1_R2278_U559, P1_INSTADDRPOINTER_REG_1__SCAN_IN, P1_R2278_U230);
  not ginst2117 (P1_R2278_U56, P1_INSTADDRPOINTER_REG_19__SCAN_IN);
  nand ginst2118 (P1_R2278_U560, P1_R2278_U56, P1_U2781);
  nand ginst2119 (P1_R2278_U561, P1_INSTADDRPOINTER_REG_19__SCAN_IN, P1_R2278_U57);
  nand ginst2120 (P1_R2278_U562, P1_R2278_U56, P1_U2781);
  nand ginst2121 (P1_R2278_U563, P1_INSTADDRPOINTER_REG_19__SCAN_IN, P1_R2278_U57);
  nand ginst2122 (P1_R2278_U564, P1_R2278_U562, P1_R2278_U563);
  nand ginst2123 (P1_R2278_U565, P1_R2278_U215, P1_R2278_U216);
  nand ginst2124 (P1_R2278_U566, P1_R2278_U297, P1_R2278_U564);
  nand ginst2125 (P1_R2278_U567, P1_R2278_U77, P1_U2782);
  nand ginst2126 (P1_R2278_U568, P1_INSTADDRPOINTER_REG_18__SCAN_IN, P1_R2278_U78);
  nand ginst2127 (P1_R2278_U569, P1_R2278_U77, P1_U2782);
  not ginst2128 (P1_R2278_U57, P1_U2781);
  nand ginst2129 (P1_R2278_U570, P1_INSTADDRPOINTER_REG_18__SCAN_IN, P1_R2278_U78);
  nand ginst2130 (P1_R2278_U571, P1_R2278_U569, P1_R2278_U570);
  nand ginst2131 (P1_R2278_U572, P1_R2278_U217, P1_R2278_U218);
  nand ginst2132 (P1_R2278_U573, P1_R2278_U294, P1_R2278_U571);
  nand ginst2133 (P1_R2278_U574, P1_R2278_U71, P1_U2783);
  nand ginst2134 (P1_R2278_U575, P1_INSTADDRPOINTER_REG_17__SCAN_IN, P1_R2278_U72);
  nand ginst2135 (P1_R2278_U576, P1_R2278_U71, P1_U2783);
  nand ginst2136 (P1_R2278_U577, P1_INSTADDRPOINTER_REG_17__SCAN_IN, P1_R2278_U72);
  nand ginst2137 (P1_R2278_U578, P1_R2278_U576, P1_R2278_U577);
  nand ginst2138 (P1_R2278_U579, P1_R2278_U219, P1_R2278_U220);
  not ginst2139 (P1_R2278_U58, P1_INSTADDRPOINTER_REG_11__SCAN_IN);
  nand ginst2140 (P1_R2278_U580, P1_R2278_U291, P1_R2278_U578);
  nand ginst2141 (P1_R2278_U581, P1_R2278_U69, P1_U2784);
  nand ginst2142 (P1_R2278_U582, P1_INSTADDRPOINTER_REG_16__SCAN_IN, P1_R2278_U70);
  nand ginst2143 (P1_R2278_U583, P1_R2278_U69, P1_U2784);
  nand ginst2144 (P1_R2278_U584, P1_INSTADDRPOINTER_REG_16__SCAN_IN, P1_R2278_U70);
  nand ginst2145 (P1_R2278_U585, P1_R2278_U583, P1_R2278_U584);
  nand ginst2146 (P1_R2278_U586, P1_R2278_U221, P1_R2278_U222);
  nand ginst2147 (P1_R2278_U587, P1_R2278_U416, P1_R2278_U585);
  nand ginst2148 (P1_R2278_U588, P1_R2278_U62, P1_U2785);
  nand ginst2149 (P1_R2278_U589, P1_INSTADDRPOINTER_REG_15__SCAN_IN, P1_R2278_U63);
  not ginst2150 (P1_R2278_U59, P1_U2789);
  nand ginst2151 (P1_R2278_U590, P1_R2278_U66, P1_U2786);
  nand ginst2152 (P1_R2278_U591, P1_INSTADDRPOINTER_REG_14__SCAN_IN, P1_R2278_U67);
  nand ginst2153 (P1_R2278_U592, P1_R2278_U590, P1_R2278_U591);
  nand ginst2154 (P1_R2278_U593, P1_R2278_U348, P1_R2278_U97);
  nand ginst2155 (P1_R2278_U594, P1_R2278_U332, P1_R2278_U592);
  nand ginst2156 (P1_R2278_U595, P1_R2278_U64, P1_U2787);
  nand ginst2157 (P1_R2278_U596, P1_INSTADDRPOINTER_REG_13__SCAN_IN, P1_R2278_U65);
  nand ginst2158 (P1_R2278_U597, P1_R2278_U595, P1_R2278_U596);
  nand ginst2159 (P1_R2278_U598, P1_R2278_U223, P1_R2278_U349);
  nand ginst2160 (P1_R2278_U599, P1_R2278_U329, P1_R2278_U597);
  and ginst2161 (P1_R2278_U6, P1_R2278_U288, P1_R2278_U292);
  not ginst2162 (P1_R2278_U60, P1_INSTADDRPOINTER_REG_10__SCAN_IN);
  nand ginst2163 (P1_R2278_U600, P1_R2278_U224, P1_R2278_U350);
  nand ginst2164 (P1_R2278_U601, P1_R2278_U124, P1_R2278_U280);
  nand ginst2165 (P1_R2278_U602, P1_R2278_U58, P1_U2789);
  nand ginst2166 (P1_R2278_U603, P1_INSTADDRPOINTER_REG_11__SCAN_IN, P1_R2278_U59);
  nand ginst2167 (P1_R2278_U604, P1_R2278_U60, P1_U2790);
  nand ginst2168 (P1_R2278_U605, P1_INSTADDRPOINTER_REG_10__SCAN_IN, P1_R2278_U61);
  nand ginst2169 (P1_R2278_U606, P1_R2278_U604, P1_R2278_U605);
  nand ginst2170 (P1_R2278_U607, P1_R2278_U225, P1_R2278_U351);
  nand ginst2171 (P1_R2278_U608, P1_R2278_U275, P1_R2278_U606);
  nand ginst2172 (P1_R2278_U609, P1_INSTADDRPOINTER_REG_0__SCAN_IN, P1_R2278_U29);
  not ginst2173 (P1_R2278_U61, P1_U2790);
  nand ginst2174 (P1_R2278_U610, P1_R2278_U30, P1_U2800);
  not ginst2175 (P1_R2278_U62, P1_INSTADDRPOINTER_REG_15__SCAN_IN);
  not ginst2176 (P1_R2278_U63, P1_U2785);
  not ginst2177 (P1_R2278_U64, P1_INSTADDRPOINTER_REG_13__SCAN_IN);
  not ginst2178 (P1_R2278_U65, P1_U2787);
  not ginst2179 (P1_R2278_U66, P1_INSTADDRPOINTER_REG_14__SCAN_IN);
  not ginst2180 (P1_R2278_U67, P1_U2786);
  nand ginst2181 (P1_R2278_U68, P1_INSTADDRPOINTER_REG_12__SCAN_IN, P1_U2788);
  not ginst2182 (P1_R2278_U69, P1_INSTADDRPOINTER_REG_16__SCAN_IN);
  and ginst2183 (P1_R2278_U7, P1_R2278_U295, P1_R2278_U6);
  not ginst2184 (P1_R2278_U70, P1_U2784);
  not ginst2185 (P1_R2278_U71, P1_INSTADDRPOINTER_REG_17__SCAN_IN);
  not ginst2186 (P1_R2278_U72, P1_U2783);
  nand ginst2187 (P1_R2278_U73, P1_R2278_U12, P1_R2278_U308, P1_R2278_U359, P1_R2278_U8);
  not ginst2188 (P1_R2278_U74, P1_INSTADDRPOINTER_REG_22__SCAN_IN);
  not ginst2189 (P1_R2278_U75, P1_U2778);
  nand ginst2190 (P1_R2278_U76, P1_INSTADDRPOINTER_REG_22__SCAN_IN, P1_U2778);
  not ginst2191 (P1_R2278_U77, P1_INSTADDRPOINTER_REG_18__SCAN_IN);
  not ginst2192 (P1_R2278_U78, P1_U2782);
  nand ginst2193 (P1_R2278_U79, P1_INSTADDRPOINTER_REG_18__SCAN_IN, P1_U2782);
  and ginst2194 (P1_R2278_U8, P1_R2278_U298, P1_R2278_U302, P1_R2278_U305);
  nand ginst2195 (P1_R2278_U80, P1_R2278_U144, P1_R2278_U8);
  not ginst2196 (P1_R2278_U81, P1_U2772);
  not ginst2197 (P1_R2278_U82, P1_INSTADDRPOINTER_REG_28__SCAN_IN);
  not ginst2198 (P1_R2278_U83, P1_INSTADDRPOINTER_REG_27__SCAN_IN);
  not ginst2199 (P1_R2278_U84, P1_U2773);
  nand ginst2200 (P1_R2278_U85, P1_INSTADDRPOINTER_REG_27__SCAN_IN, P1_U2773);
  nand ginst2201 (P1_R2278_U86, P1_R2278_U322, P1_R2278_U379);
  nand ginst2202 (P1_R2278_U87, P1_R2278_U392, P1_R2278_U92, P1_R2278_U93);
  not ginst2203 (P1_R2278_U88, P1_U2770);
  not ginst2204 (P1_R2278_U89, P1_INSTADDRPOINTER_REG_30__SCAN_IN);
  and ginst2205 (P1_R2278_U9, P1_R2278_U308, P1_R2278_U8);
  not ginst2206 (P1_R2278_U90, P1_U2771);
  not ginst2207 (P1_R2278_U91, P1_INSTADDRPOINTER_REG_29__SCAN_IN);
  nand ginst2208 (P1_R2278_U92, P1_R2278_U11, P1_R2278_U143);
  nand ginst2209 (P1_R2278_U93, P1_R2278_U11, P1_R2278_U321, P1_R2278_U377);
  nand ginst2210 (P1_R2278_U94, P1_R2278_U132, P1_R2278_U372);
  nand ginst2211 (P1_R2278_U95, P1_R2278_U136, P1_R2278_U368);
  nand ginst2212 (P1_R2278_U96, P1_R2278_U11, P1_R2278_U321, P1_R2278_U378);
  nand ginst2213 (P1_R2278_U97, P1_R2278_U229, P1_R2278_U331);
  nand ginst2214 (P1_R2278_U98, P1_R2278_U138, P1_R2278_U354);
  nand ginst2215 (P1_R2278_U99, P1_R2278_U609, P1_R2278_U610);
  nand ginst2216 (P1_R2337_U10, P1_PHYADDRPOINTER_REG_4__SCAN_IN, P1_R2337_U95);
  not ginst2217 (P1_R2337_U100, P1_R2337_U19);
  not ginst2218 (P1_R2337_U101, P1_R2337_U20);
  not ginst2219 (P1_R2337_U102, P1_R2337_U22);
  not ginst2220 (P1_R2337_U103, P1_R2337_U24);
  not ginst2221 (P1_R2337_U104, P1_R2337_U26);
  not ginst2222 (P1_R2337_U105, P1_R2337_U28);
  not ginst2223 (P1_R2337_U106, P1_R2337_U30);
  not ginst2224 (P1_R2337_U107, P1_R2337_U32);
  not ginst2225 (P1_R2337_U108, P1_R2337_U34);
  not ginst2226 (P1_R2337_U109, P1_R2337_U36);
  not ginst2227 (P1_R2337_U11, P1_PHYADDRPOINTER_REG_5__SCAN_IN);
  not ginst2228 (P1_R2337_U110, P1_R2337_U38);
  not ginst2229 (P1_R2337_U111, P1_R2337_U40);
  not ginst2230 (P1_R2337_U112, P1_R2337_U42);
  not ginst2231 (P1_R2337_U113, P1_R2337_U44);
  not ginst2232 (P1_R2337_U114, P1_R2337_U46);
  not ginst2233 (P1_R2337_U115, P1_R2337_U48);
  not ginst2234 (P1_R2337_U116, P1_R2337_U50);
  not ginst2235 (P1_R2337_U117, P1_R2337_U52);
  not ginst2236 (P1_R2337_U118, P1_R2337_U54);
  not ginst2237 (P1_R2337_U119, P1_R2337_U56);
  nand ginst2238 (P1_R2337_U12, P1_PHYADDRPOINTER_REG_5__SCAN_IN, P1_R2337_U96);
  not ginst2239 (P1_R2337_U120, P1_R2337_U58);
  not ginst2240 (P1_R2337_U121, P1_R2337_U60);
  not ginst2241 (P1_R2337_U122, P1_R2337_U93);
  nand ginst2242 (P1_R2337_U123, P1_PHYADDRPOINTER_REG_9__SCAN_IN, P1_R2337_U19);
  nand ginst2243 (P1_R2337_U124, P1_R2337_U100, P1_R2337_U18);
  nand ginst2244 (P1_R2337_U125, P1_PHYADDRPOINTER_REG_8__SCAN_IN, P1_R2337_U16);
  nand ginst2245 (P1_R2337_U126, P1_R2337_U17, P1_R2337_U99);
  nand ginst2246 (P1_R2337_U127, P1_PHYADDRPOINTER_REG_7__SCAN_IN, P1_R2337_U14);
  nand ginst2247 (P1_R2337_U128, P1_R2337_U15, P1_R2337_U98);
  nand ginst2248 (P1_R2337_U129, P1_PHYADDRPOINTER_REG_6__SCAN_IN, P1_R2337_U12);
  not ginst2249 (P1_R2337_U13, P1_PHYADDRPOINTER_REG_6__SCAN_IN);
  nand ginst2250 (P1_R2337_U130, P1_R2337_U13, P1_R2337_U97);
  nand ginst2251 (P1_R2337_U131, P1_PHYADDRPOINTER_REG_5__SCAN_IN, P1_R2337_U10);
  nand ginst2252 (P1_R2337_U132, P1_R2337_U11, P1_R2337_U96);
  nand ginst2253 (P1_R2337_U133, P1_PHYADDRPOINTER_REG_4__SCAN_IN, P1_R2337_U8);
  nand ginst2254 (P1_R2337_U134, P1_R2337_U9, P1_R2337_U95);
  nand ginst2255 (P1_R2337_U135, P1_PHYADDRPOINTER_REG_3__SCAN_IN, P1_R2337_U6);
  nand ginst2256 (P1_R2337_U136, P1_R2337_U7, P1_R2337_U94);
  nand ginst2257 (P1_R2337_U137, P1_PHYADDRPOINTER_REG_31__SCAN_IN, P1_R2337_U93);
  nand ginst2258 (P1_R2337_U138, P1_R2337_U122, P1_R2337_U92);
  nand ginst2259 (P1_R2337_U139, P1_PHYADDRPOINTER_REG_30__SCAN_IN, P1_R2337_U60);
  nand ginst2260 (P1_R2337_U14, P1_PHYADDRPOINTER_REG_6__SCAN_IN, P1_R2337_U97);
  nand ginst2261 (P1_R2337_U140, P1_R2337_U121, P1_R2337_U61);
  nand ginst2262 (P1_R2337_U141, P1_PHYADDRPOINTER_REG_2__SCAN_IN, P1_R2337_U4);
  nand ginst2263 (P1_R2337_U142, P1_PHYADDRPOINTER_REG_1__SCAN_IN, P1_R2337_U5);
  nand ginst2264 (P1_R2337_U143, P1_PHYADDRPOINTER_REG_29__SCAN_IN, P1_R2337_U58);
  nand ginst2265 (P1_R2337_U144, P1_R2337_U120, P1_R2337_U59);
  nand ginst2266 (P1_R2337_U145, P1_PHYADDRPOINTER_REG_28__SCAN_IN, P1_R2337_U56);
  nand ginst2267 (P1_R2337_U146, P1_R2337_U119, P1_R2337_U57);
  nand ginst2268 (P1_R2337_U147, P1_PHYADDRPOINTER_REG_27__SCAN_IN, P1_R2337_U54);
  nand ginst2269 (P1_R2337_U148, P1_R2337_U118, P1_R2337_U55);
  nand ginst2270 (P1_R2337_U149, P1_PHYADDRPOINTER_REG_26__SCAN_IN, P1_R2337_U52);
  not ginst2271 (P1_R2337_U15, P1_PHYADDRPOINTER_REG_7__SCAN_IN);
  nand ginst2272 (P1_R2337_U150, P1_R2337_U117, P1_R2337_U53);
  nand ginst2273 (P1_R2337_U151, P1_PHYADDRPOINTER_REG_25__SCAN_IN, P1_R2337_U50);
  nand ginst2274 (P1_R2337_U152, P1_R2337_U116, P1_R2337_U51);
  nand ginst2275 (P1_R2337_U153, P1_PHYADDRPOINTER_REG_24__SCAN_IN, P1_R2337_U48);
  nand ginst2276 (P1_R2337_U154, P1_R2337_U115, P1_R2337_U49);
  nand ginst2277 (P1_R2337_U155, P1_PHYADDRPOINTER_REG_23__SCAN_IN, P1_R2337_U46);
  nand ginst2278 (P1_R2337_U156, P1_R2337_U114, P1_R2337_U47);
  nand ginst2279 (P1_R2337_U157, P1_PHYADDRPOINTER_REG_22__SCAN_IN, P1_R2337_U44);
  nand ginst2280 (P1_R2337_U158, P1_R2337_U113, P1_R2337_U45);
  nand ginst2281 (P1_R2337_U159, P1_PHYADDRPOINTER_REG_21__SCAN_IN, P1_R2337_U42);
  nand ginst2282 (P1_R2337_U16, P1_PHYADDRPOINTER_REG_7__SCAN_IN, P1_R2337_U98);
  nand ginst2283 (P1_R2337_U160, P1_R2337_U112, P1_R2337_U43);
  nand ginst2284 (P1_R2337_U161, P1_PHYADDRPOINTER_REG_20__SCAN_IN, P1_R2337_U40);
  nand ginst2285 (P1_R2337_U162, P1_R2337_U111, P1_R2337_U41);
  nand ginst2286 (P1_R2337_U163, P1_PHYADDRPOINTER_REG_19__SCAN_IN, P1_R2337_U38);
  nand ginst2287 (P1_R2337_U164, P1_R2337_U110, P1_R2337_U39);
  nand ginst2288 (P1_R2337_U165, P1_PHYADDRPOINTER_REG_18__SCAN_IN, P1_R2337_U36);
  nand ginst2289 (P1_R2337_U166, P1_R2337_U109, P1_R2337_U37);
  nand ginst2290 (P1_R2337_U167, P1_PHYADDRPOINTER_REG_17__SCAN_IN, P1_R2337_U34);
  nand ginst2291 (P1_R2337_U168, P1_R2337_U108, P1_R2337_U35);
  nand ginst2292 (P1_R2337_U169, P1_PHYADDRPOINTER_REG_16__SCAN_IN, P1_R2337_U32);
  not ginst2293 (P1_R2337_U17, P1_PHYADDRPOINTER_REG_8__SCAN_IN);
  nand ginst2294 (P1_R2337_U170, P1_R2337_U107, P1_R2337_U33);
  nand ginst2295 (P1_R2337_U171, P1_PHYADDRPOINTER_REG_15__SCAN_IN, P1_R2337_U30);
  nand ginst2296 (P1_R2337_U172, P1_R2337_U106, P1_R2337_U31);
  nand ginst2297 (P1_R2337_U173, P1_PHYADDRPOINTER_REG_14__SCAN_IN, P1_R2337_U28);
  nand ginst2298 (P1_R2337_U174, P1_R2337_U105, P1_R2337_U29);
  nand ginst2299 (P1_R2337_U175, P1_PHYADDRPOINTER_REG_13__SCAN_IN, P1_R2337_U26);
  nand ginst2300 (P1_R2337_U176, P1_R2337_U104, P1_R2337_U27);
  nand ginst2301 (P1_R2337_U177, P1_PHYADDRPOINTER_REG_12__SCAN_IN, P1_R2337_U24);
  nand ginst2302 (P1_R2337_U178, P1_R2337_U103, P1_R2337_U25);
  nand ginst2303 (P1_R2337_U179, P1_PHYADDRPOINTER_REG_11__SCAN_IN, P1_R2337_U22);
  not ginst2304 (P1_R2337_U18, P1_PHYADDRPOINTER_REG_9__SCAN_IN);
  nand ginst2305 (P1_R2337_U180, P1_R2337_U102, P1_R2337_U23);
  nand ginst2306 (P1_R2337_U181, P1_PHYADDRPOINTER_REG_10__SCAN_IN, P1_R2337_U20);
  nand ginst2307 (P1_R2337_U182, P1_R2337_U101, P1_R2337_U21);
  nand ginst2308 (P1_R2337_U19, P1_PHYADDRPOINTER_REG_8__SCAN_IN, P1_R2337_U99);
  nand ginst2309 (P1_R2337_U20, P1_PHYADDRPOINTER_REG_9__SCAN_IN, P1_R2337_U100);
  not ginst2310 (P1_R2337_U21, P1_PHYADDRPOINTER_REG_10__SCAN_IN);
  nand ginst2311 (P1_R2337_U22, P1_PHYADDRPOINTER_REG_10__SCAN_IN, P1_R2337_U101);
  not ginst2312 (P1_R2337_U23, P1_PHYADDRPOINTER_REG_11__SCAN_IN);
  nand ginst2313 (P1_R2337_U24, P1_PHYADDRPOINTER_REG_11__SCAN_IN, P1_R2337_U102);
  not ginst2314 (P1_R2337_U25, P1_PHYADDRPOINTER_REG_12__SCAN_IN);
  nand ginst2315 (P1_R2337_U26, P1_PHYADDRPOINTER_REG_12__SCAN_IN, P1_R2337_U103);
  not ginst2316 (P1_R2337_U27, P1_PHYADDRPOINTER_REG_13__SCAN_IN);
  nand ginst2317 (P1_R2337_U28, P1_PHYADDRPOINTER_REG_13__SCAN_IN, P1_R2337_U104);
  not ginst2318 (P1_R2337_U29, P1_PHYADDRPOINTER_REG_14__SCAN_IN);
  nand ginst2319 (P1_R2337_U30, P1_PHYADDRPOINTER_REG_14__SCAN_IN, P1_R2337_U105);
  not ginst2320 (P1_R2337_U31, P1_PHYADDRPOINTER_REG_15__SCAN_IN);
  nand ginst2321 (P1_R2337_U32, P1_PHYADDRPOINTER_REG_15__SCAN_IN, P1_R2337_U106);
  not ginst2322 (P1_R2337_U33, P1_PHYADDRPOINTER_REG_16__SCAN_IN);
  nand ginst2323 (P1_R2337_U34, P1_PHYADDRPOINTER_REG_16__SCAN_IN, P1_R2337_U107);
  not ginst2324 (P1_R2337_U35, P1_PHYADDRPOINTER_REG_17__SCAN_IN);
  nand ginst2325 (P1_R2337_U36, P1_PHYADDRPOINTER_REG_17__SCAN_IN, P1_R2337_U108);
  not ginst2326 (P1_R2337_U37, P1_PHYADDRPOINTER_REG_18__SCAN_IN);
  nand ginst2327 (P1_R2337_U38, P1_PHYADDRPOINTER_REG_18__SCAN_IN, P1_R2337_U109);
  not ginst2328 (P1_R2337_U39, P1_PHYADDRPOINTER_REG_19__SCAN_IN);
  not ginst2329 (P1_R2337_U4, P1_PHYADDRPOINTER_REG_1__SCAN_IN);
  nand ginst2330 (P1_R2337_U40, P1_PHYADDRPOINTER_REG_19__SCAN_IN, P1_R2337_U110);
  not ginst2331 (P1_R2337_U41, P1_PHYADDRPOINTER_REG_20__SCAN_IN);
  nand ginst2332 (P1_R2337_U42, P1_PHYADDRPOINTER_REG_20__SCAN_IN, P1_R2337_U111);
  not ginst2333 (P1_R2337_U43, P1_PHYADDRPOINTER_REG_21__SCAN_IN);
  nand ginst2334 (P1_R2337_U44, P1_PHYADDRPOINTER_REG_21__SCAN_IN, P1_R2337_U112);
  not ginst2335 (P1_R2337_U45, P1_PHYADDRPOINTER_REG_22__SCAN_IN);
  nand ginst2336 (P1_R2337_U46, P1_PHYADDRPOINTER_REG_22__SCAN_IN, P1_R2337_U113);
  not ginst2337 (P1_R2337_U47, P1_PHYADDRPOINTER_REG_23__SCAN_IN);
  nand ginst2338 (P1_R2337_U48, P1_PHYADDRPOINTER_REG_23__SCAN_IN, P1_R2337_U114);
  not ginst2339 (P1_R2337_U49, P1_PHYADDRPOINTER_REG_24__SCAN_IN);
  not ginst2340 (P1_R2337_U5, P1_PHYADDRPOINTER_REG_2__SCAN_IN);
  nand ginst2341 (P1_R2337_U50, P1_PHYADDRPOINTER_REG_24__SCAN_IN, P1_R2337_U115);
  not ginst2342 (P1_R2337_U51, P1_PHYADDRPOINTER_REG_25__SCAN_IN);
  nand ginst2343 (P1_R2337_U52, P1_PHYADDRPOINTER_REG_25__SCAN_IN, P1_R2337_U116);
  not ginst2344 (P1_R2337_U53, P1_PHYADDRPOINTER_REG_26__SCAN_IN);
  nand ginst2345 (P1_R2337_U54, P1_PHYADDRPOINTER_REG_26__SCAN_IN, P1_R2337_U117);
  not ginst2346 (P1_R2337_U55, P1_PHYADDRPOINTER_REG_27__SCAN_IN);
  nand ginst2347 (P1_R2337_U56, P1_PHYADDRPOINTER_REG_27__SCAN_IN, P1_R2337_U118);
  not ginst2348 (P1_R2337_U57, P1_PHYADDRPOINTER_REG_28__SCAN_IN);
  nand ginst2349 (P1_R2337_U58, P1_PHYADDRPOINTER_REG_28__SCAN_IN, P1_R2337_U119);
  not ginst2350 (P1_R2337_U59, P1_PHYADDRPOINTER_REG_29__SCAN_IN);
  nand ginst2351 (P1_R2337_U6, P1_PHYADDRPOINTER_REG_2__SCAN_IN, P1_PHYADDRPOINTER_REG_1__SCAN_IN);
  nand ginst2352 (P1_R2337_U60, P1_PHYADDRPOINTER_REG_29__SCAN_IN, P1_R2337_U120);
  not ginst2353 (P1_R2337_U61, P1_PHYADDRPOINTER_REG_30__SCAN_IN);
  nand ginst2354 (P1_R2337_U62, P1_R2337_U123, P1_R2337_U124);
  nand ginst2355 (P1_R2337_U63, P1_R2337_U125, P1_R2337_U126);
  nand ginst2356 (P1_R2337_U64, P1_R2337_U127, P1_R2337_U128);
  nand ginst2357 (P1_R2337_U65, P1_R2337_U129, P1_R2337_U130);
  nand ginst2358 (P1_R2337_U66, P1_R2337_U131, P1_R2337_U132);
  nand ginst2359 (P1_R2337_U67, P1_R2337_U133, P1_R2337_U134);
  nand ginst2360 (P1_R2337_U68, P1_R2337_U135, P1_R2337_U136);
  nand ginst2361 (P1_R2337_U69, P1_R2337_U137, P1_R2337_U138);
  not ginst2362 (P1_R2337_U7, P1_PHYADDRPOINTER_REG_3__SCAN_IN);
  nand ginst2363 (P1_R2337_U70, P1_R2337_U139, P1_R2337_U140);
  nand ginst2364 (P1_R2337_U71, P1_R2337_U141, P1_R2337_U142);
  nand ginst2365 (P1_R2337_U72, P1_R2337_U143, P1_R2337_U144);
  nand ginst2366 (P1_R2337_U73, P1_R2337_U145, P1_R2337_U146);
  nand ginst2367 (P1_R2337_U74, P1_R2337_U147, P1_R2337_U148);
  nand ginst2368 (P1_R2337_U75, P1_R2337_U149, P1_R2337_U150);
  nand ginst2369 (P1_R2337_U76, P1_R2337_U151, P1_R2337_U152);
  nand ginst2370 (P1_R2337_U77, P1_R2337_U153, P1_R2337_U154);
  nand ginst2371 (P1_R2337_U78, P1_R2337_U155, P1_R2337_U156);
  nand ginst2372 (P1_R2337_U79, P1_R2337_U157, P1_R2337_U158);
  nand ginst2373 (P1_R2337_U8, P1_PHYADDRPOINTER_REG_3__SCAN_IN, P1_R2337_U94);
  nand ginst2374 (P1_R2337_U80, P1_R2337_U159, P1_R2337_U160);
  nand ginst2375 (P1_R2337_U81, P1_R2337_U161, P1_R2337_U162);
  nand ginst2376 (P1_R2337_U82, P1_R2337_U163, P1_R2337_U164);
  nand ginst2377 (P1_R2337_U83, P1_R2337_U165, P1_R2337_U166);
  nand ginst2378 (P1_R2337_U84, P1_R2337_U167, P1_R2337_U168);
  nand ginst2379 (P1_R2337_U85, P1_R2337_U169, P1_R2337_U170);
  nand ginst2380 (P1_R2337_U86, P1_R2337_U171, P1_R2337_U172);
  nand ginst2381 (P1_R2337_U87, P1_R2337_U173, P1_R2337_U174);
  nand ginst2382 (P1_R2337_U88, P1_R2337_U175, P1_R2337_U176);
  nand ginst2383 (P1_R2337_U89, P1_R2337_U177, P1_R2337_U178);
  not ginst2384 (P1_R2337_U9, P1_PHYADDRPOINTER_REG_4__SCAN_IN);
  nand ginst2385 (P1_R2337_U90, P1_R2337_U179, P1_R2337_U180);
  nand ginst2386 (P1_R2337_U91, P1_R2337_U181, P1_R2337_U182);
  not ginst2387 (P1_R2337_U92, P1_PHYADDRPOINTER_REG_31__SCAN_IN);
  nand ginst2388 (P1_R2337_U93, P1_PHYADDRPOINTER_REG_30__SCAN_IN, P1_R2337_U121);
  not ginst2389 (P1_R2337_U94, P1_R2337_U6);
  not ginst2390 (P1_R2337_U95, P1_R2337_U8);
  not ginst2391 (P1_R2337_U96, P1_R2337_U10);
  not ginst2392 (P1_R2337_U97, P1_R2337_U12);
  not ginst2393 (P1_R2337_U98, P1_R2337_U14);
  not ginst2394 (P1_R2337_U99, P1_R2337_U16);
  and ginst2395 (P1_R2358_U10, P1_R2358_U292, P1_R2358_U9);
  and ginst2396 (P1_R2358_U100, P1_R2358_U284, P1_R2358_U285);
  nand ginst2397 (P1_R2358_U101, P1_R2358_U590, P1_R2358_U591);
  and ginst2398 (P1_R2358_U102, P1_R2358_U282, P1_R2358_U283);
  nand ginst2399 (P1_R2358_U103, P1_R2358_U592, P1_R2358_U593);
  and ginst2400 (P1_R2358_U104, P1_R2358_U280, P1_R2358_U281);
  nand ginst2401 (P1_R2358_U105, P1_R2358_U594, P1_R2358_U595);
  and ginst2402 (P1_R2358_U106, P1_R2358_U205, P1_R2358_U206);
  nand ginst2403 (P1_R2358_U107, P1_R2358_U596, P1_R2358_U597);
  and ginst2404 (P1_R2358_U108, P1_R2358_U278, P1_R2358_U47);
  nand ginst2405 (P1_R2358_U109, P1_R2358_U598, P1_R2358_U599);
  and ginst2406 (P1_R2358_U11, P1_R2358_U457, P1_R2358_U458);
  and ginst2407 (P1_R2358_U110, P1_R2358_U276, P1_R2358_U277);
  nand ginst2408 (P1_R2358_U111, P1_R2358_U600, P1_R2358_U601);
  and ginst2409 (P1_R2358_U112, P1_R2358_U274, P1_R2358_U275);
  nand ginst2410 (P1_R2358_U113, P1_R2358_U602, P1_R2358_U603);
  and ginst2411 (P1_R2358_U114, P1_R2358_U272, P1_R2358_U51);
  nand ginst2412 (P1_R2358_U115, P1_R2358_U604, P1_R2358_U605);
  and ginst2413 (P1_R2358_U116, P1_R2358_U258, P1_R2358_U59);
  nand ginst2414 (P1_R2358_U117, P1_R2358_U606, P1_R2358_U607);
  and ginst2415 (P1_R2358_U118, P1_R2358_U259, P1_R2358_U57);
  nand ginst2416 (P1_R2358_U119, P1_R2358_U608, P1_R2358_U609);
  and ginst2417 (P1_R2358_U12, P1_R2358_U480, P1_R2358_U481);
  and ginst2418 (P1_R2358_U120, P1_R2358_U205, P1_R2358_U208);
  and ginst2419 (P1_R2358_U121, P1_R2358_U202, P1_R2358_U204);
  and ginst2420 (P1_R2358_U122, P1_R2358_U216, P1_R2358_U217);
  and ginst2421 (P1_R2358_U123, P1_R2358_U203, P1_R2358_U204);
  and ginst2422 (P1_R2358_U124, P1_R2358_U229, P1_R2358_U54);
  and ginst2423 (P1_R2358_U125, P1_R2358_U262, P1_R2358_U265);
  and ginst2424 (P1_R2358_U126, P1_R2358_U255, P1_R2358_U258, P1_R2358_U259, P1_R2358_U356);
  and ginst2425 (P1_R2358_U127, P1_R2358_U256, P1_R2358_U353, P1_R2358_U354, P1_R2358_U355);
  and ginst2426 (P1_R2358_U128, P1_R2358_U276, P1_R2358_U5);
  and ginst2427 (P1_R2358_U129, P1_R2358_U277, P1_R2358_U361);
  and ginst2428 (P1_R2358_U13, P1_R2358_U554, P1_R2358_U555);
  and ginst2429 (P1_R2358_U130, P1_R2358_U284, P1_R2358_U7);
  and ginst2430 (P1_R2358_U131, P1_R2358_U285, P1_R2358_U366);
  and ginst2431 (P1_R2358_U132, P1_R2358_U10, P1_R2358_U294);
  and ginst2432 (P1_R2358_U133, P1_R2358_U295, P1_R2358_U373);
  and ginst2433 (P1_R2358_U134, P1_R2358_U305, P1_R2358_U561);
  and ginst2434 (P1_R2358_U135, P1_R2358_U13, P1_R2358_U304);
  and ginst2435 (P1_R2358_U136, P1_R2358_U180, P1_R2358_U374);
  and ginst2436 (P1_R2358_U137, P1_R2358_U289, P1_R2358_U367);
  and ginst2437 (P1_R2358_U138, P1_R2358_U281, P1_R2358_U362);
  and ginst2438 (P1_R2358_U139, P1_R2358_U256, P1_R2358_U257);
  and ginst2439 (P1_R2358_U14, P1_R2358_U329, P1_R2358_U330);
  and ginst2440 (P1_R2358_U140, P1_R2358_U316, P1_R2358_U61);
  and ginst2441 (P1_R2358_U141, P1_R2358_U264, P1_R2358_U265);
  and ginst2442 (P1_R2358_U142, P1_R2358_U263, P1_R2358_U326);
  not ginst2443 (P1_R2358_U143, P1_U2618);
  not ginst2444 (P1_R2358_U144, P1_U2615);
  not ginst2445 (P1_R2358_U145, P1_U2614);
  not ginst2446 (P1_R2358_U146, P1_U2667);
  not ginst2447 (P1_R2358_U147, P1_U2668);
  not ginst2448 (P1_R2358_U148, P1_U2670);
  not ginst2449 (P1_R2358_U149, P1_U2671);
  and ginst2450 (P1_R2358_U15, P1_R2358_U325, P1_R2358_U327);
  not ginst2451 (P1_R2358_U150, P1_U2672);
  not ginst2452 (P1_R2358_U151, P1_U2669);
  not ginst2453 (P1_R2358_U152, P1_U2617);
  nand ginst2454 (P1_R2358_U153, P1_R2358_U228, P1_R2358_U230);
  nand ginst2455 (P1_R2358_U154, P1_R2358_U216, P1_R2358_U224, P1_R2358_U226);
  nand ginst2456 (P1_R2358_U155, P1_R2358_U234, P1_R2358_U28);
  nand ginst2457 (P1_R2358_U156, P1_R2358_U203, P1_R2358_U213);
  not ginst2458 (P1_R2358_U157, P1_U2611);
  not ginst2459 (P1_R2358_U158, P1_U2612);
  not ginst2460 (P1_R2358_U159, P1_U2613);
  and ginst2461 (P1_R2358_U16, P1_R2358_U319, P1_R2358_U320);
  not ginst2462 (P1_R2358_U160, P1_U2616);
  not ginst2463 (P1_R2358_U161, P1_U2610);
  not ginst2464 (P1_R2358_U162, P1_U2609);
  not ginst2465 (P1_R2358_U163, P1_U2666);
  not ginst2466 (P1_R2358_U164, P1_U2665);
  not ginst2467 (P1_R2358_U165, P1_U2664);
  not ginst2468 (P1_R2358_U166, P1_U2660);
  not ginst2469 (P1_R2358_U167, P1_U2661);
  not ginst2470 (P1_R2358_U168, P1_U2663);
  not ginst2471 (P1_R2358_U169, P1_U2662);
  and ginst2472 (P1_R2358_U17, P1_R2358_U315, P1_R2358_U317);
  not ginst2473 (P1_R2358_U170, P1_U2655);
  not ginst2474 (P1_R2358_U171, P1_U2656);
  not ginst2475 (P1_R2358_U172, P1_U2657);
  not ginst2476 (P1_R2358_U173, P1_U2659);
  not ginst2477 (P1_R2358_U174, P1_U2658);
  not ginst2478 (P1_R2358_U175, P1_U2654);
  not ginst2479 (P1_R2358_U176, P1_U2653);
  not ginst2480 (P1_R2358_U177, P1_U2651);
  not ginst2481 (P1_R2358_U178, P1_U2652);
  nand ginst2482 (P1_R2358_U179, P1_R2358_U564, P1_U2621);
  and ginst2483 (P1_R2358_U18, P1_R2358_U307, P1_R2358_U308);
  and ginst2484 (P1_R2358_U180, P1_R2358_U567, P1_R2358_U568);
  and ginst2485 (P1_R2358_U181, P1_R2358_U569, P1_R2358_U570);
  nand ginst2486 (P1_R2358_U182, P1_R2358_U179, P1_R2358_U302);
  nand ginst2487 (P1_R2358_U183, P1_R2358_U297, P1_R2358_U298);
  nand ginst2488 (P1_R2358_U184, P1_R2358_U133, P1_R2358_U383);
  nand ginst2489 (P1_R2358_U185, P1_R2358_U372, P1_R2358_U381);
  nand ginst2490 (P1_R2358_U186, P1_R2358_U370, P1_R2358_U379);
  nand ginst2491 (P1_R2358_U187, P1_R2358_U137, P1_R2358_U377);
  nand ginst2492 (P1_R2358_U188, P1_R2358_U375, P1_R2358_U42);
  nand ginst2493 (P1_R2358_U189, P1_R2358_U131, P1_R2358_U385);
  and ginst2494 (P1_R2358_U19, P1_R2358_U252, P1_R2358_U254);
  nand ginst2495 (P1_R2358_U190, P1_R2358_U365, P1_R2358_U387);
  nand ginst2496 (P1_R2358_U191, P1_R2358_U138, P1_R2358_U389);
  nand ginst2497 (P1_R2358_U192, P1_R2358_U391, P1_R2358_U47);
  nand ginst2498 (P1_R2358_U193, P1_R2358_U209, P1_R2358_U246);
  nand ginst2499 (P1_R2358_U194, P1_R2358_U129, P1_R2358_U393);
  nand ginst2500 (P1_R2358_U195, P1_R2358_U359, P1_R2358_U395);
  nand ginst2501 (P1_R2358_U196, P1_R2358_U397, P1_R2358_U51);
  nand ginst2502 (P1_R2358_U197, P1_R2358_U127, P1_R2358_U201);
  nand ginst2503 (P1_R2358_U198, P1_R2358_U309, P1_R2358_U57);
  nand ginst2504 (P1_R2358_U199, P1_R2358_U264, P1_R2358_U267, P1_R2358_U268);
  and ginst2505 (P1_R2358_U20, P1_R2358_U244, P1_R2358_U245);
  nand ginst2506 (P1_R2358_U200, P1_R2358_U208, P1_R2358_U209);
  nand ginst2507 (P1_R2358_U201, P1_R2358_U126, P1_R2358_U199);
  nand ginst2508 (P1_R2358_U202, P1_R2358_U30, P1_R2358_U435, P1_R2358_U436);
  nand ginst2509 (P1_R2358_U203, P1_R2358_U441, P1_U2647);
  nand ginst2510 (P1_R2358_U204, P1_R2358_U32, P1_R2358_U437, P1_R2358_U438);
  nand ginst2511 (P1_R2358_U205, P1_R2358_U29, P1_R2358_U431, P1_R2358_U432);
  nand ginst2512 (P1_R2358_U206, P1_R2358_U427, P1_U2649);
  nand ginst2513 (P1_R2358_U207, P1_R2358_U424, P1_U2648);
  nand ginst2514 (P1_R2358_U208, P1_R2358_U31, P1_R2358_U433, P1_R2358_U434);
  nand ginst2515 (P1_R2358_U209, P1_R2358_U430, P1_U2650);
  and ginst2516 (P1_R2358_U21, P1_R2358_U240, P1_R2358_U242);
  nand ginst2517 (P1_R2358_U210, P1_R2358_U209, P1_R2358_U23);
  nand ginst2518 (P1_R2358_U211, P1_R2358_U120, P1_R2358_U210);
  nand ginst2519 (P1_R2358_U212, P1_R2358_U206, P1_R2358_U207, P1_R2358_U211);
  nand ginst2520 (P1_R2358_U213, P1_R2358_U121, P1_R2358_U212);
  not ginst2521 (P1_R2358_U214, P1_R2358_U156);
  nand ginst2522 (P1_R2358_U215, P1_R2358_U408, P1_U2644);
  nand ginst2523 (P1_R2358_U216, P1_R2358_U421, P1_U2643);
  nand ginst2524 (P1_R2358_U217, P1_R2358_U24, P1_R2358_U404, P1_R2358_U405);
  nand ginst2525 (P1_R2358_U218, P1_R2358_U25, P1_R2358_U417, P1_R2358_U418);
  nand ginst2526 (P1_R2358_U219, P1_R2358_U26, P1_R2358_U409, P1_R2358_U410);
  and ginst2527 (P1_R2358_U22, P1_R2358_U136, P1_R2358_U565, P1_R2358_U566);
  nand ginst2528 (P1_R2358_U220, P1_R2358_U416, P1_U2645);
  not ginst2529 (P1_R2358_U221, P1_R2358_U28);
  nand ginst2530 (P1_R2358_U222, P1_R2358_U219, P1_R2358_U221);
  nand ginst2531 (P1_R2358_U223, P1_R2358_U215, P1_R2358_U220, P1_R2358_U222);
  nand ginst2532 (P1_R2358_U224, P1_R2358_U217, P1_R2358_U218, P1_R2358_U223);
  nand ginst2533 (P1_R2358_U225, P1_R2358_U27, P1_R2358_U442, P1_R2358_U443);
  nand ginst2534 (P1_R2358_U226, P1_R2358_U156, P1_R2358_U217, P1_R2358_U218, P1_R2358_U219, P1_R2358_U225);
  not ginst2535 (P1_R2358_U227, P1_R2358_U154);
  nand ginst2536 (P1_R2358_U228, P1_R2358_U448, P1_U2642);
  nand ginst2537 (P1_R2358_U229, P1_R2358_U33, P1_R2358_U444, P1_R2358_U445);
  not ginst2538 (P1_R2358_U23, P1_U2352);
  nand ginst2539 (P1_R2358_U230, P1_R2358_U154, P1_R2358_U229);
  not ginst2540 (P1_R2358_U231, P1_R2358_U153);
  not ginst2541 (P1_R2358_U232, P1_R2358_U54);
  nand ginst2542 (P1_R2358_U233, P1_R2358_U403, P1_U2641);
  nand ginst2543 (P1_R2358_U234, P1_R2358_U156, P1_R2358_U225);
  not ginst2544 (P1_R2358_U235, P1_R2358_U155);
  nand ginst2545 (P1_R2358_U236, P1_R2358_U155, P1_R2358_U219);
  not ginst2546 (P1_R2358_U237, P1_R2358_U35);
  not ginst2547 (P1_R2358_U238, P1_R2358_U36);
  nand ginst2548 (P1_R2358_U239, P1_R2358_U215, P1_R2358_U36);
  not ginst2549 (P1_R2358_U24, P1_U2643);
  nand ginst2550 (P1_R2358_U240, P1_R2358_U122, P1_R2358_U239);
  nand ginst2551 (P1_R2358_U241, P1_R2358_U216, P1_R2358_U217);
  nand ginst2552 (P1_R2358_U242, P1_R2358_U215, P1_R2358_U241, P1_R2358_U36);
  nand ginst2553 (P1_R2358_U243, P1_R2358_U215, P1_R2358_U218);
  nand ginst2554 (P1_R2358_U244, P1_R2358_U237, P1_R2358_U243);
  nand ginst2555 (P1_R2358_U245, P1_R2358_U215, P1_R2358_U238);
  nand ginst2556 (P1_R2358_U246, P1_R2358_U208, P1_U2352);
  not ginst2557 (P1_R2358_U247, P1_R2358_U193);
  nand ginst2558 (P1_R2358_U248, P1_R2358_U193, P1_R2358_U205);
  not ginst2559 (P1_R2358_U249, P1_R2358_U65);
  not ginst2560 (P1_R2358_U25, P1_U2644);
  not ginst2561 (P1_R2358_U250, P1_R2358_U66);
  nand ginst2562 (P1_R2358_U251, P1_R2358_U207, P1_R2358_U66);
  nand ginst2563 (P1_R2358_U252, P1_R2358_U123, P1_R2358_U251);
  nand ginst2564 (P1_R2358_U253, P1_R2358_U203, P1_R2358_U204);
  nand ginst2565 (P1_R2358_U254, P1_R2358_U207, P1_R2358_U253, P1_R2358_U66);
  nand ginst2566 (P1_R2358_U255, P1_R2358_U459, P1_R2358_U460, P1_R2358_U60);
  nand ginst2567 (P1_R2358_U256, P1_R2358_U474, P1_U2635);
  nand ginst2568 (P1_R2358_U257, P1_R2358_U11, P1_R2358_U55);
  nand ginst2569 (P1_R2358_U258, P1_R2358_U467, P1_R2358_U468, P1_R2358_U58);
  nand ginst2570 (P1_R2358_U259, P1_R2358_U485, P1_R2358_U486, P1_R2358_U56);
  not ginst2571 (P1_R2358_U26, P1_U2645);
  not ginst2572 (P1_R2358_U260, P1_R2358_U59);
  not ginst2573 (P1_R2358_U261, P1_R2358_U61);
  nand ginst2574 (P1_R2358_U262, P1_R2358_U475, P1_R2358_U476, P1_R2358_U53);
  nand ginst2575 (P1_R2358_U263, P1_R2358_U479, P1_U2640);
  nand ginst2576 (P1_R2358_U264, P1_R2358_U484, P1_U2639);
  nand ginst2577 (P1_R2358_U265, P1_R2358_U12, P1_R2358_U52);
  nand ginst2578 (P1_R2358_U266, P1_R2358_U228, P1_R2358_U233, P1_R2358_U263);
  nand ginst2579 (P1_R2358_U267, P1_R2358_U262, P1_R2358_U266, P1_R2358_U357, P1_R2358_U360);
  nand ginst2580 (P1_R2358_U268, P1_R2358_U124, P1_R2358_U125, P1_R2358_U154);
  not ginst2581 (P1_R2358_U269, P1_R2358_U199);
  not ginst2582 (P1_R2358_U27, P1_U2646);
  not ginst2583 (P1_R2358_U270, P1_R2358_U57);
  not ginst2584 (P1_R2358_U271, P1_R2358_U197);
  nand ginst2585 (P1_R2358_U272, P1_R2358_U487, P1_R2358_U488, P1_R2358_U50);
  not ginst2586 (P1_R2358_U273, P1_R2358_U51);
  nand ginst2587 (P1_R2358_U274, P1_R2358_U489, P1_R2358_U49, P1_R2358_U490);
  nand ginst2588 (P1_R2358_U275, P1_R2358_U498, P1_U2633);
  nand ginst2589 (P1_R2358_U276, P1_R2358_U48, P1_R2358_U491, P1_R2358_U492);
  nand ginst2590 (P1_R2358_U277, P1_R2358_U495, P1_U2632);
  nand ginst2591 (P1_R2358_U278, P1_R2358_U46, P1_R2358_U506, P1_R2358_U507);
  not ginst2592 (P1_R2358_U279, P1_R2358_U47);
  nand ginst2593 (P1_R2358_U28, P1_R2358_U413, P1_U2646);
  nand ginst2594 (P1_R2358_U280, P1_R2358_U45, P1_R2358_U508, P1_R2358_U509);
  nand ginst2595 (P1_R2358_U281, P1_R2358_U518, P1_U2630);
  nand ginst2596 (P1_R2358_U282, P1_R2358_U44, P1_R2358_U504, P1_R2358_U505);
  nand ginst2597 (P1_R2358_U283, P1_R2358_U515, P1_U2629);
  nand ginst2598 (P1_R2358_U284, P1_R2358_U43, P1_R2358_U502, P1_R2358_U503);
  nand ginst2599 (P1_R2358_U285, P1_R2358_U512, P1_U2628);
  nand ginst2600 (P1_R2358_U286, P1_R2358_U41, P1_R2358_U528, P1_R2358_U529);
  not ginst2601 (P1_R2358_U287, P1_R2358_U42);
  nand ginst2602 (P1_R2358_U288, P1_R2358_U40, P1_R2358_U530, P1_R2358_U531);
  nand ginst2603 (P1_R2358_U289, P1_R2358_U543, P1_U2626);
  not ginst2604 (P1_R2358_U29, P1_U2649);
  nand ginst2605 (P1_R2358_U290, P1_R2358_U39, P1_R2358_U526, P1_R2358_U527);
  nand ginst2606 (P1_R2358_U291, P1_R2358_U540, P1_U2625);
  nand ginst2607 (P1_R2358_U292, P1_R2358_U38, P1_R2358_U524, P1_R2358_U525);
  nand ginst2608 (P1_R2358_U293, P1_R2358_U537, P1_U2624);
  nand ginst2609 (P1_R2358_U294, P1_R2358_U37, P1_R2358_U522, P1_R2358_U523);
  nand ginst2610 (P1_R2358_U295, P1_R2358_U534, P1_U2623);
  nand ginst2611 (P1_R2358_U296, P1_R2358_U547, P1_R2358_U548, P1_R2358_U62);
  nand ginst2612 (P1_R2358_U297, P1_R2358_U551, P1_U2622);
  nand ginst2613 (P1_R2358_U298, P1_R2358_U184, P1_R2358_U296);
  not ginst2614 (P1_R2358_U299, P1_R2358_U183);
  not ginst2615 (P1_R2358_U30, P1_U2648);
  nand ginst2616 (P1_R2358_U300, P1_R2358_U552, P1_R2358_U553, P1_R2358_U64);
  not ginst2617 (P1_R2358_U301, P1_R2358_U179);
  nand ginst2618 (P1_R2358_U302, P1_R2358_U183, P1_R2358_U300);
  not ginst2619 (P1_R2358_U303, P1_R2358_U182);
  nand ginst2620 (P1_R2358_U304, P1_R2358_U75, P1_U2620);
  nand ginst2621 (P1_R2358_U305, P1_R2358_U558, P1_R2358_U63);
  nand ginst2622 (P1_R2358_U306, P1_R2358_U202, P1_R2358_U207);
  nand ginst2623 (P1_R2358_U307, P1_R2358_U249, P1_R2358_U306);
  nand ginst2624 (P1_R2358_U308, P1_R2358_U207, P1_R2358_U250);
  nand ginst2625 (P1_R2358_U309, P1_R2358_U199, P1_R2358_U259);
  not ginst2626 (P1_R2358_U31, P1_U2650);
  not ginst2627 (P1_R2358_U310, P1_R2358_U198);
  nand ginst2628 (P1_R2358_U311, P1_R2358_U198, P1_R2358_U258);
  not ginst2629 (P1_R2358_U312, P1_R2358_U71);
  not ginst2630 (P1_R2358_U313, P1_R2358_U72);
  nand ginst2631 (P1_R2358_U314, P1_R2358_U61, P1_R2358_U72);
  nand ginst2632 (P1_R2358_U315, P1_R2358_U139, P1_R2358_U314);
  nand ginst2633 (P1_R2358_U316, P1_R2358_U256, P1_R2358_U257);
  nand ginst2634 (P1_R2358_U317, P1_R2358_U140, P1_R2358_U72);
  nand ginst2635 (P1_R2358_U318, P1_R2358_U255, P1_R2358_U61);
  nand ginst2636 (P1_R2358_U319, P1_R2358_U312, P1_R2358_U318);
  not ginst2637 (P1_R2358_U32, P1_U2647);
  nand ginst2638 (P1_R2358_U320, P1_R2358_U313, P1_R2358_U61);
  nand ginst2639 (P1_R2358_U321, P1_R2358_U153, P1_R2358_U54);
  not ginst2640 (P1_R2358_U322, P1_R2358_U73);
  not ginst2641 (P1_R2358_U323, P1_R2358_U74);
  nand ginst2642 (P1_R2358_U324, P1_R2358_U263, P1_R2358_U74);
  nand ginst2643 (P1_R2358_U325, P1_R2358_U141, P1_R2358_U324);
  nand ginst2644 (P1_R2358_U326, P1_R2358_U264, P1_R2358_U265);
  nand ginst2645 (P1_R2358_U327, P1_R2358_U142, P1_R2358_U74);
  nand ginst2646 (P1_R2358_U328, P1_R2358_U262, P1_R2358_U263);
  nand ginst2647 (P1_R2358_U329, P1_R2358_U322, P1_R2358_U328);
  not ginst2648 (P1_R2358_U33, P1_U2642);
  nand ginst2649 (P1_R2358_U330, P1_R2358_U263, P1_R2358_U323);
  not ginst2650 (P1_R2358_U331, P1_R2358_U200);
  nand ginst2651 (P1_R2358_U332, P1_R2358_U233, P1_R2358_U54);
  nand ginst2652 (P1_R2358_U333, P1_R2358_U228, P1_R2358_U229);
  nand ginst2653 (P1_R2358_U334, P1_R2358_U219, P1_R2358_U220);
  nand ginst2654 (P1_R2358_U335, P1_R2358_U225, P1_R2358_U28);
  nand ginst2655 (P1_R2358_U336, P1_R2358_U179, P1_R2358_U300);
  nand ginst2656 (P1_R2358_U337, P1_R2358_U296, P1_R2358_U297);
  nand ginst2657 (P1_R2358_U338, P1_R2358_U294, P1_R2358_U295);
  nand ginst2658 (P1_R2358_U339, P1_R2358_U292, P1_R2358_U293);
  not ginst2659 (P1_R2358_U34, P1_U2641);
  nand ginst2660 (P1_R2358_U340, P1_R2358_U290, P1_R2358_U291);
  nand ginst2661 (P1_R2358_U341, P1_R2358_U288, P1_R2358_U289);
  nand ginst2662 (P1_R2358_U342, P1_R2358_U286, P1_R2358_U42);
  nand ginst2663 (P1_R2358_U343, P1_R2358_U284, P1_R2358_U285);
  nand ginst2664 (P1_R2358_U344, P1_R2358_U282, P1_R2358_U283);
  nand ginst2665 (P1_R2358_U345, P1_R2358_U280, P1_R2358_U281);
  nand ginst2666 (P1_R2358_U346, P1_R2358_U205, P1_R2358_U206);
  nand ginst2667 (P1_R2358_U347, P1_R2358_U278, P1_R2358_U47);
  nand ginst2668 (P1_R2358_U348, P1_R2358_U276, P1_R2358_U277);
  nand ginst2669 (P1_R2358_U349, P1_R2358_U274, P1_R2358_U275);
  nand ginst2670 (P1_R2358_U35, P1_R2358_U220, P1_R2358_U236);
  nand ginst2671 (P1_R2358_U350, P1_R2358_U272, P1_R2358_U51);
  nand ginst2672 (P1_R2358_U351, P1_R2358_U258, P1_R2358_U59);
  nand ginst2673 (P1_R2358_U352, P1_R2358_U259, P1_R2358_U57);
  nand ginst2674 (P1_R2358_U353, P1_R2358_U255, P1_R2358_U257, P1_R2358_U258, P1_R2358_U270);
  nand ginst2675 (P1_R2358_U354, P1_R2358_U255, P1_R2358_U257, P1_R2358_U260);
  nand ginst2676 (P1_R2358_U355, P1_R2358_U257, P1_R2358_U261);
  nand ginst2677 (P1_R2358_U356, P1_R2358_U11, P1_R2358_U55);
  nand ginst2678 (P1_R2358_U357, P1_R2358_U232, P1_R2358_U263);
  nand ginst2679 (P1_R2358_U358, P1_R2358_U273, P1_R2358_U274);
  not ginst2680 (P1_R2358_U359, P1_R2358_U70);
  nand ginst2681 (P1_R2358_U36, P1_R2358_U218, P1_R2358_U35);
  nand ginst2682 (P1_R2358_U360, P1_R2358_U12, P1_R2358_U52);
  nand ginst2683 (P1_R2358_U361, P1_R2358_U276, P1_R2358_U70);
  nand ginst2684 (P1_R2358_U362, P1_R2358_U279, P1_R2358_U280);
  nand ginst2685 (P1_R2358_U363, P1_R2358_U281, P1_R2358_U362);
  nand ginst2686 (P1_R2358_U364, P1_R2358_U282, P1_R2358_U363);
  not ginst2687 (P1_R2358_U365, P1_R2358_U69);
  nand ginst2688 (P1_R2358_U366, P1_R2358_U284, P1_R2358_U69);
  nand ginst2689 (P1_R2358_U367, P1_R2358_U287, P1_R2358_U288);
  nand ginst2690 (P1_R2358_U368, P1_R2358_U289, P1_R2358_U367);
  nand ginst2691 (P1_R2358_U369, P1_R2358_U290, P1_R2358_U368);
  not ginst2692 (P1_R2358_U37, P1_U2623);
  not ginst2693 (P1_R2358_U370, P1_R2358_U68);
  nand ginst2694 (P1_R2358_U371, P1_R2358_U292, P1_R2358_U68);
  not ginst2695 (P1_R2358_U372, P1_R2358_U67);
  nand ginst2696 (P1_R2358_U373, P1_R2358_U294, P1_R2358_U67);
  nand ginst2697 (P1_R2358_U374, P1_R2358_U134, P1_R2358_U183, P1_R2358_U300);
  nand ginst2698 (P1_R2358_U375, P1_R2358_U189, P1_R2358_U286);
  not ginst2699 (P1_R2358_U376, P1_R2358_U188);
  nand ginst2700 (P1_R2358_U377, P1_R2358_U189, P1_R2358_U8);
  not ginst2701 (P1_R2358_U378, P1_R2358_U187);
  nand ginst2702 (P1_R2358_U379, P1_R2358_U189, P1_R2358_U9);
  not ginst2703 (P1_R2358_U38, P1_U2624);
  not ginst2704 (P1_R2358_U380, P1_R2358_U186);
  nand ginst2705 (P1_R2358_U381, P1_R2358_U10, P1_R2358_U189);
  not ginst2706 (P1_R2358_U382, P1_R2358_U185);
  nand ginst2707 (P1_R2358_U383, P1_R2358_U132, P1_R2358_U189);
  not ginst2708 (P1_R2358_U384, P1_R2358_U184);
  nand ginst2709 (P1_R2358_U385, P1_R2358_U130, P1_R2358_U194);
  not ginst2710 (P1_R2358_U386, P1_R2358_U189);
  nand ginst2711 (P1_R2358_U387, P1_R2358_U194, P1_R2358_U7);
  not ginst2712 (P1_R2358_U388, P1_R2358_U190);
  nand ginst2713 (P1_R2358_U389, P1_R2358_U194, P1_R2358_U6);
  not ginst2714 (P1_R2358_U39, P1_U2625);
  not ginst2715 (P1_R2358_U390, P1_R2358_U191);
  nand ginst2716 (P1_R2358_U391, P1_R2358_U194, P1_R2358_U278);
  not ginst2717 (P1_R2358_U392, P1_R2358_U192);
  nand ginst2718 (P1_R2358_U393, P1_R2358_U128, P1_R2358_U197);
  not ginst2719 (P1_R2358_U394, P1_R2358_U194);
  nand ginst2720 (P1_R2358_U395, P1_R2358_U197, P1_R2358_U5);
  not ginst2721 (P1_R2358_U396, P1_R2358_U195);
  nand ginst2722 (P1_R2358_U397, P1_R2358_U197, P1_R2358_U272);
  not ginst2723 (P1_R2358_U398, P1_R2358_U196);
  nand ginst2724 (P1_R2358_U399, P1_R2358_U143, P1_U2352);
  not ginst2725 (P1_R2358_U40, P1_U2626);
  nand ginst2726 (P1_R2358_U400, P1_R2358_U23, P1_U2618);
  nand ginst2727 (P1_R2358_U401, P1_R2358_U143, P1_U2352);
  nand ginst2728 (P1_R2358_U402, P1_R2358_U23, P1_U2618);
  nand ginst2729 (P1_R2358_U403, P1_R2358_U401, P1_R2358_U402);
  nand ginst2730 (P1_R2358_U404, P1_R2358_U144, P1_U2352);
  nand ginst2731 (P1_R2358_U405, P1_R2358_U23, P1_U2615);
  nand ginst2732 (P1_R2358_U406, P1_R2358_U145, P1_U2352);
  nand ginst2733 (P1_R2358_U407, P1_R2358_U23, P1_U2614);
  nand ginst2734 (P1_R2358_U408, P1_R2358_U406, P1_R2358_U407);
  nand ginst2735 (P1_R2358_U409, P1_R2358_U146, P1_U2352);
  not ginst2736 (P1_R2358_U41, P1_U2627);
  nand ginst2737 (P1_R2358_U410, P1_R2358_U23, P1_U2667);
  nand ginst2738 (P1_R2358_U411, P1_R2358_U147, P1_U2352);
  nand ginst2739 (P1_R2358_U412, P1_R2358_U23, P1_U2668);
  nand ginst2740 (P1_R2358_U413, P1_R2358_U411, P1_R2358_U412);
  nand ginst2741 (P1_R2358_U414, P1_R2358_U146, P1_U2352);
  nand ginst2742 (P1_R2358_U415, P1_R2358_U23, P1_U2667);
  nand ginst2743 (P1_R2358_U416, P1_R2358_U414, P1_R2358_U415);
  nand ginst2744 (P1_R2358_U417, P1_R2358_U145, P1_U2352);
  nand ginst2745 (P1_R2358_U418, P1_R2358_U23, P1_U2614);
  nand ginst2746 (P1_R2358_U419, P1_R2358_U144, P1_U2352);
  nand ginst2747 (P1_R2358_U42, P1_R2358_U546, P1_U2627);
  nand ginst2748 (P1_R2358_U420, P1_R2358_U23, P1_U2615);
  nand ginst2749 (P1_R2358_U421, P1_R2358_U419, P1_R2358_U420);
  nand ginst2750 (P1_R2358_U422, P1_R2358_U148, P1_U2352);
  nand ginst2751 (P1_R2358_U423, P1_R2358_U23, P1_U2670);
  nand ginst2752 (P1_R2358_U424, P1_R2358_U422, P1_R2358_U423);
  nand ginst2753 (P1_R2358_U425, P1_R2358_U149, P1_U2352);
  nand ginst2754 (P1_R2358_U426, P1_R2358_U23, P1_U2671);
  nand ginst2755 (P1_R2358_U427, P1_R2358_U425, P1_R2358_U426);
  nand ginst2756 (P1_R2358_U428, P1_R2358_U150, P1_U2352);
  nand ginst2757 (P1_R2358_U429, P1_R2358_U23, P1_U2672);
  not ginst2758 (P1_R2358_U43, P1_U2628);
  nand ginst2759 (P1_R2358_U430, P1_R2358_U428, P1_R2358_U429);
  nand ginst2760 (P1_R2358_U431, P1_R2358_U149, P1_U2352);
  nand ginst2761 (P1_R2358_U432, P1_R2358_U23, P1_U2671);
  nand ginst2762 (P1_R2358_U433, P1_R2358_U150, P1_U2352);
  nand ginst2763 (P1_R2358_U434, P1_R2358_U23, P1_U2672);
  nand ginst2764 (P1_R2358_U435, P1_R2358_U148, P1_U2352);
  nand ginst2765 (P1_R2358_U436, P1_R2358_U23, P1_U2670);
  nand ginst2766 (P1_R2358_U437, P1_R2358_U151, P1_U2352);
  nand ginst2767 (P1_R2358_U438, P1_R2358_U23, P1_U2669);
  nand ginst2768 (P1_R2358_U439, P1_R2358_U151, P1_U2352);
  not ginst2769 (P1_R2358_U44, P1_U2629);
  nand ginst2770 (P1_R2358_U440, P1_R2358_U23, P1_U2669);
  nand ginst2771 (P1_R2358_U441, P1_R2358_U439, P1_R2358_U440);
  nand ginst2772 (P1_R2358_U442, P1_R2358_U147, P1_U2352);
  nand ginst2773 (P1_R2358_U443, P1_R2358_U23, P1_U2668);
  nand ginst2774 (P1_R2358_U444, P1_R2358_U152, P1_U2352);
  nand ginst2775 (P1_R2358_U445, P1_R2358_U23, P1_U2617);
  nand ginst2776 (P1_R2358_U446, P1_R2358_U152, P1_U2352);
  nand ginst2777 (P1_R2358_U447, P1_R2358_U23, P1_U2617);
  nand ginst2778 (P1_R2358_U448, P1_R2358_U446, P1_R2358_U447);
  nand ginst2779 (P1_R2358_U449, P1_R2358_U153, P1_R2358_U332);
  not ginst2780 (P1_R2358_U45, P1_U2630);
  nand ginst2781 (P1_R2358_U450, P1_R2358_U231, P1_R2358_U77);
  nand ginst2782 (P1_R2358_U451, P1_R2358_U154, P1_R2358_U333);
  nand ginst2783 (P1_R2358_U452, P1_R2358_U227, P1_R2358_U79);
  nand ginst2784 (P1_R2358_U453, P1_R2358_U155, P1_R2358_U334);
  nand ginst2785 (P1_R2358_U454, P1_R2358_U235, P1_R2358_U81);
  nand ginst2786 (P1_R2358_U455, P1_R2358_U156, P1_R2358_U335);
  nand ginst2787 (P1_R2358_U456, P1_R2358_U214, P1_R2358_U83);
  nand ginst2788 (P1_R2358_U457, P1_R2358_U157, P1_U2352);
  nand ginst2789 (P1_R2358_U458, P1_R2358_U23, P1_U2611);
  nand ginst2790 (P1_R2358_U459, P1_R2358_U158, P1_U2352);
  not ginst2791 (P1_R2358_U46, P1_U2631);
  nand ginst2792 (P1_R2358_U460, P1_R2358_U23, P1_U2612);
  nand ginst2793 (P1_R2358_U461, P1_R2358_U159, P1_U2352);
  nand ginst2794 (P1_R2358_U462, P1_R2358_U23, P1_U2613);
  nand ginst2795 (P1_R2358_U463, P1_R2358_U461, P1_R2358_U462);
  nand ginst2796 (P1_R2358_U464, P1_R2358_U158, P1_U2352);
  nand ginst2797 (P1_R2358_U465, P1_R2358_U23, P1_U2612);
  nand ginst2798 (P1_R2358_U466, P1_R2358_U464, P1_R2358_U465);
  nand ginst2799 (P1_R2358_U467, P1_R2358_U159, P1_U2352);
  nand ginst2800 (P1_R2358_U468, P1_R2358_U23, P1_U2613);
  nand ginst2801 (P1_R2358_U469, P1_R2358_U160, P1_U2352);
  nand ginst2802 (P1_R2358_U47, P1_R2358_U521, P1_U2631);
  nand ginst2803 (P1_R2358_U470, P1_R2358_U23, P1_U2616);
  nand ginst2804 (P1_R2358_U471, P1_R2358_U469, P1_R2358_U470);
  nand ginst2805 (P1_R2358_U472, P1_R2358_U157, P1_U2352);
  nand ginst2806 (P1_R2358_U473, P1_R2358_U23, P1_U2611);
  nand ginst2807 (P1_R2358_U474, P1_R2358_U472, P1_R2358_U473);
  nand ginst2808 (P1_R2358_U475, P1_R2358_U161, P1_U2352);
  nand ginst2809 (P1_R2358_U476, P1_R2358_U23, P1_U2610);
  nand ginst2810 (P1_R2358_U477, P1_R2358_U161, P1_U2352);
  nand ginst2811 (P1_R2358_U478, P1_R2358_U23, P1_U2610);
  nand ginst2812 (P1_R2358_U479, P1_R2358_U477, P1_R2358_U478);
  not ginst2813 (P1_R2358_U48, P1_U2632);
  nand ginst2814 (P1_R2358_U480, P1_R2358_U162, P1_U2352);
  nand ginst2815 (P1_R2358_U481, P1_R2358_U23, P1_U2609);
  nand ginst2816 (P1_R2358_U482, P1_R2358_U162, P1_U2352);
  nand ginst2817 (P1_R2358_U483, P1_R2358_U23, P1_U2609);
  nand ginst2818 (P1_R2358_U484, P1_R2358_U482, P1_R2358_U483);
  nand ginst2819 (P1_R2358_U485, P1_R2358_U160, P1_U2352);
  nand ginst2820 (P1_R2358_U486, P1_R2358_U23, P1_U2616);
  nand ginst2821 (P1_R2358_U487, P1_R2358_U163, P1_U2352);
  nand ginst2822 (P1_R2358_U488, P1_R2358_U23, P1_U2666);
  nand ginst2823 (P1_R2358_U489, P1_R2358_U164, P1_U2352);
  not ginst2824 (P1_R2358_U49, P1_U2633);
  nand ginst2825 (P1_R2358_U490, P1_R2358_U23, P1_U2665);
  nand ginst2826 (P1_R2358_U491, P1_R2358_U165, P1_U2352);
  nand ginst2827 (P1_R2358_U492, P1_R2358_U23, P1_U2664);
  nand ginst2828 (P1_R2358_U493, P1_R2358_U165, P1_U2352);
  nand ginst2829 (P1_R2358_U494, P1_R2358_U23, P1_U2664);
  nand ginst2830 (P1_R2358_U495, P1_R2358_U493, P1_R2358_U494);
  nand ginst2831 (P1_R2358_U496, P1_R2358_U164, P1_U2352);
  nand ginst2832 (P1_R2358_U497, P1_R2358_U23, P1_U2665);
  nand ginst2833 (P1_R2358_U498, P1_R2358_U496, P1_R2358_U497);
  nand ginst2834 (P1_R2358_U499, P1_R2358_U163, P1_U2352);
  and ginst2835 (P1_R2358_U5, P1_R2358_U272, P1_R2358_U274);
  not ginst2836 (P1_R2358_U50, P1_U2634);
  nand ginst2837 (P1_R2358_U500, P1_R2358_U23, P1_U2666);
  nand ginst2838 (P1_R2358_U501, P1_R2358_U499, P1_R2358_U500);
  nand ginst2839 (P1_R2358_U502, P1_R2358_U166, P1_U2352);
  nand ginst2840 (P1_R2358_U503, P1_R2358_U23, P1_U2660);
  nand ginst2841 (P1_R2358_U504, P1_R2358_U167, P1_U2352);
  nand ginst2842 (P1_R2358_U505, P1_R2358_U23, P1_U2661);
  nand ginst2843 (P1_R2358_U506, P1_R2358_U168, P1_U2352);
  nand ginst2844 (P1_R2358_U507, P1_R2358_U23, P1_U2663);
  nand ginst2845 (P1_R2358_U508, P1_R2358_U169, P1_U2352);
  nand ginst2846 (P1_R2358_U509, P1_R2358_U23, P1_U2662);
  nand ginst2847 (P1_R2358_U51, P1_R2358_U501, P1_U2634);
  nand ginst2848 (P1_R2358_U510, P1_R2358_U166, P1_U2352);
  nand ginst2849 (P1_R2358_U511, P1_R2358_U23, P1_U2660);
  nand ginst2850 (P1_R2358_U512, P1_R2358_U510, P1_R2358_U511);
  nand ginst2851 (P1_R2358_U513, P1_R2358_U167, P1_U2352);
  nand ginst2852 (P1_R2358_U514, P1_R2358_U23, P1_U2661);
  nand ginst2853 (P1_R2358_U515, P1_R2358_U513, P1_R2358_U514);
  nand ginst2854 (P1_R2358_U516, P1_R2358_U169, P1_U2352);
  nand ginst2855 (P1_R2358_U517, P1_R2358_U23, P1_U2662);
  nand ginst2856 (P1_R2358_U518, P1_R2358_U516, P1_R2358_U517);
  nand ginst2857 (P1_R2358_U519, P1_R2358_U168, P1_U2352);
  not ginst2858 (P1_R2358_U52, P1_U2639);
  nand ginst2859 (P1_R2358_U520, P1_R2358_U23, P1_U2663);
  nand ginst2860 (P1_R2358_U521, P1_R2358_U519, P1_R2358_U520);
  nand ginst2861 (P1_R2358_U522, P1_R2358_U170, P1_U2352);
  nand ginst2862 (P1_R2358_U523, P1_R2358_U23, P1_U2655);
  nand ginst2863 (P1_R2358_U524, P1_R2358_U171, P1_U2352);
  nand ginst2864 (P1_R2358_U525, P1_R2358_U23, P1_U2656);
  nand ginst2865 (P1_R2358_U526, P1_R2358_U172, P1_U2352);
  nand ginst2866 (P1_R2358_U527, P1_R2358_U23, P1_U2657);
  nand ginst2867 (P1_R2358_U528, P1_R2358_U173, P1_U2352);
  nand ginst2868 (P1_R2358_U529, P1_R2358_U23, P1_U2659);
  not ginst2869 (P1_R2358_U53, P1_U2640);
  nand ginst2870 (P1_R2358_U530, P1_R2358_U174, P1_U2352);
  nand ginst2871 (P1_R2358_U531, P1_R2358_U23, P1_U2658);
  nand ginst2872 (P1_R2358_U532, P1_R2358_U170, P1_U2352);
  nand ginst2873 (P1_R2358_U533, P1_R2358_U23, P1_U2655);
  nand ginst2874 (P1_R2358_U534, P1_R2358_U532, P1_R2358_U533);
  nand ginst2875 (P1_R2358_U535, P1_R2358_U171, P1_U2352);
  nand ginst2876 (P1_R2358_U536, P1_R2358_U23, P1_U2656);
  nand ginst2877 (P1_R2358_U537, P1_R2358_U535, P1_R2358_U536);
  nand ginst2878 (P1_R2358_U538, P1_R2358_U172, P1_U2352);
  nand ginst2879 (P1_R2358_U539, P1_R2358_U23, P1_U2657);
  nand ginst2880 (P1_R2358_U54, P1_R2358_U34, P1_R2358_U399, P1_R2358_U400);
  nand ginst2881 (P1_R2358_U540, P1_R2358_U538, P1_R2358_U539);
  nand ginst2882 (P1_R2358_U541, P1_R2358_U174, P1_U2352);
  nand ginst2883 (P1_R2358_U542, P1_R2358_U23, P1_U2658);
  nand ginst2884 (P1_R2358_U543, P1_R2358_U541, P1_R2358_U542);
  nand ginst2885 (P1_R2358_U544, P1_R2358_U173, P1_U2352);
  nand ginst2886 (P1_R2358_U545, P1_R2358_U23, P1_U2659);
  nand ginst2887 (P1_R2358_U546, P1_R2358_U544, P1_R2358_U545);
  nand ginst2888 (P1_R2358_U547, P1_R2358_U175, P1_U2352);
  nand ginst2889 (P1_R2358_U548, P1_R2358_U23, P1_U2654);
  nand ginst2890 (P1_R2358_U549, P1_R2358_U175, P1_U2352);
  not ginst2891 (P1_R2358_U55, P1_U2635);
  nand ginst2892 (P1_R2358_U550, P1_R2358_U23, P1_U2654);
  nand ginst2893 (P1_R2358_U551, P1_R2358_U549, P1_R2358_U550);
  nand ginst2894 (P1_R2358_U552, P1_R2358_U176, P1_U2352);
  nand ginst2895 (P1_R2358_U553, P1_R2358_U23, P1_U2653);
  nand ginst2896 (P1_R2358_U554, P1_R2358_U177, P1_U2352);
  nand ginst2897 (P1_R2358_U555, P1_R2358_U23, P1_U2651);
  nand ginst2898 (P1_R2358_U556, P1_R2358_U178, P1_U2352);
  nand ginst2899 (P1_R2358_U557, P1_R2358_U23, P1_U2652);
  not ginst2900 (P1_R2358_U558, P1_R2358_U75);
  nand ginst2901 (P1_R2358_U559, P1_R2358_U177, P1_U2352);
  not ginst2902 (P1_R2358_U56, P1_U2638);
  nand ginst2903 (P1_R2358_U560, P1_R2358_U23, P1_U2651);
  nand ginst2904 (P1_R2358_U561, P1_R2358_U559, P1_R2358_U560);
  nand ginst2905 (P1_R2358_U562, P1_R2358_U176, P1_U2352);
  nand ginst2906 (P1_R2358_U563, P1_R2358_U23, P1_U2653);
  nand ginst2907 (P1_R2358_U564, P1_R2358_U562, P1_R2358_U563);
  nand ginst2908 (P1_R2358_U565, P1_R2358_U135, P1_R2358_U179, P1_R2358_U302);
  nand ginst2909 (P1_R2358_U566, P1_R2358_U301, P1_R2358_U305, P1_R2358_U561);
  nand ginst2910 (P1_R2358_U567, P1_R2358_U13, P1_R2358_U558, P1_R2358_U63);
  nand ginst2911 (P1_R2358_U568, P1_R2358_U561, P1_R2358_U75, P1_U2620);
  nand ginst2912 (P1_R2358_U569, P1_R2358_U558, P1_U2620);
  nand ginst2913 (P1_R2358_U57, P1_R2358_U471, P1_U2638);
  nand ginst2914 (P1_R2358_U570, P1_R2358_U63, P1_R2358_U75);
  nand ginst2915 (P1_R2358_U571, P1_R2358_U558, P1_U2620);
  nand ginst2916 (P1_R2358_U572, P1_R2358_U63, P1_R2358_U75);
  nand ginst2917 (P1_R2358_U573, P1_R2358_U571, P1_R2358_U572);
  nand ginst2918 (P1_R2358_U574, P1_R2358_U181, P1_R2358_U182);
  nand ginst2919 (P1_R2358_U575, P1_R2358_U303, P1_R2358_U573);
  nand ginst2920 (P1_R2358_U576, P1_R2358_U183, P1_R2358_U336);
  nand ginst2921 (P1_R2358_U577, P1_R2358_U299, P1_R2358_U86);
  nand ginst2922 (P1_R2358_U578, P1_R2358_U184, P1_R2358_U337);
  nand ginst2923 (P1_R2358_U579, P1_R2358_U384, P1_R2358_U88);
  not ginst2924 (P1_R2358_U58, P1_U2637);
  nand ginst2925 (P1_R2358_U580, P1_R2358_U185, P1_R2358_U338);
  nand ginst2926 (P1_R2358_U581, P1_R2358_U382, P1_R2358_U90);
  nand ginst2927 (P1_R2358_U582, P1_R2358_U186, P1_R2358_U339);
  nand ginst2928 (P1_R2358_U583, P1_R2358_U380, P1_R2358_U92);
  nand ginst2929 (P1_R2358_U584, P1_R2358_U187, P1_R2358_U340);
  nand ginst2930 (P1_R2358_U585, P1_R2358_U378, P1_R2358_U94);
  nand ginst2931 (P1_R2358_U586, P1_R2358_U188, P1_R2358_U341);
  nand ginst2932 (P1_R2358_U587, P1_R2358_U376, P1_R2358_U96);
  nand ginst2933 (P1_R2358_U588, P1_R2358_U189, P1_R2358_U342);
  nand ginst2934 (P1_R2358_U589, P1_R2358_U386, P1_R2358_U98);
  nand ginst2935 (P1_R2358_U59, P1_R2358_U463, P1_U2637);
  nand ginst2936 (P1_R2358_U590, P1_R2358_U190, P1_R2358_U343);
  nand ginst2937 (P1_R2358_U591, P1_R2358_U100, P1_R2358_U388);
  nand ginst2938 (P1_R2358_U592, P1_R2358_U191, P1_R2358_U344);
  nand ginst2939 (P1_R2358_U593, P1_R2358_U102, P1_R2358_U390);
  nand ginst2940 (P1_R2358_U594, P1_R2358_U192, P1_R2358_U345);
  nand ginst2941 (P1_R2358_U595, P1_R2358_U104, P1_R2358_U392);
  nand ginst2942 (P1_R2358_U596, P1_R2358_U193, P1_R2358_U346);
  nand ginst2943 (P1_R2358_U597, P1_R2358_U106, P1_R2358_U247);
  nand ginst2944 (P1_R2358_U598, P1_R2358_U194, P1_R2358_U347);
  nand ginst2945 (P1_R2358_U599, P1_R2358_U108, P1_R2358_U394);
  and ginst2946 (P1_R2358_U6, P1_R2358_U278, P1_R2358_U280);
  not ginst2947 (P1_R2358_U60, P1_U2636);
  nand ginst2948 (P1_R2358_U600, P1_R2358_U195, P1_R2358_U348);
  nand ginst2949 (P1_R2358_U601, P1_R2358_U110, P1_R2358_U396);
  nand ginst2950 (P1_R2358_U602, P1_R2358_U196, P1_R2358_U349);
  nand ginst2951 (P1_R2358_U603, P1_R2358_U112, P1_R2358_U398);
  nand ginst2952 (P1_R2358_U604, P1_R2358_U197, P1_R2358_U350);
  nand ginst2953 (P1_R2358_U605, P1_R2358_U114, P1_R2358_U271);
  nand ginst2954 (P1_R2358_U606, P1_R2358_U198, P1_R2358_U351);
  nand ginst2955 (P1_R2358_U607, P1_R2358_U116, P1_R2358_U310);
  nand ginst2956 (P1_R2358_U608, P1_R2358_U199, P1_R2358_U352);
  nand ginst2957 (P1_R2358_U609, P1_R2358_U118, P1_R2358_U269);
  nand ginst2958 (P1_R2358_U61, P1_R2358_U466, P1_U2636);
  nand ginst2959 (P1_R2358_U610, P1_R2358_U200, P1_U2352);
  nand ginst2960 (P1_R2358_U611, P1_R2358_U23, P1_R2358_U331);
  not ginst2961 (P1_R2358_U62, P1_U2622);
  not ginst2962 (P1_R2358_U63, P1_U2620);
  not ginst2963 (P1_R2358_U64, P1_U2621);
  nand ginst2964 (P1_R2358_U65, P1_R2358_U206, P1_R2358_U248);
  nand ginst2965 (P1_R2358_U66, P1_R2358_U202, P1_R2358_U65);
  nand ginst2966 (P1_R2358_U67, P1_R2358_U293, P1_R2358_U371);
  nand ginst2967 (P1_R2358_U68, P1_R2358_U291, P1_R2358_U369);
  nand ginst2968 (P1_R2358_U69, P1_R2358_U283, P1_R2358_U364);
  and ginst2969 (P1_R2358_U7, P1_R2358_U282, P1_R2358_U6);
  nand ginst2970 (P1_R2358_U70, P1_R2358_U275, P1_R2358_U358);
  nand ginst2971 (P1_R2358_U71, P1_R2358_U311, P1_R2358_U59);
  nand ginst2972 (P1_R2358_U72, P1_R2358_U255, P1_R2358_U71);
  nand ginst2973 (P1_R2358_U73, P1_R2358_U233, P1_R2358_U321);
  nand ginst2974 (P1_R2358_U74, P1_R2358_U262, P1_R2358_U73);
  nand ginst2975 (P1_R2358_U75, P1_R2358_U556, P1_R2358_U557);
  nand ginst2976 (P1_R2358_U76, P1_R2358_U610, P1_R2358_U611);
  and ginst2977 (P1_R2358_U77, P1_R2358_U233, P1_R2358_U54);
  nand ginst2978 (P1_R2358_U78, P1_R2358_U449, P1_R2358_U450);
  and ginst2979 (P1_R2358_U79, P1_R2358_U228, P1_R2358_U229);
  and ginst2980 (P1_R2358_U8, P1_R2358_U286, P1_R2358_U288);
  nand ginst2981 (P1_R2358_U80, P1_R2358_U451, P1_R2358_U452);
  and ginst2982 (P1_R2358_U81, P1_R2358_U219, P1_R2358_U220);
  nand ginst2983 (P1_R2358_U82, P1_R2358_U453, P1_R2358_U454);
  and ginst2984 (P1_R2358_U83, P1_R2358_U225, P1_R2358_U28);
  nand ginst2985 (P1_R2358_U84, P1_R2358_U455, P1_R2358_U456);
  nand ginst2986 (P1_R2358_U85, P1_R2358_U574, P1_R2358_U575);
  and ginst2987 (P1_R2358_U86, P1_R2358_U179, P1_R2358_U300);
  nand ginst2988 (P1_R2358_U87, P1_R2358_U576, P1_R2358_U577);
  and ginst2989 (P1_R2358_U88, P1_R2358_U296, P1_R2358_U297);
  nand ginst2990 (P1_R2358_U89, P1_R2358_U578, P1_R2358_U579);
  and ginst2991 (P1_R2358_U9, P1_R2358_U290, P1_R2358_U8);
  and ginst2992 (P1_R2358_U90, P1_R2358_U294, P1_R2358_U295);
  nand ginst2993 (P1_R2358_U91, P1_R2358_U580, P1_R2358_U581);
  and ginst2994 (P1_R2358_U92, P1_R2358_U292, P1_R2358_U293);
  nand ginst2995 (P1_R2358_U93, P1_R2358_U582, P1_R2358_U583);
  and ginst2996 (P1_R2358_U94, P1_R2358_U290, P1_R2358_U291);
  nand ginst2997 (P1_R2358_U95, P1_R2358_U584, P1_R2358_U585);
  and ginst2998 (P1_R2358_U96, P1_R2358_U288, P1_R2358_U289);
  nand ginst2999 (P1_R2358_U97, P1_R2358_U586, P1_R2358_U587);
  and ginst3000 (P1_R2358_U98, P1_R2358_U286, P1_R2358_U42);
  nand ginst3001 (P1_R2358_U99, P1_R2358_U588, P1_R2358_U589);
  not ginst3002 (P1_R584_U6, P1_U2676);
  not ginst3003 (P1_R584_U7, P1_U2677);
  not ginst3004 (P1_R584_U8, P1_U2674);
  not ginst3005 (P1_R584_U9, P1_U2675);
  not ginst3006 (P1_SUB_357_U10, P1_U3227);
  not ginst3007 (P1_SUB_357_U11, P1_U3230);
  not ginst3008 (P1_SUB_357_U12, P1_U3229);
  not ginst3009 (P1_SUB_357_U13, P1_U3231);
  not ginst3010 (P1_SUB_357_U6, P1_U3233);
  not ginst3011 (P1_SUB_357_U7, P1_U3228);
  not ginst3012 (P1_SUB_357_U8, P1_U3234);
  not ginst3013 (P1_SUB_357_U9, P1_U3232);
  not ginst3014 (P1_SUB_450_U10, P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN);
  not ginst3015 (P1_SUB_450_U11, P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN);
  not ginst3016 (P1_SUB_450_U12, P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN);
  not ginst3017 (P1_SUB_450_U13, P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN);
  not ginst3018 (P1_SUB_450_U14, P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN);
  not ginst3019 (P1_SUB_450_U15, P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN);
  nand ginst3020 (P1_SUB_450_U16, P1_SUB_450_U40, P1_SUB_450_U41);
  not ginst3021 (P1_SUB_450_U17, P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN);
  not ginst3022 (P1_SUB_450_U18, P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN);
  nand ginst3023 (P1_SUB_450_U19, P1_SUB_450_U50, P1_SUB_450_U51);
  nand ginst3024 (P1_SUB_450_U20, P1_SUB_450_U55, P1_SUB_450_U56);
  nand ginst3025 (P1_SUB_450_U21, P1_SUB_450_U60, P1_SUB_450_U61);
  nand ginst3026 (P1_SUB_450_U22, P1_SUB_450_U65, P1_SUB_450_U66);
  nand ginst3027 (P1_SUB_450_U23, P1_SUB_450_U47, P1_SUB_450_U48);
  nand ginst3028 (P1_SUB_450_U24, P1_SUB_450_U52, P1_SUB_450_U53);
  nand ginst3029 (P1_SUB_450_U25, P1_SUB_450_U57, P1_SUB_450_U58);
  nand ginst3030 (P1_SUB_450_U26, P1_SUB_450_U62, P1_SUB_450_U63);
  nand ginst3031 (P1_SUB_450_U27, P1_SUB_450_U36, P1_SUB_450_U37);
  nand ginst3032 (P1_SUB_450_U28, P1_SUB_450_U32, P1_SUB_450_U33);
  not ginst3033 (P1_SUB_450_U29, P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN);
  not ginst3034 (P1_SUB_450_U30, P1_SUB_450_U9);
  nand ginst3035 (P1_SUB_450_U31, P1_SUB_450_U10, P1_SUB_450_U30);
  nand ginst3036 (P1_SUB_450_U32, P1_SUB_450_U29, P1_SUB_450_U31);
  nand ginst3037 (P1_SUB_450_U33, P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN, P1_SUB_450_U9);
  not ginst3038 (P1_SUB_450_U34, P1_SUB_450_U28);
  nand ginst3039 (P1_SUB_450_U35, P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN, P1_SUB_450_U12);
  nand ginst3040 (P1_SUB_450_U36, P1_SUB_450_U28, P1_SUB_450_U35);
  nand ginst3041 (P1_SUB_450_U37, P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN, P1_SUB_450_U11);
  not ginst3042 (P1_SUB_450_U38, P1_SUB_450_U27);
  nand ginst3043 (P1_SUB_450_U39, P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P1_SUB_450_U14);
  nand ginst3044 (P1_SUB_450_U40, P1_SUB_450_U27, P1_SUB_450_U39);
  nand ginst3045 (P1_SUB_450_U41, P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN, P1_SUB_450_U13);
  not ginst3046 (P1_SUB_450_U42, P1_SUB_450_U16);
  nand ginst3047 (P1_SUB_450_U43, P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN, P1_SUB_450_U17);
  nand ginst3048 (P1_SUB_450_U44, P1_SUB_450_U42, P1_SUB_450_U43);
  nand ginst3049 (P1_SUB_450_U45, P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN, P1_SUB_450_U15);
  nand ginst3050 (P1_SUB_450_U46, P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P1_SUB_450_U8);
  nand ginst3051 (P1_SUB_450_U47, P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN, P1_SUB_450_U15);
  nand ginst3052 (P1_SUB_450_U48, P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN, P1_SUB_450_U17);
  not ginst3053 (P1_SUB_450_U49, P1_SUB_450_U23);
  nand ginst3054 (P1_SUB_450_U50, P1_SUB_450_U42, P1_SUB_450_U49);
  nand ginst3055 (P1_SUB_450_U51, P1_SUB_450_U16, P1_SUB_450_U23);
  nand ginst3056 (P1_SUB_450_U52, P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P1_SUB_450_U14);
  nand ginst3057 (P1_SUB_450_U53, P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN, P1_SUB_450_U13);
  not ginst3058 (P1_SUB_450_U54, P1_SUB_450_U24);
  nand ginst3059 (P1_SUB_450_U55, P1_SUB_450_U38, P1_SUB_450_U54);
  nand ginst3060 (P1_SUB_450_U56, P1_SUB_450_U24, P1_SUB_450_U27);
  nand ginst3061 (P1_SUB_450_U57, P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN, P1_SUB_450_U12);
  nand ginst3062 (P1_SUB_450_U58, P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN, P1_SUB_450_U11);
  not ginst3063 (P1_SUB_450_U59, P1_SUB_450_U25);
  nand ginst3064 (P1_SUB_450_U6, P1_SUB_450_U44, P1_SUB_450_U45);
  nand ginst3065 (P1_SUB_450_U60, P1_SUB_450_U34, P1_SUB_450_U59);
  nand ginst3066 (P1_SUB_450_U61, P1_SUB_450_U25, P1_SUB_450_U28);
  nand ginst3067 (P1_SUB_450_U62, P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P1_SUB_450_U10);
  nand ginst3068 (P1_SUB_450_U63, P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN, P1_SUB_450_U29);
  not ginst3069 (P1_SUB_450_U64, P1_SUB_450_U26);
  nand ginst3070 (P1_SUB_450_U65, P1_SUB_450_U30, P1_SUB_450_U64);
  nand ginst3071 (P1_SUB_450_U66, P1_SUB_450_U26, P1_SUB_450_U9);
  nand ginst3072 (P1_SUB_450_U7, P1_SUB_450_U46, P1_SUB_450_U9);
  not ginst3073 (P1_SUB_450_U8, P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN);
  nand ginst3074 (P1_SUB_450_U9, P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN, P1_SUB_450_U18);
  nand ginst3075 (P1_SUB_580_U10, P1_INSTADDRPOINTER_REG_0__SCAN_IN, P1_SUB_580_U7);
  nand ginst3076 (P1_SUB_580_U6, P1_SUB_580_U10, P1_SUB_580_U9);
  not ginst3077 (P1_SUB_580_U7, P1_INSTADDRPOINTER_REG_1__SCAN_IN);
  not ginst3078 (P1_SUB_580_U8, P1_INSTADDRPOINTER_REG_0__SCAN_IN);
  nand ginst3079 (P1_SUB_580_U9, P1_INSTADDRPOINTER_REG_1__SCAN_IN, P1_SUB_580_U8);
  nor ginst3080 (P1_U2352, P1_STATEBS16_REG_SCAN_IN, P1_STATE2_REG_2__SCAN_IN);
  and ginst3081 (P1_U2353, P1_STATE2_REG_2__SCAN_IN, P1_U4231);
  and ginst3082 (P1_U2354, P1_U4265, P1_U4477);
  and ginst3083 (P1_U2355, P1_U2450, P1_U3234);
  and ginst3084 (P1_U2356, P1_R2238_U6, P1_U4192);
  and ginst3085 (P1_U2357, P1_R2167_U17, P1_U3865, P1_U5959);
  and ginst3086 (P1_U2358, P1_U2388, P1_U4224);
  and ginst3087 (P1_U2359, P1_STATE2_REG_2__SCAN_IN, P1_U3431);
  and ginst3088 (P1_U2360, P1_STATE2_REG_2__SCAN_IN, P1_U3414);
  and ginst3089 (P1_U2361, P1_STATE2_REG_3__SCAN_IN, P1_U4224);
  and ginst3090 (P1_U2362, P1_U2359, P1_U4208);
  and ginst3091 (P1_U2363, P1_U2359, P1_U4210);
  and ginst3092 (P1_U2364, P1_U3416, P1_U3864);
  and ginst3093 (P1_U2365, P1_U3416, P1_U4261);
  and ginst3094 (P1_U2366, P1_STATE2_REG_1__SCAN_IN, P1_U3430, P1_U3431);
  and ginst3095 (P1_U2367, P1_STATE2_REG_1__SCAN_IN, P1_R2337_U69, P1_U3431);
  and ginst3096 (P1_U2368, P1_STATE2_REG_0__SCAN_IN, P1_U4235);
  and ginst3097 (P1_U2369, P1_U2362, P1_U4497);
  and ginst3098 (P1_U2370, P1_U3263, P1_U3414);
  and ginst3099 (P1_U2371, P1_U4222, P1_U4449);
  and ginst3100 (P1_U2372, P1_STATE2_REG_0__SCAN_IN, P1_U3416);
  and ginst3101 (P1_U2373, P1_STATE2_REG_3__SCAN_IN, P1_U3431);
  and ginst3102 (P1_U2374, P1_U2360, P1_U4214);
  and ginst3103 (P1_U2375, P1_U2360, P1_U4216);
  and ginst3104 (P1_U2376, P1_U3416, P1_U5798);
  and ginst3105 (P1_U2377, P1_U3414, P1_U3762);
  and ginst3106 (P1_U2378, P1_U2360, P1_U5569);
  and ginst3107 (P1_U2379, P1_U2363, P1_U3280);
  and ginst3108 (P1_U2380, P1_U2360, P1_U7608);
  and ginst3109 (P1_U2381, P1_U2357, P1_U3271);
  and ginst3110 (P1_U2382, P1_U2357, P1_U4477);
  and ginst3111 (P1_U2383, P1_U3391, P1_U4222);
  and ginst3112 (P1_U2384, P1_STATE2_REG_0__SCAN_IN, P1_U3417);
  and ginst3113 (P1_U2385, P1_U3294, P1_U3417);
  and ginst3114 (P1_U2386, P1_U3423, P1_U4223);
  and ginst3115 (P1_U2387, P1_U3884, P1_U4223);
  and ginst3116 (P1_U2388, P1_STATEBS16_REG_SCAN_IN, P1_U4209);
  and ginst3117 (P1_U2389, P1_U2452, P1_U7494);
  and ginst3118 (P1_U2390, P1_U4224, U346);
  and ginst3119 (P1_U2391, P1_U4224, U335);
  and ginst3120 (P1_U2392, P1_U4224, U324);
  and ginst3121 (P1_U2393, P1_U4224, U321);
  and ginst3122 (P1_U2394, P1_U4224, U320);
  and ginst3123 (P1_U2395, P1_U4224, U319);
  and ginst3124 (P1_U2396, P1_U4224, U318);
  and ginst3125 (P1_U2397, P1_U4224, U317);
  and ginst3126 (P1_U2398, P1_U2358, U330);
  and ginst3127 (P1_U2399, P1_U2358, U339);
  and ginst3128 (P1_U2400, P1_U2358, U329);
  and ginst3129 (P1_U2401, P1_U2358, U338);
  and ginst3130 (P1_U2402, P1_U2358, U328);
  and ginst3131 (P1_U2403, P1_U2358, U337);
  and ginst3132 (P1_U2404, P1_U2358, U327);
  and ginst3133 (P1_U2405, P1_U2358, U336);
  and ginst3134 (P1_U2406, P1_U2358, U326);
  and ginst3135 (P1_U2407, P1_U2358, U334);
  and ginst3136 (P1_U2408, P1_U2358, U325);
  and ginst3137 (P1_U2409, P1_U2358, U333);
  and ginst3138 (P1_U2410, P1_U2358, U323);
  and ginst3139 (P1_U2411, P1_U2358, U332);
  and ginst3140 (P1_U2412, P1_U2358, U322);
  and ginst3141 (P1_U2413, P1_U2358, U331);
  and ginst3142 (P1_U2414, P1_U2361, P1_U3271);
  and ginst3143 (P1_U2415, P1_U2361, P1_U3391);
  and ginst3144 (P1_U2416, P1_U2361, P1_U3277);
  and ginst3145 (P1_U2417, P1_U2361, P1_U3284);
  and ginst3146 (P1_U2418, P1_U2361, P1_U3283);
  and ginst3147 (P1_U2419, P1_U2361, P1_U3278);
  and ginst3148 (P1_U2420, P1_U2361, P1_U4173);
  and ginst3149 (P1_U2421, P1_U2361, P1_U4171);
  and ginst3150 (P1_U2422, P1_U4223, P1_U5461);
  and ginst3151 (P1_U2423, P1_U4223, P1_U4231);
  and ginst3152 (P1_U2424, P1_U2384, P1_U3284);
  and ginst3153 (P1_U2425, P1_U2368, P1_U2448);
  and ginst3154 (P1_U2426, P1_U3431, P1_U3889);
  nor ginst3155 (P1_U2427, P1_STATE2_REG_3__SCAN_IN, P1_STATE2_REG_1__SCAN_IN);
  and ginst3156 (P1_U2428, P1_STATE2_REG_2__SCAN_IN, P1_STATE2_REG_1__SCAN_IN);
  and ginst3157 (P1_U2429, P1_U3431, P1_U6366);
  and ginst3158 (P1_U2430, P1_STATE2_REG_1__SCAN_IN, P1_U3387);
  and ginst3159 (P1_U2431, P1_U4199, P1_U7494);
  and ginst3160 (P1_U2432, P1_U3360, P1_U3455);
  and ginst3161 (P1_U2433, P1_U3455, P1_U4540);
  and ginst3162 (P1_U2434, P1_U3360, P1_U7696);
  and ginst3163 (P1_U2435, P1_U4540, P1_U7696);
  and ginst3164 (P1_U2436, P1_U3235, P1_U3301);
  and ginst3165 (P1_U2437, P1_U3301, P1_U4543);
  and ginst3166 (P1_U2438, P1_R2182_U25, P1_R2182_U42);
  and ginst3167 (P1_U2439, P1_R2182_U42, P1_U3316);
  and ginst3168 (P1_U2440, P1_R2182_U25, P1_U3317);
  nor ginst3169 (P1_U2441, P1_R2182_U25, P1_R2182_U42);
  and ginst3170 (P1_U2442, P1_R2182_U33, P1_R2182_U34);
  and ginst3171 (P1_U2443, P1_R2182_U33, P1_U3318);
  and ginst3172 (P1_U2444, P1_R2182_U34, P1_U3319);
  nor ginst3173 (P1_U2445, P1_R2182_U33, P1_R2182_U34);
  and ginst3174 (P1_U2446, P1_STATE2_REG_1__SCAN_IN, P1_U3471);
  and ginst3175 (P1_U2447, P1_U2452, P1_U3577);
  and ginst3176 (P1_U2448, P1_R2167_U17, P1_U3284);
  and ginst3177 (P1_U2449, P1_U3271, P1_U4494);
  and ginst3178 (P1_U2450, P1_STATE2_REG_0__SCAN_IN, P1_U4400);
  and ginst3179 (P1_U2451, P1_STATE2_REG_0__SCAN_IN, P1_U4251);
  and ginst3180 (P1_U2452, P1_U3277, P1_U3391, P1_U4173, P1_U4400);
  and ginst3181 (P1_U2453, P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN, P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN, P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN);
  and ginst3182 (P1_U2454, P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P1_U3266);
  and ginst3183 (P1_U2455, P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN, P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P1_U3266);
  and ginst3184 (P1_U2456, P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN, P1_U3265);
  and ginst3185 (P1_U2457, P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN, P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN, P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P1_U3265);
  and ginst3186 (P1_U2458, P1_U3507, P1_U4378);
  and ginst3187 (P1_U2459, P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN, P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P1_U3264);
  and ginst3188 (P1_U2460, P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P1_U3264, P1_U3266);
  and ginst3189 (P1_U2461, P1_U3505, P1_U3506);
  and ginst3190 (P1_U2462, P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN, P1_U3264, P1_U3265);
  and ginst3191 (P1_U2463, P1_U3503, P1_U3504);
  and ginst3192 (P1_U2464, P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P1_U4380);
  and ginst3193 (P1_U2465, P1_U3501, P1_U3502);
  and ginst3194 (P1_U2466, P1_U3499, P1_U3500);
  and ginst3195 (P1_U2467, P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN, P1_U3270, P1_U4378);
  and ginst3196 (P1_U2468, P1_U3497, P1_U3498);
  nor ginst3197 (P1_U2469, P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN, P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN);
  and ginst3198 (P1_U2470, P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P1_U2469, P1_U3266);
  and ginst3199 (P1_U2471, P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN, P1_U2469, P1_U3265);
  and ginst3200 (P1_U2472, P1_U3270, P1_U4380);
  and ginst3201 (P1_U2473, P1_U3406, P1_U7679, P1_U7680);
  and ginst3202 (P1_U2474, P1_R2144_U49, P1_U3312);
  and ginst3203 (P1_U2475, P1_U3358, P1_U3454);
  and ginst3204 (P1_U2476, P1_R2144_U49, P1_R2144_U8);
  and ginst3205 (P1_U2477, P1_U2476, P1_U4528);
  and ginst3206 (P1_U2478, P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN, P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN);
  and ginst3207 (P1_U2479, P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN, P1_U3303);
  and ginst3208 (P1_U2480, P1_U3315, P1_U4548);
  and ginst3209 (P1_U2481, P1_U2476, P1_U4524);
  and ginst3210 (P1_U2482, P1_U3327, P1_U4606);
  and ginst3211 (P1_U2483, P1_U2476, P1_U4525);
  and ginst3212 (P1_U2484, P1_U3334, P1_U4665);
  and ginst3213 (P1_U2485, P1_R2144_U43, P1_U4526);
  nor ginst3214 (P1_U2486, P1_R2144_U43, P1_R2144_U50);
  and ginst3215 (P1_U2487, P1_U2476, P1_U2486);
  nor ginst3216 (P1_U2488, P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN);
  and ginst3217 (P1_U2489, P1_U3338, P1_U4722);
  and ginst3218 (P1_U2490, P1_U3358, P1_U7693);
  and ginst3219 (P1_U2491, P1_U4528, P1_U4529);
  and ginst3220 (P1_U2492, P1_U3343, P1_U4780);
  and ginst3221 (P1_U2493, P1_U4524, P1_U4529);
  and ginst3222 (P1_U2494, P1_U3347, P1_U4837);
  and ginst3223 (P1_U2495, P1_U4525, P1_U4529);
  and ginst3224 (P1_U2496, P1_U3350, P1_U4895);
  and ginst3225 (P1_U2497, P1_U2486, P1_U4529);
  and ginst3226 (P1_U2498, P1_U3354, P1_U4952);
  and ginst3227 (P1_U2499, P1_U3454, P1_U4531);
  and ginst3228 (P1_U2500, P1_U3357, P1_U3359);
  and ginst3229 (P1_U2501, P1_U2474, P1_U4524);
  and ginst3230 (P1_U2502, P1_U3364, P1_U5065);
  and ginst3231 (P1_U2503, P1_U2474, P1_U4525);
  and ginst3232 (P1_U2504, P1_U3367, P1_U5123);
  and ginst3233 (P1_U2505, P1_U2474, P1_U2486);
  and ginst3234 (P1_U2506, P1_U3371, P1_U5180);
  and ginst3235 (P1_U2507, P1_U4531, P1_U7693);
  nor ginst3236 (P1_U2508, P1_R2144_U49, P1_R2144_U8);
  and ginst3237 (P1_U2509, P1_U2508, P1_U4528);
  nor ginst3238 (P1_U2510, P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN, P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN);
  and ginst3239 (P1_U2511, P1_U3374, P1_U5238);
  and ginst3240 (P1_U2512, P1_U2508, P1_U4524);
  and ginst3241 (P1_U2513, P1_U3378, P1_U5295);
  and ginst3242 (P1_U2514, P1_U2508, P1_U4525);
  and ginst3243 (P1_U2515, P1_U3381, P1_U5353);
  and ginst3244 (P1_U2516, P1_U2486, P1_U2508);
  and ginst3245 (P1_U2517, P1_U3385, P1_U5410);
  and ginst3246 (P1_U2518, P1_U5468, P1_U7699, P1_U7700);
  and ginst3247 (P1_U2519, P1_U3744, P1_U5499);
  and ginst3248 (P1_U2520, P1_U3446, P1_U4219);
  and ginst3249 (P1_U2521, P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN, P1_U3402);
  and ginst3250 (P1_U2522, P1_U5483, P1_U5511);
  and ginst3251 (P1_U2523, P1_U2521, P1_U2522);
  and ginst3252 (P1_U2524, P1_U3266, P1_U3402);
  and ginst3253 (P1_U2525, P1_U2522, P1_U2524);
  and ginst3254 (P1_U2526, P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN, P1_U5519);
  and ginst3255 (P1_U2527, P1_U2522, P1_U2526);
  and ginst3256 (P1_U2528, P1_U3266, P1_U5519);
  and ginst3257 (P1_U2529, P1_U2522, P1_U2528);
  and ginst3258 (P1_U2530, P1_U3401, P1_U5483);
  and ginst3259 (P1_U2531, P1_U2521, P1_U2530);
  and ginst3260 (P1_U2532, P1_U2524, P1_U2530);
  and ginst3261 (P1_U2533, P1_U2526, P1_U2530);
  and ginst3262 (P1_U2534, P1_U2528, P1_U2530);
  and ginst3263 (P1_U2535, P1_U3438, P1_U5511);
  and ginst3264 (P1_U2536, P1_U2521, P1_U2535);
  and ginst3265 (P1_U2537, P1_U2524, P1_U2535);
  and ginst3266 (P1_U2538, P1_U2526, P1_U2535);
  and ginst3267 (P1_U2539, P1_U2528, P1_U2535);
  and ginst3268 (P1_U2540, P1_U3401, P1_U3438);
  and ginst3269 (P1_U2541, P1_U2521, P1_U2540);
  and ginst3270 (P1_U2542, P1_U2524, P1_U2540);
  and ginst3271 (P1_U2543, P1_U2526, P1_U2540);
  and ginst3272 (P1_U2544, P1_U2528, P1_U2540);
  and ginst3273 (P1_U2545, P1_U5480, P1_U7720);
  and ginst3274 (P1_U2546, P1_U2454, P1_U2545);
  and ginst3275 (P1_U2547, P1_U2545, P1_U3498);
  and ginst3276 (P1_U2548, P1_U2545, P1_U4378);
  and ginst3277 (P1_U2549, P1_U2456, P1_U2545);
  and ginst3278 (P1_U2550, P1_U3456, P1_U5480);
  and ginst3279 (P1_U2551, P1_U2454, P1_U2550);
  and ginst3280 (P1_U2552, P1_U2550, P1_U3498);
  and ginst3281 (P1_U2553, P1_U2550, P1_U4378);
  and ginst3282 (P1_U2554, P1_U2456, P1_U2550);
  and ginst3283 (P1_U2555, P1_U3442, P1_U7720);
  and ginst3284 (P1_U2556, P1_U2454, P1_U2555);
  and ginst3285 (P1_U2557, P1_U2555, P1_U3498);
  and ginst3286 (P1_U2558, P1_U2555, P1_U4378);
  and ginst3287 (P1_U2559, P1_U2456, P1_U2555);
  and ginst3288 (P1_U2560, P1_U3442, P1_U3456);
  and ginst3289 (P1_U2561, P1_U2454, P1_U2560);
  and ginst3290 (P1_U2562, P1_U2560, P1_U3498);
  and ginst3291 (P1_U2563, P1_U2560, P1_U4378);
  and ginst3292 (P1_U2564, P1_U2456, P1_U2560);
  and ginst3293 (P1_U2565, P1_U4379, P1_U7065);
  and ginst3294 (P1_U2566, P1_U2460, P1_U7065);
  and ginst3295 (P1_U2567, P1_U2462, P1_U7065);
  and ginst3296 (P1_U2568, P1_U4380, P1_U7065);
  and ginst3297 (P1_U2569, P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN, P1_U7065);
  and ginst3298 (P1_U2570, P1_U2569, P1_U3498);
  and ginst3299 (P1_U2571, P1_U2454, P1_U2569);
  and ginst3300 (P1_U2572, P1_U2456, P1_U2569);
  and ginst3301 (P1_U2573, P1_U2569, P1_U4378);
  and ginst3302 (P1_U2574, P1_U3445, P1_U4379);
  and ginst3303 (P1_U2575, P1_U2460, P1_U3445);
  and ginst3304 (P1_U2576, P1_U2462, P1_U3445);
  and ginst3305 (P1_U2577, P1_U3445, P1_U4380);
  and ginst3306 (P1_U2578, P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN, P1_U3445);
  and ginst3307 (P1_U2579, P1_U2578, P1_U3498);
  and ginst3308 (P1_U2580, P1_U2454, P1_U2578);
  and ginst3309 (P1_U2581, P1_U2456, P1_U2578);
  and ginst3310 (P1_U2582, P1_U2578, P1_U4378);
  and ginst3311 (P1_U2583, P1_U4184, P1_U7790);
  and ginst3312 (P1_U2584, P1_U2524, P1_U2583);
  and ginst3313 (P1_U2585, P1_U2521, P1_U2583);
  and ginst3314 (P1_U2586, P1_U2528, P1_U2583);
  and ginst3315 (P1_U2587, P1_U2526, P1_U2583);
  and ginst3316 (P1_U2588, P1_U3452, P1_U7790);
  and ginst3317 (P1_U2589, P1_U2524, P1_U2588);
  and ginst3318 (P1_U2590, P1_U2521, P1_U2588);
  and ginst3319 (P1_U2591, P1_U2528, P1_U2588);
  and ginst3320 (P1_U2592, P1_U2526, P1_U2588);
  and ginst3321 (P1_U2593, P1_U3457, P1_U4184);
  and ginst3322 (P1_U2594, P1_U2524, P1_U2593);
  and ginst3323 (P1_U2595, P1_U2521, P1_U2593);
  and ginst3324 (P1_U2596, P1_U2528, P1_U2593);
  and ginst3325 (P1_U2597, P1_U2526, P1_U2593);
  and ginst3326 (P1_U2598, P1_U3452, P1_U3457);
  and ginst3327 (P1_U2599, P1_U2524, P1_U2598);
  and ginst3328 (P1_U2600, P1_U2521, P1_U2598);
  and ginst3329 (P1_U2601, P1_U2528, P1_U2598);
  and ginst3330 (P1_U2602, P1_U2526, P1_U2598);
  and ginst3331 (P1_U2603, P1_STATE2_REG_0__SCAN_IN, P1_U3389);
  and ginst3332 (P1_U2604, P1_EBX_REG_31__SCAN_IN, P1_U2379);
  and ginst3333 (P1_U2605, P1_U2607, P1_U3530, P1_U3531, P1_U3532, P1_U3533);
  and ginst3334 (P1_U2606, P1_U3427, P1_U7504);
  and ginst3335 (P1_U2607, P1_U7671, P1_U7672);
  and ginst3336 (P1_U2608, P1_U7786, P1_U7787);
  nand ginst3337 (P1_U2609, P1_U6853, P1_U6854, P1_U6855);
  nand ginst3338 (P1_U2610, P1_U4026, P1_U6856);
  nand ginst3339 (P1_U2611, P1_U6841, P1_U6842, P1_U6843);
  nand ginst3340 (P1_U2612, P1_U6844, P1_U6845, P1_U6846);
  nand ginst3341 (P1_U2613, P1_U6847, P1_U6848, P1_U6849);
  nand ginst3342 (P1_U2614, P1_U4005, P1_U6756);
  nand ginst3343 (P1_U2615, P1_U4004, P1_U6753);
  nand ginst3344 (P1_U2616, P1_U6850, P1_U6851, P1_U6852);
  nand ginst3345 (P1_U2617, P1_U4003, P1_U6750);
  nand ginst3346 (P1_U2618, P1_U4002, P1_U6747);
  and ginst3347 (P1_U2620, P1_R2144_U145, P1_U6746);
  and ginst3348 (P1_U2621, P1_R2144_U145, P1_U6746);
  and ginst3349 (P1_U2622, P1_R2144_U145, P1_U6746);
  and ginst3350 (P1_U2623, P1_R2144_U145, P1_U6746);
  and ginst3351 (P1_U2624, P1_R2144_U145, P1_U6746);
  and ginst3352 (P1_U2625, P1_R2144_U145, P1_U6746);
  and ginst3353 (P1_U2626, P1_R2144_U145, P1_U6746);
  and ginst3354 (P1_U2627, P1_R2144_U145, P1_U6746);
  and ginst3355 (P1_U2628, P1_R2144_U145, P1_U6746);
  and ginst3356 (P1_U2629, P1_R2144_U145, P1_U6746);
  and ginst3357 (P1_U2630, P1_R2144_U145, P1_U6746);
  and ginst3358 (P1_U2631, P1_R2144_U145, P1_U6746);
  and ginst3359 (P1_U2632, P1_R2144_U145, P1_U6746);
  and ginst3360 (P1_U2633, P1_R2144_U145, P1_U6746);
  and ginst3361 (P1_U2634, P1_R2144_U11, P1_U6746);
  and ginst3362 (P1_U2635, P1_R2144_U37, P1_U6746);
  and ginst3363 (P1_U2636, P1_R2144_U38, P1_U6746);
  and ginst3364 (P1_U2637, P1_R2144_U39, P1_U6746);
  and ginst3365 (P1_U2638, P1_R2144_U40, P1_U6746);
  and ginst3366 (P1_U2639, P1_R2144_U41, P1_U6746);
  and ginst3367 (P1_U2640, P1_R2144_U42, P1_U6746);
  and ginst3368 (P1_U2641, P1_R2144_U30, P1_U6746);
  and ginst3369 (P1_U2642, P1_R2144_U80, P1_U6746);
  and ginst3370 (P1_U2643, P1_R2144_U10, P1_U6746);
  and ginst3371 (P1_U2644, P1_R2144_U9, P1_U6746);
  and ginst3372 (P1_U2645, P1_R2144_U45, P1_U6746);
  and ginst3373 (P1_U2646, P1_R2144_U47, P1_U6746);
  and ginst3374 (P1_U2647, P1_R2144_U8, P1_U6746);
  nand ginst3375 (P1_U2648, P1_U3440, P1_U6869);
  and ginst3376 (P1_U2649, P1_R2144_U50, P1_U6746);
  and ginst3377 (P1_U2650, P1_STATE2_REG_2__SCAN_IN, P1_U6870);
  nand ginst3378 (P1_U2651, P1_U6768, P1_U6769, P1_U6770);
  nand ginst3379 (P1_U2652, P1_U4009, P1_U6771);
  nand ginst3380 (P1_U2653, P1_U4011, P1_U6780);
  nand ginst3381 (P1_U2654, P1_U4012, P1_U6784);
  nand ginst3382 (P1_U2655, P1_U4013, P1_U6788);
  nand ginst3383 (P1_U2656, P1_U4014, P1_U6792);
  nand ginst3384 (P1_U2657, P1_U4015, P1_U6796);
  nand ginst3385 (P1_U2658, P1_U4016, P1_U6800);
  nand ginst3386 (P1_U2659, P1_U4017, P1_U6804);
  nand ginst3387 (P1_U2660, P1_U4018, P1_U6808);
  nand ginst3388 (P1_U2661, P1_U4019, P1_U6812);
  nand ginst3389 (P1_U2662, P1_U4020, P1_U6816);
  nand ginst3390 (P1_U2663, P1_U4022, P1_U6825);
  nand ginst3391 (P1_U2664, P1_U4023, P1_U6829);
  nand ginst3392 (P1_U2665, P1_U4024, P1_U6833);
  nand ginst3393 (P1_U2666, P1_U4025, P1_U6837);
  nand ginst3394 (P1_U2667, P1_U4006, P1_U6759);
  nand ginst3395 (P1_U2668, P1_U4008, P1_U6763, P1_U6766, P1_U6767);
  nand ginst3396 (P1_U2669, P1_U4010, P1_U6775, P1_U6778, P1_U6779);
  nand ginst3397 (P1_U2670, P1_U4021, P1_U6820, P1_U6823, P1_U6824);
  nand ginst3398 (P1_U2671, P1_U4027, P1_U6859, P1_U6862, P1_U6863);
  nand ginst3399 (P1_U2672, P1_U6864, P1_U6865, P1_U6866, P1_U6867, P1_U6868);
  nand ginst3400 (P1_U2673, P1_U7457, P1_U7458);
  nand ginst3401 (P1_U2674, P1_U7459, P1_U7460);
  nand ginst3402 (P1_U2675, P1_U4168, P1_U7463);
  nand ginst3403 (P1_U2676, P1_U4169, P1_U7466);
  nand ginst3404 (P1_U2677, P1_U7467, P1_U7793, P1_U7794);
  nand ginst3405 (P1_U2678, P1_U3284, P1_U7456);
  nand ginst3406 (P1_U2679, P1_U7404, P1_U7405);
  nand ginst3407 (P1_U2680, P1_U7406, P1_U7407);
  nand ginst3408 (P1_U2681, P1_U7410, P1_U7411);
  nand ginst3409 (P1_U2682, P1_U7412, P1_U7413);
  nand ginst3410 (P1_U2683, P1_U7414, P1_U7415);
  nand ginst3411 (P1_U2684, P1_U7416, P1_U7417);
  nand ginst3412 (P1_U2685, P1_U7418, P1_U7419);
  nand ginst3413 (P1_U2686, P1_U7420, P1_U7421);
  nand ginst3414 (P1_U2687, P1_U7422, P1_U7423);
  nand ginst3415 (P1_U2688, P1_U7424, P1_U7425);
  nand ginst3416 (P1_U2689, P1_U7426, P1_U7427);
  nand ginst3417 (P1_U2690, P1_U7428, P1_U7429);
  nand ginst3418 (P1_U2691, P1_U7432, P1_U7433);
  nand ginst3419 (P1_U2692, P1_U7434, P1_U7435);
  nand ginst3420 (P1_U2693, P1_U7436, P1_U7437);
  nand ginst3421 (P1_U2694, P1_U7438, P1_U7439);
  nand ginst3422 (P1_U2695, P1_U7440, P1_U7441);
  nand ginst3423 (P1_U2696, P1_U7442, P1_U7443);
  nand ginst3424 (P1_U2697, P1_U7444, P1_U7445);
  nand ginst3425 (P1_U2698, P1_U7446, P1_U7447);
  nand ginst3426 (P1_U2699, P1_U7448, P1_U7449);
  nand ginst3427 (P1_U2700, P1_U7450, P1_U7451);
  nand ginst3428 (P1_U2701, P1_U7392, P1_U7393);
  nand ginst3429 (P1_U2702, P1_U7394, P1_U7395);
  nand ginst3430 (P1_U2703, P1_U7396, P1_U7397);
  nand ginst3431 (P1_U2704, P1_U7398, P1_U7399);
  nand ginst3432 (P1_U2705, P1_U7400, P1_U7401);
  nand ginst3433 (P1_U2706, P1_U7402, P1_U7403);
  nand ginst3434 (P1_U2707, P1_U7408, P1_U7409);
  nand ginst3435 (P1_U2708, P1_U7430, P1_U7431);
  nand ginst3436 (P1_U2709, P1_U7452, P1_U7453);
  nand ginst3437 (P1_U2710, P1_U7454, P1_U7455);
  nand ginst3438 (P1_U2711, P1_U7376, P1_U7377);
  nand ginst3439 (P1_U2712, P1_U7378, P1_U7379);
  nand ginst3440 (P1_U2713, P1_U4165, P1_U4239);
  nand ginst3441 (P1_U2714, P1_U3434, P1_U4166, P1_U7385, P1_U7386);
  nand ginst3442 (P1_U2715, P1_U4167, P1_U4239);
  nand ginst3443 (P1_U2716, P1_U7364, P1_U7365);
  nand ginst3444 (P1_U2717, P1_U7366, P1_U7367);
  nand ginst3445 (P1_U2718, P1_U4161, P1_U7368);
  nand ginst3446 (P1_U2719, P1_U4162, P1_U7370);
  nand ginst3447 (P1_U2720, P1_U4163, P1_U7372);
  nand ginst3448 (P1_U2721, P1_U4164, P1_U7374);
  nand ginst3449 (P1_U2722, P1_U4159, P1_U4192);
  and ginst3450 (P1_U2723, P1_U7083, P1_U7236);
  and ginst3451 (P1_U2724, P1_U7083, P1_U7253);
  and ginst3452 (P1_U2725, P1_U7083, P1_U7270);
  and ginst3453 (P1_U2726, P1_U7083, P1_U7620);
  and ginst3454 (P1_U2727, P1_U7083, P1_U7302);
  and ginst3455 (P1_U2728, P1_U7083, P1_U7319);
  and ginst3456 (P1_U2729, P1_U7083, P1_U7336);
  and ginst3457 (P1_U2730, P1_U7083, P1_U7353);
  nand ginst3458 (P1_U2731, P1_U2606, P1_U7354);
  and ginst3459 (P1_U2732, P1_U7082, P1_U7083);
  and ginst3460 (P1_U2733, P1_U7083, P1_U7114);
  and ginst3461 (P1_U2734, P1_U7083, P1_U7131);
  and ginst3462 (P1_U2735, P1_U7083, P1_U7618);
  and ginst3463 (P1_U2736, P1_U7083, P1_U7163);
  and ginst3464 (P1_U2737, P1_U7083, P1_U7180);
  and ginst3465 (P1_U2738, P1_U7083, P1_U7197);
  and ginst3466 (P1_U2739, P1_U7083, P1_U7214);
  and ginst3467 (P1_U2740, P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN, P1_U7063);
  nand ginst3468 (P1_U2741, P1_U4078, P1_U7096);
  and ginst3469 (P1_U2742, P1_U7491, P1_U7492);
  and ginst3470 (P1_U2743, P1_U7470, P1_U7506);
  and ginst3471 (P1_U2744, P1_U7478, P1_U7479);
  nand ginst3472 (P1_U2745, P1_U7047, P1_U7048);
  nand ginst3473 (P1_U2746, P1_U7049, P1_U7050);
  nand ginst3474 (P1_U2747, P1_U7051, P1_U7052);
  nand ginst3475 (P1_U2748, P1_U7053, P1_U7616);
  nand ginst3476 (P1_U2749, P1_U7054, P1_U7055);
  nand ginst3477 (P1_U2750, P1_U7056, P1_U7057);
  nand ginst3478 (P1_U2751, P1_U4061, P1_U7058);
  nand ginst3479 (P1_U2752, P1_U4062, P1_U7060, P1_U7061);
  and ginst3480 (P1_U2753, P1_U6909, P1_U6957);
  and ginst3481 (P1_U2754, P1_U6909, P1_U6974);
  and ginst3482 (P1_U2755, P1_U6909, P1_U6991);
  and ginst3483 (P1_U2756, P1_U6909, P1_U7615);
  and ginst3484 (P1_U2757, P1_U6909, P1_U7023);
  and ginst3485 (P1_U2758, P1_U6909, P1_U7040);
  and ginst3486 (P1_U2759, P1_U6908, P1_U6909);
  and ginst3487 (P1_U2760, P1_U6909, P1_U6926);
  nand ginst3488 (P1_U2761, P1_U6927, P1_U6928);
  nand ginst3489 (P1_U2762, P1_U6929, P1_U6930);
  nand ginst3490 (P1_U2763, P1_U6931, P1_U6932);
  nand ginst3491 (P1_U2764, P1_U6933, P1_U6934);
  nand ginst3492 (P1_U2765, P1_U6935, P1_U6936, P1_U6937);
  nand ginst3493 (P1_U2766, P1_U6938, P1_U6939, P1_U6940);
  nand ginst3494 (P1_U2767, P1_U7041, P1_U7042, P1_U7043);
  nand ginst3495 (P1_U2768, P1_U7044, P1_U7045, P1_U7046);
  and ginst3496 (P1_U2769, P1_R2144_U145, P1_U4159);
  and ginst3497 (P1_U2770, P1_R2144_U145, P1_U4159);
  and ginst3498 (P1_U2771, P1_R2144_U145, P1_U4159);
  and ginst3499 (P1_U2772, P1_R2144_U145, P1_U4159);
  and ginst3500 (P1_U2773, P1_R2144_U145, P1_U4159);
  and ginst3501 (P1_U2774, P1_R2144_U145, P1_U4159);
  and ginst3502 (P1_U2775, P1_R2144_U145, P1_U4159);
  and ginst3503 (P1_U2776, P1_R2144_U145, P1_U4159);
  and ginst3504 (P1_U2777, P1_R2144_U145, P1_U4159);
  and ginst3505 (P1_U2778, P1_R2144_U145, P1_U4159);
  and ginst3506 (P1_U2779, P1_R2144_U145, P1_U4159);
  and ginst3507 (P1_U2780, P1_R2144_U145, P1_U4159);
  and ginst3508 (P1_U2781, P1_R2144_U145, P1_U4159);
  and ginst3509 (P1_U2782, P1_R2144_U145, P1_U4159);
  and ginst3510 (P1_U2783, P1_R2144_U145, P1_U4159);
  and ginst3511 (P1_U2784, P1_R2144_U11, P1_U4159);
  and ginst3512 (P1_U2785, P1_R2144_U37, P1_U4159);
  and ginst3513 (P1_U2786, P1_R2144_U38, P1_U4159);
  and ginst3514 (P1_U2787, P1_R2144_U39, P1_U4159);
  and ginst3515 (P1_U2788, P1_R2144_U40, P1_U4159);
  and ginst3516 (P1_U2789, P1_R2144_U41, P1_U4159);
  and ginst3517 (P1_U2790, P1_R2144_U42, P1_U4159);
  and ginst3518 (P1_U2791, P1_R2144_U30, P1_U4159);
  nand ginst3519 (P1_U2792, P1_U6871, P1_U6872);
  nand ginst3520 (P1_U2793, P1_U6873, P1_U6874);
  nand ginst3521 (P1_U2794, P1_U6875, P1_U6876);
  nand ginst3522 (P1_U2795, P1_U6877, P1_U6878);
  nand ginst3523 (P1_U2796, P1_U6879, P1_U6880);
  nand ginst3524 (P1_U2797, P1_U6881, P1_U6882);
  nand ginst3525 (P1_U2798, P1_U6883, P1_U6884, P1_U6885);
  nand ginst3526 (P1_U2799, P1_U4028, P1_U6886, P1_U6887);
  nand ginst3527 (P1_U2800, P1_U6889, P1_U6890, P1_U6891);
  nand ginst3528 (P1_U2801, P1_U3432, P1_U6617, P1_U7498);
  nand ginst3529 (P1_U2802, P1_U6613, P1_U7650);
  nand ginst3530 (P1_U2803, P1_U6611, P1_U6612);
  nand ginst3531 (P1_U2804, P1_U4243, P1_U7768, P1_U7769);
  nand ginst3532 (P1_U2805, P1_U4243, P1_U7764, P1_U7765);
  nand ginst3533 (P1_U2806, P1_U4248, P1_U6601);
  nand ginst3534 (P1_U2807, P1_U4240, P1_U7756, P1_U7757);
  nand ginst3535 (P1_U2808, P1_U4240, P1_U7746, P1_U7747);
  nand ginst3536 (P1_U2809, P1_U3948, P1_U3949, P1_U6591, P1_U6593, P1_U6595);
  nand ginst3537 (P1_U2810, P1_U3946, P1_U3947, P1_U6584, P1_U6586, P1_U6588);
  nand ginst3538 (P1_U2811, P1_U3944, P1_U3945, P1_U6577, P1_U6579, P1_U6581);
  nand ginst3539 (P1_U2812, P1_U3942, P1_U3943, P1_U6570, P1_U6572, P1_U6574);
  nand ginst3540 (P1_U2813, P1_U3940, P1_U3941, P1_U6563, P1_U6565, P1_U6567);
  nand ginst3541 (P1_U2814, P1_U3938, P1_U3939, P1_U6556, P1_U6558, P1_U6560);
  nand ginst3542 (P1_U2815, P1_U3936, P1_U3937, P1_U6549, P1_U6551, P1_U6553);
  nand ginst3543 (P1_U2816, P1_U3934, P1_U3935, P1_U6542, P1_U6544, P1_U6546);
  nand ginst3544 (P1_U2817, P1_U3932, P1_U3933, P1_U6535, P1_U6537, P1_U6539);
  nand ginst3545 (P1_U2818, P1_U3930, P1_U3931, P1_U6528, P1_U6530, P1_U6532);
  nand ginst3546 (P1_U2819, P1_U3928, P1_U3929, P1_U6521, P1_U6523, P1_U6525);
  nand ginst3547 (P1_U2820, P1_U3926, P1_U3927, P1_U6514, P1_U6516, P1_U6518);
  nand ginst3548 (P1_U2821, P1_U3924, P1_U3925, P1_U6507, P1_U6509, P1_U6511);
  nand ginst3549 (P1_U2822, P1_U3922, P1_U3923, P1_U6500, P1_U6502, P1_U6504);
  nand ginst3550 (P1_U2823, P1_U3920, P1_U3921, P1_U6493, P1_U6495, P1_U6497);
  nand ginst3551 (P1_U2824, P1_U3918, P1_U3919, P1_U6487, P1_U6488, P1_U6490);
  nand ginst3552 (P1_U2825, P1_U3916, P1_U3917, P1_U6480, P1_U6481, P1_U6483);
  nand ginst3553 (P1_U2826, P1_U3914, P1_U3915, P1_U6473, P1_U6474, P1_U6476);
  nand ginst3554 (P1_U2827, P1_U3912, P1_U3913, P1_U6466, P1_U6467, P1_U6469);
  nand ginst3555 (P1_U2828, P1_U3910, P1_U3911, P1_U6459, P1_U6460, P1_U6462);
  nand ginst3556 (P1_U2829, P1_U3908, P1_U3909, P1_U6452, P1_U6453, P1_U6455);
  nand ginst3557 (P1_U2830, P1_U3906, P1_U3907, P1_U6445, P1_U6446, P1_U6448);
  nand ginst3558 (P1_U2831, P1_U3904, P1_U3905, P1_U6438, P1_U6439, P1_U6441);
  nand ginst3559 (P1_U2832, P1_U3902, P1_U3903, P1_U6431, P1_U6432, P1_U6434);
  nand ginst3560 (P1_U2833, P1_U3900, P1_U3901, P1_U6424, P1_U6425, P1_U6427);
  nand ginst3561 (P1_U2834, P1_U3898, P1_U3899, P1_U6417, P1_U6418, P1_U6420);
  nand ginst3562 (P1_U2835, P1_U3896, P1_U3897, P1_U6409, P1_U6410);
  nand ginst3563 (P1_U2836, P1_U3894, P1_U3895, P1_U6401, P1_U6402, P1_U6403);
  nand ginst3564 (P1_U2837, P1_U3893, P1_U6392, P1_U6393, P1_U6394);
  nand ginst3565 (P1_U2838, P1_U3892, P1_U6384, P1_U6385, P1_U6386);
  nand ginst3566 (P1_U2839, P1_U3891, P1_U6376, P1_U6377, P1_U6378);
  nand ginst3567 (P1_U2840, P1_U3890, P1_U6368, P1_U6369, P1_U6370);
  nand ginst3568 (P1_U2841, P1_U6358, P1_U6359);
  nand ginst3569 (P1_U2842, P1_U6355, P1_U6356, P1_U6357);
  nand ginst3570 (P1_U2843, P1_U6352, P1_U6353, P1_U6354);
  nand ginst3571 (P1_U2844, P1_U6349, P1_U6350, P1_U6351);
  nand ginst3572 (P1_U2845, P1_U6346, P1_U6347, P1_U6348);
  nand ginst3573 (P1_U2846, P1_U6343, P1_U6344, P1_U6345);
  nand ginst3574 (P1_U2847, P1_U6340, P1_U6341, P1_U6342);
  nand ginst3575 (P1_U2848, P1_U6337, P1_U6338, P1_U6339);
  nand ginst3576 (P1_U2849, P1_U6334, P1_U6335, P1_U6336);
  nand ginst3577 (P1_U2850, P1_U6331, P1_U6332, P1_U6333);
  nand ginst3578 (P1_U2851, P1_U6328, P1_U6329, P1_U6330);
  nand ginst3579 (P1_U2852, P1_U6325, P1_U6326, P1_U6327);
  nand ginst3580 (P1_U2853, P1_U6322, P1_U6323, P1_U6324);
  nand ginst3581 (P1_U2854, P1_U6319, P1_U6320, P1_U6321);
  nand ginst3582 (P1_U2855, P1_U6316, P1_U6317, P1_U6318);
  nand ginst3583 (P1_U2856, P1_U6313, P1_U6314, P1_U6315);
  nand ginst3584 (P1_U2857, P1_U6310, P1_U6311, P1_U6312);
  nand ginst3585 (P1_U2858, P1_U6307, P1_U6308, P1_U6309);
  nand ginst3586 (P1_U2859, P1_U6304, P1_U6305, P1_U6306);
  nand ginst3587 (P1_U2860, P1_U6301, P1_U6302, P1_U6303);
  nand ginst3588 (P1_U2861, P1_U6298, P1_U6299, P1_U6300);
  nand ginst3589 (P1_U2862, P1_U6295, P1_U6296, P1_U6297);
  nand ginst3590 (P1_U2863, P1_U6292, P1_U6293, P1_U6294);
  nand ginst3591 (P1_U2864, P1_U6289, P1_U6290, P1_U6291);
  nand ginst3592 (P1_U2865, P1_U6286, P1_U6287, P1_U6288);
  nand ginst3593 (P1_U2866, P1_U6283, P1_U6284, P1_U6285);
  nand ginst3594 (P1_U2867, P1_U6280, P1_U6281, P1_U6282);
  nand ginst3595 (P1_U2868, P1_U6277, P1_U6278, P1_U6279);
  nand ginst3596 (P1_U2869, P1_U6274, P1_U6275, P1_U6276);
  nand ginst3597 (P1_U2870, P1_U6271, P1_U6272, P1_U6273);
  nand ginst3598 (P1_U2871, P1_U6268, P1_U6269, P1_U6270);
  nand ginst3599 (P1_U2872, P1_U6265, P1_U6266, P1_U6267);
  nand ginst3600 (P1_U2873, P1_U4176, P1_U6262);
  nand ginst3601 (P1_U2874, P1_U6258, P1_U6259, P1_U6260, P1_U6261);
  nand ginst3602 (P1_U2875, P1_U6254, P1_U6255, P1_U6256, P1_U6257);
  nand ginst3603 (P1_U2876, P1_U6250, P1_U6251, P1_U6252, P1_U6253);
  nand ginst3604 (P1_U2877, P1_U6246, P1_U6247, P1_U6248, P1_U6249);
  nand ginst3605 (P1_U2878, P1_U6242, P1_U6243, P1_U6244, P1_U6245);
  nand ginst3606 (P1_U2879, P1_U6238, P1_U6239, P1_U6240, P1_U6241);
  nand ginst3607 (P1_U2880, P1_U6234, P1_U6235, P1_U6236, P1_U6237);
  nand ginst3608 (P1_U2881, P1_U6230, P1_U6231, P1_U6232, P1_U6233);
  nand ginst3609 (P1_U2882, P1_U6226, P1_U6227, P1_U6228, P1_U6229);
  nand ginst3610 (P1_U2883, P1_U6222, P1_U6223, P1_U6224, P1_U6225);
  nand ginst3611 (P1_U2884, P1_U6218, P1_U6219, P1_U6220, P1_U6221);
  nand ginst3612 (P1_U2885, P1_U6214, P1_U6215, P1_U6216, P1_U6217);
  nand ginst3613 (P1_U2886, P1_U6210, P1_U6211, P1_U6212, P1_U6213);
  nand ginst3614 (P1_U2887, P1_U6206, P1_U6207, P1_U6208, P1_U6209);
  nand ginst3615 (P1_U2888, P1_U6202, P1_U6203, P1_U6204, P1_U6205);
  nand ginst3616 (P1_U2889, P1_U6199, P1_U6200, P1_U6201);
  nand ginst3617 (P1_U2890, P1_U6196, P1_U6197, P1_U6198);
  nand ginst3618 (P1_U2891, P1_U6193, P1_U6194, P1_U6195);
  nand ginst3619 (P1_U2892, P1_U6190, P1_U6191, P1_U6192);
  nand ginst3620 (P1_U2893, P1_U6187, P1_U6188, P1_U6189);
  nand ginst3621 (P1_U2894, P1_U6184, P1_U6185, P1_U6186);
  nand ginst3622 (P1_U2895, P1_U6181, P1_U6182, P1_U6183);
  nand ginst3623 (P1_U2896, P1_U6178, P1_U6179, P1_U6180);
  nand ginst3624 (P1_U2897, P1_U6175, P1_U6176, P1_U6177);
  nand ginst3625 (P1_U2898, P1_U6172, P1_U6173, P1_U6174);
  nand ginst3626 (P1_U2899, P1_U6169, P1_U6170, P1_U6171);
  nand ginst3627 (P1_U2900, P1_U6166, P1_U6167, P1_U6168);
  nand ginst3628 (P1_U2901, P1_U6163, P1_U6164, P1_U6165);
  nand ginst3629 (P1_U2902, P1_U6160, P1_U6161, P1_U6162);
  nand ginst3630 (P1_U2903, P1_U6157, P1_U6158, P1_U6159);
  nand ginst3631 (P1_U2904, P1_U6154, P1_U6155, P1_U6156);
  and ginst3632 (P1_U2905, P1_DATAO_REG_31__SCAN_IN, P1_U6055);
  nand ginst3633 (P1_U2906, P1_U3882, P1_U6146);
  nand ginst3634 (P1_U2907, P1_U3881, P1_U6143);
  nand ginst3635 (P1_U2908, P1_U3880, P1_U6140);
  nand ginst3636 (P1_U2909, P1_U3879, P1_U6137);
  nand ginst3637 (P1_U2910, P1_U3878, P1_U6134);
  nand ginst3638 (P1_U2911, P1_U3877, P1_U6131);
  nand ginst3639 (P1_U2912, P1_U3876, P1_U6128);
  nand ginst3640 (P1_U2913, P1_U3875, P1_U6125);
  nand ginst3641 (P1_U2914, P1_U3874, P1_U6122);
  nand ginst3642 (P1_U2915, P1_U3873, P1_U6119);
  nand ginst3643 (P1_U2916, P1_U3872, P1_U6116);
  nand ginst3644 (P1_U2917, P1_U3871, P1_U6113);
  nand ginst3645 (P1_U2918, P1_U3870, P1_U6110);
  nand ginst3646 (P1_U2919, P1_U3869, P1_U6107);
  nand ginst3647 (P1_U2920, P1_U3868, P1_U6104);
  nand ginst3648 (P1_U2921, P1_U6101, P1_U6102, P1_U6103);
  nand ginst3649 (P1_U2922, P1_U6098, P1_U6099, P1_U6100);
  nand ginst3650 (P1_U2923, P1_U6095, P1_U6096, P1_U6097);
  nand ginst3651 (P1_U2924, P1_U6092, P1_U6093, P1_U6094);
  nand ginst3652 (P1_U2925, P1_U6089, P1_U6090, P1_U6091);
  nand ginst3653 (P1_U2926, P1_U6086, P1_U6087, P1_U6088);
  nand ginst3654 (P1_U2927, P1_U6083, P1_U6084, P1_U6085);
  nand ginst3655 (P1_U2928, P1_U6080, P1_U6081, P1_U6082);
  nand ginst3656 (P1_U2929, P1_U6077, P1_U6078, P1_U6079);
  nand ginst3657 (P1_U2930, P1_U6074, P1_U6075, P1_U6076);
  nand ginst3658 (P1_U2931, P1_U6071, P1_U6072, P1_U6073);
  nand ginst3659 (P1_U2932, P1_U6068, P1_U6069, P1_U6070);
  nand ginst3660 (P1_U2933, P1_U6065, P1_U6066, P1_U6067);
  nand ginst3661 (P1_U2934, P1_U6062, P1_U6063, P1_U6064);
  nand ginst3662 (P1_U2935, P1_U6059, P1_U6060, P1_U6061);
  nand ginst3663 (P1_U2936, P1_U6056, P1_U6057, P1_U6058);
  nand ginst3664 (P1_U2937, P1_U7540, P1_U7542);
  nand ginst3665 (P1_U2938, P1_U7539, P1_U7544);
  nand ginst3666 (P1_U2939, P1_U7538, P1_U7546);
  nand ginst3667 (P1_U2940, P1_U7537, P1_U7548);
  nand ginst3668 (P1_U2941, P1_U7536, P1_U7550);
  nand ginst3669 (P1_U2942, P1_U7535, P1_U7552);
  nand ginst3670 (P1_U2943, P1_U7534, P1_U7554);
  nand ginst3671 (P1_U2944, P1_U7533, P1_U7556);
  nand ginst3672 (P1_U2945, P1_U7532, P1_U7558);
  nand ginst3673 (P1_U2946, P1_U7531, P1_U7560);
  nand ginst3674 (P1_U2947, P1_U7530, P1_U7562);
  nand ginst3675 (P1_U2948, P1_U7529, P1_U7564);
  nand ginst3676 (P1_U2949, P1_U7528, P1_U7566);
  nand ginst3677 (P1_U2950, P1_U7527, P1_U7568);
  nand ginst3678 (P1_U2951, P1_U7526, P1_U7570);
  nand ginst3679 (P1_U2952, P1_U7525, P1_U7572);
  nand ginst3680 (P1_U2953, P1_U7524, P1_U7574);
  nand ginst3681 (P1_U2954, P1_U7523, P1_U7576);
  nand ginst3682 (P1_U2955, P1_U7522, P1_U7578);
  nand ginst3683 (P1_U2956, P1_U7521, P1_U7580);
  nand ginst3684 (P1_U2957, P1_U7520, P1_U7582);
  nand ginst3685 (P1_U2958, P1_U7519, P1_U7584);
  nand ginst3686 (P1_U2959, P1_U7518, P1_U7586);
  nand ginst3687 (P1_U2960, P1_U7517, P1_U7588);
  nand ginst3688 (P1_U2961, P1_U7516, P1_U7590);
  nand ginst3689 (P1_U2962, P1_U7515, P1_U7592);
  nand ginst3690 (P1_U2963, P1_U7514, P1_U7594);
  nand ginst3691 (P1_U2964, P1_U7513, P1_U7596);
  nand ginst3692 (P1_U2965, P1_U7512, P1_U7598);
  nand ginst3693 (P1_U2966, P1_U7511, P1_U7600);
  nand ginst3694 (P1_U2967, P1_U7510, P1_U7602);
  nand ginst3695 (P1_U2968, P1_U5954, P1_U5955, P1_U5956, P1_U5957, P1_U5958);
  nand ginst3696 (P1_U2969, P1_U5949, P1_U5950, P1_U5951, P1_U5952, P1_U5953);
  nand ginst3697 (P1_U2970, P1_U5944, P1_U5945, P1_U5946, P1_U5947, P1_U5948);
  nand ginst3698 (P1_U2971, P1_U5939, P1_U5940, P1_U5941, P1_U5942, P1_U5943);
  nand ginst3699 (P1_U2972, P1_U5934, P1_U5935, P1_U5936, P1_U5937, P1_U5938);
  nand ginst3700 (P1_U2973, P1_U5929, P1_U5930, P1_U5931, P1_U5932, P1_U5933);
  nand ginst3701 (P1_U2974, P1_U5924, P1_U5925, P1_U5926, P1_U5927, P1_U5928);
  nand ginst3702 (P1_U2975, P1_U5919, P1_U5920, P1_U5921, P1_U5922, P1_U5923);
  nand ginst3703 (P1_U2976, P1_U5914, P1_U5915, P1_U5916, P1_U5917, P1_U5918);
  nand ginst3704 (P1_U2977, P1_U5909, P1_U5910, P1_U5911, P1_U5912, P1_U5913);
  nand ginst3705 (P1_U2978, P1_U5904, P1_U5905, P1_U5906, P1_U5907, P1_U5908);
  nand ginst3706 (P1_U2979, P1_U5899, P1_U5900, P1_U5901, P1_U5902, P1_U5903);
  nand ginst3707 (P1_U2980, P1_U5894, P1_U5895, P1_U5896, P1_U5897, P1_U5898);
  nand ginst3708 (P1_U2981, P1_U5889, P1_U5890, P1_U5891, P1_U5892, P1_U5893);
  nand ginst3709 (P1_U2982, P1_U5884, P1_U5885, P1_U5886, P1_U5887, P1_U5888);
  nand ginst3710 (P1_U2983, P1_U5879, P1_U5880, P1_U5881, P1_U5882, P1_U5883);
  nand ginst3711 (P1_U2984, P1_U5874, P1_U5875, P1_U5876, P1_U5877, P1_U5878);
  nand ginst3712 (P1_U2985, P1_U5869, P1_U5870, P1_U5871, P1_U5872, P1_U5873);
  nand ginst3713 (P1_U2986, P1_U5864, P1_U5865, P1_U5866, P1_U5867, P1_U5868);
  nand ginst3714 (P1_U2987, P1_U5859, P1_U5860, P1_U5861, P1_U5862, P1_U5863);
  nand ginst3715 (P1_U2988, P1_U5854, P1_U5855, P1_U5856, P1_U5857, P1_U5858);
  nand ginst3716 (P1_U2989, P1_U5849, P1_U5850, P1_U5851, P1_U5852, P1_U5853);
  nand ginst3717 (P1_U2990, P1_U5844, P1_U5845, P1_U5846, P1_U5847, P1_U5848);
  nand ginst3718 (P1_U2991, P1_U5839, P1_U5840, P1_U5841, P1_U5842, P1_U5843);
  nand ginst3719 (P1_U2992, P1_U5834, P1_U5835, P1_U5836, P1_U5837, P1_U5838);
  nand ginst3720 (P1_U2993, P1_U5829, P1_U5830, P1_U5831, P1_U5832, P1_U5833);
  nand ginst3721 (P1_U2994, P1_U5824, P1_U5825, P1_U5826, P1_U5827, P1_U5828);
  nand ginst3722 (P1_U2995, P1_U5819, P1_U5820, P1_U5821, P1_U5822, P1_U5823);
  nand ginst3723 (P1_U2996, P1_U5814, P1_U5815, P1_U5816, P1_U5817, P1_U5818);
  nand ginst3724 (P1_U2997, P1_U5809, P1_U5810, P1_U5811, P1_U5812, P1_U5813);
  nand ginst3725 (P1_U2998, P1_U5804, P1_U5805, P1_U5806, P1_U5807, P1_U5808);
  nand ginst3726 (P1_U2999, P1_U5799, P1_U5800, P1_U5801, P1_U5802, P1_U5803);
  nand ginst3727 (P1_U3000, P1_U3859, P1_U3861, P1_U5787, P1_U5789);
  nand ginst3728 (P1_U3001, P1_U3856, P1_U3858, P1_U5780, P1_U5782);
  nand ginst3729 (P1_U3002, P1_U3853, P1_U3855, P1_U5773, P1_U5775);
  nand ginst3730 (P1_U3003, P1_U3850, P1_U3852, P1_U5766, P1_U5768);
  nand ginst3731 (P1_U3004, P1_U3847, P1_U3849, P1_U5759, P1_U5761);
  nand ginst3732 (P1_U3005, P1_U3844, P1_U3846, P1_U5752, P1_U5754);
  nand ginst3733 (P1_U3006, P1_U3841, P1_U3843, P1_U5745, P1_U5747);
  nand ginst3734 (P1_U3007, P1_U3838, P1_U3840, P1_U5738, P1_U5740);
  nand ginst3735 (P1_U3008, P1_U3835, P1_U3837, P1_U5731, P1_U5733);
  nand ginst3736 (P1_U3009, P1_U3832, P1_U3834, P1_U5724, P1_U5726);
  nand ginst3737 (P1_U3010, P1_U3829, P1_U3831, P1_U5717, P1_U5719);
  nand ginst3738 (P1_U3011, P1_U3826, P1_U3828, P1_U5710, P1_U5712);
  nand ginst3739 (P1_U3012, P1_U3823, P1_U3825, P1_U5703, P1_U5705);
  nand ginst3740 (P1_U3013, P1_U3820, P1_U3822, P1_U5696, P1_U5698);
  nand ginst3741 (P1_U3014, P1_U3817, P1_U3819, P1_U5689, P1_U5691);
  nand ginst3742 (P1_U3015, P1_U3814, P1_U3816, P1_U5682, P1_U5684);
  nand ginst3743 (P1_U3016, P1_U3811, P1_U3813, P1_U5675, P1_U5677);
  nand ginst3744 (P1_U3017, P1_U3808, P1_U3810, P1_U5668, P1_U5670);
  nand ginst3745 (P1_U3018, P1_U3805, P1_U3807, P1_U5661, P1_U5663);
  nand ginst3746 (P1_U3019, P1_U3802, P1_U3804, P1_U5656);
  nand ginst3747 (P1_U3020, P1_U3799, P1_U3801, P1_U5649);
  nand ginst3748 (P1_U3021, P1_U3796, P1_U3798, P1_U5642);
  nand ginst3749 (P1_U3022, P1_U3793, P1_U3795, P1_U5635);
  nand ginst3750 (P1_U3023, P1_U3790, P1_U3792, P1_U5628);
  nand ginst3751 (P1_U3024, P1_U3787, P1_U3789, P1_U5621);
  nand ginst3752 (P1_U3025, P1_U3784, P1_U3786, P1_U5614);
  nand ginst3753 (P1_U3026, P1_U3781, P1_U3783, P1_U5607);
  nand ginst3754 (P1_U3027, P1_U3778, P1_U3780, P1_U5600);
  nand ginst3755 (P1_U3028, P1_U3775, P1_U3776);
  nand ginst3756 (P1_U3029, P1_U3771, P1_U3772, P1_U3774);
  nand ginst3757 (P1_U3030, P1_U3767, P1_U3768, P1_U3770);
  nand ginst3758 (P1_U3031, P1_U3763, P1_U3764, P1_U3766);
  and ginst3759 (P1_U3032, P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN, P1_U5537);
  nand ginst3760 (P1_U3033, P1_U3730, P1_U5459, P1_U5460);
  nand ginst3761 (P1_U3034, P1_U3729, P1_U5454, P1_U5455);
  nand ginst3762 (P1_U3035, P1_U3728, P1_U5449, P1_U5450);
  nand ginst3763 (P1_U3036, P1_U3727, P1_U5444, P1_U5445);
  nand ginst3764 (P1_U3037, P1_U3726, P1_U5440, P1_U7612);
  nand ginst3765 (P1_U3038, P1_U3725, P1_U5435, P1_U5436);
  nand ginst3766 (P1_U3039, P1_U3724, P1_U5430, P1_U5431);
  nand ginst3767 (P1_U3040, P1_U3723, P1_U5425, P1_U5426);
  nand ginst3768 (P1_U3041, P1_U3721, P1_U5403, P1_U5404);
  nand ginst3769 (P1_U3042, P1_U3720, P1_U5398, P1_U5399);
  nand ginst3770 (P1_U3043, P1_U3719, P1_U5393, P1_U5394);
  nand ginst3771 (P1_U3044, P1_U3718, P1_U5388, P1_U5389);
  nand ginst3772 (P1_U3045, P1_U3717, P1_U5383, P1_U5384);
  nand ginst3773 (P1_U3046, P1_U3716, P1_U5378, P1_U5379);
  nand ginst3774 (P1_U3047, P1_U3715, P1_U5373, P1_U5374);
  nand ginst3775 (P1_U3048, P1_U3714, P1_U5368, P1_U5369);
  nand ginst3776 (P1_U3049, P1_U3712, P1_U5345, P1_U5346);
  nand ginst3777 (P1_U3050, P1_U3711, P1_U5340, P1_U5341);
  nand ginst3778 (P1_U3051, P1_U3710, P1_U5335, P1_U5336);
  nand ginst3779 (P1_U3052, P1_U3709, P1_U5330, P1_U5331);
  nand ginst3780 (P1_U3053, P1_U3708, P1_U5325, P1_U5326);
  nand ginst3781 (P1_U3054, P1_U3707, P1_U5320, P1_U5321);
  nand ginst3782 (P1_U3055, P1_U3706, P1_U5315, P1_U5316);
  nand ginst3783 (P1_U3056, P1_U3705, P1_U5310, P1_U5311);
  nand ginst3784 (P1_U3057, P1_U3703, P1_U5288, P1_U5289);
  nand ginst3785 (P1_U3058, P1_U3702, P1_U5283, P1_U5284);
  nand ginst3786 (P1_U3059, P1_U3701, P1_U5278, P1_U5279);
  nand ginst3787 (P1_U3060, P1_U3700, P1_U5273, P1_U5274);
  nand ginst3788 (P1_U3061, P1_U3699, P1_U5268, P1_U5269);
  nand ginst3789 (P1_U3062, P1_U3698, P1_U5263, P1_U5264);
  nand ginst3790 (P1_U3063, P1_U3697, P1_U5258, P1_U5259);
  nand ginst3791 (P1_U3064, P1_U3696, P1_U5253, P1_U5254);
  nand ginst3792 (P1_U3065, P1_U3694, P1_U5230, P1_U5231);
  nand ginst3793 (P1_U3066, P1_U3693, P1_U5225, P1_U5226);
  nand ginst3794 (P1_U3067, P1_U3692, P1_U5220, P1_U5221);
  nand ginst3795 (P1_U3068, P1_U3691, P1_U5215, P1_U5216);
  nand ginst3796 (P1_U3069, P1_U3690, P1_U5210, P1_U5211);
  nand ginst3797 (P1_U3070, P1_U3689, P1_U5205, P1_U5206);
  nand ginst3798 (P1_U3071, P1_U3688, P1_U5200, P1_U5201);
  nand ginst3799 (P1_U3072, P1_U3687, P1_U5195, P1_U5196);
  nand ginst3800 (P1_U3073, P1_U3685, P1_U5173, P1_U5174);
  nand ginst3801 (P1_U3074, P1_U3684, P1_U5168, P1_U5169);
  nand ginst3802 (P1_U3075, P1_U3683, P1_U5163, P1_U5164);
  nand ginst3803 (P1_U3076, P1_U3682, P1_U5158, P1_U5159);
  nand ginst3804 (P1_U3077, P1_U3681, P1_U5153, P1_U5154);
  nand ginst3805 (P1_U3078, P1_U3680, P1_U5148, P1_U5149);
  nand ginst3806 (P1_U3079, P1_U3679, P1_U5143, P1_U5144);
  nand ginst3807 (P1_U3080, P1_U3678, P1_U5138, P1_U5139);
  nand ginst3808 (P1_U3081, P1_U3676, P1_U5115, P1_U5116);
  nand ginst3809 (P1_U3082, P1_U3675, P1_U5110, P1_U5111);
  nand ginst3810 (P1_U3083, P1_U3674, P1_U5105, P1_U5106);
  nand ginst3811 (P1_U3084, P1_U3673, P1_U5100, P1_U5101);
  nand ginst3812 (P1_U3085, P1_U3672, P1_U5095, P1_U5096);
  nand ginst3813 (P1_U3086, P1_U3671, P1_U5090, P1_U5091);
  nand ginst3814 (P1_U3087, P1_U3670, P1_U5085, P1_U5086);
  nand ginst3815 (P1_U3088, P1_U3669, P1_U5080, P1_U5081);
  nand ginst3816 (P1_U3089, P1_U3667, P1_U5058, P1_U5059);
  nand ginst3817 (P1_U3090, P1_U3666, P1_U5053, P1_U5054);
  nand ginst3818 (P1_U3091, P1_U3665, P1_U5048, P1_U5049);
  nand ginst3819 (P1_U3092, P1_U3664, P1_U5043, P1_U5044);
  nand ginst3820 (P1_U3093, P1_U3663, P1_U5038, P1_U5039);
  nand ginst3821 (P1_U3094, P1_U3662, P1_U5033, P1_U5034);
  nand ginst3822 (P1_U3095, P1_U3661, P1_U5028, P1_U5029);
  nand ginst3823 (P1_U3096, P1_U3660, P1_U5023, P1_U5024);
  nand ginst3824 (P1_U3097, P1_U3658, P1_U5002, P1_U5003);
  nand ginst3825 (P1_U3098, P1_U3657, P1_U4997, P1_U4998);
  nand ginst3826 (P1_U3099, P1_U3656, P1_U4992, P1_U4993);
  nand ginst3827 (P1_U3100, P1_U3655, P1_U4987, P1_U4988);
  nand ginst3828 (P1_U3101, P1_U3654, P1_U4982, P1_U4983);
  nand ginst3829 (P1_U3102, P1_U3653, P1_U4977, P1_U4978);
  nand ginst3830 (P1_U3103, P1_U3652, P1_U4972, P1_U4973);
  nand ginst3831 (P1_U3104, P1_U3651, P1_U4967, P1_U4968);
  nand ginst3832 (P1_U3105, P1_U3649, P1_U4945, P1_U4946);
  nand ginst3833 (P1_U3106, P1_U3648, P1_U4940, P1_U4941);
  nand ginst3834 (P1_U3107, P1_U3647, P1_U4935, P1_U4936);
  nand ginst3835 (P1_U3108, P1_U3646, P1_U4930, P1_U4931);
  nand ginst3836 (P1_U3109, P1_U3645, P1_U4925, P1_U4926);
  nand ginst3837 (P1_U3110, P1_U3644, P1_U4920, P1_U4921);
  nand ginst3838 (P1_U3111, P1_U3643, P1_U4915, P1_U4916);
  nand ginst3839 (P1_U3112, P1_U3642, P1_U4910, P1_U4911);
  nand ginst3840 (P1_U3113, P1_U3640, P1_U4887, P1_U4888);
  nand ginst3841 (P1_U3114, P1_U3639, P1_U4882, P1_U4883);
  nand ginst3842 (P1_U3115, P1_U3638, P1_U4877, P1_U4878);
  nand ginst3843 (P1_U3116, P1_U3637, P1_U4872, P1_U4873);
  nand ginst3844 (P1_U3117, P1_U3636, P1_U4867, P1_U4868);
  nand ginst3845 (P1_U3118, P1_U3635, P1_U4862, P1_U4863);
  nand ginst3846 (P1_U3119, P1_U3634, P1_U4857, P1_U4858);
  nand ginst3847 (P1_U3120, P1_U3633, P1_U4852, P1_U4853);
  nand ginst3848 (P1_U3121, P1_U3631, P1_U4830, P1_U4831);
  nand ginst3849 (P1_U3122, P1_U3630, P1_U4825, P1_U4826);
  nand ginst3850 (P1_U3123, P1_U3629, P1_U4820, P1_U4821);
  nand ginst3851 (P1_U3124, P1_U3628, P1_U4815, P1_U4816);
  nand ginst3852 (P1_U3125, P1_U3627, P1_U4810, P1_U4811);
  nand ginst3853 (P1_U3126, P1_U3626, P1_U4805, P1_U4806);
  nand ginst3854 (P1_U3127, P1_U3625, P1_U4800, P1_U4801);
  nand ginst3855 (P1_U3128, P1_U3624, P1_U4795, P1_U4796);
  nand ginst3856 (P1_U3129, P1_U3622, P1_U4772, P1_U4773);
  nand ginst3857 (P1_U3130, P1_U3621, P1_U4767, P1_U4768);
  nand ginst3858 (P1_U3131, P1_U3620, P1_U4762, P1_U4763);
  nand ginst3859 (P1_U3132, P1_U3619, P1_U4757, P1_U4758);
  nand ginst3860 (P1_U3133, P1_U3618, P1_U4752, P1_U4753);
  nand ginst3861 (P1_U3134, P1_U3617, P1_U4747, P1_U4748);
  nand ginst3862 (P1_U3135, P1_U3616, P1_U4742, P1_U4743);
  nand ginst3863 (P1_U3136, P1_U3615, P1_U4737, P1_U4738);
  nand ginst3864 (P1_U3137, P1_U3613, P1_U4715, P1_U4716);
  nand ginst3865 (P1_U3138, P1_U3612, P1_U4710, P1_U4711);
  nand ginst3866 (P1_U3139, P1_U3611, P1_U4705, P1_U4706);
  nand ginst3867 (P1_U3140, P1_U3610, P1_U4700, P1_U4701);
  nand ginst3868 (P1_U3141, P1_U3609, P1_U4695, P1_U4696);
  nand ginst3869 (P1_U3142, P1_U3608, P1_U4690, P1_U4691);
  nand ginst3870 (P1_U3143, P1_U3607, P1_U4685, P1_U4686);
  nand ginst3871 (P1_U3144, P1_U3606, P1_U4680, P1_U4681);
  nand ginst3872 (P1_U3145, P1_U3604, P1_U4656, P1_U4657);
  nand ginst3873 (P1_U3146, P1_U3603, P1_U4651, P1_U4652);
  nand ginst3874 (P1_U3147, P1_U3602, P1_U4646, P1_U4647);
  nand ginst3875 (P1_U3148, P1_U3601, P1_U4641, P1_U4642);
  xor ginst3876 (P1_U3149, P1_U3149_in, flip_signal);
  nand ginst3877 (P1_U3149_in, P1_U3600, P1_U4636, P1_U4637);
  nand ginst3878 (P1_U3150, P1_U3599, P1_U4631, P1_U4632);
  nand ginst3879 (P1_U3151, P1_U3598, P1_U4626, P1_U4627);
  nand ginst3880 (P1_U3152, P1_U3597, P1_U4621, P1_U4622);
  nand ginst3881 (P1_U3153, P1_U3595, P1_U4598, P1_U4599);
  nand ginst3882 (P1_U3154, P1_U3594, P1_U4593, P1_U4594);
  nand ginst3883 (P1_U3155, P1_U3593, P1_U4588, P1_U4589);
  nand ginst3884 (P1_U3156, P1_U3592, P1_U4583, P1_U4584);
  nand ginst3885 (P1_U3157, P1_U3591, P1_U4578, P1_U4579);
  nand ginst3886 (P1_U3158, P1_U3590, P1_U4573, P1_U4574);
  nand ginst3887 (P1_U3159, P1_U3589, P1_U4568, P1_U4569);
  nand ginst3888 (P1_U3160, P1_U3588, P1_U4563, P1_U4564);
  nand ginst3889 (P1_U3161, P1_U3586, P1_U7689, P1_U7690);
  nand ginst3890 (P1_U3162, P1_U4244, P1_U4518, P1_U4519, P1_U4520);
  nand ginst3891 (P1_U3163, P1_U3582, P1_U4516);
  and ginst3892 (P1_U3164, P1_DATAWIDTH_REG_31__SCAN_IN, P1_U7650);
  and ginst3893 (P1_U3165, P1_DATAWIDTH_REG_30__SCAN_IN, P1_U7650);
  and ginst3894 (P1_U3166, P1_DATAWIDTH_REG_29__SCAN_IN, P1_U7650);
  and ginst3895 (P1_U3167, P1_DATAWIDTH_REG_28__SCAN_IN, P1_U7650);
  and ginst3896 (P1_U3168, P1_DATAWIDTH_REG_27__SCAN_IN, P1_U7650);
  and ginst3897 (P1_U3169, P1_DATAWIDTH_REG_26__SCAN_IN, P1_U7650);
  and ginst3898 (P1_U3170, P1_DATAWIDTH_REG_25__SCAN_IN, P1_U7650);
  and ginst3899 (P1_U3171, P1_DATAWIDTH_REG_24__SCAN_IN, P1_U7650);
  and ginst3900 (P1_U3172, P1_DATAWIDTH_REG_23__SCAN_IN, P1_U7650);
  and ginst3901 (P1_U3173, P1_DATAWIDTH_REG_22__SCAN_IN, P1_U7650);
  and ginst3902 (P1_U3174, P1_DATAWIDTH_REG_21__SCAN_IN, P1_U7650);
  and ginst3903 (P1_U3175, P1_DATAWIDTH_REG_20__SCAN_IN, P1_U7650);
  and ginst3904 (P1_U3176, P1_DATAWIDTH_REG_19__SCAN_IN, P1_U7650);
  and ginst3905 (P1_U3177, P1_DATAWIDTH_REG_18__SCAN_IN, P1_U7650);
  and ginst3906 (P1_U3178, P1_DATAWIDTH_REG_17__SCAN_IN, P1_U7650);
  and ginst3907 (P1_U3179, P1_DATAWIDTH_REG_16__SCAN_IN, P1_U7650);
  and ginst3908 (P1_U3180, P1_DATAWIDTH_REG_15__SCAN_IN, P1_U7650);
  and ginst3909 (P1_U3181, P1_DATAWIDTH_REG_14__SCAN_IN, P1_U7650);
  and ginst3910 (P1_U3182, P1_DATAWIDTH_REG_13__SCAN_IN, P1_U7650);
  and ginst3911 (P1_U3183, P1_DATAWIDTH_REG_12__SCAN_IN, P1_U7650);
  and ginst3912 (P1_U3184, P1_DATAWIDTH_REG_11__SCAN_IN, P1_U7650);
  and ginst3913 (P1_U3185, P1_DATAWIDTH_REG_10__SCAN_IN, P1_U7650);
  and ginst3914 (P1_U3186, P1_DATAWIDTH_REG_9__SCAN_IN, P1_U7650);
  and ginst3915 (P1_U3187, P1_DATAWIDTH_REG_8__SCAN_IN, P1_U7650);
  and ginst3916 (P1_U3188, P1_DATAWIDTH_REG_7__SCAN_IN, P1_U7650);
  and ginst3917 (P1_U3189, P1_DATAWIDTH_REG_6__SCAN_IN, P1_U7650);
  and ginst3918 (P1_U3190, P1_DATAWIDTH_REG_5__SCAN_IN, P1_U7650);
  and ginst3919 (P1_U3191, P1_DATAWIDTH_REG_4__SCAN_IN, P1_U7650);
  and ginst3920 (P1_U3192, P1_DATAWIDTH_REG_3__SCAN_IN, P1_U7650);
  and ginst3921 (P1_U3193, P1_DATAWIDTH_REG_2__SCAN_IN, P1_U7650);
  nand ginst3922 (P1_U3194, P1_U4375, P1_U7646, P1_U7647);
  nand ginst3923 (P1_U3195, P1_U3495, P1_U7644, P1_U7645);
  nand ginst3924 (P1_U3196, P1_U3494, P1_U4369);
  nand ginst3925 (P1_U3197, P1_U4354, P1_U4355, P1_U4356);
  nand ginst3926 (P1_U3198, P1_U4351, P1_U4352, P1_U4353);
  nand ginst3927 (P1_U3199, P1_U4348, P1_U4349, P1_U4350);
  nand ginst3928 (P1_U3200, P1_U4345, P1_U4346, P1_U4347);
  nand ginst3929 (P1_U3201, P1_U4342, P1_U4343, P1_U4344);
  nand ginst3930 (P1_U3202, P1_U4339, P1_U4340, P1_U4341);
  nand ginst3931 (P1_U3203, P1_U4336, P1_U4337, P1_U4338);
  nand ginst3932 (P1_U3204, P1_U4333, P1_U4334, P1_U4335);
  nand ginst3933 (P1_U3205, P1_U4330, P1_U4331, P1_U4332);
  nand ginst3934 (P1_U3206, P1_U4327, P1_U4328, P1_U4329);
  nand ginst3935 (P1_U3207, P1_U4324, P1_U4325, P1_U4326);
  nand ginst3936 (P1_U3208, P1_U4321, P1_U4322, P1_U4323);
  nand ginst3937 (P1_U3209, P1_U4318, P1_U4319, P1_U4320);
  nand ginst3938 (P1_U3210, P1_U4315, P1_U4316, P1_U4317);
  nand ginst3939 (P1_U3211, P1_U4312, P1_U4313, P1_U4314);
  nand ginst3940 (P1_U3212, P1_U4309, P1_U4310, P1_U4311);
  nand ginst3941 (P1_U3213, P1_U4306, P1_U4307, P1_U4308);
  nand ginst3942 (P1_U3214, P1_U4303, P1_U4304, P1_U4305);
  nand ginst3943 (P1_U3215, P1_U4300, P1_U4301, P1_U4302);
  nand ginst3944 (P1_U3216, P1_U4297, P1_U4298, P1_U4299);
  nand ginst3945 (P1_U3217, P1_U4294, P1_U4295, P1_U4296);
  nand ginst3946 (P1_U3218, P1_U4291, P1_U4292, P1_U4293);
  nand ginst3947 (P1_U3219, P1_U4288, P1_U4289, P1_U4290);
  nand ginst3948 (P1_U3220, P1_U4285, P1_U4286, P1_U4287);
  nand ginst3949 (P1_U3221, P1_U4282, P1_U4283, P1_U4284);
  nand ginst3950 (P1_U3222, P1_U4279, P1_U4280, P1_U4281);
  nand ginst3951 (P1_U3223, P1_U4276, P1_U4277, P1_U4278);
  nand ginst3952 (P1_U3224, P1_U4273, P1_U4274, P1_U4275);
  nand ginst3953 (P1_U3225, P1_U4270, P1_U4271, P1_U4272);
  nand ginst3954 (P1_U3226, P1_U4267, P1_U4268, P1_U4269);
  nand ginst3955 (P1_U3227, P1_U3998, P1_U3999, P1_U4000, P1_U4001);
  nand ginst3956 (P1_U3228, P1_U3994, P1_U3995, P1_U3996, P1_U3997);
  nand ginst3957 (P1_U3229, P1_U3990, P1_U3991, P1_U3992, P1_U3993);
  nand ginst3958 (P1_U3230, P1_U3986, P1_U3987, P1_U3988, P1_U3989);
  nand ginst3959 (P1_U3231, P1_U3982, P1_U3983, P1_U3984, P1_U3985);
  nand ginst3960 (P1_U3232, P1_U3978, P1_U3979, P1_U3980, P1_U3981);
  nand ginst3961 (P1_U3233, P1_U3974, P1_U3975, P1_U3976, P1_U3977);
  nand ginst3962 (P1_U3234, P1_U3970, P1_U3971, P1_U3972, P1_U3973);
  nand ginst3963 (P1_U3235, P1_U3323, P1_U3329);
  nand ginst3964 (P1_U3236, P1_U2432, P1_U3235);
  nand ginst3965 (P1_U3237, P1_U2432, P1_U4543);
  nand ginst3966 (P1_U3238, P1_U2434, P1_U3235);
  nand ginst3967 (P1_U3239, P1_U2434, P1_U4543);
  nand ginst3968 (P1_U3240, P1_U2433, P1_U3235);
  nand ginst3969 (P1_U3241, P1_U2433, P1_U4543);
  nand ginst3970 (P1_U3242, P1_U2435, P1_U3235);
  nand ginst3971 (P1_U3243, P1_U2435, P1_U4543);
  nand ginst3972 (P1_U3244, P1_U3391, P1_U3394, P1_U5463);
  nand ginst3973 (P1_U3245, P1_U5464, P1_U7086);
  nand ginst3974 (P1_U3246, P1_U4156, P1_U4158, P1_U7791, P1_U7792);
  not ginst3975 (P1_U3247, P1_REQUESTPENDING_REG_SCAN_IN);
  not ginst3976 (P1_U3248, P1_STATE_REG_1__SCAN_IN);
  nand ginst3977 (P1_U3249, P1_STATE_REG_1__SCAN_IN, P1_U3258);
  nand ginst3978 (P1_U3250, P1_U3251, P1_U4221);
  not ginst3979 (P1_U3251, P1_STATE_REG_2__SCAN_IN);
  nand ginst3980 (P1_U3252, P1_STATE_REG_2__SCAN_IN, P1_U4221);
  not ginst3981 (P1_U3253, P1_REIP_REG_1__SCAN_IN);
  nand ginst3982 (P1_U3254, P1_STATE_REG_1__SCAN_IN, P1_U3251);
  or ginst3983 (P1_U3255, P1_STATE_REG_2__SCAN_IN, P1_STATE_REG_1__SCAN_IN);
  not ginst3984 (P1_U3256, HOLD);
  not ginst3985 (P1_U3257, U210);
  not ginst3986 (P1_U3258, P1_STATE_REG_0__SCAN_IN);
  nand ginst3987 (P1_U3259, P1_STATE_REG_0__SCAN_IN, P1_U3260);
  nand ginst3988 (P1_U3260, P1_REQUESTPENDING_REG_SCAN_IN, P1_U3256);
  or ginst3989 (P1_U3261, HOLD, P1_REQUESTPENDING_REG_SCAN_IN);
  not ginst3990 (P1_U3262, P1_STATE2_REG_1__SCAN_IN);
  not ginst3991 (P1_U3263, P1_STATE2_REG_2__SCAN_IN);
  not ginst3992 (P1_U3264, P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN);
  not ginst3993 (P1_U3265, P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN);
  not ginst3994 (P1_U3266, P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN);
  nand ginst3995 (P1_U3267, P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN, P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN, P1_U3270);
  or ginst3996 (P1_U3268, P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN, P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN);
  or ginst3997 (P1_U3269, P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN, P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN);
  not ginst3998 (P1_U3270, P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN);
  nand ginst3999 (P1_U3271, P1_U3564, P1_U3565, P1_U3566, P1_U3567);
  nand ginst4000 (P1_U3272, P1_U3258, P1_U4496);
  not ginst4001 (P1_U3273, P1_R2167_U17);
  nand ginst4002 (P1_U3274, P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN, P1_U3270);
  nand ginst4003 (P1_U3275, P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN, P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN);
  nand ginst4004 (P1_U3276, P1_U3516, P1_U3517, P1_U3518, P1_U3519);
  nand ginst4005 (P1_U3277, P1_U3536, P1_U3537, P1_U3538, P1_U3539, P1_U4170);
  nand ginst4006 (P1_U3278, P1_U3554, P1_U3555, P1_U3556, P1_U3557);
  nand ginst4007 (P1_U3279, P1_U3558, P1_U3559);
  or ginst4008 (P1_U3280, P1_STATEBS16_REG_SCAN_IN, U210);
  nand ginst4009 (P1_U3281, P1_R2167_U17, P1_U4497);
  nand ginst4010 (P1_U3282, P1_U3284, P1_U4477);
  nand ginst4011 (P1_U3283, P1_U3508, P1_U3509, P1_U3510, P1_U3511);
  nand ginst4012 (P1_U3284, P1_U3560, P1_U3561, P1_U3562, P1_U3563);
  nand ginst4013 (P1_U3285, P1_U2473, P1_U4501);
  nand ginst4014 (P1_U3286, P1_U2389, P1_U3283);
  nand ginst4015 (P1_U3287, P1_U4477, P1_U4494);
  nand ginst4016 (P1_U3288, P1_U2447, P1_U4249);
  nand ginst4017 (P1_U3289, P1_U3278, P1_U3391, P1_U4173, P1_U4460);
  nand ginst4018 (P1_U3290, P1_U3271, P1_U3283);
  nand ginst4019 (P1_U3291, P1_U3284, P1_U4190);
  nand ginst4020 (P1_U3292, P1_U2431, P1_U4256);
  nand ginst4021 (P1_U3293, P1_LT_563_U6, P1_U4178, P1_U4225, P1_U4509, P1_U7626);
  not ginst4022 (P1_U3294, P1_STATE2_REG_0__SCAN_IN);
  nand ginst4023 (P1_U3295, P1_STATE2_REG_0__SCAN_IN, P1_U7604);
  not ginst4024 (P1_U3296, P1_STATE2_REG_3__SCAN_IN);
  nand ginst4025 (P1_U3297, P1_STATE2_REG_2__SCAN_IN, P1_U3262);
  or ginst4026 (P1_U3298, P1_STATE2_REG_2__SCAN_IN, P1_STATE2_REG_1__SCAN_IN);
  nand ginst4027 (P1_U3299, P1_STATE2_REG_3__SCAN_IN, P1_R2167_U17);
  nand ginst4028 (P1_U3300, P1_U3294, P1_U4547);
  not ginst4029 (P1_U3301, P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN);
  not ginst4030 (P1_U3302, P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN);
  not ginst4031 (P1_U3303, P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN);
  not ginst4032 (P1_U3304, P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN);
  nand ginst4033 (P1_U3305, P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN);
  nand ginst4034 (P1_U3306, P1_U2478, P1_U4533);
  or ginst4035 (P1_U3307, P1_STATE2_REG_3__SCAN_IN, P1_STATE2_REG_2__SCAN_IN);
  not ginst4036 (P1_U3308, P1_STATEBS16_REG_SCAN_IN);
  not ginst4037 (P1_U3309, P1_R2144_U43);
  not ginst4038 (P1_U3310, P1_R2144_U50);
  not ginst4039 (P1_U3311, P1_R2144_U49);
  not ginst4040 (P1_U3312, P1_R2144_U8);
  nand ginst4041 (P1_U3313, P1_R2144_U43, P1_R2144_U50);
  nand ginst4042 (P1_U3314, P1_U3309, P1_U3332);
  nand ginst4043 (P1_U3315, P1_U2475, P1_U4527);
  not ginst4044 (P1_U3316, P1_R2182_U25);
  not ginst4045 (P1_U3317, P1_R2182_U42);
  not ginst4046 (P1_U3318, P1_R2182_U34);
  not ginst4047 (P1_U3319, P1_R2182_U33);
  nand ginst4048 (P1_U3320, P1_U3308, P1_U4209);
  nand ginst4049 (P1_U3321, P1_U3306, P1_U4535);
  nand ginst4050 (P1_U3322, P1_U3306, P1_U4544);
  nand ginst4051 (P1_U3323, P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN, P1_U3301);
  nand ginst4052 (P1_U3324, P1_U2478, P1_U4542);
  nand ginst4053 (P1_U3325, P1_R2144_U50, P1_U3309);
  nand ginst4054 (P1_U3326, P1_R2144_U43, P1_U3332);
  nand ginst4055 (P1_U3327, P1_U2475, P1_U4600);
  nand ginst4056 (P1_U3328, P1_U3324, P1_U4603);
  nand ginst4057 (P1_U3329, P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P1_U3302);
  nand ginst4058 (P1_U3330, P1_U2478, P1_U4541);
  nand ginst4059 (P1_U3331, P1_R2144_U43, P1_U3310);
  nand ginst4060 (P1_U3332, P1_U3325, P1_U3331);
  nand ginst4061 (P1_U3333, P1_U3309, P1_U4526);
  nand ginst4062 (P1_U3334, P1_U2475, P1_U4658);
  nand ginst4063 (P1_U3335, P1_U3330, P1_U4661);
  nand ginst4064 (P1_U3336, P1_U3330, P1_U4663);
  nand ginst4065 (P1_U3337, P1_U2478, P1_U2488);
  nand ginst4066 (P1_U3338, P1_U2475, P1_U2485);
  nand ginst4067 (P1_U3339, P1_U3337, P1_U4719);
  nand ginst4068 (P1_U3340, P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN, P1_U3304);
  nand ginst4069 (P1_U3341, P1_U4533, P1_U4538);
  nand ginst4070 (P1_U3342, P1_R2144_U8, P1_U3311);
  nand ginst4071 (P1_U3343, P1_U2490, P1_U4527);
  nand ginst4072 (P1_U3344, P1_U3341, P1_U4776);
  nand ginst4073 (P1_U3345, P1_U3341, P1_U4778);
  nand ginst4074 (P1_U3346, P1_U4538, P1_U4542);
  nand ginst4075 (P1_U3347, P1_U2490, P1_U4600);
  nand ginst4076 (P1_U3348, P1_U3346, P1_U4834);
  nand ginst4077 (P1_U3349, P1_U4538, P1_U4541);
  nand ginst4078 (P1_U3350, P1_U2490, P1_U4658);
  nand ginst4079 (P1_U3351, P1_U3349, P1_U4891);
  nand ginst4080 (P1_U3352, P1_U3349, P1_U4893);
  nand ginst4081 (P1_U3353, P1_U2488, P1_U4538);
  nand ginst4082 (P1_U3354, P1_U2485, P1_U2490);
  nand ginst4083 (P1_U3355, P1_U3353, P1_U4949);
  nand ginst4084 (P1_U3356, P1_U2479, P1_U4533);
  nand ginst4085 (P1_U3357, P1_U2474, P1_U4528);
  nand ginst4086 (P1_U3358, P1_U3342, P1_U3357, P1_U4530);
  nand ginst4087 (P1_U3359, P1_U2499, P1_U4527);
  nand ginst4088 (P1_U3360, P1_U3340, P1_U3356, P1_U4539);
  nand ginst4089 (P1_U3361, P1_U3356, P1_U5005);
  nand ginst4090 (P1_U3362, P1_U3356, P1_U5007);
  nand ginst4091 (P1_U3363, P1_U2479, P1_U4542);
  nand ginst4092 (P1_U3364, P1_U2499, P1_U4600);
  nand ginst4093 (P1_U3365, P1_U3363, P1_U5062);
  nand ginst4094 (P1_U3366, P1_U2479, P1_U4541);
  nand ginst4095 (P1_U3367, P1_U2499, P1_U4658);
  nand ginst4096 (P1_U3368, P1_U3366, P1_U5119);
  nand ginst4097 (P1_U3369, P1_U3366, P1_U5121);
  nand ginst4098 (P1_U3370, P1_U2479, P1_U2488);
  nand ginst4099 (P1_U3371, P1_U2485, P1_U2499);
  nand ginst4100 (P1_U3372, P1_U3370, P1_U5177);
  nand ginst4101 (P1_U3373, P1_U2510, P1_U4533);
  nand ginst4102 (P1_U3374, P1_U2507, P1_U4527);
  nand ginst4103 (P1_U3375, P1_U3373, P1_U5234);
  nand ginst4104 (P1_U3376, P1_U3373, P1_U5236);
  nand ginst4105 (P1_U3377, P1_U2510, P1_U4542);
  nand ginst4106 (P1_U3378, P1_U2507, P1_U4600);
  nand ginst4107 (P1_U3379, P1_U3377, P1_U5292);
  nand ginst4108 (P1_U3380, P1_U2510, P1_U4541);
  nand ginst4109 (P1_U3381, P1_U2507, P1_U4658);
  nand ginst4110 (P1_U3382, P1_U3380, P1_U5349);
  nand ginst4111 (P1_U3383, P1_U3380, P1_U5351);
  nand ginst4112 (P1_U3384, P1_U2488, P1_U2510);
  nand ginst4113 (P1_U3385, P1_U2485, P1_U2507);
  nand ginst4114 (P1_U3386, P1_U3384, P1_U5407);
  not ginst4115 (P1_U3387, P1_FLUSH_REG_SCAN_IN);
  not ginst4116 (P1_U3388, P1_GTE_485_U6);
  nand ginst4117 (P1_U3389, P1_U3278, P1_U3284);
  nand ginst4118 (P1_U3390, P1_U3271, P1_U3284);
  nand ginst4119 (P1_U3391, P1_U3512, P1_U3513, P1_U3514, P1_U3515);
  nand ginst4120 (P1_U3392, P1_U5489, P1_U5490, P1_U7628);
  nand ginst4121 (P1_U3393, P1_U3284, P1_U4399);
  nand ginst4122 (P1_U3394, P1_U2605, P1_U3277);
  nand ginst4123 (P1_U3395, P1_U4399, P1_U4494, P1_U7494);
  nand ginst4124 (P1_U3396, P1_U3741, P1_U4247);
  nand ginst4125 (P1_U3397, P1_U2605, P1_U4399, P1_U4477, P1_U4494, P1_U7494);
  nand ginst4126 (P1_U3398, P1_U2605, P1_U4171, P1_U4400, P1_U4449, P1_U4460);
  nand ginst4127 (P1_U3399, P1_U4199, P1_U4234, P1_U4477);
  nand ginst4128 (P1_U3400, P1_U2447, P1_U2449);
  nand ginst4129 (P1_U3401, P1_U3444, P1_U5510);
  nand ginst4130 (P1_U3402, P1_U3269, P1_U3275);
  not ginst4131 (P1_U3403, P1_LT_589_U6);
  nand ginst4132 (P1_U3404, P1_U3300, P1_U4242, P1_U5536);
  nand ginst4133 (P1_U3405, P1_STATE2_REG_0__SCAN_IN, P1_U3278, P1_U3284);
  nand ginst4134 (P1_U3406, P1_U3271, P1_U3273);
  nand ginst4135 (P1_U3407, P1_U3277, P1_U3391);
  nand ginst4136 (P1_U3408, P1_U2427, P1_U3294);
  nand ginst4137 (P1_U3409, P1_U3391, P1_U4460);
  nand ginst4138 (P1_U3410, P1_U3278, P1_U4253);
  nand ginst4139 (P1_U3411, P1_U2452, P1_U4190);
  nand ginst4140 (P1_U3412, P1_STATE2_REG_2__SCAN_IN, P1_U3271);
  not ginst4141 (P1_U3413, P1_REIP_REG_0__SCAN_IN);
  nand ginst4142 (P1_U3414, P1_U3756, P1_U5562);
  nand ginst4143 (P1_U3415, P1_U4173, P1_U4400);
  nand ginst4144 (P1_U3416, P1_U3863, P1_U4248);
  nand ginst4145 (P1_U3417, P1_U6053, P1_U6054);
  nand ginst4146 (P1_U3418, P1_STATE2_REG_0__SCAN_IN, P1_U4494);
  nand ginst4147 (P1_U3419, P1_U4399, P1_U7494);
  nand ginst4148 (P1_U3420, P1_U4206, P1_U4477);
  nand ginst4149 (P1_U3421, P1_U2431, P1_U4194);
  nand ginst4150 (P1_U3422, P1_STATE2_REG_0__SCAN_IN, P1_U4210);
  nand ginst4151 (P1_U3423, P1_U3391, P1_U4503);
  nand ginst4152 (P1_U3424, P1_U4235, P1_U6153);
  nand ginst4153 (P1_U3425, P1_STATE2_REG_0__SCAN_IN, P1_U4216);
  nand ginst4154 (P1_U3426, P1_U4235, P1_U6264);
  nand ginst4155 (P1_U3427, P1_STATE2_REG_0__SCAN_IN, P1_U2452, P1_U3886, P1_U4249);
  nand ginst4156 (P1_U3428, P1_U2447, P1_U3866);
  not ginst4157 (P1_U3429, P1_EBX_REG_31__SCAN_IN);
  not ginst4158 (P1_U3430, P1_R2337_U69);
  nand ginst4159 (P1_U3431, P1_U3887, P1_U4228);
  nand ginst4160 (P1_U3432, P1_U3262, P1_U4209);
  nand ginst4161 (P1_U3433, P1_U3952, P1_U3955, P1_U3958, P1_U3962);
  nand ginst4162 (P1_U3434, P1_U3271, P1_U4206);
  not ginst4163 (P1_U3435, P1_CODEFETCH_REG_SCAN_IN);
  not ginst4164 (P1_U3436, P1_READREQUEST_REG_SCAN_IN);
  nand ginst4165 (P1_U3437, P1_U2447, P1_U4498);
  nand ginst4166 (P1_U3438, P1_U3267, P1_U5482);
  nand ginst4167 (P1_U3439, P1_STATE2_REG_2__SCAN_IN, P1_U4449);
  nand ginst4168 (P1_U3440, P1_STATEBS16_REG_SCAN_IN, P1_U3263);
  not ginst4169 (P1_U3441, P1_U3234);
  nand ginst4170 (P1_U3442, P1_U5478, P1_U5479);
  nand ginst4171 (P1_U3443, P1_U2450, P1_U3441);
  nand ginst4172 (P1_U3444, P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN, P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P1_U3264);
  nand ginst4173 (P1_U3445, P1_U3274, P1_U7064);
  nand ginst4174 (P1_U3446, P1_U4197, P1_U4234);
  nand ginst4175 (P1_U3447, P1_U4231, P1_U4250, P1_U4400);
  nand ginst4176 (P1_U3448, P1_U3278, P1_U4231, P1_U4250);
  nand ginst4177 (P1_U3449, P1_U4477, P1_U4496);
  nand ginst4178 (P1_U3450, P1_U4074, P1_U4075, P1_U4077, P1_U7093);
  nand ginst4179 (P1_U3451, P1_U4254, P1_U4266);
  nand ginst4180 (P1_U3452, P1_U3268, P1_U4183);
  nand ginst4181 (P1_U3453, P1_STATE2_REG_0__SCAN_IN, P1_U2605);
  nand ginst4182 (P1_U3454, P1_U7691, P1_U7692);
  nand ginst4183 (P1_U3455, P1_U7694, P1_U7695);
  nand ginst4184 (P1_U3456, P1_U7718, P1_U7719);
  nand ginst4185 (P1_U3457, P1_U7788, P1_U7789);
  nand ginst4186 (P1_U3458, P1_U7633, P1_U7634);
  nand ginst4187 (P1_U3459, P1_U7635, P1_U7636);
  nand ginst4188 (P1_U3460, P1_U7637, P1_U7638);
  nand ginst4189 (P1_U3461, P1_U7639, P1_U7640);
  nand ginst4190 (P1_U3462, P1_U7648, P1_U7649);
  and ginst4191 (P1_U3463, P1_U3255, P1_U4179);
  nand ginst4192 (P1_U3464, P1_U7651, P1_U7652);
  nand ginst4193 (P1_U3465, P1_U7653, P1_U7654);
  nand ginst4194 (P1_U3466, P1_U7685, P1_U7686);
  and ginst4195 (P1_U3467, P1_R2182_U24, P1_U2427, P1_U4215);
  nand ginst4196 (P1_U3468, P1_U7701, P1_U7702);
  nand ginst4197 (P1_U3469, P1_U7708, P1_U7709);
  nand ginst4198 (P1_U3470, P1_U7710, P1_U7711);
  nand ginst4199 (P1_U3471, P1_U7713, P1_U7714);
  nand ginst4200 (P1_U3472, P1_U7721, P1_U7722);
  nand ginst4201 (P1_U3473, P1_U7723, P1_U7724);
  nand ginst4202 (P1_U3474, P1_U7727, P1_U7728);
  nand ginst4203 (P1_U3475, P1_U7729, P1_U7730);
  nand ginst4204 (P1_U3476, P1_U7734, P1_U7735);
  nand ginst4205 (P1_U3477, P1_U7736, P1_U7737);
  nand ginst4206 (P1_U3478, P1_U7738, P1_U7739);
  and ginst4207 (P1_U3479, P1_R2358_U22, P1_U4449);
  nor ginst4208 (P1_U3480, P1_REIP_REG_1__SCAN_IN, P1_DATAWIDTH_REG_1__SCAN_IN);
  nand ginst4209 (P1_U3481, P1_U7754, P1_U7755);
  nand ginst4210 (P1_U3482, P1_U7758, P1_U7759);
  nand ginst4211 (P1_U3483, P1_U7760, P1_U7761);
  nand ginst4212 (P1_U3484, P1_U7762, P1_U7763);
  nand ginst4213 (P1_U3485, P1_U7766, P1_U7767);
  nand ginst4214 (P1_U3486, P1_U7770, P1_U7771);
  nand ginst4215 (P1_U3487, P1_U7772, P1_U7773);
  and ginst4216 (P1_U3488, P1_R2182_U24, P1_U4215);
  nand ginst4217 (P1_U3489, P1_U7774, P1_U7775);
  nand ginst4218 (P1_U3490, P1_U7776, P1_U7777);
  nand ginst4219 (P1_U3491, P1_U7778, P1_U7779);
  nand ginst4220 (P1_U3492, P1_U7780, P1_U7781);
  nand ginst4221 (P1_U3493, P1_U7782, P1_U7783);
  and ginst4222 (P1_U3494, P1_U3252, P1_U4368);
  and ginst4223 (P1_U3495, P1_U3250, P1_U4370);
  and ginst4224 (P1_U3496, P1_REQUESTPENDING_REG_SCAN_IN, P1_STATE_REG_0__SCAN_IN);
  nor ginst4225 (P1_U3497, P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN, P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN);
  and ginst4226 (P1_U3498, P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN, P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN);
  nor ginst4227 (P1_U3499, P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN);
  and ginst4228 (P1_U3500, P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN, P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN);
  nor ginst4229 (P1_U3501, P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN, P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN);
  and ginst4230 (P1_U3502, P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN);
  nor ginst4231 (P1_U3503, P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN);
  and ginst4232 (P1_U3504, P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN, P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN);
  nor ginst4233 (P1_U3505, P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN, P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN);
  and ginst4234 (P1_U3506, P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN);
  and ginst4235 (P1_U3507, P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN, P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN);
  and ginst4236 (P1_U3508, P1_U4383, P1_U4384, P1_U4385, P1_U4386);
  and ginst4237 (P1_U3509, P1_U4387, P1_U4388, P1_U4389, P1_U4390);
  and ginst4238 (P1_U3510, P1_U4391, P1_U4392, P1_U4393, P1_U4394);
  and ginst4239 (P1_U3511, P1_U4395, P1_U4396, P1_U4397, P1_U4398);
  and ginst4240 (P1_U3512, P1_U4433, P1_U4434, P1_U4435, P1_U4436);
  and ginst4241 (P1_U3513, P1_U4437, P1_U4438, P1_U4439, P1_U4440);
  and ginst4242 (P1_U3514, P1_U4441, P1_U4442, P1_U4443, P1_U4444);
  and ginst4243 (P1_U3515, P1_U4445, P1_U4446, P1_U4447, P1_U4448);
  and ginst4244 (P1_U3516, P1_U4416, P1_U4417, P1_U4418, P1_U4419);
  and ginst4245 (P1_U3517, P1_U4420, P1_U4421, P1_U4422, P1_U4423);
  and ginst4246 (P1_U3518, P1_U4424, P1_U4425, P1_U4426, P1_U4427);
  and ginst4247 (P1_U3519, P1_U4428, P1_U4429, P1_U4430, P1_U4431);
  nor ginst4248 (P1_U3520, P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN);
  and ginst4249 (P1_U3521, P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN, P1_INSTQUEUE_REG_5__5__SCAN_IN);
  nor ginst4250 (P1_U3522, P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN, P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN);
  and ginst4251 (P1_U3523, P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P1_INSTQUEUE_REG_6__5__SCAN_IN);
  and ginst4252 (P1_U3524, P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P1_INSTQUEUE_REG_8__5__SCAN_IN);
  nor ginst4253 (P1_U3525, P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN, P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN);
  and ginst4254 (P1_U3526, P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P1_INSTQUEUE_REG_10__5__SCAN_IN);
  and ginst4255 (P1_U3527, P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P1_INSTQUEUE_REG_12__5__SCAN_IN);
  nor ginst4256 (P1_U3528, P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN);
  and ginst4257 (P1_U3529, P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN, P1_INSTQUEUE_REG_9__5__SCAN_IN);
  and ginst4258 (P1_U3530, P1_U4401, P1_U4402, P1_U4403, P1_U4404);
  and ginst4259 (P1_U3531, P1_U4405, P1_U4406, P1_U4407, P1_U4408);
  and ginst4260 (P1_U3532, P1_U4409, P1_U4410, P1_U4411, P1_U4412);
  and ginst4261 (P1_U3533, P1_U4413, P1_U4414);
  nor ginst4262 (P1_U3534, P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN, P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN);
  and ginst4263 (P1_U3535, P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN, P1_INSTQUEUE_REG_3__6__SCAN_IN);
  and ginst4264 (P1_U3536, P1_U4450, P1_U4451, P1_U4452, P1_U4453);
  and ginst4265 (P1_U3537, P1_U4454, P1_U4455, P1_U4456);
  and ginst4266 (P1_U3538, P1_U4457, P1_U4458, P1_U4459);
  and ginst4267 (P1_U3539, P1_U7675, P1_U7676, P1_U7677, P1_U7678);
  nor ginst4268 (P1_U3540, P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN, P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN);
  and ginst4269 (P1_U3541, P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN, P1_INSTQUEUE_REG_1__4__SCAN_IN);
  nor ginst4270 (P1_U3542, P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN, P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN);
  and ginst4271 (P1_U3543, P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN, P1_INSTQUEUE_REG_4__4__SCAN_IN);
  nor ginst4272 (P1_U3544, P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN, P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN);
  and ginst4273 (P1_U3545, P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN, P1_INSTQUEUE_REG_12__4__SCAN_IN);
  and ginst4274 (P1_U3546, P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN, P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN);
  and ginst4275 (P1_U3547, P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P1_INSTQUEUE_REG_13__4__SCAN_IN);
  nor ginst4276 (P1_U3548, P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN, P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN);
  and ginst4277 (P1_U3549, P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN, P1_INSTQUEUE_REG_6__4__SCAN_IN);
  and ginst4278 (P1_U3550, P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN);
  and ginst4279 (P1_U3551, P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P1_INSTQUEUE_REG_14__4__SCAN_IN);
  nor ginst4280 (P1_U3552, P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN);
  and ginst4281 (P1_U3553, P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P1_INSTQUEUE_REG_9__4__SCAN_IN);
  and ginst4282 (P1_U3554, P1_U7655, P1_U7656, P1_U7657, P1_U7658);
  and ginst4283 (P1_U3555, P1_U7659, P1_U7660, P1_U7661, P1_U7662);
  and ginst4284 (P1_U3556, P1_U7663, P1_U7664, P1_U7665, P1_U7666);
  and ginst4285 (P1_U3557, P1_U7667, P1_U7668, P1_U7669, P1_U7670);
  and ginst4286 (P1_U3558, P1_U3283, P1_U3391, P1_U7494);
  and ginst4287 (P1_U3559, P1_U2605, P1_U4400, P1_U4460);
  and ginst4288 (P1_U3560, P1_U4478, P1_U4479, P1_U4480, P1_U4481);
  and ginst4289 (P1_U3561, P1_U4482, P1_U4483, P1_U4484, P1_U4485);
  and ginst4290 (P1_U3562, P1_U4486, P1_U4487, P1_U4488, P1_U4489);
  and ginst4291 (P1_U3563, P1_U4490, P1_U4491, P1_U4492, P1_U4493);
  and ginst4292 (P1_U3564, P1_U4461, P1_U4462, P1_U4463, P1_U4464);
  and ginst4293 (P1_U3565, P1_U4465, P1_U4466, P1_U4467, P1_U4468);
  and ginst4294 (P1_U3566, P1_U4469, P1_U4470, P1_U4471, P1_U4472);
  and ginst4295 (P1_U3567, P1_U4473, P1_U4474, P1_U4475, P1_U4476);
  and ginst4296 (P1_U3568, P1_U4208, P1_U4377);
  and ginst4297 (P1_U3569, P1_U4416, P1_U4417, P1_U4418, P1_U4419);
  and ginst4298 (P1_U3570, P1_U4420, P1_U4421, P1_U4422, P1_U4423);
  and ginst4299 (P1_U3571, P1_U4424, P1_U4425, P1_U4426, P1_U4427);
  and ginst4300 (P1_U3572, P1_U4428, P1_U4429, P1_U4430, P1_U4431);
  and ginst4301 (P1_U3573, P1_U4401, P1_U4402, P1_U4403, P1_U4404);
  and ginst4302 (P1_U3574, P1_U4405, P1_U4406, P1_U4407, P1_U4408);
  and ginst4303 (P1_U3575, P1_U4409, P1_U4410, P1_U4411, P1_U4412);
  and ginst4304 (P1_U3576, P1_U4413, P1_U4414);
  and ginst4305 (P1_U3577, P1_U4171, P1_U4399);
  and ginst4306 (P1_U3578, P1_U3283, P1_U4249);
  and ginst4307 (P1_U3579, P1_U3283, P1_U3284, P1_U4400, P1_U7494);
  and ginst4308 (P1_U3580, P1_U3400, P1_U4217);
  and ginst4309 (P1_U3581, P1_STATE2_REG_2__SCAN_IN, P1_U7603);
  and ginst4310 (P1_U3582, P1_U3297, P1_U4515);
  and ginst4311 (P1_U3583, P1_U2427, P1_U3257);
  and ginst4312 (P1_U3584, P1_STATE2_REG_3__SCAN_IN, P1_STATE2_REG_0__SCAN_IN);
  and ginst4313 (P1_U3585, P1_U4241, P1_U4246);
  and ginst4314 (P1_U3586, P1_U3585, P1_U4523);
  and ginst4315 (P1_U3587, P1_U4224, P1_U4552, P1_U4553);
  and ginst4316 (P1_U3588, P1_U4560, P1_U4561, P1_U4562);
  and ginst4317 (P1_U3589, P1_U4565, P1_U4566, P1_U4567);
  and ginst4318 (P1_U3590, P1_U4570, P1_U4571, P1_U4572);
  and ginst4319 (P1_U3591, P1_U4575, P1_U4576, P1_U4577);
  and ginst4320 (P1_U3592, P1_U4580, P1_U4581, P1_U4582);
  and ginst4321 (P1_U3593, P1_U4585, P1_U4586, P1_U4587);
  and ginst4322 (P1_U3594, P1_U4590, P1_U4591, P1_U4592);
  and ginst4323 (P1_U3595, P1_U4595, P1_U4596, P1_U4597);
  and ginst4324 (P1_U3596, P1_U4224, P1_U4610, P1_U4611);
  and ginst4325 (P1_U3597, P1_U4618, P1_U4619, P1_U4620);
  and ginst4326 (P1_U3598, P1_U4623, P1_U4624, P1_U4625);
  and ginst4327 (P1_U3599, P1_U4628, P1_U4629, P1_U4630);
  and ginst4328 (P1_U3600, P1_U4633, P1_U4634, P1_U4635);
  and ginst4329 (P1_U3601, P1_U4638, P1_U4639, P1_U4640);
  and ginst4330 (P1_U3602, P1_U4643, P1_U4644, P1_U4645);
  and ginst4331 (P1_U3603, P1_U4648, P1_U4649, P1_U4650);
  and ginst4332 (P1_U3604, P1_U4653, P1_U4654, P1_U4655);
  and ginst4333 (P1_U3605, P1_U4224, P1_U4669, P1_U4670);
  and ginst4334 (P1_U3606, P1_U4677, P1_U4678, P1_U4679);
  and ginst4335 (P1_U3607, P1_U4682, P1_U4683, P1_U4684);
  and ginst4336 (P1_U3608, P1_U4687, P1_U4688, P1_U4689);
  and ginst4337 (P1_U3609, P1_U4692, P1_U4693, P1_U4694);
  and ginst4338 (P1_U3610, P1_U4697, P1_U4698, P1_U4699);
  and ginst4339 (P1_U3611, P1_U4702, P1_U4703, P1_U4704);
  and ginst4340 (P1_U3612, P1_U4707, P1_U4708, P1_U4709);
  and ginst4341 (P1_U3613, P1_U4712, P1_U4713, P1_U4714);
  and ginst4342 (P1_U3614, P1_U4224, P1_U4726, P1_U4727);
  and ginst4343 (P1_U3615, P1_U4734, P1_U4735, P1_U4736);
  and ginst4344 (P1_U3616, P1_U4739, P1_U4740, P1_U4741);
  and ginst4345 (P1_U3617, P1_U4744, P1_U4745, P1_U4746);
  and ginst4346 (P1_U3618, P1_U4749, P1_U4750, P1_U4751);
  and ginst4347 (P1_U3619, P1_U4754, P1_U4755, P1_U4756);
  and ginst4348 (P1_U3620, P1_U4759, P1_U4760, P1_U4761);
  and ginst4349 (P1_U3621, P1_U4764, P1_U4765, P1_U4766);
  and ginst4350 (P1_U3622, P1_U4769, P1_U4770, P1_U4771);
  and ginst4351 (P1_U3623, P1_U4224, P1_U4784, P1_U4785);
  and ginst4352 (P1_U3624, P1_U4792, P1_U4793, P1_U4794);
  and ginst4353 (P1_U3625, P1_U4797, P1_U4798, P1_U4799);
  and ginst4354 (P1_U3626, P1_U4802, P1_U4803, P1_U4804);
  and ginst4355 (P1_U3627, P1_U4807, P1_U4808, P1_U4809);
  and ginst4356 (P1_U3628, P1_U4812, P1_U4813, P1_U4814);
  and ginst4357 (P1_U3629, P1_U4817, P1_U4818, P1_U4819);
  and ginst4358 (P1_U3630, P1_U4822, P1_U4823, P1_U4824);
  and ginst4359 (P1_U3631, P1_U4827, P1_U4828, P1_U4829);
  and ginst4360 (P1_U3632, P1_U4224, P1_U4841, P1_U4842);
  and ginst4361 (P1_U3633, P1_U4849, P1_U4850, P1_U4851);
  and ginst4362 (P1_U3634, P1_U4854, P1_U4855, P1_U4856);
  and ginst4363 (P1_U3635, P1_U4859, P1_U4860, P1_U4861);
  and ginst4364 (P1_U3636, P1_U4864, P1_U4865, P1_U4866);
  and ginst4365 (P1_U3637, P1_U4869, P1_U4870, P1_U4871);
  and ginst4366 (P1_U3638, P1_U4874, P1_U4875, P1_U4876);
  and ginst4367 (P1_U3639, P1_U4879, P1_U4880, P1_U4881);
  and ginst4368 (P1_U3640, P1_U4884, P1_U4885, P1_U4886);
  and ginst4369 (P1_U3641, P1_U4224, P1_U4899, P1_U4900);
  and ginst4370 (P1_U3642, P1_U4907, P1_U4908, P1_U4909);
  and ginst4371 (P1_U3643, P1_U4912, P1_U4913, P1_U4914);
  and ginst4372 (P1_U3644, P1_U4917, P1_U4918, P1_U4919);
  and ginst4373 (P1_U3645, P1_U4922, P1_U4923, P1_U4924);
  and ginst4374 (P1_U3646, P1_U4927, P1_U4928, P1_U4929);
  and ginst4375 (P1_U3647, P1_U4932, P1_U4933, P1_U4934);
  and ginst4376 (P1_U3648, P1_U4937, P1_U4938, P1_U4939);
  and ginst4377 (P1_U3649, P1_U4942, P1_U4943, P1_U4944);
  and ginst4378 (P1_U3650, P1_U4224, P1_U4956, P1_U4957);
  and ginst4379 (P1_U3651, P1_U4964, P1_U4965, P1_U4966);
  and ginst4380 (P1_U3652, P1_U4969, P1_U4970, P1_U4971);
  and ginst4381 (P1_U3653, P1_U4974, P1_U4975, P1_U4976);
  and ginst4382 (P1_U3654, P1_U4979, P1_U4980, P1_U4981);
  and ginst4383 (P1_U3655, P1_U4984, P1_U4985, P1_U4986);
  and ginst4384 (P1_U3656, P1_U4989, P1_U4990, P1_U4991);
  and ginst4385 (P1_U3657, P1_U4994, P1_U4995, P1_U4996);
  and ginst4386 (P1_U3658, P1_U4999, P1_U5000, P1_U5001);
  and ginst4387 (P1_U3659, P1_U4224, P1_U5012, P1_U5013);
  and ginst4388 (P1_U3660, P1_U5020, P1_U5021, P1_U5022);
  and ginst4389 (P1_U3661, P1_U5025, P1_U5026, P1_U5027);
  and ginst4390 (P1_U3662, P1_U5030, P1_U5031, P1_U5032);
  and ginst4391 (P1_U3663, P1_U5035, P1_U5036, P1_U5037);
  and ginst4392 (P1_U3664, P1_U5040, P1_U5041, P1_U5042);
  and ginst4393 (P1_U3665, P1_U5045, P1_U5046, P1_U5047);
  and ginst4394 (P1_U3666, P1_U5050, P1_U5051, P1_U5052);
  and ginst4395 (P1_U3667, P1_U5055, P1_U5056, P1_U5057);
  and ginst4396 (P1_U3668, P1_U4224, P1_U5069, P1_U5070);
  and ginst4397 (P1_U3669, P1_U5077, P1_U5078, P1_U5079);
  and ginst4398 (P1_U3670, P1_U5082, P1_U5083, P1_U5084);
  and ginst4399 (P1_U3671, P1_U5087, P1_U5088, P1_U5089);
  and ginst4400 (P1_U3672, P1_U5092, P1_U5093, P1_U5094);
  and ginst4401 (P1_U3673, P1_U5097, P1_U5098, P1_U5099);
  and ginst4402 (P1_U3674, P1_U5102, P1_U5103, P1_U5104);
  and ginst4403 (P1_U3675, P1_U5107, P1_U5108, P1_U5109);
  and ginst4404 (P1_U3676, P1_U5112, P1_U5113, P1_U5114);
  and ginst4405 (P1_U3677, P1_U4224, P1_U5127, P1_U5128);
  and ginst4406 (P1_U3678, P1_U5135, P1_U5136, P1_U5137);
  and ginst4407 (P1_U3679, P1_U5140, P1_U5141, P1_U5142);
  and ginst4408 (P1_U3680, P1_U5145, P1_U5146, P1_U5147);
  and ginst4409 (P1_U3681, P1_U5150, P1_U5151, P1_U5152);
  and ginst4410 (P1_U3682, P1_U5155, P1_U5156, P1_U5157);
  and ginst4411 (P1_U3683, P1_U5160, P1_U5161, P1_U5162);
  and ginst4412 (P1_U3684, P1_U5165, P1_U5166, P1_U5167);
  and ginst4413 (P1_U3685, P1_U5170, P1_U5171, P1_U5172);
  and ginst4414 (P1_U3686, P1_U4224, P1_U5184, P1_U5185);
  and ginst4415 (P1_U3687, P1_U5192, P1_U5193, P1_U5194);
  and ginst4416 (P1_U3688, P1_U5197, P1_U5198, P1_U5199);
  and ginst4417 (P1_U3689, P1_U5202, P1_U5203, P1_U5204);
  and ginst4418 (P1_U3690, P1_U5207, P1_U5208, P1_U5209);
  and ginst4419 (P1_U3691, P1_U5212, P1_U5213, P1_U5214);
  and ginst4420 (P1_U3692, P1_U5217, P1_U5218, P1_U5219);
  and ginst4421 (P1_U3693, P1_U5222, P1_U5223, P1_U5224);
  and ginst4422 (P1_U3694, P1_U5227, P1_U5228, P1_U5229);
  and ginst4423 (P1_U3695, P1_U4224, P1_U5242, P1_U5243);
  and ginst4424 (P1_U3696, P1_U5250, P1_U5251, P1_U5252);
  and ginst4425 (P1_U3697, P1_U5255, P1_U5256, P1_U5257);
  and ginst4426 (P1_U3698, P1_U5260, P1_U5261, P1_U5262);
  and ginst4427 (P1_U3699, P1_U5265, P1_U5266, P1_U5267);
  and ginst4428 (P1_U3700, P1_U5270, P1_U5271, P1_U5272);
  and ginst4429 (P1_U3701, P1_U5275, P1_U5276, P1_U5277);
  and ginst4430 (P1_U3702, P1_U5280, P1_U5281, P1_U5282);
  and ginst4431 (P1_U3703, P1_U5285, P1_U5286, P1_U5287);
  and ginst4432 (P1_U3704, P1_U4224, P1_U5299, P1_U5300);
  and ginst4433 (P1_U3705, P1_U5307, P1_U5308, P1_U5309);
  and ginst4434 (P1_U3706, P1_U5312, P1_U5313, P1_U5314);
  and ginst4435 (P1_U3707, P1_U5317, P1_U5318, P1_U5319);
  and ginst4436 (P1_U3708, P1_U5322, P1_U5323, P1_U5324);
  and ginst4437 (P1_U3709, P1_U5327, P1_U5328, P1_U5329);
  and ginst4438 (P1_U3710, P1_U5332, P1_U5333, P1_U5334);
  and ginst4439 (P1_U3711, P1_U5337, P1_U5338, P1_U5339);
  and ginst4440 (P1_U3712, P1_U5342, P1_U5343, P1_U5344);
  and ginst4441 (P1_U3713, P1_U4224, P1_U5357, P1_U5358);
  and ginst4442 (P1_U3714, P1_U5365, P1_U5366, P1_U5367);
  and ginst4443 (P1_U3715, P1_U5370, P1_U5371, P1_U5372);
  and ginst4444 (P1_U3716, P1_U5375, P1_U5376, P1_U5377);
  and ginst4445 (P1_U3717, P1_U5380, P1_U5381, P1_U5382);
  and ginst4446 (P1_U3718, P1_U5385, P1_U5386, P1_U5387);
  and ginst4447 (P1_U3719, P1_U5390, P1_U5391, P1_U5392);
  and ginst4448 (P1_U3720, P1_U5395, P1_U5396, P1_U5397);
  and ginst4449 (P1_U3721, P1_U5400, P1_U5401, P1_U5402);
  and ginst4450 (P1_U3722, P1_U4224, P1_U5414, P1_U5415);
  and ginst4451 (P1_U3723, P1_U5422, P1_U5423, P1_U5424);
  and ginst4452 (P1_U3724, P1_U5427, P1_U5428, P1_U5429);
  and ginst4453 (P1_U3725, P1_U5432, P1_U5433, P1_U5434);
  and ginst4454 (P1_U3726, P1_U5437, P1_U5438, P1_U5439);
  and ginst4455 (P1_U3727, P1_U5441, P1_U5442, P1_U5443);
  and ginst4456 (P1_U3728, P1_U5446, P1_U5447, P1_U5448);
  and ginst4457 (P1_U3729, P1_U5451, P1_U5452, P1_U5453);
  and ginst4458 (P1_U3730, P1_U5456, P1_U5457, P1_U5458);
  and ginst4459 (P1_U3731, P1_FLUSH_REG_SCAN_IN, P1_STATE2_REG_0__SCAN_IN);
  and ginst4460 (P1_U3732, P1_U4399, P1_U4494);
  and ginst4461 (P1_U3733, P1_U3257, P1_U4497);
  and ginst4462 (P1_U3734, P1_U3257, P1_U4210);
  and ginst4463 (P1_U3735, P1_U4217, P1_U7496);
  and ginst4464 (P1_U3736, P1_U5471, P1_U5472);
  and ginst4465 (P1_U3737, P1_U3736, P1_U5470);
  and ginst4466 (P1_U3738, P1_U2518, P1_U3737);
  and ginst4467 (P1_U3739, P1_U4242, P1_U5475);
  and ginst4468 (P1_U3740, P1_U5485, P1_U5486);
  and ginst4469 (P1_U3741, P1_U4400, P1_U4449);
  and ginst4470 (P1_U3742, P1_U3393, P1_U5496);
  and ginst4471 (P1_U3743, P1_U5497, P1_U5498);
  and ginst4472 (P1_U3744, P1_U3742, P1_U3743, P1_U5500, P1_U7627);
  and ginst4473 (P1_U3745, P1_U3397, P1_U4263);
  and ginst4474 (P1_U3746, P1_U2520, P1_U3279, P1_U3288, P1_U3411, P1_U3745);
  and ginst4475 (P1_U3747, P1_U3748, P1_U5502);
  and ginst4476 (P1_U3748, P1_U5504, P1_U5505);
  and ginst4477 (P1_U3749, P1_U5513, P1_U7716, P1_U7717);
  and ginst4478 (P1_U3750, P1_U5522, P1_U5524);
  and ginst4479 (P1_U3751, P1_U5543, P1_U5544);
  and ginst4480 (P1_U3752, P1_U5547, P1_U5548);
  and ginst4481 (P1_U3753, P1_U5552, P1_U5553);
  and ginst4482 (P1_U3754, P1_U3257, P1_U5558);
  and ginst4483 (P1_U3755, P1_U3284, P1_U3407);
  and ginst4484 (P1_U3756, P1_U5561, P1_U5563);
  and ginst4485 (P1_U3757, P1_U3398, P1_U3399, P1_U5567);
  and ginst4486 (P1_U3758, P1_U2520, P1_U3757, P1_U5568);
  and ginst4487 (P1_U3759, P1_U3284, P1_U4186);
  and ginst4488 (P1_U3760, P1_U3288, P1_U3448, P1_U4217);
  and ginst4489 (P1_U3761, P1_U5566, P1_U7507);
  and ginst4490 (P1_U3762, P1_STATE2_REG_2__SCAN_IN, P1_U7508);
  and ginst4491 (P1_U3763, P1_U5570, P1_U5571);
  and ginst4492 (P1_U3764, P1_U5572, P1_U5573);
  and ginst4493 (P1_U3765, P1_U5575, P1_U5576);
  and ginst4494 (P1_U3766, P1_U3765, P1_U5574);
  and ginst4495 (P1_U3767, P1_U5577, P1_U5578);
  and ginst4496 (P1_U3768, P1_U5579, P1_U5580);
  and ginst4497 (P1_U3769, P1_U5582, P1_U5583);
  and ginst4498 (P1_U3770, P1_U3769, P1_U5581);
  and ginst4499 (P1_U3771, P1_U5584, P1_U5585);
  and ginst4500 (P1_U3772, P1_U5586, P1_U5587);
  and ginst4501 (P1_U3773, P1_U5589, P1_U5590);
  and ginst4502 (P1_U3774, P1_U3773, P1_U5588);
  and ginst4503 (P1_U3775, P1_U5591, P1_U5592, P1_U5594);
  and ginst4504 (P1_U3776, P1_U3777, P1_U5593, P1_U5595);
  and ginst4505 (P1_U3777, P1_U5596, P1_U5597);
  and ginst4506 (P1_U3778, P1_U5598, P1_U5599, P1_U5601);
  and ginst4507 (P1_U3779, P1_U5603, P1_U5604);
  and ginst4508 (P1_U3780, P1_U3779, P1_U5602);
  and ginst4509 (P1_U3781, P1_U5605, P1_U5606, P1_U5608);
  and ginst4510 (P1_U3782, P1_U5610, P1_U5611);
  and ginst4511 (P1_U3783, P1_U3782, P1_U5609);
  and ginst4512 (P1_U3784, P1_U5612, P1_U5613, P1_U5615);
  and ginst4513 (P1_U3785, P1_U5617, P1_U5618);
  and ginst4514 (P1_U3786, P1_U3785, P1_U5616);
  and ginst4515 (P1_U3787, P1_U5619, P1_U5620, P1_U5622);
  and ginst4516 (P1_U3788, P1_U5624, P1_U5625);
  and ginst4517 (P1_U3789, P1_U3788, P1_U5623);
  and ginst4518 (P1_U3790, P1_U5626, P1_U5627, P1_U5629);
  and ginst4519 (P1_U3791, P1_U5631, P1_U5632);
  and ginst4520 (P1_U3792, P1_U3791, P1_U5630);
  and ginst4521 (P1_U3793, P1_U5633, P1_U5634, P1_U5636);
  and ginst4522 (P1_U3794, P1_U5638, P1_U5639);
  and ginst4523 (P1_U3795, P1_U3794, P1_U5637);
  and ginst4524 (P1_U3796, P1_U5640, P1_U5641, P1_U5643);
  and ginst4525 (P1_U3797, P1_U5645, P1_U5646);
  and ginst4526 (P1_U3798, P1_U3797, P1_U5644);
  and ginst4527 (P1_U3799, P1_U5647, P1_U5648, P1_U5650);
  and ginst4528 (P1_U3800, P1_U5652, P1_U5653);
  and ginst4529 (P1_U3801, P1_U3800, P1_U5651);
  and ginst4530 (P1_U3802, P1_U5654, P1_U5655, P1_U5657);
  and ginst4531 (P1_U3803, P1_U5659, P1_U5660);
  and ginst4532 (P1_U3804, P1_U3803, P1_U5658);
  and ginst4533 (P1_U3805, P1_U5662, P1_U5664);
  and ginst4534 (P1_U3806, P1_U5666, P1_U5667);
  and ginst4535 (P1_U3807, P1_U3806, P1_U5665);
  and ginst4536 (P1_U3808, P1_U5669, P1_U5671);
  and ginst4537 (P1_U3809, P1_U5673, P1_U5674);
  and ginst4538 (P1_U3810, P1_U3809, P1_U5672);
  and ginst4539 (P1_U3811, P1_U5676, P1_U5678);
  and ginst4540 (P1_U3812, P1_U5680, P1_U5681);
  and ginst4541 (P1_U3813, P1_U3812, P1_U5679);
  and ginst4542 (P1_U3814, P1_U5683, P1_U5685);
  and ginst4543 (P1_U3815, P1_U5687, P1_U5688);
  and ginst4544 (P1_U3816, P1_U3815, P1_U5686);
  and ginst4545 (P1_U3817, P1_U5690, P1_U5692);
  and ginst4546 (P1_U3818, P1_U5694, P1_U5695);
  and ginst4547 (P1_U3819, P1_U3818, P1_U5693);
  and ginst4548 (P1_U3820, P1_U5697, P1_U5699);
  and ginst4549 (P1_U3821, P1_U5701, P1_U5702);
  and ginst4550 (P1_U3822, P1_U3821, P1_U5700);
  and ginst4551 (P1_U3823, P1_U5704, P1_U5706);
  and ginst4552 (P1_U3824, P1_U5708, P1_U5709);
  and ginst4553 (P1_U3825, P1_U3824, P1_U5707);
  and ginst4554 (P1_U3826, P1_U5711, P1_U5713);
  and ginst4555 (P1_U3827, P1_U5715, P1_U5716);
  and ginst4556 (P1_U3828, P1_U3827, P1_U5714);
  and ginst4557 (P1_U3829, P1_U5718, P1_U5720);
  and ginst4558 (P1_U3830, P1_U5722, P1_U5723);
  and ginst4559 (P1_U3831, P1_U3830, P1_U5721);
  and ginst4560 (P1_U3832, P1_U5725, P1_U5727);
  and ginst4561 (P1_U3833, P1_U5729, P1_U5730);
  and ginst4562 (P1_U3834, P1_U3833, P1_U5728);
  and ginst4563 (P1_U3835, P1_U5732, P1_U5734);
  and ginst4564 (P1_U3836, P1_U5736, P1_U5737);
  and ginst4565 (P1_U3837, P1_U3836, P1_U5735);
  and ginst4566 (P1_U3838, P1_U5739, P1_U5741);
  and ginst4567 (P1_U3839, P1_U5743, P1_U5744);
  and ginst4568 (P1_U3840, P1_U3839, P1_U5742);
  and ginst4569 (P1_U3841, P1_U5746, P1_U5748);
  and ginst4570 (P1_U3842, P1_U5750, P1_U5751);
  and ginst4571 (P1_U3843, P1_U3842, P1_U5749);
  and ginst4572 (P1_U3844, P1_U5753, P1_U5755);
  and ginst4573 (P1_U3845, P1_U5757, P1_U5758);
  and ginst4574 (P1_U3846, P1_U3845, P1_U5756);
  and ginst4575 (P1_U3847, P1_U5760, P1_U5762);
  and ginst4576 (P1_U3848, P1_U5764, P1_U5765);
  and ginst4577 (P1_U3849, P1_U3848, P1_U5763);
  and ginst4578 (P1_U3850, P1_U5767, P1_U5769);
  and ginst4579 (P1_U3851, P1_U5771, P1_U5772);
  and ginst4580 (P1_U3852, P1_U3851, P1_U5770);
  and ginst4581 (P1_U3853, P1_U5774, P1_U5776);
  and ginst4582 (P1_U3854, P1_U5778, P1_U5779);
  and ginst4583 (P1_U3855, P1_U3854, P1_U5777);
  and ginst4584 (P1_U3856, P1_U5781, P1_U5783);
  and ginst4585 (P1_U3857, P1_U5785, P1_U5786);
  and ginst4586 (P1_U3858, P1_U3857, P1_U5784);
  and ginst4587 (P1_U3859, P1_U5788, P1_U5790);
  and ginst4588 (P1_U3860, P1_U5792, P1_U5793);
  and ginst4589 (P1_U3861, P1_U3860, P1_U5791);
  and ginst4590 (P1_U3862, P1_U3262, P1_U3283, P1_U7494);
  and ginst4591 (P1_U3863, P1_U3408, P1_U5794);
  and ginst4592 (P1_U3864, P1_STATEBS16_REG_SCAN_IN, P1_STATE2_REG_1__SCAN_IN);
  and ginst4593 (P1_U3865, P1_U2368, P1_U3284);
  and ginst4594 (P1_U3866, P1_STATE2_REG_0__SCAN_IN, P1_U2449);
  and ginst4595 (P1_U3867, P1_U2368, P1_U4208);
  and ginst4596 (P1_U3868, P1_U6105, P1_U6106);
  and ginst4597 (P1_U3869, P1_U6108, P1_U6109);
  and ginst4598 (P1_U3870, P1_U6111, P1_U6112);
  and ginst4599 (P1_U3871, P1_U6114, P1_U6115);
  and ginst4600 (P1_U3872, P1_U6117, P1_U6118);
  and ginst4601 (P1_U3873, P1_U6120, P1_U6121);
  and ginst4602 (P1_U3874, P1_U6123, P1_U6124);
  and ginst4603 (P1_U3875, P1_U6126, P1_U6127);
  and ginst4604 (P1_U3876, P1_U6129, P1_U6130);
  and ginst4605 (P1_U3877, P1_U6132, P1_U6133);
  and ginst4606 (P1_U3878, P1_U6135, P1_U6136);
  and ginst4607 (P1_U3879, P1_U6138, P1_U6139);
  and ginst4608 (P1_U3880, P1_U6141, P1_U6142);
  and ginst4609 (P1_U3881, P1_U6144, P1_U6145);
  and ginst4610 (P1_U3882, P1_U6147, P1_U6148);
  and ginst4611 (P1_U3883, P1_U6150, P1_U6151);
  and ginst4612 (P1_U3884, P1_U2605, P1_U3391);
  and ginst4613 (P1_U3885, P1_STATE2_REG_0__SCAN_IN, P1_U3271, P1_U7494);
  and ginst4614 (P1_U3886, P1_U4171, P1_U4399);
  and ginst4615 (P1_U3887, P1_U4241, P1_U4244, P1_U6362);
  nor ginst4616 (P1_U3888, P1_STATEBS16_REG_SCAN_IN, U210);
  and ginst4617 (P1_U3889, P1_U4186, P1_U4494);
  and ginst4618 (P1_U3890, P1_U6371, P1_U6372, P1_U6373, P1_U6374, P1_U6375);
  and ginst4619 (P1_U3891, P1_U6379, P1_U6380, P1_U6381, P1_U6382, P1_U6383);
  and ginst4620 (P1_U3892, P1_U6387, P1_U6388, P1_U6389, P1_U6390, P1_U6391);
  and ginst4621 (P1_U3893, P1_U6395, P1_U6396, P1_U6397, P1_U6398, P1_U6399);
  and ginst4622 (P1_U3894, P1_U4227, P1_U6400);
  and ginst4623 (P1_U3895, P1_U6404, P1_U6405, P1_U6406, P1_U6407);
  and ginst4624 (P1_U3896, P1_U4227, P1_U6408);
  and ginst4625 (P1_U3897, P1_U6411, P1_U6412, P1_U6413, P1_U6414, P1_U6415);
  and ginst4626 (P1_U3898, P1_U4227, P1_U6416);
  and ginst4627 (P1_U3899, P1_U6419, P1_U6421, P1_U6422);
  and ginst4628 (P1_U3900, P1_U4227, P1_U6423);
  and ginst4629 (P1_U3901, P1_U6426, P1_U6428, P1_U6429);
  and ginst4630 (P1_U3902, P1_U4227, P1_U6430);
  and ginst4631 (P1_U3903, P1_U6433, P1_U6435, P1_U6436);
  and ginst4632 (P1_U3904, P1_U4227, P1_U6437);
  and ginst4633 (P1_U3905, P1_U6440, P1_U6442, P1_U6443);
  and ginst4634 (P1_U3906, P1_U4227, P1_U6444);
  and ginst4635 (P1_U3907, P1_U6447, P1_U6449, P1_U6450);
  and ginst4636 (P1_U3908, P1_U4227, P1_U6451);
  and ginst4637 (P1_U3909, P1_U6454, P1_U6456, P1_U6457);
  and ginst4638 (P1_U3910, P1_U4227, P1_U6458);
  and ginst4639 (P1_U3911, P1_U6461, P1_U6463, P1_U6464);
  and ginst4640 (P1_U3912, P1_U4227, P1_U6465);
  and ginst4641 (P1_U3913, P1_U6468, P1_U6470, P1_U6471);
  and ginst4642 (P1_U3914, P1_U4227, P1_U6472);
  and ginst4643 (P1_U3915, P1_U6475, P1_U6477, P1_U6478);
  and ginst4644 (P1_U3916, P1_U4227, P1_U6479);
  and ginst4645 (P1_U3917, P1_U6482, P1_U6484, P1_U6485);
  and ginst4646 (P1_U3918, P1_U4227, P1_U6486);
  and ginst4647 (P1_U3919, P1_U6489, P1_U6491, P1_U6492);
  and ginst4648 (P1_U3920, P1_U4227, P1_U6494);
  and ginst4649 (P1_U3921, P1_U6496, P1_U6498, P1_U6499);
  and ginst4650 (P1_U3922, P1_U4227, P1_U6501);
  and ginst4651 (P1_U3923, P1_U6503, P1_U6505, P1_U6506);
  and ginst4652 (P1_U3924, P1_U4227, P1_U6508);
  and ginst4653 (P1_U3925, P1_U6510, P1_U6512, P1_U6513);
  and ginst4654 (P1_U3926, P1_U6515, P1_U6517);
  and ginst4655 (P1_U3927, P1_U6519, P1_U6520);
  and ginst4656 (P1_U3928, P1_U6522, P1_U6524);
  and ginst4657 (P1_U3929, P1_U6526, P1_U6527);
  and ginst4658 (P1_U3930, P1_U6529, P1_U6531);
  and ginst4659 (P1_U3931, P1_U6533, P1_U6534);
  and ginst4660 (P1_U3932, P1_U6536, P1_U6538);
  and ginst4661 (P1_U3933, P1_U6540, P1_U6541);
  and ginst4662 (P1_U3934, P1_U6543, P1_U6545);
  and ginst4663 (P1_U3935, P1_U6547, P1_U6548);
  and ginst4664 (P1_U3936, P1_U6550, P1_U6552);
  and ginst4665 (P1_U3937, P1_U6554, P1_U6555);
  and ginst4666 (P1_U3938, P1_U6557, P1_U6559);
  and ginst4667 (P1_U3939, P1_U6561, P1_U6562);
  and ginst4668 (P1_U3940, P1_U6564, P1_U6566);
  and ginst4669 (P1_U3941, P1_U6568, P1_U6569);
  and ginst4670 (P1_U3942, P1_U6571, P1_U6573);
  and ginst4671 (P1_U3943, P1_U6575, P1_U6576);
  and ginst4672 (P1_U3944, P1_U6578, P1_U6580);
  and ginst4673 (P1_U3945, P1_U6582, P1_U6583);
  and ginst4674 (P1_U3946, P1_U6585, P1_U6587);
  and ginst4675 (P1_U3947, P1_U6589, P1_U6590);
  and ginst4676 (P1_U3948, P1_U6592, P1_U6594);
  and ginst4677 (P1_U3949, P1_U6596, P1_U6597);
  nor ginst4678 (P1_U3950, P1_DATAWIDTH_REG_2__SCAN_IN, P1_DATAWIDTH_REG_3__SCAN_IN, P1_DATAWIDTH_REG_4__SCAN_IN, P1_DATAWIDTH_REG_5__SCAN_IN);
  nor ginst4679 (P1_U3951, P1_DATAWIDTH_REG_6__SCAN_IN, P1_DATAWIDTH_REG_7__SCAN_IN, P1_DATAWIDTH_REG_8__SCAN_IN, P1_DATAWIDTH_REG_9__SCAN_IN);
  and ginst4680 (P1_U3952, P1_U3950, P1_U3951);
  nor ginst4681 (P1_U3953, P1_DATAWIDTH_REG_10__SCAN_IN, P1_DATAWIDTH_REG_11__SCAN_IN, P1_DATAWIDTH_REG_12__SCAN_IN, P1_DATAWIDTH_REG_13__SCAN_IN);
  nor ginst4682 (P1_U3954, P1_DATAWIDTH_REG_14__SCAN_IN, P1_DATAWIDTH_REG_15__SCAN_IN, P1_DATAWIDTH_REG_16__SCAN_IN, P1_DATAWIDTH_REG_17__SCAN_IN);
  and ginst4683 (P1_U3955, P1_U3953, P1_U3954);
  nor ginst4684 (P1_U3956, P1_DATAWIDTH_REG_18__SCAN_IN, P1_DATAWIDTH_REG_19__SCAN_IN, P1_DATAWIDTH_REG_20__SCAN_IN, P1_DATAWIDTH_REG_21__SCAN_IN);
  nor ginst4685 (P1_U3957, P1_DATAWIDTH_REG_22__SCAN_IN, P1_DATAWIDTH_REG_23__SCAN_IN, P1_DATAWIDTH_REG_24__SCAN_IN, P1_DATAWIDTH_REG_25__SCAN_IN);
  and ginst4686 (P1_U3958, P1_U3956, P1_U3957);
  nor ginst4687 (P1_U3959, P1_DATAWIDTH_REG_26__SCAN_IN, P1_DATAWIDTH_REG_27__SCAN_IN);
  nor ginst4688 (P1_U3960, P1_DATAWIDTH_REG_28__SCAN_IN, P1_DATAWIDTH_REG_29__SCAN_IN);
  nor ginst4689 (P1_U3961, P1_DATAWIDTH_REG_30__SCAN_IN, P1_DATAWIDTH_REG_31__SCAN_IN);
  and ginst4690 (P1_U3962, P1_U3959, P1_U3960, P1_U3961, P1_U6598);
  nor ginst4691 (P1_U3963, P1_REIP_REG_0__SCAN_IN, P1_DATAWIDTH_REG_0__SCAN_IN, P1_DATAWIDTH_REG_1__SCAN_IN);
  and ginst4692 (P1_U3964, P1_STATE2_REG_2__SCAN_IN, P1_U3257);
  and ginst4693 (P1_U3965, P1_U3298, P1_U6608);
  nor ginst4694 (P1_U3966, P1_STATE2_REG_0__SCAN_IN, U210);
  and ginst4695 (P1_U3967, P1_U3307, P1_U3408, P1_U6602);
  and ginst4696 (P1_U3968, P1_STATE2_REG_2__SCAN_IN, P1_U3287);
  and ginst4697 (P1_U3969, P1_U4206, P1_U4235);
  and ginst4698 (P1_U3970, P1_U6618, P1_U6619, P1_U6620, P1_U6621);
  and ginst4699 (P1_U3971, P1_U6622, P1_U6623, P1_U6624, P1_U6625);
  and ginst4700 (P1_U3972, P1_U6626, P1_U6627, P1_U6628, P1_U6629);
  and ginst4701 (P1_U3973, P1_U6630, P1_U6631, P1_U6632, P1_U6633);
  and ginst4702 (P1_U3974, P1_U6634, P1_U6635, P1_U6636, P1_U6637);
  and ginst4703 (P1_U3975, P1_U6638, P1_U6639, P1_U6640, P1_U6641);
  and ginst4704 (P1_U3976, P1_U6642, P1_U6643, P1_U6644, P1_U6645);
  and ginst4705 (P1_U3977, P1_U6646, P1_U6647, P1_U6648, P1_U6649);
  and ginst4706 (P1_U3978, P1_U6650, P1_U6651, P1_U6652, P1_U6653);
  and ginst4707 (P1_U3979, P1_U6654, P1_U6655, P1_U6656, P1_U6657);
  and ginst4708 (P1_U3980, P1_U6658, P1_U6659, P1_U6660, P1_U6661);
  and ginst4709 (P1_U3981, P1_U6662, P1_U6663, P1_U6664, P1_U6665);
  and ginst4710 (P1_U3982, P1_U6666, P1_U6667, P1_U6668, P1_U6669);
  and ginst4711 (P1_U3983, P1_U6670, P1_U6671, P1_U6672, P1_U6673);
  and ginst4712 (P1_U3984, P1_U6674, P1_U6675, P1_U6676, P1_U6677);
  and ginst4713 (P1_U3985, P1_U6678, P1_U6679, P1_U6680, P1_U7613);
  and ginst4714 (P1_U3986, P1_U6681, P1_U6682, P1_U6683, P1_U6684);
  and ginst4715 (P1_U3987, P1_U6685, P1_U6686, P1_U6687, P1_U6688);
  and ginst4716 (P1_U3988, P1_U6689, P1_U6690, P1_U6691, P1_U6692);
  and ginst4717 (P1_U3989, P1_U6693, P1_U6694, P1_U6695, P1_U6696);
  and ginst4718 (P1_U3990, P1_U6697, P1_U6698, P1_U6699, P1_U6700);
  and ginst4719 (P1_U3991, P1_U6701, P1_U6702, P1_U6703, P1_U6704);
  and ginst4720 (P1_U3992, P1_U6705, P1_U6706, P1_U6707, P1_U6708);
  and ginst4721 (P1_U3993, P1_U6709, P1_U6710, P1_U6711, P1_U6712);
  and ginst4722 (P1_U3994, P1_U6713, P1_U6714, P1_U6715, P1_U6716);
  and ginst4723 (P1_U3995, P1_U6717, P1_U6718, P1_U6719, P1_U6720);
  and ginst4724 (P1_U3996, P1_U6721, P1_U6722, P1_U6723, P1_U6724);
  and ginst4725 (P1_U3997, P1_U6725, P1_U6726, P1_U6727, P1_U6728);
  and ginst4726 (P1_U3998, P1_U6729, P1_U6730, P1_U6731, P1_U6732);
  and ginst4727 (P1_U3999, P1_U6733, P1_U6734, P1_U6735, P1_U6736);
  and ginst4728 (P1_U4000, P1_U6737, P1_U6738, P1_U6739, P1_U6740);
  and ginst4729 (P1_U4001, P1_U6741, P1_U6742, P1_U6743, P1_U6744);
  and ginst4730 (P1_U4002, P1_U6748, P1_U6749);
  and ginst4731 (P1_U4003, P1_U6751, P1_U6752);
  and ginst4732 (P1_U4004, P1_U6754, P1_U6755);
  and ginst4733 (P1_U4005, P1_U6757, P1_U6758);
  and ginst4734 (P1_U4006, P1_U4007, P1_U6760);
  and ginst4735 (P1_U4007, P1_U6761, P1_U6762);
  and ginst4736 (P1_U4008, P1_U6764, P1_U6765);
  and ginst4737 (P1_U4009, P1_U6772, P1_U6773, P1_U6774);
  and ginst4738 (P1_U4010, P1_U6776, P1_U6777);
  and ginst4739 (P1_U4011, P1_U6781, P1_U6782, P1_U6783);
  and ginst4740 (P1_U4012, P1_U6785, P1_U6786, P1_U6787);
  and ginst4741 (P1_U4013, P1_U6789, P1_U6790, P1_U6791);
  and ginst4742 (P1_U4014, P1_U6793, P1_U6794, P1_U6795);
  and ginst4743 (P1_U4015, P1_U6797, P1_U6798, P1_U6799);
  and ginst4744 (P1_U4016, P1_U6801, P1_U6802, P1_U6803);
  and ginst4745 (P1_U4017, P1_U6805, P1_U6806, P1_U6807);
  and ginst4746 (P1_U4018, P1_U6809, P1_U6810, P1_U6811);
  and ginst4747 (P1_U4019, P1_U6813, P1_U6814, P1_U6815);
  and ginst4748 (P1_U4020, P1_U6817, P1_U6818, P1_U6819);
  and ginst4749 (P1_U4021, P1_U6821, P1_U6822);
  and ginst4750 (P1_U4022, P1_U6826, P1_U6827, P1_U6828);
  and ginst4751 (P1_U4023, P1_U6830, P1_U6831, P1_U6832);
  and ginst4752 (P1_U4024, P1_U6834, P1_U6835, P1_U6836);
  and ginst4753 (P1_U4025, P1_U6838, P1_U6839, P1_U6840);
  and ginst4754 (P1_U4026, P1_U6857, P1_U6858);
  and ginst4755 (P1_U4027, P1_U6860, P1_U6861);
  and ginst4756 (P1_U4028, P1_U3283, P1_U6888, P1_U7494);
  and ginst4757 (P1_U4029, P1_U6892, P1_U6893, P1_U6894, P1_U6895);
  and ginst4758 (P1_U4030, P1_U6896, P1_U6897, P1_U6898, P1_U6899);
  and ginst4759 (P1_U4031, P1_U6900, P1_U6901, P1_U6902, P1_U6903);
  and ginst4760 (P1_U4032, P1_U6904, P1_U6905, P1_U6906, P1_U6907);
  and ginst4761 (P1_U4033, P1_U6910, P1_U6911, P1_U6912, P1_U6913);
  and ginst4762 (P1_U4034, P1_U6914, P1_U6915, P1_U6916, P1_U6917);
  and ginst4763 (P1_U4035, P1_U6918, P1_U6919, P1_U6920, P1_U6921);
  and ginst4764 (P1_U4036, P1_U6922, P1_U6923, P1_U6924, P1_U6925);
  and ginst4765 (P1_U4037, P1_U6941, P1_U6942, P1_U6943, P1_U6944);
  and ginst4766 (P1_U4038, P1_U6945, P1_U6946, P1_U6947, P1_U6948);
  and ginst4767 (P1_U4039, P1_U6949, P1_U6950, P1_U6951, P1_U6952);
  and ginst4768 (P1_U4040, P1_U6953, P1_U6954, P1_U6955, P1_U6956);
  and ginst4769 (P1_U4041, P1_U6958, P1_U6959, P1_U6960, P1_U6961);
  and ginst4770 (P1_U4042, P1_U6962, P1_U6963, P1_U6964, P1_U6965);
  and ginst4771 (P1_U4043, P1_U6966, P1_U6967, P1_U6968, P1_U6969);
  and ginst4772 (P1_U4044, P1_U6970, P1_U6971, P1_U6972, P1_U6973);
  and ginst4773 (P1_U4045, P1_U6975, P1_U6976, P1_U6977, P1_U6978);
  and ginst4774 (P1_U4046, P1_U6979, P1_U6980, P1_U6981, P1_U6982);
  and ginst4775 (P1_U4047, P1_U6983, P1_U6984, P1_U6985, P1_U6986);
  and ginst4776 (P1_U4048, P1_U6987, P1_U6988, P1_U6989, P1_U6990);
  and ginst4777 (P1_U4049, P1_U6992, P1_U6993, P1_U6994, P1_U6995);
  and ginst4778 (P1_U4050, P1_U6996, P1_U6997, P1_U6998, P1_U6999);
  and ginst4779 (P1_U4051, P1_U7000, P1_U7001, P1_U7002, P1_U7003);
  and ginst4780 (P1_U4052, P1_U7004, P1_U7005, P1_U7006, P1_U7614);
  and ginst4781 (P1_U4053, P1_U7007, P1_U7008, P1_U7009, P1_U7010);
  and ginst4782 (P1_U4054, P1_U7011, P1_U7012, P1_U7013, P1_U7014);
  and ginst4783 (P1_U4055, P1_U7015, P1_U7016, P1_U7017, P1_U7018);
  and ginst4784 (P1_U4056, P1_U7019, P1_U7020, P1_U7021, P1_U7022);
  and ginst4785 (P1_U4057, P1_U7024, P1_U7025, P1_U7026, P1_U7027);
  and ginst4786 (P1_U4058, P1_U7028, P1_U7029, P1_U7030, P1_U7031);
  and ginst4787 (P1_U4059, P1_U7032, P1_U7033, P1_U7034, P1_U7035);
  and ginst4788 (P1_U4060, P1_U7036, P1_U7037, P1_U7038, P1_U7039);
  and ginst4789 (P1_U4061, P1_U3443, P1_U7059);
  and ginst4790 (P1_U4062, P1_STATE2_REG_0__SCAN_IN, P1_U7062);
  and ginst4791 (P1_U4063, P1_U7066, P1_U7067, P1_U7068, P1_U7069);
  and ginst4792 (P1_U4064, P1_U7070, P1_U7071, P1_U7072, P1_U7073);
  and ginst4793 (P1_U4065, P1_U7074, P1_U7075, P1_U7076, P1_U7077);
  and ginst4794 (P1_U4066, P1_U7078, P1_U7079, P1_U7080, P1_U7081);
  and ginst4795 (P1_U4067, P1_STATE2_REG_0__SCAN_IN, P1_U4256);
  and ginst4796 (P1_U4068, P1_U4401, P1_U4403, P1_U4404, P1_U4405);
  and ginst4797 (P1_U4069, P1_U4406, P1_U4407, P1_U4408);
  and ginst4798 (P1_U4070, P1_U4409, P1_U4410, P1_U4411, P1_U4412);
  and ginst4799 (P1_U4071, P1_U4413, P1_U4414);
  and ginst4800 (P1_U4072, P1_U3391, P1_U4400);
  and ginst4801 (P1_U4073, P1_STATE2_REG_0__SCAN_IN, P1_U3284);
  and ginst4802 (P1_U4074, P1_U7089, P1_U7090);
  and ginst4803 (P1_U4075, P1_U3434, P1_U7472, P1_U7473);
  and ginst4804 (P1_U4076, P1_U7474, P1_U7475, P1_U7476);
  and ginst4805 (P1_U4077, P1_U2606, P1_U4076, P1_U7477);
  and ginst4806 (P1_U4078, P1_U7095, P1_U7097);
  and ginst4807 (P1_U4079, P1_U7098, P1_U7099, P1_U7100, P1_U7101);
  and ginst4808 (P1_U4080, P1_U7102, P1_U7103, P1_U7104, P1_U7105);
  and ginst4809 (P1_U4081, P1_U7106, P1_U7107, P1_U7108, P1_U7109);
  and ginst4810 (P1_U4082, P1_U7110, P1_U7111, P1_U7112, P1_U7113);
  and ginst4811 (P1_U4083, P1_U7115, P1_U7116, P1_U7117, P1_U7118);
  and ginst4812 (P1_U4084, P1_U7119, P1_U7120, P1_U7121, P1_U7122);
  and ginst4813 (P1_U4085, P1_U7123, P1_U7124, P1_U7125, P1_U7126);
  and ginst4814 (P1_U4086, P1_U7127, P1_U7128, P1_U7129, P1_U7130);
  and ginst4815 (P1_U4087, P1_U7132, P1_U7133, P1_U7134, P1_U7135);
  and ginst4816 (P1_U4088, P1_U7136, P1_U7137, P1_U7138, P1_U7139);
  and ginst4817 (P1_U4089, P1_U7140, P1_U7141, P1_U7142, P1_U7143);
  and ginst4818 (P1_U4090, P1_U7144, P1_U7145);
  and ginst4819 (P1_U4091, P1_U4090, P1_U7146, P1_U7617);
  and ginst4820 (P1_U4092, P1_U7147, P1_U7148, P1_U7149, P1_U7150);
  and ginst4821 (P1_U4093, P1_U7151, P1_U7152, P1_U7153, P1_U7154);
  and ginst4822 (P1_U4094, P1_U7155, P1_U7156, P1_U7157, P1_U7158);
  and ginst4823 (P1_U4095, P1_U7159, P1_U7160, P1_U7161, P1_U7162);
  and ginst4824 (P1_U4096, P1_U7164, P1_U7165, P1_U7166, P1_U7167);
  and ginst4825 (P1_U4097, P1_U7168, P1_U7169, P1_U7170, P1_U7171);
  and ginst4826 (P1_U4098, P1_U7172, P1_U7173, P1_U7174, P1_U7175);
  and ginst4827 (P1_U4099, P1_U7176, P1_U7177, P1_U7178, P1_U7179);
  and ginst4828 (P1_U4100, P1_U7181, P1_U7182, P1_U7183, P1_U7184);
  and ginst4829 (P1_U4101, P1_U7185, P1_U7186, P1_U7187, P1_U7188);
  and ginst4830 (P1_U4102, P1_U7189, P1_U7190, P1_U7191, P1_U7192);
  and ginst4831 (P1_U4103, P1_U7193, P1_U7194, P1_U7195, P1_U7196);
  and ginst4832 (P1_U4104, P1_U7198, P1_U7199, P1_U7200, P1_U7201);
  and ginst4833 (P1_U4105, P1_U7202, P1_U7203, P1_U7204, P1_U7205);
  and ginst4834 (P1_U4106, P1_U7206, P1_U7207, P1_U7208, P1_U7209);
  and ginst4835 (P1_U4107, P1_U7210, P1_U7211, P1_U7212, P1_U7213);
  and ginst4836 (P1_U4108, P1_U3264, P1_U7215);
  and ginst4837 (P1_U4109, P1_U7215, P1_U7216);
  and ginst4838 (P1_U4110, P1_U3265, P1_U7217);
  and ginst4839 (P1_U4111, P1_U3427, P1_U7089);
  and ginst4840 (P1_U4112, P1_U7217, P1_U7218);
  and ginst4841 (P1_U4113, P1_U4112, P1_U7472, P1_U7473);
  and ginst4842 (P1_U4114, P1_U3434, P1_U4111, P1_U4113, P1_U7090);
  and ginst4843 (P1_U4115, P1_U7474, P1_U7476, P1_U7480, P1_U7486);
  and ginst4844 (P1_U4116, P1_U7487, P1_U7488, P1_U7489, P1_U7505);
  and ginst4845 (P1_U4117, P1_U7089, P1_U7090);
  and ginst4846 (P1_U4118, P1_U3434, P1_U7472, P1_U7473);
  and ginst4847 (P1_U4119, P1_U7474, P1_U7475, P1_U7476);
  and ginst4848 (P1_U4120, P1_U2606, P1_U2608, P1_U4119, P1_U7477);
  and ginst4849 (P1_U4121, P1_U7220, P1_U7221, P1_U7222, P1_U7223);
  and ginst4850 (P1_U4122, P1_U7224, P1_U7225, P1_U7226, P1_U7227);
  and ginst4851 (P1_U4123, P1_U7228, P1_U7229, P1_U7230, P1_U7231);
  and ginst4852 (P1_U4124, P1_U7232, P1_U7233, P1_U7234, P1_U7235);
  and ginst4853 (P1_U4125, P1_U7237, P1_U7238, P1_U7239, P1_U7240);
  and ginst4854 (P1_U4126, P1_U7241, P1_U7242, P1_U7243, P1_U7244);
  and ginst4855 (P1_U4127, P1_U7245, P1_U7246, P1_U7247, P1_U7248);
  and ginst4856 (P1_U4128, P1_U7249, P1_U7250, P1_U7251, P1_U7252);
  and ginst4857 (P1_U4129, P1_U7254, P1_U7255, P1_U7256, P1_U7257);
  and ginst4858 (P1_U4130, P1_U7258, P1_U7259, P1_U7260, P1_U7261);
  and ginst4859 (P1_U4131, P1_U7262, P1_U7263, P1_U7264, P1_U7265);
  and ginst4860 (P1_U4132, P1_U7266, P1_U7267, P1_U7268, P1_U7269);
  and ginst4861 (P1_U4133, P1_U7271, P1_U7272, P1_U7273, P1_U7274);
  and ginst4862 (P1_U4134, P1_U7275, P1_U7276, P1_U7277, P1_U7278);
  and ginst4863 (P1_U4135, P1_U7279, P1_U7280, P1_U7281, P1_U7282);
  and ginst4864 (P1_U4136, P1_U7283, P1_U7284, P1_U7285, P1_U7619);
  and ginst4865 (P1_U4137, P1_U7286, P1_U7287, P1_U7288, P1_U7289);
  and ginst4866 (P1_U4138, P1_U7290, P1_U7291, P1_U7292, P1_U7293);
  and ginst4867 (P1_U4139, P1_U7294, P1_U7295, P1_U7296, P1_U7297);
  and ginst4868 (P1_U4140, P1_U7298, P1_U7299, P1_U7300, P1_U7301);
  and ginst4869 (P1_U4141, P1_U7303, P1_U7304, P1_U7305, P1_U7306);
  and ginst4870 (P1_U4142, P1_U7307, P1_U7308, P1_U7309, P1_U7310);
  and ginst4871 (P1_U4143, P1_U7311, P1_U7312, P1_U7313, P1_U7314);
  and ginst4872 (P1_U4144, P1_U7315, P1_U7316, P1_U7317, P1_U7318);
  and ginst4873 (P1_U4145, P1_U7320, P1_U7321, P1_U7322, P1_U7323);
  and ginst4874 (P1_U4146, P1_U7324, P1_U7325, P1_U7326, P1_U7327);
  and ginst4875 (P1_U4147, P1_U7328, P1_U7329, P1_U7330, P1_U7331);
  and ginst4876 (P1_U4148, P1_U7332, P1_U7333, P1_U7334, P1_U7335);
  and ginst4877 (P1_U4149, P1_U7337, P1_U7338, P1_U7339, P1_U7340);
  and ginst4878 (P1_U4150, P1_U7341, P1_U7342, P1_U7343, P1_U7344);
  and ginst4879 (P1_U4151, P1_U7345, P1_U7346, P1_U7347, P1_U7348);
  and ginst4880 (P1_U4152, P1_U7349, P1_U7350, P1_U7351, P1_U7352);
  and ginst4881 (P1_U4153, P1_U3284, P1_U3419);
  and ginst4882 (P1_U4154, P1_U3283, P1_U3391);
  and ginst4883 (P1_U4155, P1_U4263, P1_U7357, P1_U7358);
  and ginst4884 (P1_U4156, P1_U4155, P1_U7359);
  and ginst4885 (P1_U4157, P1_STATE2_REG_0__SCAN_IN, P1_U2427);
  and ginst4886 (P1_U4158, P1_U4157, P1_U7360);
  and ginst4887 (P1_U4159, P1_U3271, P1_U4173);
  and ginst4888 (P1_U4160, P1_STATE2_REG_0__SCAN_IN, P1_U4173);
  and ginst4889 (P1_U4161, P1_STATE2_REG_0__SCAN_IN, P1_U7369);
  and ginst4890 (P1_U4162, P1_U2603, P1_U7371);
  and ginst4891 (P1_U4163, P1_STATE2_REG_0__SCAN_IN, P1_U7373);
  and ginst4892 (P1_U4164, P1_U2603, P1_U7375);
  and ginst4893 (P1_U4165, P1_U7382, P1_U7383);
  and ginst4894 (P1_U4166, P1_U3453, P1_U7384);
  and ginst4895 (P1_U4167, P1_U7387, P1_U7388, P1_U7389);
  and ginst4896 (P1_U4168, P1_U7461, P1_U7462);
  and ginst4897 (P1_U4169, P1_U7464, P1_U7465);
  and ginst4898 (P1_U4170, P1_U7673, P1_U7674);
  nand ginst4899 (P1_U4171, P1_U3569, P1_U3570, P1_U3571, P1_U3572);
  nand ginst4900 (P1_U4172, P1_U3739, P1_U5474);
  nand ginst4901 (P1_U4173, P1_U2607, P1_U3573, P1_U3574, P1_U3575, P1_U3576);
  not ginst4902 (P1_U4174, P1_INSTADDRPOINTER_REG_31__SCAN_IN);
  and ginst4903 (P1_U4175, P1_U7725, P1_U7726);
  and ginst4904 (P1_U4176, P1_U7744, P1_U7745);
  nand ginst4905 (P1_U4177, P1_U2368, P1_U3285);
  nand ginst4906 (P1_U4178, P1_U3391, P1_U4508);
  not ginst4907 (P1_U4179, BS16);
  nand ginst4908 (P1_U4180, P1_U3967, P1_U4228);
  nand ginst4909 (P1_U4181, P1_U3432, P1_U4228);
  nand ginst4910 (P1_U4182, P1_U3738, P1_U7697, P1_U7698);
  nand ginst4911 (P1_U4183, P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN, P1_U3269);
  not ginst4912 (P1_U4184, P1_U3452);
  nand ginst4913 (P1_U4185, HOLD, P1_U3257);
  not ginst4914 (P1_U4186, P1_U3412);
  not ginst4915 (P1_U4187, P1_U3440);
  not ginst4916 (P1_U4188, P1_U3439);
  not ginst4917 (P1_U4189, P1_U3393);
  not ginst4918 (P1_U4190, P1_U3290);
  not ginst4919 (P1_U4191, P1_U3449);
  not ginst4920 (P1_U4192, P1_U3405);
  not ginst4921 (P1_U4193, P1_U3434);
  not ginst4922 (P1_U4194, P1_U3420);
  nand ginst4923 (P1_U4195, P1_U3271, P1_U4265);
  nand ginst4924 (P1_U4196, P1_U2605, P1_U4460);
  not ginst4925 (P1_U4197, P1_U3396);
  not ginst4926 (P1_U4198, P1_U3425);
  not ginst4927 (P1_U4199, P1_U3289);
  not ginst4928 (P1_U4200, P1_U3421);
  not ginst4929 (P1_U4201, P1_U3422);
  not ginst4930 (P1_U4202, P1_U3428);
  not ginst4931 (P1_U4203, P1_U3408);
  not ginst4932 (P1_U4204, P1_U3427);
  nand ginst4933 (P1_U4205, P1_U3885, P1_U4189, P1_U4197);
  not ginst4934 (P1_U4206, P1_U3418);
  not ginst4935 (P1_U4207, P1_U3443);
  not ginst4936 (P1_U4208, P1_U3282);
  not ginst4937 (P1_U4209, P1_U3307);
  not ginst4938 (P1_U4210, P1_U3390);
  not ginst4939 (P1_U4211, P1_U3446);
  not ginst4940 (P1_U4212, P1_U3447);
  not ginst4941 (P1_U4213, P1_U3448);
  not ginst4942 (P1_U4214, P1_U3400);
  not ginst4943 (P1_U4215, P1_U3288);
  not ginst4944 (P1_U4216, P1_U3292);
  nand ginst4945 (P1_U4217, P1_U2431, P1_U3578);
  not ginst4946 (P1_U4218, P1_U3399);
  nand ginst4947 (P1_U4219, P1_U3271, P1_U4449);
  not ginst4948 (P1_U4220, P1_U3433);
  not ginst4949 (P1_U4221, P1_U3249);
  not ginst4950 (P1_U4222, P1_U3426);
  not ginst4951 (P1_U4223, P1_U3424);
  not ginst4952 (P1_U4224, P1_U3300);
  not ginst4953 (P1_U4225, P1_LT_563_1260_U6);
  not ginst4954 (P1_U4226, P1_U3320);
  nand ginst4955 (P1_U4227, P1_U3431, P1_U4255);
  nand ginst4956 (P1_U4228, P1_U4235, P1_U7500);
  nand ginst4957 (P1_U4229, P1_U2362, P1_U3272);
  nand ginst4958 (P1_U4230, P1_U2363, P1_U4377);
  not ginst4959 (P1_U4231, P1_U3407);
  not ginst4960 (P1_U4232, P1_U3252);
  not ginst4961 (P1_U4233, P1_U3250);
  not ginst4962 (P1_U4234, P1_U3395);
  not ginst4963 (P1_U4235, P1_U3297);
  not ginst4964 (P1_U4236, P1_U3398);
  not ginst4965 (P1_U4237, P1_U4178);
  not ginst4966 (P1_U4238, P1_U3357);
  nand ginst4967 (P1_U4239, P1_U4477, P1_U7381);
  nand ginst4968 (P1_U4240, P1_U3963, P1_U4220);
  nand ginst4969 (P1_U4241, P1_U3584, P1_U4261);
  nand ginst4970 (P1_U4242, P1_U2428, P1_U3731);
  nand ginst4971 (P1_U4243, P1_U3258, P1_U4364);
  nand ginst4972 (P1_U4244, P1_STATE2_REG_1__SCAN_IN, P1_U2352, P1_U3294);
  nand ginst4973 (P1_U4245, P1_U2428, P1_U3403);
  nand ginst4974 (P1_U4246, P1_STATE2_REG_0__SCAN_IN, P1_U3263, U210);
  not ginst4975 (P1_U4247, P1_U3394);
  nand ginst4976 (P1_U4248, P1_U2353, P1_U2448, P1_U2451, P1_U3862);
  not ginst4977 (P1_U4249, P1_U3287);
  not ginst4978 (P1_U4250, P1_U3397);
  not ginst4979 (P1_U4251, P1_U3415);
  not ginst4980 (P1_U4252, P1_U3299);
  not ginst4981 (P1_U4253, P1_U3409);
  not ginst4982 (P1_U4254, P1_U3419);
  not ginst4983 (P1_U4255, P1_U3432);
  not ginst4984 (P1_U4256, P1_U3291);
  not ginst4985 (P1_U4257, P1_U3389);
  not ginst4986 (P1_U4258, P1_U3254);
  not ginst4987 (P1_U4259, P1_U3281);
  not ginst4988 (P1_U4260, P1_U3406);
  not ginst4989 (P1_U4261, P1_U3298);
  not ginst4990 (P1_U4262, P1_U3286);
  nand ginst4991 (P1_U4263, P1_U4236, P1_U4399);
  not ginst4992 (P1_U4264, P1_U3411);
  not ginst4993 (P1_U4265, P1_U3453);
  not ginst4994 (P1_U4266, P1_U3410);
  nand ginst4995 (P1_U4267, P1_REIP_REG_31__SCAN_IN, P1_U4233);
  nand ginst4996 (P1_U4268, P1_REIP_REG_30__SCAN_IN, P1_U4232);
  nand ginst4997 (P1_U4269, P1_ADDRESS_REG_29__SCAN_IN, P1_U3249);
  nand ginst4998 (P1_U4270, P1_REIP_REG_30__SCAN_IN, P1_U4233);
  nand ginst4999 (P1_U4271, P1_REIP_REG_29__SCAN_IN, P1_U4232);
  nand ginst5000 (P1_U4272, P1_ADDRESS_REG_28__SCAN_IN, P1_U3249);
  nand ginst5001 (P1_U4273, P1_REIP_REG_29__SCAN_IN, P1_U4233);
  nand ginst5002 (P1_U4274, P1_REIP_REG_28__SCAN_IN, P1_U4232);
  nand ginst5003 (P1_U4275, P1_ADDRESS_REG_27__SCAN_IN, P1_U3249);
  nand ginst5004 (P1_U4276, P1_REIP_REG_28__SCAN_IN, P1_U4233);
  nand ginst5005 (P1_U4277, P1_REIP_REG_27__SCAN_IN, P1_U4232);
  nand ginst5006 (P1_U4278, P1_ADDRESS_REG_26__SCAN_IN, P1_U3249);
  nand ginst5007 (P1_U4279, P1_REIP_REG_27__SCAN_IN, P1_U4233);
  nand ginst5008 (P1_U4280, P1_REIP_REG_26__SCAN_IN, P1_U4232);
  nand ginst5009 (P1_U4281, P1_ADDRESS_REG_25__SCAN_IN, P1_U3249);
  nand ginst5010 (P1_U4282, P1_REIP_REG_26__SCAN_IN, P1_U4233);
  nand ginst5011 (P1_U4283, P1_REIP_REG_25__SCAN_IN, P1_U4232);
  nand ginst5012 (P1_U4284, P1_ADDRESS_REG_24__SCAN_IN, P1_U3249);
  nand ginst5013 (P1_U4285, P1_REIP_REG_25__SCAN_IN, P1_U4233);
  nand ginst5014 (P1_U4286, P1_REIP_REG_24__SCAN_IN, P1_U4232);
  nand ginst5015 (P1_U4287, P1_ADDRESS_REG_23__SCAN_IN, P1_U3249);
  nand ginst5016 (P1_U4288, P1_REIP_REG_24__SCAN_IN, P1_U4233);
  nand ginst5017 (P1_U4289, P1_REIP_REG_23__SCAN_IN, P1_U4232);
  nand ginst5018 (P1_U4290, P1_ADDRESS_REG_22__SCAN_IN, P1_U3249);
  nand ginst5019 (P1_U4291, P1_REIP_REG_23__SCAN_IN, P1_U4233);
  nand ginst5020 (P1_U4292, P1_REIP_REG_22__SCAN_IN, P1_U4232);
  nand ginst5021 (P1_U4293, P1_ADDRESS_REG_21__SCAN_IN, P1_U3249);
  nand ginst5022 (P1_U4294, P1_REIP_REG_22__SCAN_IN, P1_U4233);
  nand ginst5023 (P1_U4295, P1_REIP_REG_21__SCAN_IN, P1_U4232);
  nand ginst5024 (P1_U4296, P1_ADDRESS_REG_20__SCAN_IN, P1_U3249);
  nand ginst5025 (P1_U4297, P1_REIP_REG_21__SCAN_IN, P1_U4233);
  nand ginst5026 (P1_U4298, P1_REIP_REG_20__SCAN_IN, P1_U4232);
  nand ginst5027 (P1_U4299, P1_ADDRESS_REG_19__SCAN_IN, P1_U3249);
  nand ginst5028 (P1_U4300, P1_REIP_REG_20__SCAN_IN, P1_U4233);
  nand ginst5029 (P1_U4301, P1_REIP_REG_19__SCAN_IN, P1_U4232);
  nand ginst5030 (P1_U4302, P1_ADDRESS_REG_18__SCAN_IN, P1_U3249);
  nand ginst5031 (P1_U4303, P1_REIP_REG_19__SCAN_IN, P1_U4233);
  nand ginst5032 (P1_U4304, P1_REIP_REG_18__SCAN_IN, P1_U4232);
  nand ginst5033 (P1_U4305, P1_ADDRESS_REG_17__SCAN_IN, P1_U3249);
  nand ginst5034 (P1_U4306, P1_REIP_REG_18__SCAN_IN, P1_U4233);
  nand ginst5035 (P1_U4307, P1_REIP_REG_17__SCAN_IN, P1_U4232);
  nand ginst5036 (P1_U4308, P1_ADDRESS_REG_16__SCAN_IN, P1_U3249);
  nand ginst5037 (P1_U4309, P1_REIP_REG_17__SCAN_IN, P1_U4233);
  nand ginst5038 (P1_U4310, P1_REIP_REG_16__SCAN_IN, P1_U4232);
  nand ginst5039 (P1_U4311, P1_ADDRESS_REG_15__SCAN_IN, P1_U3249);
  nand ginst5040 (P1_U4312, P1_REIP_REG_16__SCAN_IN, P1_U4233);
  nand ginst5041 (P1_U4313, P1_REIP_REG_15__SCAN_IN, P1_U4232);
  nand ginst5042 (P1_U4314, P1_ADDRESS_REG_14__SCAN_IN, P1_U3249);
  nand ginst5043 (P1_U4315, P1_REIP_REG_15__SCAN_IN, P1_U4233);
  nand ginst5044 (P1_U4316, P1_REIP_REG_14__SCAN_IN, P1_U4232);
  nand ginst5045 (P1_U4317, P1_ADDRESS_REG_13__SCAN_IN, P1_U3249);
  nand ginst5046 (P1_U4318, P1_REIP_REG_14__SCAN_IN, P1_U4233);
  nand ginst5047 (P1_U4319, P1_REIP_REG_13__SCAN_IN, P1_U4232);
  nand ginst5048 (P1_U4320, P1_ADDRESS_REG_12__SCAN_IN, P1_U3249);
  nand ginst5049 (P1_U4321, P1_REIP_REG_13__SCAN_IN, P1_U4233);
  nand ginst5050 (P1_U4322, P1_REIP_REG_12__SCAN_IN, P1_U4232);
  nand ginst5051 (P1_U4323, P1_ADDRESS_REG_11__SCAN_IN, P1_U3249);
  nand ginst5052 (P1_U4324, P1_REIP_REG_12__SCAN_IN, P1_U4233);
  nand ginst5053 (P1_U4325, P1_REIP_REG_11__SCAN_IN, P1_U4232);
  nand ginst5054 (P1_U4326, P1_ADDRESS_REG_10__SCAN_IN, P1_U3249);
  nand ginst5055 (P1_U4327, P1_REIP_REG_11__SCAN_IN, P1_U4233);
  nand ginst5056 (P1_U4328, P1_REIP_REG_10__SCAN_IN, P1_U4232);
  nand ginst5057 (P1_U4329, P1_ADDRESS_REG_9__SCAN_IN, P1_U3249);
  nand ginst5058 (P1_U4330, P1_REIP_REG_10__SCAN_IN, P1_U4233);
  nand ginst5059 (P1_U4331, P1_REIP_REG_9__SCAN_IN, P1_U4232);
  nand ginst5060 (P1_U4332, P1_ADDRESS_REG_8__SCAN_IN, P1_U3249);
  nand ginst5061 (P1_U4333, P1_REIP_REG_9__SCAN_IN, P1_U4233);
  nand ginst5062 (P1_U4334, P1_REIP_REG_8__SCAN_IN, P1_U4232);
  nand ginst5063 (P1_U4335, P1_ADDRESS_REG_7__SCAN_IN, P1_U3249);
  nand ginst5064 (P1_U4336, P1_REIP_REG_8__SCAN_IN, P1_U4233);
  nand ginst5065 (P1_U4337, P1_REIP_REG_7__SCAN_IN, P1_U4232);
  nand ginst5066 (P1_U4338, P1_ADDRESS_REG_6__SCAN_IN, P1_U3249);
  nand ginst5067 (P1_U4339, P1_REIP_REG_7__SCAN_IN, P1_U4233);
  nand ginst5068 (P1_U4340, P1_REIP_REG_6__SCAN_IN, P1_U4232);
  nand ginst5069 (P1_U4341, P1_ADDRESS_REG_5__SCAN_IN, P1_U3249);
  nand ginst5070 (P1_U4342, P1_REIP_REG_6__SCAN_IN, P1_U4233);
  nand ginst5071 (P1_U4343, P1_REIP_REG_5__SCAN_IN, P1_U4232);
  nand ginst5072 (P1_U4344, P1_ADDRESS_REG_4__SCAN_IN, P1_U3249);
  nand ginst5073 (P1_U4345, P1_REIP_REG_5__SCAN_IN, P1_U4233);
  nand ginst5074 (P1_U4346, P1_REIP_REG_4__SCAN_IN, P1_U4232);
  nand ginst5075 (P1_U4347, P1_ADDRESS_REG_3__SCAN_IN, P1_U3249);
  nand ginst5076 (P1_U4348, P1_REIP_REG_4__SCAN_IN, P1_U4233);
  nand ginst5077 (P1_U4349, P1_REIP_REG_3__SCAN_IN, P1_U4232);
  nand ginst5078 (P1_U4350, P1_ADDRESS_REG_2__SCAN_IN, P1_U3249);
  nand ginst5079 (P1_U4351, P1_REIP_REG_3__SCAN_IN, P1_U4233);
  nand ginst5080 (P1_U4352, P1_REIP_REG_2__SCAN_IN, P1_U4232);
  nand ginst5081 (P1_U4353, P1_ADDRESS_REG_1__SCAN_IN, P1_U3249);
  nand ginst5082 (P1_U4354, P1_REIP_REG_2__SCAN_IN, P1_U4233);
  nand ginst5083 (P1_U4355, P1_REIP_REG_1__SCAN_IN, P1_U4232);
  nand ginst5084 (P1_U4356, P1_ADDRESS_REG_0__SCAN_IN, P1_U3249);
  not ginst5085 (P1_U4357, P1_U3260);
  nand ginst5086 (P1_U4358, P1_U3257, P1_U4357);
  nand ginst5087 (P1_U4359, NA, P1_U4258);
  not ginst5088 (P1_U4360, P1_U3261);
  nand ginst5089 (P1_U4361, P1_U3257, P1_U4360);
  or ginst5090 (P1_U4362, NA, P1_STATE_REG_0__SCAN_IN);
  nand ginst5091 (P1_U4363, P1_U4362, P1_U7622, P1_U7623);
  not ginst5092 (P1_U4364, P1_U3255);
  nand ginst5093 (P1_U4365, HOLD, P1_U3247, P1_U4364);
  nand ginst5094 (P1_U4366, P1_STATE_REG_1__SCAN_IN, P1_U3261, U210);
  nand ginst5095 (P1_U4367, P1_U4365, P1_U4366);
  nand ginst5096 (P1_U4368, P1_STATE_REG_0__SCAN_IN, P1_U4359, P1_U4367);
  nand ginst5097 (P1_U4369, P1_STATE_REG_2__SCAN_IN, P1_U4363);
  nand ginst5098 (P1_U4370, P1_U4221, U210);
  nand ginst5099 (P1_U4371, P1_U3496, P1_U7625);
  nand ginst5100 (P1_U4372, P1_STATE_REG_2__SCAN_IN, P1_U3260);
  nand ginst5101 (P1_U4373, NA, P1_U3258);
  nand ginst5102 (P1_U4374, P1_U4372, P1_U4373);
  nand ginst5103 (P1_U4375, P1_U3248, P1_U4374);
  nand ginst5104 (P1_U4376, P1_U3255, P1_U4179);
  not ginst5105 (P1_U4377, P1_U3280);
  not ginst5106 (P1_U4378, P1_U3269);
  not ginst5107 (P1_U4379, P1_U3444);
  not ginst5108 (P1_U4380, P1_U3268);
  not ginst5109 (P1_U4381, P1_U3274);
  not ginst5110 (P1_U4382, P1_U3267);
  nand ginst5111 (P1_U4383, P1_INSTQUEUE_REG_7__3__SCAN_IN, P1_U4382);
  nand ginst5112 (P1_U4384, P1_INSTQUEUE_REG_0__3__SCAN_IN, P1_U2472);
  nand ginst5113 (P1_U4385, P1_INSTQUEUE_REG_1__3__SCAN_IN, P1_U2471);
  nand ginst5114 (P1_U4386, P1_INSTQUEUE_REG_2__3__SCAN_IN, P1_U2470);
  nand ginst5115 (P1_U4387, P1_INSTQUEUE_REG_3__3__SCAN_IN, P1_U2468);
  nand ginst5116 (P1_U4388, P1_INSTQUEUE_REG_4__3__SCAN_IN, P1_U2467);
  nand ginst5117 (P1_U4389, P1_INSTQUEUE_REG_5__3__SCAN_IN, P1_U2466);
  nand ginst5118 (P1_U4390, P1_INSTQUEUE_REG_6__3__SCAN_IN, P1_U2465);
  nand ginst5119 (P1_U4391, P1_INSTQUEUE_REG_8__3__SCAN_IN, P1_U2464);
  nand ginst5120 (P1_U4392, P1_INSTQUEUE_REG_9__3__SCAN_IN, P1_U2463);
  nand ginst5121 (P1_U4393, P1_INSTQUEUE_REG_10__3__SCAN_IN, P1_U2461);
  nand ginst5122 (P1_U4394, P1_INSTQUEUE_REG_11__3__SCAN_IN, P1_U2459);
  nand ginst5123 (P1_U4395, P1_INSTQUEUE_REG_12__3__SCAN_IN, P1_U2458);
  nand ginst5124 (P1_U4396, P1_INSTQUEUE_REG_13__3__SCAN_IN, P1_U2457);
  nand ginst5125 (P1_U4397, P1_INSTQUEUE_REG_14__3__SCAN_IN, P1_U2455);
  nand ginst5126 (P1_U4398, P1_INSTQUEUE_REG_15__3__SCAN_IN, P1_U2453);
  not ginst5127 (P1_U4399, P1_U3283);
  not ginst5128 (P1_U4400, P1_U3278);
  nand ginst5129 (P1_U4401, P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN, P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN, P1_INSTQUEUE_REG_7__5__SCAN_IN, P1_U3270);
  nand ginst5130 (P1_U4402, P1_INSTQUEUE_REG_0__5__SCAN_IN, P1_U3270, P1_U4380);
  nand ginst5131 (P1_U4403, P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN, P1_INSTQUEUE_REG_1__5__SCAN_IN, P1_U2469, P1_U3265);
  nand ginst5132 (P1_U4404, P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P1_INSTQUEUE_REG_2__5__SCAN_IN, P1_U2469, P1_U3266);
  nand ginst5133 (P1_U4405, P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN, P1_INSTQUEUE_REG_4__5__SCAN_IN, P1_U3270, P1_U4378);
  nand ginst5134 (P1_U4406, P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN, P1_U3520, P1_U3521);
  nand ginst5135 (P1_U4407, P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN, P1_U3522, P1_U3523);
  nand ginst5136 (P1_U4408, P1_U3524, P1_U4380);
  nand ginst5137 (P1_U4409, P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P1_U3525, P1_U3526);
  nand ginst5138 (P1_U4410, P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN, P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P1_INSTQUEUE_REG_11__5__SCAN_IN, P1_U3264);
  nand ginst5139 (P1_U4411, P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN, P1_U3527, P1_U4378);
  nand ginst5140 (P1_U4412, P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN, P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN, P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P1_INSTQUEUE_REG_13__5__SCAN_IN, P1_U3265);
  nand ginst5141 (P1_U4413, P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN, P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P1_INSTQUEUE_REG_14__5__SCAN_IN, P1_U3266);
  nand ginst5142 (P1_U4414, P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN, P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN, P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P1_INSTQUEUE_REG_15__5__SCAN_IN);
  not ginst5143 (P1_U4415, P1_U4173);
  nand ginst5144 (P1_U4416, P1_INSTQUEUE_REG_7__2__SCAN_IN, P1_U4382);
  nand ginst5145 (P1_U4417, P1_INSTQUEUE_REG_0__2__SCAN_IN, P1_U2472);
  nand ginst5146 (P1_U4418, P1_INSTQUEUE_REG_1__2__SCAN_IN, P1_U2471);
  nand ginst5147 (P1_U4419, P1_INSTQUEUE_REG_2__2__SCAN_IN, P1_U2470);
  nand ginst5148 (P1_U4420, P1_INSTQUEUE_REG_3__2__SCAN_IN, P1_U2468);
  nand ginst5149 (P1_U4421, P1_INSTQUEUE_REG_4__2__SCAN_IN, P1_U2467);
  nand ginst5150 (P1_U4422, P1_INSTQUEUE_REG_5__2__SCAN_IN, P1_U2466);
  nand ginst5151 (P1_U4423, P1_INSTQUEUE_REG_6__2__SCAN_IN, P1_U2465);
  nand ginst5152 (P1_U4424, P1_INSTQUEUE_REG_8__2__SCAN_IN, P1_U2464);
  nand ginst5153 (P1_U4425, P1_INSTQUEUE_REG_9__2__SCAN_IN, P1_U2463);
  nand ginst5154 (P1_U4426, P1_INSTQUEUE_REG_10__2__SCAN_IN, P1_U2461);
  nand ginst5155 (P1_U4427, P1_INSTQUEUE_REG_11__2__SCAN_IN, P1_U2459);
  nand ginst5156 (P1_U4428, P1_INSTQUEUE_REG_12__2__SCAN_IN, P1_U2458);
  nand ginst5157 (P1_U4429, P1_INSTQUEUE_REG_13__2__SCAN_IN, P1_U2457);
  nand ginst5158 (P1_U4430, P1_INSTQUEUE_REG_14__2__SCAN_IN, P1_U2455);
  nand ginst5159 (P1_U4431, P1_INSTQUEUE_REG_15__2__SCAN_IN, P1_U2453);
  not ginst5160 (P1_U4432, P1_U4171);
  nand ginst5161 (P1_U4433, P1_INSTQUEUE_REG_7__7__SCAN_IN, P1_U4382);
  nand ginst5162 (P1_U4434, P1_INSTQUEUE_REG_0__7__SCAN_IN, P1_U2472);
  nand ginst5163 (P1_U4435, P1_INSTQUEUE_REG_1__7__SCAN_IN, P1_U2471);
  nand ginst5164 (P1_U4436, P1_INSTQUEUE_REG_2__7__SCAN_IN, P1_U2470);
  nand ginst5165 (P1_U4437, P1_INSTQUEUE_REG_3__7__SCAN_IN, P1_U2468);
  nand ginst5166 (P1_U4438, P1_INSTQUEUE_REG_4__7__SCAN_IN, P1_U2467);
  nand ginst5167 (P1_U4439, P1_INSTQUEUE_REG_5__7__SCAN_IN, P1_U2466);
  nand ginst5168 (P1_U4440, P1_INSTQUEUE_REG_6__7__SCAN_IN, P1_U2465);
  nand ginst5169 (P1_U4441, P1_INSTQUEUE_REG_8__7__SCAN_IN, P1_U2464);
  nand ginst5170 (P1_U4442, P1_INSTQUEUE_REG_9__7__SCAN_IN, P1_U2463);
  nand ginst5171 (P1_U4443, P1_INSTQUEUE_REG_10__7__SCAN_IN, P1_U2461);
  nand ginst5172 (P1_U4444, P1_INSTQUEUE_REG_11__7__SCAN_IN, P1_U2459);
  nand ginst5173 (P1_U4445, P1_INSTQUEUE_REG_12__7__SCAN_IN, P1_U2458);
  nand ginst5174 (P1_U4446, P1_INSTQUEUE_REG_13__7__SCAN_IN, P1_U2457);
  nand ginst5175 (P1_U4447, P1_INSTQUEUE_REG_14__7__SCAN_IN, P1_U2455);
  nand ginst5176 (P1_U4448, P1_INSTQUEUE_REG_15__7__SCAN_IN, P1_U2453);
  not ginst5177 (P1_U4449, P1_U3391);
  nand ginst5178 (P1_U4450, P1_INSTQUEUE_REG_7__6__SCAN_IN, P1_U3498, P1_U4381);
  nand ginst5179 (P1_U4451, P1_INSTQUEUE_REG_1__6__SCAN_IN, P1_U2456, P1_U2469);
  nand ginst5180 (P1_U4452, P1_INSTQUEUE_REG_2__6__SCAN_IN, P1_U2454, P1_U2469);
  nand ginst5181 (P1_U4453, P1_INSTQUEUE_REG_4__6__SCAN_IN, P1_U4378, P1_U4381);
  nand ginst5182 (P1_U4454, P1_INSTQUEUE_REG_5__6__SCAN_IN, P1_U2456, P1_U4381);
  nand ginst5183 (P1_U4455, P1_INSTQUEUE_REG_6__6__SCAN_IN, P1_U2454, P1_U4381);
  nand ginst5184 (P1_U4456, P1_INSTQUEUE_REG_12__6__SCAN_IN, P1_U3507, P1_U4378);
  nand ginst5185 (P1_U4457, P1_INSTQUEUE_REG_13__6__SCAN_IN, P1_U2456, P1_U3507);
  nand ginst5186 (P1_U4458, P1_INSTQUEUE_REG_14__6__SCAN_IN, P1_U2454, P1_U3507);
  nand ginst5187 (P1_U4459, P1_INSTQUEUE_REG_15__6__SCAN_IN, P1_U3498, P1_U3507);
  not ginst5188 (P1_U4460, P1_U3277);
  nand ginst5189 (P1_U4461, P1_INSTQUEUE_REG_7__1__SCAN_IN, P1_U4382);
  nand ginst5190 (P1_U4462, P1_INSTQUEUE_REG_0__1__SCAN_IN, P1_U2472);
  nand ginst5191 (P1_U4463, P1_INSTQUEUE_REG_1__1__SCAN_IN, P1_U2471);
  nand ginst5192 (P1_U4464, P1_INSTQUEUE_REG_2__1__SCAN_IN, P1_U2470);
  nand ginst5193 (P1_U4465, P1_INSTQUEUE_REG_3__1__SCAN_IN, P1_U2468);
  nand ginst5194 (P1_U4466, P1_INSTQUEUE_REG_4__1__SCAN_IN, P1_U2467);
  nand ginst5195 (P1_U4467, P1_INSTQUEUE_REG_5__1__SCAN_IN, P1_U2466);
  nand ginst5196 (P1_U4468, P1_INSTQUEUE_REG_6__1__SCAN_IN, P1_U2465);
  nand ginst5197 (P1_U4469, P1_INSTQUEUE_REG_8__1__SCAN_IN, P1_U2464);
  nand ginst5198 (P1_U4470, P1_INSTQUEUE_REG_9__1__SCAN_IN, P1_U2463);
  nand ginst5199 (P1_U4471, P1_INSTQUEUE_REG_10__1__SCAN_IN, P1_U2461);
  nand ginst5200 (P1_U4472, P1_INSTQUEUE_REG_11__1__SCAN_IN, P1_U2459);
  nand ginst5201 (P1_U4473, P1_INSTQUEUE_REG_12__1__SCAN_IN, P1_U2458);
  nand ginst5202 (P1_U4474, P1_INSTQUEUE_REG_13__1__SCAN_IN, P1_U2457);
  nand ginst5203 (P1_U4475, P1_INSTQUEUE_REG_14__1__SCAN_IN, P1_U2455);
  nand ginst5204 (P1_U4476, P1_INSTQUEUE_REG_15__1__SCAN_IN, P1_U2453);
  not ginst5205 (P1_U4477, P1_U3271);
  nand ginst5206 (P1_U4478, P1_INSTQUEUE_REG_7__0__SCAN_IN, P1_U4382);
  nand ginst5207 (P1_U4479, P1_INSTQUEUE_REG_0__0__SCAN_IN, P1_U2472);
  nand ginst5208 (P1_U4480, P1_INSTQUEUE_REG_1__0__SCAN_IN, P1_U2471);
  nand ginst5209 (P1_U4481, P1_INSTQUEUE_REG_2__0__SCAN_IN, P1_U2470);
  nand ginst5210 (P1_U4482, P1_INSTQUEUE_REG_3__0__SCAN_IN, P1_U2468);
  nand ginst5211 (P1_U4483, P1_INSTQUEUE_REG_4__0__SCAN_IN, P1_U2467);
  nand ginst5212 (P1_U4484, P1_INSTQUEUE_REG_5__0__SCAN_IN, P1_U2466);
  nand ginst5213 (P1_U4485, P1_INSTQUEUE_REG_6__0__SCAN_IN, P1_U2465);
  nand ginst5214 (P1_U4486, P1_INSTQUEUE_REG_8__0__SCAN_IN, P1_U2464);
  nand ginst5215 (P1_U4487, P1_INSTQUEUE_REG_9__0__SCAN_IN, P1_U2463);
  nand ginst5216 (P1_U4488, P1_INSTQUEUE_REG_10__0__SCAN_IN, P1_U2461);
  nand ginst5217 (P1_U4489, P1_INSTQUEUE_REG_11__0__SCAN_IN, P1_U2459);
  nand ginst5218 (P1_U4490, P1_INSTQUEUE_REG_12__0__SCAN_IN, P1_U2458);
  nand ginst5219 (P1_U4491, P1_INSTQUEUE_REG_13__0__SCAN_IN, P1_U2457);
  nand ginst5220 (P1_U4492, P1_INSTQUEUE_REG_14__0__SCAN_IN, P1_U2455);
  nand ginst5221 (P1_U4493, P1_INSTQUEUE_REG_15__0__SCAN_IN, P1_U2453);
  not ginst5222 (P1_U4494, P1_U3284);
  nand ginst5223 (P1_U4495, P1_STATE_REG_2__SCAN_IN, P1_U3248);
  nand ginst5224 (P1_U4496, P1_U3254, P1_U4495);
  not ginst5225 (P1_U4497, P1_U3272);
  nand ginst5226 (P1_U4498, P1_U3388, P1_U4477);
  not ginst5227 (P1_U4499, P1_U3437);
  nand ginst5228 (P1_U4500, P1_U3272, P1_U3287, P1_U3390);
  nand ginst5229 (P1_U4501, P1_U3257, P1_U4500);
  not ginst5230 (P1_U4502, P1_U3285);
  nand ginst5231 (P1_U4503, P1_U4173, P1_U4460);
  nand ginst5232 (P1_U4504, P1_U3286, P1_U4196);
  nand ginst5233 (P1_U4505, P1_U3579, P1_U4504);
  nand ginst5234 (P1_U4506, P1_U3580, P1_U4505);
  nand ginst5235 (P1_U4507, P1_U3388, P1_U4215);
  nand ginst5236 (P1_U4508, P1_U4507, P1_U7681, P1_U7682);
  nand ginst5237 (P1_U4509, P1_U2448, P1_U4262);
  or ginst5238 (P1_U4510, P1_MORE_REG_SCAN_IN, P1_FLUSH_REG_SCAN_IN);
  not ginst5239 (P1_U4511, P1_U3293);
  nand ginst5240 (P1_U4512, P1_U3262, P1_U4511);
  nand ginst5241 (P1_U4513, P1_STATE2_REG_1__SCAN_IN, U210);
  not ginst5242 (P1_U4514, P1_U3295);
  nand ginst5243 (P1_U4515, P1_STATE2_REG_1__SCAN_IN, P1_U7687, P1_U7688);
  nand ginst5244 (P1_U4516, P1_STATE2_REG_2__SCAN_IN, P1_U3295);
  nand ginst5245 (P1_U4517, P1_U4246, P1_U7604);
  nand ginst5246 (P1_U4518, P1_U3583, P1_U4514);
  nand ginst5247 (P1_U4519, P1_STATE2_REG_1__SCAN_IN, P1_U4517);
  nand ginst5248 (P1_U4520, P1_U2368, P1_U7604);
  nand ginst5249 (P1_U4521, P1_U4252, P1_U4261);
  nand ginst5250 (P1_U4522, P1_U4245, P1_U7604);
  nand ginst5251 (P1_U4523, P1_U2368, P1_U3293);
  not ginst5252 (P1_U4524, P1_U3325);
  not ginst5253 (P1_U4525, P1_U3331);
  not ginst5254 (P1_U4526, P1_U3332);
  not ginst5255 (P1_U4527, P1_U3314);
  not ginst5256 (P1_U4528, P1_U3313);
  not ginst5257 (P1_U4529, P1_U3342);
  nand ginst5258 (P1_U4530, P1_R2144_U8, P1_U3313);
  not ginst5259 (P1_U4531, P1_U3358);
  not ginst5260 (P1_U4532, P1_U3315);
  not ginst5261 (P1_U4533, P1_U3305);
  not ginst5262 (P1_U4534, P1_U3306);
  nand ginst5263 (P1_U4535, P1_U2438, P1_U2442);
  not ginst5264 (P1_U4536, P1_U3321);
  not ginst5265 (P1_U4537, P1_U3356);
  not ginst5266 (P1_U4538, P1_U3340);
  nand ginst5267 (P1_U4539, P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN, P1_U3305);
  not ginst5268 (P1_U4540, P1_U3360);
  not ginst5269 (P1_U4541, P1_U3329);
  not ginst5270 (P1_U4542, P1_U3323);
  not ginst5271 (P1_U4543, P1_U3235);
  nand ginst5272 (P1_U4544, P1_U2432, P1_U2436);
  not ginst5273 (P1_U4545, P1_U3322);
  nand ginst5274 (P1_U4546, P1_STATE2_REG_1__SCAN_IN, P1_U3263);
  nand ginst5275 (P1_U4547, P1_U3297, P1_U3299, P1_U4546);
  nand ginst5276 (P1_U4548, P1_U2476, P1_U4528);
  nand ginst5277 (P1_U4549, P1_U2358, P1_U2480);
  nand ginst5278 (P1_U4550, P1_U3320, P1_U4549);
  nand ginst5279 (P1_U4551, P1_U4536, P1_U4550);
  nand ginst5280 (P1_U4552, P1_STATE2_REG_3__SCAN_IN, P1_U3306);
  nand ginst5281 (P1_U4553, P1_STATE2_REG_2__SCAN_IN, P1_U4545);
  nand ginst5282 (P1_U4554, P1_U3587, P1_U4551);
  nand ginst5283 (P1_U4555, P1_U2388, P1_U2480);
  nand ginst5284 (P1_U4556, P1_U3320, P1_U4555);
  nand ginst5285 (P1_U4557, P1_U3321, P1_U4556);
  nand ginst5286 (P1_U4558, P1_STATE2_REG_2__SCAN_IN, P1_U3322);
  nand ginst5287 (P1_U4559, P1_U4557, P1_U4558);
  nand ginst5288 (P1_U4560, P1_U2415, P1_U4534);
  nand ginst5289 (P1_U4561, P1_U2413, P1_U2477);
  nand ginst5290 (P1_U4562, P1_U2412, P1_U4532);
  nand ginst5291 (P1_U4563, P1_U2397, P1_U4559);
  nand ginst5292 (P1_U4564, P1_INSTQUEUE_REG_15__7__SCAN_IN, P1_U4554);
  nand ginst5293 (P1_U4565, P1_U2416, P1_U4534);
  nand ginst5294 (P1_U4566, P1_U2411, P1_U2477);
  nand ginst5295 (P1_U4567, P1_U2410, P1_U4532);
  nand ginst5296 (P1_U4568, P1_U2396, P1_U4559);
  nand ginst5297 (P1_U4569, P1_INSTQUEUE_REG_15__6__SCAN_IN, P1_U4554);
  nand ginst5298 (P1_U4570, P1_U2420, P1_U4534);
  nand ginst5299 (P1_U4571, P1_U2409, P1_U2477);
  nand ginst5300 (P1_U4572, P1_U2408, P1_U4532);
  nand ginst5301 (P1_U4573, P1_U2395, P1_U4559);
  nand ginst5302 (P1_U4574, P1_INSTQUEUE_REG_15__5__SCAN_IN, P1_U4554);
  nand ginst5303 (P1_U4575, P1_U2419, P1_U4534);
  nand ginst5304 (P1_U4576, P1_U2407, P1_U2477);
  nand ginst5305 (P1_U4577, P1_U2406, P1_U4532);
  nand ginst5306 (P1_U4578, P1_U2394, P1_U4559);
  nand ginst5307 (P1_U4579, P1_INSTQUEUE_REG_15__4__SCAN_IN, P1_U4554);
  nand ginst5308 (P1_U4580, P1_U2418, P1_U4534);
  nand ginst5309 (P1_U4581, P1_U2405, P1_U2477);
  nand ginst5310 (P1_U4582, P1_U2404, P1_U4532);
  nand ginst5311 (P1_U4583, P1_U2393, P1_U4559);
  nand ginst5312 (P1_U4584, P1_INSTQUEUE_REG_15__3__SCAN_IN, P1_U4554);
  nand ginst5313 (P1_U4585, P1_U2421, P1_U4534);
  nand ginst5314 (P1_U4586, P1_U2403, P1_U2477);
  nand ginst5315 (P1_U4587, P1_U2402, P1_U4532);
  nand ginst5316 (P1_U4588, P1_U2392, P1_U4559);
  nand ginst5317 (P1_U4589, P1_INSTQUEUE_REG_15__2__SCAN_IN, P1_U4554);
  nand ginst5318 (P1_U4590, P1_U2414, P1_U4534);
  nand ginst5319 (P1_U4591, P1_U2401, P1_U2477);
  nand ginst5320 (P1_U4592, P1_U2400, P1_U4532);
  nand ginst5321 (P1_U4593, P1_U2391, P1_U4559);
  nand ginst5322 (P1_U4594, P1_INSTQUEUE_REG_15__1__SCAN_IN, P1_U4554);
  nand ginst5323 (P1_U4595, P1_U2417, P1_U4534);
  nand ginst5324 (P1_U4596, P1_U2399, P1_U2477);
  nand ginst5325 (P1_U4597, P1_U2398, P1_U4532);
  nand ginst5326 (P1_U4598, P1_U2390, P1_U4559);
  nand ginst5327 (P1_U4599, P1_INSTQUEUE_REG_15__0__SCAN_IN, P1_U4554);
  not ginst5328 (P1_U4600, P1_U3326);
  not ginst5329 (P1_U4601, P1_U3327);
  not ginst5330 (P1_U4602, P1_U3324);
  nand ginst5331 (P1_U4603, P1_U2438, P1_U2443);
  not ginst5332 (P1_U4604, P1_U3328);
  not ginst5333 (P1_U4605, P1_U3236);
  nand ginst5334 (P1_U4606, P1_U2476, P1_U4524);
  nand ginst5335 (P1_U4607, P1_U2358, P1_U2482);
  nand ginst5336 (P1_U4608, P1_U3320, P1_U4607);
  nand ginst5337 (P1_U4609, P1_U4604, P1_U4608);
  nand ginst5338 (P1_U4610, P1_STATE2_REG_3__SCAN_IN, P1_U3324);
  nand ginst5339 (P1_U4611, P1_STATE2_REG_2__SCAN_IN, P1_U3236);
  nand ginst5340 (P1_U4612, P1_U3596, P1_U4609);
  nand ginst5341 (P1_U4613, P1_U2388, P1_U2482);
  nand ginst5342 (P1_U4614, P1_U3320, P1_U4613);
  nand ginst5343 (P1_U4615, P1_U3328, P1_U4614);
  nand ginst5344 (P1_U4616, P1_STATE2_REG_2__SCAN_IN, P1_U4605);
  nand ginst5345 (P1_U4617, P1_U4615, P1_U4616);
  nand ginst5346 (P1_U4618, P1_U2415, P1_U4602);
  nand ginst5347 (P1_U4619, P1_U2413, P1_U2481);
  nand ginst5348 (P1_U4620, P1_U2412, P1_U4601);
  nand ginst5349 (P1_U4621, P1_U2397, P1_U4617);
  nand ginst5350 (P1_U4622, P1_INSTQUEUE_REG_14__7__SCAN_IN, P1_U4612);
  nand ginst5351 (P1_U4623, P1_U2416, P1_U4602);
  nand ginst5352 (P1_U4624, P1_U2411, P1_U2481);
  nand ginst5353 (P1_U4625, P1_U2410, P1_U4601);
  nand ginst5354 (P1_U4626, P1_U2396, P1_U4617);
  nand ginst5355 (P1_U4627, P1_INSTQUEUE_REG_14__6__SCAN_IN, P1_U4612);
  nand ginst5356 (P1_U4628, P1_U2420, P1_U4602);
  nand ginst5357 (P1_U4629, P1_U2409, P1_U2481);
  nand ginst5358 (P1_U4630, P1_U2408, P1_U4601);
  nand ginst5359 (P1_U4631, P1_U2395, P1_U4617);
  nand ginst5360 (P1_U4632, P1_INSTQUEUE_REG_14__5__SCAN_IN, P1_U4612);
  nand ginst5361 (P1_U4633, P1_U2419, P1_U4602);
  nand ginst5362 (P1_U4634, P1_U2407, P1_U2481);
  nand ginst5363 (P1_U4635, P1_U2406, P1_U4601);
  nand ginst5364 (P1_U4636, P1_U2394, P1_U4617);
  nand ginst5365 (P1_U4637, P1_INSTQUEUE_REG_14__4__SCAN_IN, P1_U4612);
  nand ginst5366 (P1_U4638, P1_U2418, P1_U4602);
  nand ginst5367 (P1_U4639, P1_U2405, P1_U2481);
  nand ginst5368 (P1_U4640, P1_U2404, P1_U4601);
  nand ginst5369 (P1_U4641, P1_U2393, P1_U4617);
  nand ginst5370 (P1_U4642, P1_INSTQUEUE_REG_14__3__SCAN_IN, P1_U4612);
  nand ginst5371 (P1_U4643, P1_U2421, P1_U4602);
  nand ginst5372 (P1_U4644, P1_U2403, P1_U2481);
  nand ginst5373 (P1_U4645, P1_U2402, P1_U4601);
  nand ginst5374 (P1_U4646, P1_U2392, P1_U4617);
  nand ginst5375 (P1_U4647, P1_INSTQUEUE_REG_14__2__SCAN_IN, P1_U4612);
  nand ginst5376 (P1_U4648, P1_U2414, P1_U4602);
  nand ginst5377 (P1_U4649, P1_U2401, P1_U2481);
  nand ginst5378 (P1_U4650, P1_U2400, P1_U4601);
  nand ginst5379 (P1_U4651, P1_U2391, P1_U4617);
  nand ginst5380 (P1_U4652, P1_INSTQUEUE_REG_14__1__SCAN_IN, P1_U4612);
  nand ginst5381 (P1_U4653, P1_U2417, P1_U4602);
  nand ginst5382 (P1_U4654, P1_U2399, P1_U2481);
  nand ginst5383 (P1_U4655, P1_U2398, P1_U4601);
  nand ginst5384 (P1_U4656, P1_U2390, P1_U4617);
  nand ginst5385 (P1_U4657, P1_INSTQUEUE_REG_14__0__SCAN_IN, P1_U4612);
  not ginst5386 (P1_U4658, P1_U3333);
  not ginst5387 (P1_U4659, P1_U3334);
  not ginst5388 (P1_U4660, P1_U3330);
  nand ginst5389 (P1_U4661, P1_U2438, P1_U2444);
  not ginst5390 (P1_U4662, P1_U3335);
  nand ginst5391 (P1_U4663, P1_U2432, P1_U2437);
  not ginst5392 (P1_U4664, P1_U3336);
  nand ginst5393 (P1_U4665, P1_U2476, P1_U4525);
  nand ginst5394 (P1_U4666, P1_U2358, P1_U2484);
  nand ginst5395 (P1_U4667, P1_U3320, P1_U4666);
  nand ginst5396 (P1_U4668, P1_U4662, P1_U4667);
  nand ginst5397 (P1_U4669, P1_STATE2_REG_3__SCAN_IN, P1_U3330);
  nand ginst5398 (P1_U4670, P1_STATE2_REG_2__SCAN_IN, P1_U4664);
  nand ginst5399 (P1_U4671, P1_U3605, P1_U4668);
  nand ginst5400 (P1_U4672, P1_U2388, P1_U2484);
  nand ginst5401 (P1_U4673, P1_U3320, P1_U4672);
  nand ginst5402 (P1_U4674, P1_U3335, P1_U4673);
  nand ginst5403 (P1_U4675, P1_STATE2_REG_2__SCAN_IN, P1_U3336);
  nand ginst5404 (P1_U4676, P1_U4674, P1_U4675);
  nand ginst5405 (P1_U4677, P1_U2415, P1_U4660);
  nand ginst5406 (P1_U4678, P1_U2413, P1_U2483);
  nand ginst5407 (P1_U4679, P1_U2412, P1_U4659);
  nand ginst5408 (P1_U4680, P1_U2397, P1_U4676);
  nand ginst5409 (P1_U4681, P1_INSTQUEUE_REG_13__7__SCAN_IN, P1_U4671);
  nand ginst5410 (P1_U4682, P1_U2416, P1_U4660);
  nand ginst5411 (P1_U4683, P1_U2411, P1_U2483);
  nand ginst5412 (P1_U4684, P1_U2410, P1_U4659);
  nand ginst5413 (P1_U4685, P1_U2396, P1_U4676);
  nand ginst5414 (P1_U4686, P1_INSTQUEUE_REG_13__6__SCAN_IN, P1_U4671);
  nand ginst5415 (P1_U4687, P1_U2420, P1_U4660);
  nand ginst5416 (P1_U4688, P1_U2409, P1_U2483);
  nand ginst5417 (P1_U4689, P1_U2408, P1_U4659);
  nand ginst5418 (P1_U4690, P1_U2395, P1_U4676);
  nand ginst5419 (P1_U4691, P1_INSTQUEUE_REG_13__5__SCAN_IN, P1_U4671);
  nand ginst5420 (P1_U4692, P1_U2419, P1_U4660);
  nand ginst5421 (P1_U4693, P1_U2407, P1_U2483);
  nand ginst5422 (P1_U4694, P1_U2406, P1_U4659);
  nand ginst5423 (P1_U4695, P1_U2394, P1_U4676);
  nand ginst5424 (P1_U4696, P1_INSTQUEUE_REG_13__4__SCAN_IN, P1_U4671);
  nand ginst5425 (P1_U4697, P1_U2418, P1_U4660);
  nand ginst5426 (P1_U4698, P1_U2405, P1_U2483);
  nand ginst5427 (P1_U4699, P1_U2404, P1_U4659);
  nand ginst5428 (P1_U4700, P1_U2393, P1_U4676);
  nand ginst5429 (P1_U4701, P1_INSTQUEUE_REG_13__3__SCAN_IN, P1_U4671);
  nand ginst5430 (P1_U4702, P1_U2421, P1_U4660);
  nand ginst5431 (P1_U4703, P1_U2403, P1_U2483);
  nand ginst5432 (P1_U4704, P1_U2402, P1_U4659);
  nand ginst5433 (P1_U4705, P1_U2392, P1_U4676);
  nand ginst5434 (P1_U4706, P1_INSTQUEUE_REG_13__2__SCAN_IN, P1_U4671);
  nand ginst5435 (P1_U4707, P1_U2414, P1_U4660);
  nand ginst5436 (P1_U4708, P1_U2401, P1_U2483);
  nand ginst5437 (P1_U4709, P1_U2400, P1_U4659);
  nand ginst5438 (P1_U4710, P1_U2391, P1_U4676);
  nand ginst5439 (P1_U4711, P1_INSTQUEUE_REG_13__1__SCAN_IN, P1_U4671);
  nand ginst5440 (P1_U4712, P1_U2417, P1_U4660);
  nand ginst5441 (P1_U4713, P1_U2399, P1_U2483);
  nand ginst5442 (P1_U4714, P1_U2398, P1_U4659);
  nand ginst5443 (P1_U4715, P1_U2390, P1_U4676);
  nand ginst5444 (P1_U4716, P1_INSTQUEUE_REG_13__0__SCAN_IN, P1_U4671);
  not ginst5445 (P1_U4717, P1_U3338);
  not ginst5446 (P1_U4718, P1_U3337);
  nand ginst5447 (P1_U4719, P1_U2438, P1_U2445);
  not ginst5448 (P1_U4720, P1_U3339);
  not ginst5449 (P1_U4721, P1_U3237);
  nand ginst5450 (P1_U4722, P1_U2476, P1_U2486);
  nand ginst5451 (P1_U4723, P1_U2358, P1_U2489);
  nand ginst5452 (P1_U4724, P1_U3320, P1_U4723);
  nand ginst5453 (P1_U4725, P1_U4720, P1_U4724);
  nand ginst5454 (P1_U4726, P1_STATE2_REG_3__SCAN_IN, P1_U3337);
  nand ginst5455 (P1_U4727, P1_STATE2_REG_2__SCAN_IN, P1_U3237);
  nand ginst5456 (P1_U4728, P1_U3614, P1_U4725);
  nand ginst5457 (P1_U4729, P1_U2388, P1_U2489);
  nand ginst5458 (P1_U4730, P1_U3320, P1_U4729);
  nand ginst5459 (P1_U4731, P1_U3339, P1_U4730);
  nand ginst5460 (P1_U4732, P1_STATE2_REG_2__SCAN_IN, P1_U4721);
  nand ginst5461 (P1_U4733, P1_U4731, P1_U4732);
  nand ginst5462 (P1_U4734, P1_U2415, P1_U4718);
  nand ginst5463 (P1_U4735, P1_U2413, P1_U2487);
  nand ginst5464 (P1_U4736, P1_U2412, P1_U4717);
  nand ginst5465 (P1_U4737, P1_U2397, P1_U4733);
  nand ginst5466 (P1_U4738, P1_INSTQUEUE_REG_12__7__SCAN_IN, P1_U4728);
  nand ginst5467 (P1_U4739, P1_U2416, P1_U4718);
  nand ginst5468 (P1_U4740, P1_U2411, P1_U2487);
  nand ginst5469 (P1_U4741, P1_U2410, P1_U4717);
  nand ginst5470 (P1_U4742, P1_U2396, P1_U4733);
  nand ginst5471 (P1_U4743, P1_INSTQUEUE_REG_12__6__SCAN_IN, P1_U4728);
  nand ginst5472 (P1_U4744, P1_U2420, P1_U4718);
  nand ginst5473 (P1_U4745, P1_U2409, P1_U2487);
  nand ginst5474 (P1_U4746, P1_U2408, P1_U4717);
  nand ginst5475 (P1_U4747, P1_U2395, P1_U4733);
  nand ginst5476 (P1_U4748, P1_INSTQUEUE_REG_12__5__SCAN_IN, P1_U4728);
  nand ginst5477 (P1_U4749, P1_U2419, P1_U4718);
  nand ginst5478 (P1_U4750, P1_U2407, P1_U2487);
  nand ginst5479 (P1_U4751, P1_U2406, P1_U4717);
  nand ginst5480 (P1_U4752, P1_U2394, P1_U4733);
  nand ginst5481 (P1_U4753, P1_INSTQUEUE_REG_12__4__SCAN_IN, P1_U4728);
  nand ginst5482 (P1_U4754, P1_U2418, P1_U4718);
  nand ginst5483 (P1_U4755, P1_U2405, P1_U2487);
  nand ginst5484 (P1_U4756, P1_U2404, P1_U4717);
  nand ginst5485 (P1_U4757, P1_U2393, P1_U4733);
  nand ginst5486 (P1_U4758, P1_INSTQUEUE_REG_12__3__SCAN_IN, P1_U4728);
  nand ginst5487 (P1_U4759, P1_U2421, P1_U4718);
  nand ginst5488 (P1_U4760, P1_U2403, P1_U2487);
  nand ginst5489 (P1_U4761, P1_U2402, P1_U4717);
  nand ginst5490 (P1_U4762, P1_U2392, P1_U4733);
  nand ginst5491 (P1_U4763, P1_INSTQUEUE_REG_12__2__SCAN_IN, P1_U4728);
  nand ginst5492 (P1_U4764, P1_U2414, P1_U4718);
  nand ginst5493 (P1_U4765, P1_U2401, P1_U2487);
  nand ginst5494 (P1_U4766, P1_U2400, P1_U4717);
  nand ginst5495 (P1_U4767, P1_U2391, P1_U4733);
  nand ginst5496 (P1_U4768, P1_INSTQUEUE_REG_12__1__SCAN_IN, P1_U4728);
  nand ginst5497 (P1_U4769, P1_U2417, P1_U4718);
  nand ginst5498 (P1_U4770, P1_U2399, P1_U2487);
  nand ginst5499 (P1_U4771, P1_U2398, P1_U4717);
  nand ginst5500 (P1_U4772, P1_U2390, P1_U4733);
  nand ginst5501 (P1_U4773, P1_INSTQUEUE_REG_12__0__SCAN_IN, P1_U4728);
  not ginst5502 (P1_U4774, P1_U3343);
  not ginst5503 (P1_U4775, P1_U3341);
  nand ginst5504 (P1_U4776, P1_U2440, P1_U2442);
  not ginst5505 (P1_U4777, P1_U3344);
  nand ginst5506 (P1_U4778, P1_U2434, P1_U2436);
  not ginst5507 (P1_U4779, P1_U3345);
  nand ginst5508 (P1_U4780, P1_U4528, P1_U4529);
  nand ginst5509 (P1_U4781, P1_U2358, P1_U2492);
  nand ginst5510 (P1_U4782, P1_U3320, P1_U4781);
  nand ginst5511 (P1_U4783, P1_U4777, P1_U4782);
  nand ginst5512 (P1_U4784, P1_STATE2_REG_3__SCAN_IN, P1_U3341);
  nand ginst5513 (P1_U4785, P1_STATE2_REG_2__SCAN_IN, P1_U4779);
  nand ginst5514 (P1_U4786, P1_U3623, P1_U4783);
  nand ginst5515 (P1_U4787, P1_U2388, P1_U2492);
  nand ginst5516 (P1_U4788, P1_U3320, P1_U4787);
  nand ginst5517 (P1_U4789, P1_U3344, P1_U4788);
  nand ginst5518 (P1_U4790, P1_STATE2_REG_2__SCAN_IN, P1_U3345);
  nand ginst5519 (P1_U4791, P1_U4789, P1_U4790);
  nand ginst5520 (P1_U4792, P1_U2415, P1_U4775);
  nand ginst5521 (P1_U4793, P1_U2413, P1_U2491);
  nand ginst5522 (P1_U4794, P1_U2412, P1_U4774);
  nand ginst5523 (P1_U4795, P1_U2397, P1_U4791);
  nand ginst5524 (P1_U4796, P1_INSTQUEUE_REG_11__7__SCAN_IN, P1_U4786);
  nand ginst5525 (P1_U4797, P1_U2416, P1_U4775);
  nand ginst5526 (P1_U4798, P1_U2411, P1_U2491);
  nand ginst5527 (P1_U4799, P1_U2410, P1_U4774);
  nand ginst5528 (P1_U4800, P1_U2396, P1_U4791);
  nand ginst5529 (P1_U4801, P1_INSTQUEUE_REG_11__6__SCAN_IN, P1_U4786);
  nand ginst5530 (P1_U4802, P1_U2420, P1_U4775);
  nand ginst5531 (P1_U4803, P1_U2409, P1_U2491);
  nand ginst5532 (P1_U4804, P1_U2408, P1_U4774);
  nand ginst5533 (P1_U4805, P1_U2395, P1_U4791);
  nand ginst5534 (P1_U4806, P1_INSTQUEUE_REG_11__5__SCAN_IN, P1_U4786);
  nand ginst5535 (P1_U4807, P1_U2419, P1_U4775);
  nand ginst5536 (P1_U4808, P1_U2407, P1_U2491);
  nand ginst5537 (P1_U4809, P1_U2406, P1_U4774);
  nand ginst5538 (P1_U4810, P1_U2394, P1_U4791);
  nand ginst5539 (P1_U4811, P1_INSTQUEUE_REG_11__4__SCAN_IN, P1_U4786);
  nand ginst5540 (P1_U4812, P1_U2418, P1_U4775);
  nand ginst5541 (P1_U4813, P1_U2405, P1_U2491);
  nand ginst5542 (P1_U4814, P1_U2404, P1_U4774);
  nand ginst5543 (P1_U4815, P1_U2393, P1_U4791);
  nand ginst5544 (P1_U4816, P1_INSTQUEUE_REG_11__3__SCAN_IN, P1_U4786);
  nand ginst5545 (P1_U4817, P1_U2421, P1_U4775);
  nand ginst5546 (P1_U4818, P1_U2403, P1_U2491);
  nand ginst5547 (P1_U4819, P1_U2402, P1_U4774);
  nand ginst5548 (P1_U4820, P1_U2392, P1_U4791);
  nand ginst5549 (P1_U4821, P1_INSTQUEUE_REG_11__2__SCAN_IN, P1_U4786);
  nand ginst5550 (P1_U4822, P1_U2414, P1_U4775);
  nand ginst5551 (P1_U4823, P1_U2401, P1_U2491);
  nand ginst5552 (P1_U4824, P1_U2400, P1_U4774);
  nand ginst5553 (P1_U4825, P1_U2391, P1_U4791);
  nand ginst5554 (P1_U4826, P1_INSTQUEUE_REG_11__1__SCAN_IN, P1_U4786);
  nand ginst5555 (P1_U4827, P1_U2417, P1_U4775);
  nand ginst5556 (P1_U4828, P1_U2399, P1_U2491);
  nand ginst5557 (P1_U4829, P1_U2398, P1_U4774);
  nand ginst5558 (P1_U4830, P1_U2390, P1_U4791);
  nand ginst5559 (P1_U4831, P1_INSTQUEUE_REG_11__0__SCAN_IN, P1_U4786);
  not ginst5560 (P1_U4832, P1_U3347);
  not ginst5561 (P1_U4833, P1_U3346);
  nand ginst5562 (P1_U4834, P1_U2440, P1_U2443);
  not ginst5563 (P1_U4835, P1_U3348);
  not ginst5564 (P1_U4836, P1_U3238);
  nand ginst5565 (P1_U4837, P1_U4524, P1_U4529);
  nand ginst5566 (P1_U4838, P1_U2358, P1_U2494);
  nand ginst5567 (P1_U4839, P1_U3320, P1_U4838);
  nand ginst5568 (P1_U4840, P1_U4835, P1_U4839);
  nand ginst5569 (P1_U4841, P1_STATE2_REG_3__SCAN_IN, P1_U3346);
  nand ginst5570 (P1_U4842, P1_STATE2_REG_2__SCAN_IN, P1_U3238);
  nand ginst5571 (P1_U4843, P1_U3632, P1_U4840);
  nand ginst5572 (P1_U4844, P1_U2388, P1_U2494);
  nand ginst5573 (P1_U4845, P1_U3320, P1_U4844);
  nand ginst5574 (P1_U4846, P1_U3348, P1_U4845);
  nand ginst5575 (P1_U4847, P1_STATE2_REG_2__SCAN_IN, P1_U4836);
  nand ginst5576 (P1_U4848, P1_U4846, P1_U4847);
  nand ginst5577 (P1_U4849, P1_U2415, P1_U4833);
  nand ginst5578 (P1_U4850, P1_U2413, P1_U2493);
  nand ginst5579 (P1_U4851, P1_U2412, P1_U4832);
  nand ginst5580 (P1_U4852, P1_U2397, P1_U4848);
  nand ginst5581 (P1_U4853, P1_INSTQUEUE_REG_10__7__SCAN_IN, P1_U4843);
  nand ginst5582 (P1_U4854, P1_U2416, P1_U4833);
  nand ginst5583 (P1_U4855, P1_U2411, P1_U2493);
  nand ginst5584 (P1_U4856, P1_U2410, P1_U4832);
  nand ginst5585 (P1_U4857, P1_U2396, P1_U4848);
  nand ginst5586 (P1_U4858, P1_INSTQUEUE_REG_10__6__SCAN_IN, P1_U4843);
  nand ginst5587 (P1_U4859, P1_U2420, P1_U4833);
  nand ginst5588 (P1_U4860, P1_U2409, P1_U2493);
  nand ginst5589 (P1_U4861, P1_U2408, P1_U4832);
  nand ginst5590 (P1_U4862, P1_U2395, P1_U4848);
  nand ginst5591 (P1_U4863, P1_INSTQUEUE_REG_10__5__SCAN_IN, P1_U4843);
  nand ginst5592 (P1_U4864, P1_U2419, P1_U4833);
  nand ginst5593 (P1_U4865, P1_U2407, P1_U2493);
  nand ginst5594 (P1_U4866, P1_U2406, P1_U4832);
  nand ginst5595 (P1_U4867, P1_U2394, P1_U4848);
  nand ginst5596 (P1_U4868, P1_INSTQUEUE_REG_10__4__SCAN_IN, P1_U4843);
  nand ginst5597 (P1_U4869, P1_U2418, P1_U4833);
  nand ginst5598 (P1_U4870, P1_U2405, P1_U2493);
  nand ginst5599 (P1_U4871, P1_U2404, P1_U4832);
  nand ginst5600 (P1_U4872, P1_U2393, P1_U4848);
  nand ginst5601 (P1_U4873, P1_INSTQUEUE_REG_10__3__SCAN_IN, P1_U4843);
  nand ginst5602 (P1_U4874, P1_U2421, P1_U4833);
  nand ginst5603 (P1_U4875, P1_U2403, P1_U2493);
  nand ginst5604 (P1_U4876, P1_U2402, P1_U4832);
  nand ginst5605 (P1_U4877, P1_U2392, P1_U4848);
  nand ginst5606 (P1_U4878, P1_INSTQUEUE_REG_10__2__SCAN_IN, P1_U4843);
  nand ginst5607 (P1_U4879, P1_U2414, P1_U4833);
  nand ginst5608 (P1_U4880, P1_U2401, P1_U2493);
  nand ginst5609 (P1_U4881, P1_U2400, P1_U4832);
  nand ginst5610 (P1_U4882, P1_U2391, P1_U4848);
  nand ginst5611 (P1_U4883, P1_INSTQUEUE_REG_10__1__SCAN_IN, P1_U4843);
  nand ginst5612 (P1_U4884, P1_U2417, P1_U4833);
  nand ginst5613 (P1_U4885, P1_U2399, P1_U2493);
  nand ginst5614 (P1_U4886, P1_U2398, P1_U4832);
  nand ginst5615 (P1_U4887, P1_U2390, P1_U4848);
  nand ginst5616 (P1_U4888, P1_INSTQUEUE_REG_10__0__SCAN_IN, P1_U4843);
  not ginst5617 (P1_U4889, P1_U3350);
  not ginst5618 (P1_U4890, P1_U3349);
  nand ginst5619 (P1_U4891, P1_U2440, P1_U2444);
  not ginst5620 (P1_U4892, P1_U3351);
  nand ginst5621 (P1_U4893, P1_U2434, P1_U2437);
  not ginst5622 (P1_U4894, P1_U3352);
  nand ginst5623 (P1_U4895, P1_U4525, P1_U4529);
  nand ginst5624 (P1_U4896, P1_U2358, P1_U2496);
  nand ginst5625 (P1_U4897, P1_U3320, P1_U4896);
  nand ginst5626 (P1_U4898, P1_U4892, P1_U4897);
  nand ginst5627 (P1_U4899, P1_STATE2_REG_3__SCAN_IN, P1_U3349);
  nand ginst5628 (P1_U4900, P1_STATE2_REG_2__SCAN_IN, P1_U4894);
  nand ginst5629 (P1_U4901, P1_U3641, P1_U4898);
  nand ginst5630 (P1_U4902, P1_U2388, P1_U2496);
  nand ginst5631 (P1_U4903, P1_U3320, P1_U4902);
  nand ginst5632 (P1_U4904, P1_U3351, P1_U4903);
  nand ginst5633 (P1_U4905, P1_STATE2_REG_2__SCAN_IN, P1_U3352);
  nand ginst5634 (P1_U4906, P1_U4904, P1_U4905);
  nand ginst5635 (P1_U4907, P1_U2415, P1_U4890);
  nand ginst5636 (P1_U4908, P1_U2413, P1_U2495);
  nand ginst5637 (P1_U4909, P1_U2412, P1_U4889);
  nand ginst5638 (P1_U4910, P1_U2397, P1_U4906);
  nand ginst5639 (P1_U4911, P1_INSTQUEUE_REG_9__7__SCAN_IN, P1_U4901);
  nand ginst5640 (P1_U4912, P1_U2416, P1_U4890);
  nand ginst5641 (P1_U4913, P1_U2411, P1_U2495);
  nand ginst5642 (P1_U4914, P1_U2410, P1_U4889);
  nand ginst5643 (P1_U4915, P1_U2396, P1_U4906);
  nand ginst5644 (P1_U4916, P1_INSTQUEUE_REG_9__6__SCAN_IN, P1_U4901);
  nand ginst5645 (P1_U4917, P1_U2420, P1_U4890);
  nand ginst5646 (P1_U4918, P1_U2409, P1_U2495);
  nand ginst5647 (P1_U4919, P1_U2408, P1_U4889);
  nand ginst5648 (P1_U4920, P1_U2395, P1_U4906);
  nand ginst5649 (P1_U4921, P1_INSTQUEUE_REG_9__5__SCAN_IN, P1_U4901);
  nand ginst5650 (P1_U4922, P1_U2419, P1_U4890);
  nand ginst5651 (P1_U4923, P1_U2407, P1_U2495);
  nand ginst5652 (P1_U4924, P1_U2406, P1_U4889);
  nand ginst5653 (P1_U4925, P1_U2394, P1_U4906);
  nand ginst5654 (P1_U4926, P1_INSTQUEUE_REG_9__4__SCAN_IN, P1_U4901);
  nand ginst5655 (P1_U4927, P1_U2418, P1_U4890);
  nand ginst5656 (P1_U4928, P1_U2405, P1_U2495);
  nand ginst5657 (P1_U4929, P1_U2404, P1_U4889);
  nand ginst5658 (P1_U4930, P1_U2393, P1_U4906);
  nand ginst5659 (P1_U4931, P1_INSTQUEUE_REG_9__3__SCAN_IN, P1_U4901);
  nand ginst5660 (P1_U4932, P1_U2421, P1_U4890);
  nand ginst5661 (P1_U4933, P1_U2403, P1_U2495);
  nand ginst5662 (P1_U4934, P1_U2402, P1_U4889);
  nand ginst5663 (P1_U4935, P1_U2392, P1_U4906);
  nand ginst5664 (P1_U4936, P1_INSTQUEUE_REG_9__2__SCAN_IN, P1_U4901);
  nand ginst5665 (P1_U4937, P1_U2414, P1_U4890);
  nand ginst5666 (P1_U4938, P1_U2401, P1_U2495);
  nand ginst5667 (P1_U4939, P1_U2400, P1_U4889);
  nand ginst5668 (P1_U4940, P1_U2391, P1_U4906);
  nand ginst5669 (P1_U4941, P1_INSTQUEUE_REG_9__1__SCAN_IN, P1_U4901);
  nand ginst5670 (P1_U4942, P1_U2417, P1_U4890);
  nand ginst5671 (P1_U4943, P1_U2399, P1_U2495);
  nand ginst5672 (P1_U4944, P1_U2398, P1_U4889);
  nand ginst5673 (P1_U4945, P1_U2390, P1_U4906);
  nand ginst5674 (P1_U4946, P1_INSTQUEUE_REG_9__0__SCAN_IN, P1_U4901);
  not ginst5675 (P1_U4947, P1_U3354);
  not ginst5676 (P1_U4948, P1_U3353);
  nand ginst5677 (P1_U4949, P1_U2440, P1_U2445);
  not ginst5678 (P1_U4950, P1_U3355);
  not ginst5679 (P1_U4951, P1_U3239);
  nand ginst5680 (P1_U4952, P1_U2486, P1_U4529);
  nand ginst5681 (P1_U4953, P1_U2358, P1_U2498);
  nand ginst5682 (P1_U4954, P1_U3320, P1_U4953);
  nand ginst5683 (P1_U4955, P1_U4950, P1_U4954);
  nand ginst5684 (P1_U4956, P1_STATE2_REG_3__SCAN_IN, P1_U3353);
  nand ginst5685 (P1_U4957, P1_STATE2_REG_2__SCAN_IN, P1_U3239);
  nand ginst5686 (P1_U4958, P1_U3650, P1_U4955);
  nand ginst5687 (P1_U4959, P1_U2388, P1_U2498);
  nand ginst5688 (P1_U4960, P1_U3320, P1_U4959);
  nand ginst5689 (P1_U4961, P1_U3355, P1_U4960);
  nand ginst5690 (P1_U4962, P1_STATE2_REG_2__SCAN_IN, P1_U4951);
  nand ginst5691 (P1_U4963, P1_U4961, P1_U4962);
  nand ginst5692 (P1_U4964, P1_U2415, P1_U4948);
  nand ginst5693 (P1_U4965, P1_U2413, P1_U2497);
  nand ginst5694 (P1_U4966, P1_U2412, P1_U4947);
  nand ginst5695 (P1_U4967, P1_U2397, P1_U4963);
  nand ginst5696 (P1_U4968, P1_INSTQUEUE_REG_8__7__SCAN_IN, P1_U4958);
  nand ginst5697 (P1_U4969, P1_U2416, P1_U4948);
  nand ginst5698 (P1_U4970, P1_U2411, P1_U2497);
  nand ginst5699 (P1_U4971, P1_U2410, P1_U4947);
  nand ginst5700 (P1_U4972, P1_U2396, P1_U4963);
  nand ginst5701 (P1_U4973, P1_INSTQUEUE_REG_8__6__SCAN_IN, P1_U4958);
  nand ginst5702 (P1_U4974, P1_U2420, P1_U4948);
  nand ginst5703 (P1_U4975, P1_U2409, P1_U2497);
  nand ginst5704 (P1_U4976, P1_U2408, P1_U4947);
  nand ginst5705 (P1_U4977, P1_U2395, P1_U4963);
  nand ginst5706 (P1_U4978, P1_INSTQUEUE_REG_8__5__SCAN_IN, P1_U4958);
  nand ginst5707 (P1_U4979, P1_U2419, P1_U4948);
  nand ginst5708 (P1_U4980, P1_U2407, P1_U2497);
  nand ginst5709 (P1_U4981, P1_U2406, P1_U4947);
  nand ginst5710 (P1_U4982, P1_U2394, P1_U4963);
  nand ginst5711 (P1_U4983, P1_INSTQUEUE_REG_8__4__SCAN_IN, P1_U4958);
  nand ginst5712 (P1_U4984, P1_U2418, P1_U4948);
  nand ginst5713 (P1_U4985, P1_U2405, P1_U2497);
  nand ginst5714 (P1_U4986, P1_U2404, P1_U4947);
  nand ginst5715 (P1_U4987, P1_U2393, P1_U4963);
  nand ginst5716 (P1_U4988, P1_INSTQUEUE_REG_8__3__SCAN_IN, P1_U4958);
  nand ginst5717 (P1_U4989, P1_U2421, P1_U4948);
  nand ginst5718 (P1_U4990, P1_U2403, P1_U2497);
  nand ginst5719 (P1_U4991, P1_U2402, P1_U4947);
  nand ginst5720 (P1_U4992, P1_U2392, P1_U4963);
  nand ginst5721 (P1_U4993, P1_INSTQUEUE_REG_8__2__SCAN_IN, P1_U4958);
  nand ginst5722 (P1_U4994, P1_U2414, P1_U4948);
  nand ginst5723 (P1_U4995, P1_U2401, P1_U2497);
  nand ginst5724 (P1_U4996, P1_U2400, P1_U4947);
  nand ginst5725 (P1_U4997, P1_U2391, P1_U4963);
  nand ginst5726 (P1_U4998, P1_INSTQUEUE_REG_8__1__SCAN_IN, P1_U4958);
  nand ginst5727 (P1_U4999, P1_U2417, P1_U4948);
  nand ginst5728 (P1_U5000, P1_U2399, P1_U2497);
  nand ginst5729 (P1_U5001, P1_U2398, P1_U4947);
  nand ginst5730 (P1_U5002, P1_U2390, P1_U4963);
  nand ginst5731 (P1_U5003, P1_INSTQUEUE_REG_8__0__SCAN_IN, P1_U4958);
  not ginst5732 (P1_U5004, P1_U3359);
  nand ginst5733 (P1_U5005, P1_U2439, P1_U2442);
  not ginst5734 (P1_U5006, P1_U3361);
  nand ginst5735 (P1_U5007, P1_U2433, P1_U2436);
  not ginst5736 (P1_U5008, P1_U3362);
  nand ginst5737 (P1_U5009, P1_U2358, P1_U2500);
  nand ginst5738 (P1_U5010, P1_U3320, P1_U5009);
  nand ginst5739 (P1_U5011, P1_U5006, P1_U5010);
  nand ginst5740 (P1_U5012, P1_STATE2_REG_3__SCAN_IN, P1_U3356);
  nand ginst5741 (P1_U5013, P1_STATE2_REG_2__SCAN_IN, P1_U5008);
  nand ginst5742 (P1_U5014, P1_U3659, P1_U5011);
  nand ginst5743 (P1_U5015, P1_U2388, P1_U2500);
  nand ginst5744 (P1_U5016, P1_U3320, P1_U5015);
  nand ginst5745 (P1_U5017, P1_U3361, P1_U5016);
  nand ginst5746 (P1_U5018, P1_STATE2_REG_2__SCAN_IN, P1_U3362);
  nand ginst5747 (P1_U5019, P1_U5017, P1_U5018);
  nand ginst5748 (P1_U5020, P1_U2415, P1_U4537);
  nand ginst5749 (P1_U5021, P1_U2413, P1_U4238);
  nand ginst5750 (P1_U5022, P1_U2412, P1_U5004);
  nand ginst5751 (P1_U5023, P1_U2397, P1_U5019);
  nand ginst5752 (P1_U5024, P1_INSTQUEUE_REG_7__7__SCAN_IN, P1_U5014);
  nand ginst5753 (P1_U5025, P1_U2416, P1_U4537);
  nand ginst5754 (P1_U5026, P1_U2411, P1_U4238);
  nand ginst5755 (P1_U5027, P1_U2410, P1_U5004);
  nand ginst5756 (P1_U5028, P1_U2396, P1_U5019);
  nand ginst5757 (P1_U5029, P1_INSTQUEUE_REG_7__6__SCAN_IN, P1_U5014);
  nand ginst5758 (P1_U5030, P1_U2420, P1_U4537);
  nand ginst5759 (P1_U5031, P1_U2409, P1_U4238);
  nand ginst5760 (P1_U5032, P1_U2408, P1_U5004);
  nand ginst5761 (P1_U5033, P1_U2395, P1_U5019);
  nand ginst5762 (P1_U5034, P1_INSTQUEUE_REG_7__5__SCAN_IN, P1_U5014);
  nand ginst5763 (P1_U5035, P1_U2419, P1_U4537);
  nand ginst5764 (P1_U5036, P1_U2407, P1_U4238);
  nand ginst5765 (P1_U5037, P1_U2406, P1_U5004);
  nand ginst5766 (P1_U5038, P1_U2394, P1_U5019);
  nand ginst5767 (P1_U5039, P1_INSTQUEUE_REG_7__4__SCAN_IN, P1_U5014);
  nand ginst5768 (P1_U5040, P1_U2418, P1_U4537);
  nand ginst5769 (P1_U5041, P1_U2405, P1_U4238);
  nand ginst5770 (P1_U5042, P1_U2404, P1_U5004);
  nand ginst5771 (P1_U5043, P1_U2393, P1_U5019);
  nand ginst5772 (P1_U5044, P1_INSTQUEUE_REG_7__3__SCAN_IN, P1_U5014);
  nand ginst5773 (P1_U5045, P1_U2421, P1_U4537);
  nand ginst5774 (P1_U5046, P1_U2403, P1_U4238);
  nand ginst5775 (P1_U5047, P1_U2402, P1_U5004);
  nand ginst5776 (P1_U5048, P1_U2392, P1_U5019);
  nand ginst5777 (P1_U5049, P1_INSTQUEUE_REG_7__2__SCAN_IN, P1_U5014);
  nand ginst5778 (P1_U5050, P1_U2414, P1_U4537);
  nand ginst5779 (P1_U5051, P1_U2401, P1_U4238);
  nand ginst5780 (P1_U5052, P1_U2400, P1_U5004);
  nand ginst5781 (P1_U5053, P1_U2391, P1_U5019);
  nand ginst5782 (P1_U5054, P1_INSTQUEUE_REG_7__1__SCAN_IN, P1_U5014);
  nand ginst5783 (P1_U5055, P1_U2417, P1_U4537);
  nand ginst5784 (P1_U5056, P1_U2399, P1_U4238);
  nand ginst5785 (P1_U5057, P1_U2398, P1_U5004);
  nand ginst5786 (P1_U5058, P1_U2390, P1_U5019);
  nand ginst5787 (P1_U5059, P1_INSTQUEUE_REG_7__0__SCAN_IN, P1_U5014);
  not ginst5788 (P1_U5060, P1_U3364);
  not ginst5789 (P1_U5061, P1_U3363);
  nand ginst5790 (P1_U5062, P1_U2439, P1_U2443);
  not ginst5791 (P1_U5063, P1_U3365);
  not ginst5792 (P1_U5064, P1_U3240);
  nand ginst5793 (P1_U5065, P1_U2474, P1_U4524);
  nand ginst5794 (P1_U5066, P1_U2358, P1_U2502);
  nand ginst5795 (P1_U5067, P1_U3320, P1_U5066);
  nand ginst5796 (P1_U5068, P1_U5063, P1_U5067);
  nand ginst5797 (P1_U5069, P1_STATE2_REG_3__SCAN_IN, P1_U3363);
  nand ginst5798 (P1_U5070, P1_STATE2_REG_2__SCAN_IN, P1_U3240);
  nand ginst5799 (P1_U5071, P1_U3668, P1_U5068);
  nand ginst5800 (P1_U5072, P1_U2388, P1_U2502);
  nand ginst5801 (P1_U5073, P1_U3320, P1_U5072);
  nand ginst5802 (P1_U5074, P1_U3365, P1_U5073);
  nand ginst5803 (P1_U5075, P1_STATE2_REG_2__SCAN_IN, P1_U5064);
  nand ginst5804 (P1_U5076, P1_U5074, P1_U5075);
  nand ginst5805 (P1_U5077, P1_U2415, P1_U5061);
  nand ginst5806 (P1_U5078, P1_U2413, P1_U2501);
  nand ginst5807 (P1_U5079, P1_U2412, P1_U5060);
  nand ginst5808 (P1_U5080, P1_U2397, P1_U5076);
  nand ginst5809 (P1_U5081, P1_INSTQUEUE_REG_6__7__SCAN_IN, P1_U5071);
  nand ginst5810 (P1_U5082, P1_U2416, P1_U5061);
  nand ginst5811 (P1_U5083, P1_U2411, P1_U2501);
  nand ginst5812 (P1_U5084, P1_U2410, P1_U5060);
  nand ginst5813 (P1_U5085, P1_U2396, P1_U5076);
  nand ginst5814 (P1_U5086, P1_INSTQUEUE_REG_6__6__SCAN_IN, P1_U5071);
  nand ginst5815 (P1_U5087, P1_U2420, P1_U5061);
  nand ginst5816 (P1_U5088, P1_U2409, P1_U2501);
  nand ginst5817 (P1_U5089, P1_U2408, P1_U5060);
  nand ginst5818 (P1_U5090, P1_U2395, P1_U5076);
  nand ginst5819 (P1_U5091, P1_INSTQUEUE_REG_6__5__SCAN_IN, P1_U5071);
  nand ginst5820 (P1_U5092, P1_U2419, P1_U5061);
  nand ginst5821 (P1_U5093, P1_U2407, P1_U2501);
  nand ginst5822 (P1_U5094, P1_U2406, P1_U5060);
  nand ginst5823 (P1_U5095, P1_U2394, P1_U5076);
  nand ginst5824 (P1_U5096, P1_INSTQUEUE_REG_6__4__SCAN_IN, P1_U5071);
  nand ginst5825 (P1_U5097, P1_U2418, P1_U5061);
  nand ginst5826 (P1_U5098, P1_U2405, P1_U2501);
  nand ginst5827 (P1_U5099, P1_U2404, P1_U5060);
  nand ginst5828 (P1_U5100, P1_U2393, P1_U5076);
  nand ginst5829 (P1_U5101, P1_INSTQUEUE_REG_6__3__SCAN_IN, P1_U5071);
  nand ginst5830 (P1_U5102, P1_U2421, P1_U5061);
  nand ginst5831 (P1_U5103, P1_U2403, P1_U2501);
  nand ginst5832 (P1_U5104, P1_U2402, P1_U5060);
  nand ginst5833 (P1_U5105, P1_U2392, P1_U5076);
  nand ginst5834 (P1_U5106, P1_INSTQUEUE_REG_6__2__SCAN_IN, P1_U5071);
  nand ginst5835 (P1_U5107, P1_U2414, P1_U5061);
  nand ginst5836 (P1_U5108, P1_U2401, P1_U2501);
  nand ginst5837 (P1_U5109, P1_U2400, P1_U5060);
  nand ginst5838 (P1_U5110, P1_U2391, P1_U5076);
  nand ginst5839 (P1_U5111, P1_INSTQUEUE_REG_6__1__SCAN_IN, P1_U5071);
  nand ginst5840 (P1_U5112, P1_U2417, P1_U5061);
  nand ginst5841 (P1_U5113, P1_U2399, P1_U2501);
  nand ginst5842 (P1_U5114, P1_U2398, P1_U5060);
  nand ginst5843 (P1_U5115, P1_U2390, P1_U5076);
  nand ginst5844 (P1_U5116, P1_INSTQUEUE_REG_6__0__SCAN_IN, P1_U5071);
  not ginst5845 (P1_U5117, P1_U3367);
  not ginst5846 (P1_U5118, P1_U3366);
  nand ginst5847 (P1_U5119, P1_U2439, P1_U2444);
  not ginst5848 (P1_U5120, P1_U3368);
  nand ginst5849 (P1_U5121, P1_U2433, P1_U2437);
  not ginst5850 (P1_U5122, P1_U3369);
  nand ginst5851 (P1_U5123, P1_U2474, P1_U4525);
  nand ginst5852 (P1_U5124, P1_U2358, P1_U2504);
  nand ginst5853 (P1_U5125, P1_U3320, P1_U5124);
  nand ginst5854 (P1_U5126, P1_U5120, P1_U5125);
  nand ginst5855 (P1_U5127, P1_STATE2_REG_3__SCAN_IN, P1_U3366);
  nand ginst5856 (P1_U5128, P1_STATE2_REG_2__SCAN_IN, P1_U5122);
  nand ginst5857 (P1_U5129, P1_U3677, P1_U5126);
  nand ginst5858 (P1_U5130, P1_U2388, P1_U2504);
  nand ginst5859 (P1_U5131, P1_U3320, P1_U5130);
  nand ginst5860 (P1_U5132, P1_U3368, P1_U5131);
  nand ginst5861 (P1_U5133, P1_STATE2_REG_2__SCAN_IN, P1_U3369);
  nand ginst5862 (P1_U5134, P1_U5132, P1_U5133);
  nand ginst5863 (P1_U5135, P1_U2415, P1_U5118);
  nand ginst5864 (P1_U5136, P1_U2413, P1_U2503);
  nand ginst5865 (P1_U5137, P1_U2412, P1_U5117);
  nand ginst5866 (P1_U5138, P1_U2397, P1_U5134);
  nand ginst5867 (P1_U5139, P1_INSTQUEUE_REG_5__7__SCAN_IN, P1_U5129);
  nand ginst5868 (P1_U5140, P1_U2416, P1_U5118);
  nand ginst5869 (P1_U5141, P1_U2411, P1_U2503);
  nand ginst5870 (P1_U5142, P1_U2410, P1_U5117);
  nand ginst5871 (P1_U5143, P1_U2396, P1_U5134);
  nand ginst5872 (P1_U5144, P1_INSTQUEUE_REG_5__6__SCAN_IN, P1_U5129);
  nand ginst5873 (P1_U5145, P1_U2420, P1_U5118);
  nand ginst5874 (P1_U5146, P1_U2409, P1_U2503);
  nand ginst5875 (P1_U5147, P1_U2408, P1_U5117);
  nand ginst5876 (P1_U5148, P1_U2395, P1_U5134);
  nand ginst5877 (P1_U5149, P1_INSTQUEUE_REG_5__5__SCAN_IN, P1_U5129);
  nand ginst5878 (P1_U5150, P1_U2419, P1_U5118);
  nand ginst5879 (P1_U5151, P1_U2407, P1_U2503);
  nand ginst5880 (P1_U5152, P1_U2406, P1_U5117);
  nand ginst5881 (P1_U5153, P1_U2394, P1_U5134);
  nand ginst5882 (P1_U5154, P1_INSTQUEUE_REG_5__4__SCAN_IN, P1_U5129);
  nand ginst5883 (P1_U5155, P1_U2418, P1_U5118);
  nand ginst5884 (P1_U5156, P1_U2405, P1_U2503);
  nand ginst5885 (P1_U5157, P1_U2404, P1_U5117);
  nand ginst5886 (P1_U5158, P1_U2393, P1_U5134);
  nand ginst5887 (P1_U5159, P1_INSTQUEUE_REG_5__3__SCAN_IN, P1_U5129);
  nand ginst5888 (P1_U5160, P1_U2421, P1_U5118);
  nand ginst5889 (P1_U5161, P1_U2403, P1_U2503);
  nand ginst5890 (P1_U5162, P1_U2402, P1_U5117);
  nand ginst5891 (P1_U5163, P1_U2392, P1_U5134);
  nand ginst5892 (P1_U5164, P1_INSTQUEUE_REG_5__2__SCAN_IN, P1_U5129);
  nand ginst5893 (P1_U5165, P1_U2414, P1_U5118);
  nand ginst5894 (P1_U5166, P1_U2401, P1_U2503);
  nand ginst5895 (P1_U5167, P1_U2400, P1_U5117);
  nand ginst5896 (P1_U5168, P1_U2391, P1_U5134);
  nand ginst5897 (P1_U5169, P1_INSTQUEUE_REG_5__1__SCAN_IN, P1_U5129);
  nand ginst5898 (P1_U5170, P1_U2417, P1_U5118);
  nand ginst5899 (P1_U5171, P1_U2399, P1_U2503);
  nand ginst5900 (P1_U5172, P1_U2398, P1_U5117);
  nand ginst5901 (P1_U5173, P1_U2390, P1_U5134);
  nand ginst5902 (P1_U5174, P1_INSTQUEUE_REG_5__0__SCAN_IN, P1_U5129);
  not ginst5903 (P1_U5175, P1_U3371);
  not ginst5904 (P1_U5176, P1_U3370);
  nand ginst5905 (P1_U5177, P1_U2439, P1_U2445);
  not ginst5906 (P1_U5178, P1_U3372);
  not ginst5907 (P1_U5179, P1_U3241);
  nand ginst5908 (P1_U5180, P1_U2474, P1_U2486);
  nand ginst5909 (P1_U5181, P1_U2358, P1_U2506);
  nand ginst5910 (P1_U5182, P1_U3320, P1_U5181);
  nand ginst5911 (P1_U5183, P1_U5178, P1_U5182);
  nand ginst5912 (P1_U5184, P1_STATE2_REG_3__SCAN_IN, P1_U3370);
  nand ginst5913 (P1_U5185, P1_STATE2_REG_2__SCAN_IN, P1_U3241);
  nand ginst5914 (P1_U5186, P1_U3686, P1_U5183);
  nand ginst5915 (P1_U5187, P1_U2388, P1_U2506);
  nand ginst5916 (P1_U5188, P1_U3320, P1_U5187);
  nand ginst5917 (P1_U5189, P1_U3372, P1_U5188);
  nand ginst5918 (P1_U5190, P1_STATE2_REG_2__SCAN_IN, P1_U5179);
  nand ginst5919 (P1_U5191, P1_U5189, P1_U5190);
  nand ginst5920 (P1_U5192, P1_U2415, P1_U5176);
  nand ginst5921 (P1_U5193, P1_U2413, P1_U2505);
  nand ginst5922 (P1_U5194, P1_U2412, P1_U5175);
  nand ginst5923 (P1_U5195, P1_U2397, P1_U5191);
  nand ginst5924 (P1_U5196, P1_INSTQUEUE_REG_4__7__SCAN_IN, P1_U5186);
  nand ginst5925 (P1_U5197, P1_U2416, P1_U5176);
  nand ginst5926 (P1_U5198, P1_U2411, P1_U2505);
  nand ginst5927 (P1_U5199, P1_U2410, P1_U5175);
  nand ginst5928 (P1_U5200, P1_U2396, P1_U5191);
  nand ginst5929 (P1_U5201, P1_INSTQUEUE_REG_4__6__SCAN_IN, P1_U5186);
  nand ginst5930 (P1_U5202, P1_U2420, P1_U5176);
  nand ginst5931 (P1_U5203, P1_U2409, P1_U2505);
  nand ginst5932 (P1_U5204, P1_U2408, P1_U5175);
  nand ginst5933 (P1_U5205, P1_U2395, P1_U5191);
  nand ginst5934 (P1_U5206, P1_INSTQUEUE_REG_4__5__SCAN_IN, P1_U5186);
  nand ginst5935 (P1_U5207, P1_U2419, P1_U5176);
  nand ginst5936 (P1_U5208, P1_U2407, P1_U2505);
  nand ginst5937 (P1_U5209, P1_U2406, P1_U5175);
  nand ginst5938 (P1_U5210, P1_U2394, P1_U5191);
  nand ginst5939 (P1_U5211, P1_INSTQUEUE_REG_4__4__SCAN_IN, P1_U5186);
  nand ginst5940 (P1_U5212, P1_U2418, P1_U5176);
  nand ginst5941 (P1_U5213, P1_U2405, P1_U2505);
  nand ginst5942 (P1_U5214, P1_U2404, P1_U5175);
  nand ginst5943 (P1_U5215, P1_U2393, P1_U5191);
  nand ginst5944 (P1_U5216, P1_INSTQUEUE_REG_4__3__SCAN_IN, P1_U5186);
  nand ginst5945 (P1_U5217, P1_U2421, P1_U5176);
  nand ginst5946 (P1_U5218, P1_U2403, P1_U2505);
  nand ginst5947 (P1_U5219, P1_U2402, P1_U5175);
  nand ginst5948 (P1_U5220, P1_U2392, P1_U5191);
  nand ginst5949 (P1_U5221, P1_INSTQUEUE_REG_4__2__SCAN_IN, P1_U5186);
  nand ginst5950 (P1_U5222, P1_U2414, P1_U5176);
  nand ginst5951 (P1_U5223, P1_U2401, P1_U2505);
  nand ginst5952 (P1_U5224, P1_U2400, P1_U5175);
  nand ginst5953 (P1_U5225, P1_U2391, P1_U5191);
  nand ginst5954 (P1_U5226, P1_INSTQUEUE_REG_4__1__SCAN_IN, P1_U5186);
  nand ginst5955 (P1_U5227, P1_U2417, P1_U5176);
  nand ginst5956 (P1_U5228, P1_U2399, P1_U2505);
  nand ginst5957 (P1_U5229, P1_U2398, P1_U5175);
  nand ginst5958 (P1_U5230, P1_U2390, P1_U5191);
  nand ginst5959 (P1_U5231, P1_INSTQUEUE_REG_4__0__SCAN_IN, P1_U5186);
  not ginst5960 (P1_U5232, P1_U3374);
  not ginst5961 (P1_U5233, P1_U3373);
  nand ginst5962 (P1_U5234, P1_U2441, P1_U2442);
  not ginst5963 (P1_U5235, P1_U3375);
  nand ginst5964 (P1_U5236, P1_U2435, P1_U2436);
  not ginst5965 (P1_U5237, P1_U3376);
  nand ginst5966 (P1_U5238, P1_U2508, P1_U4528);
  nand ginst5967 (P1_U5239, P1_U2358, P1_U2511);
  nand ginst5968 (P1_U5240, P1_U3320, P1_U5239);
  nand ginst5969 (P1_U5241, P1_U5235, P1_U5240);
  nand ginst5970 (P1_U5242, P1_STATE2_REG_3__SCAN_IN, P1_U3373);
  nand ginst5971 (P1_U5243, P1_STATE2_REG_2__SCAN_IN, P1_U5237);
  nand ginst5972 (P1_U5244, P1_U3695, P1_U5241);
  nand ginst5973 (P1_U5245, P1_U2388, P1_U2511);
  nand ginst5974 (P1_U5246, P1_U3320, P1_U5245);
  nand ginst5975 (P1_U5247, P1_U3375, P1_U5246);
  nand ginst5976 (P1_U5248, P1_STATE2_REG_2__SCAN_IN, P1_U3376);
  nand ginst5977 (P1_U5249, P1_U5247, P1_U5248);
  nand ginst5978 (P1_U5250, P1_U2415, P1_U5233);
  nand ginst5979 (P1_U5251, P1_U2413, P1_U2509);
  nand ginst5980 (P1_U5252, P1_U2412, P1_U5232);
  nand ginst5981 (P1_U5253, P1_U2397, P1_U5249);
  nand ginst5982 (P1_U5254, P1_INSTQUEUE_REG_3__7__SCAN_IN, P1_U5244);
  nand ginst5983 (P1_U5255, P1_U2416, P1_U5233);
  nand ginst5984 (P1_U5256, P1_U2411, P1_U2509);
  nand ginst5985 (P1_U5257, P1_U2410, P1_U5232);
  nand ginst5986 (P1_U5258, P1_U2396, P1_U5249);
  nand ginst5987 (P1_U5259, P1_INSTQUEUE_REG_3__6__SCAN_IN, P1_U5244);
  nand ginst5988 (P1_U5260, P1_U2420, P1_U5233);
  nand ginst5989 (P1_U5261, P1_U2409, P1_U2509);
  nand ginst5990 (P1_U5262, P1_U2408, P1_U5232);
  nand ginst5991 (P1_U5263, P1_U2395, P1_U5249);
  nand ginst5992 (P1_U5264, P1_INSTQUEUE_REG_3__5__SCAN_IN, P1_U5244);
  nand ginst5993 (P1_U5265, P1_U2419, P1_U5233);
  nand ginst5994 (P1_U5266, P1_U2407, P1_U2509);
  nand ginst5995 (P1_U5267, P1_U2406, P1_U5232);
  nand ginst5996 (P1_U5268, P1_U2394, P1_U5249);
  nand ginst5997 (P1_U5269, P1_INSTQUEUE_REG_3__4__SCAN_IN, P1_U5244);
  nand ginst5998 (P1_U5270, P1_U2418, P1_U5233);
  nand ginst5999 (P1_U5271, P1_U2405, P1_U2509);
  nand ginst6000 (P1_U5272, P1_U2404, P1_U5232);
  nand ginst6001 (P1_U5273, P1_U2393, P1_U5249);
  nand ginst6002 (P1_U5274, P1_INSTQUEUE_REG_3__3__SCAN_IN, P1_U5244);
  nand ginst6003 (P1_U5275, P1_U2421, P1_U5233);
  nand ginst6004 (P1_U5276, P1_U2403, P1_U2509);
  nand ginst6005 (P1_U5277, P1_U2402, P1_U5232);
  nand ginst6006 (P1_U5278, P1_U2392, P1_U5249);
  nand ginst6007 (P1_U5279, P1_INSTQUEUE_REG_3__2__SCAN_IN, P1_U5244);
  nand ginst6008 (P1_U5280, P1_U2414, P1_U5233);
  nand ginst6009 (P1_U5281, P1_U2401, P1_U2509);
  nand ginst6010 (P1_U5282, P1_U2400, P1_U5232);
  nand ginst6011 (P1_U5283, P1_U2391, P1_U5249);
  nand ginst6012 (P1_U5284, P1_INSTQUEUE_REG_3__1__SCAN_IN, P1_U5244);
  nand ginst6013 (P1_U5285, P1_U2417, P1_U5233);
  nand ginst6014 (P1_U5286, P1_U2399, P1_U2509);
  nand ginst6015 (P1_U5287, P1_U2398, P1_U5232);
  nand ginst6016 (P1_U5288, P1_U2390, P1_U5249);
  nand ginst6017 (P1_U5289, P1_INSTQUEUE_REG_3__0__SCAN_IN, P1_U5244);
  not ginst6018 (P1_U5290, P1_U3378);
  not ginst6019 (P1_U5291, P1_U3377);
  nand ginst6020 (P1_U5292, P1_U2441, P1_U2443);
  not ginst6021 (P1_U5293, P1_U3379);
  not ginst6022 (P1_U5294, P1_U3242);
  nand ginst6023 (P1_U5295, P1_U2508, P1_U4524);
  nand ginst6024 (P1_U5296, P1_U2358, P1_U2513);
  nand ginst6025 (P1_U5297, P1_U3320, P1_U5296);
  nand ginst6026 (P1_U5298, P1_U5293, P1_U5297);
  nand ginst6027 (P1_U5299, P1_STATE2_REG_3__SCAN_IN, P1_U3377);
  nand ginst6028 (P1_U5300, P1_STATE2_REG_2__SCAN_IN, P1_U3242);
  nand ginst6029 (P1_U5301, P1_U3704, P1_U5298);
  nand ginst6030 (P1_U5302, P1_U2388, P1_U2513);
  nand ginst6031 (P1_U5303, P1_U3320, P1_U5302);
  nand ginst6032 (P1_U5304, P1_U3379, P1_U5303);
  nand ginst6033 (P1_U5305, P1_STATE2_REG_2__SCAN_IN, P1_U5294);
  nand ginst6034 (P1_U5306, P1_U5304, P1_U5305);
  nand ginst6035 (P1_U5307, P1_U2415, P1_U5291);
  nand ginst6036 (P1_U5308, P1_U2413, P1_U2512);
  nand ginst6037 (P1_U5309, P1_U2412, P1_U5290);
  nand ginst6038 (P1_U5310, P1_U2397, P1_U5306);
  nand ginst6039 (P1_U5311, P1_INSTQUEUE_REG_2__7__SCAN_IN, P1_U5301);
  nand ginst6040 (P1_U5312, P1_U2416, P1_U5291);
  nand ginst6041 (P1_U5313, P1_U2411, P1_U2512);
  nand ginst6042 (P1_U5314, P1_U2410, P1_U5290);
  nand ginst6043 (P1_U5315, P1_U2396, P1_U5306);
  nand ginst6044 (P1_U5316, P1_INSTQUEUE_REG_2__6__SCAN_IN, P1_U5301);
  nand ginst6045 (P1_U5317, P1_U2420, P1_U5291);
  nand ginst6046 (P1_U5318, P1_U2409, P1_U2512);
  nand ginst6047 (P1_U5319, P1_U2408, P1_U5290);
  nand ginst6048 (P1_U5320, P1_U2395, P1_U5306);
  nand ginst6049 (P1_U5321, P1_INSTQUEUE_REG_2__5__SCAN_IN, P1_U5301);
  nand ginst6050 (P1_U5322, P1_U2419, P1_U5291);
  nand ginst6051 (P1_U5323, P1_U2407, P1_U2512);
  nand ginst6052 (P1_U5324, P1_U2406, P1_U5290);
  nand ginst6053 (P1_U5325, P1_U2394, P1_U5306);
  nand ginst6054 (P1_U5326, P1_INSTQUEUE_REG_2__4__SCAN_IN, P1_U5301);
  nand ginst6055 (P1_U5327, P1_U2418, P1_U5291);
  nand ginst6056 (P1_U5328, P1_U2405, P1_U2512);
  nand ginst6057 (P1_U5329, P1_U2404, P1_U5290);
  nand ginst6058 (P1_U5330, P1_U2393, P1_U5306);
  nand ginst6059 (P1_U5331, P1_INSTQUEUE_REG_2__3__SCAN_IN, P1_U5301);
  nand ginst6060 (P1_U5332, P1_U2421, P1_U5291);
  nand ginst6061 (P1_U5333, P1_U2403, P1_U2512);
  nand ginst6062 (P1_U5334, P1_U2402, P1_U5290);
  nand ginst6063 (P1_U5335, P1_U2392, P1_U5306);
  nand ginst6064 (P1_U5336, P1_INSTQUEUE_REG_2__2__SCAN_IN, P1_U5301);
  nand ginst6065 (P1_U5337, P1_U2414, P1_U5291);
  nand ginst6066 (P1_U5338, P1_U2401, P1_U2512);
  nand ginst6067 (P1_U5339, P1_U2400, P1_U5290);
  nand ginst6068 (P1_U5340, P1_U2391, P1_U5306);
  nand ginst6069 (P1_U5341, P1_INSTQUEUE_REG_2__1__SCAN_IN, P1_U5301);
  nand ginst6070 (P1_U5342, P1_U2417, P1_U5291);
  nand ginst6071 (P1_U5343, P1_U2399, P1_U2512);
  nand ginst6072 (P1_U5344, P1_U2398, P1_U5290);
  nand ginst6073 (P1_U5345, P1_U2390, P1_U5306);
  nand ginst6074 (P1_U5346, P1_INSTQUEUE_REG_2__0__SCAN_IN, P1_U5301);
  not ginst6075 (P1_U5347, P1_U3381);
  not ginst6076 (P1_U5348, P1_U3380);
  nand ginst6077 (P1_U5349, P1_U2441, P1_U2444);
  not ginst6078 (P1_U5350, P1_U3382);
  nand ginst6079 (P1_U5351, P1_U2435, P1_U2437);
  not ginst6080 (P1_U5352, P1_U3383);
  nand ginst6081 (P1_U5353, P1_U2508, P1_U4525);
  nand ginst6082 (P1_U5354, P1_U2358, P1_U2515);
  nand ginst6083 (P1_U5355, P1_U3320, P1_U5354);
  nand ginst6084 (P1_U5356, P1_U5350, P1_U5355);
  nand ginst6085 (P1_U5357, P1_STATE2_REG_3__SCAN_IN, P1_U3380);
  nand ginst6086 (P1_U5358, P1_STATE2_REG_2__SCAN_IN, P1_U5352);
  nand ginst6087 (P1_U5359, P1_U3713, P1_U5356);
  nand ginst6088 (P1_U5360, P1_U2388, P1_U2515);
  nand ginst6089 (P1_U5361, P1_U3320, P1_U5360);
  nand ginst6090 (P1_U5362, P1_U3382, P1_U5361);
  nand ginst6091 (P1_U5363, P1_STATE2_REG_2__SCAN_IN, P1_U3383);
  nand ginst6092 (P1_U5364, P1_U5362, P1_U5363);
  nand ginst6093 (P1_U5365, P1_U2415, P1_U5348);
  nand ginst6094 (P1_U5366, P1_U2413, P1_U2514);
  nand ginst6095 (P1_U5367, P1_U2412, P1_U5347);
  nand ginst6096 (P1_U5368, P1_U2397, P1_U5364);
  nand ginst6097 (P1_U5369, P1_INSTQUEUE_REG_1__7__SCAN_IN, P1_U5359);
  nand ginst6098 (P1_U5370, P1_U2416, P1_U5348);
  nand ginst6099 (P1_U5371, P1_U2411, P1_U2514);
  nand ginst6100 (P1_U5372, P1_U2410, P1_U5347);
  nand ginst6101 (P1_U5373, P1_U2396, P1_U5364);
  nand ginst6102 (P1_U5374, P1_INSTQUEUE_REG_1__6__SCAN_IN, P1_U5359);
  nand ginst6103 (P1_U5375, P1_U2420, P1_U5348);
  nand ginst6104 (P1_U5376, P1_U2409, P1_U2514);
  nand ginst6105 (P1_U5377, P1_U2408, P1_U5347);
  nand ginst6106 (P1_U5378, P1_U2395, P1_U5364);
  nand ginst6107 (P1_U5379, P1_INSTQUEUE_REG_1__5__SCAN_IN, P1_U5359);
  nand ginst6108 (P1_U5380, P1_U2419, P1_U5348);
  nand ginst6109 (P1_U5381, P1_U2407, P1_U2514);
  nand ginst6110 (P1_U5382, P1_U2406, P1_U5347);
  nand ginst6111 (P1_U5383, P1_U2394, P1_U5364);
  nand ginst6112 (P1_U5384, P1_INSTQUEUE_REG_1__4__SCAN_IN, P1_U5359);
  nand ginst6113 (P1_U5385, P1_U2418, P1_U5348);
  nand ginst6114 (P1_U5386, P1_U2405, P1_U2514);
  nand ginst6115 (P1_U5387, P1_U2404, P1_U5347);
  nand ginst6116 (P1_U5388, P1_U2393, P1_U5364);
  nand ginst6117 (P1_U5389, P1_INSTQUEUE_REG_1__3__SCAN_IN, P1_U5359);
  nand ginst6118 (P1_U5390, P1_U2421, P1_U5348);
  nand ginst6119 (P1_U5391, P1_U2403, P1_U2514);
  nand ginst6120 (P1_U5392, P1_U2402, P1_U5347);
  nand ginst6121 (P1_U5393, P1_U2392, P1_U5364);
  nand ginst6122 (P1_U5394, P1_INSTQUEUE_REG_1__2__SCAN_IN, P1_U5359);
  nand ginst6123 (P1_U5395, P1_U2414, P1_U5348);
  nand ginst6124 (P1_U5396, P1_U2401, P1_U2514);
  nand ginst6125 (P1_U5397, P1_U2400, P1_U5347);
  nand ginst6126 (P1_U5398, P1_U2391, P1_U5364);
  nand ginst6127 (P1_U5399, P1_INSTQUEUE_REG_1__1__SCAN_IN, P1_U5359);
  nand ginst6128 (P1_U5400, P1_U2417, P1_U5348);
  nand ginst6129 (P1_U5401, P1_U2399, P1_U2514);
  nand ginst6130 (P1_U5402, P1_U2398, P1_U5347);
  nand ginst6131 (P1_U5403, P1_U2390, P1_U5364);
  nand ginst6132 (P1_U5404, P1_INSTQUEUE_REG_1__0__SCAN_IN, P1_U5359);
  not ginst6133 (P1_U5405, P1_U3385);
  not ginst6134 (P1_U5406, P1_U3384);
  nand ginst6135 (P1_U5407, P1_U2441, P1_U2445);
  not ginst6136 (P1_U5408, P1_U3386);
  not ginst6137 (P1_U5409, P1_U3243);
  nand ginst6138 (P1_U5410, P1_U2486, P1_U2508);
  nand ginst6139 (P1_U5411, P1_U2358, P1_U2517);
  nand ginst6140 (P1_U5412, P1_U3320, P1_U5411);
  nand ginst6141 (P1_U5413, P1_U5408, P1_U5412);
  nand ginst6142 (P1_U5414, P1_STATE2_REG_3__SCAN_IN, P1_U3384);
  nand ginst6143 (P1_U5415, P1_STATE2_REG_2__SCAN_IN, P1_U3243);
  nand ginst6144 (P1_U5416, P1_U3722, P1_U5413);
  nand ginst6145 (P1_U5417, P1_U2388, P1_U2517);
  nand ginst6146 (P1_U5418, P1_U3320, P1_U5417);
  nand ginst6147 (P1_U5419, P1_U3386, P1_U5418);
  nand ginst6148 (P1_U5420, P1_STATE2_REG_2__SCAN_IN, P1_U5409);
  nand ginst6149 (P1_U5421, P1_U5419, P1_U5420);
  nand ginst6150 (P1_U5422, P1_U2415, P1_U5406);
  nand ginst6151 (P1_U5423, P1_U2413, P1_U2516);
  nand ginst6152 (P1_U5424, P1_U2412, P1_U5405);
  nand ginst6153 (P1_U5425, P1_U2397, P1_U5421);
  nand ginst6154 (P1_U5426, P1_INSTQUEUE_REG_0__7__SCAN_IN, P1_U5416);
  nand ginst6155 (P1_U5427, P1_U2416, P1_U5406);
  nand ginst6156 (P1_U5428, P1_U2411, P1_U2516);
  nand ginst6157 (P1_U5429, P1_U2410, P1_U5405);
  nand ginst6158 (P1_U5430, P1_U2396, P1_U5421);
  nand ginst6159 (P1_U5431, P1_INSTQUEUE_REG_0__6__SCAN_IN, P1_U5416);
  nand ginst6160 (P1_U5432, P1_U2420, P1_U5406);
  nand ginst6161 (P1_U5433, P1_U2409, P1_U2516);
  nand ginst6162 (P1_U5434, P1_U2408, P1_U5405);
  nand ginst6163 (P1_U5435, P1_U2395, P1_U5421);
  nand ginst6164 (P1_U5436, P1_INSTQUEUE_REG_0__5__SCAN_IN, P1_U5416);
  nand ginst6165 (P1_U5437, P1_U2419, P1_U5406);
  nand ginst6166 (P1_U5438, P1_U2407, P1_U2516);
  nand ginst6167 (P1_U5439, P1_U2406, P1_U5405);
  nand ginst6168 (P1_U5440, P1_U2394, P1_U5421);
  nand ginst6169 (P1_U5441, P1_U2418, P1_U5406);
  nand ginst6170 (P1_U5442, P1_U2405, P1_U2516);
  nand ginst6171 (P1_U5443, P1_U2404, P1_U5405);
  nand ginst6172 (P1_U5444, P1_U2393, P1_U5421);
  nand ginst6173 (P1_U5445, P1_INSTQUEUE_REG_0__3__SCAN_IN, P1_U5416);
  nand ginst6174 (P1_U5446, P1_U2421, P1_U5406);
  nand ginst6175 (P1_U5447, P1_U2403, P1_U2516);
  nand ginst6176 (P1_U5448, P1_U2402, P1_U5405);
  nand ginst6177 (P1_U5449, P1_U2392, P1_U5421);
  nand ginst6178 (P1_U5450, P1_INSTQUEUE_REG_0__2__SCAN_IN, P1_U5416);
  nand ginst6179 (P1_U5451, P1_U2414, P1_U5406);
  nand ginst6180 (P1_U5452, P1_U2401, P1_U2516);
  nand ginst6181 (P1_U5453, P1_U2400, P1_U5405);
  nand ginst6182 (P1_U5454, P1_U2391, P1_U5421);
  nand ginst6183 (P1_U5455, P1_INSTQUEUE_REG_0__1__SCAN_IN, P1_U5416);
  nand ginst6184 (P1_U5456, P1_U2417, P1_U5406);
  nand ginst6185 (P1_U5457, P1_U2399, P1_U2516);
  nand ginst6186 (P1_U5458, P1_U2398, P1_U5405);
  nand ginst6187 (P1_U5459, P1_U2390, P1_U5421);
  nand ginst6188 (P1_U5460, P1_INSTQUEUE_REG_0__0__SCAN_IN, P1_U5416);
  not ginst6189 (P1_U5461, P1_U3423);
  nand ginst6190 (P1_U5462, P1_U3391, P1_U3394, P1_U4503);
  nand ginst6191 (P1_U5463, P1_U4173, P1_U4400, P1_U4460);
  not ginst6192 (P1_U5464, P1_U3244);
  nand ginst6193 (P1_U5465, P1_U3289, P1_U4494);
  nand ginst6194 (P1_U5466, P1_U3283, P1_U5464, P1_U5465);
  nand ginst6195 (P1_U5467, P1_U2452, P1_U3732);
  nand ginst6196 (P1_U5468, P1_U4208, P1_U5462);
  nand ginst6197 (P1_U5469, P1_U3733, P1_U7609);
  nand ginst6198 (P1_U5470, P1_GTE_485_U6, P1_U3257, P1_U4215);
  nand ginst6199 (P1_U5471, P1_U2449, P1_U7494);
  nand ginst6200 (P1_U5472, P1_U4257, P1_U4503);
  not ginst6201 (P1_U5473, P1_U4182);
  nand ginst6202 (P1_U5474, P1_U2368, P1_U4182);
  nand ginst6203 (P1_U5475, P1_STATE2_REG_3__SCAN_IN, P1_U3294);
  not ginst6204 (P1_U5476, P1_U4172);
  nand ginst6205 (P1_U5477, P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN);
  nand ginst6206 (P1_U5478, P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P1_U5477);
  nand ginst6207 (P1_U5479, P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P1_U4381);
  not ginst6208 (P1_U5480, P1_U3442);
  nand ginst6209 (P1_U5481, P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN, P1_U3498);
  nand ginst6210 (P1_U5482, P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P1_U5481);
  not ginst6211 (P1_U5483, P1_U3438);
  nand ginst6212 (P1_U5484, P1_U3264, P1_U3275);
  nand ginst6213 (P1_U5485, P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P1_U5484);
  nand ginst6214 (P1_U5486, P1_U2469, P1_U3275);
  nand ginst6215 (P1_U5487, P1_U3290, P1_U4494);
  nand ginst6216 (P1_U5488, P1_U2605, P1_U4400);
  nand ginst6217 (P1_U5489, P1_U7494, P1_U7703, P1_U7704);
  nand ginst6218 (P1_U5490, P1_U4449, P1_U5488);
  nand ginst6219 (P1_U5491, P1_U3394, P1_U3409, P1_U4400);
  nand ginst6220 (P1_U5492, P1_U4171, P1_U5491);
  nand ginst6221 (P1_U5493, P1_U5492, P1_U7629);
  nand ginst6222 (P1_U5494, P1_U4171, P1_U4460);
  nand ginst6223 (P1_U5495, P1_U3395, P1_U5494);
  nand ginst6224 (P1_U5496, P1_U4208, P1_U5462);
  nand ginst6225 (P1_U5497, P1_U4257, P1_U4503);
  nand ginst6226 (P1_U5498, P1_U3271, P1_U5495);
  nand ginst6227 (P1_U5499, P1_U4494, P1_U7707);
  nand ginst6228 (P1_U5500, P1_U3244, P1_U4190);
  nand ginst6229 (P1_U5501, P1_U3292, P1_U4217);
  nand ginst6230 (P1_U5502, P1_U3740, P1_U5501);
  nand ginst6231 (P1_U5503, P1_R2182_U25, P1_U7509);
  nand ginst6232 (P1_U5504, P1_U3438, P1_U4218);
  nand ginst6233 (P1_U5505, P1_U3442, P1_U4214);
  nand ginst6234 (P1_U5506, P1_U3747, P1_U5503);
  nand ginst6235 (P1_U5507, P1_U3438, P1_U4252);
  nand ginst6236 (P1_U5508, P1_U2427, P1_U5506);
  nand ginst6237 (P1_U5509, P1_U5507, P1_U5508);
  nand ginst6238 (P1_U5510, P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN, P1_U3275);
  not ginst6239 (P1_U5511, P1_U3401);
  nand ginst6240 (P1_U5512, P1_R2182_U42, P1_U7509);
  nand ginst6241 (P1_U5513, P1_U3456, P1_U4214);
  nand ginst6242 (P1_U5514, P1_U3749, P1_U5512);
  nand ginst6243 (P1_U5515, P1_U2446, P1_U3470);
  nand ginst6244 (P1_U5516, P1_U3401, P1_U4252);
  nand ginst6245 (P1_U5517, P1_U2427, P1_U5514);
  nand ginst6246 (P1_U5518, P1_U5515, P1_U5516, P1_U5517);
  not ginst6247 (P1_U5519, P1_U3402);
  nand ginst6248 (P1_U5520, P1_U2431, P1_U4249);
  nand ginst6249 (P1_U5521, P1_U3292, P1_U5520);
  nand ginst6250 (P1_U5522, P1_U5519, P1_U5521);
  nand ginst6251 (P1_U5523, P1_R2182_U33, P1_U7509);
  nand ginst6252 (P1_U5524, P1_U3265, P1_U4214);
  nand ginst6253 (P1_U5525, P1_U3750, P1_U5523);
  nand ginst6254 (P1_U5526, P1_U2446, P1_U7712);
  nand ginst6255 (P1_U5527, P1_U4252, P1_U5519);
  nand ginst6256 (P1_U5528, P1_U2427, P1_U5525);
  nand ginst6257 (P1_U5529, P1_U5526, P1_U5527, P1_U5528);
  nand ginst6258 (P1_U5530, P1_R2182_U34, P1_U7509);
  nand ginst6259 (P1_U5531, P1_U4175, P1_U5530);
  nand ginst6260 (P1_U5532, P1_U3266, P1_U4252);
  nand ginst6261 (P1_U5533, P1_U2427, P1_U5531);
  nand ginst6262 (P1_U5534, P1_STATE2_REG_1__SCAN_IN, P1_U7715);
  nand ginst6263 (P1_U5535, P1_U5532, P1_U5533, P1_U5534);
  nand ginst6264 (P1_U5536, P1_STATE2_REG_0__SCAN_IN, P1_LT_589_U6, P1_U2428);
  not ginst6265 (P1_U5537, P1_U3404);
  nand ginst6266 (P1_U5538, P1_STATE2_REG_1__SCAN_IN, P1_U3296);
  nand ginst6267 (P1_U5539, P1_U3454, P1_U4527);
  nand ginst6268 (P1_U5540, P1_U3358, P1_U5539);
  nand ginst6269 (P1_U5541, P1_U3359, P1_U5540);
  nand ginst6270 (P1_U5542, P1_U2388, P1_U5541);
  nand ginst6271 (P1_U5543, P1_R2182_U25, P1_U5538);
  nand ginst6272 (P1_U5544, P1_R2144_U8, P1_U4226);
  nand ginst6273 (P1_U5545, P1_U3751, P1_U5542);
  nand ginst6274 (P1_U5546, P1_U2388, P1_U7733);
  nand ginst6275 (P1_U5547, P1_R2182_U42, P1_U5538);
  nand ginst6276 (P1_U5548, P1_R2144_U49, P1_U4226);
  nand ginst6277 (P1_U5549, P1_U3752, P1_U5546);
  nand ginst6278 (P1_U5550, P1_U3326, P1_U3333);
  nand ginst6279 (P1_U5551, P1_U2388, P1_U5550);
  nand ginst6280 (P1_U5552, P1_R2182_U33, P1_U5538);
  nand ginst6281 (P1_U5553, P1_R2144_U50, P1_U4226);
  nand ginst6282 (P1_U5554, P1_U3753, P1_U5551);
  nand ginst6283 (P1_U5555, P1_R2182_U34, P1_U5538);
  nand ginst6284 (P1_U5556, P1_R2144_U43, P1_U4209);
  nand ginst6285 (P1_U5557, P1_U4245, P1_U5555, P1_U5556);
  nand ginst6286 (P1_U5558, P1_U3272, P1_U4477);
  nand ginst6287 (P1_U5559, P1_U2431, P1_U4260);
  nand ginst6288 (P1_U5560, P1_U2518, P1_U5559, P1_U7742, P1_U7743);
  nand ginst6289 (P1_U5561, P1_U4192, P1_U4235, P1_U4503);
  nand ginst6290 (P1_U5562, P1_U2368, P1_U5560);
  nand ginst6291 (P1_U5563, P1_U3263, P1_U4203);
  not ginst6292 (P1_U5564, P1_U3414);
  nand ginst6293 (P1_U5565, P1_U4208, P1_U4262);
  nand ginst6294 (P1_U5566, P1_U2389, P1_U4256);
  nand ginst6295 (P1_U5567, P1_U4250, P1_U4266);
  nand ginst6296 (P1_U5568, P1_U4264, P1_U4494);
  nand ginst6297 (P1_U5569, P1_U2519, P1_U3758);
  nand ginst6298 (P1_U5570, P1_R2099_U86, P1_U2380);
  nand ginst6299 (P1_U5571, P1_R2027_U5, P1_U2378);
  nand ginst6300 (P1_U5572, P1_R2278_U99, P1_U2377);
  nand ginst6301 (P1_U5573, P1_ADD_405_U4, P1_U2375);
  nand ginst6302 (P1_U5574, P1_INSTADDRPOINTER_REG_0__SCAN_IN, P1_U2374);
  nand ginst6303 (P1_U5575, P1_REIP_REG_0__SCAN_IN, P1_U2370);
  nand ginst6304 (P1_U5576, P1_INSTADDRPOINTER_REG_0__SCAN_IN, P1_U5564);
  nand ginst6305 (P1_U5577, P1_R2099_U87, P1_U2380);
  nand ginst6306 (P1_U5578, P1_R2027_U71, P1_U2378);
  nand ginst6307 (P1_U5579, P1_R2278_U19, P1_U2377);
  nand ginst6308 (P1_U5580, P1_ADD_405_U85, P1_U2375);
  nand ginst6309 (P1_U5581, P1_ADD_515_U4, P1_U2374);
  nand ginst6310 (P1_U5582, P1_REIP_REG_1__SCAN_IN, P1_U2370);
  nand ginst6311 (P1_U5583, P1_INSTADDRPOINTER_REG_1__SCAN_IN, P1_U5564);
  nand ginst6312 (P1_U5584, P1_R2099_U138, P1_U2380);
  nand ginst6313 (P1_U5585, P1_R2027_U60, P1_U2378);
  nand ginst6314 (P1_U5586, P1_R2278_U107, P1_U2377);
  nand ginst6315 (P1_U5587, P1_ADD_405_U5, P1_U2375);
  nand ginst6316 (P1_U5588, P1_ADD_515_U67, P1_U2374);
  nand ginst6317 (P1_U5589, P1_REIP_REG_2__SCAN_IN, P1_U2370);
  nand ginst6318 (P1_U5590, P1_INSTADDRPOINTER_REG_2__SCAN_IN, P1_U5564);
  nand ginst6319 (P1_U5591, P1_R2099_U42, P1_U2380);
  nand ginst6320 (P1_U5592, P1_R2027_U57, P1_U2378);
  nand ginst6321 (P1_U5593, P1_R2278_U105, P1_U2377);
  nand ginst6322 (P1_U5594, P1_ADD_405_U95, P1_U2375);
  nand ginst6323 (P1_U5595, P1_ADD_515_U85, P1_U2374);
  nand ginst6324 (P1_U5596, P1_REIP_REG_3__SCAN_IN, P1_U2370);
  nand ginst6325 (P1_U5597, P1_INSTADDRPOINTER_REG_3__SCAN_IN, P1_U5564);
  nand ginst6326 (P1_U5598, P1_R2099_U41, P1_U2380);
  nand ginst6327 (P1_U5599, P1_R2027_U56, P1_U2378);
  nand ginst6328 (P1_U5600, P1_R2278_U104, P1_U2377);
  nand ginst6329 (P1_U5601, P1_ADD_405_U76, P1_U2375);
  nand ginst6330 (P1_U5602, P1_ADD_515_U76, P1_U2374);
  nand ginst6331 (P1_U5603, P1_REIP_REG_4__SCAN_IN, P1_U2370);
  nand ginst6332 (P1_U5604, P1_INSTADDRPOINTER_REG_4__SCAN_IN, P1_U5564);
  nand ginst6333 (P1_U5605, P1_R2099_U40, P1_U2380);
  nand ginst6334 (P1_U5606, P1_R2027_U55, P1_U2378);
  nand ginst6335 (P1_U5607, P1_R2278_U17, P1_U2377);
  nand ginst6336 (P1_U5608, P1_ADD_405_U79, P1_U2375);
  nand ginst6337 (P1_U5609, P1_ADD_515_U79, P1_U2374);
  nand ginst6338 (P1_U5610, P1_REIP_REG_5__SCAN_IN, P1_U2370);
  nand ginst6339 (P1_U5611, P1_INSTADDRPOINTER_REG_5__SCAN_IN, P1_U5564);
  nand ginst6340 (P1_U5612, P1_R2099_U39, P1_U2380);
  nand ginst6341 (P1_U5613, P1_R2027_U54, P1_U2378);
  nand ginst6342 (P1_U5614, P1_R2278_U103, P1_U2377);
  nand ginst6343 (P1_U5615, P1_ADD_405_U63, P1_U2375);
  nand ginst6344 (P1_U5616, P1_ADD_515_U62, P1_U2374);
  nand ginst6345 (P1_U5617, P1_REIP_REG_6__SCAN_IN, P1_U2370);
  nand ginst6346 (P1_U5618, P1_INSTADDRPOINTER_REG_6__SCAN_IN, P1_U5564);
  nand ginst6347 (P1_U5619, P1_R2099_U38, P1_U2380);
  nand ginst6348 (P1_U5620, P1_R2027_U53, P1_U2378);
  nand ginst6349 (P1_U5621, P1_R2278_U18, P1_U2377);
  nand ginst6350 (P1_U5622, P1_ADD_405_U89, P1_U2375);
  nand ginst6351 (P1_U5623, P1_ADD_515_U89, P1_U2374);
  nand ginst6352 (P1_U5624, P1_REIP_REG_7__SCAN_IN, P1_U2370);
  nand ginst6353 (P1_U5625, P1_INSTADDRPOINTER_REG_7__SCAN_IN, P1_U5564);
  nand ginst6354 (P1_U5626, P1_R2099_U37, P1_U2380);
  nand ginst6355 (P1_U5627, P1_R2027_U52, P1_U2378);
  nand ginst6356 (P1_U5628, P1_R2278_U102, P1_U2377);
  nand ginst6357 (P1_U5629, P1_ADD_405_U80, P1_U2375);
  nand ginst6358 (P1_U5630, P1_ADD_515_U80, P1_U2374);
  nand ginst6359 (P1_U5631, P1_REIP_REG_8__SCAN_IN, P1_U2370);
  nand ginst6360 (P1_U5632, P1_INSTADDRPOINTER_REG_8__SCAN_IN, P1_U5564);
  nand ginst6361 (P1_U5633, P1_R2099_U36, P1_U2380);
  nand ginst6362 (P1_U5634, P1_R2027_U51, P1_U2378);
  nand ginst6363 (P1_U5635, P1_R2278_U101, P1_U2377);
  nand ginst6364 (P1_U5636, P1_ADD_405_U70, P1_U2375);
  nand ginst6365 (P1_U5637, P1_ADD_515_U70, P1_U2374);
  nand ginst6366 (P1_U5638, P1_REIP_REG_9__SCAN_IN, P1_U2370);
  nand ginst6367 (P1_U5639, P1_INSTADDRPOINTER_REG_9__SCAN_IN, P1_U5564);
  nand ginst6368 (P1_U5640, P1_R2099_U85, P1_U2380);
  nand ginst6369 (P1_U5641, P1_R2027_U81, P1_U2378);
  nand ginst6370 (P1_U5642, P1_R2278_U126, P1_U2377);
  nand ginst6371 (P1_U5643, P1_ADD_405_U83, P1_U2375);
  nand ginst6372 (P1_U5644, P1_ADD_515_U83, P1_U2374);
  nand ginst6373 (P1_U5645, P1_REIP_REG_10__SCAN_IN, P1_U2370);
  nand ginst6374 (P1_U5646, P1_INSTADDRPOINTER_REG_10__SCAN_IN, P1_U5564);
  nand ginst6375 (P1_U5647, P1_R2099_U84, P1_U2380);
  nand ginst6376 (P1_U5648, P1_R2027_U80, P1_U2378);
  nand ginst6377 (P1_U5649, P1_R2278_U15, P1_U2377);
  nand ginst6378 (P1_U5650, P1_ADD_405_U73, P1_U2375);
  nand ginst6379 (P1_U5651, P1_ADD_515_U73, P1_U2374);
  nand ginst6380 (P1_U5652, P1_REIP_REG_11__SCAN_IN, P1_U2370);
  nand ginst6381 (P1_U5653, P1_INSTADDRPOINTER_REG_11__SCAN_IN, P1_U5564);
  nand ginst6382 (P1_U5654, P1_R2099_U83, P1_U2380);
  nand ginst6383 (P1_U5655, P1_R2027_U79, P1_U2378);
  nand ginst6384 (P1_U5656, P1_R2278_U125, P1_U2377);
  nand ginst6385 (P1_U5657, P1_ADD_405_U88, P1_U2375);
  nand ginst6386 (P1_U5658, P1_ADD_515_U88, P1_U2374);
  nand ginst6387 (P1_U5659, P1_REIP_REG_12__SCAN_IN, P1_U2370);
  nand ginst6388 (P1_U5660, P1_INSTADDRPOINTER_REG_12__SCAN_IN, P1_U5564);
  nand ginst6389 (P1_U5661, P1_R2099_U82, P1_U2380);
  nand ginst6390 (P1_U5662, P1_R2027_U78, P1_U2378);
  nand ginst6391 (P1_U5663, P1_R2278_U123, P1_U2377);
  nand ginst6392 (P1_U5664, P1_ADD_405_U69, P1_U2375);
  nand ginst6393 (P1_U5665, P1_ADD_515_U69, P1_U2374);
  nand ginst6394 (P1_U5666, P1_REIP_REG_13__SCAN_IN, P1_U2370);
  nand ginst6395 (P1_U5667, P1_INSTADDRPOINTER_REG_13__SCAN_IN, P1_U5564);
  nand ginst6396 (P1_U5668, P1_R2099_U81, P1_U2380);
  nand ginst6397 (P1_U5669, P1_R2027_U77, P1_U2378);
  nand ginst6398 (P1_U5670, P1_R2278_U122, P1_U2377);
  nand ginst6399 (P1_U5671, P1_ADD_405_U78, P1_U2375);
  nand ginst6400 (P1_U5672, P1_ADD_515_U78, P1_U2374);
  nand ginst6401 (P1_U5673, P1_REIP_REG_14__SCAN_IN, P1_U2370);
  nand ginst6402 (P1_U5674, P1_INSTADDRPOINTER_REG_14__SCAN_IN, P1_U5564);
  nand ginst6403 (P1_U5675, P1_R2099_U80, P1_U2380);
  nand ginst6404 (P1_U5676, P1_R2027_U76, P1_U2378);
  nand ginst6405 (P1_U5677, P1_R2278_U20, P1_U2377);
  nand ginst6406 (P1_U5678, P1_ADD_405_U75, P1_U2375);
  nand ginst6407 (P1_U5679, P1_ADD_515_U75, P1_U2374);
  nand ginst6408 (P1_U5680, P1_REIP_REG_15__SCAN_IN, P1_U2370);
  nand ginst6409 (P1_U5681, P1_INSTADDRPOINTER_REG_15__SCAN_IN, P1_U5564);
  nand ginst6410 (P1_U5682, P1_R2099_U79, P1_U2380);
  nand ginst6411 (P1_U5683, P1_R2027_U75, P1_U2378);
  nand ginst6412 (P1_U5684, P1_R2278_U121, P1_U2377);
  nand ginst6413 (P1_U5685, P1_ADD_405_U91, P1_U2375);
  nand ginst6414 (P1_U5686, P1_ADD_515_U91, P1_U2374);
  nand ginst6415 (P1_U5687, P1_REIP_REG_16__SCAN_IN, P1_U2370);
  nand ginst6416 (P1_U5688, P1_INSTADDRPOINTER_REG_16__SCAN_IN, P1_U5564);
  nand ginst6417 (P1_U5689, P1_R2099_U78, P1_U2380);
  nand ginst6418 (P1_U5690, P1_R2027_U74, P1_U2378);
  nand ginst6419 (P1_U5691, P1_R2278_U120, P1_U2377);
  nand ginst6420 (P1_U5692, P1_ADD_405_U67, P1_U2375);
  nand ginst6421 (P1_U5693, P1_ADD_515_U66, P1_U2374);
  nand ginst6422 (P1_U5694, P1_REIP_REG_17__SCAN_IN, P1_U2370);
  nand ginst6423 (P1_U5695, P1_INSTADDRPOINTER_REG_17__SCAN_IN, P1_U5564);
  nand ginst6424 (P1_U5696, P1_R2099_U77, P1_U2380);
  nand ginst6425 (P1_U5697, P1_R2027_U73, P1_U2378);
  nand ginst6426 (P1_U5698, P1_R2278_U119, P1_U2377);
  nand ginst6427 (P1_U5699, P1_ADD_405_U72, P1_U2375);
  nand ginst6428 (P1_U5700, P1_ADD_515_U72, P1_U2374);
  nand ginst6429 (P1_U5701, P1_REIP_REG_18__SCAN_IN, P1_U2370);
  nand ginst6430 (P1_U5702, P1_INSTADDRPOINTER_REG_18__SCAN_IN, P1_U5564);
  nand ginst6431 (P1_U5703, P1_R2099_U76, P1_U2380);
  nand ginst6432 (P1_U5704, P1_R2027_U72, P1_U2378);
  nand ginst6433 (P1_U5705, P1_R2278_U118, P1_U2377);
  nand ginst6434 (P1_U5706, P1_ADD_405_U82, P1_U2375);
  nand ginst6435 (P1_U5707, P1_ADD_515_U82, P1_U2374);
  nand ginst6436 (P1_U5708, P1_REIP_REG_19__SCAN_IN, P1_U2370);
  nand ginst6437 (P1_U5709, P1_INSTADDRPOINTER_REG_19__SCAN_IN, P1_U5564);
  nand ginst6438 (P1_U5710, P1_R2099_U75, P1_U2380);
  nand ginst6439 (P1_U5711, P1_R2027_U70, P1_U2378);
  nand ginst6440 (P1_U5712, P1_R2278_U117, P1_U2377);
  nand ginst6441 (P1_U5713, P1_ADD_405_U68, P1_U2375);
  nand ginst6442 (P1_U5714, P1_ADD_515_U68, P1_U2374);
  nand ginst6443 (P1_U5715, P1_REIP_REG_20__SCAN_IN, P1_U2370);
  nand ginst6444 (P1_U5716, P1_INSTADDRPOINTER_REG_20__SCAN_IN, P1_U5564);
  nand ginst6445 (P1_U5717, P1_R2099_U74, P1_U2380);
  nand ginst6446 (P1_U5718, P1_R2027_U69, P1_U2378);
  nand ginst6447 (P1_U5719, P1_R2278_U116, P1_U2377);
  nand ginst6448 (P1_U5720, P1_ADD_405_U87, P1_U2375);
  nand ginst6449 (P1_U5721, P1_ADD_515_U87, P1_U2374);
  nand ginst6450 (P1_U5722, P1_REIP_REG_21__SCAN_IN, P1_U2370);
  nand ginst6451 (P1_U5723, P1_INSTADDRPOINTER_REG_21__SCAN_IN, P1_U5564);
  nand ginst6452 (P1_U5724, P1_R2099_U73, P1_U2380);
  nand ginst6453 (P1_U5725, P1_R2027_U68, P1_U2378);
  nand ginst6454 (P1_U5726, P1_R2278_U115, P1_U2377);
  nand ginst6455 (P1_U5727, P1_ADD_405_U71, P1_U2375);
  nand ginst6456 (P1_U5728, P1_ADD_515_U71, P1_U2374);
  nand ginst6457 (P1_U5729, P1_REIP_REG_22__SCAN_IN, P1_U2370);
  nand ginst6458 (P1_U5730, P1_INSTADDRPOINTER_REG_22__SCAN_IN, P1_U5564);
  nand ginst6459 (P1_U5731, P1_R2099_U72, P1_U2380);
  nand ginst6460 (P1_U5732, P1_R2027_U67, P1_U2378);
  nand ginst6461 (P1_U5733, P1_R2278_U114, P1_U2377);
  nand ginst6462 (P1_U5734, P1_ADD_405_U81, P1_U2375);
  nand ginst6463 (P1_U5735, P1_ADD_515_U81, P1_U2374);
  nand ginst6464 (P1_U5736, P1_REIP_REG_23__SCAN_IN, P1_U2370);
  nand ginst6465 (P1_U5737, P1_INSTADDRPOINTER_REG_23__SCAN_IN, P1_U5564);
  nand ginst6466 (P1_U5738, P1_R2099_U71, P1_U2380);
  nand ginst6467 (P1_U5739, P1_R2027_U66, P1_U2378);
  nand ginst6468 (P1_U5740, P1_R2278_U113, P1_U2377);
  nand ginst6469 (P1_U5741, P1_ADD_405_U66, P1_U2375);
  nand ginst6470 (P1_U5742, P1_ADD_515_U65, P1_U2374);
  nand ginst6471 (P1_U5743, P1_REIP_REG_24__SCAN_IN, P1_U2370);
  nand ginst6472 (P1_U5744, P1_INSTADDRPOINTER_REG_24__SCAN_IN, P1_U5564);
  nand ginst6473 (P1_U5745, P1_R2099_U70, P1_U2380);
  nand ginst6474 (P1_U5746, P1_R2027_U65, P1_U2378);
  nand ginst6475 (P1_U5747, P1_R2278_U112, P1_U2377);
  nand ginst6476 (P1_U5748, P1_ADD_405_U90, P1_U2375);
  nand ginst6477 (P1_U5749, P1_ADD_515_U90, P1_U2374);
  nand ginst6478 (P1_U5750, P1_REIP_REG_25__SCAN_IN, P1_U2370);
  nand ginst6479 (P1_U5751, P1_INSTADDRPOINTER_REG_25__SCAN_IN, P1_U5564);
  nand ginst6480 (P1_U5752, P1_R2099_U69, P1_U2380);
  nand ginst6481 (P1_U5753, P1_R2027_U64, P1_U2378);
  nand ginst6482 (P1_U5754, P1_R2278_U111, P1_U2377);
  nand ginst6483 (P1_U5755, P1_ADD_405_U74, P1_U2375);
  nand ginst6484 (P1_U5756, P1_ADD_515_U74, P1_U2374);
  nand ginst6485 (P1_U5757, P1_REIP_REG_26__SCAN_IN, P1_U2370);
  nand ginst6486 (P1_U5758, P1_INSTADDRPOINTER_REG_26__SCAN_IN, P1_U5564);
  nand ginst6487 (P1_U5759, P1_R2099_U68, P1_U2380);
  nand ginst6488 (P1_U5760, P1_R2027_U63, P1_U2378);
  nand ginst6489 (P1_U5761, P1_R2278_U110, P1_U2377);
  nand ginst6490 (P1_U5762, P1_ADD_405_U77, P1_U2375);
  nand ginst6491 (P1_U5763, P1_ADD_515_U77, P1_U2374);
  nand ginst6492 (P1_U5764, P1_REIP_REG_27__SCAN_IN, P1_U2370);
  nand ginst6493 (P1_U5765, P1_INSTADDRPOINTER_REG_27__SCAN_IN, P1_U5564);
  nand ginst6494 (P1_U5766, P1_R2099_U67, P1_U2380);
  nand ginst6495 (P1_U5767, P1_R2027_U62, P1_U2378);
  nand ginst6496 (P1_U5768, P1_R2278_U109, P1_U2377);
  nand ginst6497 (P1_U5769, P1_ADD_405_U86, P1_U2375);
  nand ginst6498 (P1_U5770, P1_ADD_515_U86, P1_U2374);
  nand ginst6499 (P1_U5771, P1_REIP_REG_28__SCAN_IN, P1_U2370);
  nand ginst6500 (P1_U5772, P1_INSTADDRPOINTER_REG_28__SCAN_IN, P1_U5564);
  nand ginst6501 (P1_U5773, P1_R2099_U66, P1_U2380);
  nand ginst6502 (P1_U5774, P1_R2027_U61, P1_U2378);
  nand ginst6503 (P1_U5775, P1_R2278_U108, P1_U2377);
  nand ginst6504 (P1_U5776, P1_ADD_405_U65, P1_U2375);
  nand ginst6505 (P1_U5777, P1_ADD_515_U64, P1_U2374);
  nand ginst6506 (P1_U5778, P1_REIP_REG_29__SCAN_IN, P1_U2370);
  nand ginst6507 (P1_U5779, P1_INSTADDRPOINTER_REG_29__SCAN_IN, P1_U5564);
  nand ginst6508 (P1_U5780, P1_R2099_U65, P1_U2380);
  nand ginst6509 (P1_U5781, P1_R2027_U59, P1_U2378);
  nand ginst6510 (P1_U5782, P1_R2278_U106, P1_U2377);
  nand ginst6511 (P1_U5783, P1_ADD_405_U64, P1_U2375);
  nand ginst6512 (P1_U5784, P1_ADD_515_U63, P1_U2374);
  nand ginst6513 (P1_U5785, P1_REIP_REG_30__SCAN_IN, P1_U2370);
  nand ginst6514 (P1_U5786, P1_INSTADDRPOINTER_REG_30__SCAN_IN, P1_U5564);
  nand ginst6515 (P1_U5787, P1_R2099_U64, P1_U2380);
  nand ginst6516 (P1_U5788, P1_R2027_U58, P1_U2378);
  nand ginst6517 (P1_U5789, P1_R2278_U16, P1_U2377);
  nand ginst6518 (P1_U5790, P1_ADD_405_U84, P1_U2375);
  nand ginst6519 (P1_U5791, P1_ADD_515_U84, P1_U2374);
  nand ginst6520 (P1_U5792, P1_REIP_REG_31__SCAN_IN, P1_U2370);
  nand ginst6521 (P1_U5793, P1_INSTADDRPOINTER_REG_31__SCAN_IN, P1_U5564);
  nand ginst6522 (P1_U5794, P1_U3294, P1_U4209);
  not ginst6523 (P1_U5795, P1_U3416);
  nand ginst6524 (P1_U5796, P1_STATE2_REG_2__SCAN_IN, P1_U3294);
  nand ginst6525 (P1_U5797, P1_STATE2_REG_1__SCAN_IN, P1_U3308);
  nand ginst6526 (P1_U5798, P1_U5796, P1_U5797);
  nand ginst6527 (P1_U5799, P1_PHYADDRPOINTER_REG_0__SCAN_IN, P1_U2376);
  nand ginst6528 (P1_U5800, P1_R2278_U99, P1_U2372);
  nand ginst6529 (P1_U5801, P1_REIP_REG_0__SCAN_IN, P1_U2365);
  nand ginst6530 (P1_U5802, P1_R2358_U76, P1_U2364);
  nand ginst6531 (P1_U5803, P1_PHYADDRPOINTER_REG_0__SCAN_IN, P1_U5795);
  nand ginst6532 (P1_U5804, P1_R2337_U4, P1_U2376);
  nand ginst6533 (P1_U5805, P1_R2278_U19, P1_U2372);
  nand ginst6534 (P1_U5806, P1_REIP_REG_1__SCAN_IN, P1_U2365);
  nand ginst6535 (P1_U5807, P1_R2358_U107, P1_U2364);
  nand ginst6536 (P1_U5808, P1_PHYADDRPOINTER_REG_1__SCAN_IN, P1_U5795);
  nand ginst6537 (P1_U5809, P1_R2337_U71, P1_U2376);
  nand ginst6538 (P1_U5810, P1_R2278_U107, P1_U2372);
  nand ginst6539 (P1_U5811, P1_REIP_REG_2__SCAN_IN, P1_U2365);
  nand ginst6540 (P1_U5812, P1_R2358_U18, P1_U2364);
  nand ginst6541 (P1_U5813, P1_PHYADDRPOINTER_REG_2__SCAN_IN, P1_U5795);
  nand ginst6542 (P1_U5814, P1_R2337_U68, P1_U2376);
  nand ginst6543 (P1_U5815, P1_R2278_U105, P1_U2372);
  nand ginst6544 (P1_U5816, P1_REIP_REG_3__SCAN_IN, P1_U2365);
  nand ginst6545 (P1_U5817, P1_R2358_U19, P1_U2364);
  nand ginst6546 (P1_U5818, P1_PHYADDRPOINTER_REG_3__SCAN_IN, P1_U5795);
  nand ginst6547 (P1_U5819, P1_R2337_U67, P1_U2376);
  nand ginst6548 (P1_U5820, P1_R2278_U104, P1_U2372);
  nand ginst6549 (P1_U5821, P1_REIP_REG_4__SCAN_IN, P1_U2365);
  nand ginst6550 (P1_U5822, P1_R2358_U84, P1_U2364);
  nand ginst6551 (P1_U5823, P1_PHYADDRPOINTER_REG_4__SCAN_IN, P1_U5795);
  nand ginst6552 (P1_U5824, P1_R2337_U66, P1_U2376);
  nand ginst6553 (P1_U5825, P1_R2278_U17, P1_U2372);
  nand ginst6554 (P1_U5826, P1_REIP_REG_5__SCAN_IN, P1_U2365);
  nand ginst6555 (P1_U5827, P1_R2358_U82, P1_U2364);
  nand ginst6556 (P1_U5828, P1_PHYADDRPOINTER_REG_5__SCAN_IN, P1_U5795);
  nand ginst6557 (P1_U5829, P1_R2337_U65, P1_U2376);
  nand ginst6558 (P1_U5830, P1_R2278_U103, P1_U2372);
  nand ginst6559 (P1_U5831, P1_REIP_REG_6__SCAN_IN, P1_U2365);
  nand ginst6560 (P1_U5832, P1_R2358_U20, P1_U2364);
  nand ginst6561 (P1_U5833, P1_PHYADDRPOINTER_REG_6__SCAN_IN, P1_U5795);
  nand ginst6562 (P1_U5834, P1_R2337_U64, P1_U2376);
  nand ginst6563 (P1_U5835, P1_R2278_U18, P1_U2372);
  nand ginst6564 (P1_U5836, P1_REIP_REG_7__SCAN_IN, P1_U2365);
  nand ginst6565 (P1_U5837, P1_R2358_U21, P1_U2364);
  nand ginst6566 (P1_U5838, P1_PHYADDRPOINTER_REG_7__SCAN_IN, P1_U5795);
  nand ginst6567 (P1_U5839, P1_R2337_U63, P1_U2376);
  nand ginst6568 (P1_U5840, P1_R2278_U102, P1_U2372);
  nand ginst6569 (P1_U5841, P1_REIP_REG_8__SCAN_IN, P1_U2365);
  nand ginst6570 (P1_U5842, P1_R2358_U80, P1_U2364);
  nand ginst6571 (P1_U5843, P1_PHYADDRPOINTER_REG_8__SCAN_IN, P1_U5795);
  nand ginst6572 (P1_U5844, P1_R2337_U62, P1_U2376);
  nand ginst6573 (P1_U5845, P1_R2278_U101, P1_U2372);
  nand ginst6574 (P1_U5846, P1_REIP_REG_9__SCAN_IN, P1_U2365);
  nand ginst6575 (P1_U5847, P1_R2358_U78, P1_U2364);
  nand ginst6576 (P1_U5848, P1_PHYADDRPOINTER_REG_9__SCAN_IN, P1_U5795);
  nand ginst6577 (P1_U5849, P1_R2337_U91, P1_U2376);
  nand ginst6578 (P1_U5850, P1_R2278_U126, P1_U2372);
  nand ginst6579 (P1_U5851, P1_REIP_REG_10__SCAN_IN, P1_U2365);
  nand ginst6580 (P1_U5852, P1_R2358_U14, P1_U2364);
  nand ginst6581 (P1_U5853, P1_PHYADDRPOINTER_REG_10__SCAN_IN, P1_U5795);
  nand ginst6582 (P1_U5854, P1_R2337_U90, P1_U2376);
  nand ginst6583 (P1_U5855, P1_R2278_U15, P1_U2372);
  nand ginst6584 (P1_U5856, P1_REIP_REG_11__SCAN_IN, P1_U2365);
  nand ginst6585 (P1_U5857, P1_R2358_U15, P1_U2364);
  nand ginst6586 (P1_U5858, P1_PHYADDRPOINTER_REG_11__SCAN_IN, P1_U5795);
  nand ginst6587 (P1_U5859, P1_R2337_U89, P1_U2376);
  nand ginst6588 (P1_U5860, P1_R2278_U125, P1_U2372);
  nand ginst6589 (P1_U5861, P1_REIP_REG_12__SCAN_IN, P1_U2365);
  nand ginst6590 (P1_U5862, P1_R2358_U119, P1_U2364);
  nand ginst6591 (P1_U5863, P1_PHYADDRPOINTER_REG_12__SCAN_IN, P1_U5795);
  nand ginst6592 (P1_U5864, P1_R2337_U88, P1_U2376);
  nand ginst6593 (P1_U5865, P1_R2278_U123, P1_U2372);
  nand ginst6594 (P1_U5866, P1_REIP_REG_13__SCAN_IN, P1_U2365);
  nand ginst6595 (P1_U5867, P1_R2358_U117, P1_U2364);
  nand ginst6596 (P1_U5868, P1_PHYADDRPOINTER_REG_13__SCAN_IN, P1_U5795);
  nand ginst6597 (P1_U5869, P1_R2337_U87, P1_U2376);
  nand ginst6598 (P1_U5870, P1_R2278_U122, P1_U2372);
  nand ginst6599 (P1_U5871, P1_REIP_REG_14__SCAN_IN, P1_U2365);
  nand ginst6600 (P1_U5872, P1_R2358_U16, P1_U2364);
  nand ginst6601 (P1_U5873, P1_PHYADDRPOINTER_REG_14__SCAN_IN, P1_U5795);
  nand ginst6602 (P1_U5874, P1_R2337_U86, P1_U2376);
  nand ginst6603 (P1_U5875, P1_R2278_U20, P1_U2372);
  nand ginst6604 (P1_U5876, P1_REIP_REG_15__SCAN_IN, P1_U2365);
  nand ginst6605 (P1_U5877, P1_R2358_U17, P1_U2364);
  nand ginst6606 (P1_U5878, P1_PHYADDRPOINTER_REG_15__SCAN_IN, P1_U5795);
  nand ginst6607 (P1_U5879, P1_R2337_U85, P1_U2376);
  nand ginst6608 (P1_U5880, P1_R2278_U121, P1_U2372);
  nand ginst6609 (P1_U5881, P1_REIP_REG_16__SCAN_IN, P1_U2365);
  nand ginst6610 (P1_U5882, P1_R2358_U115, P1_U2364);
  nand ginst6611 (P1_U5883, P1_PHYADDRPOINTER_REG_16__SCAN_IN, P1_U5795);
  nand ginst6612 (P1_U5884, P1_R2337_U84, P1_U2376);
  nand ginst6613 (P1_U5885, P1_R2278_U120, P1_U2372);
  nand ginst6614 (P1_U5886, P1_REIP_REG_17__SCAN_IN, P1_U2365);
  nand ginst6615 (P1_U5887, P1_R2358_U113, P1_U2364);
  nand ginst6616 (P1_U5888, P1_PHYADDRPOINTER_REG_17__SCAN_IN, P1_U5795);
  nand ginst6617 (P1_U5889, P1_R2337_U83, P1_U2376);
  nand ginst6618 (P1_U5890, P1_R2278_U119, P1_U2372);
  nand ginst6619 (P1_U5891, P1_REIP_REG_18__SCAN_IN, P1_U2365);
  nand ginst6620 (P1_U5892, P1_R2358_U111, P1_U2364);
  nand ginst6621 (P1_U5893, P1_PHYADDRPOINTER_REG_18__SCAN_IN, P1_U5795);
  nand ginst6622 (P1_U5894, P1_R2337_U82, P1_U2376);
  nand ginst6623 (P1_U5895, P1_R2278_U118, P1_U2372);
  nand ginst6624 (P1_U5896, P1_REIP_REG_19__SCAN_IN, P1_U2365);
  nand ginst6625 (P1_U5897, P1_R2358_U109, P1_U2364);
  nand ginst6626 (P1_U5898, P1_PHYADDRPOINTER_REG_19__SCAN_IN, P1_U5795);
  nand ginst6627 (P1_U5899, P1_R2337_U81, P1_U2376);
  nand ginst6628 (P1_U5900, P1_R2278_U117, P1_U2372);
  nand ginst6629 (P1_U5901, P1_REIP_REG_20__SCAN_IN, P1_U2365);
  nand ginst6630 (P1_U5902, P1_R2358_U105, P1_U2364);
  nand ginst6631 (P1_U5903, P1_PHYADDRPOINTER_REG_20__SCAN_IN, P1_U5795);
  nand ginst6632 (P1_U5904, P1_R2337_U80, P1_U2376);
  nand ginst6633 (P1_U5905, P1_R2278_U116, P1_U2372);
  nand ginst6634 (P1_U5906, P1_REIP_REG_21__SCAN_IN, P1_U2365);
  nand ginst6635 (P1_U5907, P1_R2358_U103, P1_U2364);
  nand ginst6636 (P1_U5908, P1_PHYADDRPOINTER_REG_21__SCAN_IN, P1_U5795);
  nand ginst6637 (P1_U5909, P1_R2337_U79, P1_U2376);
  nand ginst6638 (P1_U5910, P1_R2278_U115, P1_U2372);
  nand ginst6639 (P1_U5911, P1_REIP_REG_22__SCAN_IN, P1_U2365);
  nand ginst6640 (P1_U5912, P1_R2358_U101, P1_U2364);
  nand ginst6641 (P1_U5913, P1_PHYADDRPOINTER_REG_22__SCAN_IN, P1_U5795);
  nand ginst6642 (P1_U5914, P1_R2337_U78, P1_U2376);
  nand ginst6643 (P1_U5915, P1_R2278_U114, P1_U2372);
  nand ginst6644 (P1_U5916, P1_REIP_REG_23__SCAN_IN, P1_U2365);
  nand ginst6645 (P1_U5917, P1_R2358_U99, P1_U2364);
  nand ginst6646 (P1_U5918, P1_PHYADDRPOINTER_REG_23__SCAN_IN, P1_U5795);
  nand ginst6647 (P1_U5919, P1_R2337_U77, P1_U2376);
  nand ginst6648 (P1_U5920, P1_R2278_U113, P1_U2372);
  nand ginst6649 (P1_U5921, P1_REIP_REG_24__SCAN_IN, P1_U2365);
  nand ginst6650 (P1_U5922, P1_R2358_U97, P1_U2364);
  nand ginst6651 (P1_U5923, P1_PHYADDRPOINTER_REG_24__SCAN_IN, P1_U5795);
  nand ginst6652 (P1_U5924, P1_R2337_U76, P1_U2376);
  nand ginst6653 (P1_U5925, P1_R2278_U112, P1_U2372);
  nand ginst6654 (P1_U5926, P1_REIP_REG_25__SCAN_IN, P1_U2365);
  nand ginst6655 (P1_U5927, P1_R2358_U95, P1_U2364);
  nand ginst6656 (P1_U5928, P1_PHYADDRPOINTER_REG_25__SCAN_IN, P1_U5795);
  nand ginst6657 (P1_U5929, P1_R2337_U75, P1_U2376);
  nand ginst6658 (P1_U5930, P1_R2278_U111, P1_U2372);
  nand ginst6659 (P1_U5931, P1_REIP_REG_26__SCAN_IN, P1_U2365);
  nand ginst6660 (P1_U5932, P1_R2358_U93, P1_U2364);
  nand ginst6661 (P1_U5933, P1_PHYADDRPOINTER_REG_26__SCAN_IN, P1_U5795);
  nand ginst6662 (P1_U5934, P1_R2337_U74, P1_U2376);
  nand ginst6663 (P1_U5935, P1_R2278_U110, P1_U2372);
  nand ginst6664 (P1_U5936, P1_REIP_REG_27__SCAN_IN, P1_U2365);
  nand ginst6665 (P1_U5937, P1_R2358_U91, P1_U2364);
  nand ginst6666 (P1_U5938, P1_PHYADDRPOINTER_REG_27__SCAN_IN, P1_U5795);
  nand ginst6667 (P1_U5939, P1_R2337_U73, P1_U2376);
  nand ginst6668 (P1_U5940, P1_R2278_U109, P1_U2372);
  nand ginst6669 (P1_U5941, P1_REIP_REG_28__SCAN_IN, P1_U2365);
  nand ginst6670 (P1_U5942, P1_R2358_U89, P1_U2364);
  nand ginst6671 (P1_U5943, P1_PHYADDRPOINTER_REG_28__SCAN_IN, P1_U5795);
  nand ginst6672 (P1_U5944, P1_R2337_U72, P1_U2376);
  nand ginst6673 (P1_U5945, P1_R2278_U108, P1_U2372);
  nand ginst6674 (P1_U5946, P1_REIP_REG_29__SCAN_IN, P1_U2365);
  nand ginst6675 (P1_U5947, P1_R2358_U87, P1_U2364);
  nand ginst6676 (P1_U5948, P1_PHYADDRPOINTER_REG_29__SCAN_IN, P1_U5795);
  nand ginst6677 (P1_U5949, P1_R2337_U70, P1_U2376);
  nand ginst6678 (P1_U5950, P1_R2278_U106, P1_U2372);
  nand ginst6679 (P1_U5951, P1_REIP_REG_30__SCAN_IN, P1_U2365);
  nand ginst6680 (P1_U5952, P1_R2358_U85, P1_U2364);
  nand ginst6681 (P1_U5953, P1_PHYADDRPOINTER_REG_30__SCAN_IN, P1_U5795);
  nand ginst6682 (P1_U5954, P1_R2337_U69, P1_U2376);
  nand ginst6683 (P1_U5955, P1_R2278_U16, P1_U2372);
  nand ginst6684 (P1_U5956, P1_REIP_REG_31__SCAN_IN, P1_U2365);
  nand ginst6685 (P1_U5957, P1_R2358_U22, P1_U2364);
  nand ginst6686 (P1_U5958, P1_PHYADDRPOINTER_REG_31__SCAN_IN, P1_U5795);
  nand ginst6687 (P1_U5959, P1_U3282, U210);
  nand ginst6688 (P1_U5960, P1_EAX_REG_15__SCAN_IN, P1_U2382);
  nand ginst6689 (P1_U5961, P1_U2381, U340);
  nand ginst6690 (P1_U5962, P1_U5960, P1_U5961);
  nand ginst6691 (P1_U5963, P1_EAX_REG_14__SCAN_IN, P1_U2382);
  nand ginst6692 (P1_U5964, P1_U2381, U341);
  nand ginst6693 (P1_U5965, P1_U5963, P1_U5964);
  nand ginst6694 (P1_U5966, P1_EAX_REG_13__SCAN_IN, P1_U2382);
  nand ginst6695 (P1_U5967, P1_U2381, U342);
  nand ginst6696 (P1_U5968, P1_U5966, P1_U5967);
  nand ginst6697 (P1_U5969, P1_EAX_REG_12__SCAN_IN, P1_U2382);
  nand ginst6698 (P1_U5970, P1_U2381, U343);
  nand ginst6699 (P1_U5971, P1_U5969, P1_U5970);
  nand ginst6700 (P1_U5972, P1_EAX_REG_11__SCAN_IN, P1_U2382);
  nand ginst6701 (P1_U5973, P1_U2381, U344);
  nand ginst6702 (P1_U5974, P1_U5972, P1_U5973);
  nand ginst6703 (P1_U5975, P1_EAX_REG_10__SCAN_IN, P1_U2382);
  nand ginst6704 (P1_U5976, P1_U2381, U345);
  nand ginst6705 (P1_U5977, P1_U5975, P1_U5976);
  nand ginst6706 (P1_U5978, P1_EAX_REG_9__SCAN_IN, P1_U2382);
  nand ginst6707 (P1_U5979, P1_U2381, U315);
  nand ginst6708 (P1_U5980, P1_U5978, P1_U5979);
  nand ginst6709 (P1_U5981, P1_EAX_REG_8__SCAN_IN, P1_U2382);
  nand ginst6710 (P1_U5982, P1_U2381, U316);
  nand ginst6711 (P1_U5983, P1_U5981, P1_U5982);
  nand ginst6712 (P1_U5984, P1_EAX_REG_7__SCAN_IN, P1_U2382);
  nand ginst6713 (P1_U5985, P1_U2381, U317);
  nand ginst6714 (P1_U5986, P1_U5984, P1_U5985);
  nand ginst6715 (P1_U5987, P1_EAX_REG_6__SCAN_IN, P1_U2382);
  nand ginst6716 (P1_U5988, P1_U2381, U318);
  nand ginst6717 (P1_U5989, P1_U5987, P1_U5988);
  nand ginst6718 (P1_U5990, P1_EAX_REG_5__SCAN_IN, P1_U2382);
  nand ginst6719 (P1_U5991, P1_U2381, U319);
  nand ginst6720 (P1_U5992, P1_U5990, P1_U5991);
  nand ginst6721 (P1_U5993, P1_EAX_REG_4__SCAN_IN, P1_U2382);
  nand ginst6722 (P1_U5994, P1_U2381, U320);
  nand ginst6723 (P1_U5995, P1_U5993, P1_U5994);
  nand ginst6724 (P1_U5996, P1_EAX_REG_3__SCAN_IN, P1_U2382);
  nand ginst6725 (P1_U5997, P1_U2381, U321);
  nand ginst6726 (P1_U5998, P1_U5996, P1_U5997);
  nand ginst6727 (P1_U5999, P1_EAX_REG_2__SCAN_IN, P1_U2382);
  nand ginst6728 (P1_U6000, P1_U2381, U324);
  nand ginst6729 (P1_U6001, P1_U5999, P1_U6000);
  nand ginst6730 (P1_U6002, P1_EAX_REG_1__SCAN_IN, P1_U2382);
  nand ginst6731 (P1_U6003, P1_U2381, U335);
  nand ginst6732 (P1_U6004, P1_U6002, P1_U6003);
  nand ginst6733 (P1_U6005, P1_EAX_REG_0__SCAN_IN, P1_U2382);
  nand ginst6734 (P1_U6006, P1_U2381, U346);
  nand ginst6735 (P1_U6007, P1_U6005, P1_U6006);
  nand ginst6736 (P1_U6008, P1_EAX_REG_30__SCAN_IN, P1_U2382);
  nand ginst6737 (P1_U6009, P1_U2381, U341);
  nand ginst6738 (P1_U6010, P1_U6008, P1_U6009);
  nand ginst6739 (P1_U6011, P1_EAX_REG_29__SCAN_IN, P1_U2382);
  nand ginst6740 (P1_U6012, P1_U2381, U342);
  nand ginst6741 (P1_U6013, P1_U6011, P1_U6012);
  nand ginst6742 (P1_U6014, P1_EAX_REG_28__SCAN_IN, P1_U2382);
  nand ginst6743 (P1_U6015, P1_U2381, U343);
  nand ginst6744 (P1_U6016, P1_U6014, P1_U6015);
  nand ginst6745 (P1_U6017, P1_EAX_REG_27__SCAN_IN, P1_U2382);
  nand ginst6746 (P1_U6018, P1_U2381, U344);
  nand ginst6747 (P1_U6019, P1_U6017, P1_U6018);
  nand ginst6748 (P1_U6020, P1_EAX_REG_26__SCAN_IN, P1_U2382);
  nand ginst6749 (P1_U6021, P1_U2381, U345);
  nand ginst6750 (P1_U6022, P1_U6020, P1_U6021);
  nand ginst6751 (P1_U6023, P1_EAX_REG_25__SCAN_IN, P1_U2382);
  nand ginst6752 (P1_U6024, P1_U2381, U315);
  nand ginst6753 (P1_U6025, P1_U6023, P1_U6024);
  nand ginst6754 (P1_U6026, P1_EAX_REG_24__SCAN_IN, P1_U2382);
  nand ginst6755 (P1_U6027, P1_U2381, U316);
  nand ginst6756 (P1_U6028, P1_U6026, P1_U6027);
  nand ginst6757 (P1_U6029, P1_EAX_REG_23__SCAN_IN, P1_U2382);
  nand ginst6758 (P1_U6030, P1_U2381, U317);
  nand ginst6759 (P1_U6031, P1_U6029, P1_U6030);
  nand ginst6760 (P1_U6032, P1_EAX_REG_22__SCAN_IN, P1_U2382);
  nand ginst6761 (P1_U6033, P1_U2381, U318);
  nand ginst6762 (P1_U6034, P1_U6032, P1_U6033);
  nand ginst6763 (P1_U6035, P1_EAX_REG_21__SCAN_IN, P1_U2382);
  nand ginst6764 (P1_U6036, P1_U2381, U319);
  nand ginst6765 (P1_U6037, P1_U6035, P1_U6036);
  nand ginst6766 (P1_U6038, P1_EAX_REG_20__SCAN_IN, P1_U2382);
  nand ginst6767 (P1_U6039, P1_U2381, U320);
  nand ginst6768 (P1_U6040, P1_U6038, P1_U6039);
  nand ginst6769 (P1_U6041, P1_EAX_REG_19__SCAN_IN, P1_U2382);
  nand ginst6770 (P1_U6042, P1_U2381, U321);
  nand ginst6771 (P1_U6043, P1_U6041, P1_U6042);
  nand ginst6772 (P1_U6044, P1_EAX_REG_18__SCAN_IN, P1_U2382);
  nand ginst6773 (P1_U6045, P1_U2381, U324);
  nand ginst6774 (P1_U6046, P1_U6044, P1_U6045);
  nand ginst6775 (P1_U6047, P1_EAX_REG_17__SCAN_IN, P1_U2382);
  nand ginst6776 (P1_U6048, P1_U2381, U335);
  nand ginst6777 (P1_U6049, P1_U6047, P1_U6048);
  nand ginst6778 (P1_U6050, P1_EAX_REG_16__SCAN_IN, P1_U2382);
  nand ginst6779 (P1_U6051, P1_U2381, U346);
  nand ginst6780 (P1_U6052, P1_U6050, P1_U6051);
  nand ginst6781 (P1_U6053, P1_U4235, P1_U4259, P1_U7606);
  nand ginst6782 (P1_U6054, P1_U2428, P1_U3294);
  not ginst6783 (P1_U6055, P1_U3417);
  nand ginst6784 (P1_U6056, P1_LWORD_REG_0__SCAN_IN, P1_U2385);
  nand ginst6785 (P1_U6057, P1_EAX_REG_0__SCAN_IN, P1_U2384);
  nand ginst6786 (P1_U6058, P1_DATAO_REG_0__SCAN_IN, P1_U6055);
  nand ginst6787 (P1_U6059, P1_LWORD_REG_1__SCAN_IN, P1_U2385);
  nand ginst6788 (P1_U6060, P1_EAX_REG_1__SCAN_IN, P1_U2384);
  nand ginst6789 (P1_U6061, P1_DATAO_REG_1__SCAN_IN, P1_U6055);
  nand ginst6790 (P1_U6062, P1_LWORD_REG_2__SCAN_IN, P1_U2385);
  nand ginst6791 (P1_U6063, P1_EAX_REG_2__SCAN_IN, P1_U2384);
  nand ginst6792 (P1_U6064, P1_DATAO_REG_2__SCAN_IN, P1_U6055);
  nand ginst6793 (P1_U6065, P1_LWORD_REG_3__SCAN_IN, P1_U2385);
  nand ginst6794 (P1_U6066, P1_EAX_REG_3__SCAN_IN, P1_U2384);
  nand ginst6795 (P1_U6067, P1_DATAO_REG_3__SCAN_IN, P1_U6055);
  nand ginst6796 (P1_U6068, P1_LWORD_REG_4__SCAN_IN, P1_U2385);
  nand ginst6797 (P1_U6069, P1_EAX_REG_4__SCAN_IN, P1_U2384);
  nand ginst6798 (P1_U6070, P1_DATAO_REG_4__SCAN_IN, P1_U6055);
  nand ginst6799 (P1_U6071, P1_LWORD_REG_5__SCAN_IN, P1_U2385);
  nand ginst6800 (P1_U6072, P1_EAX_REG_5__SCAN_IN, P1_U2384);
  nand ginst6801 (P1_U6073, P1_DATAO_REG_5__SCAN_IN, P1_U6055);
  nand ginst6802 (P1_U6074, P1_LWORD_REG_6__SCAN_IN, P1_U2385);
  nand ginst6803 (P1_U6075, P1_EAX_REG_6__SCAN_IN, P1_U2384);
  nand ginst6804 (P1_U6076, P1_DATAO_REG_6__SCAN_IN, P1_U6055);
  nand ginst6805 (P1_U6077, P1_LWORD_REG_7__SCAN_IN, P1_U2385);
  nand ginst6806 (P1_U6078, P1_EAX_REG_7__SCAN_IN, P1_U2384);
  nand ginst6807 (P1_U6079, P1_DATAO_REG_7__SCAN_IN, P1_U6055);
  nand ginst6808 (P1_U6080, P1_LWORD_REG_8__SCAN_IN, P1_U2385);
  nand ginst6809 (P1_U6081, P1_EAX_REG_8__SCAN_IN, P1_U2384);
  nand ginst6810 (P1_U6082, P1_DATAO_REG_8__SCAN_IN, P1_U6055);
  nand ginst6811 (P1_U6083, P1_LWORD_REG_9__SCAN_IN, P1_U2385);
  nand ginst6812 (P1_U6084, P1_EAX_REG_9__SCAN_IN, P1_U2384);
  nand ginst6813 (P1_U6085, P1_DATAO_REG_9__SCAN_IN, P1_U6055);
  nand ginst6814 (P1_U6086, P1_LWORD_REG_10__SCAN_IN, P1_U2385);
  nand ginst6815 (P1_U6087, P1_EAX_REG_10__SCAN_IN, P1_U2384);
  nand ginst6816 (P1_U6088, P1_DATAO_REG_10__SCAN_IN, P1_U6055);
  nand ginst6817 (P1_U6089, P1_LWORD_REG_11__SCAN_IN, P1_U2385);
  nand ginst6818 (P1_U6090, P1_EAX_REG_11__SCAN_IN, P1_U2384);
  nand ginst6819 (P1_U6091, P1_DATAO_REG_11__SCAN_IN, P1_U6055);
  nand ginst6820 (P1_U6092, P1_LWORD_REG_12__SCAN_IN, P1_U2385);
  nand ginst6821 (P1_U6093, P1_EAX_REG_12__SCAN_IN, P1_U2384);
  nand ginst6822 (P1_U6094, P1_DATAO_REG_12__SCAN_IN, P1_U6055);
  nand ginst6823 (P1_U6095, P1_LWORD_REG_13__SCAN_IN, P1_U2385);
  nand ginst6824 (P1_U6096, P1_EAX_REG_13__SCAN_IN, P1_U2384);
  nand ginst6825 (P1_U6097, P1_DATAO_REG_13__SCAN_IN, P1_U6055);
  nand ginst6826 (P1_U6098, P1_LWORD_REG_14__SCAN_IN, P1_U2385);
  nand ginst6827 (P1_U6099, P1_EAX_REG_14__SCAN_IN, P1_U2384);
  nand ginst6828 (P1_U6100, P1_DATAO_REG_14__SCAN_IN, P1_U6055);
  nand ginst6829 (P1_U6101, P1_LWORD_REG_15__SCAN_IN, P1_U2385);
  nand ginst6830 (P1_U6102, P1_EAX_REG_15__SCAN_IN, P1_U2384);
  nand ginst6831 (P1_U6103, P1_DATAO_REG_15__SCAN_IN, P1_U6055);
  nand ginst6832 (P1_U6104, P1_EAX_REG_16__SCAN_IN, P1_U2424);
  nand ginst6833 (P1_U6105, P1_UWORD_REG_0__SCAN_IN, P1_U2385);
  nand ginst6834 (P1_U6106, P1_DATAO_REG_16__SCAN_IN, P1_U6055);
  nand ginst6835 (P1_U6107, P1_EAX_REG_17__SCAN_IN, P1_U2424);
  nand ginst6836 (P1_U6108, P1_UWORD_REG_1__SCAN_IN, P1_U2385);
  nand ginst6837 (P1_U6109, P1_DATAO_REG_17__SCAN_IN, P1_U6055);
  nand ginst6838 (P1_U6110, P1_EAX_REG_18__SCAN_IN, P1_U2424);
  nand ginst6839 (P1_U6111, P1_UWORD_REG_2__SCAN_IN, P1_U2385);
  nand ginst6840 (P1_U6112, P1_DATAO_REG_18__SCAN_IN, P1_U6055);
  nand ginst6841 (P1_U6113, P1_EAX_REG_19__SCAN_IN, P1_U2424);
  nand ginst6842 (P1_U6114, P1_UWORD_REG_3__SCAN_IN, P1_U2385);
  nand ginst6843 (P1_U6115, P1_DATAO_REG_19__SCAN_IN, P1_U6055);
  nand ginst6844 (P1_U6116, P1_EAX_REG_20__SCAN_IN, P1_U2424);
  nand ginst6845 (P1_U6117, P1_UWORD_REG_4__SCAN_IN, P1_U2385);
  nand ginst6846 (P1_U6118, P1_DATAO_REG_20__SCAN_IN, P1_U6055);
  nand ginst6847 (P1_U6119, P1_EAX_REG_21__SCAN_IN, P1_U2424);
  nand ginst6848 (P1_U6120, P1_UWORD_REG_5__SCAN_IN, P1_U2385);
  nand ginst6849 (P1_U6121, P1_DATAO_REG_21__SCAN_IN, P1_U6055);
  nand ginst6850 (P1_U6122, P1_EAX_REG_22__SCAN_IN, P1_U2424);
  nand ginst6851 (P1_U6123, P1_UWORD_REG_6__SCAN_IN, P1_U2385);
  nand ginst6852 (P1_U6124, P1_DATAO_REG_22__SCAN_IN, P1_U6055);
  nand ginst6853 (P1_U6125, P1_EAX_REG_23__SCAN_IN, P1_U2424);
  nand ginst6854 (P1_U6126, P1_UWORD_REG_7__SCAN_IN, P1_U2385);
  nand ginst6855 (P1_U6127, P1_DATAO_REG_23__SCAN_IN, P1_U6055);
  nand ginst6856 (P1_U6128, P1_EAX_REG_24__SCAN_IN, P1_U2424);
  nand ginst6857 (P1_U6129, P1_UWORD_REG_8__SCAN_IN, P1_U2385);
  nand ginst6858 (P1_U6130, P1_DATAO_REG_24__SCAN_IN, P1_U6055);
  nand ginst6859 (P1_U6131, P1_EAX_REG_25__SCAN_IN, P1_U2424);
  nand ginst6860 (P1_U6132, P1_UWORD_REG_9__SCAN_IN, P1_U2385);
  nand ginst6861 (P1_U6133, P1_DATAO_REG_25__SCAN_IN, P1_U6055);
  nand ginst6862 (P1_U6134, P1_EAX_REG_26__SCAN_IN, P1_U2424);
  nand ginst6863 (P1_U6135, P1_UWORD_REG_10__SCAN_IN, P1_U2385);
  nand ginst6864 (P1_U6136, P1_DATAO_REG_26__SCAN_IN, P1_U6055);
  nand ginst6865 (P1_U6137, P1_EAX_REG_27__SCAN_IN, P1_U2424);
  nand ginst6866 (P1_U6138, P1_UWORD_REG_11__SCAN_IN, P1_U2385);
  nand ginst6867 (P1_U6139, P1_DATAO_REG_27__SCAN_IN, P1_U6055);
  nand ginst6868 (P1_U6140, P1_EAX_REG_28__SCAN_IN, P1_U2424);
  nand ginst6869 (P1_U6141, P1_UWORD_REG_12__SCAN_IN, P1_U2385);
  nand ginst6870 (P1_U6142, P1_DATAO_REG_28__SCAN_IN, P1_U6055);
  nand ginst6871 (P1_U6143, P1_EAX_REG_29__SCAN_IN, P1_U2424);
  nand ginst6872 (P1_U6144, P1_UWORD_REG_13__SCAN_IN, P1_U2385);
  nand ginst6873 (P1_U6145, P1_DATAO_REG_29__SCAN_IN, P1_U6055);
  nand ginst6874 (P1_U6146, P1_EAX_REG_30__SCAN_IN, P1_U2424);
  nand ginst6875 (P1_U6147, P1_UWORD_REG_14__SCAN_IN, P1_U2385);
  nand ginst6876 (P1_U6148, P1_DATAO_REG_30__SCAN_IN, P1_U6055);
  nand ginst6877 (P1_U6149, P1_GTE_485_U6, P1_U2447, P1_U4194);
  nand ginst6878 (P1_U6150, P1_U4194, P1_U4197, P1_U4254);
  nand ginst6879 (P1_U6151, P1_R2167_U17, P1_U3283, P1_U4200);
  nand ginst6880 (P1_U6152, P1_U3257, P1_U7503);
  nand ginst6881 (P1_U6153, P1_U3883, P1_U6152);
  nand ginst6882 (P1_U6154, P1_U2422, U346);
  nand ginst6883 (P1_U6155, P1_R2358_U76, P1_U2386);
  nand ginst6884 (P1_U6156, P1_EAX_REG_0__SCAN_IN, P1_U3424);
  nand ginst6885 (P1_U6157, P1_U2422, U335);
  nand ginst6886 (P1_U6158, P1_R2358_U107, P1_U2386);
  nand ginst6887 (P1_U6159, P1_EAX_REG_1__SCAN_IN, P1_U3424);
  nand ginst6888 (P1_U6160, P1_U2422, U324);
  nand ginst6889 (P1_U6161, P1_R2358_U18, P1_U2386);
  nand ginst6890 (P1_U6162, P1_EAX_REG_2__SCAN_IN, P1_U3424);
  nand ginst6891 (P1_U6163, P1_U2422, U321);
  nand ginst6892 (P1_U6164, P1_R2358_U19, P1_U2386);
  nand ginst6893 (P1_U6165, P1_EAX_REG_3__SCAN_IN, P1_U3424);
  nand ginst6894 (P1_U6166, P1_U2422, U320);
  nand ginst6895 (P1_U6167, P1_R2358_U84, P1_U2386);
  nand ginst6896 (P1_U6168, P1_EAX_REG_4__SCAN_IN, P1_U3424);
  nand ginst6897 (P1_U6169, P1_U2422, U319);
  nand ginst6898 (P1_U6170, P1_R2358_U82, P1_U2386);
  nand ginst6899 (P1_U6171, P1_EAX_REG_5__SCAN_IN, P1_U3424);
  nand ginst6900 (P1_U6172, P1_U2422, U318);
  nand ginst6901 (P1_U6173, P1_R2358_U20, P1_U2386);
  nand ginst6902 (P1_U6174, P1_EAX_REG_6__SCAN_IN, P1_U3424);
  nand ginst6903 (P1_U6175, P1_U2422, U317);
  nand ginst6904 (P1_U6176, P1_R2358_U21, P1_U2386);
  nand ginst6905 (P1_U6177, P1_EAX_REG_7__SCAN_IN, P1_U3424);
  nand ginst6906 (P1_U6178, P1_U2422, U316);
  nand ginst6907 (P1_U6179, P1_R2358_U80, P1_U2386);
  nand ginst6908 (P1_U6180, P1_EAX_REG_8__SCAN_IN, P1_U3424);
  nand ginst6909 (P1_U6181, P1_U2422, U315);
  nand ginst6910 (P1_U6182, P1_R2358_U78, P1_U2386);
  nand ginst6911 (P1_U6183, P1_EAX_REG_9__SCAN_IN, P1_U3424);
  nand ginst6912 (P1_U6184, P1_U2422, U345);
  nand ginst6913 (P1_U6185, P1_R2358_U14, P1_U2386);
  nand ginst6914 (P1_U6186, P1_EAX_REG_10__SCAN_IN, P1_U3424);
  nand ginst6915 (P1_U6187, P1_U2422, U344);
  nand ginst6916 (P1_U6188, P1_R2358_U15, P1_U2386);
  nand ginst6917 (P1_U6189, P1_EAX_REG_11__SCAN_IN, P1_U3424);
  nand ginst6918 (P1_U6190, P1_U2422, U343);
  nand ginst6919 (P1_U6191, P1_R2358_U119, P1_U2386);
  nand ginst6920 (P1_U6192, P1_EAX_REG_12__SCAN_IN, P1_U3424);
  nand ginst6921 (P1_U6193, P1_U2422, U342);
  nand ginst6922 (P1_U6194, P1_R2358_U117, P1_U2386);
  nand ginst6923 (P1_U6195, P1_EAX_REG_13__SCAN_IN, P1_U3424);
  nand ginst6924 (P1_U6196, P1_U2422, U341);
  nand ginst6925 (P1_U6197, P1_R2358_U16, P1_U2386);
  nand ginst6926 (P1_U6198, P1_EAX_REG_14__SCAN_IN, P1_U3424);
  nand ginst6927 (P1_U6199, P1_U2422, U340);
  nand ginst6928 (P1_U6200, P1_R2358_U17, P1_U2386);
  nand ginst6929 (P1_U6201, P1_EAX_REG_15__SCAN_IN, P1_U3424);
  nand ginst6930 (P1_U6202, P1_U2423, U339);
  nand ginst6931 (P1_U6203, P1_U2387, U346);
  nand ginst6932 (P1_U6204, P1_R2358_U115, P1_U2386);
  nand ginst6933 (P1_U6205, P1_EAX_REG_16__SCAN_IN, P1_U3424);
  nand ginst6934 (P1_U6206, P1_U2423, U338);
  nand ginst6935 (P1_U6207, P1_U2387, U335);
  nand ginst6936 (P1_U6208, P1_R2358_U113, P1_U2386);
  nand ginst6937 (P1_U6209, P1_EAX_REG_17__SCAN_IN, P1_U3424);
  nand ginst6938 (P1_U6210, P1_U2423, U337);
  nand ginst6939 (P1_U6211, P1_U2387, U324);
  nand ginst6940 (P1_U6212, P1_R2358_U111, P1_U2386);
  nand ginst6941 (P1_U6213, P1_EAX_REG_18__SCAN_IN, P1_U3424);
  nand ginst6942 (P1_U6214, P1_U2423, U336);
  nand ginst6943 (P1_U6215, P1_U2387, U321);
  nand ginst6944 (P1_U6216, P1_R2358_U109, P1_U2386);
  nand ginst6945 (P1_U6217, P1_EAX_REG_19__SCAN_IN, P1_U3424);
  nand ginst6946 (P1_U6218, P1_U2423, U334);
  nand ginst6947 (P1_U6219, P1_U2387, U320);
  nand ginst6948 (P1_U6220, P1_R2358_U105, P1_U2386);
  nand ginst6949 (P1_U6221, P1_EAX_REG_20__SCAN_IN, P1_U3424);
  nand ginst6950 (P1_U6222, P1_U2423, U333);
  nand ginst6951 (P1_U6223, P1_U2387, U319);
  nand ginst6952 (P1_U6224, P1_R2358_U103, P1_U2386);
  nand ginst6953 (P1_U6225, P1_EAX_REG_21__SCAN_IN, P1_U3424);
  nand ginst6954 (P1_U6226, P1_U2423, U332);
  nand ginst6955 (P1_U6227, P1_U2387, U318);
  nand ginst6956 (P1_U6228, P1_R2358_U101, P1_U2386);
  nand ginst6957 (P1_U6229, P1_EAX_REG_22__SCAN_IN, P1_U3424);
  nand ginst6958 (P1_U6230, P1_U2423, U331);
  nand ginst6959 (P1_U6231, P1_U2387, U317);
  nand ginst6960 (P1_U6232, P1_R2358_U99, P1_U2386);
  nand ginst6961 (P1_U6233, P1_EAX_REG_23__SCAN_IN, P1_U3424);
  nand ginst6962 (P1_U6234, P1_U2423, U330);
  nand ginst6963 (P1_U6235, P1_U2387, U316);
  nand ginst6964 (P1_U6236, P1_R2358_U97, P1_U2386);
  nand ginst6965 (P1_U6237, P1_EAX_REG_24__SCAN_IN, P1_U3424);
  nand ginst6966 (P1_U6238, P1_U2423, U329);
  nand ginst6967 (P1_U6239, P1_U2387, U315);
  nand ginst6968 (P1_U6240, P1_R2358_U95, P1_U2386);
  nand ginst6969 (P1_U6241, P1_EAX_REG_25__SCAN_IN, P1_U3424);
  nand ginst6970 (P1_U6242, P1_U2423, U328);
  nand ginst6971 (P1_U6243, P1_U2387, U345);
  nand ginst6972 (P1_U6244, P1_R2358_U93, P1_U2386);
  nand ginst6973 (P1_U6245, P1_EAX_REG_26__SCAN_IN, P1_U3424);
  nand ginst6974 (P1_U6246, P1_U2423, U327);
  nand ginst6975 (P1_U6247, P1_U2387, U344);
  nand ginst6976 (P1_U6248, P1_R2358_U91, P1_U2386);
  nand ginst6977 (P1_U6249, P1_EAX_REG_27__SCAN_IN, P1_U3424);
  nand ginst6978 (P1_U6250, P1_U2423, U326);
  nand ginst6979 (P1_U6251, P1_U2387, U343);
  nand ginst6980 (P1_U6252, P1_R2358_U89, P1_U2386);
  nand ginst6981 (P1_U6253, P1_EAX_REG_28__SCAN_IN, P1_U3424);
  nand ginst6982 (P1_U6254, P1_U2423, U325);
  nand ginst6983 (P1_U6255, P1_U2387, U342);
  nand ginst6984 (P1_U6256, P1_R2358_U87, P1_U2386);
  nand ginst6985 (P1_U6257, P1_EAX_REG_29__SCAN_IN, P1_U3424);
  nand ginst6986 (P1_U6258, P1_U2423, U323);
  nand ginst6987 (P1_U6259, P1_U2387, U341);
  nand ginst6988 (P1_U6260, P1_R2358_U85, P1_U2386);
  nand ginst6989 (P1_U6261, P1_EAX_REG_30__SCAN_IN, P1_U3424);
  nand ginst6990 (P1_U6262, P1_U2423, U322);
  nand ginst6991 (P1_U6263, P1_U3273, P1_U4198);
  nand ginst6992 (P1_U6264, P1_U4205, P1_U6263);
  nand ginst6993 (P1_U6265, P1_R2358_U76, P1_U2383);
  nand ginst6994 (P1_U6266, P1_R2099_U86, P1_U2371);
  nand ginst6995 (P1_U6267, P1_EBX_REG_0__SCAN_IN, P1_U3426);
  nand ginst6996 (P1_U6268, P1_R2358_U107, P1_U2383);
  nand ginst6997 (P1_U6269, P1_R2099_U87, P1_U2371);
  nand ginst6998 (P1_U6270, P1_EBX_REG_1__SCAN_IN, P1_U3426);
  nand ginst6999 (P1_U6271, P1_R2358_U18, P1_U2383);
  nand ginst7000 (P1_U6272, P1_R2099_U138, P1_U2371);
  nand ginst7001 (P1_U6273, P1_EBX_REG_2__SCAN_IN, P1_U3426);
  nand ginst7002 (P1_U6274, P1_R2358_U19, P1_U2383);
  nand ginst7003 (P1_U6275, P1_R2099_U42, P1_U2371);
  nand ginst7004 (P1_U6276, P1_EBX_REG_3__SCAN_IN, P1_U3426);
  nand ginst7005 (P1_U6277, P1_R2358_U84, P1_U2383);
  nand ginst7006 (P1_U6278, P1_R2099_U41, P1_U2371);
  nand ginst7007 (P1_U6279, P1_EBX_REG_4__SCAN_IN, P1_U3426);
  nand ginst7008 (P1_U6280, P1_R2358_U82, P1_U2383);
  nand ginst7009 (P1_U6281, P1_R2099_U40, P1_U2371);
  nand ginst7010 (P1_U6282, P1_EBX_REG_5__SCAN_IN, P1_U3426);
  nand ginst7011 (P1_U6283, P1_R2358_U20, P1_U2383);
  nand ginst7012 (P1_U6284, P1_R2099_U39, P1_U2371);
  nand ginst7013 (P1_U6285, P1_EBX_REG_6__SCAN_IN, P1_U3426);
  nand ginst7014 (P1_U6286, P1_R2358_U21, P1_U2383);
  nand ginst7015 (P1_U6287, P1_R2099_U38, P1_U2371);
  nand ginst7016 (P1_U6288, P1_EBX_REG_7__SCAN_IN, P1_U3426);
  nand ginst7017 (P1_U6289, P1_R2358_U80, P1_U2383);
  nand ginst7018 (P1_U6290, P1_R2099_U37, P1_U2371);
  nand ginst7019 (P1_U6291, P1_EBX_REG_8__SCAN_IN, P1_U3426);
  nand ginst7020 (P1_U6292, P1_R2358_U78, P1_U2383);
  nand ginst7021 (P1_U6293, P1_R2099_U36, P1_U2371);
  nand ginst7022 (P1_U6294, P1_EBX_REG_9__SCAN_IN, P1_U3426);
  nand ginst7023 (P1_U6295, P1_R2358_U14, P1_U2383);
  nand ginst7024 (P1_U6296, P1_R2099_U85, P1_U2371);
  nand ginst7025 (P1_U6297, P1_EBX_REG_10__SCAN_IN, P1_U3426);
  nand ginst7026 (P1_U6298, P1_R2358_U15, P1_U2383);
  nand ginst7027 (P1_U6299, P1_R2099_U84, P1_U2371);
  nand ginst7028 (P1_U6300, P1_EBX_REG_11__SCAN_IN, P1_U3426);
  nand ginst7029 (P1_U6301, P1_R2358_U119, P1_U2383);
  nand ginst7030 (P1_U6302, P1_R2099_U83, P1_U2371);
  nand ginst7031 (P1_U6303, P1_EBX_REG_12__SCAN_IN, P1_U3426);
  nand ginst7032 (P1_U6304, P1_R2358_U117, P1_U2383);
  nand ginst7033 (P1_U6305, P1_R2099_U82, P1_U2371);
  nand ginst7034 (P1_U6306, P1_EBX_REG_13__SCAN_IN, P1_U3426);
  nand ginst7035 (P1_U6307, P1_R2358_U16, P1_U2383);
  nand ginst7036 (P1_U6308, P1_R2099_U81, P1_U2371);
  nand ginst7037 (P1_U6309, P1_EBX_REG_14__SCAN_IN, P1_U3426);
  nand ginst7038 (P1_U6310, P1_R2358_U17, P1_U2383);
  nand ginst7039 (P1_U6311, P1_R2099_U80, P1_U2371);
  nand ginst7040 (P1_U6312, P1_EBX_REG_15__SCAN_IN, P1_U3426);
  nand ginst7041 (P1_U6313, P1_R2358_U115, P1_U2383);
  nand ginst7042 (P1_U6314, P1_R2099_U79, P1_U2371);
  nand ginst7043 (P1_U6315, P1_EBX_REG_16__SCAN_IN, P1_U3426);
  nand ginst7044 (P1_U6316, P1_R2358_U113, P1_U2383);
  nand ginst7045 (P1_U6317, P1_R2099_U78, P1_U2371);
  nand ginst7046 (P1_U6318, P1_EBX_REG_17__SCAN_IN, P1_U3426);
  nand ginst7047 (P1_U6319, P1_R2358_U111, P1_U2383);
  nand ginst7048 (P1_U6320, P1_R2099_U77, P1_U2371);
  nand ginst7049 (P1_U6321, P1_EBX_REG_18__SCAN_IN, P1_U3426);
  nand ginst7050 (P1_U6322, P1_R2358_U109, P1_U2383);
  nand ginst7051 (P1_U6323, P1_R2099_U76, P1_U2371);
  nand ginst7052 (P1_U6324, P1_EBX_REG_19__SCAN_IN, P1_U3426);
  nand ginst7053 (P1_U6325, P1_R2358_U105, P1_U2383);
  nand ginst7054 (P1_U6326, P1_R2099_U75, P1_U2371);
  nand ginst7055 (P1_U6327, P1_EBX_REG_20__SCAN_IN, P1_U3426);
  nand ginst7056 (P1_U6328, P1_R2358_U103, P1_U2383);
  nand ginst7057 (P1_U6329, P1_R2099_U74, P1_U2371);
  nand ginst7058 (P1_U6330, P1_EBX_REG_21__SCAN_IN, P1_U3426);
  nand ginst7059 (P1_U6331, P1_R2358_U101, P1_U2383);
  nand ginst7060 (P1_U6332, P1_R2099_U73, P1_U2371);
  nand ginst7061 (P1_U6333, P1_EBX_REG_22__SCAN_IN, P1_U3426);
  nand ginst7062 (P1_U6334, P1_R2358_U99, P1_U2383);
  nand ginst7063 (P1_U6335, P1_R2099_U72, P1_U2371);
  nand ginst7064 (P1_U6336, P1_EBX_REG_23__SCAN_IN, P1_U3426);
  nand ginst7065 (P1_U6337, P1_R2358_U97, P1_U2383);
  nand ginst7066 (P1_U6338, P1_R2099_U71, P1_U2371);
  nand ginst7067 (P1_U6339, P1_EBX_REG_24__SCAN_IN, P1_U3426);
  nand ginst7068 (P1_U6340, P1_R2358_U95, P1_U2383);
  nand ginst7069 (P1_U6341, P1_R2099_U70, P1_U2371);
  nand ginst7070 (P1_U6342, P1_EBX_REG_25__SCAN_IN, P1_U3426);
  nand ginst7071 (P1_U6343, P1_R2358_U93, P1_U2383);
  nand ginst7072 (P1_U6344, P1_R2099_U69, P1_U2371);
  nand ginst7073 (P1_U6345, P1_EBX_REG_26__SCAN_IN, P1_U3426);
  nand ginst7074 (P1_U6346, P1_R2358_U91, P1_U2383);
  nand ginst7075 (P1_U6347, P1_R2099_U68, P1_U2371);
  nand ginst7076 (P1_U6348, P1_EBX_REG_27__SCAN_IN, P1_U3426);
  nand ginst7077 (P1_U6349, P1_R2358_U89, P1_U2383);
  nand ginst7078 (P1_U6350, P1_R2099_U67, P1_U2371);
  nand ginst7079 (P1_U6351, P1_EBX_REG_28__SCAN_IN, P1_U3426);
  nand ginst7080 (P1_U6352, P1_R2358_U87, P1_U2383);
  nand ginst7081 (P1_U6353, P1_R2099_U66, P1_U2371);
  nand ginst7082 (P1_U6354, P1_EBX_REG_29__SCAN_IN, P1_U3426);
  nand ginst7083 (P1_U6355, P1_R2358_U85, P1_U2383);
  nand ginst7084 (P1_U6356, P1_R2099_U65, P1_U2371);
  nand ginst7085 (P1_U6357, P1_EBX_REG_30__SCAN_IN, P1_U3426);
  nand ginst7086 (P1_U6358, P1_R2099_U64, P1_U2371);
  nand ginst7087 (P1_U6359, P1_EBX_REG_31__SCAN_IN, P1_U3426);
  nand ginst7088 (P1_U6360, P1_GTE_485_U6, P1_U4204);
  nand ginst7089 (P1_U6361, P1_R2167_U17, P1_U4202);
  nand ginst7090 (P1_U6362, P1_U3263, P1_U4203);
  not ginst7091 (P1_U6363, P1_U3431);
  nand ginst7092 (P1_U6364, P1_STATE2_REG_2__SCAN_IN, P1_U4249);
  nand ginst7093 (P1_U6365, P1_STATE2_REG_1__SCAN_IN, P1_R2337_U69);
  nand ginst7094 (P1_U6366, P1_U6364, P1_U6365);
  or ginst7095 (P1_U6367, P1_STATEBS16_REG_SCAN_IN, U210);
  nand ginst7096 (P1_U6368, P1_R2099_U86, P1_U2604);
  nand ginst7097 (P1_U6369, P1_REIP_REG_0__SCAN_IN, P1_U7485);
  nand ginst7098 (P1_U6370, P1_EBX_REG_0__SCAN_IN, P1_U7484);
  nand ginst7099 (P1_U6371, P1_R2358_U76, P1_U2429);
  nand ginst7100 (P1_U6372, P1_R2182_U34, P1_U2426);
  nand ginst7101 (P1_U6373, P1_PHYADDRPOINTER_REG_0__SCAN_IN, P1_U2373);
  nand ginst7102 (P1_U6374, P1_PHYADDRPOINTER_REG_0__SCAN_IN, P1_U2366);
  nand ginst7103 (P1_U6375, P1_REIP_REG_0__SCAN_IN, P1_U6363);
  nand ginst7104 (P1_U6376, P1_R2099_U87, P1_U2604);
  nand ginst7105 (P1_U6377, P1_R2096_U4, P1_U7485);
  nand ginst7106 (P1_U6378, P1_EBX_REG_1__SCAN_IN, P1_U7484);
  nand ginst7107 (P1_U6379, P1_R2358_U107, P1_U2429);
  nand ginst7108 (P1_U6380, P1_R2182_U33, P1_U2426);
  nand ginst7109 (P1_U6381, P1_PHYADDRPOINTER_REG_1__SCAN_IN, P1_U2373);
  nand ginst7110 (P1_U6382, P1_R2337_U4, P1_U2366);
  nand ginst7111 (P1_U6383, P1_REIP_REG_1__SCAN_IN, P1_U6363);
  nand ginst7112 (P1_U6384, P1_R2099_U138, P1_U2604);
  nand ginst7113 (P1_U6385, P1_R2096_U71, P1_U7485);
  nand ginst7114 (P1_U6386, P1_EBX_REG_2__SCAN_IN, P1_U7484);
  nand ginst7115 (P1_U6387, P1_R2358_U18, P1_U2429);
  nand ginst7116 (P1_U6388, P1_R2182_U42, P1_U2426);
  nand ginst7117 (P1_U6389, P1_PHYADDRPOINTER_REG_2__SCAN_IN, P1_U2373);
  nand ginst7118 (P1_U6390, P1_R2337_U71, P1_U2366);
  nand ginst7119 (P1_U6391, P1_REIP_REG_2__SCAN_IN, P1_U6363);
  nand ginst7120 (P1_U6392, P1_R2099_U42, P1_U2604);
  nand ginst7121 (P1_U6393, P1_R2096_U68, P1_U7485);
  nand ginst7122 (P1_U6394, P1_EBX_REG_3__SCAN_IN, P1_U7484);
  nand ginst7123 (P1_U6395, P1_R2358_U19, P1_U2429);
  nand ginst7124 (P1_U6396, P1_R2182_U25, P1_U2426);
  nand ginst7125 (P1_U6397, P1_PHYADDRPOINTER_REG_3__SCAN_IN, P1_U2373);
  nand ginst7126 (P1_U6398, P1_R2337_U68, P1_U2366);
  nand ginst7127 (P1_U6399, P1_REIP_REG_3__SCAN_IN, P1_U6363);
  nand ginst7128 (P1_U6400, P1_R2099_U41, P1_U2604);
  nand ginst7129 (P1_U6401, P1_R2096_U67, P1_U7485);
  nand ginst7130 (P1_U6402, P1_EBX_REG_4__SCAN_IN, P1_U7484);
  nand ginst7131 (P1_U6403, P1_R2358_U84, P1_U2429);
  nand ginst7132 (P1_U6404, P1_R2182_U24, P1_U2426);
  nand ginst7133 (P1_U6405, P1_PHYADDRPOINTER_REG_4__SCAN_IN, P1_U2373);
  nand ginst7134 (P1_U6406, P1_R2337_U67, P1_U2366);
  nand ginst7135 (P1_U6407, P1_REIP_REG_4__SCAN_IN, P1_U6363);
  nand ginst7136 (P1_U6408, P1_R2099_U40, P1_U2604);
  nand ginst7137 (P1_U6409, P1_R2096_U66, P1_U7485);
  nand ginst7138 (P1_U6410, P1_EBX_REG_5__SCAN_IN, P1_U7484);
  nand ginst7139 (P1_U6411, P1_R2358_U82, P1_U2429);
  nand ginst7140 (P1_U6412, P1_R2182_U5, P1_U2426);
  nand ginst7141 (P1_U6413, P1_PHYADDRPOINTER_REG_5__SCAN_IN, P1_U2373);
  nand ginst7142 (P1_U6414, P1_R2337_U66, P1_U2366);
  nand ginst7143 (P1_U6415, P1_REIP_REG_5__SCAN_IN, P1_U6363);
  nand ginst7144 (P1_U6416, P1_R2099_U39, P1_U2604);
  nand ginst7145 (P1_U6417, P1_R2096_U65, P1_U7485);
  nand ginst7146 (P1_U6418, P1_EBX_REG_6__SCAN_IN, P1_U7484);
  nand ginst7147 (P1_U6419, P1_PHYADDRPOINTER_REG_6__SCAN_IN, P1_U2373);
  nand ginst7148 (P1_U6420, P1_R2358_U20, P1_U2367);
  nand ginst7149 (P1_U6421, P1_R2337_U65, P1_U2366);
  nand ginst7150 (P1_U6422, P1_REIP_REG_6__SCAN_IN, P1_U6363);
  nand ginst7151 (P1_U6423, P1_R2099_U38, P1_U2604);
  nand ginst7152 (P1_U6424, P1_R2096_U64, P1_U7485);
  nand ginst7153 (P1_U6425, P1_EBX_REG_7__SCAN_IN, P1_U7484);
  nand ginst7154 (P1_U6426, P1_PHYADDRPOINTER_REG_7__SCAN_IN, P1_U2373);
  nand ginst7155 (P1_U6427, P1_R2358_U21, P1_U2367);
  nand ginst7156 (P1_U6428, P1_R2337_U64, P1_U2366);
  nand ginst7157 (P1_U6429, P1_REIP_REG_7__SCAN_IN, P1_U6363);
  nand ginst7158 (P1_U6430, P1_R2099_U37, P1_U2604);
  nand ginst7159 (P1_U6431, P1_R2096_U63, P1_U7485);
  nand ginst7160 (P1_U6432, P1_EBX_REG_8__SCAN_IN, P1_U7484);
  nand ginst7161 (P1_U6433, P1_PHYADDRPOINTER_REG_8__SCAN_IN, P1_U2373);
  nand ginst7162 (P1_U6434, P1_R2358_U80, P1_U2367);
  nand ginst7163 (P1_U6435, P1_R2337_U63, P1_U2366);
  nand ginst7164 (P1_U6436, P1_REIP_REG_8__SCAN_IN, P1_U6363);
  nand ginst7165 (P1_U6437, P1_R2099_U36, P1_U2604);
  nand ginst7166 (P1_U6438, P1_R2096_U62, P1_U7485);
  nand ginst7167 (P1_U6439, P1_EBX_REG_9__SCAN_IN, P1_U7484);
  nand ginst7168 (P1_U6440, P1_PHYADDRPOINTER_REG_9__SCAN_IN, P1_U2373);
  nand ginst7169 (P1_U6441, P1_R2358_U78, P1_U2367);
  nand ginst7170 (P1_U6442, P1_R2337_U62, P1_U2366);
  nand ginst7171 (P1_U6443, P1_REIP_REG_9__SCAN_IN, P1_U6363);
  nand ginst7172 (P1_U6444, P1_R2099_U85, P1_U2604);
  nand ginst7173 (P1_U6445, P1_R2096_U91, P1_U7485);
  nand ginst7174 (P1_U6446, P1_EBX_REG_10__SCAN_IN, P1_U7484);
  nand ginst7175 (P1_U6447, P1_PHYADDRPOINTER_REG_10__SCAN_IN, P1_U2373);
  nand ginst7176 (P1_U6448, P1_R2358_U14, P1_U2367);
  nand ginst7177 (P1_U6449, P1_R2337_U91, P1_U2366);
  nand ginst7178 (P1_U6450, P1_REIP_REG_10__SCAN_IN, P1_U6363);
  nand ginst7179 (P1_U6451, P1_R2099_U84, P1_U2604);
  nand ginst7180 (P1_U6452, P1_R2096_U90, P1_U7485);
  nand ginst7181 (P1_U6453, P1_EBX_REG_11__SCAN_IN, P1_U7484);
  nand ginst7182 (P1_U6454, P1_PHYADDRPOINTER_REG_11__SCAN_IN, P1_U2373);
  nand ginst7183 (P1_U6455, P1_R2358_U15, P1_U2367);
  nand ginst7184 (P1_U6456, P1_R2337_U90, P1_U2366);
  nand ginst7185 (P1_U6457, P1_REIP_REG_11__SCAN_IN, P1_U6363);
  nand ginst7186 (P1_U6458, P1_R2099_U83, P1_U2604);
  nand ginst7187 (P1_U6459, P1_R2096_U89, P1_U7485);
  nand ginst7188 (P1_U6460, P1_EBX_REG_12__SCAN_IN, P1_U7484);
  nand ginst7189 (P1_U6461, P1_PHYADDRPOINTER_REG_12__SCAN_IN, P1_U2373);
  nand ginst7190 (P1_U6462, P1_R2358_U119, P1_U2367);
  nand ginst7191 (P1_U6463, P1_R2337_U89, P1_U2366);
  nand ginst7192 (P1_U6464, P1_REIP_REG_12__SCAN_IN, P1_U6363);
  nand ginst7193 (P1_U6465, P1_R2099_U82, P1_U2604);
  nand ginst7194 (P1_U6466, P1_R2096_U88, P1_U7485);
  nand ginst7195 (P1_U6467, P1_EBX_REG_13__SCAN_IN, P1_U7484);
  nand ginst7196 (P1_U6468, P1_PHYADDRPOINTER_REG_13__SCAN_IN, P1_U2373);
  nand ginst7197 (P1_U6469, P1_R2358_U117, P1_U2367);
  nand ginst7198 (P1_U6470, P1_R2337_U88, P1_U2366);
  nand ginst7199 (P1_U6471, P1_REIP_REG_13__SCAN_IN, P1_U6363);
  nand ginst7200 (P1_U6472, P1_R2099_U81, P1_U2604);
  nand ginst7201 (P1_U6473, P1_R2096_U87, P1_U7485);
  nand ginst7202 (P1_U6474, P1_EBX_REG_14__SCAN_IN, P1_U7484);
  nand ginst7203 (P1_U6475, P1_PHYADDRPOINTER_REG_14__SCAN_IN, P1_U2373);
  nand ginst7204 (P1_U6476, P1_R2358_U16, P1_U2367);
  nand ginst7205 (P1_U6477, P1_R2337_U87, P1_U2366);
  nand ginst7206 (P1_U6478, P1_REIP_REG_14__SCAN_IN, P1_U6363);
  nand ginst7207 (P1_U6479, P1_R2099_U80, P1_U2604);
  nand ginst7208 (P1_U6480, P1_R2096_U86, P1_U7485);
  nand ginst7209 (P1_U6481, P1_EBX_REG_15__SCAN_IN, P1_U7484);
  nand ginst7210 (P1_U6482, P1_PHYADDRPOINTER_REG_15__SCAN_IN, P1_U2373);
  nand ginst7211 (P1_U6483, P1_R2358_U17, P1_U2367);
  nand ginst7212 (P1_U6484, P1_R2337_U86, P1_U2366);
  nand ginst7213 (P1_U6485, P1_REIP_REG_15__SCAN_IN, P1_U6363);
  nand ginst7214 (P1_U6486, P1_R2099_U79, P1_U2604);
  nand ginst7215 (P1_U6487, P1_R2096_U85, P1_U7485);
  nand ginst7216 (P1_U6488, P1_EBX_REG_16__SCAN_IN, P1_U7484);
  nand ginst7217 (P1_U6489, P1_PHYADDRPOINTER_REG_16__SCAN_IN, P1_U2373);
  nand ginst7218 (P1_U6490, P1_R2358_U115, P1_U2367);
  nand ginst7219 (P1_U6491, P1_R2337_U85, P1_U2366);
  nand ginst7220 (P1_U6492, P1_REIP_REG_16__SCAN_IN, P1_U6363);
  nand ginst7221 (P1_U6493, P1_R2099_U78, P1_U2604);
  nand ginst7222 (P1_U6494, P1_R2096_U84, P1_U7485);
  nand ginst7223 (P1_U6495, P1_EBX_REG_17__SCAN_IN, P1_U7484);
  nand ginst7224 (P1_U6496, P1_PHYADDRPOINTER_REG_17__SCAN_IN, P1_U2373);
  nand ginst7225 (P1_U6497, P1_R2358_U113, P1_U2367);
  nand ginst7226 (P1_U6498, P1_R2337_U84, P1_U2366);
  nand ginst7227 (P1_U6499, P1_REIP_REG_17__SCAN_IN, P1_U6363);
  nand ginst7228 (P1_U6500, P1_R2099_U77, P1_U2604);
  nand ginst7229 (P1_U6501, P1_R2096_U83, P1_U7485);
  nand ginst7230 (P1_U6502, P1_EBX_REG_18__SCAN_IN, P1_U7484);
  nand ginst7231 (P1_U6503, P1_PHYADDRPOINTER_REG_18__SCAN_IN, P1_U2373);
  nand ginst7232 (P1_U6504, P1_R2358_U111, P1_U2367);
  nand ginst7233 (P1_U6505, P1_R2337_U83, P1_U2366);
  nand ginst7234 (P1_U6506, P1_REIP_REG_18__SCAN_IN, P1_U6363);
  nand ginst7235 (P1_U6507, P1_R2099_U76, P1_U2604);
  nand ginst7236 (P1_U6508, P1_R2096_U82, P1_U7485);
  nand ginst7237 (P1_U6509, P1_EBX_REG_19__SCAN_IN, P1_U7484);
  nand ginst7238 (P1_U6510, P1_PHYADDRPOINTER_REG_19__SCAN_IN, P1_U2373);
  nand ginst7239 (P1_U6511, P1_R2358_U109, P1_U2367);
  nand ginst7240 (P1_U6512, P1_R2337_U82, P1_U2366);
  nand ginst7241 (P1_U6513, P1_REIP_REG_19__SCAN_IN, P1_U6363);
  nand ginst7242 (P1_U6514, P1_R2099_U75, P1_U2604);
  nand ginst7243 (P1_U6515, P1_R2096_U81, P1_U7485);
  nand ginst7244 (P1_U6516, P1_EBX_REG_20__SCAN_IN, P1_U7484);
  nand ginst7245 (P1_U6517, P1_PHYADDRPOINTER_REG_20__SCAN_IN, P1_U2373);
  nand ginst7246 (P1_U6518, P1_R2358_U105, P1_U2367);
  nand ginst7247 (P1_U6519, P1_R2337_U81, P1_U2366);
  nand ginst7248 (P1_U6520, P1_REIP_REG_20__SCAN_IN, P1_U6363);
  nand ginst7249 (P1_U6521, P1_R2099_U74, P1_U2604);
  nand ginst7250 (P1_U6522, P1_R2096_U80, P1_U7485);
  nand ginst7251 (P1_U6523, P1_EBX_REG_21__SCAN_IN, P1_U7484);
  nand ginst7252 (P1_U6524, P1_PHYADDRPOINTER_REG_21__SCAN_IN, P1_U2373);
  nand ginst7253 (P1_U6525, P1_R2358_U103, P1_U2367);
  nand ginst7254 (P1_U6526, P1_R2337_U80, P1_U2366);
  nand ginst7255 (P1_U6527, P1_REIP_REG_21__SCAN_IN, P1_U6363);
  nand ginst7256 (P1_U6528, P1_R2099_U73, P1_U2604);
  nand ginst7257 (P1_U6529, P1_R2096_U79, P1_U7485);
  nand ginst7258 (P1_U6530, P1_EBX_REG_22__SCAN_IN, P1_U7484);
  nand ginst7259 (P1_U6531, P1_PHYADDRPOINTER_REG_22__SCAN_IN, P1_U2373);
  nand ginst7260 (P1_U6532, P1_R2358_U101, P1_U2367);
  nand ginst7261 (P1_U6533, P1_R2337_U79, P1_U2366);
  nand ginst7262 (P1_U6534, P1_REIP_REG_22__SCAN_IN, P1_U6363);
  nand ginst7263 (P1_U6535, P1_R2099_U72, P1_U2604);
  nand ginst7264 (P1_U6536, P1_R2096_U78, P1_U7485);
  nand ginst7265 (P1_U6537, P1_EBX_REG_23__SCAN_IN, P1_U7484);
  nand ginst7266 (P1_U6538, P1_PHYADDRPOINTER_REG_23__SCAN_IN, P1_U2373);
  nand ginst7267 (P1_U6539, P1_R2358_U99, P1_U2367);
  nand ginst7268 (P1_U6540, P1_R2337_U78, P1_U2366);
  nand ginst7269 (P1_U6541, P1_REIP_REG_23__SCAN_IN, P1_U6363);
  nand ginst7270 (P1_U6542, P1_R2099_U71, P1_U2604);
  nand ginst7271 (P1_U6543, P1_R2096_U77, P1_U7485);
  nand ginst7272 (P1_U6544, P1_EBX_REG_24__SCAN_IN, P1_U7484);
  nand ginst7273 (P1_U6545, P1_PHYADDRPOINTER_REG_24__SCAN_IN, P1_U2373);
  nand ginst7274 (P1_U6546, P1_R2358_U97, P1_U2367);
  nand ginst7275 (P1_U6547, P1_R2337_U77, P1_U2366);
  nand ginst7276 (P1_U6548, P1_REIP_REG_24__SCAN_IN, P1_U6363);
  nand ginst7277 (P1_U6549, P1_R2099_U70, P1_U2604);
  nand ginst7278 (P1_U6550, P1_R2096_U76, P1_U7485);
  nand ginst7279 (P1_U6551, P1_EBX_REG_25__SCAN_IN, P1_U7484);
  nand ginst7280 (P1_U6552, P1_PHYADDRPOINTER_REG_25__SCAN_IN, P1_U2373);
  nand ginst7281 (P1_U6553, P1_R2358_U95, P1_U2367);
  nand ginst7282 (P1_U6554, P1_R2337_U76, P1_U2366);
  nand ginst7283 (P1_U6555, P1_REIP_REG_25__SCAN_IN, P1_U6363);
  nand ginst7284 (P1_U6556, P1_R2099_U69, P1_U2604);
  nand ginst7285 (P1_U6557, P1_R2096_U75, P1_U7485);
  nand ginst7286 (P1_U6558, P1_EBX_REG_26__SCAN_IN, P1_U7484);
  nand ginst7287 (P1_U6559, P1_PHYADDRPOINTER_REG_26__SCAN_IN, P1_U2373);
  nand ginst7288 (P1_U6560, P1_R2358_U93, P1_U2367);
  nand ginst7289 (P1_U6561, P1_R2337_U75, P1_U2366);
  nand ginst7290 (P1_U6562, P1_REIP_REG_26__SCAN_IN, P1_U6363);
  nand ginst7291 (P1_U6563, P1_R2099_U68, P1_U2604);
  nand ginst7292 (P1_U6564, P1_R2096_U74, P1_U7485);
  nand ginst7293 (P1_U6565, P1_EBX_REG_27__SCAN_IN, P1_U7484);
  nand ginst7294 (P1_U6566, P1_PHYADDRPOINTER_REG_27__SCAN_IN, P1_U2373);
  nand ginst7295 (P1_U6567, P1_R2358_U91, P1_U2367);
  nand ginst7296 (P1_U6568, P1_R2337_U74, P1_U2366);
  nand ginst7297 (P1_U6569, P1_REIP_REG_27__SCAN_IN, P1_U6363);
  nand ginst7298 (P1_U6570, P1_R2099_U67, P1_U2604);
  nand ginst7299 (P1_U6571, P1_R2096_U73, P1_U7485);
  nand ginst7300 (P1_U6572, P1_EBX_REG_28__SCAN_IN, P1_U7484);
  nand ginst7301 (P1_U6573, P1_PHYADDRPOINTER_REG_28__SCAN_IN, P1_U2373);
  nand ginst7302 (P1_U6574, P1_R2358_U89, P1_U2367);
  nand ginst7303 (P1_U6575, P1_R2337_U73, P1_U2366);
  nand ginst7304 (P1_U6576, P1_REIP_REG_28__SCAN_IN, P1_U6363);
  nand ginst7305 (P1_U6577, P1_R2099_U66, P1_U2604);
  nand ginst7306 (P1_U6578, P1_R2096_U72, P1_U7485);
  nand ginst7307 (P1_U6579, P1_EBX_REG_29__SCAN_IN, P1_U7484);
  nand ginst7308 (P1_U6580, P1_PHYADDRPOINTER_REG_29__SCAN_IN, P1_U2373);
  nand ginst7309 (P1_U6581, P1_R2358_U87, P1_U2367);
  nand ginst7310 (P1_U6582, P1_R2337_U72, P1_U2366);
  nand ginst7311 (P1_U6583, P1_REIP_REG_29__SCAN_IN, P1_U6363);
  nand ginst7312 (P1_U6584, P1_R2099_U65, P1_U2604);
  nand ginst7313 (P1_U6585, P1_R2096_U70, P1_U7485);
  nand ginst7314 (P1_U6586, P1_EBX_REG_30__SCAN_IN, P1_U7484);
  nand ginst7315 (P1_U6587, P1_PHYADDRPOINTER_REG_30__SCAN_IN, P1_U2373);
  nand ginst7316 (P1_U6588, P1_R2358_U85, P1_U2367);
  nand ginst7317 (P1_U6589, P1_R2337_U70, P1_U2366);
  nand ginst7318 (P1_U6590, P1_REIP_REG_30__SCAN_IN, P1_U6363);
  nand ginst7319 (P1_U6591, P1_R2099_U64, P1_U2604);
  nand ginst7320 (P1_U6592, P1_R2096_U69, P1_U7485);
  nand ginst7321 (P1_U6593, P1_EBX_REG_31__SCAN_IN, P1_U7484);
  nand ginst7322 (P1_U6594, P1_PHYADDRPOINTER_REG_31__SCAN_IN, P1_U2373);
  nand ginst7323 (P1_U6595, P1_R2358_U22, P1_U2367);
  nand ginst7324 (P1_U6596, P1_R2337_U69, P1_U2366);
  nand ginst7325 (P1_U6597, P1_REIP_REG_31__SCAN_IN, P1_U6363);
  nand ginst7326 (P1_U6598, P1_DATAWIDTH_REG_0__SCAN_IN, P1_DATAWIDTH_REG_1__SCAN_IN);
  or ginst7327 (P1_U6599, P1_REIP_REG_1__SCAN_IN, P1_REIP_REG_0__SCAN_IN);
  not ginst7328 (P1_U6600, P1_U4177);
  nand ginst7329 (P1_U6601, P1_FLUSH_REG_SCAN_IN, P1_U4177);
  nand ginst7330 (P1_U6602, P1_U2428, P1_U3966);
  not ginst7331 (P1_U6603, P1_U4180);
  nand ginst7332 (P1_U6604, P1_STATEBS16_REG_SCAN_IN, P1_U4497);
  nand ginst7333 (P1_U6605, P1_U4208, P1_U6604);
  nand ginst7334 (P1_U6606, P1_U3964, P1_U6605);
  nand ginst7335 (P1_U6607, P1_STATE2_REG_0__SCAN_IN, P1_U6606);
  nand ginst7336 (P1_U6608, P1_U3272, P1_U4193);
  nand ginst7337 (P1_U6609, P1_U3965, P1_U6607);
  nand ginst7338 (P1_U6610, P1_U2368, P1_U2473);
  nand ginst7339 (P1_U6611, P1_CODEFETCH_REG_SCAN_IN, P1_U6610);
  nand ginst7340 (P1_U6612, P1_STATE2_REG_0__SCAN_IN, P1_U4255);
  nand ginst7341 (P1_U6613, P1_ADS_N_REG_SCAN_IN, P1_STATE_REG_0__SCAN_IN);
  not ginst7342 (P1_U6614, P1_U4181);
  nand ginst7343 (P1_U6615, P1_U3291, P1_U3968);
  nand ginst7344 (P1_U6616, P1_U3406, P1_U3969, P1_U4499);
  nand ginst7345 (P1_U6617, P1_MEMORYFETCH_REG_SCAN_IN, P1_U6616);
  nand ginst7346 (P1_U6618, P1_INSTQUEUE_REG_15__7__SCAN_IN, P1_U2544);
  nand ginst7347 (P1_U6619, P1_INSTQUEUE_REG_14__7__SCAN_IN, P1_U2543);
  nand ginst7348 (P1_U6620, P1_INSTQUEUE_REG_13__7__SCAN_IN, P1_U2542);
  nand ginst7349 (P1_U6621, P1_INSTQUEUE_REG_12__7__SCAN_IN, P1_U2541);
  nand ginst7350 (P1_U6622, P1_INSTQUEUE_REG_11__7__SCAN_IN, P1_U2539);
  nand ginst7351 (P1_U6623, P1_INSTQUEUE_REG_10__7__SCAN_IN, P1_U2538);
  nand ginst7352 (P1_U6624, P1_INSTQUEUE_REG_9__7__SCAN_IN, P1_U2537);
  nand ginst7353 (P1_U6625, P1_INSTQUEUE_REG_8__7__SCAN_IN, P1_U2536);
  nand ginst7354 (P1_U6626, P1_INSTQUEUE_REG_7__7__SCAN_IN, P1_U2534);
  nand ginst7355 (P1_U6627, P1_INSTQUEUE_REG_6__7__SCAN_IN, P1_U2533);
  nand ginst7356 (P1_U6628, P1_INSTQUEUE_REG_5__7__SCAN_IN, P1_U2532);
  nand ginst7357 (P1_U6629, P1_INSTQUEUE_REG_4__7__SCAN_IN, P1_U2531);
  nand ginst7358 (P1_U6630, P1_INSTQUEUE_REG_3__7__SCAN_IN, P1_U2529);
  nand ginst7359 (P1_U6631, P1_INSTQUEUE_REG_2__7__SCAN_IN, P1_U2527);
  nand ginst7360 (P1_U6632, P1_INSTQUEUE_REG_1__7__SCAN_IN, P1_U2525);
  nand ginst7361 (P1_U6633, P1_INSTQUEUE_REG_0__7__SCAN_IN, P1_U2523);
  nand ginst7362 (P1_U6634, P1_INSTQUEUE_REG_15__6__SCAN_IN, P1_U2544);
  nand ginst7363 (P1_U6635, P1_INSTQUEUE_REG_14__6__SCAN_IN, P1_U2543);
  nand ginst7364 (P1_U6636, P1_INSTQUEUE_REG_13__6__SCAN_IN, P1_U2542);
  nand ginst7365 (P1_U6637, P1_INSTQUEUE_REG_12__6__SCAN_IN, P1_U2541);
  nand ginst7366 (P1_U6638, P1_INSTQUEUE_REG_11__6__SCAN_IN, P1_U2539);
  nand ginst7367 (P1_U6639, P1_INSTQUEUE_REG_10__6__SCAN_IN, P1_U2538);
  nand ginst7368 (P1_U6640, P1_INSTQUEUE_REG_9__6__SCAN_IN, P1_U2537);
  nand ginst7369 (P1_U6641, P1_INSTQUEUE_REG_8__6__SCAN_IN, P1_U2536);
  nand ginst7370 (P1_U6642, P1_INSTQUEUE_REG_7__6__SCAN_IN, P1_U2534);
  nand ginst7371 (P1_U6643, P1_INSTQUEUE_REG_6__6__SCAN_IN, P1_U2533);
  nand ginst7372 (P1_U6644, P1_INSTQUEUE_REG_5__6__SCAN_IN, P1_U2532);
  nand ginst7373 (P1_U6645, P1_INSTQUEUE_REG_4__6__SCAN_IN, P1_U2531);
  nand ginst7374 (P1_U6646, P1_INSTQUEUE_REG_3__6__SCAN_IN, P1_U2529);
  nand ginst7375 (P1_U6647, P1_INSTQUEUE_REG_2__6__SCAN_IN, P1_U2527);
  nand ginst7376 (P1_U6648, P1_INSTQUEUE_REG_1__6__SCAN_IN, P1_U2525);
  nand ginst7377 (P1_U6649, P1_INSTQUEUE_REG_0__6__SCAN_IN, P1_U2523);
  nand ginst7378 (P1_U6650, P1_INSTQUEUE_REG_15__5__SCAN_IN, P1_U2544);
  nand ginst7379 (P1_U6651, P1_INSTQUEUE_REG_14__5__SCAN_IN, P1_U2543);
  nand ginst7380 (P1_U6652, P1_INSTQUEUE_REG_13__5__SCAN_IN, P1_U2542);
  nand ginst7381 (P1_U6653, P1_INSTQUEUE_REG_12__5__SCAN_IN, P1_U2541);
  nand ginst7382 (P1_U6654, P1_INSTQUEUE_REG_11__5__SCAN_IN, P1_U2539);
  nand ginst7383 (P1_U6655, P1_INSTQUEUE_REG_10__5__SCAN_IN, P1_U2538);
  nand ginst7384 (P1_U6656, P1_INSTQUEUE_REG_9__5__SCAN_IN, P1_U2537);
  nand ginst7385 (P1_U6657, P1_INSTQUEUE_REG_8__5__SCAN_IN, P1_U2536);
  nand ginst7386 (P1_U6658, P1_INSTQUEUE_REG_7__5__SCAN_IN, P1_U2534);
  nand ginst7387 (P1_U6659, P1_INSTQUEUE_REG_6__5__SCAN_IN, P1_U2533);
  nand ginst7388 (P1_U6660, P1_INSTQUEUE_REG_5__5__SCAN_IN, P1_U2532);
  nand ginst7389 (P1_U6661, P1_INSTQUEUE_REG_4__5__SCAN_IN, P1_U2531);
  nand ginst7390 (P1_U6662, P1_INSTQUEUE_REG_3__5__SCAN_IN, P1_U2529);
  nand ginst7391 (P1_U6663, P1_INSTQUEUE_REG_2__5__SCAN_IN, P1_U2527);
  nand ginst7392 (P1_U6664, P1_INSTQUEUE_REG_1__5__SCAN_IN, P1_U2525);
  nand ginst7393 (P1_U6665, P1_INSTQUEUE_REG_0__5__SCAN_IN, P1_U2523);
  nand ginst7394 (P1_U6666, P1_INSTQUEUE_REG_15__4__SCAN_IN, P1_U2544);
  nand ginst7395 (P1_U6667, P1_INSTQUEUE_REG_14__4__SCAN_IN, P1_U2543);
  nand ginst7396 (P1_U6668, P1_INSTQUEUE_REG_13__4__SCAN_IN, P1_U2542);
  nand ginst7397 (P1_U6669, P1_INSTQUEUE_REG_12__4__SCAN_IN, P1_U2541);
  nand ginst7398 (P1_U6670, P1_INSTQUEUE_REG_11__4__SCAN_IN, P1_U2539);
  nand ginst7399 (P1_U6671, P1_INSTQUEUE_REG_10__4__SCAN_IN, P1_U2538);
  nand ginst7400 (P1_U6672, P1_INSTQUEUE_REG_9__4__SCAN_IN, P1_U2537);
  nand ginst7401 (P1_U6673, P1_INSTQUEUE_REG_8__4__SCAN_IN, P1_U2536);
  nand ginst7402 (P1_U6674, P1_INSTQUEUE_REG_7__4__SCAN_IN, P1_U2534);
  nand ginst7403 (P1_U6675, P1_INSTQUEUE_REG_6__4__SCAN_IN, P1_U2533);
  nand ginst7404 (P1_U6676, P1_INSTQUEUE_REG_5__4__SCAN_IN, P1_U2532);
  nand ginst7405 (P1_U6677, P1_INSTQUEUE_REG_4__4__SCAN_IN, P1_U2531);
  nand ginst7406 (P1_U6678, P1_INSTQUEUE_REG_3__4__SCAN_IN, P1_U2529);
  nand ginst7407 (P1_U6679, P1_INSTQUEUE_REG_2__4__SCAN_IN, P1_U2527);
  nand ginst7408 (P1_U6680, P1_INSTQUEUE_REG_1__4__SCAN_IN, P1_U2525);
  nand ginst7409 (P1_U6681, P1_INSTQUEUE_REG_15__3__SCAN_IN, P1_U2544);
  nand ginst7410 (P1_U6682, P1_INSTQUEUE_REG_14__3__SCAN_IN, P1_U2543);
  nand ginst7411 (P1_U6683, P1_INSTQUEUE_REG_13__3__SCAN_IN, P1_U2542);
  nand ginst7412 (P1_U6684, P1_INSTQUEUE_REG_12__3__SCAN_IN, P1_U2541);
  nand ginst7413 (P1_U6685, P1_INSTQUEUE_REG_11__3__SCAN_IN, P1_U2539);
  nand ginst7414 (P1_U6686, P1_INSTQUEUE_REG_10__3__SCAN_IN, P1_U2538);
  nand ginst7415 (P1_U6687, P1_INSTQUEUE_REG_9__3__SCAN_IN, P1_U2537);
  nand ginst7416 (P1_U6688, P1_INSTQUEUE_REG_8__3__SCAN_IN, P1_U2536);
  nand ginst7417 (P1_U6689, P1_INSTQUEUE_REG_7__3__SCAN_IN, P1_U2534);
  nand ginst7418 (P1_U6690, P1_INSTQUEUE_REG_6__3__SCAN_IN, P1_U2533);
  nand ginst7419 (P1_U6691, P1_INSTQUEUE_REG_5__3__SCAN_IN, P1_U2532);
  nand ginst7420 (P1_U6692, P1_INSTQUEUE_REG_4__3__SCAN_IN, P1_U2531);
  nand ginst7421 (P1_U6693, P1_INSTQUEUE_REG_3__3__SCAN_IN, P1_U2529);
  nand ginst7422 (P1_U6694, P1_INSTQUEUE_REG_2__3__SCAN_IN, P1_U2527);
  nand ginst7423 (P1_U6695, P1_INSTQUEUE_REG_1__3__SCAN_IN, P1_U2525);
  nand ginst7424 (P1_U6696, P1_INSTQUEUE_REG_0__3__SCAN_IN, P1_U2523);
  nand ginst7425 (P1_U6697, P1_INSTQUEUE_REG_15__2__SCAN_IN, P1_U2544);
  nand ginst7426 (P1_U6698, P1_INSTQUEUE_REG_14__2__SCAN_IN, P1_U2543);
  nand ginst7427 (P1_U6699, P1_INSTQUEUE_REG_13__2__SCAN_IN, P1_U2542);
  nand ginst7428 (P1_U6700, P1_INSTQUEUE_REG_12__2__SCAN_IN, P1_U2541);
  nand ginst7429 (P1_U6701, P1_INSTQUEUE_REG_11__2__SCAN_IN, P1_U2539);
  nand ginst7430 (P1_U6702, P1_INSTQUEUE_REG_10__2__SCAN_IN, P1_U2538);
  nand ginst7431 (P1_U6703, P1_INSTQUEUE_REG_9__2__SCAN_IN, P1_U2537);
  nand ginst7432 (P1_U6704, P1_INSTQUEUE_REG_8__2__SCAN_IN, P1_U2536);
  nand ginst7433 (P1_U6705, P1_INSTQUEUE_REG_7__2__SCAN_IN, P1_U2534);
  nand ginst7434 (P1_U6706, P1_INSTQUEUE_REG_6__2__SCAN_IN, P1_U2533);
  nand ginst7435 (P1_U6707, P1_INSTQUEUE_REG_5__2__SCAN_IN, P1_U2532);
  nand ginst7436 (P1_U6708, P1_INSTQUEUE_REG_4__2__SCAN_IN, P1_U2531);
  nand ginst7437 (P1_U6709, P1_INSTQUEUE_REG_3__2__SCAN_IN, P1_U2529);
  nand ginst7438 (P1_U6710, P1_INSTQUEUE_REG_2__2__SCAN_IN, P1_U2527);
  nand ginst7439 (P1_U6711, P1_INSTQUEUE_REG_1__2__SCAN_IN, P1_U2525);
  nand ginst7440 (P1_U6712, P1_INSTQUEUE_REG_0__2__SCAN_IN, P1_U2523);
  nand ginst7441 (P1_U6713, P1_INSTQUEUE_REG_15__1__SCAN_IN, P1_U2544);
  nand ginst7442 (P1_U6714, P1_INSTQUEUE_REG_14__1__SCAN_IN, P1_U2543);
  nand ginst7443 (P1_U6715, P1_INSTQUEUE_REG_13__1__SCAN_IN, P1_U2542);
  nand ginst7444 (P1_U6716, P1_INSTQUEUE_REG_12__1__SCAN_IN, P1_U2541);
  nand ginst7445 (P1_U6717, P1_INSTQUEUE_REG_11__1__SCAN_IN, P1_U2539);
  nand ginst7446 (P1_U6718, P1_INSTQUEUE_REG_10__1__SCAN_IN, P1_U2538);
  nand ginst7447 (P1_U6719, P1_INSTQUEUE_REG_9__1__SCAN_IN, P1_U2537);
  nand ginst7448 (P1_U6720, P1_INSTQUEUE_REG_8__1__SCAN_IN, P1_U2536);
  nand ginst7449 (P1_U6721, P1_INSTQUEUE_REG_7__1__SCAN_IN, P1_U2534);
  nand ginst7450 (P1_U6722, P1_INSTQUEUE_REG_6__1__SCAN_IN, P1_U2533);
  nand ginst7451 (P1_U6723, P1_INSTQUEUE_REG_5__1__SCAN_IN, P1_U2532);
  nand ginst7452 (P1_U6724, P1_INSTQUEUE_REG_4__1__SCAN_IN, P1_U2531);
  nand ginst7453 (P1_U6725, P1_INSTQUEUE_REG_3__1__SCAN_IN, P1_U2529);
  nand ginst7454 (P1_U6726, P1_INSTQUEUE_REG_2__1__SCAN_IN, P1_U2527);
  nand ginst7455 (P1_U6727, P1_INSTQUEUE_REG_1__1__SCAN_IN, P1_U2525);
  nand ginst7456 (P1_U6728, P1_INSTQUEUE_REG_0__1__SCAN_IN, P1_U2523);
  nand ginst7457 (P1_U6729, P1_INSTQUEUE_REG_15__0__SCAN_IN, P1_U2544);
  nand ginst7458 (P1_U6730, P1_INSTQUEUE_REG_14__0__SCAN_IN, P1_U2543);
  nand ginst7459 (P1_U6731, P1_INSTQUEUE_REG_13__0__SCAN_IN, P1_U2542);
  nand ginst7460 (P1_U6732, P1_INSTQUEUE_REG_12__0__SCAN_IN, P1_U2541);
  nand ginst7461 (P1_U6733, P1_INSTQUEUE_REG_11__0__SCAN_IN, P1_U2539);
  nand ginst7462 (P1_U6734, P1_INSTQUEUE_REG_10__0__SCAN_IN, P1_U2538);
  nand ginst7463 (P1_U6735, P1_INSTQUEUE_REG_9__0__SCAN_IN, P1_U2537);
  nand ginst7464 (P1_U6736, P1_INSTQUEUE_REG_8__0__SCAN_IN, P1_U2536);
  nand ginst7465 (P1_U6737, P1_INSTQUEUE_REG_7__0__SCAN_IN, P1_U2534);
  nand ginst7466 (P1_U6738, P1_INSTQUEUE_REG_6__0__SCAN_IN, P1_U2533);
  nand ginst7467 (P1_U6739, P1_INSTQUEUE_REG_5__0__SCAN_IN, P1_U2532);
  nand ginst7468 (P1_U6740, P1_INSTQUEUE_REG_4__0__SCAN_IN, P1_U2531);
  nand ginst7469 (P1_U6741, P1_INSTQUEUE_REG_3__0__SCAN_IN, P1_U2529);
  nand ginst7470 (P1_U6742, P1_INSTQUEUE_REG_2__0__SCAN_IN, P1_U2527);
  nand ginst7471 (P1_U6743, P1_INSTQUEUE_REG_1__0__SCAN_IN, P1_U2525);
  nand ginst7472 (P1_U6744, P1_INSTQUEUE_REG_0__0__SCAN_IN, P1_U2523);
  nand ginst7473 (P1_U6745, P1_STATE2_REG_2__SCAN_IN, P1_U4460);
  nand ginst7474 (P1_U6746, P1_U3412, P1_U6745);
  nand ginst7475 (P1_U6747, P1_EAX_REG_9__SCAN_IN, P1_U4188);
  nand ginst7476 (P1_U6748, P1_PHYADDRPOINTER_REG_9__SCAN_IN, P1_U4187);
  nand ginst7477 (P1_U6749, P1_R2337_U62, P1_U2352);
  nand ginst7478 (P1_U6750, P1_EAX_REG_8__SCAN_IN, P1_U4188);
  nand ginst7479 (P1_U6751, P1_PHYADDRPOINTER_REG_8__SCAN_IN, P1_U4187);
  nand ginst7480 (P1_U6752, P1_R2337_U63, P1_U2352);
  nand ginst7481 (P1_U6753, P1_EAX_REG_7__SCAN_IN, P1_U4188);
  nand ginst7482 (P1_U6754, P1_PHYADDRPOINTER_REG_7__SCAN_IN, P1_U4187);
  nand ginst7483 (P1_U6755, P1_R2337_U64, P1_U2352);
  nand ginst7484 (P1_U6756, P1_EAX_REG_6__SCAN_IN, P1_U4188);
  nand ginst7485 (P1_U6757, P1_PHYADDRPOINTER_REG_6__SCAN_IN, P1_U4187);
  nand ginst7486 (P1_U6758, P1_R2337_U65, P1_U2352);
  nand ginst7487 (P1_U6759, P1_R2182_U5, P1_U6746);
  nand ginst7488 (P1_U6760, P1_EAX_REG_5__SCAN_IN, P1_U4188);
  nand ginst7489 (P1_U6761, P1_PHYADDRPOINTER_REG_5__SCAN_IN, P1_U4187);
  nand ginst7490 (P1_U6762, P1_R2337_U66, P1_U2352);
  nand ginst7491 (P1_U6763, P1_R2182_U24, P1_U6746);
  nand ginst7492 (P1_U6764, P1_EAX_REG_4__SCAN_IN, P1_U4188);
  nand ginst7493 (P1_U6765, P1_PHYADDRPOINTER_REG_4__SCAN_IN, P1_U4187);
  nand ginst7494 (P1_U6766, P1_R2337_U67, P1_U2352);
  nand ginst7495 (P1_U6767, P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN, P1_U2353);
  nand ginst7496 (P1_U6768, P1_EAX_REG_31__SCAN_IN, P1_U4188);
  nand ginst7497 (P1_U6769, P1_PHYADDRPOINTER_REG_31__SCAN_IN, P1_U4187);
  nand ginst7498 (P1_U6770, P1_R2337_U69, P1_U2352);
  nand ginst7499 (P1_U6771, P1_R2182_U26, P1_U6746);
  nand ginst7500 (P1_U6772, P1_EAX_REG_30__SCAN_IN, P1_U4188);
  nand ginst7501 (P1_U6773, P1_PHYADDRPOINTER_REG_30__SCAN_IN, P1_U4187);
  nand ginst7502 (P1_U6774, P1_R2337_U70, P1_U2352);
  nand ginst7503 (P1_U6775, P1_R2182_U25, P1_U6746);
  nand ginst7504 (P1_U6776, P1_EAX_REG_3__SCAN_IN, P1_U4188);
  nand ginst7505 (P1_U6777, P1_PHYADDRPOINTER_REG_3__SCAN_IN, P1_U4187);
  nand ginst7506 (P1_U6778, P1_R2337_U68, P1_U2352);
  nand ginst7507 (P1_U6779, P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P1_U2353);
  nand ginst7508 (P1_U6780, P1_R2182_U27, P1_U6746);
  nand ginst7509 (P1_U6781, P1_EAX_REG_29__SCAN_IN, P1_U4188);
  nand ginst7510 (P1_U6782, P1_PHYADDRPOINTER_REG_29__SCAN_IN, P1_U4187);
  nand ginst7511 (P1_U6783, P1_R2337_U72, P1_U2352);
  nand ginst7512 (P1_U6784, P1_R2182_U28, P1_U6746);
  nand ginst7513 (P1_U6785, P1_EAX_REG_28__SCAN_IN, P1_U4188);
  nand ginst7514 (P1_U6786, P1_PHYADDRPOINTER_REG_28__SCAN_IN, P1_U4187);
  nand ginst7515 (P1_U6787, P1_R2337_U73, P1_U2352);
  nand ginst7516 (P1_U6788, P1_R2182_U29, P1_U6746);
  nand ginst7517 (P1_U6789, P1_EAX_REG_27__SCAN_IN, P1_U4188);
  nand ginst7518 (P1_U6790, P1_PHYADDRPOINTER_REG_27__SCAN_IN, P1_U4187);
  nand ginst7519 (P1_U6791, P1_R2337_U74, P1_U2352);
  nand ginst7520 (P1_U6792, P1_R2182_U30, P1_U6746);
  nand ginst7521 (P1_U6793, P1_EAX_REG_26__SCAN_IN, P1_U4188);
  nand ginst7522 (P1_U6794, P1_PHYADDRPOINTER_REG_26__SCAN_IN, P1_U4187);
  nand ginst7523 (P1_U6795, P1_R2337_U75, P1_U2352);
  nand ginst7524 (P1_U6796, P1_R2182_U31, P1_U6746);
  nand ginst7525 (P1_U6797, P1_EAX_REG_25__SCAN_IN, P1_U4188);
  nand ginst7526 (P1_U6798, P1_PHYADDRPOINTER_REG_25__SCAN_IN, P1_U4187);
  nand ginst7527 (P1_U6799, P1_R2337_U76, P1_U2352);
  nand ginst7528 (P1_U6800, P1_R2182_U32, P1_U6746);
  nand ginst7529 (P1_U6801, P1_EAX_REG_24__SCAN_IN, P1_U4188);
  nand ginst7530 (P1_U6802, P1_PHYADDRPOINTER_REG_24__SCAN_IN, P1_U4187);
  nand ginst7531 (P1_U6803, P1_R2337_U77, P1_U2352);
  nand ginst7532 (P1_U6804, P1_R2182_U6, P1_U6746);
  nand ginst7533 (P1_U6805, P1_EAX_REG_23__SCAN_IN, P1_U4188);
  nand ginst7534 (P1_U6806, P1_PHYADDRPOINTER_REG_23__SCAN_IN, P1_U4187);
  nand ginst7535 (P1_U6807, P1_R2337_U78, P1_U2352);
  nand ginst7536 (P1_U6808, P1_U2724, P1_U6746);
  nand ginst7537 (P1_U6809, P1_EAX_REG_22__SCAN_IN, P1_U4188);
  nand ginst7538 (P1_U6810, P1_PHYADDRPOINTER_REG_22__SCAN_IN, P1_U4187);
  nand ginst7539 (P1_U6811, P1_R2337_U79, P1_U2352);
  nand ginst7540 (P1_U6812, P1_U2725, P1_U6746);
  nand ginst7541 (P1_U6813, P1_EAX_REG_21__SCAN_IN, P1_U4188);
  nand ginst7542 (P1_U6814, P1_PHYADDRPOINTER_REG_21__SCAN_IN, P1_U4187);
  nand ginst7543 (P1_U6815, P1_R2337_U80, P1_U2352);
  nand ginst7544 (P1_U6816, P1_U2726, P1_U6746);
  nand ginst7545 (P1_U6817, P1_EAX_REG_20__SCAN_IN, P1_U4188);
  nand ginst7546 (P1_U6818, P1_PHYADDRPOINTER_REG_20__SCAN_IN, P1_U4187);
  nand ginst7547 (P1_U6819, P1_R2337_U81, P1_U2352);
  nand ginst7548 (P1_U6820, P1_R2182_U42, P1_U6746);
  nand ginst7549 (P1_U6821, P1_EAX_REG_2__SCAN_IN, P1_U4188);
  nand ginst7550 (P1_U6822, P1_PHYADDRPOINTER_REG_2__SCAN_IN, P1_U4187);
  nand ginst7551 (P1_U6823, P1_R2337_U71, P1_U2352);
  nand ginst7552 (P1_U6824, P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN, P1_U2353);
  nand ginst7553 (P1_U6825, P1_U2727, P1_U6746);
  nand ginst7554 (P1_U6826, P1_EAX_REG_19__SCAN_IN, P1_U4188);
  nand ginst7555 (P1_U6827, P1_PHYADDRPOINTER_REG_19__SCAN_IN, P1_U4187);
  nand ginst7556 (P1_U6828, P1_R2337_U82, P1_U2352);
  nand ginst7557 (P1_U6829, P1_U2728, P1_U6746);
  nand ginst7558 (P1_U6830, P1_EAX_REG_18__SCAN_IN, P1_U4188);
  nand ginst7559 (P1_U6831, P1_PHYADDRPOINTER_REG_18__SCAN_IN, P1_U4187);
  nand ginst7560 (P1_U6832, P1_R2337_U83, P1_U2352);
  nand ginst7561 (P1_U6833, P1_U2729, P1_U6746);
  nand ginst7562 (P1_U6834, P1_EAX_REG_17__SCAN_IN, P1_U4188);
  nand ginst7563 (P1_U6835, P1_PHYADDRPOINTER_REG_17__SCAN_IN, P1_U4187);
  nand ginst7564 (P1_U6836, P1_R2337_U84, P1_U2352);
  nand ginst7565 (P1_U6837, P1_U2730, P1_U6746);
  nand ginst7566 (P1_U6838, P1_EAX_REG_16__SCAN_IN, P1_U4188);
  nand ginst7567 (P1_U6839, P1_PHYADDRPOINTER_REG_16__SCAN_IN, P1_U4187);
  nand ginst7568 (P1_U6840, P1_R2337_U85, P1_U2352);
  nand ginst7569 (P1_U6841, P1_EAX_REG_15__SCAN_IN, P1_U4188);
  nand ginst7570 (P1_U6842, P1_PHYADDRPOINTER_REG_15__SCAN_IN, P1_U4187);
  nand ginst7571 (P1_U6843, P1_R2337_U86, P1_U2352);
  nand ginst7572 (P1_U6844, P1_EAX_REG_14__SCAN_IN, P1_U4188);
  nand ginst7573 (P1_U6845, P1_PHYADDRPOINTER_REG_14__SCAN_IN, P1_U4187);
  nand ginst7574 (P1_U6846, P1_R2337_U87, P1_U2352);
  nand ginst7575 (P1_U6847, P1_EAX_REG_13__SCAN_IN, P1_U4188);
  nand ginst7576 (P1_U6848, P1_PHYADDRPOINTER_REG_13__SCAN_IN, P1_U4187);
  nand ginst7577 (P1_U6849, P1_R2337_U88, P1_U2352);
  nand ginst7578 (P1_U6850, P1_EAX_REG_12__SCAN_IN, P1_U4188);
  nand ginst7579 (P1_U6851, P1_PHYADDRPOINTER_REG_12__SCAN_IN, P1_U4187);
  nand ginst7580 (P1_U6852, P1_R2337_U89, P1_U2352);
  nand ginst7581 (P1_U6853, P1_EAX_REG_11__SCAN_IN, P1_U4188);
  nand ginst7582 (P1_U6854, P1_PHYADDRPOINTER_REG_11__SCAN_IN, P1_U4187);
  nand ginst7583 (P1_U6855, P1_R2337_U90, P1_U2352);
  nand ginst7584 (P1_U6856, P1_EAX_REG_10__SCAN_IN, P1_U4188);
  nand ginst7585 (P1_U6857, P1_PHYADDRPOINTER_REG_10__SCAN_IN, P1_U4187);
  nand ginst7586 (P1_U6858, P1_R2337_U91, P1_U2352);
  nand ginst7587 (P1_U6859, P1_R2182_U33, P1_U6746);
  nand ginst7588 (P1_U6860, P1_EAX_REG_1__SCAN_IN, P1_U4188);
  nand ginst7589 (P1_U6861, P1_PHYADDRPOINTER_REG_1__SCAN_IN, P1_U4187);
  nand ginst7590 (P1_U6862, P1_R2337_U4, P1_U2352);
  nand ginst7591 (P1_U6863, P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P1_U2353);
  nand ginst7592 (P1_U6864, P1_R2182_U34, P1_U6746);
  nand ginst7593 (P1_U6865, P1_EAX_REG_0__SCAN_IN, P1_U4188);
  nand ginst7594 (P1_U6866, P1_PHYADDRPOINTER_REG_0__SCAN_IN, P1_U4187);
  nand ginst7595 (P1_U6867, P1_PHYADDRPOINTER_REG_0__SCAN_IN, P1_U2352);
  nand ginst7596 (P1_U6868, P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN, P1_U2353);
  nand ginst7597 (P1_U6869, P1_R2144_U49, P1_U6746);
  nand ginst7598 (P1_U6870, P1_U3309, P1_U3439, P1_U4460);
  nand ginst7599 (P1_U6871, P1_R2144_U80, P1_U4159);
  nand ginst7600 (P1_U6872, P1_ADD_371_U6, P1_U4208);
  nand ginst7601 (P1_U6873, P1_R2144_U10, P1_U4159);
  nand ginst7602 (P1_U6874, P1_ADD_371_U21, P1_U4208);
  nand ginst7603 (P1_U6875, P1_R2144_U9, P1_U4159);
  nand ginst7604 (P1_U6876, P1_ADD_371_U17, P1_U4208);
  nand ginst7605 (P1_U6877, P1_R2144_U45, P1_U4159);
  nand ginst7606 (P1_U6878, P1_ADD_371_U19, P1_U4208);
  nand ginst7607 (P1_U6879, P1_R2144_U47, P1_U4159);
  nand ginst7608 (P1_U6880, P1_ADD_371_U18, P1_U4208);
  nand ginst7609 (P1_U6881, P1_R2144_U8, P1_U4159);
  nand ginst7610 (P1_U6882, P1_ADD_371_U24, P1_U4208);
  nand ginst7611 (P1_U6883, P1_R2144_U49, P1_U4159);
  nand ginst7612 (P1_U6884, P1_ADD_371_U5, P1_U4208);
  nand ginst7613 (P1_U6885, P1_U3283, P1_U4494);
  nand ginst7614 (P1_U6886, P1_R2144_U50, P1_U4159);
  nand ginst7615 (P1_U6887, P1_ADD_371_U20, P1_U4208);
  nand ginst7616 (P1_U6888, P1_U2605, P1_U3284);
  nand ginst7617 (P1_U6889, P1_R2144_U43, P1_U4159);
  nand ginst7618 (P1_U6890, P1_ADD_371_U4, P1_U4208);
  nand ginst7619 (P1_U6891, P1_U3283, P1_U4494);
  nand ginst7620 (P1_U6892, P1_INSTQUEUE_REG_15__1__SCAN_IN, P1_U2564);
  nand ginst7621 (P1_U6893, P1_INSTQUEUE_REG_14__1__SCAN_IN, P1_U2563);
  nand ginst7622 (P1_U6894, P1_INSTQUEUE_REG_13__1__SCAN_IN, P1_U2562);
  nand ginst7623 (P1_U6895, P1_INSTQUEUE_REG_12__1__SCAN_IN, P1_U2561);
  nand ginst7624 (P1_U6896, P1_INSTQUEUE_REG_11__1__SCAN_IN, P1_U2559);
  nand ginst7625 (P1_U6897, P1_INSTQUEUE_REG_10__1__SCAN_IN, P1_U2558);
  nand ginst7626 (P1_U6898, P1_INSTQUEUE_REG_9__1__SCAN_IN, P1_U2557);
  nand ginst7627 (P1_U6899, P1_INSTQUEUE_REG_8__1__SCAN_IN, P1_U2556);
  nand ginst7628 (P1_U6900, P1_INSTQUEUE_REG_7__1__SCAN_IN, P1_U2554);
  nand ginst7629 (P1_U6901, P1_INSTQUEUE_REG_6__1__SCAN_IN, P1_U2553);
  nand ginst7630 (P1_U6902, P1_INSTQUEUE_REG_5__1__SCAN_IN, P1_U2552);
  nand ginst7631 (P1_U6903, P1_INSTQUEUE_REG_4__1__SCAN_IN, P1_U2551);
  nand ginst7632 (P1_U6904, P1_INSTQUEUE_REG_3__1__SCAN_IN, P1_U2549);
  nand ginst7633 (P1_U6905, P1_INSTQUEUE_REG_2__1__SCAN_IN, P1_U2548);
  nand ginst7634 (P1_U6906, P1_INSTQUEUE_REG_1__1__SCAN_IN, P1_U2547);
  nand ginst7635 (P1_U6907, P1_INSTQUEUE_REG_0__1__SCAN_IN, P1_U2546);
  nand ginst7636 (P1_U6908, P1_U4029, P1_U4030, P1_U4031, P1_U4032);
  nand ginst7637 (P1_U6909, P1_U3405, P1_U3418);
  nand ginst7638 (P1_U6910, P1_INSTQUEUE_REG_15__0__SCAN_IN, P1_U2564);
  nand ginst7639 (P1_U6911, P1_INSTQUEUE_REG_14__0__SCAN_IN, P1_U2563);
  nand ginst7640 (P1_U6912, P1_INSTQUEUE_REG_13__0__SCAN_IN, P1_U2562);
  nand ginst7641 (P1_U6913, P1_INSTQUEUE_REG_12__0__SCAN_IN, P1_U2561);
  nand ginst7642 (P1_U6914, P1_INSTQUEUE_REG_11__0__SCAN_IN, P1_U2559);
  nand ginst7643 (P1_U6915, P1_INSTQUEUE_REG_10__0__SCAN_IN, P1_U2558);
  nand ginst7644 (P1_U6916, P1_INSTQUEUE_REG_9__0__SCAN_IN, P1_U2557);
  nand ginst7645 (P1_U6917, P1_INSTQUEUE_REG_8__0__SCAN_IN, P1_U2556);
  nand ginst7646 (P1_U6918, P1_INSTQUEUE_REG_7__0__SCAN_IN, P1_U2554);
  nand ginst7647 (P1_U6919, P1_INSTQUEUE_REG_6__0__SCAN_IN, P1_U2553);
  nand ginst7648 (P1_U6920, P1_INSTQUEUE_REG_5__0__SCAN_IN, P1_U2552);
  nand ginst7649 (P1_U6921, P1_INSTQUEUE_REG_4__0__SCAN_IN, P1_U2551);
  nand ginst7650 (P1_U6922, P1_INSTQUEUE_REG_3__0__SCAN_IN, P1_U2549);
  nand ginst7651 (P1_U6923, P1_INSTQUEUE_REG_2__0__SCAN_IN, P1_U2548);
  nand ginst7652 (P1_U6924, P1_INSTQUEUE_REG_1__0__SCAN_IN, P1_U2547);
  nand ginst7653 (P1_U6925, P1_INSTQUEUE_REG_0__0__SCAN_IN, P1_U2546);
  nand ginst7654 (P1_U6926, P1_U4033, P1_U4034, P1_U4035, P1_U4036);
  nand ginst7655 (P1_U6927, P1_U3234, P1_U4207);
  nand ginst7656 (P1_U6928, P1_SUB_357_U8, P1_U2355);
  nand ginst7657 (P1_U6929, P1_U3233, P1_U4207);
  nand ginst7658 (P1_U6930, P1_SUB_357_U6, P1_U2355);
  nand ginst7659 (P1_U6931, P1_U3232, P1_U4207);
  nand ginst7660 (P1_U6932, P1_SUB_357_U9, P1_U2355);
  nand ginst7661 (P1_U6933, P1_U3231, P1_U4207);
  nand ginst7662 (P1_U6934, P1_SUB_357_U13, P1_U2355);
  nand ginst7663 (P1_U6935, P1_U3230, P1_U4207);
  nand ginst7664 (P1_U6936, P1_SUB_357_U11, P1_U2355);
  nand ginst7665 (P1_U6937, P1_R2182_U25, P1_U3294);
  nand ginst7666 (P1_U6938, P1_U3229, P1_U4207);
  nand ginst7667 (P1_U6939, P1_SUB_357_U12, P1_U2355);
  nand ginst7668 (P1_U6940, P1_R2182_U42, P1_U3294);
  nand ginst7669 (P1_U6941, P1_INSTQUEUE_REG_15__7__SCAN_IN, P1_U2564);
  nand ginst7670 (P1_U6942, P1_INSTQUEUE_REG_14__7__SCAN_IN, P1_U2563);
  nand ginst7671 (P1_U6943, P1_INSTQUEUE_REG_13__7__SCAN_IN, P1_U2562);
  nand ginst7672 (P1_U6944, P1_INSTQUEUE_REG_12__7__SCAN_IN, P1_U2561);
  nand ginst7673 (P1_U6945, P1_INSTQUEUE_REG_11__7__SCAN_IN, P1_U2559);
  nand ginst7674 (P1_U6946, P1_INSTQUEUE_REG_10__7__SCAN_IN, P1_U2558);
  nand ginst7675 (P1_U6947, P1_INSTQUEUE_REG_9__7__SCAN_IN, P1_U2557);
  nand ginst7676 (P1_U6948, P1_INSTQUEUE_REG_8__7__SCAN_IN, P1_U2556);
  nand ginst7677 (P1_U6949, P1_INSTQUEUE_REG_7__7__SCAN_IN, P1_U2554);
  nand ginst7678 (P1_U6950, P1_INSTQUEUE_REG_6__7__SCAN_IN, P1_U2553);
  nand ginst7679 (P1_U6951, P1_INSTQUEUE_REG_5__7__SCAN_IN, P1_U2552);
  nand ginst7680 (P1_U6952, P1_INSTQUEUE_REG_4__7__SCAN_IN, P1_U2551);
  nand ginst7681 (P1_U6953, P1_INSTQUEUE_REG_3__7__SCAN_IN, P1_U2549);
  nand ginst7682 (P1_U6954, P1_INSTQUEUE_REG_2__7__SCAN_IN, P1_U2548);
  nand ginst7683 (P1_U6955, P1_INSTQUEUE_REG_1__7__SCAN_IN, P1_U2547);
  nand ginst7684 (P1_U6956, P1_INSTQUEUE_REG_0__7__SCAN_IN, P1_U2546);
  nand ginst7685 (P1_U6957, P1_U4037, P1_U4038, P1_U4039, P1_U4040);
  nand ginst7686 (P1_U6958, P1_INSTQUEUE_REG_15__6__SCAN_IN, P1_U2564);
  nand ginst7687 (P1_U6959, P1_INSTQUEUE_REG_14__6__SCAN_IN, P1_U2563);
  nand ginst7688 (P1_U6960, P1_INSTQUEUE_REG_13__6__SCAN_IN, P1_U2562);
  nand ginst7689 (P1_U6961, P1_INSTQUEUE_REG_12__6__SCAN_IN, P1_U2561);
  nand ginst7690 (P1_U6962, P1_INSTQUEUE_REG_11__6__SCAN_IN, P1_U2559);
  nand ginst7691 (P1_U6963, P1_INSTQUEUE_REG_10__6__SCAN_IN, P1_U2558);
  nand ginst7692 (P1_U6964, P1_INSTQUEUE_REG_9__6__SCAN_IN, P1_U2557);
  nand ginst7693 (P1_U6965, P1_INSTQUEUE_REG_8__6__SCAN_IN, P1_U2556);
  nand ginst7694 (P1_U6966, P1_INSTQUEUE_REG_7__6__SCAN_IN, P1_U2554);
  nand ginst7695 (P1_U6967, P1_INSTQUEUE_REG_6__6__SCAN_IN, P1_U2553);
  nand ginst7696 (P1_U6968, P1_INSTQUEUE_REG_5__6__SCAN_IN, P1_U2552);
  nand ginst7697 (P1_U6969, P1_INSTQUEUE_REG_4__6__SCAN_IN, P1_U2551);
  nand ginst7698 (P1_U6970, P1_INSTQUEUE_REG_3__6__SCAN_IN, P1_U2549);
  nand ginst7699 (P1_U6971, P1_INSTQUEUE_REG_2__6__SCAN_IN, P1_U2548);
  nand ginst7700 (P1_U6972, P1_INSTQUEUE_REG_1__6__SCAN_IN, P1_U2547);
  nand ginst7701 (P1_U6973, P1_INSTQUEUE_REG_0__6__SCAN_IN, P1_U2546);
  nand ginst7702 (P1_U6974, P1_U4041, P1_U4042, P1_U4043, P1_U4044);
  nand ginst7703 (P1_U6975, P1_INSTQUEUE_REG_15__5__SCAN_IN, P1_U2564);
  nand ginst7704 (P1_U6976, P1_INSTQUEUE_REG_14__5__SCAN_IN, P1_U2563);
  nand ginst7705 (P1_U6977, P1_INSTQUEUE_REG_13__5__SCAN_IN, P1_U2562);
  nand ginst7706 (P1_U6978, P1_INSTQUEUE_REG_12__5__SCAN_IN, P1_U2561);
  nand ginst7707 (P1_U6979, P1_INSTQUEUE_REG_11__5__SCAN_IN, P1_U2559);
  nand ginst7708 (P1_U6980, P1_INSTQUEUE_REG_10__5__SCAN_IN, P1_U2558);
  nand ginst7709 (P1_U6981, P1_INSTQUEUE_REG_9__5__SCAN_IN, P1_U2557);
  nand ginst7710 (P1_U6982, P1_INSTQUEUE_REG_8__5__SCAN_IN, P1_U2556);
  nand ginst7711 (P1_U6983, P1_INSTQUEUE_REG_7__5__SCAN_IN, P1_U2554);
  nand ginst7712 (P1_U6984, P1_INSTQUEUE_REG_6__5__SCAN_IN, P1_U2553);
  nand ginst7713 (P1_U6985, P1_INSTQUEUE_REG_5__5__SCAN_IN, P1_U2552);
  nand ginst7714 (P1_U6986, P1_INSTQUEUE_REG_4__5__SCAN_IN, P1_U2551);
  nand ginst7715 (P1_U6987, P1_INSTQUEUE_REG_3__5__SCAN_IN, P1_U2549);
  nand ginst7716 (P1_U6988, P1_INSTQUEUE_REG_2__5__SCAN_IN, P1_U2548);
  nand ginst7717 (P1_U6989, P1_INSTQUEUE_REG_1__5__SCAN_IN, P1_U2547);
  nand ginst7718 (P1_U6990, P1_INSTQUEUE_REG_0__5__SCAN_IN, P1_U2546);
  nand ginst7719 (P1_U6991, P1_U4045, P1_U4046, P1_U4047, P1_U4048);
  nand ginst7720 (P1_U6992, P1_INSTQUEUE_REG_15__4__SCAN_IN, P1_U2564);
  nand ginst7721 (P1_U6993, P1_INSTQUEUE_REG_14__4__SCAN_IN, P1_U2563);
  nand ginst7722 (P1_U6994, P1_INSTQUEUE_REG_13__4__SCAN_IN, P1_U2562);
  nand ginst7723 (P1_U6995, P1_INSTQUEUE_REG_12__4__SCAN_IN, P1_U2561);
  nand ginst7724 (P1_U6996, P1_INSTQUEUE_REG_11__4__SCAN_IN, P1_U2559);
  nand ginst7725 (P1_U6997, P1_INSTQUEUE_REG_10__4__SCAN_IN, P1_U2558);
  nand ginst7726 (P1_U6998, P1_INSTQUEUE_REG_9__4__SCAN_IN, P1_U2557);
  nand ginst7727 (P1_U6999, P1_INSTQUEUE_REG_8__4__SCAN_IN, P1_U2556);
  nand ginst7728 (P1_U7000, P1_INSTQUEUE_REG_7__4__SCAN_IN, P1_U2554);
  nand ginst7729 (P1_U7001, P1_INSTQUEUE_REG_6__4__SCAN_IN, P1_U2553);
  nand ginst7730 (P1_U7002, P1_INSTQUEUE_REG_5__4__SCAN_IN, P1_U2552);
  nand ginst7731 (P1_U7003, P1_INSTQUEUE_REG_4__4__SCAN_IN, P1_U2551);
  nand ginst7732 (P1_U7004, P1_INSTQUEUE_REG_3__4__SCAN_IN, P1_U2549);
  nand ginst7733 (P1_U7005, P1_INSTQUEUE_REG_2__4__SCAN_IN, P1_U2548);
  nand ginst7734 (P1_U7006, P1_INSTQUEUE_REG_1__4__SCAN_IN, P1_U2547);
  nand ginst7735 (P1_U7007, P1_INSTQUEUE_REG_15__3__SCAN_IN, P1_U2564);
  nand ginst7736 (P1_U7008, P1_INSTQUEUE_REG_14__3__SCAN_IN, P1_U2563);
  nand ginst7737 (P1_U7009, P1_INSTQUEUE_REG_13__3__SCAN_IN, P1_U2562);
  nand ginst7738 (P1_U7010, P1_INSTQUEUE_REG_12__3__SCAN_IN, P1_U2561);
  nand ginst7739 (P1_U7011, P1_INSTQUEUE_REG_11__3__SCAN_IN, P1_U2559);
  nand ginst7740 (P1_U7012, P1_INSTQUEUE_REG_10__3__SCAN_IN, P1_U2558);
  nand ginst7741 (P1_U7013, P1_INSTQUEUE_REG_9__3__SCAN_IN, P1_U2557);
  nand ginst7742 (P1_U7014, P1_INSTQUEUE_REG_8__3__SCAN_IN, P1_U2556);
  nand ginst7743 (P1_U7015, P1_INSTQUEUE_REG_7__3__SCAN_IN, P1_U2554);
  nand ginst7744 (P1_U7016, P1_INSTQUEUE_REG_6__3__SCAN_IN, P1_U2553);
  nand ginst7745 (P1_U7017, P1_INSTQUEUE_REG_5__3__SCAN_IN, P1_U2552);
  nand ginst7746 (P1_U7018, P1_INSTQUEUE_REG_4__3__SCAN_IN, P1_U2551);
  nand ginst7747 (P1_U7019, P1_INSTQUEUE_REG_3__3__SCAN_IN, P1_U2549);
  nand ginst7748 (P1_U7020, P1_INSTQUEUE_REG_2__3__SCAN_IN, P1_U2548);
  nand ginst7749 (P1_U7021, P1_INSTQUEUE_REG_1__3__SCAN_IN, P1_U2547);
  nand ginst7750 (P1_U7022, P1_INSTQUEUE_REG_0__3__SCAN_IN, P1_U2546);
  nand ginst7751 (P1_U7023, P1_U4053, P1_U4054, P1_U4055, P1_U4056);
  nand ginst7752 (P1_U7024, P1_INSTQUEUE_REG_15__2__SCAN_IN, P1_U2564);
  nand ginst7753 (P1_U7025, P1_INSTQUEUE_REG_14__2__SCAN_IN, P1_U2563);
  nand ginst7754 (P1_U7026, P1_INSTQUEUE_REG_13__2__SCAN_IN, P1_U2562);
  nand ginst7755 (P1_U7027, P1_INSTQUEUE_REG_12__2__SCAN_IN, P1_U2561);
  nand ginst7756 (P1_U7028, P1_INSTQUEUE_REG_11__2__SCAN_IN, P1_U2559);
  nand ginst7757 (P1_U7029, P1_INSTQUEUE_REG_10__2__SCAN_IN, P1_U2558);
  nand ginst7758 (P1_U7030, P1_INSTQUEUE_REG_9__2__SCAN_IN, P1_U2557);
  nand ginst7759 (P1_U7031, P1_INSTQUEUE_REG_8__2__SCAN_IN, P1_U2556);
  nand ginst7760 (P1_U7032, P1_INSTQUEUE_REG_7__2__SCAN_IN, P1_U2554);
  nand ginst7761 (P1_U7033, P1_INSTQUEUE_REG_6__2__SCAN_IN, P1_U2553);
  nand ginst7762 (P1_U7034, P1_INSTQUEUE_REG_5__2__SCAN_IN, P1_U2552);
  nand ginst7763 (P1_U7035, P1_INSTQUEUE_REG_4__2__SCAN_IN, P1_U2551);
  nand ginst7764 (P1_U7036, P1_INSTQUEUE_REG_3__2__SCAN_IN, P1_U2549);
  nand ginst7765 (P1_U7037, P1_INSTQUEUE_REG_2__2__SCAN_IN, P1_U2548);
  nand ginst7766 (P1_U7038, P1_INSTQUEUE_REG_1__2__SCAN_IN, P1_U2547);
  nand ginst7767 (P1_U7039, P1_INSTQUEUE_REG_0__2__SCAN_IN, P1_U2546);
  nand ginst7768 (P1_U7040, P1_U4057, P1_U4058, P1_U4059, P1_U4060);
  nand ginst7769 (P1_U7041, P1_U3228, P1_U4207);
  nand ginst7770 (P1_U7042, P1_SUB_357_U7, P1_U2355);
  nand ginst7771 (P1_U7043, P1_R2182_U33, P1_U3294);
  nand ginst7772 (P1_U7044, P1_U3227, P1_U4207);
  nand ginst7773 (P1_U7045, P1_SUB_357_U10, P1_U2355);
  nand ginst7774 (P1_U7046, P1_R2182_U34, P1_U3294);
  nand ginst7775 (P1_U7047, P1_U3234, P1_U4206);
  nand ginst7776 (P1_U7048, P1_INSTQUEUE_REG_0__7__SCAN_IN, P1_U4192);
  nand ginst7777 (P1_U7049, P1_U3233, P1_U4206);
  nand ginst7778 (P1_U7050, P1_INSTQUEUE_REG_0__6__SCAN_IN, P1_U4192);
  nand ginst7779 (P1_U7051, P1_U3232, P1_U4206);
  nand ginst7780 (P1_U7052, P1_INSTQUEUE_REG_0__5__SCAN_IN, P1_U4192);
  nand ginst7781 (P1_U7053, P1_U3231, P1_U4206);
  nand ginst7782 (P1_U7054, P1_U3230, P1_U4206);
  nand ginst7783 (P1_U7055, P1_INSTQUEUE_REG_0__3__SCAN_IN, P1_U4192);
  nand ginst7784 (P1_U7056, P1_U3229, P1_U4206);
  nand ginst7785 (P1_U7057, P1_INSTQUEUE_REG_0__2__SCAN_IN, P1_U4192);
  nand ginst7786 (P1_U7058, P1_U3228, P1_U4206);
  nand ginst7787 (P1_U7059, P1_INSTQUEUE_REG_0__1__SCAN_IN, P1_U4192);
  nand ginst7788 (P1_U7060, P1_U3227, P1_U4206);
  nand ginst7789 (P1_U7061, P1_U3234, P1_U4400);
  nand ginst7790 (P1_U7062, P1_INSTQUEUE_REG_0__0__SCAN_IN, P1_U4192);
  nand ginst7791 (P1_U7063, P1_U3427, P1_U3428);
  nand ginst7792 (P1_U7064, P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P1_U3264);
  not ginst7793 (P1_U7065, P1_U3445);
  nand ginst7794 (P1_U7066, P1_INSTQUEUE_REG_8__7__SCAN_IN, P1_U2582);
  nand ginst7795 (P1_U7067, P1_INSTQUEUE_REG_9__7__SCAN_IN, P1_U2581);
  nand ginst7796 (P1_U7068, P1_INSTQUEUE_REG_10__7__SCAN_IN, P1_U2580);
  nand ginst7797 (P1_U7069, P1_INSTQUEUE_REG_11__7__SCAN_IN, P1_U2579);
  nand ginst7798 (P1_U7070, P1_INSTQUEUE_REG_12__7__SCAN_IN, P1_U2577);
  nand ginst7799 (P1_U7071, P1_INSTQUEUE_REG_13__7__SCAN_IN, P1_U2576);
  nand ginst7800 (P1_U7072, P1_INSTQUEUE_REG_14__7__SCAN_IN, P1_U2575);
  nand ginst7801 (P1_U7073, P1_INSTQUEUE_REG_15__7__SCAN_IN, P1_U2574);
  nand ginst7802 (P1_U7074, P1_INSTQUEUE_REG_0__7__SCAN_IN, P1_U2573);
  nand ginst7803 (P1_U7075, P1_INSTQUEUE_REG_1__7__SCAN_IN, P1_U2572);
  nand ginst7804 (P1_U7076, P1_INSTQUEUE_REG_2__7__SCAN_IN, P1_U2571);
  nand ginst7805 (P1_U7077, P1_INSTQUEUE_REG_3__7__SCAN_IN, P1_U2570);
  nand ginst7806 (P1_U7078, P1_INSTQUEUE_REG_4__7__SCAN_IN, P1_U2568);
  nand ginst7807 (P1_U7079, P1_INSTQUEUE_REG_5__7__SCAN_IN, P1_U2567);
  nand ginst7808 (P1_U7080, P1_INSTQUEUE_REG_6__7__SCAN_IN, P1_U2566);
  nand ginst7809 (P1_U7081, P1_INSTQUEUE_REG_7__7__SCAN_IN, P1_U2565);
  nand ginst7810 (P1_U7082, P1_U4063, P1_U4064, P1_U4065, P1_U4066);
  nand ginst7811 (P1_U7083, P1_U3421, P1_U3425);
  nand ginst7812 (P1_U7084, P1_U4073, P1_U4191);
  nand ginst7813 (P1_U7085, P1_U3422, P1_U7084);
  nand ginst7814 (P1_U7086, P1_U3278, P1_U4503);
  not ginst7815 (P1_U7087, P1_U3245);
  nand ginst7816 (P1_U7088, P1_U3394, P1_U4154, P1_U4400, P1_U4503);
  nand ginst7817 (P1_U7089, P1_STATE2_REG_0__SCAN_IN, P1_U4189);
  nand ginst7818 (P1_U7090, P1_U3245, P1_U4067);
  not ginst7819 (P1_U7091, P1_U3451);
  nand ginst7820 (P1_U7092, P1_U3451, P1_U5492, P1_U7629);
  nand ginst7821 (P1_U7093, P1_U4194, P1_U7092);
  not ginst7822 (P1_U7094, P1_U3450);
  nand ginst7823 (P1_U7095, P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN, P1_U3297);
  nand ginst7824 (P1_U7096, P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P1_U3450);
  nand ginst7825 (P1_U7097, P1_U3360, P1_U4203);
  nand ginst7826 (P1_U7098, P1_INSTQUEUE_REG_8__6__SCAN_IN, P1_U2582);
  nand ginst7827 (P1_U7099, P1_INSTQUEUE_REG_9__6__SCAN_IN, P1_U2581);
  nand ginst7828 (P1_U7100, P1_INSTQUEUE_REG_10__6__SCAN_IN, P1_U2580);
  nand ginst7829 (P1_U7101, P1_INSTQUEUE_REG_11__6__SCAN_IN, P1_U2579);
  nand ginst7830 (P1_U7102, P1_INSTQUEUE_REG_12__6__SCAN_IN, P1_U2577);
  nand ginst7831 (P1_U7103, P1_INSTQUEUE_REG_13__6__SCAN_IN, P1_U2576);
  nand ginst7832 (P1_U7104, P1_INSTQUEUE_REG_14__6__SCAN_IN, P1_U2575);
  nand ginst7833 (P1_U7105, P1_INSTQUEUE_REG_15__6__SCAN_IN, P1_U2574);
  nand ginst7834 (P1_U7106, P1_INSTQUEUE_REG_0__6__SCAN_IN, P1_U2573);
  nand ginst7835 (P1_U7107, P1_INSTQUEUE_REG_1__6__SCAN_IN, P1_U2572);
  nand ginst7836 (P1_U7108, P1_INSTQUEUE_REG_2__6__SCAN_IN, P1_U2571);
  nand ginst7837 (P1_U7109, P1_INSTQUEUE_REG_3__6__SCAN_IN, P1_U2570);
  nand ginst7838 (P1_U7110, P1_INSTQUEUE_REG_4__6__SCAN_IN, P1_U2568);
  nand ginst7839 (P1_U7111, P1_INSTQUEUE_REG_5__6__SCAN_IN, P1_U2567);
  nand ginst7840 (P1_U7112, P1_INSTQUEUE_REG_6__6__SCAN_IN, P1_U2566);
  nand ginst7841 (P1_U7113, P1_INSTQUEUE_REG_7__6__SCAN_IN, P1_U2565);
  nand ginst7842 (P1_U7114, P1_U4079, P1_U4080, P1_U4081, P1_U4082);
  nand ginst7843 (P1_U7115, P1_INSTQUEUE_REG_8__5__SCAN_IN, P1_U2582);
  nand ginst7844 (P1_U7116, P1_INSTQUEUE_REG_9__5__SCAN_IN, P1_U2581);
  nand ginst7845 (P1_U7117, P1_INSTQUEUE_REG_10__5__SCAN_IN, P1_U2580);
  nand ginst7846 (P1_U7118, P1_INSTQUEUE_REG_11__5__SCAN_IN, P1_U2579);
  nand ginst7847 (P1_U7119, P1_INSTQUEUE_REG_12__5__SCAN_IN, P1_U2577);
  nand ginst7848 (P1_U7120, P1_INSTQUEUE_REG_13__5__SCAN_IN, P1_U2576);
  nand ginst7849 (P1_U7121, P1_INSTQUEUE_REG_14__5__SCAN_IN, P1_U2575);
  nand ginst7850 (P1_U7122, P1_INSTQUEUE_REG_15__5__SCAN_IN, P1_U2574);
  nand ginst7851 (P1_U7123, P1_INSTQUEUE_REG_0__5__SCAN_IN, P1_U2573);
  nand ginst7852 (P1_U7124, P1_INSTQUEUE_REG_1__5__SCAN_IN, P1_U2572);
  nand ginst7853 (P1_U7125, P1_INSTQUEUE_REG_2__5__SCAN_IN, P1_U2571);
  nand ginst7854 (P1_U7126, P1_INSTQUEUE_REG_3__5__SCAN_IN, P1_U2570);
  nand ginst7855 (P1_U7127, P1_INSTQUEUE_REG_4__5__SCAN_IN, P1_U2568);
  nand ginst7856 (P1_U7128, P1_INSTQUEUE_REG_5__5__SCAN_IN, P1_U2567);
  nand ginst7857 (P1_U7129, P1_INSTQUEUE_REG_6__5__SCAN_IN, P1_U2566);
  nand ginst7858 (P1_U7130, P1_INSTQUEUE_REG_7__5__SCAN_IN, P1_U2565);
  nand ginst7859 (P1_U7131, P1_U4083, P1_U4084, P1_U4085, P1_U4086);
  nand ginst7860 (P1_U7132, P1_INSTQUEUE_REG_8__4__SCAN_IN, P1_U2582);
  nand ginst7861 (P1_U7133, P1_INSTQUEUE_REG_9__4__SCAN_IN, P1_U2581);
  nand ginst7862 (P1_U7134, P1_INSTQUEUE_REG_10__4__SCAN_IN, P1_U2580);
  nand ginst7863 (P1_U7135, P1_INSTQUEUE_REG_11__4__SCAN_IN, P1_U2579);
  nand ginst7864 (P1_U7136, P1_INSTQUEUE_REG_12__4__SCAN_IN, P1_U2577);
  nand ginst7865 (P1_U7137, P1_INSTQUEUE_REG_13__4__SCAN_IN, P1_U2576);
  nand ginst7866 (P1_U7138, P1_INSTQUEUE_REG_14__4__SCAN_IN, P1_U2575);
  nand ginst7867 (P1_U7139, P1_INSTQUEUE_REG_15__4__SCAN_IN, P1_U2574);
  nand ginst7868 (P1_U7140, P1_INSTQUEUE_REG_1__4__SCAN_IN, P1_U2572);
  nand ginst7869 (P1_U7141, P1_INSTQUEUE_REG_2__4__SCAN_IN, P1_U2571);
  nand ginst7870 (P1_U7142, P1_INSTQUEUE_REG_3__4__SCAN_IN, P1_U2570);
  nand ginst7871 (P1_U7143, P1_INSTQUEUE_REG_4__4__SCAN_IN, P1_U2568);
  nand ginst7872 (P1_U7144, P1_INSTQUEUE_REG_5__4__SCAN_IN, P1_U2567);
  nand ginst7873 (P1_U7145, P1_INSTQUEUE_REG_6__4__SCAN_IN, P1_U2566);
  nand ginst7874 (P1_U7146, P1_INSTQUEUE_REG_7__4__SCAN_IN, P1_U2565);
  nand ginst7875 (P1_U7147, P1_INSTQUEUE_REG_8__3__SCAN_IN, P1_U2582);
  nand ginst7876 (P1_U7148, P1_INSTQUEUE_REG_9__3__SCAN_IN, P1_U2581);
  nand ginst7877 (P1_U7149, P1_INSTQUEUE_REG_10__3__SCAN_IN, P1_U2580);
  nand ginst7878 (P1_U7150, P1_INSTQUEUE_REG_11__3__SCAN_IN, P1_U2579);
  nand ginst7879 (P1_U7151, P1_INSTQUEUE_REG_12__3__SCAN_IN, P1_U2577);
  nand ginst7880 (P1_U7152, P1_INSTQUEUE_REG_13__3__SCAN_IN, P1_U2576);
  nand ginst7881 (P1_U7153, P1_INSTQUEUE_REG_14__3__SCAN_IN, P1_U2575);
  nand ginst7882 (P1_U7154, P1_INSTQUEUE_REG_15__3__SCAN_IN, P1_U2574);
  nand ginst7883 (P1_U7155, P1_INSTQUEUE_REG_0__3__SCAN_IN, P1_U2573);
  nand ginst7884 (P1_U7156, P1_INSTQUEUE_REG_1__3__SCAN_IN, P1_U2572);
  nand ginst7885 (P1_U7157, P1_INSTQUEUE_REG_2__3__SCAN_IN, P1_U2571);
  nand ginst7886 (P1_U7158, P1_INSTQUEUE_REG_3__3__SCAN_IN, P1_U2570);
  nand ginst7887 (P1_U7159, P1_INSTQUEUE_REG_4__3__SCAN_IN, P1_U2568);
  nand ginst7888 (P1_U7160, P1_INSTQUEUE_REG_5__3__SCAN_IN, P1_U2567);
  nand ginst7889 (P1_U7161, P1_INSTQUEUE_REG_6__3__SCAN_IN, P1_U2566);
  nand ginst7890 (P1_U7162, P1_INSTQUEUE_REG_7__3__SCAN_IN, P1_U2565);
  nand ginst7891 (P1_U7163, P1_U4092, P1_U4093, P1_U4094, P1_U4095);
  nand ginst7892 (P1_U7164, P1_INSTQUEUE_REG_8__2__SCAN_IN, P1_U2582);
  nand ginst7893 (P1_U7165, P1_INSTQUEUE_REG_9__2__SCAN_IN, P1_U2581);
  nand ginst7894 (P1_U7166, P1_INSTQUEUE_REG_10__2__SCAN_IN, P1_U2580);
  nand ginst7895 (P1_U7167, P1_INSTQUEUE_REG_11__2__SCAN_IN, P1_U2579);
  nand ginst7896 (P1_U7168, P1_INSTQUEUE_REG_12__2__SCAN_IN, P1_U2577);
  nand ginst7897 (P1_U7169, P1_INSTQUEUE_REG_13__2__SCAN_IN, P1_U2576);
  nand ginst7898 (P1_U7170, P1_INSTQUEUE_REG_14__2__SCAN_IN, P1_U2575);
  nand ginst7899 (P1_U7171, P1_INSTQUEUE_REG_15__2__SCAN_IN, P1_U2574);
  nand ginst7900 (P1_U7172, P1_INSTQUEUE_REG_0__2__SCAN_IN, P1_U2573);
  nand ginst7901 (P1_U7173, P1_INSTQUEUE_REG_1__2__SCAN_IN, P1_U2572);
  nand ginst7902 (P1_U7174, P1_INSTQUEUE_REG_2__2__SCAN_IN, P1_U2571);
  nand ginst7903 (P1_U7175, P1_INSTQUEUE_REG_3__2__SCAN_IN, P1_U2570);
  nand ginst7904 (P1_U7176, P1_INSTQUEUE_REG_4__2__SCAN_IN, P1_U2568);
  nand ginst7905 (P1_U7177, P1_INSTQUEUE_REG_5__2__SCAN_IN, P1_U2567);
  nand ginst7906 (P1_U7178, P1_INSTQUEUE_REG_6__2__SCAN_IN, P1_U2566);
  nand ginst7907 (P1_U7179, P1_INSTQUEUE_REG_7__2__SCAN_IN, P1_U2565);
  nand ginst7908 (P1_U7180, P1_U4096, P1_U4097, P1_U4098, P1_U4099);
  nand ginst7909 (P1_U7181, P1_INSTQUEUE_REG_8__1__SCAN_IN, P1_U2582);
  nand ginst7910 (P1_U7182, P1_INSTQUEUE_REG_9__1__SCAN_IN, P1_U2581);
  nand ginst7911 (P1_U7183, P1_INSTQUEUE_REG_10__1__SCAN_IN, P1_U2580);
  nand ginst7912 (P1_U7184, P1_INSTQUEUE_REG_11__1__SCAN_IN, P1_U2579);
  nand ginst7913 (P1_U7185, P1_INSTQUEUE_REG_12__1__SCAN_IN, P1_U2577);
  nand ginst7914 (P1_U7186, P1_INSTQUEUE_REG_13__1__SCAN_IN, P1_U2576);
  nand ginst7915 (P1_U7187, P1_INSTQUEUE_REG_14__1__SCAN_IN, P1_U2575);
  nand ginst7916 (P1_U7188, P1_INSTQUEUE_REG_15__1__SCAN_IN, P1_U2574);
  nand ginst7917 (P1_U7189, P1_INSTQUEUE_REG_0__1__SCAN_IN, P1_U2573);
  nand ginst7918 (P1_U7190, P1_INSTQUEUE_REG_1__1__SCAN_IN, P1_U2572);
  nand ginst7919 (P1_U7191, P1_INSTQUEUE_REG_2__1__SCAN_IN, P1_U2571);
  nand ginst7920 (P1_U7192, P1_INSTQUEUE_REG_3__1__SCAN_IN, P1_U2570);
  nand ginst7921 (P1_U7193, P1_INSTQUEUE_REG_4__1__SCAN_IN, P1_U2568);
  nand ginst7922 (P1_U7194, P1_INSTQUEUE_REG_5__1__SCAN_IN, P1_U2567);
  nand ginst7923 (P1_U7195, P1_INSTQUEUE_REG_6__1__SCAN_IN, P1_U2566);
  nand ginst7924 (P1_U7196, P1_INSTQUEUE_REG_7__1__SCAN_IN, P1_U2565);
  nand ginst7925 (P1_U7197, P1_U4100, P1_U4101, P1_U4102, P1_U4103);
  nand ginst7926 (P1_U7198, P1_INSTQUEUE_REG_8__0__SCAN_IN, P1_U2582);
  nand ginst7927 (P1_U7199, P1_INSTQUEUE_REG_9__0__SCAN_IN, P1_U2581);
  nand ginst7928 (P1_U7200, P1_INSTQUEUE_REG_10__0__SCAN_IN, P1_U2580);
  nand ginst7929 (P1_U7201, P1_INSTQUEUE_REG_11__0__SCAN_IN, P1_U2579);
  nand ginst7930 (P1_U7202, P1_INSTQUEUE_REG_12__0__SCAN_IN, P1_U2577);
  nand ginst7931 (P1_U7203, P1_INSTQUEUE_REG_13__0__SCAN_IN, P1_U2576);
  nand ginst7932 (P1_U7204, P1_INSTQUEUE_REG_14__0__SCAN_IN, P1_U2575);
  nand ginst7933 (P1_U7205, P1_INSTQUEUE_REG_15__0__SCAN_IN, P1_U2574);
  nand ginst7934 (P1_U7206, P1_INSTQUEUE_REG_0__0__SCAN_IN, P1_U2573);
  nand ginst7935 (P1_U7207, P1_INSTQUEUE_REG_1__0__SCAN_IN, P1_U2572);
  nand ginst7936 (P1_U7208, P1_INSTQUEUE_REG_2__0__SCAN_IN, P1_U2571);
  nand ginst7937 (P1_U7209, P1_INSTQUEUE_REG_3__0__SCAN_IN, P1_U2570);
  nand ginst7938 (P1_U7210, P1_INSTQUEUE_REG_4__0__SCAN_IN, P1_U2568);
  nand ginst7939 (P1_U7211, P1_INSTQUEUE_REG_5__0__SCAN_IN, P1_U2567);
  nand ginst7940 (P1_U7212, P1_INSTQUEUE_REG_6__0__SCAN_IN, P1_U2566);
  nand ginst7941 (P1_U7213, P1_INSTQUEUE_REG_7__0__SCAN_IN, P1_U2565);
  nand ginst7942 (P1_U7214, P1_U4104, P1_U4105, P1_U4106, P1_U4107);
  nand ginst7943 (P1_U7215, P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN, P1_U3297);
  nand ginst7944 (P1_U7216, P1_U3455, P1_U4203);
  nand ginst7945 (P1_U7217, P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN, P1_U3297);
  nand ginst7946 (P1_U7218, P1_U3235, P1_U4203);
  not ginst7947 (P1_U7219, P1_U4183);
  nand ginst7948 (P1_U7220, P1_INSTQUEUE_REG_8__7__SCAN_IN, P1_U2602);
  nand ginst7949 (P1_U7221, P1_INSTQUEUE_REG_9__7__SCAN_IN, P1_U2601);
  nand ginst7950 (P1_U7222, P1_INSTQUEUE_REG_10__7__SCAN_IN, P1_U2600);
  nand ginst7951 (P1_U7223, P1_INSTQUEUE_REG_11__7__SCAN_IN, P1_U2599);
  nand ginst7952 (P1_U7224, P1_INSTQUEUE_REG_12__7__SCAN_IN, P1_U2597);
  nand ginst7953 (P1_U7225, P1_INSTQUEUE_REG_13__7__SCAN_IN, P1_U2596);
  nand ginst7954 (P1_U7226, P1_INSTQUEUE_REG_14__7__SCAN_IN, P1_U2595);
  nand ginst7955 (P1_U7227, P1_INSTQUEUE_REG_15__7__SCAN_IN, P1_U2594);
  nand ginst7956 (P1_U7228, P1_INSTQUEUE_REG_0__7__SCAN_IN, P1_U2592);
  nand ginst7957 (P1_U7229, P1_INSTQUEUE_REG_1__7__SCAN_IN, P1_U2591);
  nand ginst7958 (P1_U7230, P1_INSTQUEUE_REG_2__7__SCAN_IN, P1_U2590);
  nand ginst7959 (P1_U7231, P1_INSTQUEUE_REG_3__7__SCAN_IN, P1_U2589);
  nand ginst7960 (P1_U7232, P1_INSTQUEUE_REG_4__7__SCAN_IN, P1_U2587);
  nand ginst7961 (P1_U7233, P1_INSTQUEUE_REG_5__7__SCAN_IN, P1_U2586);
  nand ginst7962 (P1_U7234, P1_INSTQUEUE_REG_6__7__SCAN_IN, P1_U2585);
  nand ginst7963 (P1_U7235, P1_INSTQUEUE_REG_7__7__SCAN_IN, P1_U2584);
  nand ginst7964 (P1_U7236, P1_U4121, P1_U4122, P1_U4123, P1_U4124);
  nand ginst7965 (P1_U7237, P1_INSTQUEUE_REG_8__6__SCAN_IN, P1_U2602);
  nand ginst7966 (P1_U7238, P1_INSTQUEUE_REG_9__6__SCAN_IN, P1_U2601);
  nand ginst7967 (P1_U7239, P1_INSTQUEUE_REG_10__6__SCAN_IN, P1_U2600);
  nand ginst7968 (P1_U7240, P1_INSTQUEUE_REG_11__6__SCAN_IN, P1_U2599);
  nand ginst7969 (P1_U7241, P1_INSTQUEUE_REG_12__6__SCAN_IN, P1_U2597);
  nand ginst7970 (P1_U7242, P1_INSTQUEUE_REG_13__6__SCAN_IN, P1_U2596);
  nand ginst7971 (P1_U7243, P1_INSTQUEUE_REG_14__6__SCAN_IN, P1_U2595);
  nand ginst7972 (P1_U7244, P1_INSTQUEUE_REG_15__6__SCAN_IN, P1_U2594);
  nand ginst7973 (P1_U7245, P1_INSTQUEUE_REG_0__6__SCAN_IN, P1_U2592);
  nand ginst7974 (P1_U7246, P1_INSTQUEUE_REG_1__6__SCAN_IN, P1_U2591);
  nand ginst7975 (P1_U7247, P1_INSTQUEUE_REG_2__6__SCAN_IN, P1_U2590);
  nand ginst7976 (P1_U7248, P1_INSTQUEUE_REG_3__6__SCAN_IN, P1_U2589);
  nand ginst7977 (P1_U7249, P1_INSTQUEUE_REG_4__6__SCAN_IN, P1_U2587);
  nand ginst7978 (P1_U7250, P1_INSTQUEUE_REG_5__6__SCAN_IN, P1_U2586);
  nand ginst7979 (P1_U7251, P1_INSTQUEUE_REG_6__6__SCAN_IN, P1_U2585);
  nand ginst7980 (P1_U7252, P1_INSTQUEUE_REG_7__6__SCAN_IN, P1_U2584);
  nand ginst7981 (P1_U7253, P1_U4125, P1_U4126, P1_U4127, P1_U4128);
  nand ginst7982 (P1_U7254, P1_INSTQUEUE_REG_8__5__SCAN_IN, P1_U2602);
  nand ginst7983 (P1_U7255, P1_INSTQUEUE_REG_9__5__SCAN_IN, P1_U2601);
  nand ginst7984 (P1_U7256, P1_INSTQUEUE_REG_10__5__SCAN_IN, P1_U2600);
  nand ginst7985 (P1_U7257, P1_INSTQUEUE_REG_11__5__SCAN_IN, P1_U2599);
  nand ginst7986 (P1_U7258, P1_INSTQUEUE_REG_12__5__SCAN_IN, P1_U2597);
  nand ginst7987 (P1_U7259, P1_INSTQUEUE_REG_13__5__SCAN_IN, P1_U2596);
  nand ginst7988 (P1_U7260, P1_INSTQUEUE_REG_14__5__SCAN_IN, P1_U2595);
  nand ginst7989 (P1_U7261, P1_INSTQUEUE_REG_15__5__SCAN_IN, P1_U2594);
  nand ginst7990 (P1_U7262, P1_INSTQUEUE_REG_0__5__SCAN_IN, P1_U2592);
  nand ginst7991 (P1_U7263, P1_INSTQUEUE_REG_1__5__SCAN_IN, P1_U2591);
  nand ginst7992 (P1_U7264, P1_INSTQUEUE_REG_2__5__SCAN_IN, P1_U2590);
  nand ginst7993 (P1_U7265, P1_INSTQUEUE_REG_3__5__SCAN_IN, P1_U2589);
  nand ginst7994 (P1_U7266, P1_INSTQUEUE_REG_4__5__SCAN_IN, P1_U2587);
  nand ginst7995 (P1_U7267, P1_INSTQUEUE_REG_5__5__SCAN_IN, P1_U2586);
  nand ginst7996 (P1_U7268, P1_INSTQUEUE_REG_6__5__SCAN_IN, P1_U2585);
  nand ginst7997 (P1_U7269, P1_INSTQUEUE_REG_7__5__SCAN_IN, P1_U2584);
  nand ginst7998 (P1_U7270, P1_U4129, P1_U4130, P1_U4131, P1_U4132);
  nand ginst7999 (P1_U7271, P1_INSTQUEUE_REG_8__4__SCAN_IN, P1_U2602);
  nand ginst8000 (P1_U7272, P1_INSTQUEUE_REG_9__4__SCAN_IN, P1_U2601);
  nand ginst8001 (P1_U7273, P1_INSTQUEUE_REG_10__4__SCAN_IN, P1_U2600);
  nand ginst8002 (P1_U7274, P1_INSTQUEUE_REG_11__4__SCAN_IN, P1_U2599);
  nand ginst8003 (P1_U7275, P1_INSTQUEUE_REG_12__4__SCAN_IN, P1_U2597);
  nand ginst8004 (P1_U7276, P1_INSTQUEUE_REG_13__4__SCAN_IN, P1_U2596);
  nand ginst8005 (P1_U7277, P1_INSTQUEUE_REG_14__4__SCAN_IN, P1_U2595);
  nand ginst8006 (P1_U7278, P1_INSTQUEUE_REG_15__4__SCAN_IN, P1_U2594);
  nand ginst8007 (P1_U7279, P1_INSTQUEUE_REG_1__4__SCAN_IN, P1_U2591);
  nand ginst8008 (P1_U7280, P1_INSTQUEUE_REG_2__4__SCAN_IN, P1_U2590);
  nand ginst8009 (P1_U7281, P1_INSTQUEUE_REG_3__4__SCAN_IN, P1_U2589);
  nand ginst8010 (P1_U7282, P1_INSTQUEUE_REG_4__4__SCAN_IN, P1_U2587);
  nand ginst8011 (P1_U7283, P1_INSTQUEUE_REG_5__4__SCAN_IN, P1_U2586);
  nand ginst8012 (P1_U7284, P1_INSTQUEUE_REG_6__4__SCAN_IN, P1_U2585);
  nand ginst8013 (P1_U7285, P1_INSTQUEUE_REG_7__4__SCAN_IN, P1_U2584);
  nand ginst8014 (P1_U7286, P1_INSTQUEUE_REG_8__3__SCAN_IN, P1_U2602);
  nand ginst8015 (P1_U7287, P1_INSTQUEUE_REG_9__3__SCAN_IN, P1_U2601);
  nand ginst8016 (P1_U7288, P1_INSTQUEUE_REG_10__3__SCAN_IN, P1_U2600);
  nand ginst8017 (P1_U7289, P1_INSTQUEUE_REG_11__3__SCAN_IN, P1_U2599);
  nand ginst8018 (P1_U7290, P1_INSTQUEUE_REG_12__3__SCAN_IN, P1_U2597);
  nand ginst8019 (P1_U7291, P1_INSTQUEUE_REG_13__3__SCAN_IN, P1_U2596);
  nand ginst8020 (P1_U7292, P1_INSTQUEUE_REG_14__3__SCAN_IN, P1_U2595);
  nand ginst8021 (P1_U7293, P1_INSTQUEUE_REG_15__3__SCAN_IN, P1_U2594);
  nand ginst8022 (P1_U7294, P1_INSTQUEUE_REG_0__3__SCAN_IN, P1_U2592);
  nand ginst8023 (P1_U7295, P1_INSTQUEUE_REG_1__3__SCAN_IN, P1_U2591);
  nand ginst8024 (P1_U7296, P1_INSTQUEUE_REG_2__3__SCAN_IN, P1_U2590);
  nand ginst8025 (P1_U7297, P1_INSTQUEUE_REG_3__3__SCAN_IN, P1_U2589);
  nand ginst8026 (P1_U7298, P1_INSTQUEUE_REG_4__3__SCAN_IN, P1_U2587);
  nand ginst8027 (P1_U7299, P1_INSTQUEUE_REG_5__3__SCAN_IN, P1_U2586);
  nand ginst8028 (P1_U7300, P1_INSTQUEUE_REG_6__3__SCAN_IN, P1_U2585);
  nand ginst8029 (P1_U7301, P1_INSTQUEUE_REG_7__3__SCAN_IN, P1_U2584);
  nand ginst8030 (P1_U7302, P1_U4137, P1_U4138, P1_U4139, P1_U4140);
  nand ginst8031 (P1_U7303, P1_INSTQUEUE_REG_8__2__SCAN_IN, P1_U2602);
  nand ginst8032 (P1_U7304, P1_INSTQUEUE_REG_9__2__SCAN_IN, P1_U2601);
  nand ginst8033 (P1_U7305, P1_INSTQUEUE_REG_10__2__SCAN_IN, P1_U2600);
  nand ginst8034 (P1_U7306, P1_INSTQUEUE_REG_11__2__SCAN_IN, P1_U2599);
  nand ginst8035 (P1_U7307, P1_INSTQUEUE_REG_12__2__SCAN_IN, P1_U2597);
  nand ginst8036 (P1_U7308, P1_INSTQUEUE_REG_13__2__SCAN_IN, P1_U2596);
  nand ginst8037 (P1_U7309, P1_INSTQUEUE_REG_14__2__SCAN_IN, P1_U2595);
  nand ginst8038 (P1_U7310, P1_INSTQUEUE_REG_15__2__SCAN_IN, P1_U2594);
  nand ginst8039 (P1_U7311, P1_INSTQUEUE_REG_0__2__SCAN_IN, P1_U2592);
  nand ginst8040 (P1_U7312, P1_INSTQUEUE_REG_1__2__SCAN_IN, P1_U2591);
  nand ginst8041 (P1_U7313, P1_INSTQUEUE_REG_2__2__SCAN_IN, P1_U2590);
  nand ginst8042 (P1_U7314, P1_INSTQUEUE_REG_3__2__SCAN_IN, P1_U2589);
  nand ginst8043 (P1_U7315, P1_INSTQUEUE_REG_4__2__SCAN_IN, P1_U2587);
  nand ginst8044 (P1_U7316, P1_INSTQUEUE_REG_5__2__SCAN_IN, P1_U2586);
  nand ginst8045 (P1_U7317, P1_INSTQUEUE_REG_6__2__SCAN_IN, P1_U2585);
  nand ginst8046 (P1_U7318, P1_INSTQUEUE_REG_7__2__SCAN_IN, P1_U2584);
  nand ginst8047 (P1_U7319, P1_U4141, P1_U4142, P1_U4143, P1_U4144);
  nand ginst8048 (P1_U7320, P1_INSTQUEUE_REG_8__1__SCAN_IN, P1_U2602);
  nand ginst8049 (P1_U7321, P1_INSTQUEUE_REG_9__1__SCAN_IN, P1_U2601);
  nand ginst8050 (P1_U7322, P1_INSTQUEUE_REG_10__1__SCAN_IN, P1_U2600);
  nand ginst8051 (P1_U7323, P1_INSTQUEUE_REG_11__1__SCAN_IN, P1_U2599);
  nand ginst8052 (P1_U7324, P1_INSTQUEUE_REG_12__1__SCAN_IN, P1_U2597);
  nand ginst8053 (P1_U7325, P1_INSTQUEUE_REG_13__1__SCAN_IN, P1_U2596);
  nand ginst8054 (P1_U7326, P1_INSTQUEUE_REG_14__1__SCAN_IN, P1_U2595);
  nand ginst8055 (P1_U7327, P1_INSTQUEUE_REG_15__1__SCAN_IN, P1_U2594);
  nand ginst8056 (P1_U7328, P1_INSTQUEUE_REG_0__1__SCAN_IN, P1_U2592);
  nand ginst8057 (P1_U7329, P1_INSTQUEUE_REG_1__1__SCAN_IN, P1_U2591);
  nand ginst8058 (P1_U7330, P1_INSTQUEUE_REG_2__1__SCAN_IN, P1_U2590);
  nand ginst8059 (P1_U7331, P1_INSTQUEUE_REG_3__1__SCAN_IN, P1_U2589);
  nand ginst8060 (P1_U7332, P1_INSTQUEUE_REG_4__1__SCAN_IN, P1_U2587);
  nand ginst8061 (P1_U7333, P1_INSTQUEUE_REG_5__1__SCAN_IN, P1_U2586);
  nand ginst8062 (P1_U7334, P1_INSTQUEUE_REG_6__1__SCAN_IN, P1_U2585);
  nand ginst8063 (P1_U7335, P1_INSTQUEUE_REG_7__1__SCAN_IN, P1_U2584);
  nand ginst8064 (P1_U7336, P1_U4145, P1_U4146, P1_U4147, P1_U4148);
  nand ginst8065 (P1_U7337, P1_INSTQUEUE_REG_8__0__SCAN_IN, P1_U2602);
  nand ginst8066 (P1_U7338, P1_INSTQUEUE_REG_9__0__SCAN_IN, P1_U2601);
  nand ginst8067 (P1_U7339, P1_INSTQUEUE_REG_10__0__SCAN_IN, P1_U2600);
  nand ginst8068 (P1_U7340, P1_INSTQUEUE_REG_11__0__SCAN_IN, P1_U2599);
  nand ginst8069 (P1_U7341, P1_INSTQUEUE_REG_12__0__SCAN_IN, P1_U2597);
  nand ginst8070 (P1_U7342, P1_INSTQUEUE_REG_13__0__SCAN_IN, P1_U2596);
  nand ginst8071 (P1_U7343, P1_INSTQUEUE_REG_14__0__SCAN_IN, P1_U2595);
  nand ginst8072 (P1_U7344, P1_INSTQUEUE_REG_15__0__SCAN_IN, P1_U2594);
  nand ginst8073 (P1_U7345, P1_INSTQUEUE_REG_0__0__SCAN_IN, P1_U2592);
  nand ginst8074 (P1_U7346, P1_INSTQUEUE_REG_1__0__SCAN_IN, P1_U2591);
  nand ginst8075 (P1_U7347, P1_INSTQUEUE_REG_2__0__SCAN_IN, P1_U2590);
  nand ginst8076 (P1_U7348, P1_INSTQUEUE_REG_3__0__SCAN_IN, P1_U2589);
  nand ginst8077 (P1_U7349, P1_INSTQUEUE_REG_4__0__SCAN_IN, P1_U2587);
  nand ginst8078 (P1_U7350, P1_INSTQUEUE_REG_5__0__SCAN_IN, P1_U2586);
  nand ginst8079 (P1_U7351, P1_INSTQUEUE_REG_6__0__SCAN_IN, P1_U2585);
  nand ginst8080 (P1_U7352, P1_INSTQUEUE_REG_7__0__SCAN_IN, P1_U2584);
  nand ginst8081 (P1_U7353, P1_U4149, P1_U4150, P1_U4151, P1_U4152);
  nand ginst8082 (P1_U7354, P1_U2354, P1_U4231, P1_U4234);
  nand ginst8083 (P1_U7355, P1_U4153, P1_U7087);
  nand ginst8084 (P1_U7356, P1_U3396, P1_U3410);
  nand ginst8085 (P1_U7357, P1_U4234, P1_U7356);
  nand ginst8086 (P1_U7358, P1_U2452, P1_U4190);
  nand ginst8087 (P1_U7359, P1_U3271, P1_U7355);
  nand ginst8088 (P1_U7360, P1_U4208, P1_U7088);
  nand ginst8089 (P1_U7361, P1_U4160, P1_U4208);
  nand ginst8090 (P1_U7362, P1_U2451, P1_U4210);
  nand ginst8091 (P1_U7363, P1_U3420, P1_U3434, P1_U4195, P1_U7361, P1_U7362);
  nand ginst8092 (P1_U7364, P1_R2238_U6, P1_U7363);
  nand ginst8093 (P1_U7365, P1_SUB_450_U6, P1_U2354);
  nand ginst8094 (P1_U7366, P1_R2238_U19, P1_U7363);
  nand ginst8095 (P1_U7367, P1_SUB_450_U19, P1_U2354);
  nand ginst8096 (P1_U7368, P1_R2238_U20, P1_U7363);
  nand ginst8097 (P1_U7369, P1_SUB_450_U20, P1_U2354);
  nand ginst8098 (P1_U7370, P1_R2238_U21, P1_U7363);
  nand ginst8099 (P1_U7371, P1_SUB_450_U21, P1_U2354);
  nand ginst8100 (P1_U7372, P1_R2238_U22, P1_U7363);
  nand ginst8101 (P1_U7373, P1_SUB_450_U22, P1_U2354);
  nand ginst8102 (P1_U7374, P1_R2238_U7, P1_U7363);
  nand ginst8103 (P1_U7375, P1_SUB_450_U7, P1_U2354);
  nand ginst8104 (P1_U7376, P1_R2238_U19, P1_U4192);
  nand ginst8105 (P1_U7377, P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN, P1_U3294);
  nand ginst8106 (P1_U7378, P1_R2238_U20, P1_U4192);
  nand ginst8107 (P1_U7379, P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P1_U3294);
  nand ginst8108 (P1_U7380, P1_STATE2_REG_0__SCAN_IN, P1_U4173);
  nand ginst8109 (P1_U7381, P1_U3420, P1_U7380);
  nand ginst8110 (P1_U7382, P1_R2238_U21, P1_U4192);
  nand ginst8111 (P1_U7383, P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN, P1_U3294);
  nand ginst8112 (P1_U7384, P1_U2450, P1_U3271);
  nand ginst8113 (P1_U7385, P1_R2238_U22, P1_U4192);
  nand ginst8114 (P1_U7386, P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P1_U3294);
  nand ginst8115 (P1_U7387, P1_U2451, P1_U3284);
  nand ginst8116 (P1_U7388, P1_R2238_U7, P1_U4192);
  nand ginst8117 (P1_U7389, P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN, P1_U3294);
  nand ginst8118 (P1_U7390, P1_U3290, P1_U3393);
  nand ginst8119 (P1_U7391, P1_U3284, P1_U3449);
  nand ginst8120 (P1_U7392, P1_INSTADDRPOINTER_REG_9__SCAN_IN, P1_U7391);
  nand ginst8121 (P1_U7393, P1_EBX_REG_9__SCAN_IN, P1_U7390);
  nand ginst8122 (P1_U7394, P1_INSTADDRPOINTER_REG_8__SCAN_IN, P1_U7391);
  nand ginst8123 (P1_U7395, P1_EBX_REG_8__SCAN_IN, P1_U7390);
  nand ginst8124 (P1_U7396, P1_INSTADDRPOINTER_REG_7__SCAN_IN, P1_U7391);
  nand ginst8125 (P1_U7397, P1_EBX_REG_7__SCAN_IN, P1_U7390);
  nand ginst8126 (P1_U7398, P1_INSTADDRPOINTER_REG_6__SCAN_IN, P1_U7391);
  nand ginst8127 (P1_U7399, P1_EBX_REG_6__SCAN_IN, P1_U7390);
  nand ginst8128 (P1_U7400, P1_INSTADDRPOINTER_REG_5__SCAN_IN, P1_U7391);
  nand ginst8129 (P1_U7401, P1_EBX_REG_5__SCAN_IN, P1_U7390);
  nand ginst8130 (P1_U7402, P1_INSTADDRPOINTER_REG_4__SCAN_IN, P1_U7391);
  nand ginst8131 (P1_U7403, P1_EBX_REG_4__SCAN_IN, P1_U7390);
  nand ginst8132 (P1_U7404, P1_INSTADDRPOINTER_REG_31__SCAN_IN, P1_U7391);
  nand ginst8133 (P1_U7405, P1_EBX_REG_31__SCAN_IN, P1_U7390);
  nand ginst8134 (P1_U7406, P1_INSTADDRPOINTER_REG_30__SCAN_IN, P1_U7391);
  nand ginst8135 (P1_U7407, P1_EBX_REG_30__SCAN_IN, P1_U7390);
  nand ginst8136 (P1_U7408, P1_INSTADDRPOINTER_REG_3__SCAN_IN, P1_U7391);
  nand ginst8137 (P1_U7409, P1_EBX_REG_3__SCAN_IN, P1_U7390);
  nand ginst8138 (P1_U7410, P1_INSTADDRPOINTER_REG_29__SCAN_IN, P1_U7391);
  nand ginst8139 (P1_U7411, P1_EBX_REG_29__SCAN_IN, P1_U7390);
  nand ginst8140 (P1_U7412, P1_INSTADDRPOINTER_REG_28__SCAN_IN, P1_U7391);
  nand ginst8141 (P1_U7413, P1_EBX_REG_28__SCAN_IN, P1_U7390);
  nand ginst8142 (P1_U7414, P1_INSTADDRPOINTER_REG_27__SCAN_IN, P1_U7391);
  nand ginst8143 (P1_U7415, P1_EBX_REG_27__SCAN_IN, P1_U7390);
  nand ginst8144 (P1_U7416, P1_INSTADDRPOINTER_REG_26__SCAN_IN, P1_U7391);
  nand ginst8145 (P1_U7417, P1_EBX_REG_26__SCAN_IN, P1_U7390);
  nand ginst8146 (P1_U7418, P1_INSTADDRPOINTER_REG_25__SCAN_IN, P1_U7391);
  nand ginst8147 (P1_U7419, P1_EBX_REG_25__SCAN_IN, P1_U7390);
  nand ginst8148 (P1_U7420, P1_INSTADDRPOINTER_REG_24__SCAN_IN, P1_U7391);
  nand ginst8149 (P1_U7421, P1_EBX_REG_24__SCAN_IN, P1_U7390);
  nand ginst8150 (P1_U7422, P1_INSTADDRPOINTER_REG_23__SCAN_IN, P1_U7391);
  nand ginst8151 (P1_U7423, P1_EBX_REG_23__SCAN_IN, P1_U7390);
  nand ginst8152 (P1_U7424, P1_INSTADDRPOINTER_REG_22__SCAN_IN, P1_U7391);
  nand ginst8153 (P1_U7425, P1_EBX_REG_22__SCAN_IN, P1_U7390);
  nand ginst8154 (P1_U7426, P1_INSTADDRPOINTER_REG_21__SCAN_IN, P1_U7391);
  nand ginst8155 (P1_U7427, P1_EBX_REG_21__SCAN_IN, P1_U7390);
  nand ginst8156 (P1_U7428, P1_INSTADDRPOINTER_REG_20__SCAN_IN, P1_U7391);
  nand ginst8157 (P1_U7429, P1_EBX_REG_20__SCAN_IN, P1_U7390);
  nand ginst8158 (P1_U7430, P1_INSTADDRPOINTER_REG_2__SCAN_IN, P1_U7391);
  nand ginst8159 (P1_U7431, P1_EBX_REG_2__SCAN_IN, P1_U7390);
  nand ginst8160 (P1_U7432, P1_INSTADDRPOINTER_REG_19__SCAN_IN, P1_U7391);
  nand ginst8161 (P1_U7433, P1_EBX_REG_19__SCAN_IN, P1_U7390);
  nand ginst8162 (P1_U7434, P1_INSTADDRPOINTER_REG_18__SCAN_IN, P1_U7391);
  nand ginst8163 (P1_U7435, P1_EBX_REG_18__SCAN_IN, P1_U7390);
  nand ginst8164 (P1_U7436, P1_INSTADDRPOINTER_REG_17__SCAN_IN, P1_U7391);
  nand ginst8165 (P1_U7437, P1_EBX_REG_17__SCAN_IN, P1_U7390);
  nand ginst8166 (P1_U7438, P1_INSTADDRPOINTER_REG_16__SCAN_IN, P1_U7391);
  nand ginst8167 (P1_U7439, P1_EBX_REG_16__SCAN_IN, P1_U7390);
  nand ginst8168 (P1_U7440, P1_INSTADDRPOINTER_REG_15__SCAN_IN, P1_U7391);
  nand ginst8169 (P1_U7441, P1_EBX_REG_15__SCAN_IN, P1_U7390);
  nand ginst8170 (P1_U7442, P1_INSTADDRPOINTER_REG_14__SCAN_IN, P1_U7391);
  nand ginst8171 (P1_U7443, P1_EBX_REG_14__SCAN_IN, P1_U7390);
  nand ginst8172 (P1_U7444, P1_INSTADDRPOINTER_REG_13__SCAN_IN, P1_U7391);
  nand ginst8173 (P1_U7445, P1_EBX_REG_13__SCAN_IN, P1_U7390);
  nand ginst8174 (P1_U7446, P1_INSTADDRPOINTER_REG_12__SCAN_IN, P1_U7391);
  nand ginst8175 (P1_U7447, P1_EBX_REG_12__SCAN_IN, P1_U7390);
  nand ginst8176 (P1_U7448, P1_INSTADDRPOINTER_REG_11__SCAN_IN, P1_U7391);
  nand ginst8177 (P1_U7449, P1_EBX_REG_11__SCAN_IN, P1_U7390);
  nand ginst8178 (P1_U7450, P1_INSTADDRPOINTER_REG_10__SCAN_IN, P1_U7391);
  nand ginst8179 (P1_U7451, P1_EBX_REG_10__SCAN_IN, P1_U7390);
  nand ginst8180 (P1_U7452, P1_INSTADDRPOINTER_REG_1__SCAN_IN, P1_U7391);
  nand ginst8181 (P1_U7453, P1_EBX_REG_1__SCAN_IN, P1_U7390);
  nand ginst8182 (P1_U7454, P1_INSTADDRPOINTER_REG_0__SCAN_IN, P1_U7391);
  nand ginst8183 (P1_U7455, P1_EBX_REG_0__SCAN_IN, P1_U7390);
  nand ginst8184 (P1_U7456, P1_U4477, P1_U4496);
  nand ginst8185 (P1_U7457, P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN, P1_U2430);
  nand ginst8186 (P1_U7458, P1_U3262, P1_U3489);
  nand ginst8187 (P1_U7459, P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P1_U2430);
  nand ginst8188 (P1_U7460, P1_U3262, P1_U3490);
  nand ginst8189 (P1_U7461, P1_FLUSH_REG_SCAN_IN, P1_U2446, P1_U3470);
  nand ginst8190 (P1_U7462, P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN, P1_U2430);
  nand ginst8191 (P1_U7463, P1_U3262, P1_U3491);
  nand ginst8192 (P1_U7464, P1_FLUSH_REG_SCAN_IN, P1_U2446, P1_U7712);
  nand ginst8193 (P1_U7465, P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P1_U2430);
  nand ginst8194 (P1_U7466, P1_U3262, P1_U3492);
  nand ginst8195 (P1_U7467, P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN, P1_U2430);
  nand ginst8196 (P1_U7468, P1_STATE_REG_0__SCAN_IN, P1_U4185);
  or ginst8197 (P1_U7469, P1_STATE2_REG_2__SCAN_IN, U210);
  nand ginst8198 (P1_U7470, P1_U4110, P1_U7218);
  nand ginst8199 (P1_U7471, P1_U3422, P1_U7084);
  nand ginst8200 (P1_U7472, P1_STATE2_REG_0__SCAN_IN, P1_U4211);
  nand ginst8201 (P1_U7473, P1_STATE2_REG_0__SCAN_IN, P1_U4212);
  nand ginst8202 (P1_U7474, P1_STATE2_REG_0__SCAN_IN, P1_U4213);
  nand ginst8203 (P1_U7475, P1_STATE2_REG_0__SCAN_IN, P1_U4236);
  nand ginst8204 (P1_U7476, P1_STATE2_REG_0__SCAN_IN, P1_U4264);
  nand ginst8205 (P1_U7477, P1_STATE2_REG_0__SCAN_IN, P1_U7632);
  nand ginst8206 (P1_U7478, P1_U2608, P1_U3266);
  nand ginst8207 (P1_U7479, P1_U4117, P1_U4118, P1_U4120, P1_U7093);
  nand ginst8208 (P1_U7480, P1_STATE2_REG_0__SCAN_IN, P1_U7632);
  nand ginst8209 (P1_U7481, P1_U2379, P1_U3429);
  nand ginst8210 (P1_U7482, P1_U2369, P1_U6367);
  nand ginst8211 (P1_U7483, P1_U2369, P1_U3888);
  nand ginst8212 (P1_U7484, P1_U4229, P1_U7481, P1_U7482);
  nand ginst8213 (P1_U7485, P1_U4230, P1_U7483);
  nand ginst8214 (P1_U7486, P1_U4171, P1_U4194, P1_U5491);
  nand ginst8215 (P1_U7487, P1_U4194, P1_U7091);
  nand ginst8216 (P1_U7488, P1_U3392, P1_U4194);
  nand ginst8217 (P1_U7489, P1_STATE2_REG_0__SCAN_IN, P1_U4236);
  nand ginst8218 (P1_U7490, P1_U4072, P1_U7784, P1_U7785);
  nand ginst8219 (P1_U7491, P1_U4108, P1_U7216);
  nand ginst8220 (P1_U7492, P1_U4109, P1_U7094);
  not ginst8221 (P1_U7493, P1_U3279);
  not ginst8222 (P1_U7494, P1_U3276);
  nand ginst8223 (P1_U7495, P1_U2607, P1_U4068, P1_U4069, P1_U4070, P1_U4071);
  nand ginst8224 (P1_U7496, P1_U3734, P1_U7493);
  nand ginst8225 (P1_U7497, P1_U3735, P1_U5469);
  nand ginst8226 (P1_U7498, P1_U2425, P1_U7493);
  nand ginst8227 (P1_U7499, P1_U2425, P1_U7493);
  nand ginst8228 (P1_U7500, P1_U6360, P1_U6361, P1_U7499);
  nand ginst8229 (P1_U7501, P1_R2167_U17, P1_U7493);
  nand ginst8230 (P1_U7502, P1_R2167_U17, P1_U4201, P1_U7493);
  nand ginst8231 (P1_U7503, P1_U6149, P1_U7502);
  nand ginst8232 (P1_U7504, P1_U7085, P1_U7493);
  nand ginst8233 (P1_U7505, P1_U7471, P1_U7493);
  nand ginst8234 (P1_U7506, P1_U4114, P1_U4115, P1_U4116);
  nand ginst8235 (P1_U7507, P1_U3759, P1_U7493);
  nand ginst8236 (P1_U7508, P1_U3760, P1_U3761, P1_U5565);
  nand ginst8237 (P1_U7509, P1_U2519, P1_U3746);
  nand ginst8238 (P1_U7510, P1_U5962, P1_U7493);
  nand ginst8239 (P1_U7511, P1_U5965, P1_U7493);
  nand ginst8240 (P1_U7512, P1_U5968, P1_U7493);
  nand ginst8241 (P1_U7513, P1_U5971, P1_U7493);
  nand ginst8242 (P1_U7514, P1_U5974, P1_U7493);
  nand ginst8243 (P1_U7515, P1_U5977, P1_U7493);
  nand ginst8244 (P1_U7516, P1_U5980, P1_U7493);
  nand ginst8245 (P1_U7517, P1_U5983, P1_U7493);
  nand ginst8246 (P1_U7518, P1_U5986, P1_U7493);
  nand ginst8247 (P1_U7519, P1_U5989, P1_U7493);
  nand ginst8248 (P1_U7520, P1_U5992, P1_U7493);
  nand ginst8249 (P1_U7521, P1_U5995, P1_U7493);
  nand ginst8250 (P1_U7522, P1_U5998, P1_U7493);
  nand ginst8251 (P1_U7523, P1_U6001, P1_U7493);
  nand ginst8252 (P1_U7524, P1_U6004, P1_U7493);
  nand ginst8253 (P1_U7525, P1_U6007, P1_U7493);
  nand ginst8254 (P1_U7526, P1_U6010, P1_U7493);
  nand ginst8255 (P1_U7527, P1_U6013, P1_U7493);
  nand ginst8256 (P1_U7528, P1_U6016, P1_U7493);
  nand ginst8257 (P1_U7529, P1_U6019, P1_U7493);
  nand ginst8258 (P1_U7530, P1_U6022, P1_U7493);
  nand ginst8259 (P1_U7531, P1_U6025, P1_U7493);
  nand ginst8260 (P1_U7532, P1_U6028, P1_U7493);
  nand ginst8261 (P1_U7533, P1_U6031, P1_U7493);
  nand ginst8262 (P1_U7534, P1_U6034, P1_U7493);
  nand ginst8263 (P1_U7535, P1_U6037, P1_U7493);
  nand ginst8264 (P1_U7536, P1_U6040, P1_U7493);
  nand ginst8265 (P1_U7537, P1_U6043, P1_U7493);
  nand ginst8266 (P1_U7538, P1_U6046, P1_U7493);
  nand ginst8267 (P1_U7539, P1_U6049, P1_U7493);
  nand ginst8268 (P1_U7540, P1_U6052, P1_U7493);
  nand ginst8269 (P1_U7541, P1_U2357, P1_U7493);
  nand ginst8270 (P1_U7542, P1_UWORD_REG_0__SCAN_IN, P1_U7541);
  nand ginst8271 (P1_U7543, P1_U2357, P1_U7493);
  nand ginst8272 (P1_U7544, P1_UWORD_REG_1__SCAN_IN, P1_U7543);
  nand ginst8273 (P1_U7545, P1_U2357, P1_U7493);
  nand ginst8274 (P1_U7546, P1_UWORD_REG_2__SCAN_IN, P1_U7545);
  nand ginst8275 (P1_U7547, P1_U2357, P1_U7493);
  nand ginst8276 (P1_U7548, P1_UWORD_REG_3__SCAN_IN, P1_U7547);
  nand ginst8277 (P1_U7549, P1_U2357, P1_U7493);
  nand ginst8278 (P1_U7550, P1_UWORD_REG_4__SCAN_IN, P1_U7549);
  nand ginst8279 (P1_U7551, P1_U2357, P1_U7493);
  nand ginst8280 (P1_U7552, P1_UWORD_REG_5__SCAN_IN, P1_U7551);
  nand ginst8281 (P1_U7553, P1_U2357, P1_U7493);
  nand ginst8282 (P1_U7554, P1_UWORD_REG_6__SCAN_IN, P1_U7553);
  nand ginst8283 (P1_U7555, P1_U2357, P1_U7493);
  nand ginst8284 (P1_U7556, P1_UWORD_REG_7__SCAN_IN, P1_U7555);
  nand ginst8285 (P1_U7557, P1_U2357, P1_U7493);
  nand ginst8286 (P1_U7558, P1_UWORD_REG_8__SCAN_IN, P1_U7557);
  nand ginst8287 (P1_U7559, P1_U2357, P1_U7493);
  nand ginst8288 (P1_U7560, P1_UWORD_REG_9__SCAN_IN, P1_U7559);
  nand ginst8289 (P1_U7561, P1_U2357, P1_U7493);
  nand ginst8290 (P1_U7562, P1_UWORD_REG_10__SCAN_IN, P1_U7561);
  nand ginst8291 (P1_U7563, P1_U2357, P1_U7493);
  nand ginst8292 (P1_U7564, P1_UWORD_REG_11__SCAN_IN, P1_U7563);
  nand ginst8293 (P1_U7565, P1_U2357, P1_U7493);
  nand ginst8294 (P1_U7566, P1_UWORD_REG_12__SCAN_IN, P1_U7565);
  nand ginst8295 (P1_U7567, P1_U2357, P1_U7493);
  nand ginst8296 (P1_U7568, P1_UWORD_REG_13__SCAN_IN, P1_U7567);
  nand ginst8297 (P1_U7569, P1_U2357, P1_U7493);
  nand ginst8298 (P1_U7570, P1_UWORD_REG_14__SCAN_IN, P1_U7569);
  nand ginst8299 (P1_U7571, P1_U2357, P1_U7493);
  nand ginst8300 (P1_U7572, P1_LWORD_REG_0__SCAN_IN, P1_U7571);
  nand ginst8301 (P1_U7573, P1_U2357, P1_U7493);
  nand ginst8302 (P1_U7574, P1_LWORD_REG_1__SCAN_IN, P1_U7573);
  nand ginst8303 (P1_U7575, P1_U2357, P1_U7493);
  nand ginst8304 (P1_U7576, P1_LWORD_REG_2__SCAN_IN, P1_U7575);
  nand ginst8305 (P1_U7577, P1_U2357, P1_U7493);
  nand ginst8306 (P1_U7578, P1_LWORD_REG_3__SCAN_IN, P1_U7577);
  nand ginst8307 (P1_U7579, P1_U2357, P1_U7493);
  nand ginst8308 (P1_U7580, P1_LWORD_REG_4__SCAN_IN, P1_U7579);
  nand ginst8309 (P1_U7581, P1_U2357, P1_U7493);
  nand ginst8310 (P1_U7582, P1_LWORD_REG_5__SCAN_IN, P1_U7581);
  nand ginst8311 (P1_U7583, P1_U2357, P1_U7493);
  nand ginst8312 (P1_U7584, P1_LWORD_REG_6__SCAN_IN, P1_U7583);
  nand ginst8313 (P1_U7585, P1_U2357, P1_U7493);
  nand ginst8314 (P1_U7586, P1_LWORD_REG_7__SCAN_IN, P1_U7585);
  nand ginst8315 (P1_U7587, P1_U2357, P1_U7493);
  nand ginst8316 (P1_U7588, P1_LWORD_REG_8__SCAN_IN, P1_U7587);
  nand ginst8317 (P1_U7589, P1_U2357, P1_U7493);
  nand ginst8318 (P1_U7590, P1_LWORD_REG_9__SCAN_IN, P1_U7589);
  nand ginst8319 (P1_U7591, P1_U2357, P1_U7493);
  nand ginst8320 (P1_U7592, P1_LWORD_REG_10__SCAN_IN, P1_U7591);
  nand ginst8321 (P1_U7593, P1_U2357, P1_U7493);
  nand ginst8322 (P1_U7594, P1_LWORD_REG_11__SCAN_IN, P1_U7593);
  nand ginst8323 (P1_U7595, P1_U2357, P1_U7493);
  nand ginst8324 (P1_U7596, P1_LWORD_REG_12__SCAN_IN, P1_U7595);
  nand ginst8325 (P1_U7597, P1_U2357, P1_U7493);
  nand ginst8326 (P1_U7598, P1_LWORD_REG_13__SCAN_IN, P1_U7597);
  nand ginst8327 (P1_U7599, P1_U2357, P1_U7493);
  nand ginst8328 (P1_U7600, P1_LWORD_REG_14__SCAN_IN, P1_U7599);
  nand ginst8329 (P1_U7601, P1_U2357, P1_U7493);
  nand ginst8330 (P1_U7602, P1_LWORD_REG_15__SCAN_IN, P1_U7601);
  nand ginst8331 (P1_U7603, P1_U3568, P1_U4259, P1_U7493);
  nand ginst8332 (P1_U7604, P1_U3581, P1_U7683, P1_U7684);
  nand ginst8333 (P1_U7605, P1_U3867, P1_U7493);
  nand ginst8334 (P1_U7606, P1_U3428, P1_U7605);
  nand ginst8335 (P1_U7607, P1_U4208, P1_U7493);
  nand ginst8336 (P1_U7608, P1_U3447, P1_U7607);
  nand ginst8337 (P1_U7609, P1_U3279, P1_U3400);
  nand ginst8338 (P1_U7610, P1_U3754, P1_U7493);
  nand ginst8339 (P1_U7611, P1_U3755, P1_U7610);
  nand ginst8340 (P1_U7612, P1_INSTQUEUE_REG_0__4__SCAN_IN, P1_U5416);
  nand ginst8341 (P1_U7613, P1_INSTQUEUE_REG_0__4__SCAN_IN, P1_U2523);
  nand ginst8342 (P1_U7614, P1_INSTQUEUE_REG_0__4__SCAN_IN, P1_U2546);
  nand ginst8343 (P1_U7615, P1_U4049, P1_U4050, P1_U4051, P1_U4052);
  nand ginst8344 (P1_U7616, P1_INSTQUEUE_REG_0__4__SCAN_IN, P1_U4192);
  nand ginst8345 (P1_U7617, P1_INSTQUEUE_REG_0__4__SCAN_IN, P1_U2573);
  nand ginst8346 (P1_U7618, P1_U4087, P1_U4088, P1_U4089, P1_U4091);
  nand ginst8347 (P1_U7619, P1_INSTQUEUE_REG_0__4__SCAN_IN, P1_U2592);
  nand ginst8348 (P1_U7620, P1_U4133, P1_U4134, P1_U4135, P1_U4136);
  not ginst8349 (P1_U7621, P1_U3259);
  nand ginst8350 (P1_U7622, P1_U3261, P1_U7621);
  nand ginst8351 (P1_U7623, P1_STATE_REG_1__SCAN_IN, P1_U4358, P1_U4361);
  nand ginst8352 (P1_U7624, P1_STATE_REG_2__SCAN_IN, P1_U7468);
  nand ginst8353 (P1_U7625, P1_STATE_REG_1__SCAN_IN, P1_U4358);
  nand ginst8354 (P1_U7626, P1_U4502, P1_U4510);
  nand ginst8355 (P1_U7627, P1_U4171, P1_U5487);
  nand ginst8356 (P1_U7628, P1_U3283, P1_U3289);
  not ginst8357 (P1_U7629, P1_U3392);
  nand ginst8358 (P1_U7630, P1_U4208, P1_U7490);
  nand ginst8359 (P1_U7631, P1_U4171, P1_U5487);
  nand ginst8360 (P1_U7632, P1_U7630, P1_U7631);
  nand ginst8361 (P1_U7633, P1_BE_N_REG_3__SCAN_IN, P1_U3249);
  nand ginst8362 (P1_U7634, P1_BYTEENABLE_REG_3__SCAN_IN, P1_U4221);
  nand ginst8363 (P1_U7635, P1_BE_N_REG_2__SCAN_IN, P1_U3249);
  nand ginst8364 (P1_U7636, P1_BYTEENABLE_REG_2__SCAN_IN, P1_U4221);
  nand ginst8365 (P1_U7637, P1_BE_N_REG_1__SCAN_IN, P1_U3249);
  nand ginst8366 (P1_U7638, P1_BYTEENABLE_REG_1__SCAN_IN, P1_U4221);
  nand ginst8367 (P1_U7639, P1_BE_N_REG_0__SCAN_IN, P1_U3249);
  nand ginst8368 (P1_U7640, P1_BYTEENABLE_REG_0__SCAN_IN, P1_U4221);
  nand ginst8369 (P1_U7641, P1_REQUESTPENDING_REG_SCAN_IN, P1_STATE_REG_0__SCAN_IN, P1_U3251);
  nand ginst8370 (P1_U7642, P1_STATE_REG_2__SCAN_IN, P1_U3259);
  nand ginst8371 (P1_U7643, P1_U7641, P1_U7642);
  nand ginst8372 (P1_U7644, P1_STATE_REG_1__SCAN_IN, P1_U4361, P1_U7624);
  nand ginst8373 (P1_U7645, P1_U3248, P1_U7643);
  nand ginst8374 (P1_U7646, P1_STATE_REG_2__SCAN_IN, P1_STATE_REG_0__SCAN_IN, P1_U3260);
  nand ginst8375 (P1_U7647, P1_U3251, P1_U4371);
  or ginst8376 (P1_U7648, P1_STATE_REG_1__SCAN_IN, P1_STATE_REG_0__SCAN_IN);
  nand ginst8377 (P1_U7649, P1_STATE_REG_0__SCAN_IN, P1_U4258);
  not ginst8378 (P1_U7650, P1_U3462);
  nand ginst8379 (P1_U7651, P1_DATAWIDTH_REG_0__SCAN_IN, P1_U7650);
  nand ginst8380 (P1_U7652, P1_U3462, P1_U3463);
  nand ginst8381 (P1_U7653, P1_U3462, P1_U4376);
  nand ginst8382 (P1_U7654, P1_DATAWIDTH_REG_1__SCAN_IN, P1_U7650);
  nand ginst8383 (P1_U7655, P1_U3265, P1_U3540, P1_U3541);
  nand ginst8384 (P1_U7656, P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN, P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN, P1_INSTQUEUE_REG_7__4__SCAN_IN, P1_U3270);
  nand ginst8385 (P1_U7657, P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN, P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN, P1_INSTQUEUE_REG_5__4__SCAN_IN, P1_U3265, P1_U3270);
  nand ginst8386 (P1_U7658, P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P1_INSTQUEUE_REG_2__4__SCAN_IN, P1_U3264, P1_U3266, P1_U3270);
  nand ginst8387 (P1_U7659, P1_U3270, P1_U3542, P1_U3543);
  nand ginst8388 (P1_U7660, P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P1_U3544, P1_U3545);
  nand ginst8389 (P1_U7661, P1_U3265, P1_U3546, P1_U3547);
  nand ginst8390 (P1_U7662, P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P1_U3548, P1_U3549);
  nand ginst8391 (P1_U7663, P1_U3266, P1_U3550, P1_U3551);
  nand ginst8392 (P1_U7664, P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN, P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN, P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P1_INSTQUEUE_REG_15__4__SCAN_IN);
  nand ginst8393 (P1_U7665, P1_INSTQUEUE_REG_0__4__SCAN_IN, P1_U3264, P1_U3265, P1_U3266, P1_U3270);
  nand ginst8394 (P1_U7666, P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P1_INSTQUEUE_REG_8__4__SCAN_IN, P1_U3264, P1_U3265, P1_U3266);
  nand ginst8395 (P1_U7667, P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P1_INSTQUEUE_REG_10__4__SCAN_IN, P1_U3264, P1_U3266);
  nand ginst8396 (P1_U7668, P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN, P1_U3552, P1_U3553);
  nand ginst8397 (P1_U7669, P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN, P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P1_INSTQUEUE_REG_3__4__SCAN_IN, P1_U3264, P1_U3270);
  nand ginst8398 (P1_U7670, P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN, P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P1_INSTQUEUE_REG_11__4__SCAN_IN, P1_U3264);
  nand ginst8399 (P1_U7671, P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN, P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P1_INSTQUEUE_REG_3__5__SCAN_IN, P1_U3264, P1_U3270);
  nand ginst8400 (P1_U7672, P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P1_U3528, P1_U3529);
  nand ginst8401 (P1_U7673, P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN, P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P1_INSTQUEUE_REG_9__6__SCAN_IN, P1_U3264, P1_U3265);
  nand ginst8402 (P1_U7674, P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P1_U3534, P1_U3535);
  nand ginst8403 (P1_U7675, P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P1_INSTQUEUE_REG_10__6__SCAN_IN, P1_U3264, P1_U3266);
  nand ginst8404 (P1_U7676, P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN, P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P1_INSTQUEUE_REG_11__6__SCAN_IN, P1_U3264);
  nand ginst8405 (P1_U7677, P1_INSTQUEUE_REG_0__6__SCAN_IN, P1_U3264, P1_U3265, P1_U3266, P1_U3270);
  nand ginst8406 (P1_U7678, P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P1_INSTQUEUE_REG_8__6__SCAN_IN, P1_U3264, P1_U3265, P1_U3266);
  nand ginst8407 (P1_U7679, P1_U3437, P1_U4494);
  nand ginst8408 (P1_U7680, P1_U3284, P1_U7501);
  nand ginst8409 (P1_U7681, P1_R2167_U17, P1_U4216);
  nand ginst8410 (P1_U7682, P1_U3273, P1_U4506);
  nand ginst8411 (P1_U7683, P1_STATE2_REG_0__SCAN_IN, P1_U4512);
  nand ginst8412 (P1_U7684, P1_U3294, P1_U4513);
  nand ginst8413 (P1_U7685, P1_STATE2_REG_3__SCAN_IN, P1_U3295);
  nand ginst8414 (P1_U7686, P1_U2428, P1_U4514);
  or ginst8415 (P1_U7687, P1_STATEBS16_REG_SCAN_IN, P1_STATE2_REG_0__SCAN_IN);
  nand ginst8416 (P1_U7688, P1_STATE2_REG_0__SCAN_IN, P1_U7469);
  nand ginst8417 (P1_U7689, P1_STATE2_REG_0__SCAN_IN, P1_U4522);
  nand ginst8418 (P1_U7690, P1_U3294, P1_U4521, P1_U7604);
  nand ginst8419 (P1_U7691, P1_R2144_U49, P1_U3313);
  nand ginst8420 (P1_U7692, P1_U3311, P1_U4528);
  not ginst8421 (P1_U7693, P1_U3454);
  nand ginst8422 (P1_U7694, P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN, P1_U3305);
  nand ginst8423 (P1_U7695, P1_U3304, P1_U4533);
  not ginst8424 (P1_U7696, P1_U3455);
  nand ginst8425 (P1_U7697, P1_U3273, P1_U4216);
  nand ginst8426 (P1_U7698, P1_R2167_U17, P1_U7497);
  nand ginst8427 (P1_U7699, P1_U4432, P1_U5466);
  nand ginst8428 (P1_U7700, P1_U4171, P1_U5467);
  nand ginst8429 (P1_U7701, P1_U3467, P1_U4172);
  nand ginst8430 (P1_U7702, P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN, P1_U5476);
  nand ginst8431 (P1_U7703, P1_U3278, P1_U4460);
  nand ginst8432 (P1_U7704, P1_U3277, P1_U4415);
  nand ginst8433 (P1_U7705, P1_U3271, P1_U3415);
  nand ginst8434 (P1_U7706, P1_U4477, P1_U5493);
  nand ginst8435 (P1_U7707, P1_U7705, P1_U7706);
  nand ginst8436 (P1_U7708, P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P1_U5476);
  nand ginst8437 (P1_U7709, P1_U4172, P1_U5509);
  nand ginst8438 (P1_U7710, P1_INSTADDRPOINTER_REG_1__SCAN_IN, P1_U4174);
  nand ginst8439 (P1_U7711, P1_INSTADDRPOINTER_REG_31__SCAN_IN, P1_SUB_580_U6);
  not ginst8440 (P1_U7712, P1_U3470);
  nand ginst8441 (P1_U7713, P1_INSTADDRPOINTER_REG_0__SCAN_IN, P1_U4174);
  nand ginst8442 (P1_U7714, P1_INSTADDRPOINTER_REG_31__SCAN_IN, P1_INSTADDRPOINTER_REG_0__SCAN_IN);
  not ginst8443 (P1_U7715, P1_U3471);
  nand ginst8444 (P1_U7716, P1_U5501, P1_U5511);
  nand ginst8445 (P1_U7717, P1_U3401, P1_U4218);
  nand ginst8446 (P1_U7718, P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P1_U3264);
  nand ginst8447 (P1_U7719, P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN, P1_U3265);
  not ginst8448 (P1_U7720, P1_U3456);
  nand ginst8449 (P1_U7721, P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN, P1_U5476);
  nand ginst8450 (P1_U7722, P1_U4172, P1_U5518);
  nand ginst8451 (P1_U7723, P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P1_U5476);
  nand ginst8452 (P1_U7724, P1_U4172, P1_U5529);
  nand ginst8453 (P1_U7725, P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN, P1_U4214);
  nand ginst8454 (P1_U7726, P1_U3266, P1_U5521);
  nand ginst8455 (P1_U7727, P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN, P1_U5476);
  nand ginst8456 (P1_U7728, P1_U4172, P1_U5535);
  nand ginst8457 (P1_U7729, P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN, P1_U5537);
  nand ginst8458 (P1_U7730, P1_U3404, P1_U5545);
  nand ginst8459 (P1_U7731, P1_U4527, P1_U7693);
  nand ginst8460 (P1_U7732, P1_U3314, P1_U3454);
  nand ginst8461 (P1_U7733, P1_U7731, P1_U7732);
  nand ginst8462 (P1_U7734, P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN, P1_U5537);
  nand ginst8463 (P1_U7735, P1_U3404, P1_U5549);
  nand ginst8464 (P1_U7736, P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN, P1_U5537);
  nand ginst8465 (P1_U7737, P1_U3404, P1_U5554);
  nand ginst8466 (P1_U7738, P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P1_U5537);
  nand ginst8467 (P1_U7739, P1_U3404, P1_U5557);
  nand ginst8468 (P1_U7740, P1_U3388, P1_U4477);
  nand ginst8469 (P1_U7741, P1_U3271, P1_U3281);
  nand ginst8470 (P1_U7742, P1_U3257, P1_U4171, P1_U7740, P1_U7741);
  nand ginst8471 (P1_U7743, P1_R2167_U17, P1_U4432, P1_U7611);
  nand ginst8472 (P1_U7744, P1_EAX_REG_31__SCAN_IN, P1_U3424);
  nand ginst8473 (P1_U7745, P1_U3479, P1_U4223);
  nand ginst8474 (P1_U7746, P1_BYTEENABLE_REG_3__SCAN_IN, P1_U3433);
  nand ginst8475 (P1_U7747, P1_U3480, P1_U4220);
  or ginst8476 (P1_U7748, P1_DATAWIDTH_REG_0__SCAN_IN, P1_DATAWIDTH_REG_1__SCAN_IN);
  nand ginst8477 (P1_U7749, P1_DATAWIDTH_REG_0__SCAN_IN, P1_U3413);
  nand ginst8478 (P1_U7750, P1_U7748, P1_U7749);
  nand ginst8479 (P1_U7751, P1_U3253, P1_U7750);
  nand ginst8480 (P1_U7752, P1_REIP_REG_1__SCAN_IN, P1_REIP_REG_0__SCAN_IN);
  nand ginst8481 (P1_U7753, P1_U7751, P1_U7752);
  nand ginst8482 (P1_U7754, P1_BYTEENABLE_REG_2__SCAN_IN, P1_U3433);
  nand ginst8483 (P1_U7755, P1_U4220, P1_U7753);
  nand ginst8484 (P1_U7756, P1_BYTEENABLE_REG_1__SCAN_IN, P1_U3433);
  nand ginst8485 (P1_U7757, P1_REIP_REG_1__SCAN_IN, P1_U4220);
  nand ginst8486 (P1_U7758, P1_BYTEENABLE_REG_0__SCAN_IN, P1_U3433);
  nand ginst8487 (P1_U7759, P1_U4220, P1_U6599);
  nand ginst8488 (P1_U7760, P1_U3436, P1_U4221);
  nand ginst8489 (P1_U7761, P1_W_R_N_REG_SCAN_IN, P1_U3249);
  nand ginst8490 (P1_U7762, P1_MORE_REG_SCAN_IN, P1_U4177);
  nand ginst8491 (P1_U7763, P1_U4237, P1_U6600);
  nand ginst8492 (P1_U7764, P1_STATEBS16_REG_SCAN_IN, P1_U7650);
  nand ginst8493 (P1_U7765, BS16, P1_U3462);
  nand ginst8494 (P1_U7766, P1_REQUESTPENDING_REG_SCAN_IN, P1_U6603);
  nand ginst8495 (P1_U7767, P1_U4180, P1_U6609);
  nand ginst8496 (P1_U7768, P1_U3435, P1_U4221);
  nand ginst8497 (P1_U7769, P1_D_C_N_REG_SCAN_IN, P1_U3249);
  nand ginst8498 (P1_U7770, P1_M_IO_N_REG_SCAN_IN, P1_U3249);
  nand ginst8499 (P1_U7771, P1_MEMORYFETCH_REG_SCAN_IN, P1_U4221);
  nand ginst8500 (P1_U7772, P1_READREQUEST_REG_SCAN_IN, P1_U6614);
  nand ginst8501 (P1_U7773, P1_U4181, P1_U6615);
  nand ginst8502 (P1_U7774, P1_U3488, P1_U4182);
  nand ginst8503 (P1_U7775, P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN, P1_U5473);
  nand ginst8504 (P1_U7776, P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P1_U5473);
  nand ginst8505 (P1_U7777, P1_U4182, P1_U5506);
  nand ginst8506 (P1_U7778, P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN, P1_U5473);
  nand ginst8507 (P1_U7779, P1_U4182, P1_U5514);
  nand ginst8508 (P1_U7780, P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P1_U5473);
  nand ginst8509 (P1_U7781, P1_U4182, P1_U5525);
  nand ginst8510 (P1_U7782, P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN, P1_U5473);
  nand ginst8511 (P1_U7783, P1_U4182, P1_U5531);
  nand ginst8512 (P1_U7784, P1_U2605, P1_U3277);
  nand ginst8513 (P1_U7785, P1_U4460, P1_U7495);
  nand ginst8514 (P1_U7786, P1_U3301, P1_U4203);
  nand ginst8515 (P1_U7787, P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P1_U3297);
  nand ginst8516 (P1_U7788, P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P1_U4183);
  nand ginst8517 (P1_U7789, P1_U3270, P1_U7219);
  not ginst8518 (P1_U7790, P1_U3457);
  nand ginst8519 (P1_U7791, P1_U3276, P1_U3284);
  nand ginst8520 (P1_U7792, P1_U4494, P1_U7707);
  nand ginst8521 (P1_U7793, P1_U3262, P1_U3493);
  nand ginst8522 (P1_U7794, P1_FLUSH_REG_SCAN_IN, P1_STATE2_REG_1__SCAN_IN, P1_U7715);
  and ginst8523 (P2_ADD_371_1212_U10, P2_INSTADDRPOINTER_REG_9__SCAN_IN, P2_INSTADDRPOINTER_REG_10__SCAN_IN, P2_INSTADDRPOINTER_REG_11__SCAN_IN, P2_INSTADDRPOINTER_REG_12__SCAN_IN);
  and ginst8524 (P2_ADD_371_1212_U100, P2_ADD_371_1212_U101, P2_ADD_371_1212_U7);
  and ginst8525 (P2_ADD_371_1212_U101, P2_INSTADDRPOINTER_REG_16__SCAN_IN, P2_INSTADDRPOINTER_REG_17__SCAN_IN);
  and ginst8526 (P2_ADD_371_1212_U102, P2_INSTADDRPOINTER_REG_11__SCAN_IN, P2_ADD_371_1212_U5);
  and ginst8527 (P2_ADD_371_1212_U103, P2_ADD_371_1212_U104, P2_ADD_371_1212_U9);
  and ginst8528 (P2_ADD_371_1212_U104, P2_INSTADDRPOINTER_REG_24__SCAN_IN, P2_INSTADDRPOINTER_REG_25__SCAN_IN);
  and ginst8529 (P2_ADD_371_1212_U105, P2_INSTADDRPOINTER_REG_14__SCAN_IN, P2_ADD_371_1212_U4);
  and ginst8530 (P2_ADD_371_1212_U106, P2_INSTADDRPOINTER_REG_30__SCAN_IN, P2_ADD_371_1212_U12);
  and ginst8531 (P2_ADD_371_1212_U107, P2_INSTADDRPOINTER_REG_30__SCAN_IN, P2_ADD_371_1212_U12);
  and ginst8532 (P2_ADD_371_1212_U108, P2_INSTADDRPOINTER_REG_27__SCAN_IN, P2_ADD_371_1212_U8);
  and ginst8533 (P2_ADD_371_1212_U109, P2_INSTADDRPOINTER_REG_24__SCAN_IN, P2_ADD_371_1212_U9);
  and ginst8534 (P2_ADD_371_1212_U11, P2_ADD_371_1212_U7, P2_ADD_371_1212_U88);
  and ginst8535 (P2_ADD_371_1212_U110, P2_ADD_371_1212_U207, P2_ADD_371_1212_U208);
  nand ginst8536 (P2_ADD_371_1212_U111, P2_ADD_371_1212_U154, P2_ADD_371_1212_U155);
  nand ginst8537 (P2_ADD_371_1212_U112, P2_ADD_371_1212_U117, P2_ADD_371_1212_U12);
  nand ginst8538 (P2_ADD_371_1212_U113, P2_ADD_371_1212_U117, P2_ADD_371_1212_U9);
  nand ginst8539 (P2_ADD_371_1212_U114, P2_ADD_371_1212_U117, P2_ADD_371_1212_U95);
  and ginst8540 (P2_ADD_371_1212_U115, P2_ADD_371_1212_U220, P2_ADD_371_1212_U221);
  nand ginst8541 (P2_ADD_371_1212_U116, P2_ADD_371_1212_U139, P2_ADD_371_1212_U67);
  nand ginst8542 (P2_ADD_371_1212_U117, P2_ADD_371_1212_U202, P2_ADD_371_1212_U86);
  and ginst8543 (P2_ADD_371_1212_U118, P2_ADD_371_1212_U227, P2_ADD_371_1212_U228);
  nand ginst8544 (P2_ADD_371_1212_U119, P2_ADD_371_1212_U100, P2_ADD_371_1212_U117);
  and ginst8545 (P2_ADD_371_1212_U12, P2_ADD_371_1212_U8, P2_ADD_371_1212_U92);
  nand ginst8546 (P2_ADD_371_1212_U120, P2_ADD_371_1212_U105, P2_ADD_371_1212_U117);
  and ginst8547 (P2_ADD_371_1212_U121, P2_ADD_371_1212_U233, P2_ADD_371_1212_U234);
  nand ginst8548 (P2_ADD_371_1212_U122, P2_ADD_371_1212_U146, P2_ADD_371_1212_U147);
  nand ginst8549 (P2_ADD_371_1212_U123, P2_ADD_371_1212_U117, P2_ADD_371_1212_U8);
  and ginst8550 (P2_ADD_371_1212_U124, P2_ADD_371_1212_U242, P2_ADD_371_1212_U243);
  nand ginst8551 (P2_ADD_371_1212_U125, P2_ADD_371_1212_U150, P2_ADD_371_1212_U151);
  and ginst8552 (P2_ADD_371_1212_U126, P2_ADD_371_1212_U249, P2_ADD_371_1212_U250);
  nand ginst8553 (P2_ADD_371_1212_U127, P2_ADD_371_1212_U162, P2_ADD_371_1212_U163);
  not ginst8554 (P2_ADD_371_1212_U128, P2_INSTADDRPOINTER_REG_31__SCAN_IN);
  and ginst8555 (P2_ADD_371_1212_U129, P2_ADD_371_1212_U258, P2_ADD_371_1212_U259);
  and ginst8556 (P2_ADD_371_1212_U13, P2_ADD_371_1212_U168, P2_ADD_371_1212_U196);
  nand ginst8557 (P2_ADD_371_1212_U130, P2_ADD_371_1212_U142, P2_ADD_371_1212_U143);
  nand ginst8558 (P2_ADD_371_1212_U131, P2_ADD_371_1212_U117, P2_ADD_371_1212_U6);
  nand ginst8559 (P2_ADD_371_1212_U132, P2_ADD_371_1212_U102, P2_ADD_371_1212_U117);
  and ginst8560 (P2_ADD_371_1212_U133, P2_ADD_371_1212_U274, P2_ADD_371_1212_U275);
  nand ginst8561 (P2_ADD_371_1212_U134, P2_ADD_371_1212_U158, P2_ADD_371_1212_U159);
  nand ginst8562 (P2_ADD_371_1212_U135, P2_ADD_371_1212_U109, P2_ADD_371_1212_U117);
  not ginst8563 (P2_ADD_371_1212_U136, P2_ADD_371_1212_U67);
  not ginst8564 (P2_ADD_371_1212_U137, P2_ADD_371_1212_U29);
  nand ginst8565 (P2_ADD_371_1212_U138, P2_ADD_371_1212_U29, P2_ADD_371_1212_U30);
  nand ginst8566 (P2_ADD_371_1212_U139, P2_INSTADDRPOINTER_REG_1__SCAN_IN, P2_ADD_371_1212_U138);
  and ginst8567 (P2_ADD_371_1212_U14, P2_ADD_371_1212_U132, P2_ADD_371_1212_U188);
  not ginst8568 (P2_ADD_371_1212_U140, P2_ADD_371_1212_U116);
  or ginst8569 (P2_ADD_371_1212_U141, P2_INSTADDRPOINTER_REG_2__SCAN_IN, P2_R2256_U22);
  nand ginst8570 (P2_ADD_371_1212_U142, P2_ADD_371_1212_U116, P2_ADD_371_1212_U141);
  nand ginst8571 (P2_ADD_371_1212_U143, P2_INSTADDRPOINTER_REG_2__SCAN_IN, P2_R2256_U22);
  not ginst8572 (P2_ADD_371_1212_U144, P2_ADD_371_1212_U130);
  or ginst8573 (P2_ADD_371_1212_U145, P2_INSTADDRPOINTER_REG_3__SCAN_IN, P2_R2256_U26);
  nand ginst8574 (P2_ADD_371_1212_U146, P2_ADD_371_1212_U130, P2_ADD_371_1212_U145);
  nand ginst8575 (P2_ADD_371_1212_U147, P2_INSTADDRPOINTER_REG_3__SCAN_IN, P2_R2256_U26);
  not ginst8576 (P2_ADD_371_1212_U148, P2_ADD_371_1212_U122);
  or ginst8577 (P2_ADD_371_1212_U149, P2_INSTADDRPOINTER_REG_4__SCAN_IN, P2_R2256_U20);
  and ginst8578 (P2_ADD_371_1212_U15, P2_ADD_371_1212_U170, P2_ADD_371_1212_U185);
  nand ginst8579 (P2_ADD_371_1212_U150, P2_ADD_371_1212_U122, P2_ADD_371_1212_U149);
  nand ginst8580 (P2_ADD_371_1212_U151, P2_INSTADDRPOINTER_REG_4__SCAN_IN, P2_R2256_U20);
  not ginst8581 (P2_ADD_371_1212_U152, P2_ADD_371_1212_U125);
  or ginst8582 (P2_ADD_371_1212_U153, P2_INSTADDRPOINTER_REG_5__SCAN_IN, P2_R2256_U19);
  nand ginst8583 (P2_ADD_371_1212_U154, P2_ADD_371_1212_U125, P2_ADD_371_1212_U153);
  nand ginst8584 (P2_ADD_371_1212_U155, P2_INSTADDRPOINTER_REG_5__SCAN_IN, P2_R2256_U19);
  not ginst8585 (P2_ADD_371_1212_U156, P2_ADD_371_1212_U111);
  or ginst8586 (P2_ADD_371_1212_U157, P2_INSTADDRPOINTER_REG_6__SCAN_IN, P2_R2256_U18);
  nand ginst8587 (P2_ADD_371_1212_U158, P2_ADD_371_1212_U111, P2_ADD_371_1212_U157);
  nand ginst8588 (P2_ADD_371_1212_U159, P2_INSTADDRPOINTER_REG_6__SCAN_IN, P2_R2256_U18);
  and ginst8589 (P2_ADD_371_1212_U16, P2_ADD_371_1212_U120, P2_ADD_371_1212_U191);
  not ginst8590 (P2_ADD_371_1212_U160, P2_ADD_371_1212_U134);
  or ginst8591 (P2_ADD_371_1212_U161, P2_INSTADDRPOINTER_REG_7__SCAN_IN, P2_R2256_U17);
  nand ginst8592 (P2_ADD_371_1212_U162, P2_ADD_371_1212_U134, P2_ADD_371_1212_U161);
  nand ginst8593 (P2_ADD_371_1212_U163, P2_INSTADDRPOINTER_REG_7__SCAN_IN, P2_R2256_U17);
  not ginst8594 (P2_ADD_371_1212_U164, P2_ADD_371_1212_U127);
  or ginst8595 (P2_ADD_371_1212_U165, P2_INSTADDRPOINTER_REG_8__SCAN_IN, P2_R2256_U5);
  nand ginst8596 (P2_ADD_371_1212_U166, P2_INSTADDRPOINTER_REG_8__SCAN_IN, P2_R2256_U5);
  not ginst8597 (P2_ADD_371_1212_U167, P2_ADD_371_1212_U117);
  nand ginst8598 (P2_ADD_371_1212_U168, P2_ADD_371_1212_U117, P2_ADD_371_1212_U5);
  not ginst8599 (P2_ADD_371_1212_U169, P2_ADD_371_1212_U132);
  and ginst8600 (P2_ADD_371_1212_U17, P2_ADD_371_1212_U114, P2_ADD_371_1212_U200);
  nand ginst8601 (P2_ADD_371_1212_U170, P2_ADD_371_1212_U117, P2_ADD_371_1212_U4);
  not ginst8602 (P2_ADD_371_1212_U171, P2_ADD_371_1212_U120);
  not ginst8603 (P2_ADD_371_1212_U172, P2_ADD_371_1212_U114);
  not ginst8604 (P2_ADD_371_1212_U173, P2_ADD_371_1212_U119);
  nand ginst8605 (P2_ADD_371_1212_U174, P2_ADD_371_1212_U117, P2_ADD_371_1212_U96);
  not ginst8606 (P2_ADD_371_1212_U175, P2_ADD_371_1212_U131);
  nand ginst8607 (P2_ADD_371_1212_U176, P2_ADD_371_1212_U117, P2_ADD_371_1212_U97);
  not ginst8608 (P2_ADD_371_1212_U177, P2_ADD_371_1212_U113);
  not ginst8609 (P2_ADD_371_1212_U178, P2_ADD_371_1212_U135);
  not ginst8610 (P2_ADD_371_1212_U179, P2_ADD_371_1212_U123);
  and ginst8611 (P2_ADD_371_1212_U18, P2_ADD_371_1212_U174, P2_ADD_371_1212_U194);
  nand ginst8612 (P2_ADD_371_1212_U180, P2_ADD_371_1212_U117, P2_ADD_371_1212_U93);
  not ginst8613 (P2_ADD_371_1212_U181, P2_ADD_371_1212_U112);
  nand ginst8614 (P2_ADD_371_1212_U182, P2_ADD_371_1212_U180, P2_ADD_371_1212_U65);
  nand ginst8615 (P2_ADD_371_1212_U183, P2_ADD_371_1212_U174, P2_ADD_371_1212_U56);
  nand ginst8616 (P2_ADD_371_1212_U184, P2_ADD_371_1212_U10, P2_ADD_371_1212_U117);
  nand ginst8617 (P2_ADD_371_1212_U185, P2_ADD_371_1212_U184, P2_ADD_371_1212_U49);
  nand ginst8618 (P2_ADD_371_1212_U186, P2_ADD_371_1212_U117, P2_ADD_371_1212_U99);
  nand ginst8619 (P2_ADD_371_1212_U187, P2_ADD_371_1212_U186, P2_ADD_371_1212_U58);
  nand ginst8620 (P2_ADD_371_1212_U188, P2_ADD_371_1212_U168, P2_ADD_371_1212_U47);
  nand ginst8621 (P2_ADD_371_1212_U189, P2_ADD_371_1212_U103, P2_ADD_371_1212_U117);
  and ginst8622 (P2_ADD_371_1212_U19, P2_ADD_371_1212_U131, P2_ADD_371_1212_U183);
  nand ginst8623 (P2_ADD_371_1212_U190, P2_ADD_371_1212_U189, P2_ADD_371_1212_U61);
  nand ginst8624 (P2_ADD_371_1212_U191, P2_ADD_371_1212_U170, P2_ADD_371_1212_U50);
  nand ginst8625 (P2_ADD_371_1212_U192, P2_ADD_371_1212_U176, P2_ADD_371_1212_U59);
  nand ginst8626 (P2_ADD_371_1212_U193, P2_ADD_371_1212_U11, P2_ADD_371_1212_U117);
  nand ginst8627 (P2_ADD_371_1212_U194, P2_ADD_371_1212_U193, P2_ADD_371_1212_U55);
  nand ginst8628 (P2_ADD_371_1212_U195, P2_INSTADDRPOINTER_REG_9__SCAN_IN, P2_ADD_371_1212_U117);
  nand ginst8629 (P2_ADD_371_1212_U196, P2_ADD_371_1212_U195, P2_ADD_371_1212_U46);
  nand ginst8630 (P2_ADD_371_1212_U197, P2_ADD_371_1212_U108, P2_ADD_371_1212_U117);
  nand ginst8631 (P2_ADD_371_1212_U198, P2_ADD_371_1212_U197, P2_ADD_371_1212_U64);
  nand ginst8632 (P2_ADD_371_1212_U199, P2_ADD_371_1212_U117, P2_ADD_371_1212_U7);
  and ginst8633 (P2_ADD_371_1212_U20, P2_ADD_371_1212_U176, P2_ADD_371_1212_U187);
  nand ginst8634 (P2_ADD_371_1212_U200, P2_ADD_371_1212_U199, P2_ADD_371_1212_U52);
  nand ginst8635 (P2_ADD_371_1212_U201, P2_ADD_371_1212_U107, P2_ADD_371_1212_U117);
  nand ginst8636 (P2_ADD_371_1212_U202, P2_ADD_371_1212_U134, P2_ADD_371_1212_U161, P2_ADD_371_1212_U165);
  nand ginst8637 (P2_ADD_371_1212_U203, P2_INSTADDRPOINTER_REG_7__SCAN_IN, P2_ADD_371_1212_U165, P2_R2256_U17);
  nand ginst8638 (P2_ADD_371_1212_U204, P2_INSTADDRPOINTER_REG_1__SCAN_IN, P2_ADD_371_1212_U136);
  nand ginst8639 (P2_ADD_371_1212_U205, P2_INSTADDRPOINTER_REG_0__SCAN_IN, P2_ADD_371_1212_U27);
  nand ginst8640 (P2_ADD_371_1212_U206, P2_ADD_371_1212_U26, P2_R2256_U21);
  nand ginst8641 (P2_ADD_371_1212_U207, P2_INSTADDRPOINTER_REG_6__SCAN_IN, P2_ADD_371_1212_U40);
  nand ginst8642 (P2_ADD_371_1212_U208, P2_ADD_371_1212_U39, P2_R2256_U18);
  nand ginst8643 (P2_ADD_371_1212_U209, P2_INSTADDRPOINTER_REG_6__SCAN_IN, P2_ADD_371_1212_U40);
  and ginst8644 (P2_ADD_371_1212_U21, P2_ADD_371_1212_U113, P2_ADD_371_1212_U192);
  nand ginst8645 (P2_ADD_371_1212_U210, P2_ADD_371_1212_U39, P2_R2256_U18);
  nand ginst8646 (P2_ADD_371_1212_U211, P2_ADD_371_1212_U209, P2_ADD_371_1212_U210);
  nand ginst8647 (P2_ADD_371_1212_U212, P2_ADD_371_1212_U110, P2_ADD_371_1212_U111);
  nand ginst8648 (P2_ADD_371_1212_U213, P2_ADD_371_1212_U156, P2_ADD_371_1212_U211);
  nand ginst8649 (P2_ADD_371_1212_U214, P2_INSTADDRPOINTER_REG_30__SCAN_IN, P2_ADD_371_1212_U112);
  nand ginst8650 (P2_ADD_371_1212_U215, P2_ADD_371_1212_U181, P2_ADD_371_1212_U66);
  nand ginst8651 (P2_ADD_371_1212_U216, P2_INSTADDRPOINTER_REG_24__SCAN_IN, P2_ADD_371_1212_U113);
  nand ginst8652 (P2_ADD_371_1212_U217, P2_ADD_371_1212_U177, P2_ADD_371_1212_U60);
  nand ginst8653 (P2_ADD_371_1212_U218, P2_INSTADDRPOINTER_REG_17__SCAN_IN, P2_ADD_371_1212_U114);
  nand ginst8654 (P2_ADD_371_1212_U219, P2_ADD_371_1212_U172, P2_ADD_371_1212_U54);
  and ginst8655 (P2_ADD_371_1212_U22, P2_ADD_371_1212_U123, P2_ADD_371_1212_U190);
  nand ginst8656 (P2_ADD_371_1212_U220, P2_INSTADDRPOINTER_REG_2__SCAN_IN, P2_ADD_371_1212_U31);
  nand ginst8657 (P2_ADD_371_1212_U221, P2_ADD_371_1212_U32, P2_R2256_U22);
  nand ginst8658 (P2_ADD_371_1212_U222, P2_INSTADDRPOINTER_REG_2__SCAN_IN, P2_ADD_371_1212_U31);
  nand ginst8659 (P2_ADD_371_1212_U223, P2_ADD_371_1212_U32, P2_R2256_U22);
  nand ginst8660 (P2_ADD_371_1212_U224, P2_ADD_371_1212_U222, P2_ADD_371_1212_U223);
  nand ginst8661 (P2_ADD_371_1212_U225, P2_ADD_371_1212_U115, P2_ADD_371_1212_U116);
  nand ginst8662 (P2_ADD_371_1212_U226, P2_ADD_371_1212_U140, P2_ADD_371_1212_U224);
  nand ginst8663 (P2_ADD_371_1212_U227, P2_INSTADDRPOINTER_REG_9__SCAN_IN, P2_ADD_371_1212_U117);
  nand ginst8664 (P2_ADD_371_1212_U228, P2_ADD_371_1212_U167, P2_ADD_371_1212_U45);
  nand ginst8665 (P2_ADD_371_1212_U229, P2_INSTADDRPOINTER_REG_18__SCAN_IN, P2_ADD_371_1212_U119);
  and ginst8666 (P2_ADD_371_1212_U23, P2_ADD_371_1212_U180, P2_ADD_371_1212_U198);
  nand ginst8667 (P2_ADD_371_1212_U230, P2_ADD_371_1212_U173, P2_ADD_371_1212_U53);
  nand ginst8668 (P2_ADD_371_1212_U231, P2_INSTADDRPOINTER_REG_15__SCAN_IN, P2_ADD_371_1212_U120);
  nand ginst8669 (P2_ADD_371_1212_U232, P2_ADD_371_1212_U171, P2_ADD_371_1212_U51);
  nand ginst8670 (P2_ADD_371_1212_U233, P2_INSTADDRPOINTER_REG_4__SCAN_IN, P2_ADD_371_1212_U35);
  nand ginst8671 (P2_ADD_371_1212_U234, P2_ADD_371_1212_U36, P2_R2256_U20);
  nand ginst8672 (P2_ADD_371_1212_U235, P2_INSTADDRPOINTER_REG_4__SCAN_IN, P2_ADD_371_1212_U35);
  nand ginst8673 (P2_ADD_371_1212_U236, P2_ADD_371_1212_U36, P2_R2256_U20);
  nand ginst8674 (P2_ADD_371_1212_U237, P2_ADD_371_1212_U235, P2_ADD_371_1212_U236);
  nand ginst8675 (P2_ADD_371_1212_U238, P2_ADD_371_1212_U121, P2_ADD_371_1212_U122);
  nand ginst8676 (P2_ADD_371_1212_U239, P2_ADD_371_1212_U148, P2_ADD_371_1212_U237);
  and ginst8677 (P2_ADD_371_1212_U24, P2_ADD_371_1212_U112, P2_ADD_371_1212_U182);
  nand ginst8678 (P2_ADD_371_1212_U240, P2_INSTADDRPOINTER_REG_27__SCAN_IN, P2_ADD_371_1212_U123);
  nand ginst8679 (P2_ADD_371_1212_U241, P2_ADD_371_1212_U179, P2_ADD_371_1212_U63);
  nand ginst8680 (P2_ADD_371_1212_U242, P2_INSTADDRPOINTER_REG_5__SCAN_IN, P2_ADD_371_1212_U37);
  nand ginst8681 (P2_ADD_371_1212_U243, P2_ADD_371_1212_U38, P2_R2256_U19);
  nand ginst8682 (P2_ADD_371_1212_U244, P2_INSTADDRPOINTER_REG_5__SCAN_IN, P2_ADD_371_1212_U37);
  nand ginst8683 (P2_ADD_371_1212_U245, P2_ADD_371_1212_U38, P2_R2256_U19);
  nand ginst8684 (P2_ADD_371_1212_U246, P2_ADD_371_1212_U244, P2_ADD_371_1212_U245);
  nand ginst8685 (P2_ADD_371_1212_U247, P2_ADD_371_1212_U124, P2_ADD_371_1212_U125);
  nand ginst8686 (P2_ADD_371_1212_U248, P2_ADD_371_1212_U152, P2_ADD_371_1212_U246);
  nand ginst8687 (P2_ADD_371_1212_U249, P2_INSTADDRPOINTER_REG_8__SCAN_IN, P2_ADD_371_1212_U41);
  nand ginst8688 (P2_ADD_371_1212_U25, P2_ADD_371_1212_U204, P2_ADD_371_1212_U268, P2_ADD_371_1212_U269);
  nand ginst8689 (P2_ADD_371_1212_U250, P2_ADD_371_1212_U42, P2_R2256_U5);
  nand ginst8690 (P2_ADD_371_1212_U251, P2_INSTADDRPOINTER_REG_8__SCAN_IN, P2_ADD_371_1212_U41);
  nand ginst8691 (P2_ADD_371_1212_U252, P2_ADD_371_1212_U42, P2_R2256_U5);
  nand ginst8692 (P2_ADD_371_1212_U253, P2_ADD_371_1212_U251, P2_ADD_371_1212_U252);
  nand ginst8693 (P2_ADD_371_1212_U254, P2_ADD_371_1212_U126, P2_ADD_371_1212_U127);
  nand ginst8694 (P2_ADD_371_1212_U255, P2_ADD_371_1212_U164, P2_ADD_371_1212_U253);
  nand ginst8695 (P2_ADD_371_1212_U256, P2_INSTADDRPOINTER_REG_31__SCAN_IN, P2_ADD_371_1212_U201);
  nand ginst8696 (P2_ADD_371_1212_U257, P2_ADD_371_1212_U106, P2_ADD_371_1212_U117, P2_ADD_371_1212_U128);
  nand ginst8697 (P2_ADD_371_1212_U258, P2_INSTADDRPOINTER_REG_3__SCAN_IN, P2_ADD_371_1212_U33);
  nand ginst8698 (P2_ADD_371_1212_U259, P2_ADD_371_1212_U34, P2_R2256_U26);
  not ginst8699 (P2_ADD_371_1212_U26, P2_INSTADDRPOINTER_REG_0__SCAN_IN);
  nand ginst8700 (P2_ADD_371_1212_U260, P2_INSTADDRPOINTER_REG_3__SCAN_IN, P2_ADD_371_1212_U33);
  nand ginst8701 (P2_ADD_371_1212_U261, P2_ADD_371_1212_U34, P2_R2256_U26);
  nand ginst8702 (P2_ADD_371_1212_U262, P2_ADD_371_1212_U260, P2_ADD_371_1212_U261);
  nand ginst8703 (P2_ADD_371_1212_U263, P2_ADD_371_1212_U129, P2_ADD_371_1212_U130);
  nand ginst8704 (P2_ADD_371_1212_U264, P2_ADD_371_1212_U144, P2_ADD_371_1212_U262);
  nand ginst8705 (P2_ADD_371_1212_U265, P2_INSTADDRPOINTER_REG_1__SCAN_IN, P2_ADD_371_1212_U29);
  nand ginst8706 (P2_ADD_371_1212_U266, P2_ADD_371_1212_U137, P2_ADD_371_1212_U28);
  nand ginst8707 (P2_ADD_371_1212_U267, P2_ADD_371_1212_U265, P2_ADD_371_1212_U266);
  nand ginst8708 (P2_ADD_371_1212_U268, P2_ADD_371_1212_U28, P2_ADD_371_1212_U29, P2_R2256_U4);
  nand ginst8709 (P2_ADD_371_1212_U269, P2_ADD_371_1212_U267, P2_ADD_371_1212_U30);
  not ginst8710 (P2_ADD_371_1212_U27, P2_R2256_U21);
  nand ginst8711 (P2_ADD_371_1212_U270, P2_INSTADDRPOINTER_REG_21__SCAN_IN, P2_ADD_371_1212_U131);
  nand ginst8712 (P2_ADD_371_1212_U271, P2_ADD_371_1212_U175, P2_ADD_371_1212_U57);
  nand ginst8713 (P2_ADD_371_1212_U272, P2_INSTADDRPOINTER_REG_12__SCAN_IN, P2_ADD_371_1212_U132);
  nand ginst8714 (P2_ADD_371_1212_U273, P2_ADD_371_1212_U169, P2_ADD_371_1212_U48);
  nand ginst8715 (P2_ADD_371_1212_U274, P2_INSTADDRPOINTER_REG_7__SCAN_IN, P2_ADD_371_1212_U43);
  nand ginst8716 (P2_ADD_371_1212_U275, P2_ADD_371_1212_U44, P2_R2256_U17);
  nand ginst8717 (P2_ADD_371_1212_U276, P2_INSTADDRPOINTER_REG_7__SCAN_IN, P2_ADD_371_1212_U43);
  nand ginst8718 (P2_ADD_371_1212_U277, P2_ADD_371_1212_U44, P2_R2256_U17);
  nand ginst8719 (P2_ADD_371_1212_U278, P2_ADD_371_1212_U276, P2_ADD_371_1212_U277);
  nand ginst8720 (P2_ADD_371_1212_U279, P2_ADD_371_1212_U133, P2_ADD_371_1212_U134);
  not ginst8721 (P2_ADD_371_1212_U28, P2_INSTADDRPOINTER_REG_1__SCAN_IN);
  nand ginst8722 (P2_ADD_371_1212_U280, P2_ADD_371_1212_U160, P2_ADD_371_1212_U278);
  nand ginst8723 (P2_ADD_371_1212_U281, P2_INSTADDRPOINTER_REG_25__SCAN_IN, P2_ADD_371_1212_U135);
  nand ginst8724 (P2_ADD_371_1212_U282, P2_ADD_371_1212_U178, P2_ADD_371_1212_U62);
  nand ginst8725 (P2_ADD_371_1212_U29, P2_INSTADDRPOINTER_REG_0__SCAN_IN, P2_R2256_U21);
  not ginst8726 (P2_ADD_371_1212_U30, P2_R2256_U4);
  not ginst8727 (P2_ADD_371_1212_U31, P2_R2256_U22);
  not ginst8728 (P2_ADD_371_1212_U32, P2_INSTADDRPOINTER_REG_2__SCAN_IN);
  not ginst8729 (P2_ADD_371_1212_U33, P2_R2256_U26);
  not ginst8730 (P2_ADD_371_1212_U34, P2_INSTADDRPOINTER_REG_3__SCAN_IN);
  not ginst8731 (P2_ADD_371_1212_U35, P2_R2256_U20);
  not ginst8732 (P2_ADD_371_1212_U36, P2_INSTADDRPOINTER_REG_4__SCAN_IN);
  not ginst8733 (P2_ADD_371_1212_U37, P2_R2256_U19);
  not ginst8734 (P2_ADD_371_1212_U38, P2_INSTADDRPOINTER_REG_5__SCAN_IN);
  not ginst8735 (P2_ADD_371_1212_U39, P2_INSTADDRPOINTER_REG_6__SCAN_IN);
  and ginst8736 (P2_ADD_371_1212_U4, P2_INSTADDRPOINTER_REG_13__SCAN_IN, P2_ADD_371_1212_U10);
  not ginst8737 (P2_ADD_371_1212_U40, P2_R2256_U18);
  not ginst8738 (P2_ADD_371_1212_U41, P2_R2256_U5);
  not ginst8739 (P2_ADD_371_1212_U42, P2_INSTADDRPOINTER_REG_8__SCAN_IN);
  not ginst8740 (P2_ADD_371_1212_U43, P2_R2256_U17);
  not ginst8741 (P2_ADD_371_1212_U44, P2_INSTADDRPOINTER_REG_7__SCAN_IN);
  not ginst8742 (P2_ADD_371_1212_U45, P2_INSTADDRPOINTER_REG_9__SCAN_IN);
  not ginst8743 (P2_ADD_371_1212_U46, P2_INSTADDRPOINTER_REG_10__SCAN_IN);
  not ginst8744 (P2_ADD_371_1212_U47, P2_INSTADDRPOINTER_REG_11__SCAN_IN);
  not ginst8745 (P2_ADD_371_1212_U48, P2_INSTADDRPOINTER_REG_12__SCAN_IN);
  not ginst8746 (P2_ADD_371_1212_U49, P2_INSTADDRPOINTER_REG_13__SCAN_IN);
  and ginst8747 (P2_ADD_371_1212_U5, P2_INSTADDRPOINTER_REG_9__SCAN_IN, P2_INSTADDRPOINTER_REG_10__SCAN_IN);
  not ginst8748 (P2_ADD_371_1212_U50, P2_INSTADDRPOINTER_REG_14__SCAN_IN);
  not ginst8749 (P2_ADD_371_1212_U51, P2_INSTADDRPOINTER_REG_15__SCAN_IN);
  not ginst8750 (P2_ADD_371_1212_U52, P2_INSTADDRPOINTER_REG_16__SCAN_IN);
  not ginst8751 (P2_ADD_371_1212_U53, P2_INSTADDRPOINTER_REG_18__SCAN_IN);
  not ginst8752 (P2_ADD_371_1212_U54, P2_INSTADDRPOINTER_REG_17__SCAN_IN);
  not ginst8753 (P2_ADD_371_1212_U55, P2_INSTADDRPOINTER_REG_19__SCAN_IN);
  not ginst8754 (P2_ADD_371_1212_U56, P2_INSTADDRPOINTER_REG_20__SCAN_IN);
  not ginst8755 (P2_ADD_371_1212_U57, P2_INSTADDRPOINTER_REG_21__SCAN_IN);
  not ginst8756 (P2_ADD_371_1212_U58, P2_INSTADDRPOINTER_REG_22__SCAN_IN);
  not ginst8757 (P2_ADD_371_1212_U59, P2_INSTADDRPOINTER_REG_23__SCAN_IN);
  and ginst8758 (P2_ADD_371_1212_U6, P2_ADD_371_1212_U11, P2_ADD_371_1212_U89);
  not ginst8759 (P2_ADD_371_1212_U60, P2_INSTADDRPOINTER_REG_24__SCAN_IN);
  not ginst8760 (P2_ADD_371_1212_U61, P2_INSTADDRPOINTER_REG_26__SCAN_IN);
  not ginst8761 (P2_ADD_371_1212_U62, P2_INSTADDRPOINTER_REG_25__SCAN_IN);
  not ginst8762 (P2_ADD_371_1212_U63, P2_INSTADDRPOINTER_REG_27__SCAN_IN);
  not ginst8763 (P2_ADD_371_1212_U64, P2_INSTADDRPOINTER_REG_28__SCAN_IN);
  not ginst8764 (P2_ADD_371_1212_U65, P2_INSTADDRPOINTER_REG_29__SCAN_IN);
  not ginst8765 (P2_ADD_371_1212_U66, P2_INSTADDRPOINTER_REG_30__SCAN_IN);
  nand ginst8766 (P2_ADD_371_1212_U67, P2_ADD_371_1212_U137, P2_R2256_U4);
  nand ginst8767 (P2_ADD_371_1212_U68, P2_ADD_371_1212_U205, P2_ADD_371_1212_U206);
  nand ginst8768 (P2_ADD_371_1212_U69, P2_ADD_371_1212_U214, P2_ADD_371_1212_U215);
  and ginst8769 (P2_ADD_371_1212_U7, P2_ADD_371_1212_U10, P2_ADD_371_1212_U87);
  nand ginst8770 (P2_ADD_371_1212_U70, P2_ADD_371_1212_U216, P2_ADD_371_1212_U217);
  nand ginst8771 (P2_ADD_371_1212_U71, P2_ADD_371_1212_U218, P2_ADD_371_1212_U219);
  nand ginst8772 (P2_ADD_371_1212_U72, P2_ADD_371_1212_U229, P2_ADD_371_1212_U230);
  nand ginst8773 (P2_ADD_371_1212_U73, P2_ADD_371_1212_U231, P2_ADD_371_1212_U232);
  nand ginst8774 (P2_ADD_371_1212_U74, P2_ADD_371_1212_U240, P2_ADD_371_1212_U241);
  nand ginst8775 (P2_ADD_371_1212_U75, P2_ADD_371_1212_U270, P2_ADD_371_1212_U271);
  nand ginst8776 (P2_ADD_371_1212_U76, P2_ADD_371_1212_U272, P2_ADD_371_1212_U273);
  nand ginst8777 (P2_ADD_371_1212_U77, P2_ADD_371_1212_U281, P2_ADD_371_1212_U282);
  nand ginst8778 (P2_ADD_371_1212_U78, P2_ADD_371_1212_U212, P2_ADD_371_1212_U213);
  nand ginst8779 (P2_ADD_371_1212_U79, P2_ADD_371_1212_U225, P2_ADD_371_1212_U226);
  and ginst8780 (P2_ADD_371_1212_U8, P2_ADD_371_1212_U9, P2_ADD_371_1212_U91);
  nand ginst8781 (P2_ADD_371_1212_U80, P2_ADD_371_1212_U238, P2_ADD_371_1212_U239);
  nand ginst8782 (P2_ADD_371_1212_U81, P2_ADD_371_1212_U247, P2_ADD_371_1212_U248);
  nand ginst8783 (P2_ADD_371_1212_U82, P2_ADD_371_1212_U254, P2_ADD_371_1212_U255);
  nand ginst8784 (P2_ADD_371_1212_U83, P2_ADD_371_1212_U256, P2_ADD_371_1212_U257);
  nand ginst8785 (P2_ADD_371_1212_U84, P2_ADD_371_1212_U263, P2_ADD_371_1212_U264);
  nand ginst8786 (P2_ADD_371_1212_U85, P2_ADD_371_1212_U279, P2_ADD_371_1212_U280);
  and ginst8787 (P2_ADD_371_1212_U86, P2_ADD_371_1212_U166, P2_ADD_371_1212_U203);
  and ginst8788 (P2_ADD_371_1212_U87, P2_INSTADDRPOINTER_REG_13__SCAN_IN, P2_INSTADDRPOINTER_REG_14__SCAN_IN, P2_INSTADDRPOINTER_REG_15__SCAN_IN);
  and ginst8789 (P2_ADD_371_1212_U88, P2_INSTADDRPOINTER_REG_16__SCAN_IN, P2_INSTADDRPOINTER_REG_17__SCAN_IN, P2_INSTADDRPOINTER_REG_18__SCAN_IN);
  and ginst8790 (P2_ADD_371_1212_U89, P2_INSTADDRPOINTER_REG_19__SCAN_IN, P2_INSTADDRPOINTER_REG_20__SCAN_IN);
  and ginst8791 (P2_ADD_371_1212_U9, P2_ADD_371_1212_U6, P2_ADD_371_1212_U90);
  and ginst8792 (P2_ADD_371_1212_U90, P2_INSTADDRPOINTER_REG_21__SCAN_IN, P2_INSTADDRPOINTER_REG_22__SCAN_IN, P2_INSTADDRPOINTER_REG_23__SCAN_IN);
  and ginst8793 (P2_ADD_371_1212_U91, P2_INSTADDRPOINTER_REG_24__SCAN_IN, P2_INSTADDRPOINTER_REG_25__SCAN_IN, P2_INSTADDRPOINTER_REG_26__SCAN_IN);
  and ginst8794 (P2_ADD_371_1212_U92, P2_INSTADDRPOINTER_REG_27__SCAN_IN, P2_INSTADDRPOINTER_REG_28__SCAN_IN, P2_INSTADDRPOINTER_REG_29__SCAN_IN);
  and ginst8795 (P2_ADD_371_1212_U93, P2_ADD_371_1212_U8, P2_ADD_371_1212_U94);
  and ginst8796 (P2_ADD_371_1212_U94, P2_INSTADDRPOINTER_REG_27__SCAN_IN, P2_INSTADDRPOINTER_REG_28__SCAN_IN);
  and ginst8797 (P2_ADD_371_1212_U95, P2_INSTADDRPOINTER_REG_16__SCAN_IN, P2_ADD_371_1212_U7);
  and ginst8798 (P2_ADD_371_1212_U96, P2_INSTADDRPOINTER_REG_19__SCAN_IN, P2_ADD_371_1212_U11);
  and ginst8799 (P2_ADD_371_1212_U97, P2_ADD_371_1212_U6, P2_ADD_371_1212_U98);
  and ginst8800 (P2_ADD_371_1212_U98, P2_INSTADDRPOINTER_REG_21__SCAN_IN, P2_INSTADDRPOINTER_REG_22__SCAN_IN);
  and ginst8801 (P2_ADD_371_1212_U99, P2_INSTADDRPOINTER_REG_21__SCAN_IN, P2_ADD_371_1212_U6);
  and ginst8802 (P2_ADD_391_1196_U10, P2_ADD_391_1196_U199, P2_ADD_391_1196_U201);
  nand ginst8803 (P2_ADD_391_1196_U100, P2_ADD_391_1196_U405, P2_ADD_391_1196_U406);
  nand ginst8804 (P2_ADD_391_1196_U101, P2_ADD_391_1196_U412, P2_ADD_391_1196_U413);
  nand ginst8805 (P2_ADD_391_1196_U102, P2_ADD_391_1196_U419, P2_ADD_391_1196_U420);
  nand ginst8806 (P2_ADD_391_1196_U103, P2_ADD_391_1196_U431, P2_ADD_391_1196_U432);
  nand ginst8807 (P2_ADD_391_1196_U104, P2_ADD_391_1196_U438, P2_ADD_391_1196_U439);
  nand ginst8808 (P2_ADD_391_1196_U105, P2_ADD_391_1196_U445, P2_ADD_391_1196_U446);
  nand ginst8809 (P2_ADD_391_1196_U106, P2_ADD_391_1196_U452, P2_ADD_391_1196_U453);
  nand ginst8810 (P2_ADD_391_1196_U107, P2_ADD_391_1196_U459, P2_ADD_391_1196_U460);
  nand ginst8811 (P2_ADD_391_1196_U108, P2_ADD_391_1196_U468, P2_ADD_391_1196_U469);
  nand ginst8812 (P2_ADD_391_1196_U109, P2_ADD_391_1196_U475, P2_ADD_391_1196_U476);
  and ginst8813 (P2_ADD_391_1196_U11, P2_ADD_391_1196_U192, P2_ADD_391_1196_U196);
  and ginst8814 (P2_ADD_391_1196_U110, P2_ADD_391_1196_U307, P2_ADD_391_1196_U308);
  and ginst8815 (P2_ADD_391_1196_U111, P2_ADD_391_1196_U309, P2_ADD_391_1196_U310);
  nand ginst8816 (P2_ADD_391_1196_U112, P2_ADD_391_1196_U186, P2_ADD_391_1196_U37);
  and ginst8817 (P2_ADD_391_1196_U113, P2_ADD_391_1196_U316, P2_ADD_391_1196_U317);
  and ginst8818 (P2_ADD_391_1196_U114, P2_ADD_391_1196_U323, P2_ADD_391_1196_U324);
  and ginst8819 (P2_ADD_391_1196_U115, P2_ADD_391_1196_U325, P2_ADD_391_1196_U326);
  nand ginst8820 (P2_ADD_391_1196_U116, P2_ADD_391_1196_U171, P2_ADD_391_1196_U172);
  and ginst8821 (P2_ADD_391_1196_U117, P2_ADD_391_1196_U332, P2_ADD_391_1196_U333);
  nand ginst8822 (P2_ADD_391_1196_U118, P2_ADD_391_1196_U167, P2_ADD_391_1196_U168);
  not ginst8823 (P2_ADD_391_1196_U119, P2_R2182_U41);
  nand ginst8824 (P2_ADD_391_1196_U12, P2_ADD_391_1196_U144, P2_ADD_391_1196_U306);
  not ginst8825 (P2_ADD_391_1196_U120, P2_R2096_U76);
  and ginst8826 (P2_ADD_391_1196_U121, P2_ADD_391_1196_U339, P2_ADD_391_1196_U340);
  and ginst8827 (P2_ADD_391_1196_U122, P2_ADD_391_1196_U344, P2_ADD_391_1196_U345);
  nand ginst8828 (P2_ADD_391_1196_U123, P2_ADD_391_1196_U143, P2_ADD_391_1196_U164);
  and ginst8829 (P2_ADD_391_1196_U124, P2_ADD_391_1196_U351, P2_ADD_391_1196_U352);
  and ginst8830 (P2_ADD_391_1196_U125, P2_ADD_391_1196_U358, P2_ADD_391_1196_U359);
  nand ginst8831 (P2_ADD_391_1196_U126, P2_ADD_391_1196_U273, P2_ADD_391_1196_U274);
  and ginst8832 (P2_ADD_391_1196_U127, P2_ADD_391_1196_U365, P2_ADD_391_1196_U366);
  nand ginst8833 (P2_ADD_391_1196_U128, P2_ADD_391_1196_U269, P2_ADD_391_1196_U270);
  and ginst8834 (P2_ADD_391_1196_U129, P2_ADD_391_1196_U372, P2_ADD_391_1196_U373);
  not ginst8835 (P2_ADD_391_1196_U13, P2_R2182_U72);
  nand ginst8836 (P2_ADD_391_1196_U130, P2_ADD_391_1196_U265, P2_ADD_391_1196_U266);
  and ginst8837 (P2_ADD_391_1196_U131, P2_ADD_391_1196_U379, P2_ADD_391_1196_U380);
  nand ginst8838 (P2_ADD_391_1196_U132, P2_ADD_391_1196_U261, P2_ADD_391_1196_U262);
  and ginst8839 (P2_ADD_391_1196_U133, P2_ADD_391_1196_U386, P2_ADD_391_1196_U387);
  nand ginst8840 (P2_ADD_391_1196_U134, P2_ADD_391_1196_U257, P2_ADD_391_1196_U258);
  and ginst8841 (P2_ADD_391_1196_U135, P2_ADD_391_1196_U393, P2_ADD_391_1196_U394);
  nand ginst8842 (P2_ADD_391_1196_U136, P2_ADD_391_1196_U253, P2_ADD_391_1196_U254);
  and ginst8843 (P2_ADD_391_1196_U137, P2_ADD_391_1196_U400, P2_ADD_391_1196_U401);
  nand ginst8844 (P2_ADD_391_1196_U138, P2_ADD_391_1196_U249, P2_ADD_391_1196_U250);
  and ginst8845 (P2_ADD_391_1196_U139, P2_ADD_391_1196_U407, P2_ADD_391_1196_U408);
  not ginst8846 (P2_ADD_391_1196_U14, P2_R2096_U71);
  nand ginst8847 (P2_ADD_391_1196_U140, P2_ADD_391_1196_U245, P2_ADD_391_1196_U246);
  and ginst8848 (P2_ADD_391_1196_U141, P2_ADD_391_1196_U414, P2_ADD_391_1196_U415);
  nand ginst8849 (P2_ADD_391_1196_U142, P2_ADD_391_1196_U241, P2_ADD_391_1196_U242);
  nand ginst8850 (P2_ADD_391_1196_U143, P2_ADD_391_1196_U162, P2_R2096_U51);
  and ginst8851 (P2_ADD_391_1196_U144, P2_ADD_391_1196_U424, P2_ADD_391_1196_U425);
  and ginst8852 (P2_ADD_391_1196_U145, P2_ADD_391_1196_U426, P2_ADD_391_1196_U427);
  nand ginst8853 (P2_ADD_391_1196_U146, P2_ADD_391_1196_U237, P2_ADD_391_1196_U238);
  and ginst8854 (P2_ADD_391_1196_U147, P2_ADD_391_1196_U433, P2_ADD_391_1196_U434);
  nand ginst8855 (P2_ADD_391_1196_U148, P2_ADD_391_1196_U233, P2_ADD_391_1196_U234);
  and ginst8856 (P2_ADD_391_1196_U149, P2_ADD_391_1196_U440, P2_ADD_391_1196_U441);
  not ginst8857 (P2_ADD_391_1196_U15, P2_R2182_U73);
  nand ginst8858 (P2_ADD_391_1196_U150, P2_ADD_391_1196_U229, P2_ADD_391_1196_U230);
  and ginst8859 (P2_ADD_391_1196_U151, P2_ADD_391_1196_U447, P2_ADD_391_1196_U448);
  nand ginst8860 (P2_ADD_391_1196_U152, P2_ADD_391_1196_U226, P2_ADD_391_1196_U83);
  and ginst8861 (P2_ADD_391_1196_U153, P2_ADD_391_1196_U454, P2_ADD_391_1196_U455);
  and ginst8862 (P2_ADD_391_1196_U154, P2_ADD_391_1196_U461, P2_ADD_391_1196_U462);
  and ginst8863 (P2_ADD_391_1196_U155, P2_ADD_391_1196_U463, P2_ADD_391_1196_U464);
  nand ginst8864 (P2_ADD_391_1196_U156, P2_ADD_391_1196_U212, P2_ADD_391_1196_U86);
  and ginst8865 (P2_ADD_391_1196_U157, P2_ADD_391_1196_U470, P2_ADD_391_1196_U471);
  nand ginst8866 (P2_ADD_391_1196_U158, P2_R2096_U97, P2_R2182_U96);
  nand ginst8867 (P2_ADD_391_1196_U159, P2_R2096_U93, P2_R2182_U92);
  not ginst8868 (P2_ADD_391_1196_U16, P2_R2096_U72);
  not ginst8869 (P2_ADD_391_1196_U160, P2_ADD_391_1196_U143);
  nand ginst8870 (P2_ADD_391_1196_U161, P2_R2096_U72, P2_R2182_U73);
  not ginst8871 (P2_ADD_391_1196_U162, P2_ADD_391_1196_U22);
  nand ginst8872 (P2_ADD_391_1196_U163, P2_ADD_391_1196_U22, P2_ADD_391_1196_U23);
  nand ginst8873 (P2_ADD_391_1196_U164, P2_ADD_391_1196_U163, P2_R2182_U68);
  not ginst8874 (P2_ADD_391_1196_U165, P2_ADD_391_1196_U123);
  or ginst8875 (P2_ADD_391_1196_U166, P2_R2096_U77, P2_R2182_U40);
  nand ginst8876 (P2_ADD_391_1196_U167, P2_ADD_391_1196_U123, P2_ADD_391_1196_U166);
  nand ginst8877 (P2_ADD_391_1196_U168, P2_R2096_U77, P2_R2182_U40);
  not ginst8878 (P2_ADD_391_1196_U169, P2_ADD_391_1196_U118);
  not ginst8879 (P2_ADD_391_1196_U17, P2_R2182_U74);
  or ginst8880 (P2_ADD_391_1196_U170, P2_R2096_U75, P2_R2182_U76);
  nand ginst8881 (P2_ADD_391_1196_U171, P2_ADD_391_1196_U118, P2_ADD_391_1196_U170);
  nand ginst8882 (P2_ADD_391_1196_U172, P2_R2096_U75, P2_R2182_U76);
  not ginst8883 (P2_ADD_391_1196_U173, P2_ADD_391_1196_U116);
  or ginst8884 (P2_ADD_391_1196_U174, P2_R2096_U74, P2_R2182_U75);
  nand ginst8885 (P2_ADD_391_1196_U175, P2_ADD_391_1196_U116, P2_ADD_391_1196_U174);
  nand ginst8886 (P2_ADD_391_1196_U176, P2_R2096_U74, P2_R2182_U75);
  not ginst8887 (P2_ADD_391_1196_U177, P2_ADD_391_1196_U38);
  or ginst8888 (P2_ADD_391_1196_U178, P2_R2096_U73, P2_R2182_U74);
  not ginst8889 (P2_ADD_391_1196_U179, P2_ADD_391_1196_U39);
  not ginst8890 (P2_ADD_391_1196_U18, P2_R2096_U73);
  nand ginst8891 (P2_ADD_391_1196_U180, P2_R2096_U73, P2_R2182_U74);
  not ginst8892 (P2_ADD_391_1196_U181, P2_ADD_391_1196_U30);
  nand ginst8893 (P2_ADD_391_1196_U182, P2_ADD_391_1196_U161, P2_ADD_391_1196_U181);
  or ginst8894 (P2_ADD_391_1196_U183, P2_R2096_U71, P2_R2182_U72);
  or ginst8895 (P2_ADD_391_1196_U184, P2_R2096_U72, P2_R2182_U73);
  not ginst8896 (P2_ADD_391_1196_U185, P2_ADD_391_1196_U37);
  nand ginst8897 (P2_ADD_391_1196_U186, P2_R2096_U71, P2_R2182_U72);
  not ginst8898 (P2_ADD_391_1196_U187, P2_ADD_391_1196_U112);
  or ginst8899 (P2_ADD_391_1196_U188, P2_R2096_U70, P2_R2182_U71);
  nand ginst8900 (P2_ADD_391_1196_U189, P2_ADD_391_1196_U112, P2_ADD_391_1196_U188);
  not ginst8901 (P2_ADD_391_1196_U19, P2_R2096_U68);
  nand ginst8902 (P2_ADD_391_1196_U190, P2_R2096_U70, P2_R2182_U71);
  not ginst8903 (P2_ADD_391_1196_U191, P2_ADD_391_1196_U35);
  nand ginst8904 (P2_ADD_391_1196_U192, P2_ADD_391_1196_U110, P2_ADD_391_1196_U191);
  or ginst8905 (P2_ADD_391_1196_U193, P2_R2096_U69, P2_R2182_U70);
  not ginst8906 (P2_ADD_391_1196_U194, P2_ADD_391_1196_U36);
  nand ginst8907 (P2_ADD_391_1196_U195, P2_R2096_U69, P2_R2182_U70);
  nand ginst8908 (P2_ADD_391_1196_U196, P2_ADD_391_1196_U194, P2_ADD_391_1196_U195);
  or ginst8909 (P2_ADD_391_1196_U197, P2_R2096_U72, P2_R2182_U73);
  nand ginst8910 (P2_ADD_391_1196_U198, P2_ADD_391_1196_U197, P2_ADD_391_1196_U30);
  nand ginst8911 (P2_ADD_391_1196_U199, P2_ADD_391_1196_U113, P2_ADD_391_1196_U161, P2_ADD_391_1196_U198);
  not ginst8912 (P2_ADD_391_1196_U20, P2_R2182_U69);
  nand ginst8913 (P2_ADD_391_1196_U200, P2_R2096_U71, P2_R2182_U72);
  nand ginst8914 (P2_ADD_391_1196_U201, P2_ADD_391_1196_U185, P2_ADD_391_1196_U200);
  or ginst8915 (P2_ADD_391_1196_U202, P2_R2096_U72, P2_R2182_U73);
  nand ginst8916 (P2_ADD_391_1196_U203, P2_ADD_391_1196_U114, P2_ADD_391_1196_U177);
  nand ginst8917 (P2_ADD_391_1196_U204, P2_R2096_U73, P2_R2182_U74);
  nand ginst8918 (P2_ADD_391_1196_U205, P2_ADD_391_1196_U179, P2_ADD_391_1196_U204);
  nand ginst8919 (P2_ADD_391_1196_U206, P2_R2096_U69, P2_R2182_U70);
  not ginst8920 (P2_ADD_391_1196_U207, P2_ADD_391_1196_U50);
  nand ginst8921 (P2_ADD_391_1196_U208, P2_ADD_391_1196_U158, P2_ADD_391_1196_U207);
  or ginst8922 (P2_ADD_391_1196_U209, P2_R2096_U96, P2_R2182_U95);
  not ginst8923 (P2_ADD_391_1196_U21, P2_R2182_U68);
  or ginst8924 (P2_ADD_391_1196_U210, P2_R2096_U97, P2_R2182_U96);
  not ginst8925 (P2_ADD_391_1196_U211, P2_ADD_391_1196_U86);
  nand ginst8926 (P2_ADD_391_1196_U212, P2_R2096_U96, P2_R2182_U95);
  not ginst8927 (P2_ADD_391_1196_U213, P2_ADD_391_1196_U156);
  or ginst8928 (P2_ADD_391_1196_U214, P2_R2096_U95, P2_R2182_U94);
  nand ginst8929 (P2_ADD_391_1196_U215, P2_ADD_391_1196_U156, P2_ADD_391_1196_U214);
  nand ginst8930 (P2_ADD_391_1196_U216, P2_R2096_U95, P2_R2182_U94);
  not ginst8931 (P2_ADD_391_1196_U217, P2_ADD_391_1196_U84);
  or ginst8932 (P2_ADD_391_1196_U218, P2_R2096_U94, P2_R2182_U93);
  not ginst8933 (P2_ADD_391_1196_U219, P2_ADD_391_1196_U85);
  nand ginst8934 (P2_ADD_391_1196_U22, P2_R2096_U68, P2_R2182_U69);
  nand ginst8935 (P2_ADD_391_1196_U220, P2_R2096_U94, P2_R2182_U93);
  not ginst8936 (P2_ADD_391_1196_U221, P2_ADD_391_1196_U53);
  nand ginst8937 (P2_ADD_391_1196_U222, P2_ADD_391_1196_U159, P2_ADD_391_1196_U221);
  or ginst8938 (P2_ADD_391_1196_U223, P2_R2096_U92, P2_R2182_U91);
  or ginst8939 (P2_ADD_391_1196_U224, P2_R2096_U93, P2_R2182_U92);
  not ginst8940 (P2_ADD_391_1196_U225, P2_ADD_391_1196_U83);
  nand ginst8941 (P2_ADD_391_1196_U226, P2_R2096_U92, P2_R2182_U91);
  not ginst8942 (P2_ADD_391_1196_U227, P2_ADD_391_1196_U152);
  or ginst8943 (P2_ADD_391_1196_U228, P2_R2096_U91, P2_R2182_U90);
  nand ginst8944 (P2_ADD_391_1196_U229, P2_ADD_391_1196_U152, P2_ADD_391_1196_U228);
  not ginst8945 (P2_ADD_391_1196_U23, P2_R2096_U51);
  nand ginst8946 (P2_ADD_391_1196_U230, P2_R2096_U91, P2_R2182_U90);
  not ginst8947 (P2_ADD_391_1196_U231, P2_ADD_391_1196_U150);
  or ginst8948 (P2_ADD_391_1196_U232, P2_R2096_U90, P2_R2182_U89);
  nand ginst8949 (P2_ADD_391_1196_U233, P2_ADD_391_1196_U150, P2_ADD_391_1196_U232);
  nand ginst8950 (P2_ADD_391_1196_U234, P2_R2096_U90, P2_R2182_U89);
  not ginst8951 (P2_ADD_391_1196_U235, P2_ADD_391_1196_U148);
  or ginst8952 (P2_ADD_391_1196_U236, P2_R2096_U89, P2_R2182_U88);
  nand ginst8953 (P2_ADD_391_1196_U237, P2_ADD_391_1196_U148, P2_ADD_391_1196_U236);
  nand ginst8954 (P2_ADD_391_1196_U238, P2_R2096_U89, P2_R2182_U88);
  not ginst8955 (P2_ADD_391_1196_U239, P2_ADD_391_1196_U146);
  not ginst8956 (P2_ADD_391_1196_U24, P2_R2182_U40);
  or ginst8957 (P2_ADD_391_1196_U240, P2_R2096_U88, P2_R2182_U87);
  nand ginst8958 (P2_ADD_391_1196_U241, P2_ADD_391_1196_U146, P2_ADD_391_1196_U240);
  nand ginst8959 (P2_ADD_391_1196_U242, P2_R2096_U88, P2_R2182_U87);
  not ginst8960 (P2_ADD_391_1196_U243, P2_ADD_391_1196_U142);
  or ginst8961 (P2_ADD_391_1196_U244, P2_R2096_U87, P2_R2182_U86);
  nand ginst8962 (P2_ADD_391_1196_U245, P2_ADD_391_1196_U142, P2_ADD_391_1196_U244);
  nand ginst8963 (P2_ADD_391_1196_U246, P2_R2096_U87, P2_R2182_U86);
  not ginst8964 (P2_ADD_391_1196_U247, P2_ADD_391_1196_U140);
  or ginst8965 (P2_ADD_391_1196_U248, P2_R2096_U86, P2_R2182_U85);
  nand ginst8966 (P2_ADD_391_1196_U249, P2_ADD_391_1196_U140, P2_ADD_391_1196_U248);
  not ginst8967 (P2_ADD_391_1196_U25, P2_R2096_U77);
  nand ginst8968 (P2_ADD_391_1196_U250, P2_R2096_U86, P2_R2182_U85);
  not ginst8969 (P2_ADD_391_1196_U251, P2_ADD_391_1196_U138);
  or ginst8970 (P2_ADD_391_1196_U252, P2_R2096_U85, P2_R2182_U84);
  nand ginst8971 (P2_ADD_391_1196_U253, P2_ADD_391_1196_U138, P2_ADD_391_1196_U252);
  nand ginst8972 (P2_ADD_391_1196_U254, P2_R2096_U85, P2_R2182_U84);
  not ginst8973 (P2_ADD_391_1196_U255, P2_ADD_391_1196_U136);
  or ginst8974 (P2_ADD_391_1196_U256, P2_R2096_U84, P2_R2182_U83);
  nand ginst8975 (P2_ADD_391_1196_U257, P2_ADD_391_1196_U136, P2_ADD_391_1196_U256);
  nand ginst8976 (P2_ADD_391_1196_U258, P2_R2096_U84, P2_R2182_U83);
  not ginst8977 (P2_ADD_391_1196_U259, P2_ADD_391_1196_U134);
  not ginst8978 (P2_ADD_391_1196_U26, P2_R2182_U76);
  or ginst8979 (P2_ADD_391_1196_U260, P2_R2096_U83, P2_R2182_U82);
  nand ginst8980 (P2_ADD_391_1196_U261, P2_ADD_391_1196_U134, P2_ADD_391_1196_U260);
  nand ginst8981 (P2_ADD_391_1196_U262, P2_R2096_U83, P2_R2182_U82);
  not ginst8982 (P2_ADD_391_1196_U263, P2_ADD_391_1196_U132);
  or ginst8983 (P2_ADD_391_1196_U264, P2_R2096_U82, P2_R2182_U81);
  nand ginst8984 (P2_ADD_391_1196_U265, P2_ADD_391_1196_U132, P2_ADD_391_1196_U264);
  nand ginst8985 (P2_ADD_391_1196_U266, P2_R2096_U82, P2_R2182_U81);
  not ginst8986 (P2_ADD_391_1196_U267, P2_ADD_391_1196_U130);
  or ginst8987 (P2_ADD_391_1196_U268, P2_R2096_U81, P2_R2182_U80);
  nand ginst8988 (P2_ADD_391_1196_U269, P2_ADD_391_1196_U130, P2_ADD_391_1196_U268);
  not ginst8989 (P2_ADD_391_1196_U27, P2_R2096_U75);
  nand ginst8990 (P2_ADD_391_1196_U270, P2_R2096_U81, P2_R2182_U80);
  not ginst8991 (P2_ADD_391_1196_U271, P2_ADD_391_1196_U128);
  or ginst8992 (P2_ADD_391_1196_U272, P2_R2096_U80, P2_R2182_U79);
  nand ginst8993 (P2_ADD_391_1196_U273, P2_ADD_391_1196_U128, P2_ADD_391_1196_U272);
  nand ginst8994 (P2_ADD_391_1196_U274, P2_R2096_U80, P2_R2182_U79);
  not ginst8995 (P2_ADD_391_1196_U275, P2_ADD_391_1196_U126);
  or ginst8996 (P2_ADD_391_1196_U276, P2_R2096_U79, P2_R2182_U78);
  nand ginst8997 (P2_ADD_391_1196_U277, P2_ADD_391_1196_U126, P2_ADD_391_1196_U276);
  nand ginst8998 (P2_ADD_391_1196_U278, P2_R2096_U79, P2_R2182_U78);
  not ginst8999 (P2_ADD_391_1196_U279, P2_ADD_391_1196_U82);
  not ginst9000 (P2_ADD_391_1196_U28, P2_R2182_U75);
  or ginst9001 (P2_ADD_391_1196_U280, P2_R2096_U78, P2_R2182_U77);
  nand ginst9002 (P2_ADD_391_1196_U281, P2_ADD_391_1196_U280, P2_ADD_391_1196_U82);
  nand ginst9003 (P2_ADD_391_1196_U282, P2_R2096_U78, P2_R2182_U77);
  nand ginst9004 (P2_ADD_391_1196_U283, P2_ADD_391_1196_U121, P2_ADD_391_1196_U281, P2_ADD_391_1196_U282);
  nand ginst9005 (P2_ADD_391_1196_U284, P2_R2096_U78, P2_R2182_U77);
  nand ginst9006 (P2_ADD_391_1196_U285, P2_ADD_391_1196_U279, P2_ADD_391_1196_U284);
  or ginst9007 (P2_ADD_391_1196_U286, P2_R2096_U78, P2_R2182_U77);
  nand ginst9008 (P2_ADD_391_1196_U287, P2_ADD_391_1196_U285, P2_ADD_391_1196_U286, P2_ADD_391_1196_U343);
  or ginst9009 (P2_ADD_391_1196_U288, P2_R2096_U93, P2_R2182_U92);
  nand ginst9010 (P2_ADD_391_1196_U289, P2_ADD_391_1196_U288, P2_ADD_391_1196_U53);
  not ginst9011 (P2_ADD_391_1196_U29, P2_R2096_U74);
  nand ginst9012 (P2_ADD_391_1196_U290, P2_ADD_391_1196_U153, P2_ADD_391_1196_U159, P2_ADD_391_1196_U289);
  nand ginst9013 (P2_ADD_391_1196_U291, P2_R2096_U92, P2_R2182_U91);
  nand ginst9014 (P2_ADD_391_1196_U292, P2_ADD_391_1196_U225, P2_ADD_391_1196_U291);
  or ginst9015 (P2_ADD_391_1196_U293, P2_R2096_U93, P2_R2182_U92);
  nand ginst9016 (P2_ADD_391_1196_U294, P2_ADD_391_1196_U154, P2_ADD_391_1196_U217);
  nand ginst9017 (P2_ADD_391_1196_U295, P2_R2096_U94, P2_R2182_U93);
  nand ginst9018 (P2_ADD_391_1196_U296, P2_ADD_391_1196_U219, P2_ADD_391_1196_U295);
  or ginst9019 (P2_ADD_391_1196_U297, P2_R2096_U97, P2_R2182_U96);
  nand ginst9020 (P2_ADD_391_1196_U298, P2_ADD_391_1196_U297, P2_ADD_391_1196_U50);
  nand ginst9021 (P2_ADD_391_1196_U299, P2_ADD_391_1196_U157, P2_ADD_391_1196_U158, P2_ADD_391_1196_U298);
  nand ginst9022 (P2_ADD_391_1196_U30, P2_ADD_391_1196_U180, P2_ADD_391_1196_U39);
  nand ginst9023 (P2_ADD_391_1196_U300, P2_R2096_U96, P2_R2182_U95);
  nand ginst9024 (P2_ADD_391_1196_U301, P2_ADD_391_1196_U211, P2_ADD_391_1196_U300);
  or ginst9025 (P2_ADD_391_1196_U302, P2_R2096_U97, P2_R2182_U96);
  nand ginst9026 (P2_ADD_391_1196_U303, P2_ADD_391_1196_U161, P2_ADD_391_1196_U202);
  nand ginst9027 (P2_ADD_391_1196_U304, P2_ADD_391_1196_U159, P2_ADD_391_1196_U293);
  nand ginst9028 (P2_ADD_391_1196_U305, P2_ADD_391_1196_U158, P2_ADD_391_1196_U302);
  nand ginst9029 (P2_ADD_391_1196_U306, P2_ADD_391_1196_U23, P2_ADD_391_1196_U423);
  nand ginst9030 (P2_ADD_391_1196_U307, P2_ADD_391_1196_U34, P2_R2096_U69);
  nand ginst9031 (P2_ADD_391_1196_U308, P2_ADD_391_1196_U33, P2_R2182_U70);
  nand ginst9032 (P2_ADD_391_1196_U309, P2_ADD_391_1196_U31, P2_R2096_U70);
  not ginst9033 (P2_ADD_391_1196_U31, P2_R2182_U71);
  nand ginst9034 (P2_ADD_391_1196_U310, P2_ADD_391_1196_U32, P2_R2182_U71);
  nand ginst9035 (P2_ADD_391_1196_U311, P2_ADD_391_1196_U31, P2_R2096_U70);
  nand ginst9036 (P2_ADD_391_1196_U312, P2_ADD_391_1196_U32, P2_R2182_U71);
  nand ginst9037 (P2_ADD_391_1196_U313, P2_ADD_391_1196_U311, P2_ADD_391_1196_U312);
  nand ginst9038 (P2_ADD_391_1196_U314, P2_ADD_391_1196_U111, P2_ADD_391_1196_U112);
  nand ginst9039 (P2_ADD_391_1196_U315, P2_ADD_391_1196_U187, P2_ADD_391_1196_U313);
  nand ginst9040 (P2_ADD_391_1196_U316, P2_ADD_391_1196_U13, P2_R2096_U71);
  nand ginst9041 (P2_ADD_391_1196_U317, P2_ADD_391_1196_U14, P2_R2182_U72);
  nand ginst9042 (P2_ADD_391_1196_U318, P2_ADD_391_1196_U15, P2_R2096_U72);
  nand ginst9043 (P2_ADD_391_1196_U319, P2_ADD_391_1196_U16, P2_R2182_U73);
  not ginst9044 (P2_ADD_391_1196_U32, P2_R2096_U70);
  nand ginst9045 (P2_ADD_391_1196_U320, P2_ADD_391_1196_U318, P2_ADD_391_1196_U319);
  nand ginst9046 (P2_ADD_391_1196_U321, P2_ADD_391_1196_U30, P2_ADD_391_1196_U303);
  nand ginst9047 (P2_ADD_391_1196_U322, P2_ADD_391_1196_U181, P2_ADD_391_1196_U320);
  nand ginst9048 (P2_ADD_391_1196_U323, P2_ADD_391_1196_U17, P2_R2096_U73);
  nand ginst9049 (P2_ADD_391_1196_U324, P2_ADD_391_1196_U18, P2_R2182_U74);
  nand ginst9050 (P2_ADD_391_1196_U325, P2_ADD_391_1196_U28, P2_R2096_U74);
  nand ginst9051 (P2_ADD_391_1196_U326, P2_ADD_391_1196_U29, P2_R2182_U75);
  nand ginst9052 (P2_ADD_391_1196_U327, P2_ADD_391_1196_U28, P2_R2096_U74);
  nand ginst9053 (P2_ADD_391_1196_U328, P2_ADD_391_1196_U29, P2_R2182_U75);
  nand ginst9054 (P2_ADD_391_1196_U329, P2_ADD_391_1196_U327, P2_ADD_391_1196_U328);
  not ginst9055 (P2_ADD_391_1196_U33, P2_R2096_U69);
  nand ginst9056 (P2_ADD_391_1196_U330, P2_ADD_391_1196_U115, P2_ADD_391_1196_U116);
  nand ginst9057 (P2_ADD_391_1196_U331, P2_ADD_391_1196_U173, P2_ADD_391_1196_U329);
  nand ginst9058 (P2_ADD_391_1196_U332, P2_ADD_391_1196_U26, P2_R2096_U75);
  nand ginst9059 (P2_ADD_391_1196_U333, P2_ADD_391_1196_U27, P2_R2182_U76);
  nand ginst9060 (P2_ADD_391_1196_U334, P2_ADD_391_1196_U26, P2_R2096_U75);
  nand ginst9061 (P2_ADD_391_1196_U335, P2_ADD_391_1196_U27, P2_R2182_U76);
  nand ginst9062 (P2_ADD_391_1196_U336, P2_ADD_391_1196_U334, P2_ADD_391_1196_U335);
  nand ginst9063 (P2_ADD_391_1196_U337, P2_ADD_391_1196_U117, P2_ADD_391_1196_U118);
  nand ginst9064 (P2_ADD_391_1196_U338, P2_ADD_391_1196_U169, P2_ADD_391_1196_U336);
  nand ginst9065 (P2_ADD_391_1196_U339, P2_ADD_391_1196_U120, P2_R2182_U41);
  not ginst9066 (P2_ADD_391_1196_U34, P2_R2182_U70);
  nand ginst9067 (P2_ADD_391_1196_U340, P2_ADD_391_1196_U119, P2_R2096_U76);
  nand ginst9068 (P2_ADD_391_1196_U341, P2_ADD_391_1196_U120, P2_R2182_U41);
  nand ginst9069 (P2_ADD_391_1196_U342, P2_ADD_391_1196_U119, P2_R2096_U76);
  nand ginst9070 (P2_ADD_391_1196_U343, P2_ADD_391_1196_U341, P2_ADD_391_1196_U342);
  nand ginst9071 (P2_ADD_391_1196_U344, P2_ADD_391_1196_U24, P2_R2096_U77);
  nand ginst9072 (P2_ADD_391_1196_U345, P2_ADD_391_1196_U25, P2_R2182_U40);
  nand ginst9073 (P2_ADD_391_1196_U346, P2_ADD_391_1196_U24, P2_R2096_U77);
  nand ginst9074 (P2_ADD_391_1196_U347, P2_ADD_391_1196_U25, P2_R2182_U40);
  nand ginst9075 (P2_ADD_391_1196_U348, P2_ADD_391_1196_U346, P2_ADD_391_1196_U347);
  nand ginst9076 (P2_ADD_391_1196_U349, P2_ADD_391_1196_U122, P2_ADD_391_1196_U123);
  nand ginst9077 (P2_ADD_391_1196_U35, P2_ADD_391_1196_U189, P2_ADD_391_1196_U190);
  nand ginst9078 (P2_ADD_391_1196_U350, P2_ADD_391_1196_U165, P2_ADD_391_1196_U348);
  nand ginst9079 (P2_ADD_391_1196_U351, P2_ADD_391_1196_U80, P2_R2182_U77);
  nand ginst9080 (P2_ADD_391_1196_U352, P2_ADD_391_1196_U81, P2_R2096_U78);
  nand ginst9081 (P2_ADD_391_1196_U353, P2_ADD_391_1196_U80, P2_R2182_U77);
  nand ginst9082 (P2_ADD_391_1196_U354, P2_ADD_391_1196_U81, P2_R2096_U78);
  nand ginst9083 (P2_ADD_391_1196_U355, P2_ADD_391_1196_U353, P2_ADD_391_1196_U354);
  nand ginst9084 (P2_ADD_391_1196_U356, P2_ADD_391_1196_U124, P2_ADD_391_1196_U82);
  nand ginst9085 (P2_ADD_391_1196_U357, P2_ADD_391_1196_U279, P2_ADD_391_1196_U355);
  nand ginst9086 (P2_ADD_391_1196_U358, P2_ADD_391_1196_U78, P2_R2182_U78);
  nand ginst9087 (P2_ADD_391_1196_U359, P2_ADD_391_1196_U79, P2_R2096_U79);
  nand ginst9088 (P2_ADD_391_1196_U36, P2_ADD_391_1196_U193, P2_ADD_391_1196_U35);
  nand ginst9089 (P2_ADD_391_1196_U360, P2_ADD_391_1196_U78, P2_R2182_U78);
  nand ginst9090 (P2_ADD_391_1196_U361, P2_ADD_391_1196_U79, P2_R2096_U79);
  nand ginst9091 (P2_ADD_391_1196_U362, P2_ADD_391_1196_U360, P2_ADD_391_1196_U361);
  nand ginst9092 (P2_ADD_391_1196_U363, P2_ADD_391_1196_U125, P2_ADD_391_1196_U126);
  nand ginst9093 (P2_ADD_391_1196_U364, P2_ADD_391_1196_U275, P2_ADD_391_1196_U362);
  nand ginst9094 (P2_ADD_391_1196_U365, P2_ADD_391_1196_U76, P2_R2096_U80);
  nand ginst9095 (P2_ADD_391_1196_U366, P2_ADD_391_1196_U77, P2_R2182_U79);
  nand ginst9096 (P2_ADD_391_1196_U367, P2_ADD_391_1196_U76, P2_R2096_U80);
  nand ginst9097 (P2_ADD_391_1196_U368, P2_ADD_391_1196_U77, P2_R2182_U79);
  nand ginst9098 (P2_ADD_391_1196_U369, P2_ADD_391_1196_U367, P2_ADD_391_1196_U368);
  nand ginst9099 (P2_ADD_391_1196_U37, P2_ADD_391_1196_U182, P2_ADD_391_1196_U183, P2_ADD_391_1196_U184);
  nand ginst9100 (P2_ADD_391_1196_U370, P2_ADD_391_1196_U127, P2_ADD_391_1196_U128);
  nand ginst9101 (P2_ADD_391_1196_U371, P2_ADD_391_1196_U271, P2_ADD_391_1196_U369);
  nand ginst9102 (P2_ADD_391_1196_U372, P2_ADD_391_1196_U74, P2_R2096_U81);
  nand ginst9103 (P2_ADD_391_1196_U373, P2_ADD_391_1196_U75, P2_R2182_U80);
  nand ginst9104 (P2_ADD_391_1196_U374, P2_ADD_391_1196_U74, P2_R2096_U81);
  nand ginst9105 (P2_ADD_391_1196_U375, P2_ADD_391_1196_U75, P2_R2182_U80);
  nand ginst9106 (P2_ADD_391_1196_U376, P2_ADD_391_1196_U374, P2_ADD_391_1196_U375);
  nand ginst9107 (P2_ADD_391_1196_U377, P2_ADD_391_1196_U129, P2_ADD_391_1196_U130);
  nand ginst9108 (P2_ADD_391_1196_U378, P2_ADD_391_1196_U267, P2_ADD_391_1196_U376);
  nand ginst9109 (P2_ADD_391_1196_U379, P2_ADD_391_1196_U72, P2_R2096_U82);
  nand ginst9110 (P2_ADD_391_1196_U38, P2_ADD_391_1196_U175, P2_ADD_391_1196_U176);
  nand ginst9111 (P2_ADD_391_1196_U380, P2_ADD_391_1196_U73, P2_R2182_U81);
  nand ginst9112 (P2_ADD_391_1196_U381, P2_ADD_391_1196_U72, P2_R2096_U82);
  nand ginst9113 (P2_ADD_391_1196_U382, P2_ADD_391_1196_U73, P2_R2182_U81);
  nand ginst9114 (P2_ADD_391_1196_U383, P2_ADD_391_1196_U381, P2_ADD_391_1196_U382);
  nand ginst9115 (P2_ADD_391_1196_U384, P2_ADD_391_1196_U131, P2_ADD_391_1196_U132);
  nand ginst9116 (P2_ADD_391_1196_U385, P2_ADD_391_1196_U263, P2_ADD_391_1196_U383);
  nand ginst9117 (P2_ADD_391_1196_U386, P2_ADD_391_1196_U70, P2_R2096_U83);
  nand ginst9118 (P2_ADD_391_1196_U387, P2_ADD_391_1196_U71, P2_R2182_U82);
  nand ginst9119 (P2_ADD_391_1196_U388, P2_ADD_391_1196_U70, P2_R2096_U83);
  nand ginst9120 (P2_ADD_391_1196_U389, P2_ADD_391_1196_U71, P2_R2182_U82);
  nand ginst9121 (P2_ADD_391_1196_U39, P2_ADD_391_1196_U178, P2_ADD_391_1196_U38);
  nand ginst9122 (P2_ADD_391_1196_U390, P2_ADD_391_1196_U388, P2_ADD_391_1196_U389);
  nand ginst9123 (P2_ADD_391_1196_U391, P2_ADD_391_1196_U133, P2_ADD_391_1196_U134);
  nand ginst9124 (P2_ADD_391_1196_U392, P2_ADD_391_1196_U259, P2_ADD_391_1196_U390);
  nand ginst9125 (P2_ADD_391_1196_U393, P2_ADD_391_1196_U68, P2_R2096_U84);
  nand ginst9126 (P2_ADD_391_1196_U394, P2_ADD_391_1196_U69, P2_R2182_U83);
  nand ginst9127 (P2_ADD_391_1196_U395, P2_ADD_391_1196_U68, P2_R2096_U84);
  nand ginst9128 (P2_ADD_391_1196_U396, P2_ADD_391_1196_U69, P2_R2182_U83);
  nand ginst9129 (P2_ADD_391_1196_U397, P2_ADD_391_1196_U395, P2_ADD_391_1196_U396);
  nand ginst9130 (P2_ADD_391_1196_U398, P2_ADD_391_1196_U135, P2_ADD_391_1196_U136);
  nand ginst9131 (P2_ADD_391_1196_U399, P2_ADD_391_1196_U255, P2_ADD_391_1196_U397);
  not ginst9132 (P2_ADD_391_1196_U40, P2_R2182_U91);
  nand ginst9133 (P2_ADD_391_1196_U400, P2_ADD_391_1196_U66, P2_R2096_U85);
  nand ginst9134 (P2_ADD_391_1196_U401, P2_ADD_391_1196_U67, P2_R2182_U84);
  nand ginst9135 (P2_ADD_391_1196_U402, P2_ADD_391_1196_U66, P2_R2096_U85);
  nand ginst9136 (P2_ADD_391_1196_U403, P2_ADD_391_1196_U67, P2_R2182_U84);
  nand ginst9137 (P2_ADD_391_1196_U404, P2_ADD_391_1196_U402, P2_ADD_391_1196_U403);
  nand ginst9138 (P2_ADD_391_1196_U405, P2_ADD_391_1196_U137, P2_ADD_391_1196_U138);
  nand ginst9139 (P2_ADD_391_1196_U406, P2_ADD_391_1196_U251, P2_ADD_391_1196_U404);
  nand ginst9140 (P2_ADD_391_1196_U407, P2_ADD_391_1196_U64, P2_R2096_U86);
  nand ginst9141 (P2_ADD_391_1196_U408, P2_ADD_391_1196_U65, P2_R2182_U85);
  nand ginst9142 (P2_ADD_391_1196_U409, P2_ADD_391_1196_U64, P2_R2096_U86);
  not ginst9143 (P2_ADD_391_1196_U41, P2_R2096_U92);
  nand ginst9144 (P2_ADD_391_1196_U410, P2_ADD_391_1196_U65, P2_R2182_U85);
  nand ginst9145 (P2_ADD_391_1196_U411, P2_ADD_391_1196_U409, P2_ADD_391_1196_U410);
  nand ginst9146 (P2_ADD_391_1196_U412, P2_ADD_391_1196_U139, P2_ADD_391_1196_U140);
  nand ginst9147 (P2_ADD_391_1196_U413, P2_ADD_391_1196_U247, P2_ADD_391_1196_U411);
  nand ginst9148 (P2_ADD_391_1196_U414, P2_ADD_391_1196_U62, P2_R2096_U87);
  nand ginst9149 (P2_ADD_391_1196_U415, P2_ADD_391_1196_U63, P2_R2182_U86);
  nand ginst9150 (P2_ADD_391_1196_U416, P2_ADD_391_1196_U62, P2_R2096_U87);
  nand ginst9151 (P2_ADD_391_1196_U417, P2_ADD_391_1196_U63, P2_R2182_U86);
  nand ginst9152 (P2_ADD_391_1196_U418, P2_ADD_391_1196_U416, P2_ADD_391_1196_U417);
  nand ginst9153 (P2_ADD_391_1196_U419, P2_ADD_391_1196_U141, P2_ADD_391_1196_U142);
  not ginst9154 (P2_ADD_391_1196_U42, P2_R2182_U92);
  nand ginst9155 (P2_ADD_391_1196_U420, P2_ADD_391_1196_U243, P2_ADD_391_1196_U418);
  nand ginst9156 (P2_ADD_391_1196_U421, P2_ADD_391_1196_U22, P2_R2182_U68);
  nand ginst9157 (P2_ADD_391_1196_U422, P2_ADD_391_1196_U162, P2_ADD_391_1196_U21);
  nand ginst9158 (P2_ADD_391_1196_U423, P2_ADD_391_1196_U421, P2_ADD_391_1196_U422);
  nand ginst9159 (P2_ADD_391_1196_U424, P2_ADD_391_1196_U21, P2_ADD_391_1196_U22, P2_R2096_U51);
  nand ginst9160 (P2_ADD_391_1196_U425, P2_ADD_391_1196_U160, P2_R2182_U68);
  nand ginst9161 (P2_ADD_391_1196_U426, P2_ADD_391_1196_U60, P2_R2096_U88);
  nand ginst9162 (P2_ADD_391_1196_U427, P2_ADD_391_1196_U61, P2_R2182_U87);
  nand ginst9163 (P2_ADD_391_1196_U428, P2_ADD_391_1196_U60, P2_R2096_U88);
  nand ginst9164 (P2_ADD_391_1196_U429, P2_ADD_391_1196_U61, P2_R2182_U87);
  not ginst9165 (P2_ADD_391_1196_U43, P2_R2096_U93);
  nand ginst9166 (P2_ADD_391_1196_U430, P2_ADD_391_1196_U428, P2_ADD_391_1196_U429);
  nand ginst9167 (P2_ADD_391_1196_U431, P2_ADD_391_1196_U145, P2_ADD_391_1196_U146);
  nand ginst9168 (P2_ADD_391_1196_U432, P2_ADD_391_1196_U239, P2_ADD_391_1196_U430);
  nand ginst9169 (P2_ADD_391_1196_U433, P2_ADD_391_1196_U58, P2_R2096_U89);
  nand ginst9170 (P2_ADD_391_1196_U434, P2_ADD_391_1196_U59, P2_R2182_U88);
  nand ginst9171 (P2_ADD_391_1196_U435, P2_ADD_391_1196_U58, P2_R2096_U89);
  nand ginst9172 (P2_ADD_391_1196_U436, P2_ADD_391_1196_U59, P2_R2182_U88);
  nand ginst9173 (P2_ADD_391_1196_U437, P2_ADD_391_1196_U435, P2_ADD_391_1196_U436);
  nand ginst9174 (P2_ADD_391_1196_U438, P2_ADD_391_1196_U147, P2_ADD_391_1196_U148);
  nand ginst9175 (P2_ADD_391_1196_U439, P2_ADD_391_1196_U235, P2_ADD_391_1196_U437);
  not ginst9176 (P2_ADD_391_1196_U44, P2_R2182_U93);
  nand ginst9177 (P2_ADD_391_1196_U440, P2_ADD_391_1196_U56, P2_R2096_U90);
  nand ginst9178 (P2_ADD_391_1196_U441, P2_ADD_391_1196_U57, P2_R2182_U89);
  nand ginst9179 (P2_ADD_391_1196_U442, P2_ADD_391_1196_U56, P2_R2096_U90);
  nand ginst9180 (P2_ADD_391_1196_U443, P2_ADD_391_1196_U57, P2_R2182_U89);
  nand ginst9181 (P2_ADD_391_1196_U444, P2_ADD_391_1196_U442, P2_ADD_391_1196_U443);
  nand ginst9182 (P2_ADD_391_1196_U445, P2_ADD_391_1196_U149, P2_ADD_391_1196_U150);
  nand ginst9183 (P2_ADD_391_1196_U446, P2_ADD_391_1196_U231, P2_ADD_391_1196_U444);
  nand ginst9184 (P2_ADD_391_1196_U447, P2_ADD_391_1196_U54, P2_R2096_U91);
  nand ginst9185 (P2_ADD_391_1196_U448, P2_ADD_391_1196_U55, P2_R2182_U90);
  nand ginst9186 (P2_ADD_391_1196_U449, P2_ADD_391_1196_U54, P2_R2096_U91);
  not ginst9187 (P2_ADD_391_1196_U45, P2_R2096_U94);
  nand ginst9188 (P2_ADD_391_1196_U450, P2_ADD_391_1196_U55, P2_R2182_U90);
  nand ginst9189 (P2_ADD_391_1196_U451, P2_ADD_391_1196_U449, P2_ADD_391_1196_U450);
  nand ginst9190 (P2_ADD_391_1196_U452, P2_ADD_391_1196_U151, P2_ADD_391_1196_U152);
  nand ginst9191 (P2_ADD_391_1196_U453, P2_ADD_391_1196_U227, P2_ADD_391_1196_U451);
  nand ginst9192 (P2_ADD_391_1196_U454, P2_ADD_391_1196_U40, P2_R2096_U92);
  nand ginst9193 (P2_ADD_391_1196_U455, P2_ADD_391_1196_U41, P2_R2182_U91);
  nand ginst9194 (P2_ADD_391_1196_U456, P2_ADD_391_1196_U42, P2_R2096_U93);
  nand ginst9195 (P2_ADD_391_1196_U457, P2_ADD_391_1196_U43, P2_R2182_U92);
  nand ginst9196 (P2_ADD_391_1196_U458, P2_ADD_391_1196_U456, P2_ADD_391_1196_U457);
  nand ginst9197 (P2_ADD_391_1196_U459, P2_ADD_391_1196_U304, P2_ADD_391_1196_U53);
  not ginst9198 (P2_ADD_391_1196_U46, P2_R2182_U95);
  nand ginst9199 (P2_ADD_391_1196_U460, P2_ADD_391_1196_U221, P2_ADD_391_1196_U458);
  nand ginst9200 (P2_ADD_391_1196_U461, P2_ADD_391_1196_U44, P2_R2096_U94);
  nand ginst9201 (P2_ADD_391_1196_U462, P2_ADD_391_1196_U45, P2_R2182_U93);
  nand ginst9202 (P2_ADD_391_1196_U463, P2_ADD_391_1196_U51, P2_R2096_U95);
  nand ginst9203 (P2_ADD_391_1196_U464, P2_ADD_391_1196_U52, P2_R2182_U94);
  nand ginst9204 (P2_ADD_391_1196_U465, P2_ADD_391_1196_U51, P2_R2096_U95);
  nand ginst9205 (P2_ADD_391_1196_U466, P2_ADD_391_1196_U52, P2_R2182_U94);
  nand ginst9206 (P2_ADD_391_1196_U467, P2_ADD_391_1196_U465, P2_ADD_391_1196_U466);
  nand ginst9207 (P2_ADD_391_1196_U468, P2_ADD_391_1196_U155, P2_ADD_391_1196_U156);
  nand ginst9208 (P2_ADD_391_1196_U469, P2_ADD_391_1196_U213, P2_ADD_391_1196_U467);
  not ginst9209 (P2_ADD_391_1196_U47, P2_R2096_U96);
  nand ginst9210 (P2_ADD_391_1196_U470, P2_ADD_391_1196_U46, P2_R2096_U96);
  nand ginst9211 (P2_ADD_391_1196_U471, P2_ADD_391_1196_U47, P2_R2182_U95);
  nand ginst9212 (P2_ADD_391_1196_U472, P2_ADD_391_1196_U48, P2_R2096_U97);
  nand ginst9213 (P2_ADD_391_1196_U473, P2_ADD_391_1196_U49, P2_R2182_U96);
  nand ginst9214 (P2_ADD_391_1196_U474, P2_ADD_391_1196_U472, P2_ADD_391_1196_U473);
  nand ginst9215 (P2_ADD_391_1196_U475, P2_ADD_391_1196_U305, P2_ADD_391_1196_U50);
  nand ginst9216 (P2_ADD_391_1196_U476, P2_ADD_391_1196_U207, P2_ADD_391_1196_U474);
  nand ginst9217 (P2_ADD_391_1196_U477, P2_ADD_391_1196_U19, P2_R2182_U69);
  nand ginst9218 (P2_ADD_391_1196_U478, P2_ADD_391_1196_U20, P2_R2096_U68);
  not ginst9219 (P2_ADD_391_1196_U48, P2_R2182_U96);
  not ginst9220 (P2_ADD_391_1196_U49, P2_R2096_U97);
  and ginst9221 (P2_ADD_391_1196_U5, P2_ADD_391_1196_U299, P2_ADD_391_1196_U301);
  nand ginst9222 (P2_ADD_391_1196_U50, P2_ADD_391_1196_U206, P2_ADD_391_1196_U36);
  not ginst9223 (P2_ADD_391_1196_U51, P2_R2182_U94);
  not ginst9224 (P2_ADD_391_1196_U52, P2_R2096_U95);
  nand ginst9225 (P2_ADD_391_1196_U53, P2_ADD_391_1196_U220, P2_ADD_391_1196_U85);
  not ginst9226 (P2_ADD_391_1196_U54, P2_R2182_U90);
  not ginst9227 (P2_ADD_391_1196_U55, P2_R2096_U91);
  not ginst9228 (P2_ADD_391_1196_U56, P2_R2182_U89);
  not ginst9229 (P2_ADD_391_1196_U57, P2_R2096_U90);
  not ginst9230 (P2_ADD_391_1196_U58, P2_R2182_U88);
  not ginst9231 (P2_ADD_391_1196_U59, P2_R2096_U89);
  and ginst9232 (P2_ADD_391_1196_U6, P2_ADD_391_1196_U294, P2_ADD_391_1196_U296);
  not ginst9233 (P2_ADD_391_1196_U60, P2_R2182_U87);
  not ginst9234 (P2_ADD_391_1196_U61, P2_R2096_U88);
  not ginst9235 (P2_ADD_391_1196_U62, P2_R2182_U86);
  not ginst9236 (P2_ADD_391_1196_U63, P2_R2096_U87);
  not ginst9237 (P2_ADD_391_1196_U64, P2_R2182_U85);
  not ginst9238 (P2_ADD_391_1196_U65, P2_R2096_U86);
  not ginst9239 (P2_ADD_391_1196_U66, P2_R2182_U84);
  not ginst9240 (P2_ADD_391_1196_U67, P2_R2096_U85);
  not ginst9241 (P2_ADD_391_1196_U68, P2_R2182_U83);
  not ginst9242 (P2_ADD_391_1196_U69, P2_R2096_U84);
  and ginst9243 (P2_ADD_391_1196_U7, P2_ADD_391_1196_U290, P2_ADD_391_1196_U292);
  not ginst9244 (P2_ADD_391_1196_U70, P2_R2182_U82);
  not ginst9245 (P2_ADD_391_1196_U71, P2_R2096_U83);
  not ginst9246 (P2_ADD_391_1196_U72, P2_R2182_U81);
  not ginst9247 (P2_ADD_391_1196_U73, P2_R2096_U82);
  not ginst9248 (P2_ADD_391_1196_U74, P2_R2182_U80);
  not ginst9249 (P2_ADD_391_1196_U75, P2_R2096_U81);
  not ginst9250 (P2_ADD_391_1196_U76, P2_R2182_U79);
  not ginst9251 (P2_ADD_391_1196_U77, P2_R2096_U80);
  not ginst9252 (P2_ADD_391_1196_U78, P2_R2096_U79);
  not ginst9253 (P2_ADD_391_1196_U79, P2_R2182_U78);
  and ginst9254 (P2_ADD_391_1196_U8, P2_ADD_391_1196_U283, P2_ADD_391_1196_U287);
  not ginst9255 (P2_ADD_391_1196_U80, P2_R2096_U78);
  not ginst9256 (P2_ADD_391_1196_U81, P2_R2182_U77);
  nand ginst9257 (P2_ADD_391_1196_U82, P2_ADD_391_1196_U277, P2_ADD_391_1196_U278);
  nand ginst9258 (P2_ADD_391_1196_U83, P2_ADD_391_1196_U222, P2_ADD_391_1196_U223, P2_ADD_391_1196_U224);
  nand ginst9259 (P2_ADD_391_1196_U84, P2_ADD_391_1196_U215, P2_ADD_391_1196_U216);
  nand ginst9260 (P2_ADD_391_1196_U85, P2_ADD_391_1196_U218, P2_ADD_391_1196_U84);
  nand ginst9261 (P2_ADD_391_1196_U86, P2_ADD_391_1196_U208, P2_ADD_391_1196_U209, P2_ADD_391_1196_U210);
  nand ginst9262 (P2_ADD_391_1196_U87, P2_ADD_391_1196_U477, P2_ADD_391_1196_U478);
  nand ginst9263 (P2_ADD_391_1196_U88, P2_ADD_391_1196_U314, P2_ADD_391_1196_U315);
  nand ginst9264 (P2_ADD_391_1196_U89, P2_ADD_391_1196_U321, P2_ADD_391_1196_U322);
  and ginst9265 (P2_ADD_391_1196_U9, P2_ADD_391_1196_U203, P2_ADD_391_1196_U205);
  nand ginst9266 (P2_ADD_391_1196_U90, P2_ADD_391_1196_U330, P2_ADD_391_1196_U331);
  nand ginst9267 (P2_ADD_391_1196_U91, P2_ADD_391_1196_U337, P2_ADD_391_1196_U338);
  nand ginst9268 (P2_ADD_391_1196_U92, P2_ADD_391_1196_U349, P2_ADD_391_1196_U350);
  nand ginst9269 (P2_ADD_391_1196_U93, P2_ADD_391_1196_U356, P2_ADD_391_1196_U357);
  nand ginst9270 (P2_ADD_391_1196_U94, P2_ADD_391_1196_U363, P2_ADD_391_1196_U364);
  nand ginst9271 (P2_ADD_391_1196_U95, P2_ADD_391_1196_U370, P2_ADD_391_1196_U371);
  nand ginst9272 (P2_ADD_391_1196_U96, P2_ADD_391_1196_U377, P2_ADD_391_1196_U378);
  nand ginst9273 (P2_ADD_391_1196_U97, P2_ADD_391_1196_U384, P2_ADD_391_1196_U385);
  nand ginst9274 (P2_ADD_391_1196_U98, P2_ADD_391_1196_U391, P2_ADD_391_1196_U392);
  nand ginst9275 (P2_ADD_391_1196_U99, P2_ADD_391_1196_U398, P2_ADD_391_1196_U399);
  nand ginst9276 (P2_ADD_394_U10, P2_INSTADDRPOINTER_REG_4__SCAN_IN, P2_ADD_394_U98);
  not ginst9277 (P2_ADD_394_U100, P2_ADD_394_U13);
  not ginst9278 (P2_ADD_394_U101, P2_ADD_394_U14);
  not ginst9279 (P2_ADD_394_U102, P2_ADD_394_U16);
  not ginst9280 (P2_ADD_394_U103, P2_ADD_394_U18);
  not ginst9281 (P2_ADD_394_U104, P2_ADD_394_U20);
  not ginst9282 (P2_ADD_394_U105, P2_ADD_394_U22);
  not ginst9283 (P2_ADD_394_U106, P2_ADD_394_U24);
  not ginst9284 (P2_ADD_394_U107, P2_ADD_394_U26);
  not ginst9285 (P2_ADD_394_U108, P2_ADD_394_U28);
  not ginst9286 (P2_ADD_394_U109, P2_ADD_394_U30);
  not ginst9287 (P2_ADD_394_U11, P2_INSTADDRPOINTER_REG_5__SCAN_IN);
  not ginst9288 (P2_ADD_394_U110, P2_ADD_394_U32);
  not ginst9289 (P2_ADD_394_U111, P2_ADD_394_U34);
  not ginst9290 (P2_ADD_394_U112, P2_ADD_394_U36);
  not ginst9291 (P2_ADD_394_U113, P2_ADD_394_U38);
  not ginst9292 (P2_ADD_394_U114, P2_ADD_394_U40);
  not ginst9293 (P2_ADD_394_U115, P2_ADD_394_U42);
  not ginst9294 (P2_ADD_394_U116, P2_ADD_394_U44);
  not ginst9295 (P2_ADD_394_U117, P2_ADD_394_U46);
  not ginst9296 (P2_ADD_394_U118, P2_ADD_394_U48);
  not ginst9297 (P2_ADD_394_U119, P2_ADD_394_U50);
  not ginst9298 (P2_ADD_394_U12, P2_INSTADDRPOINTER_REG_6__SCAN_IN);
  not ginst9299 (P2_ADD_394_U120, P2_ADD_394_U52);
  not ginst9300 (P2_ADD_394_U121, P2_ADD_394_U54);
  not ginst9301 (P2_ADD_394_U122, P2_ADD_394_U56);
  not ginst9302 (P2_ADD_394_U123, P2_ADD_394_U58);
  not ginst9303 (P2_ADD_394_U124, P2_ADD_394_U61);
  nand ginst9304 (P2_ADD_394_U125, P2_INSTADDRPOINTER_REG_0__SCAN_IN, P2_INSTADDRPOINTER_REG_1__SCAN_IN, P2_INSTADDRPOINTER_REG_2__SCAN_IN);
  not ginst9305 (P2_ADD_394_U126, P2_ADD_394_U93);
  nand ginst9306 (P2_ADD_394_U127, P2_INSTADDRPOINTER_REG_6__SCAN_IN, P2_ADD_394_U13);
  nand ginst9307 (P2_ADD_394_U128, P2_ADD_394_U100, P2_ADD_394_U12);
  nand ginst9308 (P2_ADD_394_U129, P2_INSTADDRPOINTER_REG_30__SCAN_IN, P2_ADD_394_U61);
  nand ginst9309 (P2_ADD_394_U13, P2_INSTADDRPOINTER_REG_5__SCAN_IN, P2_ADD_394_U99);
  nand ginst9310 (P2_ADD_394_U130, P2_ADD_394_U124, P2_ADD_394_U60);
  nand ginst9311 (P2_ADD_394_U131, P2_INSTADDRPOINTER_REG_29__SCAN_IN, P2_ADD_394_U58);
  nand ginst9312 (P2_ADD_394_U132, P2_ADD_394_U123, P2_ADD_394_U59);
  nand ginst9313 (P2_ADD_394_U133, P2_INSTADDRPOINTER_REG_24__SCAN_IN, P2_ADD_394_U48);
  nand ginst9314 (P2_ADD_394_U134, P2_ADD_394_U118, P2_ADD_394_U49);
  nand ginst9315 (P2_ADD_394_U135, P2_INSTADDRPOINTER_REG_17__SCAN_IN, P2_ADD_394_U34);
  nand ginst9316 (P2_ADD_394_U136, P2_ADD_394_U111, P2_ADD_394_U35);
  nand ginst9317 (P2_ADD_394_U137, P2_INSTADDRPOINTER_REG_20__SCAN_IN, P2_ADD_394_U40);
  nand ginst9318 (P2_ADD_394_U138, P2_ADD_394_U114, P2_ADD_394_U41);
  nand ginst9319 (P2_ADD_394_U139, P2_INSTADDRPOINTER_REG_13__SCAN_IN, P2_ADD_394_U26);
  nand ginst9320 (P2_ADD_394_U14, P2_INSTADDRPOINTER_REG_6__SCAN_IN, P2_ADD_394_U100);
  nand ginst9321 (P2_ADD_394_U140, P2_ADD_394_U107, P2_ADD_394_U27);
  nand ginst9322 (P2_ADD_394_U141, P2_INSTADDRPOINTER_REG_9__SCAN_IN, P2_ADD_394_U18);
  nand ginst9323 (P2_ADD_394_U142, P2_ADD_394_U103, P2_ADD_394_U19);
  nand ginst9324 (P2_ADD_394_U143, P2_INSTADDRPOINTER_REG_22__SCAN_IN, P2_ADD_394_U44);
  nand ginst9325 (P2_ADD_394_U144, P2_ADD_394_U116, P2_ADD_394_U45);
  nand ginst9326 (P2_ADD_394_U145, P2_INSTADDRPOINTER_REG_18__SCAN_IN, P2_ADD_394_U36);
  nand ginst9327 (P2_ADD_394_U146, P2_ADD_394_U112, P2_ADD_394_U37);
  nand ginst9328 (P2_ADD_394_U147, P2_INSTADDRPOINTER_REG_11__SCAN_IN, P2_ADD_394_U22);
  nand ginst9329 (P2_ADD_394_U148, P2_ADD_394_U105, P2_ADD_394_U23);
  nand ginst9330 (P2_ADD_394_U149, P2_INSTADDRPOINTER_REG_26__SCAN_IN, P2_ADD_394_U52);
  not ginst9331 (P2_ADD_394_U15, P2_INSTADDRPOINTER_REG_7__SCAN_IN);
  nand ginst9332 (P2_ADD_394_U150, P2_ADD_394_U120, P2_ADD_394_U53);
  nand ginst9333 (P2_ADD_394_U151, P2_INSTADDRPOINTER_REG_15__SCAN_IN, P2_ADD_394_U30);
  nand ginst9334 (P2_ADD_394_U152, P2_ADD_394_U109, P2_ADD_394_U31);
  nand ginst9335 (P2_ADD_394_U153, P2_INSTADDRPOINTER_REG_4__SCAN_IN, P2_ADD_394_U8);
  nand ginst9336 (P2_ADD_394_U154, P2_ADD_394_U9, P2_ADD_394_U98);
  nand ginst9337 (P2_ADD_394_U155, P2_INSTADDRPOINTER_REG_27__SCAN_IN, P2_ADD_394_U54);
  nand ginst9338 (P2_ADD_394_U156, P2_ADD_394_U121, P2_ADD_394_U55);
  nand ginst9339 (P2_ADD_394_U157, P2_INSTADDRPOINTER_REG_14__SCAN_IN, P2_ADD_394_U28);
  nand ginst9340 (P2_ADD_394_U158, P2_ADD_394_U108, P2_ADD_394_U29);
  nand ginst9341 (P2_ADD_394_U159, P2_INSTADDRPOINTER_REG_5__SCAN_IN, P2_ADD_394_U10);
  nand ginst9342 (P2_ADD_394_U16, P2_INSTADDRPOINTER_REG_7__SCAN_IN, P2_ADD_394_U101);
  nand ginst9343 (P2_ADD_394_U160, P2_ADD_394_U11, P2_ADD_394_U99);
  nand ginst9344 (P2_ADD_394_U161, P2_INSTADDRPOINTER_REG_8__SCAN_IN, P2_ADD_394_U16);
  nand ginst9345 (P2_ADD_394_U162, P2_ADD_394_U102, P2_ADD_394_U17);
  nand ginst9346 (P2_ADD_394_U163, P2_INSTADDRPOINTER_REG_23__SCAN_IN, P2_ADD_394_U46);
  nand ginst9347 (P2_ADD_394_U164, P2_ADD_394_U117, P2_ADD_394_U47);
  nand ginst9348 (P2_ADD_394_U165, P2_INSTADDRPOINTER_REG_19__SCAN_IN, P2_ADD_394_U38);
  nand ginst9349 (P2_ADD_394_U166, P2_ADD_394_U113, P2_ADD_394_U39);
  nand ginst9350 (P2_ADD_394_U167, P2_INSTADDRPOINTER_REG_10__SCAN_IN, P2_ADD_394_U20);
  nand ginst9351 (P2_ADD_394_U168, P2_ADD_394_U104, P2_ADD_394_U21);
  nand ginst9352 (P2_ADD_394_U169, P2_INSTADDRPOINTER_REG_31__SCAN_IN, P2_ADD_394_U93);
  not ginst9353 (P2_ADD_394_U17, P2_INSTADDRPOINTER_REG_8__SCAN_IN);
  nand ginst9354 (P2_ADD_394_U170, P2_ADD_394_U126, P2_ADD_394_U92);
  nand ginst9355 (P2_ADD_394_U171, P2_INSTADDRPOINTER_REG_3__SCAN_IN, P2_ADD_394_U94);
  nand ginst9356 (P2_ADD_394_U172, P2_ADD_394_U7, P2_ADD_394_U97);
  nand ginst9357 (P2_ADD_394_U173, P2_INSTADDRPOINTER_REG_1__SCAN_IN, P2_ADD_394_U4);
  nand ginst9358 (P2_ADD_394_U174, P2_INSTADDRPOINTER_REG_0__SCAN_IN, P2_ADD_394_U6);
  nand ginst9359 (P2_ADD_394_U175, P2_INSTADDRPOINTER_REG_28__SCAN_IN, P2_ADD_394_U56);
  nand ginst9360 (P2_ADD_394_U176, P2_ADD_394_U122, P2_ADD_394_U57);
  nand ginst9361 (P2_ADD_394_U177, P2_INSTADDRPOINTER_REG_21__SCAN_IN, P2_ADD_394_U42);
  nand ginst9362 (P2_ADD_394_U178, P2_ADD_394_U115, P2_ADD_394_U43);
  nand ginst9363 (P2_ADD_394_U179, P2_INSTADDRPOINTER_REG_12__SCAN_IN, P2_ADD_394_U24);
  nand ginst9364 (P2_ADD_394_U18, P2_INSTADDRPOINTER_REG_8__SCAN_IN, P2_ADD_394_U102);
  nand ginst9365 (P2_ADD_394_U180, P2_ADD_394_U106, P2_ADD_394_U25);
  nand ginst9366 (P2_ADD_394_U181, P2_INSTADDRPOINTER_REG_7__SCAN_IN, P2_ADD_394_U14);
  nand ginst9367 (P2_ADD_394_U182, P2_ADD_394_U101, P2_ADD_394_U15);
  nand ginst9368 (P2_ADD_394_U183, P2_INSTADDRPOINTER_REG_25__SCAN_IN, P2_ADD_394_U50);
  nand ginst9369 (P2_ADD_394_U184, P2_ADD_394_U119, P2_ADD_394_U51);
  nand ginst9370 (P2_ADD_394_U185, P2_INSTADDRPOINTER_REG_16__SCAN_IN, P2_ADD_394_U32);
  nand ginst9371 (P2_ADD_394_U186, P2_ADD_394_U110, P2_ADD_394_U33);
  not ginst9372 (P2_ADD_394_U19, P2_INSTADDRPOINTER_REG_9__SCAN_IN);
  nand ginst9373 (P2_ADD_394_U20, P2_INSTADDRPOINTER_REG_9__SCAN_IN, P2_ADD_394_U103);
  not ginst9374 (P2_ADD_394_U21, P2_INSTADDRPOINTER_REG_10__SCAN_IN);
  nand ginst9375 (P2_ADD_394_U22, P2_INSTADDRPOINTER_REG_10__SCAN_IN, P2_ADD_394_U104);
  not ginst9376 (P2_ADD_394_U23, P2_INSTADDRPOINTER_REG_11__SCAN_IN);
  nand ginst9377 (P2_ADD_394_U24, P2_INSTADDRPOINTER_REG_11__SCAN_IN, P2_ADD_394_U105);
  not ginst9378 (P2_ADD_394_U25, P2_INSTADDRPOINTER_REG_12__SCAN_IN);
  nand ginst9379 (P2_ADD_394_U26, P2_INSTADDRPOINTER_REG_12__SCAN_IN, P2_ADD_394_U106);
  not ginst9380 (P2_ADD_394_U27, P2_INSTADDRPOINTER_REG_13__SCAN_IN);
  nand ginst9381 (P2_ADD_394_U28, P2_INSTADDRPOINTER_REG_13__SCAN_IN, P2_ADD_394_U107);
  not ginst9382 (P2_ADD_394_U29, P2_INSTADDRPOINTER_REG_14__SCAN_IN);
  nand ginst9383 (P2_ADD_394_U30, P2_INSTADDRPOINTER_REG_14__SCAN_IN, P2_ADD_394_U108);
  not ginst9384 (P2_ADD_394_U31, P2_INSTADDRPOINTER_REG_15__SCAN_IN);
  nand ginst9385 (P2_ADD_394_U32, P2_INSTADDRPOINTER_REG_15__SCAN_IN, P2_ADD_394_U109);
  not ginst9386 (P2_ADD_394_U33, P2_INSTADDRPOINTER_REG_16__SCAN_IN);
  nand ginst9387 (P2_ADD_394_U34, P2_INSTADDRPOINTER_REG_16__SCAN_IN, P2_ADD_394_U110);
  not ginst9388 (P2_ADD_394_U35, P2_INSTADDRPOINTER_REG_17__SCAN_IN);
  nand ginst9389 (P2_ADD_394_U36, P2_INSTADDRPOINTER_REG_17__SCAN_IN, P2_ADD_394_U111);
  not ginst9390 (P2_ADD_394_U37, P2_INSTADDRPOINTER_REG_18__SCAN_IN);
  nand ginst9391 (P2_ADD_394_U38, P2_INSTADDRPOINTER_REG_18__SCAN_IN, P2_ADD_394_U112);
  not ginst9392 (P2_ADD_394_U39, P2_INSTADDRPOINTER_REG_19__SCAN_IN);
  not ginst9393 (P2_ADD_394_U4, P2_INSTADDRPOINTER_REG_0__SCAN_IN);
  nand ginst9394 (P2_ADD_394_U40, P2_INSTADDRPOINTER_REG_19__SCAN_IN, P2_ADD_394_U113);
  not ginst9395 (P2_ADD_394_U41, P2_INSTADDRPOINTER_REG_20__SCAN_IN);
  nand ginst9396 (P2_ADD_394_U42, P2_INSTADDRPOINTER_REG_20__SCAN_IN, P2_ADD_394_U114);
  not ginst9397 (P2_ADD_394_U43, P2_INSTADDRPOINTER_REG_21__SCAN_IN);
  nand ginst9398 (P2_ADD_394_U44, P2_INSTADDRPOINTER_REG_21__SCAN_IN, P2_ADD_394_U115);
  not ginst9399 (P2_ADD_394_U45, P2_INSTADDRPOINTER_REG_22__SCAN_IN);
  nand ginst9400 (P2_ADD_394_U46, P2_INSTADDRPOINTER_REG_22__SCAN_IN, P2_ADD_394_U116);
  not ginst9401 (P2_ADD_394_U47, P2_INSTADDRPOINTER_REG_23__SCAN_IN);
  nand ginst9402 (P2_ADD_394_U48, P2_INSTADDRPOINTER_REG_23__SCAN_IN, P2_ADD_394_U117);
  not ginst9403 (P2_ADD_394_U49, P2_INSTADDRPOINTER_REG_24__SCAN_IN);
  nand ginst9404 (P2_ADD_394_U5, P2_ADD_394_U125, P2_ADD_394_U94);
  nand ginst9405 (P2_ADD_394_U50, P2_INSTADDRPOINTER_REG_24__SCAN_IN, P2_ADD_394_U118);
  not ginst9406 (P2_ADD_394_U51, P2_INSTADDRPOINTER_REG_25__SCAN_IN);
  nand ginst9407 (P2_ADD_394_U52, P2_INSTADDRPOINTER_REG_25__SCAN_IN, P2_ADD_394_U119);
  not ginst9408 (P2_ADD_394_U53, P2_INSTADDRPOINTER_REG_26__SCAN_IN);
  nand ginst9409 (P2_ADD_394_U54, P2_INSTADDRPOINTER_REG_26__SCAN_IN, P2_ADD_394_U120);
  not ginst9410 (P2_ADD_394_U55, P2_INSTADDRPOINTER_REG_27__SCAN_IN);
  nand ginst9411 (P2_ADD_394_U56, P2_INSTADDRPOINTER_REG_27__SCAN_IN, P2_ADD_394_U121);
  not ginst9412 (P2_ADD_394_U57, P2_INSTADDRPOINTER_REG_28__SCAN_IN);
  nand ginst9413 (P2_ADD_394_U58, P2_INSTADDRPOINTER_REG_28__SCAN_IN, P2_ADD_394_U122);
  not ginst9414 (P2_ADD_394_U59, P2_INSTADDRPOINTER_REG_29__SCAN_IN);
  not ginst9415 (P2_ADD_394_U6, P2_INSTADDRPOINTER_REG_1__SCAN_IN);
  not ginst9416 (P2_ADD_394_U60, P2_INSTADDRPOINTER_REG_30__SCAN_IN);
  nand ginst9417 (P2_ADD_394_U61, P2_INSTADDRPOINTER_REG_29__SCAN_IN, P2_ADD_394_U123);
  not ginst9418 (P2_ADD_394_U62, P2_INSTADDRPOINTER_REG_2__SCAN_IN);
  nand ginst9419 (P2_ADD_394_U63, P2_ADD_394_U127, P2_ADD_394_U128);
  nand ginst9420 (P2_ADD_394_U64, P2_ADD_394_U129, P2_ADD_394_U130);
  nand ginst9421 (P2_ADD_394_U65, P2_ADD_394_U131, P2_ADD_394_U132);
  nand ginst9422 (P2_ADD_394_U66, P2_ADD_394_U133, P2_ADD_394_U134);
  nand ginst9423 (P2_ADD_394_U67, P2_ADD_394_U135, P2_ADD_394_U136);
  nand ginst9424 (P2_ADD_394_U68, P2_ADD_394_U137, P2_ADD_394_U138);
  nand ginst9425 (P2_ADD_394_U69, P2_ADD_394_U139, P2_ADD_394_U140);
  not ginst9426 (P2_ADD_394_U7, P2_INSTADDRPOINTER_REG_3__SCAN_IN);
  nand ginst9427 (P2_ADD_394_U70, P2_ADD_394_U141, P2_ADD_394_U142);
  nand ginst9428 (P2_ADD_394_U71, P2_ADD_394_U143, P2_ADD_394_U144);
  nand ginst9429 (P2_ADD_394_U72, P2_ADD_394_U145, P2_ADD_394_U146);
  nand ginst9430 (P2_ADD_394_U73, P2_ADD_394_U147, P2_ADD_394_U148);
  nand ginst9431 (P2_ADD_394_U74, P2_ADD_394_U149, P2_ADD_394_U150);
  nand ginst9432 (P2_ADD_394_U75, P2_ADD_394_U151, P2_ADD_394_U152);
  nand ginst9433 (P2_ADD_394_U76, P2_ADD_394_U153, P2_ADD_394_U154);
  nand ginst9434 (P2_ADD_394_U77, P2_ADD_394_U155, P2_ADD_394_U156);
  nand ginst9435 (P2_ADD_394_U78, P2_ADD_394_U157, P2_ADD_394_U158);
  nand ginst9436 (P2_ADD_394_U79, P2_ADD_394_U159, P2_ADD_394_U160);
  nand ginst9437 (P2_ADD_394_U8, P2_INSTADDRPOINTER_REG_3__SCAN_IN, P2_ADD_394_U94);
  nand ginst9438 (P2_ADD_394_U80, P2_ADD_394_U161, P2_ADD_394_U162);
  nand ginst9439 (P2_ADD_394_U81, P2_ADD_394_U163, P2_ADD_394_U164);
  nand ginst9440 (P2_ADD_394_U82, P2_ADD_394_U165, P2_ADD_394_U166);
  nand ginst9441 (P2_ADD_394_U83, P2_ADD_394_U167, P2_ADD_394_U168);
  nand ginst9442 (P2_ADD_394_U84, P2_ADD_394_U169, P2_ADD_394_U170);
  nand ginst9443 (P2_ADD_394_U85, P2_ADD_394_U173, P2_ADD_394_U174);
  nand ginst9444 (P2_ADD_394_U86, P2_ADD_394_U175, P2_ADD_394_U176);
  nand ginst9445 (P2_ADD_394_U87, P2_ADD_394_U177, P2_ADD_394_U178);
  nand ginst9446 (P2_ADD_394_U88, P2_ADD_394_U179, P2_ADD_394_U180);
  nand ginst9447 (P2_ADD_394_U89, P2_ADD_394_U181, P2_ADD_394_U182);
  not ginst9448 (P2_ADD_394_U9, P2_INSTADDRPOINTER_REG_4__SCAN_IN);
  nand ginst9449 (P2_ADD_394_U90, P2_ADD_394_U183, P2_ADD_394_U184);
  nand ginst9450 (P2_ADD_394_U91, P2_ADD_394_U185, P2_ADD_394_U186);
  not ginst9451 (P2_ADD_394_U92, P2_INSTADDRPOINTER_REG_31__SCAN_IN);
  nand ginst9452 (P2_ADD_394_U93, P2_INSTADDRPOINTER_REG_30__SCAN_IN, P2_ADD_394_U124);
  nand ginst9453 (P2_ADD_394_U94, P2_ADD_394_U62, P2_ADD_394_U96);
  and ginst9454 (P2_ADD_394_U95, P2_ADD_394_U171, P2_ADD_394_U172);
  nand ginst9455 (P2_ADD_394_U96, P2_INSTADDRPOINTER_REG_0__SCAN_IN, P2_INSTADDRPOINTER_REG_1__SCAN_IN);
  not ginst9456 (P2_ADD_394_U97, P2_ADD_394_U94);
  not ginst9457 (P2_ADD_394_U98, P2_ADD_394_U8);
  not ginst9458 (P2_ADD_394_U99, P2_ADD_394_U10);
  nand ginst9459 (P2_ADD_402_1132_U10, P2_ADD_402_1132_U29, P2_U2593);
  not ginst9460 (P2_ADD_402_1132_U11, P2_U2594);
  nand ginst9461 (P2_ADD_402_1132_U12, P2_ADD_402_1132_U30, P2_U2594);
  not ginst9462 (P2_ADD_402_1132_U13, P2_U2595);
  nand ginst9463 (P2_ADD_402_1132_U14, P2_ADD_402_1132_U31, P2_U2595);
  not ginst9464 (P2_ADD_402_1132_U15, P2_U2596);
  nand ginst9465 (P2_ADD_402_1132_U16, P2_ADD_402_1132_U32, P2_U2596);
  not ginst9466 (P2_ADD_402_1132_U17, P2_U2597);
  nand ginst9467 (P2_ADD_402_1132_U18, P2_ADD_402_1132_U35, P2_ADD_402_1132_U36);
  nand ginst9468 (P2_ADD_402_1132_U19, P2_ADD_402_1132_U37, P2_ADD_402_1132_U38);
  nand ginst9469 (P2_ADD_402_1132_U20, P2_ADD_402_1132_U39, P2_ADD_402_1132_U40);
  nand ginst9470 (P2_ADD_402_1132_U21, P2_ADD_402_1132_U41, P2_ADD_402_1132_U42);
  nand ginst9471 (P2_ADD_402_1132_U22, P2_ADD_402_1132_U43, P2_ADD_402_1132_U44);
  nand ginst9472 (P2_ADD_402_1132_U23, P2_ADD_402_1132_U45, P2_ADD_402_1132_U46);
  nand ginst9473 (P2_ADD_402_1132_U24, P2_ADD_402_1132_U47, P2_ADD_402_1132_U48);
  nand ginst9474 (P2_ADD_402_1132_U25, P2_ADD_402_1132_U49, P2_ADD_402_1132_U50);
  not ginst9475 (P2_ADD_402_1132_U26, P2_U2598);
  nand ginst9476 (P2_ADD_402_1132_U27, P2_ADD_402_1132_U33, P2_U2597);
  not ginst9477 (P2_ADD_402_1132_U28, P2_ADD_402_1132_U6);
  not ginst9478 (P2_ADD_402_1132_U29, P2_ADD_402_1132_U8);
  not ginst9479 (P2_ADD_402_1132_U30, P2_ADD_402_1132_U10);
  not ginst9480 (P2_ADD_402_1132_U31, P2_ADD_402_1132_U12);
  not ginst9481 (P2_ADD_402_1132_U32, P2_ADD_402_1132_U14);
  not ginst9482 (P2_ADD_402_1132_U33, P2_ADD_402_1132_U16);
  not ginst9483 (P2_ADD_402_1132_U34, P2_ADD_402_1132_U27);
  nand ginst9484 (P2_ADD_402_1132_U35, P2_ADD_402_1132_U27, P2_U2598);
  nand ginst9485 (P2_ADD_402_1132_U36, P2_ADD_402_1132_U26, P2_ADD_402_1132_U34);
  nand ginst9486 (P2_ADD_402_1132_U37, P2_ADD_402_1132_U16, P2_U2597);
  nand ginst9487 (P2_ADD_402_1132_U38, P2_ADD_402_1132_U17, P2_ADD_402_1132_U33);
  nand ginst9488 (P2_ADD_402_1132_U39, P2_ADD_402_1132_U6, P2_U2592);
  not ginst9489 (P2_ADD_402_1132_U4, P2_U2606);
  nand ginst9490 (P2_ADD_402_1132_U40, P2_ADD_402_1132_U28, P2_ADD_402_1132_U7);
  nand ginst9491 (P2_ADD_402_1132_U41, P2_ADD_402_1132_U10, P2_U2594);
  nand ginst9492 (P2_ADD_402_1132_U42, P2_ADD_402_1132_U11, P2_ADD_402_1132_U30);
  nand ginst9493 (P2_ADD_402_1132_U43, P2_ADD_402_1132_U12, P2_U2595);
  nand ginst9494 (P2_ADD_402_1132_U44, P2_ADD_402_1132_U13, P2_ADD_402_1132_U31);
  nand ginst9495 (P2_ADD_402_1132_U45, P2_ADD_402_1132_U4, P2_U2591);
  nand ginst9496 (P2_ADD_402_1132_U46, P2_ADD_402_1132_U5, P2_U2606);
  nand ginst9497 (P2_ADD_402_1132_U47, P2_ADD_402_1132_U14, P2_U2596);
  nand ginst9498 (P2_ADD_402_1132_U48, P2_ADD_402_1132_U15, P2_ADD_402_1132_U32);
  nand ginst9499 (P2_ADD_402_1132_U49, P2_ADD_402_1132_U8, P2_U2593);
  not ginst9500 (P2_ADD_402_1132_U5, P2_U2591);
  nand ginst9501 (P2_ADD_402_1132_U50, P2_ADD_402_1132_U29, P2_ADD_402_1132_U9);
  nand ginst9502 (P2_ADD_402_1132_U6, P2_U2591, P2_U2606);
  not ginst9503 (P2_ADD_402_1132_U7, P2_U2592);
  nand ginst9504 (P2_ADD_402_1132_U8, P2_ADD_402_1132_U28, P2_U2592);
  not ginst9505 (P2_ADD_402_1132_U9, P2_U2593);
  nor ginst9506 (P2_GTE_370_U6, P2_GTE_370_U8, P2_R2219_U25);
  and ginst9507 (P2_GTE_370_U7, P2_GTE_370_U9, P2_R2219_U29);
  nor ginst9508 (P2_GTE_370_U8, P2_GTE_370_U7, P2_R2219_U26, P2_R2219_U27, P2_R2219_U28);
  or ginst9509 (P2_GTE_370_U9, P2_R2219_U30, P2_R2219_U8);
  or ginst9510 (P2_LT_563_1260_U6, P2_LT_563_1260_U7, P2_U3617);
  nor ginst9511 (P2_LT_563_1260_U7, P2_SUB_563_U6, P2_SUB_563_U7);
  not ginst9512 (P2_LT_563_U10, P2_U3619);
  not ginst9513 (P2_LT_563_U11, P2_U3618);
  not ginst9514 (P2_LT_563_U12, P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN);
  not ginst9515 (P2_LT_563_U13, P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN);
  not ginst9516 (P2_LT_563_U14, P2_U3617);
  not ginst9517 (P2_LT_563_U15, P2_U3621);
  nand ginst9518 (P2_LT_563_U16, P2_LT_563_U8, P2_U3620);
  nand ginst9519 (P2_LT_563_U17, P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P2_LT_563_U15, P2_LT_563_U16);
  nand ginst9520 (P2_LT_563_U18, P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN, P2_LT_563_U7);
  nand ginst9521 (P2_LT_563_U19, P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN, P2_LT_563_U10);
  nand ginst9522 (P2_LT_563_U20, P2_LT_563_U17, P2_LT_563_U18, P2_LT_563_U19);
  nand ginst9523 (P2_LT_563_U21, P2_LT_563_U9, P2_U3619);
  nand ginst9524 (P2_LT_563_U22, P2_LT_563_U12, P2_U3618);
  nand ginst9525 (P2_LT_563_U23, P2_LT_563_U20, P2_LT_563_U21, P2_LT_563_U22);
  nand ginst9526 (P2_LT_563_U24, P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN, P2_LT_563_U11);
  nand ginst9527 (P2_LT_563_U25, P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN, P2_LT_563_U14);
  nand ginst9528 (P2_LT_563_U26, P2_LT_563_U23, P2_LT_563_U24, P2_LT_563_U25);
  nand ginst9529 (P2_LT_563_U27, P2_LT_563_U13, P2_U3617);
  and ginst9530 (P2_LT_563_U6, P2_LT_563_U26, P2_LT_563_U27);
  not ginst9531 (P2_LT_563_U7, P2_U3620);
  not ginst9532 (P2_LT_563_U8, P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN);
  not ginst9533 (P2_LT_563_U9, P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN);
  and ginst9534 (P2_R1957_U10, P2_R1957_U118, P2_R1957_U31);
  not ginst9535 (P2_R1957_U100, P2_R1957_U34);
  not ginst9536 (P2_R1957_U101, P2_R1957_U35);
  not ginst9537 (P2_R1957_U102, P2_R1957_U36);
  not ginst9538 (P2_R1957_U103, P2_R1957_U37);
  or ginst9539 (P2_R1957_U104, P2_U3682, P2_U3683);
  nand ginst9540 (P2_R1957_U105, P2_R1957_U104, P2_U3671);
  nand ginst9541 (P2_R1957_U106, P2_R1957_U36, P2_U3661);
  nand ginst9542 (P2_R1957_U107, P2_R1957_U101, P2_R1957_U63);
  nand ginst9543 (P2_R1957_U108, P2_R1957_U107, P2_U3662);
  nand ginst9544 (P2_R1957_U109, P2_R1957_U100, P2_R1957_U65);
  and ginst9545 (P2_R1957_U11, P2_R1957_U116, P2_R1957_U32);
  nand ginst9546 (P2_R1957_U110, P2_R1957_U109, P2_U3664);
  nand ginst9547 (P2_R1957_U111, P2_R1957_U67, P2_R1957_U99);
  nand ginst9548 (P2_R1957_U112, P2_R1957_U111, P2_U3666);
  nand ginst9549 (P2_R1957_U113, P2_R1957_U69, P2_R1957_U98);
  nand ginst9550 (P2_R1957_U114, P2_R1957_U113, P2_U3668);
  nand ginst9551 (P2_R1957_U115, P2_R1957_U73, P2_R1957_U97);
  nand ginst9552 (P2_R1957_U116, P2_R1957_U115, P2_U3670);
  nand ginst9553 (P2_R1957_U117, P2_R1957_U75, P2_R1957_U96);
  nand ginst9554 (P2_R1957_U118, P2_R1957_U117, P2_U3673);
  nand ginst9555 (P2_R1957_U119, P2_R1957_U77, P2_R1957_U95);
  and ginst9556 (P2_R1957_U12, P2_R1957_U114, P2_R1957_U33);
  nand ginst9557 (P2_R1957_U120, P2_R1957_U119, P2_U3675);
  nand ginst9558 (P2_R1957_U121, P2_R1957_U79, P2_R1957_U94);
  nand ginst9559 (P2_R1957_U122, P2_R1957_U121, P2_U3677);
  nand ginst9560 (P2_R1957_U123, P2_R1957_U81, P2_R1957_U93);
  nand ginst9561 (P2_R1957_U124, P2_R1957_U123, P2_U3679);
  nand ginst9562 (P2_R1957_U125, P2_R1957_U52, P2_R1957_U86);
  nand ginst9563 (P2_R1957_U126, P2_R1957_U125, P2_U3681);
  nand ginst9564 (P2_R1957_U127, P2_R1957_U103, P2_R1957_U61);
  nand ginst9565 (P2_R1957_U128, P2_R1957_U24, P2_U3653);
  nand ginst9566 (P2_R1957_U129, P2_R1957_U52, P2_R1957_U86);
  and ginst9567 (P2_R1957_U13, P2_R1957_U112, P2_R1957_U34);
  nand ginst9568 (P2_R1957_U130, P2_R1957_U23, P2_U3655);
  nand ginst9569 (P2_R1957_U131, P2_R1957_U54, P2_R1957_U85);
  nand ginst9570 (P2_R1957_U132, P2_R1957_U22, P2_U3657);
  nand ginst9571 (P2_R1957_U133, P2_R1957_U56, P2_R1957_U84);
  nand ginst9572 (P2_R1957_U134, P2_R1957_U21, P2_U3660);
  nand ginst9573 (P2_R1957_U135, P2_R1957_U58, P2_R1957_U83);
  nand ginst9574 (P2_R1957_U136, P2_R1957_U127, P2_R1957_U60);
  nand ginst9575 (P2_R1957_U137, P2_R1957_U103, P2_R1957_U61, P2_U3647);
  nand ginst9576 (P2_R1957_U138, P2_R1957_U37, P2_U3659);
  nand ginst9577 (P2_R1957_U139, P2_R1957_U103, P2_R1957_U61);
  and ginst9578 (P2_R1957_U14, P2_R1957_U110, P2_R1957_U35);
  nand ginst9579 (P2_R1957_U140, P2_R1957_U35, P2_U3663);
  nand ginst9580 (P2_R1957_U141, P2_R1957_U101, P2_R1957_U63);
  nand ginst9581 (P2_R1957_U142, P2_R1957_U34, P2_U3665);
  nand ginst9582 (P2_R1957_U143, P2_R1957_U100, P2_R1957_U65);
  nand ginst9583 (P2_R1957_U144, P2_R1957_U33, P2_U3667);
  nand ginst9584 (P2_R1957_U145, P2_R1957_U67, P2_R1957_U99);
  nand ginst9585 (P2_R1957_U146, P2_R1957_U32, P2_U3669);
  nand ginst9586 (P2_R1957_U147, P2_R1957_U69, P2_R1957_U98);
  nand ginst9587 (P2_R1957_U148, P2_R1957_U72, P2_U3682);
  nand ginst9588 (P2_R1957_U149, P2_R1957_U71, P2_U3683);
  and ginst9589 (P2_R1957_U15, P2_R1957_U108, P2_R1957_U36);
  nand ginst9590 (P2_R1957_U150, P2_R1957_U31, P2_U3672);
  nand ginst9591 (P2_R1957_U151, P2_R1957_U73, P2_R1957_U97);
  nand ginst9592 (P2_R1957_U152, P2_R1957_U30, P2_U3674);
  nand ginst9593 (P2_R1957_U153, P2_R1957_U75, P2_R1957_U96);
  nand ginst9594 (P2_R1957_U154, P2_R1957_U29, P2_U3676);
  nand ginst9595 (P2_R1957_U155, P2_R1957_U77, P2_R1957_U95);
  nand ginst9596 (P2_R1957_U156, P2_R1957_U28, P2_U3678);
  nand ginst9597 (P2_R1957_U157, P2_R1957_U79, P2_R1957_U94);
  nand ginst9598 (P2_R1957_U158, P2_R1957_U27, P2_U3680);
  nand ginst9599 (P2_R1957_U159, P2_R1957_U81, P2_R1957_U93);
  and ginst9600 (P2_R1957_U16, P2_R1957_U106, P2_R1957_U37);
  and ginst9601 (P2_R1957_U17, P2_R1957_U105, P2_R1957_U21);
  and ginst9602 (P2_R1957_U18, P2_R1957_U22, P2_R1957_U92);
  and ginst9603 (P2_R1957_U19, P2_R1957_U23, P2_R1957_U90);
  and ginst9604 (P2_R1957_U20, P2_R1957_U24, P2_R1957_U88);
  or ginst9605 (P2_R1957_U21, P2_U3671, P2_U3682, P2_U3683);
  nand ginst9606 (P2_R1957_U22, P2_R1957_U51, P2_R1957_U83);
  nand ginst9607 (P2_R1957_U23, P2_R1957_U26, P2_R1957_U56, P2_R1957_U84);
  nand ginst9608 (P2_R1957_U24, P2_R1957_U25, P2_R1957_U54, P2_R1957_U85);
  not ginst9609 (P2_R1957_U25, P2_U3654);
  not ginst9610 (P2_R1957_U26, P2_U3656);
  nand ginst9611 (P2_R1957_U27, P2_R1957_U48, P2_R1957_U52, P2_R1957_U86);
  nand ginst9612 (P2_R1957_U28, P2_R1957_U47, P2_R1957_U81, P2_R1957_U93);
  nand ginst9613 (P2_R1957_U29, P2_R1957_U46, P2_R1957_U79, P2_R1957_U94);
  nand ginst9614 (P2_R1957_U30, P2_R1957_U45, P2_R1957_U77, P2_R1957_U95);
  nand ginst9615 (P2_R1957_U31, P2_R1957_U44, P2_R1957_U75, P2_R1957_U96);
  nand ginst9616 (P2_R1957_U32, P2_R1957_U43, P2_R1957_U73, P2_R1957_U97);
  nand ginst9617 (P2_R1957_U33, P2_R1957_U42, P2_R1957_U69, P2_R1957_U98);
  nand ginst9618 (P2_R1957_U34, P2_R1957_U41, P2_R1957_U67, P2_R1957_U99);
  nand ginst9619 (P2_R1957_U35, P2_R1957_U100, P2_R1957_U40, P2_R1957_U65);
  nand ginst9620 (P2_R1957_U36, P2_R1957_U101, P2_R1957_U39, P2_R1957_U63);
  nand ginst9621 (P2_R1957_U37, P2_R1957_U102, P2_R1957_U38);
  not ginst9622 (P2_R1957_U38, P2_U3661);
  not ginst9623 (P2_R1957_U39, P2_U3662);
  not ginst9624 (P2_R1957_U40, P2_U3664);
  not ginst9625 (P2_R1957_U41, P2_U3666);
  not ginst9626 (P2_R1957_U42, P2_U3668);
  not ginst9627 (P2_R1957_U43, P2_U3670);
  not ginst9628 (P2_R1957_U44, P2_U3673);
  not ginst9629 (P2_R1957_U45, P2_U3675);
  not ginst9630 (P2_R1957_U46, P2_U3677);
  not ginst9631 (P2_R1957_U47, P2_U3679);
  not ginst9632 (P2_R1957_U48, P2_U3681);
  nand ginst9633 (P2_R1957_U49, P2_R1957_U148, P2_R1957_U149);
  nand ginst9634 (P2_R1957_U50, P2_R1957_U136, P2_R1957_U137);
  nor ginst9635 (P2_R1957_U51, P2_U3658, P2_U3660);
  not ginst9636 (P2_R1957_U52, P2_U3653);
  and ginst9637 (P2_R1957_U53, P2_R1957_U128, P2_R1957_U129);
  not ginst9638 (P2_R1957_U54, P2_U3655);
  and ginst9639 (P2_R1957_U55, P2_R1957_U130, P2_R1957_U131);
  not ginst9640 (P2_R1957_U56, P2_U3657);
  and ginst9641 (P2_R1957_U57, P2_R1957_U132, P2_R1957_U133);
  not ginst9642 (P2_R1957_U58, P2_U3660);
  and ginst9643 (P2_R1957_U59, P2_R1957_U134, P2_R1957_U135);
  and ginst9644 (P2_R1957_U6, P2_R1957_U126, P2_R1957_U27);
  not ginst9645 (P2_R1957_U60, P2_U3647);
  not ginst9646 (P2_R1957_U61, P2_U3659);
  and ginst9647 (P2_R1957_U62, P2_R1957_U138, P2_R1957_U139);
  not ginst9648 (P2_R1957_U63, P2_U3663);
  and ginst9649 (P2_R1957_U64, P2_R1957_U140, P2_R1957_U141);
  not ginst9650 (P2_R1957_U65, P2_U3665);
  and ginst9651 (P2_R1957_U66, P2_R1957_U142, P2_R1957_U143);
  not ginst9652 (P2_R1957_U67, P2_U3667);
  and ginst9653 (P2_R1957_U68, P2_R1957_U144, P2_R1957_U145);
  not ginst9654 (P2_R1957_U69, P2_U3669);
  and ginst9655 (P2_R1957_U7, P2_R1957_U124, P2_R1957_U28);
  and ginst9656 (P2_R1957_U70, P2_R1957_U146, P2_R1957_U147);
  not ginst9657 (P2_R1957_U71, P2_U3682);
  not ginst9658 (P2_R1957_U72, P2_U3683);
  not ginst9659 (P2_R1957_U73, P2_U3672);
  and ginst9660 (P2_R1957_U74, P2_R1957_U150, P2_R1957_U151);
  not ginst9661 (P2_R1957_U75, P2_U3674);
  and ginst9662 (P2_R1957_U76, P2_R1957_U152, P2_R1957_U153);
  not ginst9663 (P2_R1957_U77, P2_U3676);
  and ginst9664 (P2_R1957_U78, P2_R1957_U154, P2_R1957_U155);
  not ginst9665 (P2_R1957_U79, P2_U3678);
  and ginst9666 (P2_R1957_U8, P2_R1957_U122, P2_R1957_U29);
  and ginst9667 (P2_R1957_U80, P2_R1957_U156, P2_R1957_U157);
  not ginst9668 (P2_R1957_U81, P2_U3680);
  and ginst9669 (P2_R1957_U82, P2_R1957_U158, P2_R1957_U159);
  not ginst9670 (P2_R1957_U83, P2_R1957_U21);
  not ginst9671 (P2_R1957_U84, P2_R1957_U22);
  not ginst9672 (P2_R1957_U85, P2_R1957_U23);
  not ginst9673 (P2_R1957_U86, P2_R1957_U24);
  nand ginst9674 (P2_R1957_U87, P2_R1957_U54, P2_R1957_U85);
  nand ginst9675 (P2_R1957_U88, P2_R1957_U87, P2_U3654);
  nand ginst9676 (P2_R1957_U89, P2_R1957_U56, P2_R1957_U84);
  and ginst9677 (P2_R1957_U9, P2_R1957_U120, P2_R1957_U30);
  nand ginst9678 (P2_R1957_U90, P2_R1957_U89, P2_U3656);
  nand ginst9679 (P2_R1957_U91, P2_R1957_U58, P2_R1957_U83);
  nand ginst9680 (P2_R1957_U92, P2_R1957_U91, P2_U3658);
  not ginst9681 (P2_R1957_U93, P2_R1957_U27);
  not ginst9682 (P2_R1957_U94, P2_R1957_U28);
  not ginst9683 (P2_R1957_U95, P2_R1957_U29);
  not ginst9684 (P2_R1957_U96, P2_R1957_U30);
  not ginst9685 (P2_R1957_U97, P2_R1957_U31);
  not ginst9686 (P2_R1957_U98, P2_R1957_U32);
  not ginst9687 (P2_R1957_U99, P2_R1957_U33);
  not ginst9688 (P2_R2027_U10, P2_INSTADDRPOINTER_REG_3__SCAN_IN);
  not ginst9689 (P2_R2027_U100, P2_R2027_U11);
  not ginst9690 (P2_R2027_U101, P2_R2027_U13);
  not ginst9691 (P2_R2027_U102, P2_R2027_U15);
  not ginst9692 (P2_R2027_U103, P2_R2027_U17);
  not ginst9693 (P2_R2027_U104, P2_R2027_U19);
  not ginst9694 (P2_R2027_U105, P2_R2027_U22);
  not ginst9695 (P2_R2027_U106, P2_R2027_U23);
  not ginst9696 (P2_R2027_U107, P2_R2027_U25);
  not ginst9697 (P2_R2027_U108, P2_R2027_U27);
  not ginst9698 (P2_R2027_U109, P2_R2027_U29);
  nand ginst9699 (P2_R2027_U11, P2_INSTADDRPOINTER_REG_3__SCAN_IN, P2_R2027_U99);
  not ginst9700 (P2_R2027_U110, P2_R2027_U31);
  not ginst9701 (P2_R2027_U111, P2_R2027_U33);
  not ginst9702 (P2_R2027_U112, P2_R2027_U35);
  not ginst9703 (P2_R2027_U113, P2_R2027_U37);
  not ginst9704 (P2_R2027_U114, P2_R2027_U39);
  not ginst9705 (P2_R2027_U115, P2_R2027_U41);
  not ginst9706 (P2_R2027_U116, P2_R2027_U43);
  not ginst9707 (P2_R2027_U117, P2_R2027_U45);
  not ginst9708 (P2_R2027_U118, P2_R2027_U47);
  not ginst9709 (P2_R2027_U119, P2_R2027_U49);
  not ginst9710 (P2_R2027_U12, P2_INSTADDRPOINTER_REG_4__SCAN_IN);
  not ginst9711 (P2_R2027_U120, P2_R2027_U51);
  not ginst9712 (P2_R2027_U121, P2_R2027_U53);
  not ginst9713 (P2_R2027_U122, P2_R2027_U55);
  not ginst9714 (P2_R2027_U123, P2_R2027_U57);
  not ginst9715 (P2_R2027_U124, P2_R2027_U59);
  not ginst9716 (P2_R2027_U125, P2_R2027_U61);
  not ginst9717 (P2_R2027_U126, P2_R2027_U63);
  not ginst9718 (P2_R2027_U127, P2_R2027_U97);
  nand ginst9719 (P2_R2027_U128, P2_INSTADDRPOINTER_REG_9__SCAN_IN, P2_R2027_U22);
  nand ginst9720 (P2_R2027_U129, P2_R2027_U105, P2_R2027_U21);
  nand ginst9721 (P2_R2027_U13, P2_INSTADDRPOINTER_REG_4__SCAN_IN, P2_R2027_U100);
  nand ginst9722 (P2_R2027_U130, P2_INSTADDRPOINTER_REG_8__SCAN_IN, P2_R2027_U19);
  nand ginst9723 (P2_R2027_U131, P2_R2027_U104, P2_R2027_U20);
  nand ginst9724 (P2_R2027_U132, P2_INSTADDRPOINTER_REG_7__SCAN_IN, P2_R2027_U17);
  nand ginst9725 (P2_R2027_U133, P2_R2027_U103, P2_R2027_U18);
  nand ginst9726 (P2_R2027_U134, P2_INSTADDRPOINTER_REG_6__SCAN_IN, P2_R2027_U15);
  nand ginst9727 (P2_R2027_U135, P2_R2027_U102, P2_R2027_U16);
  nand ginst9728 (P2_R2027_U136, P2_INSTADDRPOINTER_REG_5__SCAN_IN, P2_R2027_U13);
  nand ginst9729 (P2_R2027_U137, P2_R2027_U101, P2_R2027_U14);
  nand ginst9730 (P2_R2027_U138, P2_INSTADDRPOINTER_REG_4__SCAN_IN, P2_R2027_U11);
  nand ginst9731 (P2_R2027_U139, P2_R2027_U100, P2_R2027_U12);
  not ginst9732 (P2_R2027_U14, P2_INSTADDRPOINTER_REG_5__SCAN_IN);
  nand ginst9733 (P2_R2027_U140, P2_INSTADDRPOINTER_REG_3__SCAN_IN, P2_R2027_U9);
  nand ginst9734 (P2_R2027_U141, P2_R2027_U10, P2_R2027_U99);
  nand ginst9735 (P2_R2027_U142, P2_INSTADDRPOINTER_REG_31__SCAN_IN, P2_R2027_U97);
  nand ginst9736 (P2_R2027_U143, P2_R2027_U127, P2_R2027_U96);
  nand ginst9737 (P2_R2027_U144, P2_INSTADDRPOINTER_REG_30__SCAN_IN, P2_R2027_U63);
  nand ginst9738 (P2_R2027_U145, P2_R2027_U126, P2_R2027_U64);
  nand ginst9739 (P2_R2027_U146, P2_INSTADDRPOINTER_REG_2__SCAN_IN, P2_R2027_U7);
  nand ginst9740 (P2_R2027_U147, P2_R2027_U8, P2_R2027_U98);
  nand ginst9741 (P2_R2027_U148, P2_INSTADDRPOINTER_REG_29__SCAN_IN, P2_R2027_U61);
  nand ginst9742 (P2_R2027_U149, P2_R2027_U125, P2_R2027_U62);
  nand ginst9743 (P2_R2027_U15, P2_INSTADDRPOINTER_REG_5__SCAN_IN, P2_R2027_U101);
  nand ginst9744 (P2_R2027_U150, P2_INSTADDRPOINTER_REG_28__SCAN_IN, P2_R2027_U59);
  nand ginst9745 (P2_R2027_U151, P2_R2027_U124, P2_R2027_U60);
  nand ginst9746 (P2_R2027_U152, P2_INSTADDRPOINTER_REG_27__SCAN_IN, P2_R2027_U57);
  nand ginst9747 (P2_R2027_U153, P2_R2027_U123, P2_R2027_U58);
  nand ginst9748 (P2_R2027_U154, P2_INSTADDRPOINTER_REG_26__SCAN_IN, P2_R2027_U55);
  nand ginst9749 (P2_R2027_U155, P2_R2027_U122, P2_R2027_U56);
  nand ginst9750 (P2_R2027_U156, P2_INSTADDRPOINTER_REG_25__SCAN_IN, P2_R2027_U53);
  nand ginst9751 (P2_R2027_U157, P2_R2027_U121, P2_R2027_U54);
  nand ginst9752 (P2_R2027_U158, P2_INSTADDRPOINTER_REG_24__SCAN_IN, P2_R2027_U51);
  nand ginst9753 (P2_R2027_U159, P2_R2027_U120, P2_R2027_U52);
  not ginst9754 (P2_R2027_U16, P2_INSTADDRPOINTER_REG_6__SCAN_IN);
  nand ginst9755 (P2_R2027_U160, P2_INSTADDRPOINTER_REG_23__SCAN_IN, P2_R2027_U49);
  nand ginst9756 (P2_R2027_U161, P2_R2027_U119, P2_R2027_U50);
  nand ginst9757 (P2_R2027_U162, P2_INSTADDRPOINTER_REG_22__SCAN_IN, P2_R2027_U47);
  nand ginst9758 (P2_R2027_U163, P2_R2027_U118, P2_R2027_U48);
  nand ginst9759 (P2_R2027_U164, P2_INSTADDRPOINTER_REG_21__SCAN_IN, P2_R2027_U45);
  nand ginst9760 (P2_R2027_U165, P2_R2027_U117, P2_R2027_U46);
  nand ginst9761 (P2_R2027_U166, P2_INSTADDRPOINTER_REG_20__SCAN_IN, P2_R2027_U43);
  nand ginst9762 (P2_R2027_U167, P2_R2027_U116, P2_R2027_U44);
  nand ginst9763 (P2_R2027_U168, P2_INSTADDRPOINTER_REG_1__SCAN_IN, P2_R2027_U5);
  nand ginst9764 (P2_R2027_U169, P2_INSTADDRPOINTER_REG_0__SCAN_IN, P2_R2027_U6);
  nand ginst9765 (P2_R2027_U17, P2_INSTADDRPOINTER_REG_6__SCAN_IN, P2_R2027_U102);
  nand ginst9766 (P2_R2027_U170, P2_INSTADDRPOINTER_REG_19__SCAN_IN, P2_R2027_U41);
  nand ginst9767 (P2_R2027_U171, P2_R2027_U115, P2_R2027_U42);
  nand ginst9768 (P2_R2027_U172, P2_INSTADDRPOINTER_REG_18__SCAN_IN, P2_R2027_U39);
  nand ginst9769 (P2_R2027_U173, P2_R2027_U114, P2_R2027_U40);
  nand ginst9770 (P2_R2027_U174, P2_INSTADDRPOINTER_REG_17__SCAN_IN, P2_R2027_U37);
  nand ginst9771 (P2_R2027_U175, P2_R2027_U113, P2_R2027_U38);
  nand ginst9772 (P2_R2027_U176, P2_INSTADDRPOINTER_REG_16__SCAN_IN, P2_R2027_U35);
  nand ginst9773 (P2_R2027_U177, P2_R2027_U112, P2_R2027_U36);
  nand ginst9774 (P2_R2027_U178, P2_INSTADDRPOINTER_REG_15__SCAN_IN, P2_R2027_U33);
  nand ginst9775 (P2_R2027_U179, P2_R2027_U111, P2_R2027_U34);
  not ginst9776 (P2_R2027_U18, P2_INSTADDRPOINTER_REG_7__SCAN_IN);
  nand ginst9777 (P2_R2027_U180, P2_INSTADDRPOINTER_REG_14__SCAN_IN, P2_R2027_U31);
  nand ginst9778 (P2_R2027_U181, P2_R2027_U110, P2_R2027_U32);
  nand ginst9779 (P2_R2027_U182, P2_INSTADDRPOINTER_REG_13__SCAN_IN, P2_R2027_U29);
  nand ginst9780 (P2_R2027_U183, P2_R2027_U109, P2_R2027_U30);
  nand ginst9781 (P2_R2027_U184, P2_INSTADDRPOINTER_REG_12__SCAN_IN, P2_R2027_U27);
  nand ginst9782 (P2_R2027_U185, P2_R2027_U108, P2_R2027_U28);
  nand ginst9783 (P2_R2027_U186, P2_INSTADDRPOINTER_REG_11__SCAN_IN, P2_R2027_U25);
  nand ginst9784 (P2_R2027_U187, P2_R2027_U107, P2_R2027_U26);
  nand ginst9785 (P2_R2027_U188, P2_INSTADDRPOINTER_REG_10__SCAN_IN, P2_R2027_U23);
  nand ginst9786 (P2_R2027_U189, P2_R2027_U106, P2_R2027_U24);
  nand ginst9787 (P2_R2027_U19, P2_INSTADDRPOINTER_REG_7__SCAN_IN, P2_R2027_U103);
  not ginst9788 (P2_R2027_U20, P2_INSTADDRPOINTER_REG_8__SCAN_IN);
  not ginst9789 (P2_R2027_U21, P2_INSTADDRPOINTER_REG_9__SCAN_IN);
  nand ginst9790 (P2_R2027_U22, P2_INSTADDRPOINTER_REG_8__SCAN_IN, P2_R2027_U104);
  nand ginst9791 (P2_R2027_U23, P2_INSTADDRPOINTER_REG_9__SCAN_IN, P2_R2027_U105);
  not ginst9792 (P2_R2027_U24, P2_INSTADDRPOINTER_REG_10__SCAN_IN);
  nand ginst9793 (P2_R2027_U25, P2_INSTADDRPOINTER_REG_10__SCAN_IN, P2_R2027_U106);
  not ginst9794 (P2_R2027_U26, P2_INSTADDRPOINTER_REG_11__SCAN_IN);
  nand ginst9795 (P2_R2027_U27, P2_INSTADDRPOINTER_REG_11__SCAN_IN, P2_R2027_U107);
  not ginst9796 (P2_R2027_U28, P2_INSTADDRPOINTER_REG_12__SCAN_IN);
  nand ginst9797 (P2_R2027_U29, P2_INSTADDRPOINTER_REG_12__SCAN_IN, P2_R2027_U108);
  not ginst9798 (P2_R2027_U30, P2_INSTADDRPOINTER_REG_13__SCAN_IN);
  nand ginst9799 (P2_R2027_U31, P2_INSTADDRPOINTER_REG_13__SCAN_IN, P2_R2027_U109);
  not ginst9800 (P2_R2027_U32, P2_INSTADDRPOINTER_REG_14__SCAN_IN);
  nand ginst9801 (P2_R2027_U33, P2_INSTADDRPOINTER_REG_14__SCAN_IN, P2_R2027_U110);
  not ginst9802 (P2_R2027_U34, P2_INSTADDRPOINTER_REG_15__SCAN_IN);
  nand ginst9803 (P2_R2027_U35, P2_INSTADDRPOINTER_REG_15__SCAN_IN, P2_R2027_U111);
  not ginst9804 (P2_R2027_U36, P2_INSTADDRPOINTER_REG_16__SCAN_IN);
  nand ginst9805 (P2_R2027_U37, P2_INSTADDRPOINTER_REG_16__SCAN_IN, P2_R2027_U112);
  not ginst9806 (P2_R2027_U38, P2_INSTADDRPOINTER_REG_17__SCAN_IN);
  nand ginst9807 (P2_R2027_U39, P2_INSTADDRPOINTER_REG_17__SCAN_IN, P2_R2027_U113);
  not ginst9808 (P2_R2027_U40, P2_INSTADDRPOINTER_REG_18__SCAN_IN);
  nand ginst9809 (P2_R2027_U41, P2_INSTADDRPOINTER_REG_18__SCAN_IN, P2_R2027_U114);
  not ginst9810 (P2_R2027_U42, P2_INSTADDRPOINTER_REG_19__SCAN_IN);
  nand ginst9811 (P2_R2027_U43, P2_INSTADDRPOINTER_REG_19__SCAN_IN, P2_R2027_U115);
  not ginst9812 (P2_R2027_U44, P2_INSTADDRPOINTER_REG_20__SCAN_IN);
  nand ginst9813 (P2_R2027_U45, P2_INSTADDRPOINTER_REG_20__SCAN_IN, P2_R2027_U116);
  not ginst9814 (P2_R2027_U46, P2_INSTADDRPOINTER_REG_21__SCAN_IN);
  nand ginst9815 (P2_R2027_U47, P2_INSTADDRPOINTER_REG_21__SCAN_IN, P2_R2027_U117);
  not ginst9816 (P2_R2027_U48, P2_INSTADDRPOINTER_REG_22__SCAN_IN);
  nand ginst9817 (P2_R2027_U49, P2_INSTADDRPOINTER_REG_22__SCAN_IN, P2_R2027_U118);
  not ginst9818 (P2_R2027_U5, P2_INSTADDRPOINTER_REG_0__SCAN_IN);
  not ginst9819 (P2_R2027_U50, P2_INSTADDRPOINTER_REG_23__SCAN_IN);
  nand ginst9820 (P2_R2027_U51, P2_INSTADDRPOINTER_REG_23__SCAN_IN, P2_R2027_U119);
  not ginst9821 (P2_R2027_U52, P2_INSTADDRPOINTER_REG_24__SCAN_IN);
  nand ginst9822 (P2_R2027_U53, P2_INSTADDRPOINTER_REG_24__SCAN_IN, P2_R2027_U120);
  not ginst9823 (P2_R2027_U54, P2_INSTADDRPOINTER_REG_25__SCAN_IN);
  nand ginst9824 (P2_R2027_U55, P2_INSTADDRPOINTER_REG_25__SCAN_IN, P2_R2027_U121);
  not ginst9825 (P2_R2027_U56, P2_INSTADDRPOINTER_REG_26__SCAN_IN);
  nand ginst9826 (P2_R2027_U57, P2_INSTADDRPOINTER_REG_26__SCAN_IN, P2_R2027_U122);
  not ginst9827 (P2_R2027_U58, P2_INSTADDRPOINTER_REG_27__SCAN_IN);
  nand ginst9828 (P2_R2027_U59, P2_INSTADDRPOINTER_REG_27__SCAN_IN, P2_R2027_U123);
  not ginst9829 (P2_R2027_U6, P2_INSTADDRPOINTER_REG_1__SCAN_IN);
  not ginst9830 (P2_R2027_U60, P2_INSTADDRPOINTER_REG_28__SCAN_IN);
  nand ginst9831 (P2_R2027_U61, P2_INSTADDRPOINTER_REG_28__SCAN_IN, P2_R2027_U124);
  not ginst9832 (P2_R2027_U62, P2_INSTADDRPOINTER_REG_29__SCAN_IN);
  nand ginst9833 (P2_R2027_U63, P2_INSTADDRPOINTER_REG_29__SCAN_IN, P2_R2027_U125);
  not ginst9834 (P2_R2027_U64, P2_INSTADDRPOINTER_REG_30__SCAN_IN);
  nand ginst9835 (P2_R2027_U65, P2_R2027_U128, P2_R2027_U129);
  nand ginst9836 (P2_R2027_U66, P2_R2027_U130, P2_R2027_U131);
  nand ginst9837 (P2_R2027_U67, P2_R2027_U132, P2_R2027_U133);
  nand ginst9838 (P2_R2027_U68, P2_R2027_U134, P2_R2027_U135);
  nand ginst9839 (P2_R2027_U69, P2_R2027_U136, P2_R2027_U137);
  nand ginst9840 (P2_R2027_U7, P2_INSTADDRPOINTER_REG_0__SCAN_IN, P2_INSTADDRPOINTER_REG_1__SCAN_IN);
  nand ginst9841 (P2_R2027_U70, P2_R2027_U138, P2_R2027_U139);
  nand ginst9842 (P2_R2027_U71, P2_R2027_U140, P2_R2027_U141);
  nand ginst9843 (P2_R2027_U72, P2_R2027_U142, P2_R2027_U143);
  nand ginst9844 (P2_R2027_U73, P2_R2027_U144, P2_R2027_U145);
  nand ginst9845 (P2_R2027_U74, P2_R2027_U146, P2_R2027_U147);
  nand ginst9846 (P2_R2027_U75, P2_R2027_U148, P2_R2027_U149);
  nand ginst9847 (P2_R2027_U76, P2_R2027_U150, P2_R2027_U151);
  nand ginst9848 (P2_R2027_U77, P2_R2027_U152, P2_R2027_U153);
  nand ginst9849 (P2_R2027_U78, P2_R2027_U154, P2_R2027_U155);
  nand ginst9850 (P2_R2027_U79, P2_R2027_U156, P2_R2027_U157);
  not ginst9851 (P2_R2027_U8, P2_INSTADDRPOINTER_REG_2__SCAN_IN);
  nand ginst9852 (P2_R2027_U80, P2_R2027_U158, P2_R2027_U159);
  nand ginst9853 (P2_R2027_U81, P2_R2027_U160, P2_R2027_U161);
  nand ginst9854 (P2_R2027_U82, P2_R2027_U162, P2_R2027_U163);
  nand ginst9855 (P2_R2027_U83, P2_R2027_U164, P2_R2027_U165);
  nand ginst9856 (P2_R2027_U84, P2_R2027_U166, P2_R2027_U167);
  nand ginst9857 (P2_R2027_U85, P2_R2027_U168, P2_R2027_U169);
  nand ginst9858 (P2_R2027_U86, P2_R2027_U170, P2_R2027_U171);
  nand ginst9859 (P2_R2027_U87, P2_R2027_U172, P2_R2027_U173);
  nand ginst9860 (P2_R2027_U88, P2_R2027_U174, P2_R2027_U175);
  nand ginst9861 (P2_R2027_U89, P2_R2027_U176, P2_R2027_U177);
  nand ginst9862 (P2_R2027_U9, P2_INSTADDRPOINTER_REG_2__SCAN_IN, P2_R2027_U98);
  nand ginst9863 (P2_R2027_U90, P2_R2027_U178, P2_R2027_U179);
  nand ginst9864 (P2_R2027_U91, P2_R2027_U180, P2_R2027_U181);
  nand ginst9865 (P2_R2027_U92, P2_R2027_U182, P2_R2027_U183);
  nand ginst9866 (P2_R2027_U93, P2_R2027_U184, P2_R2027_U185);
  nand ginst9867 (P2_R2027_U94, P2_R2027_U186, P2_R2027_U187);
  nand ginst9868 (P2_R2027_U95, P2_R2027_U188, P2_R2027_U189);
  not ginst9869 (P2_R2027_U96, P2_INSTADDRPOINTER_REG_31__SCAN_IN);
  nand ginst9870 (P2_R2027_U97, P2_INSTADDRPOINTER_REG_30__SCAN_IN, P2_R2027_U126);
  not ginst9871 (P2_R2027_U98, P2_R2027_U7);
  not ginst9872 (P2_R2027_U99, P2_R2027_U9);
  nor ginst9873 (P2_R2088_U6, P2_R2088_U7, P2_U3648);
  nor ginst9874 (P2_R2088_U7, P2_U3648, P2_U3649, P2_U3650, P2_U3651, P2_U3652);
  and ginst9875 (P2_R2096_U10, P2_R2096_U9, P2_U2626);
  and ginst9876 (P2_R2096_U100, P2_R2096_U175, P2_R2096_U176);
  nand ginst9877 (P2_R2096_U101, P2_R2096_U137, P2_R2096_U138);
  and ginst9878 (P2_R2096_U102, P2_R2096_U182, P2_R2096_U183);
  nand ginst9879 (P2_R2096_U103, P2_R2096_U133, P2_R2096_U134);
  and ginst9880 (P2_R2096_U104, P2_R2096_U189, P2_R2096_U190);
  nand ginst9881 (P2_R2096_U105, P2_R2096_U129, P2_R2096_U130);
  and ginst9882 (P2_R2096_U106, P2_R2096_U196, P2_R2096_U197);
  nand ginst9883 (P2_R2096_U107, P2_R2096_U125, P2_R2096_U126);
  and ginst9884 (P2_R2096_U108, P2_R2096_U203, P2_R2096_U204);
  nand ginst9885 (P2_R2096_U109, P2_R2096_U121, P2_R2096_U122);
  and ginst9886 (P2_R2096_U11, P2_R2096_U10, P2_U2625);
  and ginst9887 (P2_R2096_U110, P2_R2096_U212, P2_R2096_U213);
  nand ginst9888 (P2_R2096_U111, P2_R2096_U113, P2_R2096_U118);
  nand ginst9889 (P2_R2096_U112, P2_U2649, P2_U2657);
  nand ginst9890 (P2_R2096_U113, P2_U2649, P2_U2656, P2_U2657);
  and ginst9891 (P2_R2096_U114, P2_R2096_U242, P2_R2096_U243);
  not ginst9892 (P2_R2096_U115, P2_R2096_U113);
  nand ginst9893 (P2_R2096_U116, P2_U2649, P2_U2657);
  nand ginst9894 (P2_R2096_U117, P2_R2096_U116, P2_R2096_U55);
  nand ginst9895 (P2_R2096_U118, P2_R2096_U117, P2_U2648);
  not ginst9896 (P2_R2096_U119, P2_R2096_U111);
  and ginst9897 (P2_R2096_U12, P2_R2096_U11, P2_U2624);
  or ginst9898 (P2_R2096_U120, P2_U2647, P2_U2655);
  nand ginst9899 (P2_R2096_U121, P2_R2096_U111, P2_R2096_U120);
  nand ginst9900 (P2_R2096_U122, P2_U2647, P2_U2655);
  not ginst9901 (P2_R2096_U123, P2_R2096_U109);
  or ginst9902 (P2_R2096_U124, P2_U2646, P2_U2654);
  nand ginst9903 (P2_R2096_U125, P2_R2096_U109, P2_R2096_U124);
  nand ginst9904 (P2_R2096_U126, P2_U2646, P2_U2654);
  not ginst9905 (P2_R2096_U127, P2_R2096_U107);
  or ginst9906 (P2_R2096_U128, P2_U2645, P2_U2653);
  nand ginst9907 (P2_R2096_U129, P2_R2096_U107, P2_R2096_U128);
  and ginst9908 (P2_R2096_U13, P2_R2096_U15, P2_U2622);
  nand ginst9909 (P2_R2096_U130, P2_U2645, P2_U2653);
  not ginst9910 (P2_R2096_U131, P2_R2096_U105);
  or ginst9911 (P2_R2096_U132, P2_U2644, P2_U2652);
  nand ginst9912 (P2_R2096_U133, P2_R2096_U105, P2_R2096_U132);
  nand ginst9913 (P2_R2096_U134, P2_U2644, P2_U2652);
  not ginst9914 (P2_R2096_U135, P2_R2096_U103);
  or ginst9915 (P2_R2096_U136, P2_U2643, P2_U2651);
  nand ginst9916 (P2_R2096_U137, P2_R2096_U103, P2_R2096_U136);
  nand ginst9917 (P2_R2096_U138, P2_U2643, P2_U2651);
  not ginst9918 (P2_R2096_U139, P2_R2096_U101);
  and ginst9919 (P2_R2096_U14, P2_R2096_U13, P2_U2621);
  or ginst9920 (P2_R2096_U140, P2_U2642, P2_U2650);
  nand ginst9921 (P2_R2096_U141, P2_R2096_U101, P2_R2096_U140);
  nand ginst9922 (P2_R2096_U142, P2_U2642, P2_U2650);
  not ginst9923 (P2_R2096_U143, P2_R2096_U99);
  not ginst9924 (P2_R2096_U144, P2_R2096_U23);
  not ginst9925 (P2_R2096_U145, P2_R2096_U4);
  not ginst9926 (P2_R2096_U146, P2_R2096_U24);
  not ginst9927 (P2_R2096_U147, P2_R2096_U19);
  not ginst9928 (P2_R2096_U148, P2_R2096_U20);
  not ginst9929 (P2_R2096_U149, P2_R2096_U21);
  and ginst9930 (P2_R2096_U15, P2_R2096_U12, P2_U2623);
  not ginst9931 (P2_R2096_U150, P2_R2096_U17);
  not ginst9932 (P2_R2096_U151, P2_R2096_U18);
  not ginst9933 (P2_R2096_U152, P2_R2096_U5);
  not ginst9934 (P2_R2096_U153, P2_R2096_U25);
  not ginst9935 (P2_R2096_U154, P2_R2096_U6);
  not ginst9936 (P2_R2096_U155, P2_R2096_U16);
  not ginst9937 (P2_R2096_U156, P2_R2096_U7);
  not ginst9938 (P2_R2096_U157, P2_R2096_U8);
  not ginst9939 (P2_R2096_U158, P2_R2096_U9);
  not ginst9940 (P2_R2096_U159, P2_R2096_U10);
  and ginst9941 (P2_R2096_U16, P2_R2096_U6, P2_U2630);
  not ginst9942 (P2_R2096_U160, P2_R2096_U11);
  not ginst9943 (P2_R2096_U161, P2_R2096_U12);
  not ginst9944 (P2_R2096_U162, P2_R2096_U15);
  not ginst9945 (P2_R2096_U163, P2_R2096_U13);
  not ginst9946 (P2_R2096_U164, P2_R2096_U14);
  not ginst9947 (P2_R2096_U165, P2_R2096_U22);
  nand ginst9948 (P2_R2096_U166, P2_R2096_U22, P2_U2619);
  nand ginst9949 (P2_R2096_U167, P2_R2096_U166, P2_R2096_U29);
  nand ginst9950 (P2_R2096_U168, P2_R2096_U22, P2_R2096_U98);
  not ginst9951 (P2_R2096_U169, P2_R2096_U112);
  and ginst9952 (P2_R2096_U17, P2_R2096_U21, P2_U2635);
  nand ginst9953 (P2_R2096_U170, P2_R2096_U241, P2_R2096_U55);
  nand ginst9954 (P2_R2096_U171, P2_R2096_U23, P2_R2096_U28);
  nand ginst9955 (P2_R2096_U172, P2_R2096_U144, P2_U2640);
  nand ginst9956 (P2_R2096_U173, P2_R2096_U37, P2_R2096_U99);
  nand ginst9957 (P2_R2096_U174, P2_R2096_U143, P2_U2641);
  nand ginst9958 (P2_R2096_U175, P2_R2096_U66, P2_U2642);
  nand ginst9959 (P2_R2096_U176, P2_R2096_U67, P2_U2650);
  nand ginst9960 (P2_R2096_U177, P2_R2096_U66, P2_U2642);
  nand ginst9961 (P2_R2096_U178, P2_R2096_U67, P2_U2650);
  nand ginst9962 (P2_R2096_U179, P2_R2096_U177, P2_R2096_U178);
  and ginst9963 (P2_R2096_U18, P2_R2096_U17, P2_U2634);
  nand ginst9964 (P2_R2096_U180, P2_R2096_U100, P2_R2096_U101);
  nand ginst9965 (P2_R2096_U181, P2_R2096_U139, P2_R2096_U179);
  nand ginst9966 (P2_R2096_U182, P2_R2096_U64, P2_U2643);
  nand ginst9967 (P2_R2096_U183, P2_R2096_U65, P2_U2651);
  nand ginst9968 (P2_R2096_U184, P2_R2096_U64, P2_U2643);
  nand ginst9969 (P2_R2096_U185, P2_R2096_U65, P2_U2651);
  nand ginst9970 (P2_R2096_U186, P2_R2096_U184, P2_R2096_U185);
  nand ginst9971 (P2_R2096_U187, P2_R2096_U102, P2_R2096_U103);
  nand ginst9972 (P2_R2096_U188, P2_R2096_U135, P2_R2096_U186);
  nand ginst9973 (P2_R2096_U189, P2_R2096_U62, P2_U2644);
  and ginst9974 (P2_R2096_U19, P2_R2096_U24, P2_U2638);
  nand ginst9975 (P2_R2096_U190, P2_R2096_U63, P2_U2652);
  nand ginst9976 (P2_R2096_U191, P2_R2096_U62, P2_U2644);
  nand ginst9977 (P2_R2096_U192, P2_R2096_U63, P2_U2652);
  nand ginst9978 (P2_R2096_U193, P2_R2096_U191, P2_R2096_U192);
  nand ginst9979 (P2_R2096_U194, P2_R2096_U104, P2_R2096_U105);
  nand ginst9980 (P2_R2096_U195, P2_R2096_U131, P2_R2096_U193);
  nand ginst9981 (P2_R2096_U196, P2_R2096_U60, P2_U2645);
  nand ginst9982 (P2_R2096_U197, P2_R2096_U61, P2_U2653);
  nand ginst9983 (P2_R2096_U198, P2_R2096_U60, P2_U2645);
  nand ginst9984 (P2_R2096_U199, P2_R2096_U61, P2_U2653);
  and ginst9985 (P2_R2096_U20, P2_R2096_U19, P2_U2637);
  nand ginst9986 (P2_R2096_U200, P2_R2096_U198, P2_R2096_U199);
  nand ginst9987 (P2_R2096_U201, P2_R2096_U106, P2_R2096_U107);
  nand ginst9988 (P2_R2096_U202, P2_R2096_U127, P2_R2096_U200);
  nand ginst9989 (P2_R2096_U203, P2_R2096_U58, P2_U2646);
  nand ginst9990 (P2_R2096_U204, P2_R2096_U59, P2_U2654);
  nand ginst9991 (P2_R2096_U205, P2_R2096_U58, P2_U2646);
  nand ginst9992 (P2_R2096_U206, P2_R2096_U59, P2_U2654);
  nand ginst9993 (P2_R2096_U207, P2_R2096_U205, P2_R2096_U206);
  nand ginst9994 (P2_R2096_U208, P2_R2096_U108, P2_R2096_U109);
  nand ginst9995 (P2_R2096_U209, P2_R2096_U123, P2_R2096_U207);
  and ginst9996 (P2_R2096_U21, P2_R2096_U20, P2_U2636);
  nand ginst9997 (P2_R2096_U210, P2_R2096_U22, P2_R2096_U30);
  nand ginst9998 (P2_R2096_U211, P2_R2096_U165, P2_U2619);
  nand ginst9999 (P2_R2096_U212, P2_R2096_U56, P2_U2647);
  nand ginst10000 (P2_R2096_U213, P2_R2096_U57, P2_U2655);
  nand ginst10001 (P2_R2096_U214, P2_R2096_U56, P2_U2647);
  nand ginst10002 (P2_R2096_U215, P2_R2096_U57, P2_U2655);
  nand ginst10003 (P2_R2096_U216, P2_R2096_U214, P2_R2096_U215);
  nand ginst10004 (P2_R2096_U217, P2_R2096_U110, P2_R2096_U111);
  nand ginst10005 (P2_R2096_U218, P2_R2096_U119, P2_R2096_U216);
  nand ginst10006 (P2_R2096_U219, P2_R2096_U14, P2_R2096_U40);
  and ginst10007 (P2_R2096_U22, P2_R2096_U14, P2_U2620);
  nand ginst10008 (P2_R2096_U220, P2_R2096_U164, P2_U2620);
  nand ginst10009 (P2_R2096_U221, P2_R2096_U13, P2_R2096_U41);
  nand ginst10010 (P2_R2096_U222, P2_R2096_U163, P2_U2621);
  nand ginst10011 (P2_R2096_U223, P2_R2096_U15, P2_R2096_U38);
  nand ginst10012 (P2_R2096_U224, P2_R2096_U162, P2_U2622);
  nand ginst10013 (P2_R2096_U225, P2_R2096_U12, P2_R2096_U42);
  nand ginst10014 (P2_R2096_U226, P2_R2096_U161, P2_U2623);
  nand ginst10015 (P2_R2096_U227, P2_R2096_U11, P2_R2096_U43);
  nand ginst10016 (P2_R2096_U228, P2_R2096_U160, P2_U2624);
  nand ginst10017 (P2_R2096_U229, P2_R2096_U10, P2_R2096_U44);
  and ginst10018 (P2_R2096_U23, P2_R2096_U99, P2_U2641);
  nand ginst10019 (P2_R2096_U230, P2_R2096_U159, P2_U2625);
  nand ginst10020 (P2_R2096_U231, P2_R2096_U45, P2_R2096_U9);
  nand ginst10021 (P2_R2096_U232, P2_R2096_U158, P2_U2626);
  nand ginst10022 (P2_R2096_U233, P2_R2096_U39, P2_R2096_U8);
  nand ginst10023 (P2_R2096_U234, P2_R2096_U157, P2_U2627);
  nand ginst10024 (P2_R2096_U235, P2_R2096_U46, P2_R2096_U7);
  nand ginst10025 (P2_R2096_U236, P2_R2096_U156, P2_U2628);
  nand ginst10026 (P2_R2096_U237, P2_R2096_U16, P2_R2096_U36);
  nand ginst10027 (P2_R2096_U238, P2_R2096_U155, P2_U2629);
  nand ginst10028 (P2_R2096_U239, P2_R2096_U112, P2_U2648);
  and ginst10029 (P2_R2096_U24, P2_R2096_U4, P2_U2639);
  nand ginst10030 (P2_R2096_U240, P2_R2096_U169, P2_R2096_U54);
  nand ginst10031 (P2_R2096_U241, P2_R2096_U239, P2_R2096_U240);
  nand ginst10032 (P2_R2096_U242, P2_R2096_U116, P2_R2096_U54, P2_U2656);
  nand ginst10033 (P2_R2096_U243, P2_R2096_U115, P2_U2648);
  nand ginst10034 (P2_R2096_U244, P2_R2096_U47, P2_R2096_U6);
  nand ginst10035 (P2_R2096_U245, P2_R2096_U154, P2_U2630);
  nand ginst10036 (P2_R2096_U246, P2_R2096_U25, P2_R2096_U26);
  nand ginst10037 (P2_R2096_U247, P2_R2096_U153, P2_U2631);
  nand ginst10038 (P2_R2096_U248, P2_R2096_U48, P2_R2096_U5);
  nand ginst10039 (P2_R2096_U249, P2_R2096_U152, P2_U2632);
  and ginst10040 (P2_R2096_U25, P2_R2096_U5, P2_U2632);
  nand ginst10041 (P2_R2096_U250, P2_R2096_U18, P2_R2096_U34);
  nand ginst10042 (P2_R2096_U251, P2_R2096_U151, P2_U2633);
  nand ginst10043 (P2_R2096_U252, P2_R2096_U17, P2_R2096_U35);
  nand ginst10044 (P2_R2096_U253, P2_R2096_U150, P2_U2634);
  nand ginst10045 (P2_R2096_U254, P2_R2096_U21, P2_R2096_U31);
  nand ginst10046 (P2_R2096_U255, P2_R2096_U149, P2_U2635);
  nand ginst10047 (P2_R2096_U256, P2_R2096_U20, P2_R2096_U32);
  nand ginst10048 (P2_R2096_U257, P2_R2096_U148, P2_U2636);
  nand ginst10049 (P2_R2096_U258, P2_R2096_U19, P2_R2096_U33);
  nand ginst10050 (P2_R2096_U259, P2_R2096_U147, P2_U2637);
  not ginst10051 (P2_R2096_U26, P2_U2631);
  nand ginst10052 (P2_R2096_U260, P2_R2096_U24, P2_R2096_U27);
  nand ginst10053 (P2_R2096_U261, P2_R2096_U146, P2_U2638);
  nand ginst10054 (P2_R2096_U262, P2_R2096_U4, P2_R2096_U49);
  nand ginst10055 (P2_R2096_U263, P2_R2096_U145, P2_U2639);
  nand ginst10056 (P2_R2096_U264, P2_R2096_U52, P2_U2649);
  nand ginst10057 (P2_R2096_U265, P2_R2096_U53, P2_U2657);
  not ginst10058 (P2_R2096_U27, P2_U2638);
  not ginst10059 (P2_R2096_U28, P2_U2640);
  not ginst10060 (P2_R2096_U29, P2_U2618);
  not ginst10061 (P2_R2096_U30, P2_U2619);
  not ginst10062 (P2_R2096_U31, P2_U2635);
  not ginst10063 (P2_R2096_U32, P2_U2636);
  not ginst10064 (P2_R2096_U33, P2_U2637);
  not ginst10065 (P2_R2096_U34, P2_U2633);
  not ginst10066 (P2_R2096_U35, P2_U2634);
  not ginst10067 (P2_R2096_U36, P2_U2629);
  not ginst10068 (P2_R2096_U37, P2_U2641);
  not ginst10069 (P2_R2096_U38, P2_U2622);
  not ginst10070 (P2_R2096_U39, P2_U2627);
  and ginst10071 (P2_R2096_U4, P2_R2096_U23, P2_U2640);
  not ginst10072 (P2_R2096_U40, P2_U2620);
  not ginst10073 (P2_R2096_U41, P2_U2621);
  not ginst10074 (P2_R2096_U42, P2_U2623);
  not ginst10075 (P2_R2096_U43, P2_U2624);
  not ginst10076 (P2_R2096_U44, P2_U2625);
  not ginst10077 (P2_R2096_U45, P2_U2626);
  not ginst10078 (P2_R2096_U46, P2_U2628);
  not ginst10079 (P2_R2096_U47, P2_U2630);
  not ginst10080 (P2_R2096_U48, P2_U2632);
  not ginst10081 (P2_R2096_U49, P2_U2639);
  and ginst10082 (P2_R2096_U5, P2_R2096_U18, P2_U2633);
  and ginst10083 (P2_R2096_U50, P2_R2096_U167, P2_R2096_U168);
  nand ginst10084 (P2_R2096_U51, P2_R2096_U114, P2_R2096_U170);
  not ginst10085 (P2_R2096_U52, P2_U2657);
  not ginst10086 (P2_R2096_U53, P2_U2649);
  not ginst10087 (P2_R2096_U54, P2_U2648);
  not ginst10088 (P2_R2096_U55, P2_U2656);
  not ginst10089 (P2_R2096_U56, P2_U2655);
  not ginst10090 (P2_R2096_U57, P2_U2647);
  not ginst10091 (P2_R2096_U58, P2_U2654);
  not ginst10092 (P2_R2096_U59, P2_U2646);
  and ginst10093 (P2_R2096_U6, P2_R2096_U25, P2_U2631);
  not ginst10094 (P2_R2096_U60, P2_U2653);
  not ginst10095 (P2_R2096_U61, P2_U2645);
  not ginst10096 (P2_R2096_U62, P2_U2652);
  not ginst10097 (P2_R2096_U63, P2_U2644);
  not ginst10098 (P2_R2096_U64, P2_U2651);
  not ginst10099 (P2_R2096_U65, P2_U2643);
  not ginst10100 (P2_R2096_U66, P2_U2650);
  not ginst10101 (P2_R2096_U67, P2_U2642);
  nand ginst10102 (P2_R2096_U68, P2_R2096_U264, P2_R2096_U265);
  nand ginst10103 (P2_R2096_U69, P2_R2096_U171, P2_R2096_U172);
  and ginst10104 (P2_R2096_U7, P2_R2096_U16, P2_U2629);
  nand ginst10105 (P2_R2096_U70, P2_R2096_U173, P2_R2096_U174);
  nand ginst10106 (P2_R2096_U71, P2_R2096_U180, P2_R2096_U181);
  nand ginst10107 (P2_R2096_U72, P2_R2096_U187, P2_R2096_U188);
  nand ginst10108 (P2_R2096_U73, P2_R2096_U194, P2_R2096_U195);
  nand ginst10109 (P2_R2096_U74, P2_R2096_U201, P2_R2096_U202);
  nand ginst10110 (P2_R2096_U75, P2_R2096_U208, P2_R2096_U209);
  nand ginst10111 (P2_R2096_U76, P2_R2096_U210, P2_R2096_U211);
  nand ginst10112 (P2_R2096_U77, P2_R2096_U217, P2_R2096_U218);
  nand ginst10113 (P2_R2096_U78, P2_R2096_U219, P2_R2096_U220);
  nand ginst10114 (P2_R2096_U79, P2_R2096_U221, P2_R2096_U222);
  and ginst10115 (P2_R2096_U8, P2_R2096_U7, P2_U2628);
  nand ginst10116 (P2_R2096_U80, P2_R2096_U223, P2_R2096_U224);
  nand ginst10117 (P2_R2096_U81, P2_R2096_U225, P2_R2096_U226);
  nand ginst10118 (P2_R2096_U82, P2_R2096_U227, P2_R2096_U228);
  nand ginst10119 (P2_R2096_U83, P2_R2096_U229, P2_R2096_U230);
  nand ginst10120 (P2_R2096_U84, P2_R2096_U231, P2_R2096_U232);
  nand ginst10121 (P2_R2096_U85, P2_R2096_U233, P2_R2096_U234);
  nand ginst10122 (P2_R2096_U86, P2_R2096_U235, P2_R2096_U236);
  nand ginst10123 (P2_R2096_U87, P2_R2096_U237, P2_R2096_U238);
  nand ginst10124 (P2_R2096_U88, P2_R2096_U244, P2_R2096_U245);
  nand ginst10125 (P2_R2096_U89, P2_R2096_U246, P2_R2096_U247);
  and ginst10126 (P2_R2096_U9, P2_R2096_U8, P2_U2627);
  nand ginst10127 (P2_R2096_U90, P2_R2096_U248, P2_R2096_U249);
  nand ginst10128 (P2_R2096_U91, P2_R2096_U250, P2_R2096_U251);
  nand ginst10129 (P2_R2096_U92, P2_R2096_U252, P2_R2096_U253);
  nand ginst10130 (P2_R2096_U93, P2_R2096_U254, P2_R2096_U255);
  nand ginst10131 (P2_R2096_U94, P2_R2096_U256, P2_R2096_U257);
  nand ginst10132 (P2_R2096_U95, P2_R2096_U258, P2_R2096_U259);
  nand ginst10133 (P2_R2096_U96, P2_R2096_U260, P2_R2096_U261);
  nand ginst10134 (P2_R2096_U97, P2_R2096_U262, P2_R2096_U263);
  and ginst10135 (P2_R2096_U98, P2_U2618, P2_U2619);
  nand ginst10136 (P2_R2096_U99, P2_R2096_U141, P2_R2096_U142);
  not ginst10137 (P2_R2099_U10, P2_U2749);
  nand ginst10138 (P2_R2099_U100, P2_R2099_U113, P2_R2099_U114);
  not ginst10139 (P2_R2099_U101, P2_U2716);
  nand ginst10140 (P2_R2099_U102, P2_R2099_U145, P2_U2717);
  and ginst10141 (P2_R2099_U103, P2_R2099_U172, P2_R2099_U173);
  nand ginst10142 (P2_R2099_U104, P2_R2099_U106, P2_R2099_U110);
  nand ginst10143 (P2_R2099_U105, P2_U2747, P2_U2751);
  nand ginst10144 (P2_R2099_U106, P2_U2746, P2_U2747, P2_U2751);
  and ginst10145 (P2_R2099_U107, P2_R2099_U202, P2_R2099_U203);
  not ginst10146 (P2_R2099_U108, P2_R2099_U106);
  nand ginst10147 (P2_R2099_U109, P2_R2099_U105, P2_R2099_U9);
  not ginst10148 (P2_R2099_U11, P2_U2745);
  nand ginst10149 (P2_R2099_U110, P2_R2099_U109, P2_U2750);
  not ginst10150 (P2_R2099_U111, P2_R2099_U104);
  or ginst10151 (P2_R2099_U112, P2_U2745, P2_U2749);
  nand ginst10152 (P2_R2099_U113, P2_R2099_U104, P2_R2099_U112);
  nand ginst10153 (P2_R2099_U114, P2_U2745, P2_U2749);
  not ginst10154 (P2_R2099_U115, P2_R2099_U100);
  or ginst10155 (P2_R2099_U116, P2_U2744, P2_U2748);
  nand ginst10156 (P2_R2099_U117, P2_R2099_U100, P2_R2099_U116);
  nand ginst10157 (P2_R2099_U118, P2_U2744, P2_U2748);
  not ginst10158 (P2_R2099_U119, P2_R2099_U97);
  not ginst10159 (P2_R2099_U12, P2_U2748);
  not ginst10160 (P2_R2099_U120, P2_R2099_U15);
  not ginst10161 (P2_R2099_U121, P2_R2099_U17);
  not ginst10162 (P2_R2099_U122, P2_R2099_U19);
  not ginst10163 (P2_R2099_U123, P2_R2099_U21);
  not ginst10164 (P2_R2099_U124, P2_R2099_U24);
  not ginst10165 (P2_R2099_U125, P2_R2099_U25);
  not ginst10166 (P2_R2099_U126, P2_R2099_U27);
  not ginst10167 (P2_R2099_U127, P2_R2099_U29);
  not ginst10168 (P2_R2099_U128, P2_R2099_U31);
  not ginst10169 (P2_R2099_U129, P2_R2099_U33);
  not ginst10170 (P2_R2099_U13, P2_U2744);
  not ginst10171 (P2_R2099_U130, P2_R2099_U35);
  not ginst10172 (P2_R2099_U131, P2_R2099_U37);
  not ginst10173 (P2_R2099_U132, P2_R2099_U39);
  not ginst10174 (P2_R2099_U133, P2_R2099_U41);
  not ginst10175 (P2_R2099_U134, P2_R2099_U43);
  not ginst10176 (P2_R2099_U135, P2_R2099_U45);
  not ginst10177 (P2_R2099_U136, P2_R2099_U47);
  not ginst10178 (P2_R2099_U137, P2_R2099_U49);
  not ginst10179 (P2_R2099_U138, P2_R2099_U51);
  not ginst10180 (P2_R2099_U139, P2_R2099_U53);
  not ginst10181 (P2_R2099_U14, P2_U2743);
  not ginst10182 (P2_R2099_U140, P2_R2099_U55);
  not ginst10183 (P2_R2099_U141, P2_R2099_U57);
  not ginst10184 (P2_R2099_U142, P2_R2099_U59);
  not ginst10185 (P2_R2099_U143, P2_R2099_U61);
  not ginst10186 (P2_R2099_U144, P2_R2099_U63);
  not ginst10187 (P2_R2099_U145, P2_R2099_U65);
  not ginst10188 (P2_R2099_U146, P2_R2099_U102);
  not ginst10189 (P2_R2099_U147, P2_R2099_U105);
  nand ginst10190 (P2_R2099_U148, P2_R2099_U201, P2_R2099_U9);
  nand ginst10191 (P2_R2099_U149, P2_R2099_U24, P2_U2738);
  nand ginst10192 (P2_R2099_U15, P2_R2099_U97, P2_U2743);
  nand ginst10193 (P2_R2099_U150, P2_R2099_U124, P2_R2099_U23);
  nand ginst10194 (P2_R2099_U151, P2_R2099_U21, P2_U2739);
  nand ginst10195 (P2_R2099_U152, P2_R2099_U123, P2_R2099_U22);
  nand ginst10196 (P2_R2099_U153, P2_R2099_U19, P2_U2740);
  nand ginst10197 (P2_R2099_U154, P2_R2099_U122, P2_R2099_U20);
  nand ginst10198 (P2_R2099_U155, P2_R2099_U17, P2_U2741);
  nand ginst10199 (P2_R2099_U156, P2_R2099_U121, P2_R2099_U18);
  nand ginst10200 (P2_R2099_U157, P2_R2099_U15, P2_U2742);
  nand ginst10201 (P2_R2099_U158, P2_R2099_U120, P2_R2099_U16);
  nand ginst10202 (P2_R2099_U159, P2_R2099_U97, P2_U2743);
  not ginst10203 (P2_R2099_U16, P2_U2742);
  nand ginst10204 (P2_R2099_U160, P2_R2099_U119, P2_R2099_U14);
  nand ginst10205 (P2_R2099_U161, P2_R2099_U12, P2_U2744);
  nand ginst10206 (P2_R2099_U162, P2_R2099_U13, P2_U2748);
  nand ginst10207 (P2_R2099_U163, P2_R2099_U12, P2_U2744);
  nand ginst10208 (P2_R2099_U164, P2_R2099_U13, P2_U2748);
  nand ginst10209 (P2_R2099_U165, P2_R2099_U163, P2_R2099_U164);
  nand ginst10210 (P2_R2099_U166, P2_R2099_U100, P2_R2099_U99);
  nand ginst10211 (P2_R2099_U167, P2_R2099_U115, P2_R2099_U165);
  nand ginst10212 (P2_R2099_U168, P2_R2099_U102, P2_U2716);
  nand ginst10213 (P2_R2099_U169, P2_R2099_U101, P2_R2099_U146);
  nand ginst10214 (P2_R2099_U17, P2_R2099_U120, P2_U2742);
  nand ginst10215 (P2_R2099_U170, P2_R2099_U65, P2_U2717);
  nand ginst10216 (P2_R2099_U171, P2_R2099_U145, P2_R2099_U66);
  nand ginst10217 (P2_R2099_U172, P2_R2099_U10, P2_U2745);
  nand ginst10218 (P2_R2099_U173, P2_R2099_U11, P2_U2749);
  nand ginst10219 (P2_R2099_U174, P2_R2099_U10, P2_U2745);
  nand ginst10220 (P2_R2099_U175, P2_R2099_U11, P2_U2749);
  nand ginst10221 (P2_R2099_U176, P2_R2099_U174, P2_R2099_U175);
  nand ginst10222 (P2_R2099_U177, P2_R2099_U103, P2_R2099_U104);
  nand ginst10223 (P2_R2099_U178, P2_R2099_U111, P2_R2099_U176);
  nand ginst10224 (P2_R2099_U179, P2_R2099_U63, P2_U2718);
  not ginst10225 (P2_R2099_U18, P2_U2741);
  nand ginst10226 (P2_R2099_U180, P2_R2099_U144, P2_R2099_U64);
  nand ginst10227 (P2_R2099_U181, P2_R2099_U61, P2_U2719);
  nand ginst10228 (P2_R2099_U182, P2_R2099_U143, P2_R2099_U62);
  nand ginst10229 (P2_R2099_U183, P2_R2099_U59, P2_U2720);
  nand ginst10230 (P2_R2099_U184, P2_R2099_U142, P2_R2099_U60);
  nand ginst10231 (P2_R2099_U185, P2_R2099_U57, P2_U2721);
  nand ginst10232 (P2_R2099_U186, P2_R2099_U141, P2_R2099_U58);
  nand ginst10233 (P2_R2099_U187, P2_R2099_U55, P2_U2722);
  nand ginst10234 (P2_R2099_U188, P2_R2099_U140, P2_R2099_U56);
  nand ginst10235 (P2_R2099_U189, P2_R2099_U53, P2_U2723);
  nand ginst10236 (P2_R2099_U19, P2_R2099_U121, P2_U2741);
  nand ginst10237 (P2_R2099_U190, P2_R2099_U139, P2_R2099_U54);
  nand ginst10238 (P2_R2099_U191, P2_R2099_U51, P2_U2724);
  nand ginst10239 (P2_R2099_U192, P2_R2099_U138, P2_R2099_U52);
  nand ginst10240 (P2_R2099_U193, P2_R2099_U49, P2_U2725);
  nand ginst10241 (P2_R2099_U194, P2_R2099_U137, P2_R2099_U50);
  nand ginst10242 (P2_R2099_U195, P2_R2099_U47, P2_U2726);
  nand ginst10243 (P2_R2099_U196, P2_R2099_U136, P2_R2099_U48);
  nand ginst10244 (P2_R2099_U197, P2_R2099_U45, P2_U2727);
  nand ginst10245 (P2_R2099_U198, P2_R2099_U135, P2_R2099_U46);
  nand ginst10246 (P2_R2099_U199, P2_R2099_U105, P2_U2750);
  not ginst10247 (P2_R2099_U20, P2_U2740);
  nand ginst10248 (P2_R2099_U200, P2_R2099_U147, P2_R2099_U8);
  nand ginst10249 (P2_R2099_U201, P2_R2099_U199, P2_R2099_U200);
  nand ginst10250 (P2_R2099_U202, P2_R2099_U105, P2_R2099_U8, P2_U2746);
  nand ginst10251 (P2_R2099_U203, P2_R2099_U108, P2_U2750);
  nand ginst10252 (P2_R2099_U204, P2_R2099_U43, P2_U2728);
  nand ginst10253 (P2_R2099_U205, P2_R2099_U134, P2_R2099_U44);
  nand ginst10254 (P2_R2099_U206, P2_R2099_U41, P2_U2729);
  nand ginst10255 (P2_R2099_U207, P2_R2099_U133, P2_R2099_U42);
  nand ginst10256 (P2_R2099_U208, P2_R2099_U39, P2_U2730);
  nand ginst10257 (P2_R2099_U209, P2_R2099_U132, P2_R2099_U40);
  nand ginst10258 (P2_R2099_U21, P2_R2099_U122, P2_U2740);
  nand ginst10259 (P2_R2099_U210, P2_R2099_U37, P2_U2731);
  nand ginst10260 (P2_R2099_U211, P2_R2099_U131, P2_R2099_U38);
  nand ginst10261 (P2_R2099_U212, P2_R2099_U35, P2_U2732);
  nand ginst10262 (P2_R2099_U213, P2_R2099_U130, P2_R2099_U36);
  nand ginst10263 (P2_R2099_U214, P2_R2099_U33, P2_U2733);
  nand ginst10264 (P2_R2099_U215, P2_R2099_U129, P2_R2099_U34);
  nand ginst10265 (P2_R2099_U216, P2_R2099_U31, P2_U2734);
  nand ginst10266 (P2_R2099_U217, P2_R2099_U128, P2_R2099_U32);
  nand ginst10267 (P2_R2099_U218, P2_R2099_U29, P2_U2735);
  nand ginst10268 (P2_R2099_U219, P2_R2099_U127, P2_R2099_U30);
  not ginst10269 (P2_R2099_U22, P2_U2739);
  nand ginst10270 (P2_R2099_U220, P2_R2099_U27, P2_U2736);
  nand ginst10271 (P2_R2099_U221, P2_R2099_U126, P2_R2099_U28);
  nand ginst10272 (P2_R2099_U222, P2_R2099_U25, P2_U2737);
  nand ginst10273 (P2_R2099_U223, P2_R2099_U125, P2_R2099_U26);
  nand ginst10274 (P2_R2099_U224, P2_R2099_U6, P2_U2751);
  nand ginst10275 (P2_R2099_U225, P2_R2099_U7, P2_U2747);
  not ginst10276 (P2_R2099_U23, P2_U2738);
  nand ginst10277 (P2_R2099_U24, P2_R2099_U123, P2_U2739);
  nand ginst10278 (P2_R2099_U25, P2_R2099_U124, P2_U2738);
  not ginst10279 (P2_R2099_U26, P2_U2737);
  nand ginst10280 (P2_R2099_U27, P2_R2099_U125, P2_U2737);
  not ginst10281 (P2_R2099_U28, P2_U2736);
  nand ginst10282 (P2_R2099_U29, P2_R2099_U126, P2_U2736);
  not ginst10283 (P2_R2099_U30, P2_U2735);
  nand ginst10284 (P2_R2099_U31, P2_R2099_U127, P2_U2735);
  not ginst10285 (P2_R2099_U32, P2_U2734);
  nand ginst10286 (P2_R2099_U33, P2_R2099_U128, P2_U2734);
  not ginst10287 (P2_R2099_U34, P2_U2733);
  nand ginst10288 (P2_R2099_U35, P2_R2099_U129, P2_U2733);
  not ginst10289 (P2_R2099_U36, P2_U2732);
  nand ginst10290 (P2_R2099_U37, P2_R2099_U130, P2_U2732);
  not ginst10291 (P2_R2099_U38, P2_U2731);
  nand ginst10292 (P2_R2099_U39, P2_R2099_U131, P2_U2731);
  not ginst10293 (P2_R2099_U40, P2_U2730);
  nand ginst10294 (P2_R2099_U41, P2_R2099_U132, P2_U2730);
  not ginst10295 (P2_R2099_U42, P2_U2729);
  nand ginst10296 (P2_R2099_U43, P2_R2099_U133, P2_U2729);
  not ginst10297 (P2_R2099_U44, P2_U2728);
  nand ginst10298 (P2_R2099_U45, P2_R2099_U134, P2_U2728);
  not ginst10299 (P2_R2099_U46, P2_U2727);
  nand ginst10300 (P2_R2099_U47, P2_R2099_U135, P2_U2727);
  not ginst10301 (P2_R2099_U48, P2_U2726);
  nand ginst10302 (P2_R2099_U49, P2_R2099_U136, P2_U2726);
  nand ginst10303 (P2_R2099_U5, P2_R2099_U107, P2_R2099_U148);
  not ginst10304 (P2_R2099_U50, P2_U2725);
  nand ginst10305 (P2_R2099_U51, P2_R2099_U137, P2_U2725);
  not ginst10306 (P2_R2099_U52, P2_U2724);
  nand ginst10307 (P2_R2099_U53, P2_R2099_U138, P2_U2724);
  not ginst10308 (P2_R2099_U54, P2_U2723);
  nand ginst10309 (P2_R2099_U55, P2_R2099_U139, P2_U2723);
  not ginst10310 (P2_R2099_U56, P2_U2722);
  nand ginst10311 (P2_R2099_U57, P2_R2099_U140, P2_U2722);
  not ginst10312 (P2_R2099_U58, P2_U2721);
  nand ginst10313 (P2_R2099_U59, P2_R2099_U141, P2_U2721);
  not ginst10314 (P2_R2099_U6, P2_U2747);
  not ginst10315 (P2_R2099_U60, P2_U2720);
  nand ginst10316 (P2_R2099_U61, P2_R2099_U142, P2_U2720);
  not ginst10317 (P2_R2099_U62, P2_U2719);
  nand ginst10318 (P2_R2099_U63, P2_R2099_U143, P2_U2719);
  not ginst10319 (P2_R2099_U64, P2_U2718);
  nand ginst10320 (P2_R2099_U65, P2_R2099_U144, P2_U2718);
  not ginst10321 (P2_R2099_U66, P2_U2717);
  nand ginst10322 (P2_R2099_U67, P2_R2099_U149, P2_R2099_U150);
  nand ginst10323 (P2_R2099_U68, P2_R2099_U151, P2_R2099_U152);
  nand ginst10324 (P2_R2099_U69, P2_R2099_U153, P2_R2099_U154);
  not ginst10325 (P2_R2099_U7, P2_U2751);
  nand ginst10326 (P2_R2099_U70, P2_R2099_U155, P2_R2099_U156);
  nand ginst10327 (P2_R2099_U71, P2_R2099_U157, P2_R2099_U158);
  nand ginst10328 (P2_R2099_U72, P2_R2099_U168, P2_R2099_U169);
  nand ginst10329 (P2_R2099_U73, P2_R2099_U170, P2_R2099_U171);
  nand ginst10330 (P2_R2099_U74, P2_R2099_U179, P2_R2099_U180);
  nand ginst10331 (P2_R2099_U75, P2_R2099_U181, P2_R2099_U182);
  nand ginst10332 (P2_R2099_U76, P2_R2099_U183, P2_R2099_U184);
  nand ginst10333 (P2_R2099_U77, P2_R2099_U185, P2_R2099_U186);
  nand ginst10334 (P2_R2099_U78, P2_R2099_U187, P2_R2099_U188);
  nand ginst10335 (P2_R2099_U79, P2_R2099_U189, P2_R2099_U190);
  not ginst10336 (P2_R2099_U8, P2_U2750);
  nand ginst10337 (P2_R2099_U80, P2_R2099_U191, P2_R2099_U192);
  nand ginst10338 (P2_R2099_U81, P2_R2099_U193, P2_R2099_U194);
  nand ginst10339 (P2_R2099_U82, P2_R2099_U195, P2_R2099_U196);
  nand ginst10340 (P2_R2099_U83, P2_R2099_U197, P2_R2099_U198);
  nand ginst10341 (P2_R2099_U84, P2_R2099_U204, P2_R2099_U205);
  nand ginst10342 (P2_R2099_U85, P2_R2099_U206, P2_R2099_U207);
  nand ginst10343 (P2_R2099_U86, P2_R2099_U208, P2_R2099_U209);
  nand ginst10344 (P2_R2099_U87, P2_R2099_U210, P2_R2099_U211);
  nand ginst10345 (P2_R2099_U88, P2_R2099_U212, P2_R2099_U213);
  nand ginst10346 (P2_R2099_U89, P2_R2099_U214, P2_R2099_U215);
  not ginst10347 (P2_R2099_U9, P2_U2746);
  nand ginst10348 (P2_R2099_U90, P2_R2099_U216, P2_R2099_U217);
  nand ginst10349 (P2_R2099_U91, P2_R2099_U218, P2_R2099_U219);
  nand ginst10350 (P2_R2099_U92, P2_R2099_U220, P2_R2099_U221);
  nand ginst10351 (P2_R2099_U93, P2_R2099_U222, P2_R2099_U223);
  nand ginst10352 (P2_R2099_U94, P2_R2099_U224, P2_R2099_U225);
  nand ginst10353 (P2_R2099_U95, P2_R2099_U166, P2_R2099_U167);
  nand ginst10354 (P2_R2099_U96, P2_R2099_U177, P2_R2099_U178);
  nand ginst10355 (P2_R2099_U97, P2_R2099_U117, P2_R2099_U118);
  and ginst10356 (P2_R2099_U98, P2_R2099_U159, P2_R2099_U160);
  and ginst10357 (P2_R2099_U99, P2_R2099_U161, P2_R2099_U162);
  not ginst10358 (P2_R2147_U10, P2_U2752);
  nand ginst10359 (P2_R2147_U11, P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN);
  nand ginst10360 (P2_R2147_U12, P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN);
  not ginst10361 (P2_R2147_U13, P2_R2147_U11);
  not ginst10362 (P2_R2147_U14, P2_R2147_U12);
  nand ginst10363 (P2_R2147_U15, P2_R2147_U11, P2_U2752);
  nand ginst10364 (P2_R2147_U16, P2_R2147_U10, P2_R2147_U13);
  nand ginst10365 (P2_R2147_U17, P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P2_R2147_U12);
  nand ginst10366 (P2_R2147_U18, P2_R2147_U14, P2_R2147_U5);
  nand ginst10367 (P2_R2147_U19, P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN, P2_R2147_U4);
  nand ginst10368 (P2_R2147_U20, P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P2_R2147_U6);
  not ginst10369 (P2_R2147_U4, P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN);
  not ginst10370 (P2_R2147_U5, P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN);
  not ginst10371 (P2_R2147_U6, P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN);
  nand ginst10372 (P2_R2147_U7, P2_R2147_U15, P2_R2147_U16);
  nand ginst10373 (P2_R2147_U8, P2_R2147_U17, P2_R2147_U18);
  nand ginst10374 (P2_R2147_U9, P2_R2147_U19, P2_R2147_U20);
  not ginst10375 (P2_R2167_U10, P2_U2705);
  not ginst10376 (P2_R2167_U11, P2_U2704);
  not ginst10377 (P2_R2167_U12, P2_U2711);
  not ginst10378 (P2_R2167_U13, P2_U2710);
  not ginst10379 (P2_R2167_U14, P2_U2703);
  not ginst10380 (P2_R2167_U15, P2_U2361);
  not ginst10381 (P2_R2167_U16, P2_U2709);
  not ginst10382 (P2_R2167_U17, P2_STATE2_REG_0__SCAN_IN);
  not ginst10383 (P2_R2167_U18, P2_U2708);
  nand ginst10384 (P2_R2167_U19, P2_U2714, P2_U2715);
  nand ginst10385 (P2_R2167_U20, P2_R2167_U19, P2_U2707);
  or ginst10386 (P2_R2167_U21, P2_U2714, P2_U2715);
  nand ginst10387 (P2_R2167_U22, P2_R2167_U8, P2_U2706);
  nand ginst10388 (P2_R2167_U23, P2_R2167_U20, P2_R2167_U21, P2_R2167_U22);
  nand ginst10389 (P2_R2167_U24, P2_R2167_U7, P2_U2713);
  nand ginst10390 (P2_R2167_U25, P2_R2167_U10, P2_U2712);
  nand ginst10391 (P2_R2167_U26, P2_R2167_U23, P2_R2167_U24, P2_R2167_U25);
  nand ginst10392 (P2_R2167_U27, P2_R2167_U9, P2_U2705);
  nand ginst10393 (P2_R2167_U28, P2_R2167_U12, P2_U2704);
  nand ginst10394 (P2_R2167_U29, P2_R2167_U26, P2_R2167_U27, P2_R2167_U28);
  nand ginst10395 (P2_R2167_U30, P2_R2167_U11, P2_U2711);
  nand ginst10396 (P2_R2167_U31, P2_R2167_U14, P2_U2710);
  nand ginst10397 (P2_R2167_U32, P2_R2167_U29, P2_R2167_U30, P2_R2167_U31);
  nand ginst10398 (P2_R2167_U33, P2_R2167_U13, P2_U2703);
  nand ginst10399 (P2_R2167_U34, P2_R2167_U16, P2_U2361);
  nand ginst10400 (P2_R2167_U35, P2_R2167_U32, P2_R2167_U33, P2_R2167_U34);
  nand ginst10401 (P2_R2167_U36, P2_R2167_U15, P2_U2709);
  nand ginst10402 (P2_R2167_U37, P2_R2167_U35, P2_R2167_U36);
  nand ginst10403 (P2_R2167_U38, P2_R2167_U37, P2_R2167_U39, P2_R2167_U40);
  nand ginst10404 (P2_R2167_U39, P2_R2167_U18, P2_U2361);
  nand ginst10405 (P2_R2167_U40, P2_R2167_U15, P2_U2708);
  nand ginst10406 (P2_R2167_U41, P2_STATE2_REG_0__SCAN_IN, P2_R2167_U18, P2_U2361);
  nand ginst10407 (P2_R2167_U42, P2_R2167_U15, P2_R2167_U17, P2_U2708);
  nand ginst10408 (P2_R2167_U6, P2_R2167_U38, P2_R2167_U41, P2_R2167_U42);
  not ginst10409 (P2_R2167_U7, P2_U2706);
  not ginst10410 (P2_R2167_U8, P2_U2713);
  not ginst10411 (P2_R2167_U9, P2_U2712);
  and ginst10412 (P2_R2182_U10, P2_R2182_U9, P2_U2674);
  and ginst10413 (P2_R2182_U100, P2_R2182_U125, P2_R2182_U191);
  nand ginst10414 (P2_R2182_U101, P2_R2182_U279, P2_R2182_U280);
  nand ginst10415 (P2_R2182_U102, P2_R2182_U134, P2_R2182_U135);
  and ginst10416 (P2_R2182_U103, P2_R2182_U203, P2_R2182_U204);
  nand ginst10417 (P2_R2182_U104, P2_R2182_U130, P2_R2182_U131);
  and ginst10418 (P2_R2182_U105, P2_R2182_U210, P2_R2182_U211);
  nand ginst10419 (P2_R2182_U106, P2_R2182_U126, P2_R2182_U127);
  not ginst10420 (P2_R2182_U107, P2_U2658);
  not ginst10421 (P2_R2182_U108, P2_U2682);
  and ginst10422 (P2_R2182_U109, P2_R2182_U224, P2_R2182_U225);
  and ginst10423 (P2_R2182_U11, P2_R2182_U13, P2_U2692);
  and ginst10424 (P2_R2182_U110, P2_R2182_U231, P2_R2182_U232);
  nand ginst10425 (P2_R2182_U111, P2_R2182_U172, P2_R2182_U173);
  and ginst10426 (P2_R2182_U112, P2_R2182_U238, P2_R2182_U239);
  nand ginst10427 (P2_R2182_U113, P2_R2182_U168, P2_R2182_U169);
  and ginst10428 (P2_R2182_U114, P2_R2182_U245, P2_R2182_U246);
  nand ginst10429 (P2_R2182_U115, P2_R2182_U164, P2_R2182_U165);
  and ginst10430 (P2_R2182_U116, P2_R2182_U252, P2_R2182_U253);
  nand ginst10431 (P2_R2182_U117, P2_R2182_U160, P2_R2182_U161);
  and ginst10432 (P2_R2182_U118, P2_R2182_U259, P2_R2182_U260);
  nand ginst10433 (P2_R2182_U119, P2_R2182_U156, P2_R2182_U157);
  and ginst10434 (P2_R2182_U12, P2_R2182_U18, P2_U2694);
  and ginst10435 (P2_R2182_U120, P2_R2182_U266, P2_R2182_U267);
  not ginst10436 (P2_R2182_U121, P2_R2182_U46);
  nand ginst10437 (P2_R2182_U122, P2_R2182_U121, P2_U2680);
  nand ginst10438 (P2_R2182_U123, P2_R2182_U122, P2_R2182_U67);
  or ginst10439 (P2_R2182_U124, P2_U2679, P2_U2700);
  nand ginst10440 (P2_R2182_U125, P2_R2182_U46, P2_R2182_U47);
  nand ginst10441 (P2_R2182_U126, P2_R2182_U123, P2_R2182_U124, P2_R2182_U125);
  nand ginst10442 (P2_R2182_U127, P2_U2679, P2_U2700);
  not ginst10443 (P2_R2182_U128, P2_R2182_U106);
  or ginst10444 (P2_R2182_U129, P2_U2678, P2_U2699);
  and ginst10445 (P2_R2182_U13, P2_R2182_U12, P2_U2693);
  nand ginst10446 (P2_R2182_U130, P2_R2182_U106, P2_R2182_U129);
  nand ginst10447 (P2_R2182_U131, P2_U2678, P2_U2699);
  not ginst10448 (P2_R2182_U132, P2_R2182_U104);
  or ginst10449 (P2_R2182_U133, P2_U2677, P2_U2698);
  nand ginst10450 (P2_R2182_U134, P2_R2182_U104, P2_R2182_U133);
  nand ginst10451 (P2_R2182_U135, P2_U2677, P2_U2698);
  not ginst10452 (P2_R2182_U136, P2_R2182_U102);
  not ginst10453 (P2_R2182_U137, P2_R2182_U21);
  not ginst10454 (P2_R2182_U138, P2_R2182_U9);
  not ginst10455 (P2_R2182_U139, P2_R2182_U10);
  and ginst10456 (P2_R2182_U14, P2_R2182_U6, P2_U2668);
  not ginst10457 (P2_R2182_U140, P2_R2182_U19);
  not ginst10458 (P2_R2182_U141, P2_R2182_U20);
  not ginst10459 (P2_R2182_U142, P2_R2182_U4);
  not ginst10460 (P2_R2182_U143, P2_R2182_U5);
  not ginst10461 (P2_R2182_U144, P2_R2182_U6);
  not ginst10462 (P2_R2182_U145, P2_R2182_U14);
  not ginst10463 (P2_R2182_U146, P2_R2182_U15);
  not ginst10464 (P2_R2182_U147, P2_R2182_U16);
  not ginst10465 (P2_R2182_U148, P2_R2182_U17);
  not ginst10466 (P2_R2182_U149, P2_R2182_U18);
  and ginst10467 (P2_R2182_U15, P2_R2182_U14, P2_U2667);
  not ginst10468 (P2_R2182_U150, P2_R2182_U12);
  not ginst10469 (P2_R2182_U151, P2_R2182_U13);
  not ginst10470 (P2_R2182_U152, P2_R2182_U11);
  not ginst10471 (P2_R2182_U153, P2_R2182_U8);
  not ginst10472 (P2_R2182_U154, P2_R2182_U7);
  or ginst10473 (P2_R2182_U155, P2_U2665, P2_U2689);
  nand ginst10474 (P2_R2182_U156, P2_R2182_U155, P2_R2182_U7);
  nand ginst10475 (P2_R2182_U157, P2_U2665, P2_U2689);
  not ginst10476 (P2_R2182_U158, P2_R2182_U119);
  or ginst10477 (P2_R2182_U159, P2_U2664, P2_U2688);
  and ginst10478 (P2_R2182_U16, P2_R2182_U15, P2_U2666);
  nand ginst10479 (P2_R2182_U160, P2_R2182_U119, P2_R2182_U159);
  nand ginst10480 (P2_R2182_U161, P2_U2664, P2_U2688);
  not ginst10481 (P2_R2182_U162, P2_R2182_U117);
  or ginst10482 (P2_R2182_U163, P2_U2663, P2_U2687);
  nand ginst10483 (P2_R2182_U164, P2_R2182_U117, P2_R2182_U163);
  nand ginst10484 (P2_R2182_U165, P2_U2663, P2_U2687);
  not ginst10485 (P2_R2182_U166, P2_R2182_U115);
  or ginst10486 (P2_R2182_U167, P2_U2662, P2_U2686);
  nand ginst10487 (P2_R2182_U168, P2_R2182_U115, P2_R2182_U167);
  nand ginst10488 (P2_R2182_U169, P2_U2662, P2_U2686);
  and ginst10489 (P2_R2182_U17, P2_R2182_U16, P2_U2696);
  not ginst10490 (P2_R2182_U170, P2_R2182_U113);
  or ginst10491 (P2_R2182_U171, P2_U2661, P2_U2685);
  nand ginst10492 (P2_R2182_U172, P2_R2182_U113, P2_R2182_U171);
  nand ginst10493 (P2_R2182_U173, P2_U2661, P2_U2685);
  not ginst10494 (P2_R2182_U174, P2_R2182_U111);
  or ginst10495 (P2_R2182_U175, P2_U2660, P2_U2684);
  nand ginst10496 (P2_R2182_U176, P2_R2182_U111, P2_R2182_U175);
  nand ginst10497 (P2_R2182_U177, P2_U2660, P2_U2684);
  not ginst10498 (P2_R2182_U178, P2_R2182_U66);
  or ginst10499 (P2_R2182_U179, P2_U2659, P2_U2683);
  and ginst10500 (P2_R2182_U18, P2_R2182_U17, P2_U2695);
  nand ginst10501 (P2_R2182_U180, P2_R2182_U179, P2_R2182_U66);
  nand ginst10502 (P2_R2182_U181, P2_U2659, P2_U2683);
  nand ginst10503 (P2_R2182_U182, P2_R2182_U180, P2_R2182_U97);
  nand ginst10504 (P2_R2182_U183, P2_U2659, P2_U2683);
  nand ginst10505 (P2_R2182_U184, P2_R2182_U178, P2_R2182_U183);
  or ginst10506 (P2_R2182_U185, P2_U2659, P2_U2683);
  nand ginst10507 (P2_R2182_U186, P2_R2182_U184, P2_R2182_U98);
  nand ginst10508 (P2_R2182_U187, P2_R2182_U46, P2_R2182_U47);
  nand ginst10509 (P2_R2182_U188, P2_R2182_U187, P2_U2701);
  nand ginst10510 (P2_R2182_U189, P2_R2182_U121, P2_U2680);
  and ginst10511 (P2_R2182_U19, P2_R2182_U10, P2_U2673);
  nand ginst10512 (P2_R2182_U190, P2_R2182_U188, P2_R2182_U99);
  nand ginst10513 (P2_R2182_U191, P2_U2679, P2_U2700);
  nand ginst10514 (P2_R2182_U192, P2_R2182_U100, P2_R2182_U123, P2_R2182_U124);
  nand ginst10515 (P2_R2182_U193, P2_R2182_U19, P2_R2182_U34);
  nand ginst10516 (P2_R2182_U194, P2_R2182_U140, P2_U2672);
  nand ginst10517 (P2_R2182_U195, P2_R2182_U10, P2_R2182_U36);
  nand ginst10518 (P2_R2182_U196, P2_R2182_U139, P2_U2673);
  nand ginst10519 (P2_R2182_U197, P2_R2182_U35, P2_R2182_U9);
  nand ginst10520 (P2_R2182_U198, P2_R2182_U138, P2_U2674);
  nand ginst10521 (P2_R2182_U199, P2_R2182_U21, P2_R2182_U22);
  and ginst10522 (P2_R2182_U20, P2_R2182_U19, P2_U2672);
  nand ginst10523 (P2_R2182_U200, P2_R2182_U137, P2_U2675);
  nand ginst10524 (P2_R2182_U201, P2_R2182_U102, P2_R2182_U24);
  nand ginst10525 (P2_R2182_U202, P2_R2182_U136, P2_U2676);
  nand ginst10526 (P2_R2182_U203, P2_R2182_U50, P2_U2677);
  nand ginst10527 (P2_R2182_U204, P2_R2182_U51, P2_U2698);
  nand ginst10528 (P2_R2182_U205, P2_R2182_U50, P2_U2677);
  nand ginst10529 (P2_R2182_U206, P2_R2182_U51, P2_U2698);
  nand ginst10530 (P2_R2182_U207, P2_R2182_U205, P2_R2182_U206);
  nand ginst10531 (P2_R2182_U208, P2_R2182_U103, P2_R2182_U104);
  nand ginst10532 (P2_R2182_U209, P2_R2182_U132, P2_R2182_U207);
  and ginst10533 (P2_R2182_U21, P2_R2182_U102, P2_U2676);
  nand ginst10534 (P2_R2182_U210, P2_R2182_U48, P2_U2678);
  nand ginst10535 (P2_R2182_U211, P2_R2182_U49, P2_U2699);
  nand ginst10536 (P2_R2182_U212, P2_R2182_U48, P2_U2678);
  nand ginst10537 (P2_R2182_U213, P2_R2182_U49, P2_U2699);
  nand ginst10538 (P2_R2182_U214, P2_R2182_U212, P2_R2182_U213);
  nand ginst10539 (P2_R2182_U215, P2_R2182_U105, P2_R2182_U106);
  nand ginst10540 (P2_R2182_U216, P2_R2182_U128, P2_R2182_U214);
  nand ginst10541 (P2_R2182_U217, P2_R2182_U108, P2_U2658);
  nand ginst10542 (P2_R2182_U218, P2_R2182_U107, P2_U2682);
  nand ginst10543 (P2_R2182_U219, P2_R2182_U108, P2_U2658);
  not ginst10544 (P2_R2182_U22, P2_U2675);
  nand ginst10545 (P2_R2182_U220, P2_R2182_U107, P2_U2682);
  nand ginst10546 (P2_R2182_U221, P2_R2182_U219, P2_R2182_U220);
  nand ginst10547 (P2_R2182_U222, P2_R2182_U42, P2_U2679);
  nand ginst10548 (P2_R2182_U223, P2_R2182_U43, P2_U2700);
  nand ginst10549 (P2_R2182_U224, P2_R2182_U64, P2_U2659);
  nand ginst10550 (P2_R2182_U225, P2_R2182_U65, P2_U2683);
  nand ginst10551 (P2_R2182_U226, P2_R2182_U64, P2_U2659);
  nand ginst10552 (P2_R2182_U227, P2_R2182_U65, P2_U2683);
  nand ginst10553 (P2_R2182_U228, P2_R2182_U226, P2_R2182_U227);
  nand ginst10554 (P2_R2182_U229, P2_R2182_U109, P2_R2182_U66);
  not ginst10555 (P2_R2182_U23, P2_U2671);
  nand ginst10556 (P2_R2182_U230, P2_R2182_U178, P2_R2182_U228);
  nand ginst10557 (P2_R2182_U231, P2_R2182_U62, P2_U2660);
  nand ginst10558 (P2_R2182_U232, P2_R2182_U63, P2_U2684);
  nand ginst10559 (P2_R2182_U233, P2_R2182_U62, P2_U2660);
  nand ginst10560 (P2_R2182_U234, P2_R2182_U63, P2_U2684);
  nand ginst10561 (P2_R2182_U235, P2_R2182_U233, P2_R2182_U234);
  nand ginst10562 (P2_R2182_U236, P2_R2182_U110, P2_R2182_U111);
  nand ginst10563 (P2_R2182_U237, P2_R2182_U174, P2_R2182_U235);
  nand ginst10564 (P2_R2182_U238, P2_R2182_U60, P2_U2661);
  nand ginst10565 (P2_R2182_U239, P2_R2182_U61, P2_U2685);
  not ginst10566 (P2_R2182_U24, P2_U2676);
  nand ginst10567 (P2_R2182_U240, P2_R2182_U60, P2_U2661);
  nand ginst10568 (P2_R2182_U241, P2_R2182_U61, P2_U2685);
  nand ginst10569 (P2_R2182_U242, P2_R2182_U240, P2_R2182_U241);
  nand ginst10570 (P2_R2182_U243, P2_R2182_U112, P2_R2182_U113);
  nand ginst10571 (P2_R2182_U244, P2_R2182_U170, P2_R2182_U242);
  nand ginst10572 (P2_R2182_U245, P2_R2182_U58, P2_U2662);
  nand ginst10573 (P2_R2182_U246, P2_R2182_U59, P2_U2686);
  nand ginst10574 (P2_R2182_U247, P2_R2182_U58, P2_U2662);
  nand ginst10575 (P2_R2182_U248, P2_R2182_U59, P2_U2686);
  nand ginst10576 (P2_R2182_U249, P2_R2182_U247, P2_R2182_U248);
  not ginst10577 (P2_R2182_U25, P2_U2666);
  nand ginst10578 (P2_R2182_U250, P2_R2182_U114, P2_R2182_U115);
  nand ginst10579 (P2_R2182_U251, P2_R2182_U166, P2_R2182_U249);
  nand ginst10580 (P2_R2182_U252, P2_R2182_U56, P2_U2663);
  nand ginst10581 (P2_R2182_U253, P2_R2182_U57, P2_U2687);
  nand ginst10582 (P2_R2182_U254, P2_R2182_U56, P2_U2663);
  nand ginst10583 (P2_R2182_U255, P2_R2182_U57, P2_U2687);
  nand ginst10584 (P2_R2182_U256, P2_R2182_U254, P2_R2182_U255);
  nand ginst10585 (P2_R2182_U257, P2_R2182_U116, P2_R2182_U117);
  nand ginst10586 (P2_R2182_U258, P2_R2182_U162, P2_R2182_U256);
  nand ginst10587 (P2_R2182_U259, P2_R2182_U54, P2_U2664);
  not ginst10588 (P2_R2182_U26, P2_U2667);
  nand ginst10589 (P2_R2182_U260, P2_R2182_U55, P2_U2688);
  nand ginst10590 (P2_R2182_U261, P2_R2182_U54, P2_U2664);
  nand ginst10591 (P2_R2182_U262, P2_R2182_U55, P2_U2688);
  nand ginst10592 (P2_R2182_U263, P2_R2182_U261, P2_R2182_U262);
  nand ginst10593 (P2_R2182_U264, P2_R2182_U118, P2_R2182_U119);
  nand ginst10594 (P2_R2182_U265, P2_R2182_U158, P2_R2182_U263);
  nand ginst10595 (P2_R2182_U266, P2_R2182_U52, P2_U2665);
  nand ginst10596 (P2_R2182_U267, P2_R2182_U53, P2_U2689);
  nand ginst10597 (P2_R2182_U268, P2_R2182_U52, P2_U2665);
  nand ginst10598 (P2_R2182_U269, P2_R2182_U53, P2_U2689);
  not ginst10599 (P2_R2182_U27, P2_U2696);
  nand ginst10600 (P2_R2182_U270, P2_R2182_U268, P2_R2182_U269);
  nand ginst10601 (P2_R2182_U271, P2_R2182_U120, P2_R2182_U7);
  nand ginst10602 (P2_R2182_U272, P2_R2182_U154, P2_R2182_U270);
  nand ginst10603 (P2_R2182_U273, P2_R2182_U37, P2_R2182_U8);
  nand ginst10604 (P2_R2182_U274, P2_R2182_U153, P2_U2690);
  nand ginst10605 (P2_R2182_U275, P2_R2182_U11, P2_R2182_U32);
  nand ginst10606 (P2_R2182_U276, P2_R2182_U152, P2_U2691);
  nand ginst10607 (P2_R2182_U277, P2_R2182_U13, P2_R2182_U31);
  nand ginst10608 (P2_R2182_U278, P2_R2182_U151, P2_U2692);
  nand ginst10609 (P2_R2182_U279, P2_R2182_U121, P2_R2182_U47);
  not ginst10610 (P2_R2182_U28, P2_U2695);
  nand ginst10611 (P2_R2182_U280, P2_R2182_U46, P2_U2680);
  not ginst10612 (P2_R2182_U281, P2_R2182_U101);
  nand ginst10613 (P2_R2182_U282, P2_R2182_U281, P2_U2701);
  nand ginst10614 (P2_R2182_U283, P2_R2182_U101, P2_R2182_U67);
  nand ginst10615 (P2_R2182_U284, P2_R2182_U12, P2_R2182_U30);
  nand ginst10616 (P2_R2182_U285, P2_R2182_U150, P2_U2693);
  nand ginst10617 (P2_R2182_U286, P2_R2182_U18, P2_R2182_U29);
  nand ginst10618 (P2_R2182_U287, P2_R2182_U149, P2_U2694);
  nand ginst10619 (P2_R2182_U288, P2_R2182_U17, P2_R2182_U28);
  nand ginst10620 (P2_R2182_U289, P2_R2182_U148, P2_U2695);
  not ginst10621 (P2_R2182_U29, P2_U2694);
  nand ginst10622 (P2_R2182_U290, P2_R2182_U16, P2_R2182_U27);
  nand ginst10623 (P2_R2182_U291, P2_R2182_U147, P2_U2696);
  nand ginst10624 (P2_R2182_U292, P2_R2182_U15, P2_R2182_U25);
  nand ginst10625 (P2_R2182_U293, P2_R2182_U146, P2_U2666);
  nand ginst10626 (P2_R2182_U294, P2_R2182_U14, P2_R2182_U26);
  nand ginst10627 (P2_R2182_U295, P2_R2182_U145, P2_U2667);
  nand ginst10628 (P2_R2182_U296, P2_R2182_U38, P2_R2182_U6);
  nand ginst10629 (P2_R2182_U297, P2_R2182_U144, P2_U2668);
  nand ginst10630 (P2_R2182_U298, P2_R2182_U39, P2_R2182_U5);
  nand ginst10631 (P2_R2182_U299, P2_R2182_U143, P2_U2669);
  not ginst10632 (P2_R2182_U30, P2_U2693);
  nand ginst10633 (P2_R2182_U300, P2_R2182_U33, P2_R2182_U4);
  nand ginst10634 (P2_R2182_U301, P2_R2182_U142, P2_U2670);
  nand ginst10635 (P2_R2182_U302, P2_R2182_U20, P2_R2182_U23);
  nand ginst10636 (P2_R2182_U303, P2_R2182_U141, P2_U2671);
  nand ginst10637 (P2_R2182_U304, P2_R2182_U44, P2_U2681);
  nand ginst10638 (P2_R2182_U305, P2_R2182_U45, P2_U2702);
  not ginst10639 (P2_R2182_U31, P2_U2692);
  not ginst10640 (P2_R2182_U32, P2_U2691);
  not ginst10641 (P2_R2182_U33, P2_U2670);
  not ginst10642 (P2_R2182_U34, P2_U2672);
  not ginst10643 (P2_R2182_U35, P2_U2674);
  not ginst10644 (P2_R2182_U36, P2_U2673);
  not ginst10645 (P2_R2182_U37, P2_U2690);
  not ginst10646 (P2_R2182_U38, P2_U2668);
  not ginst10647 (P2_R2182_U39, P2_U2669);
  and ginst10648 (P2_R2182_U4, P2_R2182_U20, P2_U2671);
  and ginst10649 (P2_R2182_U40, P2_R2182_U190, P2_R2182_U192);
  and ginst10650 (P2_R2182_U41, P2_R2182_U182, P2_R2182_U186);
  not ginst10651 (P2_R2182_U42, P2_U2700);
  not ginst10652 (P2_R2182_U43, P2_U2679);
  not ginst10653 (P2_R2182_U44, P2_U2702);
  not ginst10654 (P2_R2182_U45, P2_U2681);
  nand ginst10655 (P2_R2182_U46, P2_U2681, P2_U2702);
  not ginst10656 (P2_R2182_U47, P2_U2680);
  not ginst10657 (P2_R2182_U48, P2_U2699);
  not ginst10658 (P2_R2182_U49, P2_U2678);
  and ginst10659 (P2_R2182_U5, P2_R2182_U4, P2_U2670);
  not ginst10660 (P2_R2182_U50, P2_U2698);
  not ginst10661 (P2_R2182_U51, P2_U2677);
  not ginst10662 (P2_R2182_U52, P2_U2689);
  not ginst10663 (P2_R2182_U53, P2_U2665);
  not ginst10664 (P2_R2182_U54, P2_U2688);
  not ginst10665 (P2_R2182_U55, P2_U2664);
  not ginst10666 (P2_R2182_U56, P2_U2687);
  not ginst10667 (P2_R2182_U57, P2_U2663);
  not ginst10668 (P2_R2182_U58, P2_U2686);
  not ginst10669 (P2_R2182_U59, P2_U2662);
  and ginst10670 (P2_R2182_U6, P2_R2182_U5, P2_U2669);
  not ginst10671 (P2_R2182_U60, P2_U2685);
  not ginst10672 (P2_R2182_U61, P2_U2661);
  not ginst10673 (P2_R2182_U62, P2_U2684);
  not ginst10674 (P2_R2182_U63, P2_U2660);
  not ginst10675 (P2_R2182_U64, P2_U2683);
  not ginst10676 (P2_R2182_U65, P2_U2659);
  nand ginst10677 (P2_R2182_U66, P2_R2182_U176, P2_R2182_U177);
  not ginst10678 (P2_R2182_U67, P2_U2701);
  nand ginst10679 (P2_R2182_U68, P2_R2182_U282, P2_R2182_U283);
  nand ginst10680 (P2_R2182_U69, P2_R2182_U304, P2_R2182_U305);
  and ginst10681 (P2_R2182_U7, P2_R2182_U8, P2_U2690);
  nand ginst10682 (P2_R2182_U70, P2_R2182_U193, P2_R2182_U194);
  nand ginst10683 (P2_R2182_U71, P2_R2182_U195, P2_R2182_U196);
  nand ginst10684 (P2_R2182_U72, P2_R2182_U197, P2_R2182_U198);
  nand ginst10685 (P2_R2182_U73, P2_R2182_U199, P2_R2182_U200);
  nand ginst10686 (P2_R2182_U74, P2_R2182_U201, P2_R2182_U202);
  nand ginst10687 (P2_R2182_U75, P2_R2182_U208, P2_R2182_U209);
  nand ginst10688 (P2_R2182_U76, P2_R2182_U215, P2_R2182_U216);
  nand ginst10689 (P2_R2182_U77, P2_R2182_U229, P2_R2182_U230);
  nand ginst10690 (P2_R2182_U78, P2_R2182_U236, P2_R2182_U237);
  nand ginst10691 (P2_R2182_U79, P2_R2182_U243, P2_R2182_U244);
  and ginst10692 (P2_R2182_U8, P2_R2182_U11, P2_U2691);
  nand ginst10693 (P2_R2182_U80, P2_R2182_U250, P2_R2182_U251);
  nand ginst10694 (P2_R2182_U81, P2_R2182_U257, P2_R2182_U258);
  nand ginst10695 (P2_R2182_U82, P2_R2182_U264, P2_R2182_U265);
  nand ginst10696 (P2_R2182_U83, P2_R2182_U271, P2_R2182_U272);
  nand ginst10697 (P2_R2182_U84, P2_R2182_U273, P2_R2182_U274);
  nand ginst10698 (P2_R2182_U85, P2_R2182_U275, P2_R2182_U276);
  nand ginst10699 (P2_R2182_U86, P2_R2182_U277, P2_R2182_U278);
  nand ginst10700 (P2_R2182_U87, P2_R2182_U284, P2_R2182_U285);
  nand ginst10701 (P2_R2182_U88, P2_R2182_U286, P2_R2182_U287);
  nand ginst10702 (P2_R2182_U89, P2_R2182_U288, P2_R2182_U289);
  and ginst10703 (P2_R2182_U9, P2_R2182_U21, P2_U2675);
  nand ginst10704 (P2_R2182_U90, P2_R2182_U290, P2_R2182_U291);
  nand ginst10705 (P2_R2182_U91, P2_R2182_U292, P2_R2182_U293);
  nand ginst10706 (P2_R2182_U92, P2_R2182_U294, P2_R2182_U295);
  nand ginst10707 (P2_R2182_U93, P2_R2182_U296, P2_R2182_U297);
  nand ginst10708 (P2_R2182_U94, P2_R2182_U298, P2_R2182_U299);
  nand ginst10709 (P2_R2182_U95, P2_R2182_U300, P2_R2182_U301);
  nand ginst10710 (P2_R2182_U96, P2_R2182_U302, P2_R2182_U303);
  and ginst10711 (P2_R2182_U97, P2_R2182_U181, P2_R2182_U217, P2_R2182_U218);
  and ginst10712 (P2_R2182_U98, P2_R2182_U185, P2_R2182_U221);
  and ginst10713 (P2_R2182_U99, P2_R2182_U189, P2_R2182_U222, P2_R2182_U223);
  not ginst10714 (P2_R2219_U10, P2_U2753);
  nand ginst10715 (P2_R2219_U100, P2_R2219_U54, P2_R2219_U99);
  nand ginst10716 (P2_R2219_U101, P2_R2219_U35, P2_R2219_U42);
  nand ginst10717 (P2_R2219_U102, P2_R2219_U18, P2_U2762);
  nand ginst10718 (P2_R2219_U103, P2_R2219_U13, P2_U2754);
  not ginst10719 (P2_R2219_U104, P2_R2219_U36);
  nand ginst10720 (P2_R2219_U105, P2_R2219_U104, P2_R2219_U51);
  nand ginst10721 (P2_R2219_U106, P2_R2219_U36, P2_R2219_U43);
  nand ginst10722 (P2_R2219_U107, P2_R2219_U17, P2_U2763);
  nand ginst10723 (P2_R2219_U108, P2_R2219_U12, P2_U2755);
  not ginst10724 (P2_R2219_U109, P2_R2219_U37);
  not ginst10725 (P2_R2219_U11, P2_U2761);
  nand ginst10726 (P2_R2219_U110, P2_R2219_U109, P2_R2219_U79);
  nand ginst10727 (P2_R2219_U111, P2_R2219_U37, P2_R2219_U44);
  nand ginst10728 (P2_R2219_U112, P2_R2219_U14, P2_U2764);
  nand ginst10729 (P2_R2219_U113, P2_R2219_U16, P2_U2756);
  not ginst10730 (P2_R2219_U114, P2_R2219_U38);
  nand ginst10731 (P2_R2219_U115, P2_R2219_U114, P2_R2219_U46);
  nand ginst10732 (P2_R2219_U116, P2_R2219_U38, P2_R2219_U45);
  not ginst10733 (P2_R2219_U12, P2_U2763);
  not ginst10734 (P2_R2219_U13, P2_U2762);
  not ginst10735 (P2_R2219_U14, P2_U2756);
  not ginst10736 (P2_R2219_U15, P2_U2765);
  not ginst10737 (P2_R2219_U16, P2_U2764);
  not ginst10738 (P2_R2219_U17, P2_U2755);
  not ginst10739 (P2_R2219_U18, P2_U2754);
  nand ginst10740 (P2_R2219_U19, P2_R2219_U72, P2_R2219_U76);
  not ginst10741 (P2_R2219_U20, P2_U2760);
  not ginst10742 (P2_R2219_U21, P2_U2759);
  not ginst10743 (P2_R2219_U22, P2_U2758);
  not ginst10744 (P2_R2219_U23, P2_U2757);
  nand ginst10745 (P2_R2219_U24, P2_R2219_U85, P2_R2219_U86);
  nand ginst10746 (P2_R2219_U25, P2_R2219_U90, P2_R2219_U91);
  nand ginst10747 (P2_R2219_U26, P2_R2219_U95, P2_R2219_U96);
  nand ginst10748 (P2_R2219_U27, P2_R2219_U100, P2_R2219_U101);
  nand ginst10749 (P2_R2219_U28, P2_R2219_U105, P2_R2219_U106);
  nand ginst10750 (P2_R2219_U29, P2_R2219_U110, P2_R2219_U111);
  nand ginst10751 (P2_R2219_U30, P2_R2219_U115, P2_R2219_U116);
  and ginst10752 (P2_R2219_U31, P2_R2219_U55, P2_R2219_U6);
  nand ginst10753 (P2_R2219_U32, P2_R2219_U82, P2_R2219_U83);
  nand ginst10754 (P2_R2219_U33, P2_R2219_U87, P2_R2219_U88);
  nand ginst10755 (P2_R2219_U34, P2_R2219_U92, P2_R2219_U93);
  nand ginst10756 (P2_R2219_U35, P2_R2219_U97, P2_R2219_U98);
  nand ginst10757 (P2_R2219_U36, P2_R2219_U102, P2_R2219_U103);
  nand ginst10758 (P2_R2219_U37, P2_R2219_U107, P2_R2219_U108);
  nand ginst10759 (P2_R2219_U38, P2_R2219_U112, P2_R2219_U113);
  nand ginst10760 (P2_R2219_U39, P2_R2219_U63, P2_R2219_U64);
  nand ginst10761 (P2_R2219_U40, P2_R2219_U59, P2_R2219_U60);
  nand ginst10762 (P2_R2219_U41, P2_R2219_U56, P2_R2219_U74, P2_R2219_U75);
  nand ginst10763 (P2_R2219_U42, P2_R2219_U19, P2_R2219_U71);
  nand ginst10764 (P2_R2219_U43, P2_R2219_U49, P2_R2219_U50);
  nand ginst10765 (P2_R2219_U44, P2_R2219_U70, P2_R2219_U78);
  nand ginst10766 (P2_R2219_U45, P2_R2219_U23, P2_U2765);
  not ginst10767 (P2_R2219_U46, P2_R2219_U45);
  nand ginst10768 (P2_R2219_U47, P2_R2219_U14, P2_U2764);
  nand ginst10769 (P2_R2219_U48, P2_R2219_U17, P2_U2763);
  nand ginst10770 (P2_R2219_U49, P2_R2219_U48, P2_R2219_U81);
  nand ginst10771 (P2_R2219_U50, P2_R2219_U12, P2_U2755);
  not ginst10772 (P2_R2219_U51, P2_R2219_U43);
  nand ginst10773 (P2_R2219_U52, P2_R2219_U18, P2_U2762);
  nand ginst10774 (P2_R2219_U53, P2_R2219_U13, P2_U2754);
  not ginst10775 (P2_R2219_U54, P2_R2219_U42);
  nand ginst10776 (P2_R2219_U55, P2_R2219_U10, P2_U2761);
  nand ginst10777 (P2_R2219_U56, P2_R2219_U11, P2_U2753);
  not ginst10778 (P2_R2219_U57, P2_R2219_U41);
  nand ginst10779 (P2_R2219_U58, P2_R2219_U9, P2_U2760);
  nand ginst10780 (P2_R2219_U59, P2_R2219_U41, P2_R2219_U58);
  and ginst10781 (P2_R2219_U6, P2_R2219_U48, P2_R2219_U52);
  nand ginst10782 (P2_R2219_U60, P2_R2219_U20, P2_U4428);
  not ginst10783 (P2_R2219_U61, P2_R2219_U40);
  nand ginst10784 (P2_R2219_U62, P2_R2219_U9, P2_U2759);
  nand ginst10785 (P2_R2219_U63, P2_R2219_U40, P2_R2219_U62);
  nand ginst10786 (P2_R2219_U64, P2_R2219_U21, P2_U4428);
  not ginst10787 (P2_R2219_U65, P2_R2219_U39);
  nand ginst10788 (P2_R2219_U66, P2_R2219_U22, P2_U4428);
  nand ginst10789 (P2_R2219_U67, P2_R2219_U9, P2_U2758);
  nand ginst10790 (P2_R2219_U68, P2_R2219_U39, P2_R2219_U67);
  nand ginst10791 (P2_R2219_U69, P2_R2219_U15, P2_U2757);
  and ginst10792 (P2_R2219_U7, P2_R2219_U66, P2_R2219_U68);
  nand ginst10793 (P2_R2219_U70, P2_R2219_U16, P2_U2756);
  nand ginst10794 (P2_R2219_U71, P2_R2219_U44, P2_R2219_U6);
  nand ginst10795 (P2_R2219_U72, P2_R2219_U50, P2_R2219_U53);
  not ginst10796 (P2_R2219_U73, P2_R2219_U19);
  nand ginst10797 (P2_R2219_U74, P2_R2219_U31, P2_R2219_U44);
  nand ginst10798 (P2_R2219_U75, P2_R2219_U55, P2_R2219_U73);
  nand ginst10799 (P2_R2219_U76, P2_R2219_U18, P2_U2762);
  nand ginst10800 (P2_R2219_U77, P2_R2219_U14, P2_U2764);
  nand ginst10801 (P2_R2219_U78, P2_R2219_U45, P2_R2219_U47);
  not ginst10802 (P2_R2219_U79, P2_R2219_U44);
  nand ginst10803 (P2_R2219_U8, P2_R2219_U45, P2_R2219_U69);
  nand ginst10804 (P2_R2219_U80, P2_R2219_U45, P2_R2219_U77);
  nand ginst10805 (P2_R2219_U81, P2_R2219_U70, P2_R2219_U80);
  nand ginst10806 (P2_R2219_U82, P2_R2219_U9, P2_U2758);
  nand ginst10807 (P2_R2219_U83, P2_R2219_U22, P2_U4428);
  not ginst10808 (P2_R2219_U84, P2_R2219_U32);
  nand ginst10809 (P2_R2219_U85, P2_R2219_U65, P2_R2219_U84);
  nand ginst10810 (P2_R2219_U86, P2_R2219_U32, P2_R2219_U39);
  nand ginst10811 (P2_R2219_U87, P2_R2219_U9, P2_U2759);
  nand ginst10812 (P2_R2219_U88, P2_R2219_U21, P2_U4428);
  not ginst10813 (P2_R2219_U89, P2_R2219_U33);
  not ginst10814 (P2_R2219_U9, P2_U4428);
  nand ginst10815 (P2_R2219_U90, P2_R2219_U61, P2_R2219_U89);
  nand ginst10816 (P2_R2219_U91, P2_R2219_U33, P2_R2219_U40);
  nand ginst10817 (P2_R2219_U92, P2_R2219_U9, P2_U2760);
  nand ginst10818 (P2_R2219_U93, P2_R2219_U20, P2_U4428);
  not ginst10819 (P2_R2219_U94, P2_R2219_U34);
  nand ginst10820 (P2_R2219_U95, P2_R2219_U57, P2_R2219_U94);
  nand ginst10821 (P2_R2219_U96, P2_R2219_U34, P2_R2219_U41);
  nand ginst10822 (P2_R2219_U97, P2_R2219_U10, P2_U2761);
  nand ginst10823 (P2_R2219_U98, P2_R2219_U11, P2_U2753);
  not ginst10824 (P2_R2219_U99, P2_R2219_U35);
  not ginst10825 (P2_R2238_U10, P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN);
  not ginst10826 (P2_R2238_U11, P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN);
  not ginst10827 (P2_R2238_U12, P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN);
  not ginst10828 (P2_R2238_U13, P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN);
  not ginst10829 (P2_R2238_U14, P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN);
  not ginst10830 (P2_R2238_U15, P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN);
  nand ginst10831 (P2_R2238_U16, P2_R2238_U40, P2_R2238_U41);
  not ginst10832 (P2_R2238_U17, P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN);
  not ginst10833 (P2_R2238_U18, P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN);
  nand ginst10834 (P2_R2238_U19, P2_R2238_U50, P2_R2238_U51);
  nand ginst10835 (P2_R2238_U20, P2_R2238_U55, P2_R2238_U56);
  nand ginst10836 (P2_R2238_U21, P2_R2238_U60, P2_R2238_U61);
  nand ginst10837 (P2_R2238_U22, P2_R2238_U65, P2_R2238_U66);
  nand ginst10838 (P2_R2238_U23, P2_R2238_U47, P2_R2238_U48);
  nand ginst10839 (P2_R2238_U24, P2_R2238_U52, P2_R2238_U53);
  nand ginst10840 (P2_R2238_U25, P2_R2238_U57, P2_R2238_U58);
  nand ginst10841 (P2_R2238_U26, P2_R2238_U62, P2_R2238_U63);
  nand ginst10842 (P2_R2238_U27, P2_R2238_U36, P2_R2238_U37);
  nand ginst10843 (P2_R2238_U28, P2_R2238_U32, P2_R2238_U33);
  not ginst10844 (P2_R2238_U29, P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN);
  not ginst10845 (P2_R2238_U30, P2_R2238_U9);
  nand ginst10846 (P2_R2238_U31, P2_R2238_U10, P2_R2238_U30);
  nand ginst10847 (P2_R2238_U32, P2_R2238_U29, P2_R2238_U31);
  nand ginst10848 (P2_R2238_U33, P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN, P2_R2238_U9);
  not ginst10849 (P2_R2238_U34, P2_R2238_U28);
  nand ginst10850 (P2_R2238_U35, P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN, P2_R2238_U12);
  nand ginst10851 (P2_R2238_U36, P2_R2238_U28, P2_R2238_U35);
  nand ginst10852 (P2_R2238_U37, P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN, P2_R2238_U11);
  not ginst10853 (P2_R2238_U38, P2_R2238_U27);
  nand ginst10854 (P2_R2238_U39, P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P2_R2238_U14);
  nand ginst10855 (P2_R2238_U40, P2_R2238_U27, P2_R2238_U39);
  nand ginst10856 (P2_R2238_U41, P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN, P2_R2238_U13);
  not ginst10857 (P2_R2238_U42, P2_R2238_U16);
  nand ginst10858 (P2_R2238_U43, P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN, P2_R2238_U17);
  nand ginst10859 (P2_R2238_U44, P2_R2238_U42, P2_R2238_U43);
  nand ginst10860 (P2_R2238_U45, P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN, P2_R2238_U15);
  nand ginst10861 (P2_R2238_U46, P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P2_R2238_U8);
  nand ginst10862 (P2_R2238_U47, P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN, P2_R2238_U15);
  nand ginst10863 (P2_R2238_U48, P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN, P2_R2238_U17);
  not ginst10864 (P2_R2238_U49, P2_R2238_U23);
  nand ginst10865 (P2_R2238_U50, P2_R2238_U42, P2_R2238_U49);
  nand ginst10866 (P2_R2238_U51, P2_R2238_U16, P2_R2238_U23);
  nand ginst10867 (P2_R2238_U52, P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P2_R2238_U14);
  nand ginst10868 (P2_R2238_U53, P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN, P2_R2238_U13);
  not ginst10869 (P2_R2238_U54, P2_R2238_U24);
  nand ginst10870 (P2_R2238_U55, P2_R2238_U38, P2_R2238_U54);
  nand ginst10871 (P2_R2238_U56, P2_R2238_U24, P2_R2238_U27);
  nand ginst10872 (P2_R2238_U57, P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN, P2_R2238_U12);
  nand ginst10873 (P2_R2238_U58, P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN, P2_R2238_U11);
  not ginst10874 (P2_R2238_U59, P2_R2238_U25);
  nand ginst10875 (P2_R2238_U6, P2_R2238_U44, P2_R2238_U45);
  nand ginst10876 (P2_R2238_U60, P2_R2238_U34, P2_R2238_U59);
  nand ginst10877 (P2_R2238_U61, P2_R2238_U25, P2_R2238_U28);
  nand ginst10878 (P2_R2238_U62, P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P2_R2238_U10);
  nand ginst10879 (P2_R2238_U63, P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN, P2_R2238_U29);
  not ginst10880 (P2_R2238_U64, P2_R2238_U26);
  nand ginst10881 (P2_R2238_U65, P2_R2238_U30, P2_R2238_U64);
  nand ginst10882 (P2_R2238_U66, P2_R2238_U26, P2_R2238_U9);
  nand ginst10883 (P2_R2238_U7, P2_R2238_U46, P2_R2238_U9);
  not ginst10884 (P2_R2238_U8, P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN);
  nand ginst10885 (P2_R2238_U9, P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN, P2_R2238_U18);
  not ginst10886 (P2_R2243_U10, P2_U3688);
  nand ginst10887 (P2_R2243_U11, P2_R2243_U10, P2_R2243_U6);
  nor ginst10888 (P2_R2243_U6, P2_U3684, P2_U3685, P2_U3686, P2_U3687);
  nor ginst10889 (P2_R2243_U7, P2_R2243_U9, P2_U3684);
  nand ginst10890 (P2_R2243_U8, P2_R2243_U11, P2_R2243_U7);
  nor ginst10891 (P2_R2243_U9, P2_U3684, P2_U3685, P2_U3686, P2_U3687, P2_U3689);
  nand ginst10892 (P2_R2256_U10, P2_R2256_U25, P2_U3626);
  not ginst10893 (P2_R2256_U11, P2_U3625);
  nand ginst10894 (P2_R2256_U12, P2_R2256_U41, P2_U3625);
  not ginst10895 (P2_R2256_U13, P2_U3624);
  nand ginst10896 (P2_R2256_U14, P2_R2256_U42, P2_U3624);
  not ginst10897 (P2_R2256_U15, P2_U3622);
  not ginst10898 (P2_R2256_U16, P2_U3623);
  nand ginst10899 (P2_R2256_U17, P2_R2256_U47, P2_R2256_U48);
  nand ginst10900 (P2_R2256_U18, P2_R2256_U49, P2_R2256_U50);
  nand ginst10901 (P2_R2256_U19, P2_R2256_U51, P2_R2256_U52);
  nand ginst10902 (P2_R2256_U20, P2_R2256_U53, P2_R2256_U54);
  nand ginst10903 (P2_R2256_U21, P2_R2256_U69, P2_R2256_U70);
  nand ginst10904 (P2_R2256_U22, P2_R2256_U62, P2_R2256_U63);
  and ginst10905 (P2_R2256_U23, P2_U3622, P2_U3623);
  nand ginst10906 (P2_R2256_U24, P2_R2256_U43, P2_U3623);
  nand ginst10907 (P2_R2256_U25, P2_R2256_U38, P2_R2256_U39);
  and ginst10908 (P2_R2256_U26, P2_R2256_U55, P2_R2256_U56);
  and ginst10909 (P2_R2256_U27, P2_R2256_U57, P2_R2256_U58);
  nand ginst10910 (P2_R2256_U28, P2_R2256_U30, P2_R2256_U35);
  nand ginst10911 (P2_R2256_U29, P2_U3629, P2_U7873);
  nand ginst10912 (P2_R2256_U30, P2_U3628, P2_U3629, P2_U7873);
  and ginst10913 (P2_R2256_U31, P2_R2256_U67, P2_R2256_U68);
  not ginst10914 (P2_R2256_U32, P2_R2256_U30);
  nand ginst10915 (P2_R2256_U33, P2_U3629, P2_U7873);
  nand ginst10916 (P2_R2256_U34, P2_R2256_U33, P2_R2256_U7);
  nand ginst10917 (P2_R2256_U35, P2_R2256_U34, P2_U2616);
  not ginst10918 (P2_R2256_U36, P2_R2256_U28);
  or ginst10919 (P2_R2256_U37, P2_U3627, P2_U7873);
  nand ginst10920 (P2_R2256_U38, P2_R2256_U28, P2_R2256_U37);
  nand ginst10921 (P2_R2256_U39, P2_U3627, P2_U7873);
  nand ginst10922 (P2_R2256_U4, P2_R2256_U31, P2_R2256_U46);
  not ginst10923 (P2_R2256_U40, P2_R2256_U25);
  not ginst10924 (P2_R2256_U41, P2_R2256_U10);
  not ginst10925 (P2_R2256_U42, P2_R2256_U12);
  not ginst10926 (P2_R2256_U43, P2_R2256_U14);
  not ginst10927 (P2_R2256_U44, P2_R2256_U24);
  not ginst10928 (P2_R2256_U45, P2_R2256_U29);
  nand ginst10929 (P2_R2256_U46, P2_R2256_U66, P2_R2256_U7);
  nand ginst10930 (P2_R2256_U47, P2_R2256_U24, P2_U3622);
  nand ginst10931 (P2_R2256_U48, P2_R2256_U15, P2_R2256_U44);
  nand ginst10932 (P2_R2256_U49, P2_R2256_U14, P2_U3623);
  and ginst10933 (P2_R2256_U5, P2_R2256_U23, P2_R2256_U43);
  nand ginst10934 (P2_R2256_U50, P2_R2256_U16, P2_R2256_U43);
  nand ginst10935 (P2_R2256_U51, P2_R2256_U12, P2_U3624);
  nand ginst10936 (P2_R2256_U52, P2_R2256_U13, P2_R2256_U42);
  nand ginst10937 (P2_R2256_U53, P2_R2256_U10, P2_U3625);
  nand ginst10938 (P2_R2256_U54, P2_R2256_U11, P2_R2256_U41);
  nand ginst10939 (P2_R2256_U55, P2_R2256_U25, P2_U3626);
  nand ginst10940 (P2_R2256_U56, P2_R2256_U40, P2_R2256_U9);
  nand ginst10941 (P2_R2256_U57, P2_R2256_U8, P2_U7873);
  nand ginst10942 (P2_R2256_U58, P2_U2616, P2_U3627);
  nand ginst10943 (P2_R2256_U59, P2_R2256_U8, P2_U7873);
  not ginst10944 (P2_R2256_U6, P2_U3629);
  nand ginst10945 (P2_R2256_U60, P2_U2616, P2_U3627);
  nand ginst10946 (P2_R2256_U61, P2_R2256_U59, P2_R2256_U60);
  nand ginst10947 (P2_R2256_U62, P2_R2256_U27, P2_R2256_U28);
  nand ginst10948 (P2_R2256_U63, P2_R2256_U36, P2_R2256_U61);
  nand ginst10949 (P2_R2256_U64, P2_R2256_U29, P2_U2616);
  nand ginst10950 (P2_R2256_U65, P2_R2256_U45, P2_U7873);
  nand ginst10951 (P2_R2256_U66, P2_R2256_U64, P2_R2256_U65);
  nand ginst10952 (P2_R2256_U67, P2_R2256_U33, P2_U3628, P2_U7873);
  nand ginst10953 (P2_R2256_U68, P2_R2256_U32, P2_U2616);
  nand ginst10954 (P2_R2256_U69, P2_R2256_U6, P2_U7873);
  not ginst10955 (P2_R2256_U7, P2_U3628);
  nand ginst10956 (P2_R2256_U70, P2_U2616, P2_U3629);
  not ginst10957 (P2_R2256_U8, P2_U3627);
  not ginst10958 (P2_R2256_U9, P2_U3626);
  and ginst10959 (P2_R2267_U10, P2_R2267_U125, P2_R2267_U35);
  nand ginst10960 (P2_R2267_U100, P2_R2267_U64, P2_R2267_U89);
  nand ginst10961 (P2_R2267_U101, P2_R2267_U100, P2_U3643);
  not ginst10962 (P2_R2267_U102, P2_R2267_U31);
  not ginst10963 (P2_R2267_U103, P2_R2267_U32);
  not ginst10964 (P2_R2267_U104, P2_R2267_U33);
  not ginst10965 (P2_R2267_U105, P2_R2267_U34);
  not ginst10966 (P2_R2267_U106, P2_R2267_U35);
  not ginst10967 (P2_R2267_U107, P2_R2267_U36);
  not ginst10968 (P2_R2267_U108, P2_R2267_U37);
  not ginst10969 (P2_R2267_U109, P2_R2267_U38);
  and ginst10970 (P2_R2267_U11, P2_R2267_U123, P2_R2267_U36);
  not ginst10971 (P2_R2267_U110, P2_R2267_U39);
  not ginst10972 (P2_R2267_U111, P2_R2267_U40);
  not ginst10973 (P2_R2267_U112, P2_R2267_U62);
  nand ginst10974 (P2_R2267_U113, P2_R2267_U40, P2_U2767);
  nand ginst10975 (P2_R2267_U114, P2_R2267_U110, P2_R2267_U66);
  nand ginst10976 (P2_R2267_U115, P2_R2267_U114, P2_U2768);
  nand ginst10977 (P2_R2267_U116, P2_R2267_U109, P2_R2267_U68);
  nand ginst10978 (P2_R2267_U117, P2_R2267_U116, P2_U2770);
  nand ginst10979 (P2_R2267_U118, P2_R2267_U108, P2_R2267_U70);
  nand ginst10980 (P2_R2267_U119, P2_R2267_U118, P2_U2772);
  and ginst10981 (P2_R2267_U12, P2_R2267_U121, P2_R2267_U37);
  nand ginst10982 (P2_R2267_U120, P2_R2267_U107, P2_R2267_U72);
  nand ginst10983 (P2_R2267_U121, P2_R2267_U120, P2_U2774);
  nand ginst10984 (P2_R2267_U122, P2_R2267_U106, P2_R2267_U74);
  nand ginst10985 (P2_R2267_U123, P2_R2267_U122, P2_U2776);
  nand ginst10986 (P2_R2267_U124, P2_R2267_U105, P2_R2267_U78);
  nand ginst10987 (P2_R2267_U125, P2_R2267_U124, P2_U2778);
  nand ginst10988 (P2_R2267_U126, P2_R2267_U104, P2_R2267_U80);
  nand ginst10989 (P2_R2267_U127, P2_R2267_U126, P2_U2780);
  nand ginst10990 (P2_R2267_U128, P2_R2267_U103, P2_R2267_U82);
  nand ginst10991 (P2_R2267_U129, P2_R2267_U128, P2_U2782);
  and ginst10992 (P2_R2267_U13, P2_R2267_U119, P2_R2267_U38);
  nand ginst10993 (P2_R2267_U130, P2_R2267_U102, P2_R2267_U84);
  nand ginst10994 (P2_R2267_U131, P2_R2267_U130, P2_U2784);
  nand ginst10995 (P2_R2267_U132, P2_R2267_U86, P2_R2267_U93);
  nand ginst10996 (P2_R2267_U133, P2_R2267_U132, P2_U2786);
  nand ginst10997 (P2_R2267_U134, P2_R2267_U22, P2_U2617);
  nand ginst10998 (P2_R2267_U135, P2_R2267_U26, P2_U2789);
  nand ginst10999 (P2_R2267_U136, P2_R2267_U55, P2_R2267_U92);
  nand ginst11000 (P2_R2267_U137, P2_R2267_U25, P2_U3640);
  nand ginst11001 (P2_R2267_U138, P2_R2267_U57, P2_R2267_U91);
  nand ginst11002 (P2_R2267_U139, P2_R2267_U24, P2_U3642);
  and ginst11003 (P2_R2267_U14, P2_R2267_U117, P2_R2267_U39);
  nand ginst11004 (P2_R2267_U140, P2_R2267_U59, P2_R2267_U90);
  nand ginst11005 (P2_R2267_U141, P2_R2267_U62, P2_U2766);
  nand ginst11006 (P2_R2267_U142, P2_R2267_U112, P2_R2267_U61);
  nand ginst11007 (P2_R2267_U143, P2_R2267_U23, P2_U3644);
  nand ginst11008 (P2_R2267_U144, P2_R2267_U64, P2_R2267_U89);
  nand ginst11009 (P2_R2267_U145, P2_R2267_U39, P2_U2769);
  nand ginst11010 (P2_R2267_U146, P2_R2267_U110, P2_R2267_U66);
  nand ginst11011 (P2_R2267_U147, P2_R2267_U38, P2_U2771);
  nand ginst11012 (P2_R2267_U148, P2_R2267_U109, P2_R2267_U68);
  nand ginst11013 (P2_R2267_U149, P2_R2267_U37, P2_U2773);
  and ginst11014 (P2_R2267_U15, P2_R2267_U115, P2_R2267_U40);
  nand ginst11015 (P2_R2267_U150, P2_R2267_U108, P2_R2267_U70);
  nand ginst11016 (P2_R2267_U151, P2_R2267_U36, P2_U2775);
  nand ginst11017 (P2_R2267_U152, P2_R2267_U107, P2_R2267_U72);
  nand ginst11018 (P2_R2267_U153, P2_R2267_U35, P2_U2777);
  nand ginst11019 (P2_R2267_U154, P2_R2267_U106, P2_R2267_U74);
  nand ginst11020 (P2_R2267_U155, P2_R2267_U77, P2_U3645);
  nand ginst11021 (P2_R2267_U156, P2_R2267_U76, P2_R2267_U88);
  nand ginst11022 (P2_R2267_U157, P2_R2267_U34, P2_U2779);
  nand ginst11023 (P2_R2267_U158, P2_R2267_U105, P2_R2267_U78);
  nand ginst11024 (P2_R2267_U159, P2_R2267_U33, P2_U2781);
  and ginst11025 (P2_R2267_U16, P2_R2267_U113, P2_R2267_U62);
  nand ginst11026 (P2_R2267_U160, P2_R2267_U104, P2_R2267_U80);
  nand ginst11027 (P2_R2267_U161, P2_R2267_U32, P2_U2783);
  nand ginst11028 (P2_R2267_U162, P2_R2267_U103, P2_R2267_U82);
  nand ginst11029 (P2_R2267_U163, P2_R2267_U31, P2_U2785);
  nand ginst11030 (P2_R2267_U164, P2_R2267_U102, P2_R2267_U84);
  nand ginst11031 (P2_R2267_U165, P2_R2267_U30, P2_U2787);
  nand ginst11032 (P2_R2267_U166, P2_R2267_U86, P2_R2267_U93);
  and ginst11033 (P2_R2267_U17, P2_R2267_U101, P2_R2267_U24);
  and ginst11034 (P2_R2267_U18, P2_R2267_U25, P2_R2267_U99);
  and ginst11035 (P2_R2267_U19, P2_R2267_U26, P2_R2267_U97);
  and ginst11036 (P2_R2267_U20, P2_R2267_U30, P2_R2267_U95);
  nand ginst11037 (P2_R2267_U21, P2_R2267_U134, P2_R2267_U77);
  not ginst11038 (P2_R2267_U22, P2_U3646);
  nand ginst11039 (P2_R2267_U23, P2_R2267_U76, P2_R2267_U77);
  nand ginst11040 (P2_R2267_U24, P2_R2267_U29, P2_R2267_U64, P2_R2267_U89);
  nand ginst11041 (P2_R2267_U25, P2_R2267_U28, P2_R2267_U59, P2_R2267_U90);
  nand ginst11042 (P2_R2267_U26, P2_R2267_U27, P2_R2267_U57, P2_R2267_U91);
  not ginst11043 (P2_R2267_U27, P2_U3639);
  not ginst11044 (P2_R2267_U28, P2_U3641);
  not ginst11045 (P2_R2267_U29, P2_U3643);
  nand ginst11046 (P2_R2267_U30, P2_R2267_U44, P2_R2267_U92);
  nand ginst11047 (P2_R2267_U31, P2_R2267_U45, P2_R2267_U93);
  nand ginst11048 (P2_R2267_U32, P2_R2267_U102, P2_R2267_U46);
  nand ginst11049 (P2_R2267_U33, P2_R2267_U103, P2_R2267_U47);
  nand ginst11050 (P2_R2267_U34, P2_R2267_U104, P2_R2267_U48);
  nand ginst11051 (P2_R2267_U35, P2_R2267_U105, P2_R2267_U49);
  nand ginst11052 (P2_R2267_U36, P2_R2267_U106, P2_R2267_U50);
  nand ginst11053 (P2_R2267_U37, P2_R2267_U107, P2_R2267_U51);
  nand ginst11054 (P2_R2267_U38, P2_R2267_U108, P2_R2267_U52);
  nand ginst11055 (P2_R2267_U39, P2_R2267_U109, P2_R2267_U53);
  nand ginst11056 (P2_R2267_U40, P2_R2267_U110, P2_R2267_U54);
  not ginst11057 (P2_R2267_U41, P2_U2767);
  not ginst11058 (P2_R2267_U42, P2_U2617);
  nand ginst11059 (P2_R2267_U43, P2_R2267_U155, P2_R2267_U156);
  nor ginst11060 (P2_R2267_U44, P2_U2788, P2_U2789);
  nor ginst11061 (P2_R2267_U45, P2_U2786, P2_U2787);
  nor ginst11062 (P2_R2267_U46, P2_U2784, P2_U2785);
  nor ginst11063 (P2_R2267_U47, P2_U2782, P2_U2783);
  nor ginst11064 (P2_R2267_U48, P2_U2780, P2_U2781);
  nor ginst11065 (P2_R2267_U49, P2_U2778, P2_U2779);
  nor ginst11066 (P2_R2267_U50, P2_U2776, P2_U2777);
  nor ginst11067 (P2_R2267_U51, P2_U2774, P2_U2775);
  nor ginst11068 (P2_R2267_U52, P2_U2772, P2_U2773);
  nor ginst11069 (P2_R2267_U53, P2_U2770, P2_U2771);
  nor ginst11070 (P2_R2267_U54, P2_U2768, P2_U2769);
  not ginst11071 (P2_R2267_U55, P2_U2789);
  and ginst11072 (P2_R2267_U56, P2_R2267_U135, P2_R2267_U136);
  not ginst11073 (P2_R2267_U57, P2_U3640);
  and ginst11074 (P2_R2267_U58, P2_R2267_U137, P2_R2267_U138);
  not ginst11075 (P2_R2267_U59, P2_U3642);
  and ginst11076 (P2_R2267_U6, P2_R2267_U133, P2_R2267_U31);
  and ginst11077 (P2_R2267_U60, P2_R2267_U139, P2_R2267_U140);
  not ginst11078 (P2_R2267_U61, P2_U2766);
  nand ginst11079 (P2_R2267_U62, P2_R2267_U111, P2_R2267_U41);
  and ginst11080 (P2_R2267_U63, P2_R2267_U141, P2_R2267_U142);
  not ginst11081 (P2_R2267_U64, P2_U3644);
  and ginst11082 (P2_R2267_U65, P2_R2267_U143, P2_R2267_U144);
  not ginst11083 (P2_R2267_U66, P2_U2769);
  and ginst11084 (P2_R2267_U67, P2_R2267_U145, P2_R2267_U146);
  not ginst11085 (P2_R2267_U68, P2_U2771);
  and ginst11086 (P2_R2267_U69, P2_R2267_U147, P2_R2267_U148);
  and ginst11087 (P2_R2267_U7, P2_R2267_U131, P2_R2267_U32);
  not ginst11088 (P2_R2267_U70, P2_U2773);
  and ginst11089 (P2_R2267_U71, P2_R2267_U149, P2_R2267_U150);
  not ginst11090 (P2_R2267_U72, P2_U2775);
  and ginst11091 (P2_R2267_U73, P2_R2267_U151, P2_R2267_U152);
  not ginst11092 (P2_R2267_U74, P2_U2777);
  and ginst11093 (P2_R2267_U75, P2_R2267_U153, P2_R2267_U154);
  not ginst11094 (P2_R2267_U76, P2_U3645);
  nand ginst11095 (P2_R2267_U77, P2_R2267_U42, P2_U3646);
  not ginst11096 (P2_R2267_U78, P2_U2779);
  and ginst11097 (P2_R2267_U79, P2_R2267_U157, P2_R2267_U158);
  and ginst11098 (P2_R2267_U8, P2_R2267_U129, P2_R2267_U33);
  not ginst11099 (P2_R2267_U80, P2_U2781);
  and ginst11100 (P2_R2267_U81, P2_R2267_U159, P2_R2267_U160);
  not ginst11101 (P2_R2267_U82, P2_U2783);
  and ginst11102 (P2_R2267_U83, P2_R2267_U161, P2_R2267_U162);
  not ginst11103 (P2_R2267_U84, P2_U2785);
  and ginst11104 (P2_R2267_U85, P2_R2267_U163, P2_R2267_U164);
  not ginst11105 (P2_R2267_U86, P2_U2787);
  and ginst11106 (P2_R2267_U87, P2_R2267_U165, P2_R2267_U166);
  not ginst11107 (P2_R2267_U88, P2_R2267_U77);
  not ginst11108 (P2_R2267_U89, P2_R2267_U23);
  and ginst11109 (P2_R2267_U9, P2_R2267_U127, P2_R2267_U34);
  not ginst11110 (P2_R2267_U90, P2_R2267_U24);
  not ginst11111 (P2_R2267_U91, P2_R2267_U25);
  not ginst11112 (P2_R2267_U92, P2_R2267_U26);
  not ginst11113 (P2_R2267_U93, P2_R2267_U30);
  nand ginst11114 (P2_R2267_U94, P2_R2267_U55, P2_R2267_U92);
  nand ginst11115 (P2_R2267_U95, P2_R2267_U94, P2_U2788);
  nand ginst11116 (P2_R2267_U96, P2_R2267_U57, P2_R2267_U91);
  nand ginst11117 (P2_R2267_U97, P2_R2267_U96, P2_U3639);
  nand ginst11118 (P2_R2267_U98, P2_R2267_U59, P2_R2267_U90);
  nand ginst11119 (P2_R2267_U99, P2_R2267_U98, P2_U3641);
  not ginst11120 (P2_R2278_U10, P2_INSTADDRPOINTER_REG_5__SCAN_IN);
  nand ginst11121 (P2_R2278_U100, P2_R2278_U470, P2_R2278_U471);
  nand ginst11122 (P2_R2278_U101, P2_R2278_U477, P2_R2278_U478);
  nand ginst11123 (P2_R2278_U102, P2_R2278_U484, P2_R2278_U485);
  nand ginst11124 (P2_R2278_U103, P2_R2278_U496, P2_R2278_U497);
  nand ginst11125 (P2_R2278_U104, P2_R2278_U503, P2_R2278_U504);
  nand ginst11126 (P2_R2278_U105, P2_R2278_U510, P2_R2278_U511);
  nand ginst11127 (P2_R2278_U106, P2_R2278_U517, P2_R2278_U518);
  nand ginst11128 (P2_R2278_U107, P2_R2278_U524, P2_R2278_U525);
  nand ginst11129 (P2_R2278_U108, P2_R2278_U531, P2_R2278_U532);
  nand ginst11130 (P2_R2278_U109, P2_R2278_U538, P2_R2278_U539);
  not ginst11131 (P2_R2278_U11, P2_U3635);
  nand ginst11132 (P2_R2278_U110, P2_R2278_U545, P2_R2278_U546);
  nand ginst11133 (P2_R2278_U111, P2_R2278_U552, P2_R2278_U553);
  nand ginst11134 (P2_R2278_U112, P2_R2278_U559, P2_R2278_U560);
  and ginst11135 (P2_R2278_U113, P2_R2278_U210, P2_R2278_U314);
  and ginst11136 (P2_R2278_U114, P2_R2278_U215, P2_R2278_U313);
  and ginst11137 (P2_R2278_U115, P2_R2278_U217, P2_R2278_U221);
  and ginst11138 (P2_R2278_U116, P2_R2278_U222, P2_R2278_U316);
  and ginst11139 (P2_R2278_U117, P2_R2278_U224, P2_R2278_U228);
  and ginst11140 (P2_R2278_U118, P2_R2278_U229, P2_R2278_U318);
  and ginst11141 (P2_R2278_U119, P2_R2278_U231, P2_R2278_U235);
  not ginst11142 (P2_R2278_U12, P2_INSTADDRPOINTER_REG_3__SCAN_IN);
  and ginst11143 (P2_R2278_U120, P2_R2278_U236, P2_R2278_U320);
  and ginst11144 (P2_R2278_U121, P2_R2278_U238, P2_R2278_U242);
  and ginst11145 (P2_R2278_U122, P2_R2278_U243, P2_R2278_U322);
  and ginst11146 (P2_R2278_U123, P2_R2278_U245, P2_R2278_U249);
  and ginst11147 (P2_R2278_U124, P2_R2278_U250, P2_R2278_U324);
  and ginst11148 (P2_R2278_U125, P2_R2278_U252, P2_R2278_U256);
  and ginst11149 (P2_R2278_U126, P2_R2278_U257, P2_R2278_U326);
  and ginst11150 (P2_R2278_U127, P2_R2278_U259, P2_R2278_U263);
  and ginst11151 (P2_R2278_U128, P2_R2278_U264, P2_R2278_U328);
  and ginst11152 (P2_R2278_U129, P2_R2278_U270, P2_R2278_U273);
  not ginst11153 (P2_R2278_U13, P2_U3638);
  and ginst11154 (P2_R2278_U130, P2_R2278_U273, P2_R2278_U331);
  and ginst11155 (P2_R2278_U131, P2_R2278_U274, P2_R2278_U334);
  and ginst11156 (P2_R2278_U132, P2_R2278_U276, P2_R2278_U280);
  and ginst11157 (P2_R2278_U133, P2_R2278_U281, P2_R2278_U336);
  and ginst11158 (P2_R2278_U134, P2_R2278_U283, P2_R2278_U287);
  and ginst11159 (P2_R2278_U135, P2_R2278_U288, P2_R2278_U338);
  and ginst11160 (P2_R2278_U136, P2_R2278_U292, P2_R2278_U296, P2_R2278_U299);
  and ginst11161 (P2_R2278_U137, P2_R2278_U300, P2_R2278_U304);
  and ginst11162 (P2_R2278_U138, P2_R2278_U302, P2_R2278_U307);
  and ginst11163 (P2_R2278_U139, P2_R2278_U138, P2_R2278_U397);
  not ginst11164 (P2_R2278_U14, P2_INSTADDRPOINTER_REG_0__SCAN_IN);
  and ginst11165 (P2_R2278_U140, P2_R2278_U300, P2_R2278_U343);
  and ginst11166 (P2_R2278_U141, P2_R2278_U142, P2_R2278_U4);
  and ginst11167 (P2_R2278_U142, P2_R2278_U304, P2_R2278_U306);
  and ginst11168 (P2_R2278_U143, P2_R2278_U292, P2_R2278_U296);
  and ginst11169 (P2_R2278_U144, P2_R2278_U266, P2_R2278_U270);
  and ginst11170 (P2_R2278_U145, P2_R2278_U346, P2_R2278_U347);
  nand ginst11171 (P2_R2278_U146, P2_R2278_U232, P2_R2278_U49);
  and ginst11172 (P2_R2278_U147, P2_R2278_U353, P2_R2278_U354);
  nand ginst11173 (P2_R2278_U148, P2_R2278_U118, P2_R2278_U317);
  and ginst11174 (P2_R2278_U149, P2_R2278_U360, P2_R2278_U361);
  nand ginst11175 (P2_R2278_U15, P2_INSTADDRPOINTER_REG_0__SCAN_IN, P2_U3638);
  nand ginst11176 (P2_R2278_U150, P2_R2278_U225, P2_R2278_U26);
  and ginst11177 (P2_R2278_U151, P2_R2278_U367, P2_R2278_U368);
  nand ginst11178 (P2_R2278_U152, P2_R2278_U116, P2_R2278_U315);
  and ginst11179 (P2_R2278_U153, P2_R2278_U374, P2_R2278_U375);
  nand ginst11180 (P2_R2278_U154, P2_R2278_U218, P2_R2278_U23);
  and ginst11181 (P2_R2278_U155, P2_R2278_U381, P2_R2278_U382);
  nand ginst11182 (P2_R2278_U156, P2_R2278_U114, P2_R2278_U312);
  and ginst11183 (P2_R2278_U157, P2_R2278_U388, P2_R2278_U389);
  nand ginst11184 (P2_R2278_U158, P2_R2278_U20, P2_R2278_U211);
  not ginst11185 (P2_R2278_U159, P2_INSTADDRPOINTER_REG_31__SCAN_IN);
  not ginst11186 (P2_R2278_U16, P2_U3637);
  not ginst11187 (P2_R2278_U160, P2_U2790);
  and ginst11188 (P2_R2278_U161, P2_R2278_U400, P2_R2278_U401);
  and ginst11189 (P2_R2278_U162, P2_R2278_U402, P2_R2278_U403);
  nand ginst11190 (P2_R2278_U163, P2_R2278_U303, P2_R2278_U304);
  and ginst11191 (P2_R2278_U164, P2_R2278_U409, P2_R2278_U410);
  nand ginst11192 (P2_R2278_U165, P2_R2278_U310, P2_R2278_U311, P2_R2278_U82);
  and ginst11193 (P2_R2278_U166, P2_R2278_U416, P2_R2278_U417);
  nand ginst11194 (P2_R2278_U167, P2_R2278_U140, P2_R2278_U342);
  and ginst11195 (P2_R2278_U168, P2_R2278_U423, P2_R2278_U424);
  nand ginst11196 (P2_R2278_U169, P2_R2278_U339, P2_R2278_U341);
  not ginst11197 (P2_R2278_U17, P2_INSTADDRPOINTER_REG_1__SCAN_IN);
  and ginst11198 (P2_R2278_U170, P2_R2278_U430, P2_R2278_U431);
  nand ginst11199 (P2_R2278_U171, P2_R2278_U293, P2_R2278_U78);
  and ginst11200 (P2_R2278_U172, P2_R2278_U437, P2_R2278_U438);
  nand ginst11201 (P2_R2278_U173, P2_R2278_U205, P2_R2278_U290, P2_R2278_U308);
  nand ginst11202 (P2_R2278_U174, P2_R2278_U135, P2_R2278_U337);
  and ginst11203 (P2_R2278_U175, P2_R2278_U451, P2_R2278_U452);
  nand ginst11204 (P2_R2278_U176, P2_R2278_U284, P2_R2278_U71);
  and ginst11205 (P2_R2278_U177, P2_R2278_U458, P2_R2278_U459);
  nand ginst11206 (P2_R2278_U178, P2_R2278_U133, P2_R2278_U335);
  and ginst11207 (P2_R2278_U179, P2_R2278_U465, P2_R2278_U466);
  not ginst11208 (P2_R2278_U18, P2_U3636);
  nand ginst11209 (P2_R2278_U180, P2_R2278_U277, P2_R2278_U68);
  and ginst11210 (P2_R2278_U181, P2_R2278_U472, P2_R2278_U473);
  nand ginst11211 (P2_R2278_U182, P2_R2278_U131, P2_R2278_U333);
  and ginst11212 (P2_R2278_U183, P2_R2278_U479, P2_R2278_U480);
  nand ginst11213 (P2_R2278_U184, P2_R2278_U329, P2_R2278_U330);
  and ginst11214 (P2_R2278_U185, P2_R2278_U491, P2_R2278_U492);
  nand ginst11215 (P2_R2278_U186, P2_R2278_U267, P2_R2278_U268);
  and ginst11216 (P2_R2278_U187, P2_R2278_U498, P2_R2278_U499);
  nand ginst11217 (P2_R2278_U188, P2_R2278_U128, P2_R2278_U327);
  and ginst11218 (P2_R2278_U189, P2_R2278_U505, P2_R2278_U506);
  not ginst11219 (P2_R2278_U19, P2_INSTADDRPOINTER_REG_2__SCAN_IN);
  nand ginst11220 (P2_R2278_U190, P2_R2278_U260, P2_R2278_U61);
  and ginst11221 (P2_R2278_U191, P2_R2278_U512, P2_R2278_U513);
  nand ginst11222 (P2_R2278_U192, P2_R2278_U126, P2_R2278_U325);
  and ginst11223 (P2_R2278_U193, P2_R2278_U519, P2_R2278_U520);
  nand ginst11224 (P2_R2278_U194, P2_R2278_U253, P2_R2278_U58);
  and ginst11225 (P2_R2278_U195, P2_R2278_U526, P2_R2278_U527);
  nand ginst11226 (P2_R2278_U196, P2_R2278_U124, P2_R2278_U323);
  and ginst11227 (P2_R2278_U197, P2_R2278_U533, P2_R2278_U534);
  nand ginst11228 (P2_R2278_U198, P2_R2278_U246, P2_R2278_U55);
  and ginst11229 (P2_R2278_U199, P2_R2278_U540, P2_R2278_U541);
  nand ginst11230 (P2_R2278_U20, P2_INSTADDRPOINTER_REG_2__SCAN_IN, P2_U3636);
  nand ginst11231 (P2_R2278_U200, P2_R2278_U122, P2_R2278_U321);
  and ginst11232 (P2_R2278_U201, P2_R2278_U547, P2_R2278_U548);
  nand ginst11233 (P2_R2278_U202, P2_R2278_U239, P2_R2278_U52);
  and ginst11234 (P2_R2278_U203, P2_R2278_U554, P2_R2278_U555);
  nand ginst11235 (P2_R2278_U204, P2_R2278_U120, P2_R2278_U319);
  nand ginst11236 (P2_R2278_U205, P2_R2278_U174, P2_U2796);
  nand ginst11237 (P2_R2278_U206, P2_R2278_U139, P2_R2278_U344);
  not ginst11238 (P2_R2278_U207, P2_R2278_U82);
  not ginst11239 (P2_R2278_U208, P2_R2278_U15);
  not ginst11240 (P2_R2278_U209, P2_R2278_U165);
  not ginst11241 (P2_R2278_U21, P2_U3634);
  or ginst11242 (P2_R2278_U210, P2_INSTADDRPOINTER_REG_2__SCAN_IN, P2_U3636);
  nand ginst11243 (P2_R2278_U211, P2_R2278_U165, P2_R2278_U210);
  not ginst11244 (P2_R2278_U212, P2_R2278_U20);
  not ginst11245 (P2_R2278_U213, P2_R2278_U158);
  or ginst11246 (P2_R2278_U214, P2_INSTADDRPOINTER_REG_3__SCAN_IN, P2_U3635);
  nand ginst11247 (P2_R2278_U215, P2_INSTADDRPOINTER_REG_3__SCAN_IN, P2_U3635);
  not ginst11248 (P2_R2278_U216, P2_R2278_U156);
  or ginst11249 (P2_R2278_U217, P2_INSTADDRPOINTER_REG_4__SCAN_IN, P2_U3634);
  nand ginst11250 (P2_R2278_U218, P2_R2278_U156, P2_R2278_U217);
  not ginst11251 (P2_R2278_U219, P2_R2278_U23);
  not ginst11252 (P2_R2278_U22, P2_INSTADDRPOINTER_REG_4__SCAN_IN);
  not ginst11253 (P2_R2278_U220, P2_R2278_U154);
  or ginst11254 (P2_R2278_U221, P2_INSTADDRPOINTER_REG_5__SCAN_IN, P2_U3633);
  nand ginst11255 (P2_R2278_U222, P2_INSTADDRPOINTER_REG_5__SCAN_IN, P2_U3633);
  not ginst11256 (P2_R2278_U223, P2_R2278_U152);
  or ginst11257 (P2_R2278_U224, P2_INSTADDRPOINTER_REG_6__SCAN_IN, P2_U3632);
  nand ginst11258 (P2_R2278_U225, P2_R2278_U152, P2_R2278_U224);
  not ginst11259 (P2_R2278_U226, P2_R2278_U26);
  not ginst11260 (P2_R2278_U227, P2_R2278_U150);
  or ginst11261 (P2_R2278_U228, P2_INSTADDRPOINTER_REG_7__SCAN_IN, P2_U3631);
  nand ginst11262 (P2_R2278_U229, P2_INSTADDRPOINTER_REG_7__SCAN_IN, P2_U3631);
  nand ginst11263 (P2_R2278_U23, P2_INSTADDRPOINTER_REG_4__SCAN_IN, P2_U3634);
  not ginst11264 (P2_R2278_U230, P2_R2278_U148);
  or ginst11265 (P2_R2278_U231, P2_INSTADDRPOINTER_REG_8__SCAN_IN, P2_U3630);
  nand ginst11266 (P2_R2278_U232, P2_R2278_U148, P2_R2278_U231);
  not ginst11267 (P2_R2278_U233, P2_R2278_U49);
  not ginst11268 (P2_R2278_U234, P2_R2278_U146);
  or ginst11269 (P2_R2278_U235, P2_INSTADDRPOINTER_REG_9__SCAN_IN, P2_U2812);
  nand ginst11270 (P2_R2278_U236, P2_INSTADDRPOINTER_REG_9__SCAN_IN, P2_U2812);
  not ginst11271 (P2_R2278_U237, P2_R2278_U204);
  or ginst11272 (P2_R2278_U238, P2_INSTADDRPOINTER_REG_10__SCAN_IN, P2_U2811);
  nand ginst11273 (P2_R2278_U239, P2_R2278_U204, P2_R2278_U238);
  not ginst11274 (P2_R2278_U24, P2_U3632);
  not ginst11275 (P2_R2278_U240, P2_R2278_U52);
  not ginst11276 (P2_R2278_U241, P2_R2278_U202);
  or ginst11277 (P2_R2278_U242, P2_INSTADDRPOINTER_REG_11__SCAN_IN, P2_U2810);
  nand ginst11278 (P2_R2278_U243, P2_INSTADDRPOINTER_REG_11__SCAN_IN, P2_U2810);
  not ginst11279 (P2_R2278_U244, P2_R2278_U200);
  or ginst11280 (P2_R2278_U245, P2_INSTADDRPOINTER_REG_12__SCAN_IN, P2_U2809);
  nand ginst11281 (P2_R2278_U246, P2_R2278_U200, P2_R2278_U245);
  not ginst11282 (P2_R2278_U247, P2_R2278_U55);
  not ginst11283 (P2_R2278_U248, P2_R2278_U198);
  or ginst11284 (P2_R2278_U249, P2_INSTADDRPOINTER_REG_13__SCAN_IN, P2_U2808);
  not ginst11285 (P2_R2278_U25, P2_INSTADDRPOINTER_REG_6__SCAN_IN);
  nand ginst11286 (P2_R2278_U250, P2_INSTADDRPOINTER_REG_13__SCAN_IN, P2_U2808);
  not ginst11287 (P2_R2278_U251, P2_R2278_U196);
  or ginst11288 (P2_R2278_U252, P2_INSTADDRPOINTER_REG_14__SCAN_IN, P2_U2807);
  nand ginst11289 (P2_R2278_U253, P2_R2278_U196, P2_R2278_U252);
  not ginst11290 (P2_R2278_U254, P2_R2278_U58);
  not ginst11291 (P2_R2278_U255, P2_R2278_U194);
  or ginst11292 (P2_R2278_U256, P2_INSTADDRPOINTER_REG_15__SCAN_IN, P2_U2806);
  nand ginst11293 (P2_R2278_U257, P2_INSTADDRPOINTER_REG_15__SCAN_IN, P2_U2806);
  not ginst11294 (P2_R2278_U258, P2_R2278_U192);
  or ginst11295 (P2_R2278_U259, P2_INSTADDRPOINTER_REG_16__SCAN_IN, P2_U2805);
  nand ginst11296 (P2_R2278_U26, P2_INSTADDRPOINTER_REG_6__SCAN_IN, P2_U3632);
  nand ginst11297 (P2_R2278_U260, P2_R2278_U192, P2_R2278_U259);
  not ginst11298 (P2_R2278_U261, P2_R2278_U61);
  not ginst11299 (P2_R2278_U262, P2_R2278_U190);
  or ginst11300 (P2_R2278_U263, P2_INSTADDRPOINTER_REG_17__SCAN_IN, P2_U2804);
  nand ginst11301 (P2_R2278_U264, P2_INSTADDRPOINTER_REG_17__SCAN_IN, P2_U2804);
  not ginst11302 (P2_R2278_U265, P2_R2278_U188);
  or ginst11303 (P2_R2278_U266, P2_INSTADDRPOINTER_REG_18__SCAN_IN, P2_U2803);
  nand ginst11304 (P2_R2278_U267, P2_R2278_U188, P2_R2278_U266);
  nand ginst11305 (P2_R2278_U268, P2_INSTADDRPOINTER_REG_18__SCAN_IN, P2_U2803);
  not ginst11306 (P2_R2278_U269, P2_R2278_U186);
  not ginst11307 (P2_R2278_U27, P2_U3630);
  or ginst11308 (P2_R2278_U270, P2_INSTADDRPOINTER_REG_19__SCAN_IN, P2_U2802);
  nand ginst11309 (P2_R2278_U271, P2_INSTADDRPOINTER_REG_19__SCAN_IN, P2_U2802);
  not ginst11310 (P2_R2278_U272, P2_R2278_U184);
  or ginst11311 (P2_R2278_U273, P2_INSTADDRPOINTER_REG_20__SCAN_IN, P2_U2801);
  nand ginst11312 (P2_R2278_U274, P2_INSTADDRPOINTER_REG_20__SCAN_IN, P2_U2801);
  not ginst11313 (P2_R2278_U275, P2_R2278_U182);
  or ginst11314 (P2_R2278_U276, P2_INSTADDRPOINTER_REG_21__SCAN_IN, P2_U2800);
  nand ginst11315 (P2_R2278_U277, P2_R2278_U182, P2_R2278_U276);
  not ginst11316 (P2_R2278_U278, P2_R2278_U68);
  not ginst11317 (P2_R2278_U279, P2_R2278_U180);
  not ginst11318 (P2_R2278_U28, P2_INSTADDRPOINTER_REG_8__SCAN_IN);
  or ginst11319 (P2_R2278_U280, P2_INSTADDRPOINTER_REG_22__SCAN_IN, P2_U2799);
  nand ginst11320 (P2_R2278_U281, P2_INSTADDRPOINTER_REG_22__SCAN_IN, P2_U2799);
  not ginst11321 (P2_R2278_U282, P2_R2278_U178);
  or ginst11322 (P2_R2278_U283, P2_INSTADDRPOINTER_REG_23__SCAN_IN, P2_U2798);
  nand ginst11323 (P2_R2278_U284, P2_R2278_U178, P2_R2278_U283);
  not ginst11324 (P2_R2278_U285, P2_R2278_U71);
  not ginst11325 (P2_R2278_U286, P2_R2278_U176);
  or ginst11326 (P2_R2278_U287, P2_INSTADDRPOINTER_REG_24__SCAN_IN, P2_U2797);
  nand ginst11327 (P2_R2278_U288, P2_INSTADDRPOINTER_REG_24__SCAN_IN, P2_U2797);
  not ginst11328 (P2_R2278_U289, P2_R2278_U174);
  not ginst11329 (P2_R2278_U29, P2_INSTADDRPOINTER_REG_9__SCAN_IN);
  nand ginst11330 (P2_R2278_U290, P2_INSTADDRPOINTER_REG_25__SCAN_IN, P2_R2278_U174);
  not ginst11331 (P2_R2278_U291, P2_R2278_U173);
  or ginst11332 (P2_R2278_U292, P2_INSTADDRPOINTER_REG_26__SCAN_IN, P2_U2795);
  nand ginst11333 (P2_R2278_U293, P2_R2278_U173, P2_R2278_U292);
  not ginst11334 (P2_R2278_U294, P2_R2278_U78);
  not ginst11335 (P2_R2278_U295, P2_R2278_U171);
  or ginst11336 (P2_R2278_U296, P2_INSTADDRPOINTER_REG_27__SCAN_IN, P2_U2794);
  nand ginst11337 (P2_R2278_U297, P2_INSTADDRPOINTER_REG_27__SCAN_IN, P2_U2794);
  not ginst11338 (P2_R2278_U298, P2_R2278_U169);
  or ginst11339 (P2_R2278_U299, P2_INSTADDRPOINTER_REG_28__SCAN_IN, P2_U2793);
  not ginst11340 (P2_R2278_U30, P2_U2812);
  nand ginst11341 (P2_R2278_U300, P2_INSTADDRPOINTER_REG_28__SCAN_IN, P2_U2793);
  not ginst11342 (P2_R2278_U301, P2_R2278_U167);
  or ginst11343 (P2_R2278_U302, P2_INSTADDRPOINTER_REG_29__SCAN_IN, P2_U2792);
  nand ginst11344 (P2_R2278_U303, P2_R2278_U167, P2_R2278_U302);
  nand ginst11345 (P2_R2278_U304, P2_INSTADDRPOINTER_REG_29__SCAN_IN, P2_U2792);
  not ginst11346 (P2_R2278_U305, P2_R2278_U163);
  nand ginst11347 (P2_R2278_U306, P2_INSTADDRPOINTER_REG_30__SCAN_IN, P2_U2791);
  or ginst11348 (P2_R2278_U307, P2_INSTADDRPOINTER_REG_30__SCAN_IN, P2_U2791);
  nand ginst11349 (P2_R2278_U308, P2_INSTADDRPOINTER_REG_25__SCAN_IN, P2_U2796);
  nand ginst11350 (P2_R2278_U309, P2_R2278_U141, P2_R2278_U303);
  not ginst11351 (P2_R2278_U31, P2_U2793);
  nand ginst11352 (P2_R2278_U310, P2_INSTADDRPOINTER_REG_1__SCAN_IN, P2_R2278_U208);
  nand ginst11353 (P2_R2278_U311, P2_INSTADDRPOINTER_REG_1__SCAN_IN, P2_U3637);
  nand ginst11354 (P2_R2278_U312, P2_R2278_U113, P2_R2278_U165);
  nand ginst11355 (P2_R2278_U313, P2_R2278_U212, P2_R2278_U214);
  or ginst11356 (P2_R2278_U314, P2_INSTADDRPOINTER_REG_3__SCAN_IN, P2_U3635);
  nand ginst11357 (P2_R2278_U315, P2_R2278_U115, P2_R2278_U156);
  nand ginst11358 (P2_R2278_U316, P2_R2278_U219, P2_R2278_U221);
  nand ginst11359 (P2_R2278_U317, P2_R2278_U117, P2_R2278_U152);
  nand ginst11360 (P2_R2278_U318, P2_R2278_U226, P2_R2278_U228);
  nand ginst11361 (P2_R2278_U319, P2_R2278_U119, P2_R2278_U148);
  not ginst11362 (P2_R2278_U32, P2_INSTADDRPOINTER_REG_28__SCAN_IN);
  nand ginst11363 (P2_R2278_U320, P2_R2278_U233, P2_R2278_U235);
  nand ginst11364 (P2_R2278_U321, P2_R2278_U121, P2_R2278_U204);
  nand ginst11365 (P2_R2278_U322, P2_R2278_U240, P2_R2278_U242);
  nand ginst11366 (P2_R2278_U323, P2_R2278_U123, P2_R2278_U200);
  nand ginst11367 (P2_R2278_U324, P2_R2278_U247, P2_R2278_U249);
  nand ginst11368 (P2_R2278_U325, P2_R2278_U125, P2_R2278_U196);
  nand ginst11369 (P2_R2278_U326, P2_R2278_U254, P2_R2278_U256);
  nand ginst11370 (P2_R2278_U327, P2_R2278_U127, P2_R2278_U192);
  nand ginst11371 (P2_R2278_U328, P2_R2278_U261, P2_R2278_U263);
  nand ginst11372 (P2_R2278_U329, P2_R2278_U144, P2_R2278_U188);
  not ginst11373 (P2_R2278_U33, P2_U2792);
  nand ginst11374 (P2_R2278_U330, P2_R2278_U331, P2_R2278_U332);
  or ginst11375 (P2_R2278_U331, P2_INSTADDRPOINTER_REG_19__SCAN_IN, P2_U2802);
  nand ginst11376 (P2_R2278_U332, P2_R2278_U268, P2_R2278_U271);
  nand ginst11377 (P2_R2278_U333, P2_R2278_U129, P2_R2278_U188, P2_R2278_U266);
  nand ginst11378 (P2_R2278_U334, P2_R2278_U130, P2_R2278_U332);
  nand ginst11379 (P2_R2278_U335, P2_R2278_U132, P2_R2278_U182);
  nand ginst11380 (P2_R2278_U336, P2_R2278_U278, P2_R2278_U280);
  nand ginst11381 (P2_R2278_U337, P2_R2278_U134, P2_R2278_U178);
  nand ginst11382 (P2_R2278_U338, P2_R2278_U285, P2_R2278_U287);
  nand ginst11383 (P2_R2278_U339, P2_R2278_U143, P2_R2278_U173);
  not ginst11384 (P2_R2278_U34, P2_INSTADDRPOINTER_REG_29__SCAN_IN);
  nand ginst11385 (P2_R2278_U340, P2_R2278_U294, P2_R2278_U296);
  not ginst11386 (P2_R2278_U341, P2_R2278_U81);
  nand ginst11387 (P2_R2278_U342, P2_R2278_U136, P2_R2278_U173);
  nand ginst11388 (P2_R2278_U343, P2_R2278_U299, P2_R2278_U81);
  nand ginst11389 (P2_R2278_U344, P2_R2278_U137, P2_R2278_U342, P2_R2278_U343);
  nand ginst11390 (P2_R2278_U345, P2_INSTADDRPOINTER_REG_1__SCAN_IN, P2_R2278_U207);
  nand ginst11391 (P2_R2278_U346, P2_INSTADDRPOINTER_REG_9__SCAN_IN, P2_R2278_U30);
  nand ginst11392 (P2_R2278_U347, P2_R2278_U29, P2_U2812);
  nand ginst11393 (P2_R2278_U348, P2_INSTADDRPOINTER_REG_9__SCAN_IN, P2_R2278_U30);
  nand ginst11394 (P2_R2278_U349, P2_R2278_U29, P2_U2812);
  not ginst11395 (P2_R2278_U35, P2_U2797);
  nand ginst11396 (P2_R2278_U350, P2_R2278_U348, P2_R2278_U349);
  nand ginst11397 (P2_R2278_U351, P2_R2278_U145, P2_R2278_U146);
  nand ginst11398 (P2_R2278_U352, P2_R2278_U234, P2_R2278_U350);
  nand ginst11399 (P2_R2278_U353, P2_INSTADDRPOINTER_REG_8__SCAN_IN, P2_R2278_U27);
  nand ginst11400 (P2_R2278_U354, P2_R2278_U28, P2_U3630);
  nand ginst11401 (P2_R2278_U355, P2_INSTADDRPOINTER_REG_8__SCAN_IN, P2_R2278_U27);
  nand ginst11402 (P2_R2278_U356, P2_R2278_U28, P2_U3630);
  nand ginst11403 (P2_R2278_U357, P2_R2278_U355, P2_R2278_U356);
  nand ginst11404 (P2_R2278_U358, P2_R2278_U147, P2_R2278_U148);
  nand ginst11405 (P2_R2278_U359, P2_R2278_U230, P2_R2278_U357);
  not ginst11406 (P2_R2278_U36, P2_INSTADDRPOINTER_REG_24__SCAN_IN);
  nand ginst11407 (P2_R2278_U360, P2_INSTADDRPOINTER_REG_7__SCAN_IN, P2_R2278_U7);
  nand ginst11408 (P2_R2278_U361, P2_R2278_U8, P2_U3631);
  nand ginst11409 (P2_R2278_U362, P2_INSTADDRPOINTER_REG_7__SCAN_IN, P2_R2278_U7);
  nand ginst11410 (P2_R2278_U363, P2_R2278_U8, P2_U3631);
  nand ginst11411 (P2_R2278_U364, P2_R2278_U362, P2_R2278_U363);
  nand ginst11412 (P2_R2278_U365, P2_R2278_U149, P2_R2278_U150);
  nand ginst11413 (P2_R2278_U366, P2_R2278_U227, P2_R2278_U364);
  nand ginst11414 (P2_R2278_U367, P2_INSTADDRPOINTER_REG_6__SCAN_IN, P2_R2278_U24);
  nand ginst11415 (P2_R2278_U368, P2_R2278_U25, P2_U3632);
  nand ginst11416 (P2_R2278_U369, P2_INSTADDRPOINTER_REG_6__SCAN_IN, P2_R2278_U24);
  not ginst11417 (P2_R2278_U37, P2_U2799);
  nand ginst11418 (P2_R2278_U370, P2_R2278_U25, P2_U3632);
  nand ginst11419 (P2_R2278_U371, P2_R2278_U369, P2_R2278_U370);
  nand ginst11420 (P2_R2278_U372, P2_R2278_U151, P2_R2278_U152);
  nand ginst11421 (P2_R2278_U373, P2_R2278_U223, P2_R2278_U371);
  nand ginst11422 (P2_R2278_U374, P2_INSTADDRPOINTER_REG_5__SCAN_IN, P2_R2278_U9);
  nand ginst11423 (P2_R2278_U375, P2_R2278_U10, P2_U3633);
  nand ginst11424 (P2_R2278_U376, P2_INSTADDRPOINTER_REG_5__SCAN_IN, P2_R2278_U9);
  nand ginst11425 (P2_R2278_U377, P2_R2278_U10, P2_U3633);
  nand ginst11426 (P2_R2278_U378, P2_R2278_U376, P2_R2278_U377);
  nand ginst11427 (P2_R2278_U379, P2_R2278_U153, P2_R2278_U154);
  not ginst11428 (P2_R2278_U38, P2_INSTADDRPOINTER_REG_22__SCAN_IN);
  nand ginst11429 (P2_R2278_U380, P2_R2278_U220, P2_R2278_U378);
  nand ginst11430 (P2_R2278_U381, P2_INSTADDRPOINTER_REG_4__SCAN_IN, P2_R2278_U21);
  nand ginst11431 (P2_R2278_U382, P2_R2278_U22, P2_U3634);
  nand ginst11432 (P2_R2278_U383, P2_INSTADDRPOINTER_REG_4__SCAN_IN, P2_R2278_U21);
  nand ginst11433 (P2_R2278_U384, P2_R2278_U22, P2_U3634);
  nand ginst11434 (P2_R2278_U385, P2_R2278_U383, P2_R2278_U384);
  nand ginst11435 (P2_R2278_U386, P2_R2278_U155, P2_R2278_U156);
  nand ginst11436 (P2_R2278_U387, P2_R2278_U216, P2_R2278_U385);
  nand ginst11437 (P2_R2278_U388, P2_INSTADDRPOINTER_REG_3__SCAN_IN, P2_R2278_U11);
  nand ginst11438 (P2_R2278_U389, P2_R2278_U12, P2_U3635);
  not ginst11439 (P2_R2278_U39, P2_U2801);
  nand ginst11440 (P2_R2278_U390, P2_INSTADDRPOINTER_REG_3__SCAN_IN, P2_R2278_U11);
  nand ginst11441 (P2_R2278_U391, P2_R2278_U12, P2_U3635);
  nand ginst11442 (P2_R2278_U392, P2_R2278_U390, P2_R2278_U391);
  nand ginst11443 (P2_R2278_U393, P2_R2278_U157, P2_R2278_U158);
  nand ginst11444 (P2_R2278_U394, P2_R2278_U213, P2_R2278_U392);
  nand ginst11445 (P2_R2278_U395, P2_INSTADDRPOINTER_REG_31__SCAN_IN, P2_R2278_U160);
  nand ginst11446 (P2_R2278_U396, P2_R2278_U159, P2_U2790);
  nand ginst11447 (P2_R2278_U397, P2_R2278_U395, P2_R2278_U396);
  nand ginst11448 (P2_R2278_U398, P2_INSTADDRPOINTER_REG_31__SCAN_IN, P2_R2278_U160);
  nand ginst11449 (P2_R2278_U399, P2_R2278_U159, P2_U2790);
  and ginst11450 (P2_R2278_U4, P2_R2278_U398, P2_R2278_U399);
  not ginst11451 (P2_R2278_U40, P2_INSTADDRPOINTER_REG_20__SCAN_IN);
  nand ginst11452 (P2_R2278_U400, P2_R2278_U4, P2_R2278_U79, P2_R2278_U80);
  nand ginst11453 (P2_R2278_U401, P2_INSTADDRPOINTER_REG_30__SCAN_IN, P2_R2278_U397, P2_U2791);
  nand ginst11454 (P2_R2278_U402, P2_INSTADDRPOINTER_REG_30__SCAN_IN, P2_R2278_U79);
  nand ginst11455 (P2_R2278_U403, P2_R2278_U80, P2_U2791);
  nand ginst11456 (P2_R2278_U404, P2_INSTADDRPOINTER_REG_30__SCAN_IN, P2_R2278_U79);
  nand ginst11457 (P2_R2278_U405, P2_R2278_U80, P2_U2791);
  nand ginst11458 (P2_R2278_U406, P2_R2278_U404, P2_R2278_U405);
  nand ginst11459 (P2_R2278_U407, P2_R2278_U162, P2_R2278_U163);
  nand ginst11460 (P2_R2278_U408, P2_R2278_U305, P2_R2278_U406);
  nand ginst11461 (P2_R2278_U409, P2_INSTADDRPOINTER_REG_2__SCAN_IN, P2_R2278_U18);
  not ginst11462 (P2_R2278_U41, P2_U2804);
  nand ginst11463 (P2_R2278_U410, P2_R2278_U19, P2_U3636);
  nand ginst11464 (P2_R2278_U411, P2_INSTADDRPOINTER_REG_2__SCAN_IN, P2_R2278_U18);
  nand ginst11465 (P2_R2278_U412, P2_R2278_U19, P2_U3636);
  nand ginst11466 (P2_R2278_U413, P2_R2278_U411, P2_R2278_U412);
  nand ginst11467 (P2_R2278_U414, P2_R2278_U164, P2_R2278_U165);
  nand ginst11468 (P2_R2278_U415, P2_R2278_U209, P2_R2278_U413);
  nand ginst11469 (P2_R2278_U416, P2_INSTADDRPOINTER_REG_29__SCAN_IN, P2_R2278_U33);
  nand ginst11470 (P2_R2278_U417, P2_R2278_U34, P2_U2792);
  nand ginst11471 (P2_R2278_U418, P2_INSTADDRPOINTER_REG_29__SCAN_IN, P2_R2278_U33);
  nand ginst11472 (P2_R2278_U419, P2_R2278_U34, P2_U2792);
  not ginst11473 (P2_R2278_U42, P2_INSTADDRPOINTER_REG_17__SCAN_IN);
  nand ginst11474 (P2_R2278_U420, P2_R2278_U418, P2_R2278_U419);
  nand ginst11475 (P2_R2278_U421, P2_R2278_U166, P2_R2278_U167);
  nand ginst11476 (P2_R2278_U422, P2_R2278_U301, P2_R2278_U420);
  nand ginst11477 (P2_R2278_U423, P2_INSTADDRPOINTER_REG_28__SCAN_IN, P2_R2278_U31);
  nand ginst11478 (P2_R2278_U424, P2_R2278_U32, P2_U2793);
  nand ginst11479 (P2_R2278_U425, P2_INSTADDRPOINTER_REG_28__SCAN_IN, P2_R2278_U31);
  nand ginst11480 (P2_R2278_U426, P2_R2278_U32, P2_U2793);
  nand ginst11481 (P2_R2278_U427, P2_R2278_U425, P2_R2278_U426);
  nand ginst11482 (P2_R2278_U428, P2_R2278_U168, P2_R2278_U169);
  nand ginst11483 (P2_R2278_U429, P2_R2278_U298, P2_R2278_U427);
  not ginst11484 (P2_R2278_U43, P2_U2806);
  nand ginst11485 (P2_R2278_U430, P2_INSTADDRPOINTER_REG_27__SCAN_IN, P2_R2278_U74);
  nand ginst11486 (P2_R2278_U431, P2_R2278_U75, P2_U2794);
  nand ginst11487 (P2_R2278_U432, P2_INSTADDRPOINTER_REG_27__SCAN_IN, P2_R2278_U74);
  nand ginst11488 (P2_R2278_U433, P2_R2278_U75, P2_U2794);
  nand ginst11489 (P2_R2278_U434, P2_R2278_U432, P2_R2278_U433);
  nand ginst11490 (P2_R2278_U435, P2_R2278_U170, P2_R2278_U171);
  nand ginst11491 (P2_R2278_U436, P2_R2278_U295, P2_R2278_U434);
  nand ginst11492 (P2_R2278_U437, P2_INSTADDRPOINTER_REG_26__SCAN_IN, P2_R2278_U76);
  nand ginst11493 (P2_R2278_U438, P2_R2278_U77, P2_U2795);
  nand ginst11494 (P2_R2278_U439, P2_INSTADDRPOINTER_REG_26__SCAN_IN, P2_R2278_U76);
  not ginst11495 (P2_R2278_U44, P2_INSTADDRPOINTER_REG_15__SCAN_IN);
  nand ginst11496 (P2_R2278_U440, P2_R2278_U77, P2_U2795);
  nand ginst11497 (P2_R2278_U441, P2_R2278_U439, P2_R2278_U440);
  nand ginst11498 (P2_R2278_U442, P2_R2278_U172, P2_R2278_U173);
  nand ginst11499 (P2_R2278_U443, P2_R2278_U291, P2_R2278_U441);
  nand ginst11500 (P2_R2278_U444, P2_INSTADDRPOINTER_REG_25__SCAN_IN, P2_R2278_U174);
  nand ginst11501 (P2_R2278_U445, P2_R2278_U289, P2_R2278_U73);
  nand ginst11502 (P2_R2278_U446, P2_INSTADDRPOINTER_REG_25__SCAN_IN, P2_R2278_U174);
  nand ginst11503 (P2_R2278_U447, P2_R2278_U289, P2_R2278_U73);
  nand ginst11504 (P2_R2278_U448, P2_R2278_U446, P2_R2278_U447);
  nand ginst11505 (P2_R2278_U449, P2_R2278_U444, P2_R2278_U445, P2_R2278_U72);
  not ginst11506 (P2_R2278_U45, P2_U2808);
  nand ginst11507 (P2_R2278_U450, P2_R2278_U448, P2_U2796);
  nand ginst11508 (P2_R2278_U451, P2_INSTADDRPOINTER_REG_24__SCAN_IN, P2_R2278_U35);
  nand ginst11509 (P2_R2278_U452, P2_R2278_U36, P2_U2797);
  nand ginst11510 (P2_R2278_U453, P2_INSTADDRPOINTER_REG_24__SCAN_IN, P2_R2278_U35);
  nand ginst11511 (P2_R2278_U454, P2_R2278_U36, P2_U2797);
  nand ginst11512 (P2_R2278_U455, P2_R2278_U453, P2_R2278_U454);
  nand ginst11513 (P2_R2278_U456, P2_R2278_U175, P2_R2278_U176);
  nand ginst11514 (P2_R2278_U457, P2_R2278_U286, P2_R2278_U455);
  nand ginst11515 (P2_R2278_U458, P2_INSTADDRPOINTER_REG_23__SCAN_IN, P2_R2278_U69);
  nand ginst11516 (P2_R2278_U459, P2_R2278_U70, P2_U2798);
  not ginst11517 (P2_R2278_U46, P2_INSTADDRPOINTER_REG_13__SCAN_IN);
  nand ginst11518 (P2_R2278_U460, P2_INSTADDRPOINTER_REG_23__SCAN_IN, P2_R2278_U69);
  nand ginst11519 (P2_R2278_U461, P2_R2278_U70, P2_U2798);
  nand ginst11520 (P2_R2278_U462, P2_R2278_U460, P2_R2278_U461);
  nand ginst11521 (P2_R2278_U463, P2_R2278_U177, P2_R2278_U178);
  nand ginst11522 (P2_R2278_U464, P2_R2278_U282, P2_R2278_U462);
  nand ginst11523 (P2_R2278_U465, P2_INSTADDRPOINTER_REG_22__SCAN_IN, P2_R2278_U37);
  nand ginst11524 (P2_R2278_U466, P2_R2278_U38, P2_U2799);
  nand ginst11525 (P2_R2278_U467, P2_INSTADDRPOINTER_REG_22__SCAN_IN, P2_R2278_U37);
  nand ginst11526 (P2_R2278_U468, P2_R2278_U38, P2_U2799);
  nand ginst11527 (P2_R2278_U469, P2_R2278_U467, P2_R2278_U468);
  not ginst11528 (P2_R2278_U47, P2_U2810);
  nand ginst11529 (P2_R2278_U470, P2_R2278_U179, P2_R2278_U180);
  nand ginst11530 (P2_R2278_U471, P2_R2278_U279, P2_R2278_U469);
  nand ginst11531 (P2_R2278_U472, P2_INSTADDRPOINTER_REG_21__SCAN_IN, P2_R2278_U66);
  nand ginst11532 (P2_R2278_U473, P2_R2278_U67, P2_U2800);
  nand ginst11533 (P2_R2278_U474, P2_INSTADDRPOINTER_REG_21__SCAN_IN, P2_R2278_U66);
  nand ginst11534 (P2_R2278_U475, P2_R2278_U67, P2_U2800);
  nand ginst11535 (P2_R2278_U476, P2_R2278_U474, P2_R2278_U475);
  nand ginst11536 (P2_R2278_U477, P2_R2278_U181, P2_R2278_U182);
  nand ginst11537 (P2_R2278_U478, P2_R2278_U275, P2_R2278_U476);
  nand ginst11538 (P2_R2278_U479, P2_INSTADDRPOINTER_REG_20__SCAN_IN, P2_R2278_U39);
  not ginst11539 (P2_R2278_U48, P2_INSTADDRPOINTER_REG_11__SCAN_IN);
  nand ginst11540 (P2_R2278_U480, P2_R2278_U40, P2_U2801);
  nand ginst11541 (P2_R2278_U481, P2_INSTADDRPOINTER_REG_20__SCAN_IN, P2_R2278_U39);
  nand ginst11542 (P2_R2278_U482, P2_R2278_U40, P2_U2801);
  nand ginst11543 (P2_R2278_U483, P2_R2278_U481, P2_R2278_U482);
  nand ginst11544 (P2_R2278_U484, P2_R2278_U183, P2_R2278_U184);
  nand ginst11545 (P2_R2278_U485, P2_R2278_U272, P2_R2278_U483);
  nand ginst11546 (P2_R2278_U486, P2_INSTADDRPOINTER_REG_1__SCAN_IN, P2_R2278_U15);
  nand ginst11547 (P2_R2278_U487, P2_R2278_U17, P2_R2278_U208);
  nand ginst11548 (P2_R2278_U488, P2_R2278_U486, P2_R2278_U487);
  nand ginst11549 (P2_R2278_U489, P2_R2278_U15, P2_R2278_U17, P2_U3637);
  nand ginst11550 (P2_R2278_U49, P2_INSTADDRPOINTER_REG_8__SCAN_IN, P2_U3630);
  nand ginst11551 (P2_R2278_U490, P2_R2278_U16, P2_R2278_U488);
  nand ginst11552 (P2_R2278_U491, P2_INSTADDRPOINTER_REG_19__SCAN_IN, P2_R2278_U62);
  nand ginst11553 (P2_R2278_U492, P2_R2278_U63, P2_U2802);
  nand ginst11554 (P2_R2278_U493, P2_INSTADDRPOINTER_REG_19__SCAN_IN, P2_R2278_U62);
  nand ginst11555 (P2_R2278_U494, P2_R2278_U63, P2_U2802);
  nand ginst11556 (P2_R2278_U495, P2_R2278_U493, P2_R2278_U494);
  nand ginst11557 (P2_R2278_U496, P2_R2278_U185, P2_R2278_U186);
  nand ginst11558 (P2_R2278_U497, P2_R2278_U269, P2_R2278_U495);
  nand ginst11559 (P2_R2278_U498, P2_INSTADDRPOINTER_REG_18__SCAN_IN, P2_R2278_U64);
  nand ginst11560 (P2_R2278_U499, P2_R2278_U65, P2_U2803);
  and ginst11561 (P2_R2278_U5, P2_R2278_U161, P2_R2278_U206, P2_R2278_U309);
  not ginst11562 (P2_R2278_U50, P2_U2811);
  nand ginst11563 (P2_R2278_U500, P2_INSTADDRPOINTER_REG_18__SCAN_IN, P2_R2278_U64);
  nand ginst11564 (P2_R2278_U501, P2_R2278_U65, P2_U2803);
  nand ginst11565 (P2_R2278_U502, P2_R2278_U500, P2_R2278_U501);
  nand ginst11566 (P2_R2278_U503, P2_R2278_U187, P2_R2278_U188);
  nand ginst11567 (P2_R2278_U504, P2_R2278_U265, P2_R2278_U502);
  nand ginst11568 (P2_R2278_U505, P2_INSTADDRPOINTER_REG_17__SCAN_IN, P2_R2278_U41);
  nand ginst11569 (P2_R2278_U506, P2_R2278_U42, P2_U2804);
  nand ginst11570 (P2_R2278_U507, P2_INSTADDRPOINTER_REG_17__SCAN_IN, P2_R2278_U41);
  nand ginst11571 (P2_R2278_U508, P2_R2278_U42, P2_U2804);
  nand ginst11572 (P2_R2278_U509, P2_R2278_U507, P2_R2278_U508);
  not ginst11573 (P2_R2278_U51, P2_INSTADDRPOINTER_REG_10__SCAN_IN);
  nand ginst11574 (P2_R2278_U510, P2_R2278_U189, P2_R2278_U190);
  nand ginst11575 (P2_R2278_U511, P2_R2278_U262, P2_R2278_U509);
  nand ginst11576 (P2_R2278_U512, P2_INSTADDRPOINTER_REG_16__SCAN_IN, P2_R2278_U59);
  nand ginst11577 (P2_R2278_U513, P2_R2278_U60, P2_U2805);
  nand ginst11578 (P2_R2278_U514, P2_INSTADDRPOINTER_REG_16__SCAN_IN, P2_R2278_U59);
  nand ginst11579 (P2_R2278_U515, P2_R2278_U60, P2_U2805);
  nand ginst11580 (P2_R2278_U516, P2_R2278_U514, P2_R2278_U515);
  nand ginst11581 (P2_R2278_U517, P2_R2278_U191, P2_R2278_U192);
  nand ginst11582 (P2_R2278_U518, P2_R2278_U258, P2_R2278_U516);
  nand ginst11583 (P2_R2278_U519, P2_INSTADDRPOINTER_REG_15__SCAN_IN, P2_R2278_U43);
  nand ginst11584 (P2_R2278_U52, P2_INSTADDRPOINTER_REG_10__SCAN_IN, P2_U2811);
  nand ginst11585 (P2_R2278_U520, P2_R2278_U44, P2_U2806);
  nand ginst11586 (P2_R2278_U521, P2_INSTADDRPOINTER_REG_15__SCAN_IN, P2_R2278_U43);
  nand ginst11587 (P2_R2278_U522, P2_R2278_U44, P2_U2806);
  nand ginst11588 (P2_R2278_U523, P2_R2278_U521, P2_R2278_U522);
  nand ginst11589 (P2_R2278_U524, P2_R2278_U193, P2_R2278_U194);
  nand ginst11590 (P2_R2278_U525, P2_R2278_U255, P2_R2278_U523);
  nand ginst11591 (P2_R2278_U526, P2_INSTADDRPOINTER_REG_14__SCAN_IN, P2_R2278_U56);
  nand ginst11592 (P2_R2278_U527, P2_R2278_U57, P2_U2807);
  nand ginst11593 (P2_R2278_U528, P2_INSTADDRPOINTER_REG_14__SCAN_IN, P2_R2278_U56);
  nand ginst11594 (P2_R2278_U529, P2_R2278_U57, P2_U2807);
  not ginst11595 (P2_R2278_U53, P2_U2809);
  nand ginst11596 (P2_R2278_U530, P2_R2278_U528, P2_R2278_U529);
  nand ginst11597 (P2_R2278_U531, P2_R2278_U195, P2_R2278_U196);
  nand ginst11598 (P2_R2278_U532, P2_R2278_U251, P2_R2278_U530);
  nand ginst11599 (P2_R2278_U533, P2_INSTADDRPOINTER_REG_13__SCAN_IN, P2_R2278_U45);
  nand ginst11600 (P2_R2278_U534, P2_R2278_U46, P2_U2808);
  nand ginst11601 (P2_R2278_U535, P2_INSTADDRPOINTER_REG_13__SCAN_IN, P2_R2278_U45);
  nand ginst11602 (P2_R2278_U536, P2_R2278_U46, P2_U2808);
  nand ginst11603 (P2_R2278_U537, P2_R2278_U535, P2_R2278_U536);
  nand ginst11604 (P2_R2278_U538, P2_R2278_U197, P2_R2278_U198);
  nand ginst11605 (P2_R2278_U539, P2_R2278_U248, P2_R2278_U537);
  not ginst11606 (P2_R2278_U54, P2_INSTADDRPOINTER_REG_12__SCAN_IN);
  nand ginst11607 (P2_R2278_U540, P2_INSTADDRPOINTER_REG_12__SCAN_IN, P2_R2278_U53);
  nand ginst11608 (P2_R2278_U541, P2_R2278_U54, P2_U2809);
  nand ginst11609 (P2_R2278_U542, P2_INSTADDRPOINTER_REG_12__SCAN_IN, P2_R2278_U53);
  nand ginst11610 (P2_R2278_U543, P2_R2278_U54, P2_U2809);
  nand ginst11611 (P2_R2278_U544, P2_R2278_U542, P2_R2278_U543);
  nand ginst11612 (P2_R2278_U545, P2_R2278_U199, P2_R2278_U200);
  nand ginst11613 (P2_R2278_U546, P2_R2278_U244, P2_R2278_U544);
  nand ginst11614 (P2_R2278_U547, P2_INSTADDRPOINTER_REG_11__SCAN_IN, P2_R2278_U47);
  nand ginst11615 (P2_R2278_U548, P2_R2278_U48, P2_U2810);
  nand ginst11616 (P2_R2278_U549, P2_INSTADDRPOINTER_REG_11__SCAN_IN, P2_R2278_U47);
  nand ginst11617 (P2_R2278_U55, P2_INSTADDRPOINTER_REG_12__SCAN_IN, P2_U2809);
  nand ginst11618 (P2_R2278_U550, P2_R2278_U48, P2_U2810);
  nand ginst11619 (P2_R2278_U551, P2_R2278_U549, P2_R2278_U550);
  nand ginst11620 (P2_R2278_U552, P2_R2278_U201, P2_R2278_U202);
  nand ginst11621 (P2_R2278_U553, P2_R2278_U241, P2_R2278_U551);
  nand ginst11622 (P2_R2278_U554, P2_INSTADDRPOINTER_REG_10__SCAN_IN, P2_R2278_U50);
  nand ginst11623 (P2_R2278_U555, P2_R2278_U51, P2_U2811);
  nand ginst11624 (P2_R2278_U556, P2_INSTADDRPOINTER_REG_10__SCAN_IN, P2_R2278_U50);
  nand ginst11625 (P2_R2278_U557, P2_R2278_U51, P2_U2811);
  nand ginst11626 (P2_R2278_U558, P2_R2278_U556, P2_R2278_U557);
  nand ginst11627 (P2_R2278_U559, P2_R2278_U203, P2_R2278_U204);
  not ginst11628 (P2_R2278_U56, P2_U2807);
  nand ginst11629 (P2_R2278_U560, P2_R2278_U237, P2_R2278_U558);
  nand ginst11630 (P2_R2278_U561, P2_INSTADDRPOINTER_REG_0__SCAN_IN, P2_R2278_U13);
  nand ginst11631 (P2_R2278_U562, P2_R2278_U14, P2_U3638);
  not ginst11632 (P2_R2278_U57, P2_INSTADDRPOINTER_REG_14__SCAN_IN);
  nand ginst11633 (P2_R2278_U58, P2_INSTADDRPOINTER_REG_14__SCAN_IN, P2_U2807);
  not ginst11634 (P2_R2278_U59, P2_U2805);
  nand ginst11635 (P2_R2278_U6, P2_R2278_U345, P2_R2278_U489, P2_R2278_U490);
  not ginst11636 (P2_R2278_U60, P2_INSTADDRPOINTER_REG_16__SCAN_IN);
  nand ginst11637 (P2_R2278_U61, P2_INSTADDRPOINTER_REG_16__SCAN_IN, P2_U2805);
  not ginst11638 (P2_R2278_U62, P2_U2802);
  not ginst11639 (P2_R2278_U63, P2_INSTADDRPOINTER_REG_19__SCAN_IN);
  not ginst11640 (P2_R2278_U64, P2_U2803);
  not ginst11641 (P2_R2278_U65, P2_INSTADDRPOINTER_REG_18__SCAN_IN);
  not ginst11642 (P2_R2278_U66, P2_U2800);
  not ginst11643 (P2_R2278_U67, P2_INSTADDRPOINTER_REG_21__SCAN_IN);
  nand ginst11644 (P2_R2278_U68, P2_INSTADDRPOINTER_REG_21__SCAN_IN, P2_U2800);
  not ginst11645 (P2_R2278_U69, P2_U2798);
  not ginst11646 (P2_R2278_U7, P2_U3631);
  not ginst11647 (P2_R2278_U70, P2_INSTADDRPOINTER_REG_23__SCAN_IN);
  nand ginst11648 (P2_R2278_U71, P2_INSTADDRPOINTER_REG_23__SCAN_IN, P2_U2798);
  not ginst11649 (P2_R2278_U72, P2_U2796);
  not ginst11650 (P2_R2278_U73, P2_INSTADDRPOINTER_REG_25__SCAN_IN);
  not ginst11651 (P2_R2278_U74, P2_U2794);
  not ginst11652 (P2_R2278_U75, P2_INSTADDRPOINTER_REG_27__SCAN_IN);
  not ginst11653 (P2_R2278_U76, P2_U2795);
  not ginst11654 (P2_R2278_U77, P2_INSTADDRPOINTER_REG_26__SCAN_IN);
  nand ginst11655 (P2_R2278_U78, P2_INSTADDRPOINTER_REG_26__SCAN_IN, P2_U2795);
  not ginst11656 (P2_R2278_U79, P2_U2791);
  not ginst11657 (P2_R2278_U8, P2_INSTADDRPOINTER_REG_7__SCAN_IN);
  not ginst11658 (P2_R2278_U80, P2_INSTADDRPOINTER_REG_30__SCAN_IN);
  nand ginst11659 (P2_R2278_U81, P2_R2278_U297, P2_R2278_U340);
  nand ginst11660 (P2_R2278_U82, P2_R2278_U208, P2_U3637);
  nand ginst11661 (P2_R2278_U83, P2_R2278_U561, P2_R2278_U562);
  nand ginst11662 (P2_R2278_U84, P2_R2278_U351, P2_R2278_U352);
  nand ginst11663 (P2_R2278_U85, P2_R2278_U358, P2_R2278_U359);
  nand ginst11664 (P2_R2278_U86, P2_R2278_U365, P2_R2278_U366);
  nand ginst11665 (P2_R2278_U87, P2_R2278_U372, P2_R2278_U373);
  nand ginst11666 (P2_R2278_U88, P2_R2278_U379, P2_R2278_U380);
  nand ginst11667 (P2_R2278_U89, P2_R2278_U386, P2_R2278_U387);
  not ginst11668 (P2_R2278_U9, P2_U3633);
  nand ginst11669 (P2_R2278_U90, P2_R2278_U393, P2_R2278_U394);
  nand ginst11670 (P2_R2278_U91, P2_R2278_U407, P2_R2278_U408);
  nand ginst11671 (P2_R2278_U92, P2_R2278_U414, P2_R2278_U415);
  nand ginst11672 (P2_R2278_U93, P2_R2278_U421, P2_R2278_U422);
  nand ginst11673 (P2_R2278_U94, P2_R2278_U428, P2_R2278_U429);
  nand ginst11674 (P2_R2278_U95, P2_R2278_U435, P2_R2278_U436);
  nand ginst11675 (P2_R2278_U96, P2_R2278_U442, P2_R2278_U443);
  nand ginst11676 (P2_R2278_U97, P2_R2278_U449, P2_R2278_U450);
  nand ginst11677 (P2_R2278_U98, P2_R2278_U456, P2_R2278_U457);
  nand ginst11678 (P2_R2278_U99, P2_R2278_U463, P2_R2278_U464);
  not ginst11679 (P2_R2337_U10, P2_PHYADDRPOINTER_REG_5__SCAN_IN);
  not ginst11680 (P2_R2337_U100, P2_R2337_U18);
  not ginst11681 (P2_R2337_U101, P2_R2337_U19);
  not ginst11682 (P2_R2337_U102, P2_R2337_U21);
  not ginst11683 (P2_R2337_U103, P2_R2337_U23);
  not ginst11684 (P2_R2337_U104, P2_R2337_U25);
  not ginst11685 (P2_R2337_U105, P2_R2337_U27);
  not ginst11686 (P2_R2337_U106, P2_R2337_U29);
  not ginst11687 (P2_R2337_U107, P2_R2337_U31);
  not ginst11688 (P2_R2337_U108, P2_R2337_U33);
  not ginst11689 (P2_R2337_U109, P2_R2337_U35);
  nand ginst11690 (P2_R2337_U11, P2_PHYADDRPOINTER_REG_5__SCAN_IN, P2_R2337_U96);
  not ginst11691 (P2_R2337_U110, P2_R2337_U37);
  not ginst11692 (P2_R2337_U111, P2_R2337_U39);
  not ginst11693 (P2_R2337_U112, P2_R2337_U41);
  not ginst11694 (P2_R2337_U113, P2_R2337_U43);
  not ginst11695 (P2_R2337_U114, P2_R2337_U45);
  not ginst11696 (P2_R2337_U115, P2_R2337_U47);
  not ginst11697 (P2_R2337_U116, P2_R2337_U49);
  not ginst11698 (P2_R2337_U117, P2_R2337_U51);
  not ginst11699 (P2_R2337_U118, P2_R2337_U53);
  not ginst11700 (P2_R2337_U119, P2_R2337_U55);
  not ginst11701 (P2_R2337_U12, P2_PHYADDRPOINTER_REG_6__SCAN_IN);
  not ginst11702 (P2_R2337_U120, P2_R2337_U57);
  not ginst11703 (P2_R2337_U121, P2_R2337_U59);
  not ginst11704 (P2_R2337_U122, P2_R2337_U93);
  nand ginst11705 (P2_R2337_U123, P2_PHYADDRPOINTER_REG_9__SCAN_IN, P2_R2337_U18);
  nand ginst11706 (P2_R2337_U124, P2_R2337_U100, P2_R2337_U17);
  nand ginst11707 (P2_R2337_U125, P2_PHYADDRPOINTER_REG_8__SCAN_IN, P2_R2337_U15);
  nand ginst11708 (P2_R2337_U126, P2_R2337_U16, P2_R2337_U99);
  nand ginst11709 (P2_R2337_U127, P2_PHYADDRPOINTER_REG_7__SCAN_IN, P2_R2337_U13);
  nand ginst11710 (P2_R2337_U128, P2_R2337_U14, P2_R2337_U98);
  nand ginst11711 (P2_R2337_U129, P2_PHYADDRPOINTER_REG_6__SCAN_IN, P2_R2337_U11);
  nand ginst11712 (P2_R2337_U13, P2_PHYADDRPOINTER_REG_6__SCAN_IN, P2_R2337_U97);
  nand ginst11713 (P2_R2337_U130, P2_R2337_U12, P2_R2337_U97);
  nand ginst11714 (P2_R2337_U131, P2_PHYADDRPOINTER_REG_5__SCAN_IN, P2_R2337_U9);
  nand ginst11715 (P2_R2337_U132, P2_R2337_U10, P2_R2337_U96);
  nand ginst11716 (P2_R2337_U133, P2_PHYADDRPOINTER_REG_4__SCAN_IN, P2_R2337_U7);
  nand ginst11717 (P2_R2337_U134, P2_R2337_U8, P2_R2337_U95);
  nand ginst11718 (P2_R2337_U135, P2_PHYADDRPOINTER_REG_3__SCAN_IN, P2_R2337_U91);
  nand ginst11719 (P2_R2337_U136, P2_R2337_U5, P2_R2337_U94);
  nand ginst11720 (P2_R2337_U137, P2_PHYADDRPOINTER_REG_31__SCAN_IN, P2_R2337_U93);
  nand ginst11721 (P2_R2337_U138, P2_R2337_U122, P2_R2337_U92);
  nand ginst11722 (P2_R2337_U139, P2_PHYADDRPOINTER_REG_30__SCAN_IN, P2_R2337_U59);
  not ginst11723 (P2_R2337_U14, P2_PHYADDRPOINTER_REG_7__SCAN_IN);
  nand ginst11724 (P2_R2337_U140, P2_R2337_U121, P2_R2337_U60);
  nand ginst11725 (P2_R2337_U141, P2_PHYADDRPOINTER_REG_2__SCAN_IN, P2_R2337_U4);
  nand ginst11726 (P2_R2337_U142, P2_PHYADDRPOINTER_REG_1__SCAN_IN, P2_R2337_U6);
  nand ginst11727 (P2_R2337_U143, P2_PHYADDRPOINTER_REG_29__SCAN_IN, P2_R2337_U57);
  nand ginst11728 (P2_R2337_U144, P2_R2337_U120, P2_R2337_U58);
  nand ginst11729 (P2_R2337_U145, P2_PHYADDRPOINTER_REG_28__SCAN_IN, P2_R2337_U55);
  nand ginst11730 (P2_R2337_U146, P2_R2337_U119, P2_R2337_U56);
  nand ginst11731 (P2_R2337_U147, P2_PHYADDRPOINTER_REG_27__SCAN_IN, P2_R2337_U53);
  nand ginst11732 (P2_R2337_U148, P2_R2337_U118, P2_R2337_U54);
  nand ginst11733 (P2_R2337_U149, P2_PHYADDRPOINTER_REG_26__SCAN_IN, P2_R2337_U51);
  nand ginst11734 (P2_R2337_U15, P2_PHYADDRPOINTER_REG_7__SCAN_IN, P2_R2337_U98);
  nand ginst11735 (P2_R2337_U150, P2_R2337_U117, P2_R2337_U52);
  nand ginst11736 (P2_R2337_U151, P2_PHYADDRPOINTER_REG_25__SCAN_IN, P2_R2337_U49);
  nand ginst11737 (P2_R2337_U152, P2_R2337_U116, P2_R2337_U50);
  nand ginst11738 (P2_R2337_U153, P2_PHYADDRPOINTER_REG_24__SCAN_IN, P2_R2337_U47);
  nand ginst11739 (P2_R2337_U154, P2_R2337_U115, P2_R2337_U48);
  nand ginst11740 (P2_R2337_U155, P2_PHYADDRPOINTER_REG_23__SCAN_IN, P2_R2337_U45);
  nand ginst11741 (P2_R2337_U156, P2_R2337_U114, P2_R2337_U46);
  nand ginst11742 (P2_R2337_U157, P2_PHYADDRPOINTER_REG_22__SCAN_IN, P2_R2337_U43);
  nand ginst11743 (P2_R2337_U158, P2_R2337_U113, P2_R2337_U44);
  nand ginst11744 (P2_R2337_U159, P2_PHYADDRPOINTER_REG_21__SCAN_IN, P2_R2337_U41);
  not ginst11745 (P2_R2337_U16, P2_PHYADDRPOINTER_REG_8__SCAN_IN);
  nand ginst11746 (P2_R2337_U160, P2_R2337_U112, P2_R2337_U42);
  nand ginst11747 (P2_R2337_U161, P2_PHYADDRPOINTER_REG_20__SCAN_IN, P2_R2337_U39);
  nand ginst11748 (P2_R2337_U162, P2_R2337_U111, P2_R2337_U40);
  nand ginst11749 (P2_R2337_U163, P2_PHYADDRPOINTER_REG_19__SCAN_IN, P2_R2337_U37);
  nand ginst11750 (P2_R2337_U164, P2_R2337_U110, P2_R2337_U38);
  nand ginst11751 (P2_R2337_U165, P2_PHYADDRPOINTER_REG_18__SCAN_IN, P2_R2337_U35);
  nand ginst11752 (P2_R2337_U166, P2_R2337_U109, P2_R2337_U36);
  nand ginst11753 (P2_R2337_U167, P2_PHYADDRPOINTER_REG_17__SCAN_IN, P2_R2337_U33);
  nand ginst11754 (P2_R2337_U168, P2_R2337_U108, P2_R2337_U34);
  nand ginst11755 (P2_R2337_U169, P2_PHYADDRPOINTER_REG_16__SCAN_IN, P2_R2337_U31);
  not ginst11756 (P2_R2337_U17, P2_PHYADDRPOINTER_REG_9__SCAN_IN);
  nand ginst11757 (P2_R2337_U170, P2_R2337_U107, P2_R2337_U32);
  nand ginst11758 (P2_R2337_U171, P2_PHYADDRPOINTER_REG_15__SCAN_IN, P2_R2337_U29);
  nand ginst11759 (P2_R2337_U172, P2_R2337_U106, P2_R2337_U30);
  nand ginst11760 (P2_R2337_U173, P2_PHYADDRPOINTER_REG_14__SCAN_IN, P2_R2337_U27);
  nand ginst11761 (P2_R2337_U174, P2_R2337_U105, P2_R2337_U28);
  nand ginst11762 (P2_R2337_U175, P2_PHYADDRPOINTER_REG_13__SCAN_IN, P2_R2337_U25);
  nand ginst11763 (P2_R2337_U176, P2_R2337_U104, P2_R2337_U26);
  nand ginst11764 (P2_R2337_U177, P2_PHYADDRPOINTER_REG_12__SCAN_IN, P2_R2337_U23);
  nand ginst11765 (P2_R2337_U178, P2_R2337_U103, P2_R2337_U24);
  nand ginst11766 (P2_R2337_U179, P2_PHYADDRPOINTER_REG_11__SCAN_IN, P2_R2337_U21);
  nand ginst11767 (P2_R2337_U18, P2_PHYADDRPOINTER_REG_8__SCAN_IN, P2_R2337_U99);
  nand ginst11768 (P2_R2337_U180, P2_R2337_U102, P2_R2337_U22);
  nand ginst11769 (P2_R2337_U181, P2_PHYADDRPOINTER_REG_10__SCAN_IN, P2_R2337_U19);
  nand ginst11770 (P2_R2337_U182, P2_R2337_U101, P2_R2337_U20);
  nand ginst11771 (P2_R2337_U19, P2_PHYADDRPOINTER_REG_9__SCAN_IN, P2_R2337_U100);
  not ginst11772 (P2_R2337_U20, P2_PHYADDRPOINTER_REG_10__SCAN_IN);
  nand ginst11773 (P2_R2337_U21, P2_PHYADDRPOINTER_REG_10__SCAN_IN, P2_R2337_U101);
  not ginst11774 (P2_R2337_U22, P2_PHYADDRPOINTER_REG_11__SCAN_IN);
  nand ginst11775 (P2_R2337_U23, P2_PHYADDRPOINTER_REG_11__SCAN_IN, P2_R2337_U102);
  not ginst11776 (P2_R2337_U24, P2_PHYADDRPOINTER_REG_12__SCAN_IN);
  nand ginst11777 (P2_R2337_U25, P2_PHYADDRPOINTER_REG_12__SCAN_IN, P2_R2337_U103);
  not ginst11778 (P2_R2337_U26, P2_PHYADDRPOINTER_REG_13__SCAN_IN);
  nand ginst11779 (P2_R2337_U27, P2_PHYADDRPOINTER_REG_13__SCAN_IN, P2_R2337_U104);
  not ginst11780 (P2_R2337_U28, P2_PHYADDRPOINTER_REG_14__SCAN_IN);
  nand ginst11781 (P2_R2337_U29, P2_PHYADDRPOINTER_REG_14__SCAN_IN, P2_R2337_U105);
  not ginst11782 (P2_R2337_U30, P2_PHYADDRPOINTER_REG_15__SCAN_IN);
  nand ginst11783 (P2_R2337_U31, P2_PHYADDRPOINTER_REG_15__SCAN_IN, P2_R2337_U106);
  not ginst11784 (P2_R2337_U32, P2_PHYADDRPOINTER_REG_16__SCAN_IN);
  nand ginst11785 (P2_R2337_U33, P2_PHYADDRPOINTER_REG_16__SCAN_IN, P2_R2337_U107);
  not ginst11786 (P2_R2337_U34, P2_PHYADDRPOINTER_REG_17__SCAN_IN);
  nand ginst11787 (P2_R2337_U35, P2_PHYADDRPOINTER_REG_17__SCAN_IN, P2_R2337_U108);
  not ginst11788 (P2_R2337_U36, P2_PHYADDRPOINTER_REG_18__SCAN_IN);
  nand ginst11789 (P2_R2337_U37, P2_PHYADDRPOINTER_REG_18__SCAN_IN, P2_R2337_U109);
  not ginst11790 (P2_R2337_U38, P2_PHYADDRPOINTER_REG_19__SCAN_IN);
  nand ginst11791 (P2_R2337_U39, P2_PHYADDRPOINTER_REG_19__SCAN_IN, P2_R2337_U110);
  not ginst11792 (P2_R2337_U4, P2_PHYADDRPOINTER_REG_1__SCAN_IN);
  not ginst11793 (P2_R2337_U40, P2_PHYADDRPOINTER_REG_20__SCAN_IN);
  nand ginst11794 (P2_R2337_U41, P2_PHYADDRPOINTER_REG_20__SCAN_IN, P2_R2337_U111);
  not ginst11795 (P2_R2337_U42, P2_PHYADDRPOINTER_REG_21__SCAN_IN);
  nand ginst11796 (P2_R2337_U43, P2_PHYADDRPOINTER_REG_21__SCAN_IN, P2_R2337_U112);
  not ginst11797 (P2_R2337_U44, P2_PHYADDRPOINTER_REG_22__SCAN_IN);
  nand ginst11798 (P2_R2337_U45, P2_PHYADDRPOINTER_REG_22__SCAN_IN, P2_R2337_U113);
  not ginst11799 (P2_R2337_U46, P2_PHYADDRPOINTER_REG_23__SCAN_IN);
  nand ginst11800 (P2_R2337_U47, P2_PHYADDRPOINTER_REG_23__SCAN_IN, P2_R2337_U114);
  not ginst11801 (P2_R2337_U48, P2_PHYADDRPOINTER_REG_24__SCAN_IN);
  nand ginst11802 (P2_R2337_U49, P2_PHYADDRPOINTER_REG_24__SCAN_IN, P2_R2337_U115);
  not ginst11803 (P2_R2337_U5, P2_PHYADDRPOINTER_REG_3__SCAN_IN);
  not ginst11804 (P2_R2337_U50, P2_PHYADDRPOINTER_REG_25__SCAN_IN);
  nand ginst11805 (P2_R2337_U51, P2_PHYADDRPOINTER_REG_25__SCAN_IN, P2_R2337_U116);
  not ginst11806 (P2_R2337_U52, P2_PHYADDRPOINTER_REG_26__SCAN_IN);
  nand ginst11807 (P2_R2337_U53, P2_PHYADDRPOINTER_REG_26__SCAN_IN, P2_R2337_U117);
  not ginst11808 (P2_R2337_U54, P2_PHYADDRPOINTER_REG_27__SCAN_IN);
  nand ginst11809 (P2_R2337_U55, P2_PHYADDRPOINTER_REG_27__SCAN_IN, P2_R2337_U118);
  not ginst11810 (P2_R2337_U56, P2_PHYADDRPOINTER_REG_28__SCAN_IN);
  nand ginst11811 (P2_R2337_U57, P2_PHYADDRPOINTER_REG_28__SCAN_IN, P2_R2337_U119);
  not ginst11812 (P2_R2337_U58, P2_PHYADDRPOINTER_REG_29__SCAN_IN);
  nand ginst11813 (P2_R2337_U59, P2_PHYADDRPOINTER_REG_29__SCAN_IN, P2_R2337_U120);
  not ginst11814 (P2_R2337_U6, P2_PHYADDRPOINTER_REG_2__SCAN_IN);
  not ginst11815 (P2_R2337_U60, P2_PHYADDRPOINTER_REG_30__SCAN_IN);
  nand ginst11816 (P2_R2337_U61, P2_R2337_U123, P2_R2337_U124);
  nand ginst11817 (P2_R2337_U62, P2_R2337_U125, P2_R2337_U126);
  nand ginst11818 (P2_R2337_U63, P2_R2337_U127, P2_R2337_U128);
  nand ginst11819 (P2_R2337_U64, P2_R2337_U129, P2_R2337_U130);
  nand ginst11820 (P2_R2337_U65, P2_R2337_U131, P2_R2337_U132);
  nand ginst11821 (P2_R2337_U66, P2_R2337_U133, P2_R2337_U134);
  nand ginst11822 (P2_R2337_U67, P2_R2337_U135, P2_R2337_U136);
  nand ginst11823 (P2_R2337_U68, P2_R2337_U137, P2_R2337_U138);
  nand ginst11824 (P2_R2337_U69, P2_R2337_U139, P2_R2337_U140);
  nand ginst11825 (P2_R2337_U7, P2_PHYADDRPOINTER_REG_1__SCAN_IN, P2_PHYADDRPOINTER_REG_2__SCAN_IN, P2_PHYADDRPOINTER_REG_3__SCAN_IN);
  nand ginst11826 (P2_R2337_U70, P2_R2337_U141, P2_R2337_U142);
  nand ginst11827 (P2_R2337_U71, P2_R2337_U143, P2_R2337_U144);
  nand ginst11828 (P2_R2337_U72, P2_R2337_U145, P2_R2337_U146);
  nand ginst11829 (P2_R2337_U73, P2_R2337_U147, P2_R2337_U148);
  nand ginst11830 (P2_R2337_U74, P2_R2337_U149, P2_R2337_U150);
  nand ginst11831 (P2_R2337_U75, P2_R2337_U151, P2_R2337_U152);
  nand ginst11832 (P2_R2337_U76, P2_R2337_U153, P2_R2337_U154);
  nand ginst11833 (P2_R2337_U77, P2_R2337_U155, P2_R2337_U156);
  nand ginst11834 (P2_R2337_U78, P2_R2337_U157, P2_R2337_U158);
  nand ginst11835 (P2_R2337_U79, P2_R2337_U159, P2_R2337_U160);
  not ginst11836 (P2_R2337_U8, P2_PHYADDRPOINTER_REG_4__SCAN_IN);
  nand ginst11837 (P2_R2337_U80, P2_R2337_U161, P2_R2337_U162);
  nand ginst11838 (P2_R2337_U81, P2_R2337_U163, P2_R2337_U164);
  nand ginst11839 (P2_R2337_U82, P2_R2337_U165, P2_R2337_U166);
  nand ginst11840 (P2_R2337_U83, P2_R2337_U167, P2_R2337_U168);
  nand ginst11841 (P2_R2337_U84, P2_R2337_U169, P2_R2337_U170);
  nand ginst11842 (P2_R2337_U85, P2_R2337_U171, P2_R2337_U172);
  nand ginst11843 (P2_R2337_U86, P2_R2337_U173, P2_R2337_U174);
  nand ginst11844 (P2_R2337_U87, P2_R2337_U175, P2_R2337_U176);
  nand ginst11845 (P2_R2337_U88, P2_R2337_U177, P2_R2337_U178);
  nand ginst11846 (P2_R2337_U89, P2_R2337_U179, P2_R2337_U180);
  nand ginst11847 (P2_R2337_U9, P2_PHYADDRPOINTER_REG_4__SCAN_IN, P2_R2337_U95);
  nand ginst11848 (P2_R2337_U90, P2_R2337_U181, P2_R2337_U182);
  nand ginst11849 (P2_R2337_U91, P2_PHYADDRPOINTER_REG_1__SCAN_IN, P2_PHYADDRPOINTER_REG_2__SCAN_IN);
  not ginst11850 (P2_R2337_U92, P2_PHYADDRPOINTER_REG_31__SCAN_IN);
  nand ginst11851 (P2_R2337_U93, P2_PHYADDRPOINTER_REG_30__SCAN_IN, P2_R2337_U121);
  not ginst11852 (P2_R2337_U94, P2_R2337_U91);
  not ginst11853 (P2_R2337_U95, P2_R2337_U7);
  not ginst11854 (P2_R2337_U96, P2_R2337_U9);
  not ginst11855 (P2_R2337_U97, P2_R2337_U11);
  not ginst11856 (P2_R2337_U98, P2_R2337_U13);
  not ginst11857 (P2_R2337_U99, P2_R2337_U15);
  not ginst11858 (P2_SUB_450_U10, P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN);
  not ginst11859 (P2_SUB_450_U11, P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN);
  not ginst11860 (P2_SUB_450_U12, P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN);
  not ginst11861 (P2_SUB_450_U13, P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN);
  nand ginst11862 (P2_SUB_450_U14, P2_SUB_450_U38, P2_SUB_450_U39);
  not ginst11863 (P2_SUB_450_U15, P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN);
  not ginst11864 (P2_SUB_450_U16, P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN);
  nand ginst11865 (P2_SUB_450_U17, P2_SUB_450_U47, P2_SUB_450_U48);
  nand ginst11866 (P2_SUB_450_U18, P2_SUB_450_U52, P2_SUB_450_U53);
  nand ginst11867 (P2_SUB_450_U19, P2_SUB_450_U57, P2_SUB_450_U58);
  nand ginst11868 (P2_SUB_450_U20, P2_SUB_450_U62, P2_SUB_450_U63);
  nand ginst11869 (P2_SUB_450_U21, P2_SUB_450_U44, P2_SUB_450_U45);
  nand ginst11870 (P2_SUB_450_U22, P2_SUB_450_U49, P2_SUB_450_U50);
  nand ginst11871 (P2_SUB_450_U23, P2_SUB_450_U54, P2_SUB_450_U55);
  nand ginst11872 (P2_SUB_450_U24, P2_SUB_450_U59, P2_SUB_450_U60);
  nand ginst11873 (P2_SUB_450_U25, P2_SUB_450_U34, P2_SUB_450_U35);
  nand ginst11874 (P2_SUB_450_U26, P2_SUB_450_U30, P2_SUB_450_U31);
  not ginst11875 (P2_SUB_450_U27, P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN);
  not ginst11876 (P2_SUB_450_U28, P2_SUB_450_U7);
  nand ginst11877 (P2_SUB_450_U29, P2_SUB_450_U28, P2_SUB_450_U8);
  nand ginst11878 (P2_SUB_450_U30, P2_SUB_450_U27, P2_SUB_450_U29);
  nand ginst11879 (P2_SUB_450_U31, P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN, P2_SUB_450_U7);
  not ginst11880 (P2_SUB_450_U32, P2_SUB_450_U26);
  nand ginst11881 (P2_SUB_450_U33, P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN, P2_SUB_450_U10);
  nand ginst11882 (P2_SUB_450_U34, P2_SUB_450_U26, P2_SUB_450_U33);
  nand ginst11883 (P2_SUB_450_U35, P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN, P2_SUB_450_U9);
  not ginst11884 (P2_SUB_450_U36, P2_SUB_450_U25);
  nand ginst11885 (P2_SUB_450_U37, P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P2_SUB_450_U12);
  nand ginst11886 (P2_SUB_450_U38, P2_SUB_450_U25, P2_SUB_450_U37);
  nand ginst11887 (P2_SUB_450_U39, P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN, P2_SUB_450_U11);
  not ginst11888 (P2_SUB_450_U40, P2_SUB_450_U14);
  nand ginst11889 (P2_SUB_450_U41, P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN, P2_SUB_450_U15);
  nand ginst11890 (P2_SUB_450_U42, P2_SUB_450_U40, P2_SUB_450_U41);
  nand ginst11891 (P2_SUB_450_U43, P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN, P2_SUB_450_U13);
  nand ginst11892 (P2_SUB_450_U44, P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN, P2_SUB_450_U13);
  nand ginst11893 (P2_SUB_450_U45, P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN, P2_SUB_450_U15);
  not ginst11894 (P2_SUB_450_U46, P2_SUB_450_U21);
  nand ginst11895 (P2_SUB_450_U47, P2_SUB_450_U40, P2_SUB_450_U46);
  nand ginst11896 (P2_SUB_450_U48, P2_SUB_450_U14, P2_SUB_450_U21);
  nand ginst11897 (P2_SUB_450_U49, P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P2_SUB_450_U12);
  nand ginst11898 (P2_SUB_450_U50, P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN, P2_SUB_450_U11);
  not ginst11899 (P2_SUB_450_U51, P2_SUB_450_U22);
  nand ginst11900 (P2_SUB_450_U52, P2_SUB_450_U36, P2_SUB_450_U51);
  nand ginst11901 (P2_SUB_450_U53, P2_SUB_450_U22, P2_SUB_450_U25);
  nand ginst11902 (P2_SUB_450_U54, P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN, P2_SUB_450_U10);
  nand ginst11903 (P2_SUB_450_U55, P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN, P2_SUB_450_U9);
  not ginst11904 (P2_SUB_450_U56, P2_SUB_450_U23);
  nand ginst11905 (P2_SUB_450_U57, P2_SUB_450_U32, P2_SUB_450_U56);
  nand ginst11906 (P2_SUB_450_U58, P2_SUB_450_U23, P2_SUB_450_U26);
  nand ginst11907 (P2_SUB_450_U59, P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P2_SUB_450_U8);
  nand ginst11908 (P2_SUB_450_U6, P2_SUB_450_U42, P2_SUB_450_U43);
  nand ginst11909 (P2_SUB_450_U60, P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN, P2_SUB_450_U27);
  not ginst11910 (P2_SUB_450_U61, P2_SUB_450_U24);
  nand ginst11911 (P2_SUB_450_U62, P2_SUB_450_U28, P2_SUB_450_U61);
  nand ginst11912 (P2_SUB_450_U63, P2_SUB_450_U24, P2_SUB_450_U7);
  nand ginst11913 (P2_SUB_450_U7, P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN, P2_SUB_450_U16);
  not ginst11914 (P2_SUB_450_U8, P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN);
  not ginst11915 (P2_SUB_450_U9, P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN);
  not ginst11916 (P2_SUB_563_U6, P2_U3618);
  not ginst11917 (P2_SUB_563_U7, P2_U3619);
  not ginst11918 (P2_SUB_589_U6, P2_U3614);
  not ginst11919 (P2_SUB_589_U7, P2_U3615);
  not ginst11920 (P2_SUB_589_U8, P2_U2813);
  not ginst11921 (P2_SUB_589_U9, P2_U3613);
  and ginst11922 (P2_U2352, P2_U2617, P2_U3300, P2_U7873);
  and ginst11923 (P2_U2353, P2_U2439, P2_U4343);
  and ginst11924 (P2_U2354, P2_STATE2_REG_0__SCAN_IN, P2_U7861, P2_U7873);
  and ginst11925 (P2_U2355, P2_U2447, P2_U7861);
  and ginst11926 (P2_U2356, P2_STATE2_REG_0__SCAN_IN, P2_U3253);
  and ginst11927 (P2_U2357, P2_U2458, P2_U3712);
  and ginst11928 (P2_U2358, P2_STATE2_REG_0__SCAN_IN, P2_U4431);
  and ginst11929 (P2_U2359, P2_U3265, P2_U4411);
  nor ginst11930 (P2_U2360, P2_STATEBS16_REG_SCAN_IN, U211);
  and ginst11931 (P2_U2361, P2_R2238_U6, P2_U2356);
  and ginst11932 (P2_U2362, P2_U2398, P2_U4443);
  and ginst11933 (P2_U2363, P2_STATE2_REG_2__SCAN_IN, P2_U3535);
  and ginst11934 (P2_U2364, P2_STATE2_REG_2__SCAN_IN, P2_U3546);
  and ginst11935 (P2_U2365, P2_STATE2_REG_3__SCAN_IN, P2_U4443);
  and ginst11936 (P2_U2366, P2_STATE2_REG_1__SCAN_IN, P2_U3546);
  and ginst11937 (P2_U2367, P2_U2364, P2_U4417);
  and ginst11938 (P2_U2368, P2_U2363, P2_U4420);
  and ginst11939 (P2_U2369, P2_U2364, P2_U4428);
  and ginst11940 (P2_U2370, P2_U2447, P2_U3537);
  and ginst11941 (P2_U2371, P2_U3537, P2_U3990);
  and ginst11942 (P2_U2372, P2_U3537, P2_U3989);
  and ginst11943 (P2_U2373, P2_U3537, P2_U4419);
  and ginst11944 (P2_U2374, P2_STATE2_REG_0__SCAN_IN, P2_U4468);
  and ginst11945 (P2_U2375, P2_U3521, P2_U4441);
  and ginst11946 (P2_U2376, P2_U2436, P2_U3873);
  and ginst11947 (P2_U2377, P2_U2367, P2_U4411);
  and ginst11948 (P2_U2378, P2_STATE2_REG_3__SCAN_IN, P2_U3546);
  and ginst11949 (P2_U2379, P2_U4440, P2_U7865);
  and ginst11950 (P2_U2380, P2_U4441, P2_U7865);
  and ginst11951 (P2_U2381, P2_U3270, P2_U3535);
  and ginst11952 (P2_U2382, P2_U2366, P2_U3647);
  and ginst11953 (P2_U2383, P2_U2366, P2_U3528);
  and ginst11954 (P2_U2384, P2_U2368, P2_U4417);
  and ginst11955 (P2_U2385, P2_U2368, P2_U4428);
  and ginst11956 (P2_U2386, P2_U2363, P2_U4436);
  and ginst11957 (P2_U2387, P2_U3537, P2_U5940);
  and ginst11958 (P2_U2388, P2_U2363, P2_U5675);
  and ginst11959 (P2_U2389, P2_U2363, P2_U5677);
  and ginst11960 (P2_U2390, P2_U2363, P2_U5679);
  and ginst11961 (P2_U2391, P2_U2369, P2_U3545);
  and ginst11962 (P2_U2392, P2_U2369, P2_U6571);
  and ginst11963 (P2_U2393, P2_U3521, P2_U4440);
  and ginst11964 (P2_U2394, P2_U2616, P2_U4442);
  and ginst11965 (P2_U2395, P2_U4442, P2_U7873);
  and ginst11966 (P2_U2396, P2_U3284, P2_U3541);
  and ginst11967 (P2_U2397, P2_U4441, P2_U4601);
  and ginst11968 (P2_U2398, P2_STATEBS16_REG_SCAN_IN, P2_U4430);
  and ginst11969 (P2_U2399, P2_U4443, U314);
  and ginst11970 (P2_U2400, P2_U4443, U303);
  and ginst11971 (P2_U2401, P2_U4443, U292);
  and ginst11972 (P2_U2402, P2_U4443, U289);
  and ginst11973 (P2_U2403, P2_U4443, U288);
  and ginst11974 (P2_U2404, P2_U4443, U287);
  and ginst11975 (P2_U2405, P2_U4443, U286);
  and ginst11976 (P2_U2406, P2_U4443, U285);
  and ginst11977 (P2_U2407, P2_U2362, U298);
  and ginst11978 (P2_U2408, P2_U2362, U307);
  and ginst11979 (P2_U2409, P2_U2362, U297);
  and ginst11980 (P2_U2410, P2_U2362, U306);
  and ginst11981 (P2_U2411, P2_U2362, U296);
  and ginst11982 (P2_U2412, P2_U2362, U305);
  and ginst11983 (P2_U2413, P2_U2362, U295);
  and ginst11984 (P2_U2414, P2_U2362, U304);
  and ginst11985 (P2_U2415, P2_U2362, U294);
  and ginst11986 (P2_U2416, P2_U2362, U302);
  and ginst11987 (P2_U2417, P2_U2362, U293);
  and ginst11988 (P2_U2418, P2_U2362, U301);
  and ginst11989 (P2_U2419, P2_U2362, U291);
  and ginst11990 (P2_U2420, P2_U2362, U300);
  and ginst11991 (P2_U2421, P2_U2362, U290);
  and ginst11992 (P2_U2422, P2_U2362, U299);
  and ginst11993 (P2_U2423, P2_U2365, P2_U3255);
  and ginst11994 (P2_U2424, P2_U2365, P2_U3278);
  and ginst11995 (P2_U2425, P2_U2365, P2_U3521);
  and ginst11996 (P2_U2426, P2_U2365, P2_U3279);
  and ginst11997 (P2_U2427, P2_U2375, P2_U3279);
  and ginst11998 (P2_U2428, P2_U2365, P2_U2616);
  and ginst11999 (P2_U2429, P2_U2365, P2_U2617);
  and ginst12000 (P2_U2430, P2_STATE2_REG_0__SCAN_IN, P2_U3541);
  and ginst12001 (P2_U2431, P2_U2365, P2_U3253);
  and ginst12002 (P2_U2432, P2_U2365, P2_U3280);
  and ginst12003 (P2_U2433, P2_U2375, P2_U3295);
  and ginst12004 (P2_U2434, P2_U2375, P2_U7869);
  and ginst12005 (P2_U2435, P2_U2356, P2_U3541);
  and ginst12006 (P2_U2436, P2_U7859, P2_U7867);
  and ginst12007 (P2_U2437, P2_U2364, P2_U7871);
  and ginst12008 (P2_U2438, P2_U3278, P2_U7859);
  and ginst12009 (P2_U2439, P2_U3521, P2_U4339);
  and ginst12010 (P2_U2440, P2_U3428, P2_U3580);
  and ginst12011 (P2_U2441, P2_U3580, P2_U4647);
  and ginst12012 (P2_U2442, P2_U3428, P2_U8067);
  and ginst12013 (P2_U2443, P2_U4647, P2_U8067);
  and ginst12014 (P2_U2444, P2_U3243, P2_U3307);
  and ginst12015 (P2_U2445, P2_U3307, P2_U4650);
  and ginst12016 (P2_U2446, P2_R2088_U6, P2_U4424);
  and ginst12017 (P2_U2447, P2_STATE2_REG_0__SCAN_IN, P2_U2616);
  and ginst12018 (P2_U2448, P2_STATE2_REG_2__SCAN_IN, P2_STATE2_REG_1__SCAN_IN);
  and ginst12019 (P2_U2449, P2_U3278, P2_U3521);
  and ginst12020 (P2_U2450, P2_U2354, P2_U7871);
  and ginst12021 (P2_U2451, P2_U2438, P2_U2457, P2_U4601);
  and ginst12022 (P2_U2452, P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P2_U3272);
  and ginst12023 (P2_U2453, P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN, P2_U3271);
  and ginst12024 (P2_U2454, P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN, P2_U3271, P2_U3272);
  and ginst12025 (P2_U2455, P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P2_U3272, P2_U3276);
  and ginst12026 (P2_U2456, P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN, P2_U3271, P2_U3276);
  and ginst12027 (P2_U2457, P2_U3255, P2_U3521);
  and ginst12028 (P2_U2458, P2_U2617, P2_U3279, P2_U7863);
  and ginst12029 (P2_U2459, P2_U4393, P2_U8052, P2_U8053);
  and ginst12030 (P2_U2460, P2_R2182_U40, P2_U3317);
  and ginst12031 (P2_U2461, P2_U3426, P2_U3579);
  and ginst12032 (P2_U2462, P2_R2182_U40, P2_R2182_U76);
  and ginst12033 (P2_U2463, P2_U2462, P2_U4637);
  and ginst12034 (P2_U2464, P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN, P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN);
  and ginst12035 (P2_U2465, P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN, P2_U3309);
  and ginst12036 (P2_U2466, P2_R2099_U95, P2_R2099_U96);
  and ginst12037 (P2_U2467, P2_R2099_U5, P2_R2099_U94);
  and ginst12038 (P2_U2468, P2_U3320, P2_U4657);
  and ginst12039 (P2_U2469, P2_U2462, P2_U4633);
  and ginst12040 (P2_U2470, P2_R2099_U5, P2_U3323);
  and ginst12041 (P2_U2471, P2_U3339, P2_U4715);
  and ginst12042 (P2_U2472, P2_U2462, P2_U4634);
  and ginst12043 (P2_U2473, P2_R2099_U94, P2_U3324);
  and ginst12044 (P2_U2474, P2_U3354, P2_U4774);
  and ginst12045 (P2_U2475, P2_R2182_U69, P2_U4635);
  nor ginst12046 (P2_U2476, P2_R2182_U68, P2_R2182_U69);
  and ginst12047 (P2_U2477, P2_U2462, P2_U2476);
  nor ginst12048 (P2_U2478, P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN, P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN);
  nor ginst12049 (P2_U2479, P2_R2099_U5, P2_R2099_U94);
  and ginst12050 (P2_U2480, P2_U3366, P2_U4831);
  and ginst12051 (P2_U2481, P2_U3426, P2_U8064);
  and ginst12052 (P2_U2482, P2_U4637, P2_U4638);
  and ginst12053 (P2_U2483, P2_R2099_U95, P2_U3322);
  and ginst12054 (P2_U2484, P2_U3379, P2_U4889);
  and ginst12055 (P2_U2485, P2_U4633, P2_U4638);
  and ginst12056 (P2_U2486, P2_U3391, P2_U4946);
  and ginst12057 (P2_U2487, P2_U4634, P2_U4638);
  and ginst12058 (P2_U2488, P2_U3402, P2_U5004);
  and ginst12059 (P2_U2489, P2_U2476, P2_U4638);
  and ginst12060 (P2_U2490, P2_U3414, P2_U5061);
  and ginst12061 (P2_U2491, P2_U3579, P2_U4640);
  and ginst12062 (P2_U2492, P2_R2099_U96, P2_U3321);
  and ginst12063 (P2_U2493, P2_U3425, P2_U3427);
  and ginst12064 (P2_U2494, P2_U2460, P2_U4633);
  and ginst12065 (P2_U2495, P2_U3440, P2_U5174);
  and ginst12066 (P2_U2496, P2_U2460, P2_U4634);
  and ginst12067 (P2_U2497, P2_U3451, P2_U5232);
  and ginst12068 (P2_U2498, P2_U2460, P2_U2476);
  and ginst12069 (P2_U2499, P2_U3463, P2_U5289);
  and ginst12070 (P2_U2500, P2_U4640, P2_U8064);
  nor ginst12071 (P2_U2501, P2_R2182_U40, P2_R2182_U76);
  and ginst12072 (P2_U2502, P2_U2501, P2_U4637);
  nor ginst12073 (P2_U2503, P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN, P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN);
  nor ginst12074 (P2_U2504, P2_R2099_U95, P2_R2099_U96);
  and ginst12075 (P2_U2505, P2_U3474, P2_U5347);
  and ginst12076 (P2_U2506, P2_U2501, P2_U4633);
  and ginst12077 (P2_U2507, P2_U3486, P2_U5404);
  and ginst12078 (P2_U2508, P2_U2501, P2_U4634);
  and ginst12079 (P2_U2509, P2_U3497, P2_U5462);
  and ginst12080 (P2_U2510, P2_U2476, P2_U2501);
  and ginst12081 (P2_U2511, P2_U3509, P2_U5519);
  and ginst12082 (P2_U2512, P2_U3869, P2_U8068, P2_U8069);
  and ginst12083 (P2_U2513, P2_U5579, P2_U5580);
  and ginst12084 (P2_U2514, P2_U3881, P2_U3882, P2_U7896);
  and ginst12085 (P2_U2515, P2_U8082, P2_U8100);
  and ginst12086 (P2_U2516, P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN, P2_U5616);
  and ginst12087 (P2_U2517, P2_U2515, P2_U2516);
  and ginst12088 (P2_U2518, P2_U3272, P2_U5616);
  and ginst12089 (P2_U2519, P2_U2515, P2_U2518);
  and ginst12090 (P2_U2520, P2_U3582, P2_U8082);
  and ginst12091 (P2_U2521, P2_U2516, P2_U2520);
  and ginst12092 (P2_U2522, P2_U2518, P2_U2520);
  and ginst12093 (P2_U2523, P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN, P2_U3530);
  and ginst12094 (P2_U2524, P2_U2515, P2_U2523);
  and ginst12095 (P2_U2525, P2_U3272, P2_U3530);
  and ginst12096 (P2_U2526, P2_U2515, P2_U2525);
  and ginst12097 (P2_U2527, P2_U2520, P2_U2523);
  and ginst12098 (P2_U2528, P2_U2520, P2_U2525);
  and ginst12099 (P2_U2529, P2_U3581, P2_U3582);
  and ginst12100 (P2_U2530, P2_U2525, P2_U2529);
  and ginst12101 (P2_U2531, P2_U2523, P2_U2529);
  and ginst12102 (P2_U2532, P2_U3581, P2_U8100);
  and ginst12103 (P2_U2533, P2_U2525, P2_U2532);
  and ginst12104 (P2_U2534, P2_U2523, P2_U2532);
  and ginst12105 (P2_U2535, P2_U2518, P2_U2529);
  and ginst12106 (P2_U2536, P2_U2516, P2_U2529);
  and ginst12107 (P2_U2537, P2_U2518, P2_U2532);
  and ginst12108 (P2_U2538, P2_U2516, P2_U2532);
  nor ginst12109 (P2_U2539, P2_R2147_U4, P2_R2147_U8);
  nor ginst12110 (P2_U2540, P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN, P2_R2147_U9);
  and ginst12111 (P2_U2541, P2_U2539, P2_U2540);
  and ginst12112 (P2_U2542, P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN, P2_U3529);
  and ginst12113 (P2_U2543, P2_U2539, P2_U2542);
  and ginst12114 (P2_U2544, P2_R2147_U4, P2_U3526);
  and ginst12115 (P2_U2545, P2_U2540, P2_U2544);
  and ginst12116 (P2_U2546, P2_U2542, P2_U2544);
  and ginst12117 (P2_U2547, P2_R2147_U9, P2_U3532);
  and ginst12118 (P2_U2548, P2_U2539, P2_U2547);
  and ginst12119 (P2_U2549, P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN, P2_R2147_U9);
  and ginst12120 (P2_U2550, P2_U2539, P2_U2549);
  and ginst12121 (P2_U2551, P2_U2544, P2_U2547);
  and ginst12122 (P2_U2552, P2_U2544, P2_U2549);
  and ginst12123 (P2_U2553, P2_R2147_U8, P2_U3531);
  and ginst12124 (P2_U2554, P2_U2540, P2_U2553);
  and ginst12125 (P2_U2555, P2_U2542, P2_U2553);
  and ginst12126 (P2_U2556, P2_R2147_U4, P2_R2147_U8);
  and ginst12127 (P2_U2557, P2_U2540, P2_U2556);
  and ginst12128 (P2_U2558, P2_U2542, P2_U2556);
  and ginst12129 (P2_U2559, P2_U2547, P2_U2553);
  and ginst12130 (P2_U2560, P2_U2549, P2_U2553);
  and ginst12131 (P2_U2561, P2_U2547, P2_U2556);
  and ginst12132 (P2_U2562, P2_U2549, P2_U2556);
  and ginst12133 (P2_U2563, P2_U3272, P2_U8100);
  and ginst12134 (P2_U2564, P2_U3583, P2_U4409);
  and ginst12135 (P2_U2565, P2_U2563, P2_U2564);
  and ginst12136 (P2_U2566, P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN, P2_U8100);
  and ginst12137 (P2_U2567, P2_U2564, P2_U2566);
  and ginst12138 (P2_U2568, P2_U3272, P2_U3582);
  and ginst12139 (P2_U2569, P2_U2564, P2_U2568);
  and ginst12140 (P2_U2570, P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN, P2_U3582);
  and ginst12141 (P2_U2571, P2_U2564, P2_U2570);
  and ginst12142 (P2_U2572, P2_U3553, P2_U3583);
  and ginst12143 (P2_U2573, P2_U2563, P2_U2572);
  and ginst12144 (P2_U2574, P2_U2566, P2_U2572);
  and ginst12145 (P2_U2575, P2_U2568, P2_U2572);
  and ginst12146 (P2_U2576, P2_U2570, P2_U2572);
  and ginst12147 (P2_U2577, P2_U4409, P2_U8149);
  and ginst12148 (P2_U2578, P2_U2563, P2_U2577);
  and ginst12149 (P2_U2579, P2_U2566, P2_U2577);
  and ginst12150 (P2_U2580, P2_U2568, P2_U2577);
  and ginst12151 (P2_U2581, P2_U2570, P2_U2577);
  and ginst12152 (P2_U2582, P2_U3553, P2_U8149);
  and ginst12153 (P2_U2583, P2_U2563, P2_U2582);
  and ginst12154 (P2_U2584, P2_U2566, P2_U2582);
  and ginst12155 (P2_U2585, P2_U2568, P2_U2582);
  and ginst12156 (P2_U2586, P2_U2570, P2_U2582);
  and ginst12157 (P2_U2587, P2_EBX_REG_31__SCAN_IN, P2_U2391);
  and ginst12158 (P2_U2588, P2_U2360, P2_U2377);
  and ginst12159 (P2_U2589, P2_U3549, P2_U3550, P2_U4457, P2_U7581);
  and ginst12160 (P2_U2590, P2_U2436, P2_U5590);
  nand ginst12161 (P2_U2591, P2_U4273, P2_U4274);
  nand ginst12162 (P2_U2592, P2_U4271, P2_U4272);
  nand ginst12163 (P2_U2593, P2_U4269, P2_U4270);
  nand ginst12164 (P2_U2594, P2_U4267, P2_U4268);
  nand ginst12165 (P2_U2595, P2_U4265, P2_U4266);
  nand ginst12166 (P2_U2596, P2_U4263, P2_U4264);
  nand ginst12167 (P2_U2597, P2_U4261, P2_U4262);
  nand ginst12168 (P2_U2598, P2_U4259, P2_U4260);
  nand ginst12169 (P2_U2599, P2_U4255, P2_U4256, P2_U4257, P2_U4258);
  nand ginst12170 (P2_U2600, P2_U4251, P2_U4252, P2_U4253, P2_U4254);
  nand ginst12171 (P2_U2601, P2_U4247, P2_U4248, P2_U4249, P2_U4250);
  nand ginst12172 (P2_U2602, P2_U4243, P2_U4244, P2_U4245, P2_U4246);
  nand ginst12173 (P2_U2603, P2_U4239, P2_U4240, P2_U4241, P2_U4242);
  nand ginst12174 (P2_U2604, P2_U4235, P2_U4236, P2_U4237, P2_U4238);
  nand ginst12175 (P2_U2605, P2_U4231, P2_U4232, P2_U4233, P2_U4234);
  nand ginst12176 (P2_U2606, P2_U4227, P2_U4228, P2_U4229, P2_U4230);
  nand ginst12177 (P2_U2607, P2_U4223, P2_U4224, P2_U4225, P2_U4226);
  nand ginst12178 (P2_U2608, P2_U4219, P2_U4220, P2_U4221, P2_U4222);
  nand ginst12179 (P2_U2609, P2_U4215, P2_U4216, P2_U4217, P2_U4218);
  nand ginst12180 (P2_U2610, P2_U4211, P2_U4212, P2_U4213, P2_U4214);
  nand ginst12181 (P2_U2611, P2_U4207, P2_U4208, P2_U4209, P2_U4210);
  nand ginst12182 (P2_U2612, P2_U4203, P2_U4204, P2_U4205, P2_U4206);
  nand ginst12183 (P2_U2613, P2_U4199, P2_U4200, P2_U4201, P2_U4202);
  nand ginst12184 (P2_U2614, P2_U4195, P2_U4196, P2_U4197, P2_U4198);
  and ginst12185 (P2_U2615, P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN, P2_U3519);
  nand ginst12186 (P2_U2616, P2_U3705, P2_U3706);
  nand ginst12187 (P2_U2617, P2_U3693, P2_U3694);
  nand ginst12188 (P2_U2618, P2_U4350, P2_U7453);
  nand ginst12189 (P2_U2619, P2_U4351, P2_U7456);
  nand ginst12190 (P2_U2620, P2_U4353, P2_U7462);
  nand ginst12191 (P2_U2621, P2_U4354, P2_U7465);
  nand ginst12192 (P2_U2622, P2_U4355, P2_U7468);
  nand ginst12193 (P2_U2623, P2_U4356, P2_U7471);
  nand ginst12194 (P2_U2624, P2_U4357, P2_U7474);
  nand ginst12195 (P2_U2625, P2_U4358, P2_U7477);
  nand ginst12196 (P2_U2626, P2_U4359, P2_U7480);
  nand ginst12197 (P2_U2627, P2_U4360, P2_U7483);
  nand ginst12198 (P2_U2628, P2_U4361, P2_U7486);
  nand ginst12199 (P2_U2629, P2_U4362, P2_U7489);
  nand ginst12200 (P2_U2630, P2_U4364, P2_U7495);
  nand ginst12201 (P2_U2631, P2_U4365, P2_U7498);
  nand ginst12202 (P2_U2632, P2_U4366, P2_U7501);
  nand ginst12203 (P2_U2633, P2_U4367, P2_U7504);
  nand ginst12204 (P2_U2634, P2_U4368, P2_U7507, P2_U7508);
  nand ginst12205 (P2_U2635, P2_U4369, P2_U7511, P2_U7512);
  nand ginst12206 (P2_U2636, P2_U4370, P2_U7515, P2_U7516);
  nand ginst12207 (P2_U2637, P2_U4371, P2_U7519, P2_U7520);
  nand ginst12208 (P2_U2638, P2_U4372, P2_U7523, P2_U7524);
  nand ginst12209 (P2_U2639, P2_U4373, P2_U7527, P2_U7528);
  nand ginst12210 (P2_U2640, P2_U4344, P2_U7433, P2_U7434);
  nand ginst12211 (P2_U2641, P2_U4345, P2_U7437, P2_U7438);
  nand ginst12212 (P2_U2642, P2_U4346, P2_U7441);
  nand ginst12213 (P2_U2643, P2_U4347, P2_U7444);
  nand ginst12214 (P2_U2644, P2_U4348, P2_U7447);
  nand ginst12215 (P2_U2645, P2_U4349, P2_U7450);
  nand ginst12216 (P2_U2646, P2_U4352, P2_U7459);
  nand ginst12217 (P2_U2647, P2_U4363, P2_U7492);
  nand ginst12218 (P2_U2648, P2_U4374, P2_U7531);
  nand ginst12219 (P2_U2649, P2_U3300, P2_U4375, P2_U7534);
  and ginst12220 (P2_U2650, P2_U2352, P2_U3242);
  and ginst12221 (P2_U2651, P2_U2352, P2_U7217);
  and ginst12222 (P2_U2652, P2_U2352, P2_U7251);
  and ginst12223 (P2_U2653, P2_U2352, P2_U7285);
  nand ginst12224 (P2_U2654, P2_U7422, P2_U7423);
  nand ginst12225 (P2_U2655, P2_U4338, P2_U7424);
  nand ginst12226 (P2_U2656, P2_U4340, P2_U7427);
  nand ginst12227 (P2_U2657, P2_U4342, P2_U7429);
  and ginst12228 (P2_U2658, P2_U2354, P2_U2598);
  and ginst12229 (P2_U2659, P2_U2354, P2_U2597);
  and ginst12230 (P2_U2660, P2_U2354, P2_U2596);
  and ginst12231 (P2_U2661, P2_U2354, P2_U2595);
  and ginst12232 (P2_U2662, P2_U2354, P2_U2594);
  and ginst12233 (P2_U2663, P2_U2354, P2_U2593);
  and ginst12234 (P2_U2664, P2_U2354, P2_U2592);
  and ginst12235 (P2_U2665, P2_U2354, P2_U2591);
  and ginst12236 (P2_U2666, P2_U2355, P2_U2614);
  and ginst12237 (P2_U2667, P2_U2355, P2_U2613);
  and ginst12238 (P2_U2668, P2_U2355, P2_U2612);
  and ginst12239 (P2_U2669, P2_U2355, P2_U2611);
  and ginst12240 (P2_U2670, P2_U2355, P2_U2610);
  and ginst12241 (P2_U2671, P2_U2355, P2_U2609);
  and ginst12242 (P2_U2672, P2_U2355, P2_U2608);
  and ginst12243 (P2_U2673, P2_U2355, P2_U2607);
  and ginst12244 (P2_U2674, P2_INSTQUEUE_REG_0__7__SCAN_IN, P2_U2355);
  and ginst12245 (P2_U2675, P2_INSTQUEUE_REG_0__6__SCAN_IN, P2_U2355);
  and ginst12246 (P2_U2676, P2_INSTQUEUE_REG_0__5__SCAN_IN, P2_U2355);
  and ginst12247 (P2_U2677, P2_INSTQUEUE_REG_0__4__SCAN_IN, P2_U2355);
  and ginst12248 (P2_U2678, P2_INSTQUEUE_REG_0__3__SCAN_IN, P2_U2355);
  and ginst12249 (P2_U2679, P2_INSTQUEUE_REG_0__2__SCAN_IN, P2_U2355);
  and ginst12250 (P2_U2680, P2_INSTQUEUE_REG_0__1__SCAN_IN, P2_U2355);
  nand ginst12251 (P2_U2681, P2_U4275, P2_U7166);
  and ginst12252 (P2_U2682, P2_ADD_402_1132_U18, P2_U2355);
  and ginst12253 (P2_U2683, P2_ADD_402_1132_U19, P2_U2355);
  and ginst12254 (P2_U2684, P2_ADD_402_1132_U24, P2_U2355);
  and ginst12255 (P2_U2685, P2_ADD_402_1132_U22, P2_U2355);
  and ginst12256 (P2_U2686, P2_ADD_402_1132_U21, P2_U2355);
  and ginst12257 (P2_U2687, P2_ADD_402_1132_U25, P2_U2355);
  and ginst12258 (P2_U2688, P2_ADD_402_1132_U20, P2_U2355);
  nand ginst12259 (P2_U2689, P2_U7141, P2_U7142);
  nand ginst12260 (P2_U2690, P2_U7143, P2_U7144);
  nand ginst12261 (P2_U2691, P2_U7145, P2_U7146);
  nand ginst12262 (P2_U2692, P2_U7147, P2_U7148);
  nand ginst12263 (P2_U2693, P2_U7152, P2_U7153);
  nand ginst12264 (P2_U2694, P2_U7154, P2_U7155);
  nand ginst12265 (P2_U2695, P2_U7156, P2_U7157);
  nand ginst12266 (P2_U2696, P2_U7158, P2_U7159);
  and ginst12267 (P2_U2698, P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN, P2_U3554);
  nand ginst12268 (P2_U2699, P2_U7138, P2_U7139, P2_U7140);
  nand ginst12269 (P2_U2700, P2_U7149, P2_U7150, P2_U7151);
  nand ginst12270 (P2_U2701, P2_U7160, P2_U7161, P2_U7162);
  nand ginst12271 (P2_U2702, P2_U7163, P2_U7164, P2_U7165);
  nand ginst12272 (P2_U2703, P2_U7726, P2_U7727);
  nand ginst12273 (P2_U2704, P2_U7728, P2_U7729);
  nand ginst12274 (P2_U2705, P2_U4390, P2_U7730);
  nand ginst12275 (P2_U2706, P2_U3550, P2_U7732, P2_U7733);
  nand ginst12276 (P2_U2707, P2_U4391, P2_U7734);
  and ginst12277 (P2_U2708, P2_R2219_U25, P2_U7723);
  and ginst12278 (P2_U2709, P2_R2219_U26, P2_U7723);
  and ginst12279 (P2_U2710, P2_R2219_U27, P2_U7723);
  nand ginst12280 (P2_U2711, P2_STATE2_REG_0__SCAN_IN, P2_U7724);
  nand ginst12281 (P2_U2712, P2_STATE2_REG_0__SCAN_IN, P2_U4407, P2_U7871);
  nand ginst12282 (P2_U2713, P2_STATE2_REG_0__SCAN_IN, P2_U7725);
  nand ginst12283 (P2_U2714, P2_STATE2_REG_0__SCAN_IN, P2_U4408, P2_U7871);
  nand ginst12284 (P2_U2715, P2_U2356, P2_U2616);
  nand ginst12285 (P2_U2716, P2_U7617, P2_U7618, P2_U7619, P2_U7620);
  nand ginst12286 (P2_U2717, P2_U7621, P2_U7622, P2_U7623, P2_U7624);
  nand ginst12287 (P2_U2718, P2_U7629, P2_U7630, P2_U7631, P2_U7632);
  nand ginst12288 (P2_U2719, P2_U7633, P2_U7634, P2_U7635, P2_U7636);
  nand ginst12289 (P2_U2720, P2_U7637, P2_U7638, P2_U7639, P2_U7640);
  nand ginst12290 (P2_U2721, P2_U7641, P2_U7642, P2_U7643, P2_U7644);
  nand ginst12291 (P2_U2722, P2_U7645, P2_U7646, P2_U7647, P2_U7648);
  nand ginst12292 (P2_U2723, P2_U7649, P2_U7650, P2_U7651, P2_U7652);
  nand ginst12293 (P2_U2724, P2_U7653, P2_U7654, P2_U7655, P2_U7656);
  nand ginst12294 (P2_U2725, P2_U7657, P2_U7658, P2_U7659, P2_U7660);
  nand ginst12295 (P2_U2726, P2_U7661, P2_U7662, P2_U7663, P2_U7664);
  nand ginst12296 (P2_U2727, P2_U7665, P2_U7666, P2_U7667, P2_U7668);
  nand ginst12297 (P2_U2728, P2_U7673, P2_U7674, P2_U7675, P2_U7676);
  nand ginst12298 (P2_U2729, P2_U7677, P2_U7678, P2_U7679, P2_U7680);
  nand ginst12299 (P2_U2730, P2_U7681, P2_U7682, P2_U7683, P2_U7684);
  nand ginst12300 (P2_U2731, P2_U7685, P2_U7686, P2_U7687, P2_U7688);
  nand ginst12301 (P2_U2732, P2_U7689, P2_U7690, P2_U7691, P2_U7692);
  nand ginst12302 (P2_U2733, P2_U7693, P2_U7694, P2_U7695, P2_U7696);
  nand ginst12303 (P2_U2734, P2_U7697, P2_U7698, P2_U7699, P2_U7700);
  nand ginst12304 (P2_U2735, P2_U7701, P2_U7702, P2_U7703, P2_U7704);
  nand ginst12305 (P2_U2736, P2_U7705, P2_U7706, P2_U7707, P2_U7708);
  nand ginst12306 (P2_U2737, P2_U7709, P2_U7710, P2_U7711, P2_U7712);
  nand ginst12307 (P2_U2738, P2_U7593, P2_U7594, P2_U7595, P2_U7596);
  nand ginst12308 (P2_U2739, P2_U7597, P2_U7598, P2_U7599, P2_U7600);
  nand ginst12309 (P2_U2740, P2_U7601, P2_U7602, P2_U7603, P2_U7604);
  nand ginst12310 (P2_U2741, P2_U7605, P2_U7606, P2_U7607, P2_U7608);
  nand ginst12311 (P2_U2742, P2_U7609, P2_U7610, P2_U7611, P2_U7612);
  nand ginst12312 (P2_U2743, P2_U7613, P2_U7614, P2_U7615, P2_U7616);
  nand ginst12313 (P2_U2744, P2_U7625, P2_U7626, P2_U7627, P2_U7628);
  nand ginst12314 (P2_U2745, P2_U7669, P2_U7670, P2_U7671, P2_U7672);
  nand ginst12315 (P2_U2746, P2_U7713, P2_U7714, P2_U7715, P2_U7716);
  nand ginst12316 (P2_U2747, P2_U4388, P2_U4389, P2_U7717, P2_U7721, P2_U7886);
  nand ginst12317 (P2_U2748, P2_U7582, P2_U7583);
  nand ginst12318 (P2_U2749, P2_U4380, P2_U7584);
  nand ginst12319 (P2_U2750, P2_U4382, P2_U7588);
  and ginst12320 (P2_U2751, P2_U7737, P2_U7888);
  and ginst12321 (P2_U2752, P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN, P2_U3280, P2_U7873);
  nand ginst12322 (P2_U2753, P2_U3286, P2_U7572);
  nand ginst12323 (P2_U2754, P2_U3286, P2_U7573);
  nand ginst12324 (P2_U2755, P2_U3286, P2_U7574);
  nand ginst12325 (P2_U2756, P2_U3286, P2_U7575);
  nand ginst12326 (P2_U2757, P2_U3286, P2_U7576);
  and ginst12327 (P2_U2758, P2_U3242, P2_U4428);
  and ginst12328 (P2_U2759, P2_U4428, P2_U7217);
  and ginst12329 (P2_U2760, P2_U4428, P2_U7251);
  nand ginst12330 (P2_U2761, P2_U7562, P2_U7563);
  nand ginst12331 (P2_U2762, P2_U7564, P2_U7565);
  nand ginst12332 (P2_U2763, P2_U7566, P2_U7567);
  nand ginst12333 (P2_U2764, P2_U7568, P2_U7569);
  nand ginst12334 (P2_U2765, P2_U7570, P2_U7571);
  nand ginst12335 (P2_U2766, P2_U4447, P2_U7539);
  nand ginst12336 (P2_U2767, P2_U4447, P2_U7540);
  nand ginst12337 (P2_U2768, P2_U4447, P2_U7541);
  nand ginst12338 (P2_U2769, P2_U4447, P2_U7542);
  nand ginst12339 (P2_U2770, P2_U4447, P2_U7543);
  nand ginst12340 (P2_U2771, P2_U4447, P2_U7544);
  nand ginst12341 (P2_U2772, P2_U4447, P2_U7545);
  nand ginst12342 (P2_U2773, P2_U4447, P2_U7546);
  nand ginst12343 (P2_U2774, P2_U4447, P2_U7547);
  nand ginst12344 (P2_U2775, P2_U4447, P2_U7548);
  nand ginst12345 (P2_U2776, P2_U4447, P2_U7549);
  nand ginst12346 (P2_U2777, P2_U4447, P2_U7550);
  nand ginst12347 (P2_U2778, P2_U4447, P2_U7551);
  nand ginst12348 (P2_U2779, P2_U4447, P2_U7552);
  nand ginst12349 (P2_U2780, P2_U4447, P2_U7553);
  nand ginst12350 (P2_U2781, P2_U4447, P2_U7554);
  nand ginst12351 (P2_U2782, P2_U4447, P2_U7555);
  nand ginst12352 (P2_U2783, P2_U4447, P2_U7556);
  nand ginst12353 (P2_U2784, P2_U4447, P2_U7557);
  nand ginst12354 (P2_U2785, P2_U4447, P2_U7558);
  nand ginst12355 (P2_U2786, P2_U4447, P2_U7559);
  nand ginst12356 (P2_U2787, P2_U4447, P2_U7560);
  nand ginst12357 (P2_U2788, P2_U4447, P2_U7537);
  nand ginst12358 (P2_U2789, P2_U4447, P2_U7538);
  and ginst12359 (P2_U2790, P2_R2267_U63, P2_U3242);
  and ginst12360 (P2_U2791, P2_R2267_U16, P2_U3242);
  and ginst12361 (P2_U2792, P2_R2267_U15, P2_U3242);
  and ginst12362 (P2_U2793, P2_R2267_U67, P2_U3242);
  and ginst12363 (P2_U2794, P2_R2267_U14, P2_U3242);
  and ginst12364 (P2_U2795, P2_R2267_U69, P2_U3242);
  and ginst12365 (P2_U2796, P2_R2267_U13, P2_U3242);
  and ginst12366 (P2_U2797, P2_R2267_U71, P2_U3242);
  and ginst12367 (P2_U2798, P2_R2267_U12, P2_U3242);
  and ginst12368 (P2_U2799, P2_R2267_U73, P2_U3242);
  and ginst12369 (P2_U2800, P2_R2267_U11, P2_U3242);
  and ginst12370 (P2_U2801, P2_R2267_U75, P2_U3242);
  and ginst12371 (P2_U2802, P2_R2267_U10, P2_U3242);
  and ginst12372 (P2_U2803, P2_R2267_U79, P2_U3242);
  and ginst12373 (P2_U2804, P2_R2267_U9, P2_U3242);
  and ginst12374 (P2_U2805, P2_R2267_U81, P2_U3242);
  and ginst12375 (P2_U2806, P2_R2267_U8, P2_U3242);
  and ginst12376 (P2_U2807, P2_R2267_U83, P2_U3242);
  and ginst12377 (P2_U2808, P2_R2267_U7, P2_U3242);
  and ginst12378 (P2_U2809, P2_R2267_U85, P2_U3242);
  and ginst12379 (P2_U2810, P2_R2267_U6, P2_U3242);
  and ginst12380 (P2_U2811, P2_R2267_U87, P2_U3242);
  and ginst12381 (P2_U2812, P2_R2267_U20, P2_U3242);
  and ginst12382 (P2_U2813, P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P2_U3519);
  nand ginst12383 (P2_U2814, P2_U4190, P2_U6861);
  nand ginst12384 (P2_U2815, P2_U6856, P2_U7917);
  nand ginst12385 (P2_U2816, P2_U6854, P2_U6855);
  nand ginst12386 (P2_U2817, P2_U4463, P2_U8139, P2_U8140);
  nand ginst12387 (P2_U2818, P2_U4463, P2_U8135, P2_U8136);
  nand ginst12388 (P2_U2819, P2_U6839, P2_U6840);
  nand ginst12389 (P2_U2820, P2_U3548, P2_U8127, P2_U8128);
  nand ginst12390 (P2_U2821, P2_U3548, P2_U4452, P2_U6837);
  nand ginst12391 (P2_U2822, P2_U4398, P2_U6836);
  nand ginst12392 (P2_U2823, P2_U4452, P2_U8123, P2_U8124);
  nand ginst12393 (P2_U2824, P2_U4168, P2_U6827, P2_U6828, P2_U6829, P2_U6830);
  nand ginst12394 (P2_U2825, P2_U4166, P2_U6819, P2_U6820, P2_U6821, P2_U6822);
  nand ginst12395 (P2_U2826, P2_U4164, P2_U6811, P2_U6812, P2_U6813, P2_U6814);
  nand ginst12396 (P2_U2827, P2_U4162, P2_U6803, P2_U6804, P2_U6805, P2_U6806);
  nand ginst12397 (P2_U2828, P2_U4160, P2_U6795, P2_U6796, P2_U6797, P2_U6798);
  nand ginst12398 (P2_U2829, P2_U4158, P2_U6787, P2_U6788, P2_U6789, P2_U6790);
  nand ginst12399 (P2_U2830, P2_U4156, P2_U6779, P2_U6780, P2_U6781, P2_U6782);
  nand ginst12400 (P2_U2831, P2_U4152, P2_U6772);
  nand ginst12401 (P2_U2832, P2_U4149, P2_U6764);
  nand ginst12402 (P2_U2833, P2_U4148, P2_U6755, P2_U6756, P2_U6757, P2_U6758);
  nand ginst12403 (P2_U2834, P2_U4144, P2_U4146);
  nand ginst12404 (P2_U2835, P2_U4141, P2_U4143);
  nand ginst12405 (P2_U2836, P2_U4138, P2_U4140);
  nand ginst12406 (P2_U2837, P2_U4134, P2_U4136);
  nand ginst12407 (P2_U2838, P2_U4130, P2_U4132);
  nand ginst12408 (P2_U2839, P2_U4126, P2_U4128);
  nand ginst12409 (P2_U2840, P2_U4122, P2_U4124);
  nand ginst12410 (P2_U2841, P2_U4118, P2_U4119, P2_U6692, P2_U6693, P2_U6696);
  nand ginst12411 (P2_U2842, P2_U4115, P2_U4116, P2_U6684, P2_U6685, P2_U6688);
  nand ginst12412 (P2_U2843, P2_U4112, P2_U4113, P2_U6676, P2_U6677, P2_U6680);
  nand ginst12413 (P2_U2844, P2_U4109, P2_U4110, P2_U6669, P2_U6670, P2_U6672);
  nand ginst12414 (P2_U2845, P2_U4106, P2_U4107, P2_U6661, P2_U6662, P2_U6664);
  nand ginst12415 (P2_U2846, P2_U4103, P2_U4104, P2_U6653, P2_U6654, P2_U6656);
  nand ginst12416 (P2_U2847, P2_U4100, P2_U4101, P2_U6645, P2_U6646, P2_U6648);
  nand ginst12417 (P2_U2848, P2_U4097, P2_U4098, P2_U6637, P2_U6638, P2_U6640);
  nand ginst12418 (P2_U2849, P2_U4094, P2_U4095, P2_U6629, P2_U6630, P2_U6632);
  nand ginst12419 (P2_U2850, P2_U4091, P2_U4093);
  nand ginst12420 (P2_U2851, P2_U4087, P2_U4089);
  nand ginst12421 (P2_U2852, P2_U4082, P2_U4084, P2_U6602, P2_U6606);
  nand ginst12422 (P2_U2853, P2_U4078, P2_U4080, P2_U6593, P2_U6597);
  nand ginst12423 (P2_U2854, P2_U4074, P2_U4076, P2_U6584, P2_U6588);
  nand ginst12424 (P2_U2855, P2_U4070, P2_U4072, P2_U6575, P2_U6579);
  nand ginst12425 (P2_U2856, P2_U6564, P2_U6565);
  nand ginst12426 (P2_U2857, P2_U6561, P2_U6562, P2_U6563);
  nand ginst12427 (P2_U2858, P2_U6558, P2_U6559, P2_U6560);
  nand ginst12428 (P2_U2859, P2_U6555, P2_U6556, P2_U6557);
  nand ginst12429 (P2_U2860, P2_U6552, P2_U6553, P2_U6554);
  nand ginst12430 (P2_U2861, P2_U6549, P2_U6550, P2_U6551);
  nand ginst12431 (P2_U2862, P2_U6546, P2_U6547, P2_U6548);
  nand ginst12432 (P2_U2863, P2_U6543, P2_U6544, P2_U6545);
  nand ginst12433 (P2_U2864, P2_U6540, P2_U6541, P2_U6542);
  nand ginst12434 (P2_U2865, P2_U6537, P2_U6538, P2_U6539);
  nand ginst12435 (P2_U2866, P2_U6534, P2_U6535, P2_U6536);
  nand ginst12436 (P2_U2867, P2_U6531, P2_U6532, P2_U6533);
  nand ginst12437 (P2_U2868, P2_U6528, P2_U6529, P2_U6530);
  nand ginst12438 (P2_U2869, P2_U6525, P2_U6526, P2_U6527);
  nand ginst12439 (P2_U2870, P2_U6522, P2_U6523, P2_U6524);
  nand ginst12440 (P2_U2871, P2_U6519, P2_U6520, P2_U6521);
  nand ginst12441 (P2_U2872, P2_U6516, P2_U6517, P2_U6518);
  nand ginst12442 (P2_U2873, P2_U6513, P2_U6514, P2_U6515);
  nand ginst12443 (P2_U2874, P2_U6510, P2_U6511, P2_U6512);
  nand ginst12444 (P2_U2875, P2_U6507, P2_U6508, P2_U6509);
  nand ginst12445 (P2_U2876, P2_U6504, P2_U6505, P2_U6506);
  nand ginst12446 (P2_U2877, P2_U6501, P2_U6502, P2_U6503);
  nand ginst12447 (P2_U2878, P2_U6498, P2_U6499, P2_U6500);
  nand ginst12448 (P2_U2879, P2_U6495, P2_U6496, P2_U6497);
  nand ginst12449 (P2_U2880, P2_U6492, P2_U6493, P2_U6494);
  nand ginst12450 (P2_U2881, P2_U6489, P2_U6490, P2_U6491);
  nand ginst12451 (P2_U2882, P2_U6486, P2_U6487, P2_U6488);
  nand ginst12452 (P2_U2883, P2_U6483, P2_U6484, P2_U6485);
  nand ginst12453 (P2_U2884, P2_U6480, P2_U6481, P2_U6482);
  nand ginst12454 (P2_U2885, P2_U6477, P2_U6478, P2_U6479);
  nand ginst12455 (P2_U2886, P2_U6474, P2_U6475, P2_U6476);
  nand ginst12456 (P2_U2887, P2_U6471, P2_U6472, P2_U6473);
  nand ginst12457 (P2_U2888, P2_U6466, P2_U6467, P2_U6468);
  nand ginst12458 (P2_U2889, P2_U6461, P2_U6462, P2_U6463, P2_U6464, P2_U6465);
  nand ginst12459 (P2_U2890, P2_U6456, P2_U6457, P2_U6458, P2_U6459, P2_U6460);
  nand ginst12460 (P2_U2891, P2_U6451, P2_U6452, P2_U6453, P2_U6454, P2_U6455);
  nand ginst12461 (P2_U2892, P2_U6446, P2_U6447, P2_U6448, P2_U6449, P2_U6450);
  nand ginst12462 (P2_U2893, P2_U6441, P2_U6442, P2_U6443, P2_U6444, P2_U6445);
  nand ginst12463 (P2_U2894, P2_U6436, P2_U6437, P2_U6438, P2_U6439, P2_U6440);
  nand ginst12464 (P2_U2895, P2_U6431, P2_U6432, P2_U6433, P2_U6434, P2_U6435);
  nand ginst12465 (P2_U2896, P2_U6426, P2_U6427, P2_U6428, P2_U6429, P2_U6430);
  nand ginst12466 (P2_U2897, P2_U6421, P2_U6422, P2_U6423, P2_U6424, P2_U6425);
  nand ginst12467 (P2_U2898, P2_U6416, P2_U6417, P2_U6418, P2_U6419, P2_U6420);
  nand ginst12468 (P2_U2899, P2_U6411, P2_U6412, P2_U6413, P2_U6414, P2_U6415);
  nand ginst12469 (P2_U2900, P2_U6406, P2_U6407, P2_U6408, P2_U6409, P2_U6410);
  nand ginst12470 (P2_U2901, P2_U6401, P2_U6402, P2_U6403, P2_U6404, P2_U6405);
  nand ginst12471 (P2_U2902, P2_U6396, P2_U6397, P2_U6398, P2_U6399, P2_U6400);
  nand ginst12472 (P2_U2903, P2_U6391, P2_U6392, P2_U6393, P2_U6394, P2_U6395);
  nand ginst12473 (P2_U2904, P2_U6387, P2_U6388, P2_U6389, P2_U6390);
  nand ginst12474 (P2_U2905, P2_U6383, P2_U6384, P2_U6385, P2_U6386);
  nand ginst12475 (P2_U2906, P2_U6379, P2_U6380, P2_U6381, P2_U6382);
  nand ginst12476 (P2_U2907, P2_U6375, P2_U6376, P2_U6377, P2_U6378);
  nand ginst12477 (P2_U2908, P2_U6371, P2_U6372, P2_U6373, P2_U6374);
  nand ginst12478 (P2_U2909, P2_U6367, P2_U6368, P2_U6369, P2_U6370);
  nand ginst12479 (P2_U2910, P2_U4068, P2_U6363, P2_U6364);
  nand ginst12480 (P2_U2911, P2_U4067, P2_U6359, P2_U6360);
  nand ginst12481 (P2_U2912, P2_U4066, P2_U6355, P2_U6356);
  nand ginst12482 (P2_U2913, P2_U4065, P2_U6351, P2_U6352);
  nand ginst12483 (P2_U2914, P2_U4064, P2_U6347, P2_U6348);
  nand ginst12484 (P2_U2915, P2_U4063, P2_U6343, P2_U6344);
  nand ginst12485 (P2_U2916, P2_U4062, P2_U6339, P2_U6340);
  nand ginst12486 (P2_U2917, P2_U4061, P2_U6335, P2_U6336);
  nand ginst12487 (P2_U2918, P2_U4060, P2_U6331, P2_U6332);
  nand ginst12488 (P2_U2919, P2_U4059, P2_U6327, P2_U6328);
  and ginst12489 (P2_U2920, P2_DATAO_REG_31__SCAN_IN, P2_U6232);
  nand ginst12490 (P2_U2921, P2_U6323, P2_U6324, P2_U6325);
  nand ginst12491 (P2_U2922, P2_U6320, P2_U6321, P2_U6322);
  nand ginst12492 (P2_U2923, P2_U6317, P2_U6318, P2_U6319);
  nand ginst12493 (P2_U2924, P2_U6314, P2_U6315, P2_U6316);
  nand ginst12494 (P2_U2925, P2_U6311, P2_U6312, P2_U6313);
  nand ginst12495 (P2_U2926, P2_U6308, P2_U6309, P2_U6310);
  nand ginst12496 (P2_U2927, P2_U6305, P2_U6306, P2_U6307);
  nand ginst12497 (P2_U2928, P2_U6302, P2_U6303, P2_U6304);
  nand ginst12498 (P2_U2929, P2_U6299, P2_U6300, P2_U6301);
  nand ginst12499 (P2_U2930, P2_U6296, P2_U6297, P2_U6298);
  nand ginst12500 (P2_U2931, P2_U6293, P2_U6294, P2_U6295);
  nand ginst12501 (P2_U2932, P2_U6290, P2_U6291, P2_U6292);
  nand ginst12502 (P2_U2933, P2_U6287, P2_U6288, P2_U6289);
  nand ginst12503 (P2_U2934, P2_U6284, P2_U6285, P2_U6286);
  nand ginst12504 (P2_U2935, P2_U6281, P2_U6282, P2_U6283);
  nand ginst12505 (P2_U2936, P2_U6278, P2_U6279, P2_U6280);
  nand ginst12506 (P2_U2937, P2_U6275, P2_U6276, P2_U6277);
  nand ginst12507 (P2_U2938, P2_U6272, P2_U6273, P2_U6274);
  nand ginst12508 (P2_U2939, P2_U6269, P2_U6270, P2_U6271);
  nand ginst12509 (P2_U2940, P2_U6266, P2_U6267, P2_U6268);
  nand ginst12510 (P2_U2941, P2_U6263, P2_U6264, P2_U6265);
  nand ginst12511 (P2_U2942, P2_U6260, P2_U6261, P2_U6262);
  nand ginst12512 (P2_U2943, P2_U6257, P2_U6258, P2_U6259);
  nand ginst12513 (P2_U2944, P2_U6254, P2_U6255, P2_U6256);
  nand ginst12514 (P2_U2945, P2_U6251, P2_U6252, P2_U6253);
  nand ginst12515 (P2_U2946, P2_U6248, P2_U6249, P2_U6250);
  nand ginst12516 (P2_U2947, P2_U6245, P2_U6246, P2_U6247);
  nand ginst12517 (P2_U2948, P2_U6242, P2_U6243, P2_U6244);
  nand ginst12518 (P2_U2949, P2_U6239, P2_U6240, P2_U6241);
  nand ginst12519 (P2_U2950, P2_U6236, P2_U6237, P2_U6238);
  nand ginst12520 (P2_U2951, P2_U6233, P2_U6234, P2_U6235);
  nand ginst12521 (P2_U2952, P2_U6224, P2_U6225, P2_U6226);
  nand ginst12522 (P2_U2953, P2_U6221, P2_U6222, P2_U6223);
  nand ginst12523 (P2_U2954, P2_U6218, P2_U6219, P2_U6220);
  nand ginst12524 (P2_U2955, P2_U6215, P2_U6216, P2_U6217);
  nand ginst12525 (P2_U2956, P2_U6212, P2_U6213, P2_U6214);
  nand ginst12526 (P2_U2957, P2_U6209, P2_U6210, P2_U6211);
  nand ginst12527 (P2_U2958, P2_U6206, P2_U6207, P2_U6208);
  nand ginst12528 (P2_U2959, P2_U6203, P2_U6204, P2_U6205);
  nand ginst12529 (P2_U2960, P2_U6200, P2_U6201, P2_U6202);
  nand ginst12530 (P2_U2961, P2_U6197, P2_U6198, P2_U6199);
  nand ginst12531 (P2_U2962, P2_U6194, P2_U6195, P2_U6196);
  nand ginst12532 (P2_U2963, P2_U6191, P2_U6192, P2_U6193);
  nand ginst12533 (P2_U2964, P2_U6188, P2_U6189, P2_U6190);
  nand ginst12534 (P2_U2965, P2_U6185, P2_U6186, P2_U6187);
  nand ginst12535 (P2_U2966, P2_U6182, P2_U6183, P2_U6184);
  nand ginst12536 (P2_U2967, P2_U6179, P2_U6180, P2_U6181);
  nand ginst12537 (P2_U2968, P2_U6176, P2_U6177, P2_U6178);
  nand ginst12538 (P2_U2969, P2_U6173, P2_U6174, P2_U6175);
  nand ginst12539 (P2_U2970, P2_U6170, P2_U6171, P2_U6172);
  nand ginst12540 (P2_U2971, P2_U6167, P2_U6168, P2_U6169);
  nand ginst12541 (P2_U2972, P2_U6164, P2_U6165, P2_U6166);
  nand ginst12542 (P2_U2973, P2_U6161, P2_U6162, P2_U6163);
  nand ginst12543 (P2_U2974, P2_U6158, P2_U6159, P2_U6160);
  nand ginst12544 (P2_U2975, P2_U6155, P2_U6156, P2_U6157);
  nand ginst12545 (P2_U2976, P2_U6152, P2_U6153, P2_U6154);
  nand ginst12546 (P2_U2977, P2_U6149, P2_U6150, P2_U6151);
  nand ginst12547 (P2_U2978, P2_U6146, P2_U6147, P2_U6148);
  nand ginst12548 (P2_U2979, P2_U6143, P2_U6144, P2_U6145);
  nand ginst12549 (P2_U2980, P2_U6140, P2_U6141, P2_U6142);
  nand ginst12550 (P2_U2981, P2_U6137, P2_U6138, P2_U6139);
  nand ginst12551 (P2_U2982, P2_U6134, P2_U6135, P2_U6136);
  nand ginst12552 (P2_U2983, P2_U4053, P2_U4054);
  nand ginst12553 (P2_U2984, P2_U4051, P2_U4052);
  nand ginst12554 (P2_U2985, P2_U4049, P2_U4050);
  nand ginst12555 (P2_U2986, P2_U4047, P2_U4048);
  nand ginst12556 (P2_U2987, P2_U4045, P2_U4046);
  nand ginst12557 (P2_U2988, P2_U4043, P2_U4044);
  nand ginst12558 (P2_U2989, P2_U4041, P2_U4042);
  nand ginst12559 (P2_U2990, P2_U4039, P2_U4040);
  nand ginst12560 (P2_U2991, P2_U4037, P2_U4038);
  nand ginst12561 (P2_U2992, P2_U4035, P2_U4036);
  nand ginst12562 (P2_U2993, P2_U4033, P2_U4034);
  nand ginst12563 (P2_U2994, P2_U4031, P2_U4032);
  nand ginst12564 (P2_U2995, P2_U4029, P2_U4030);
  nand ginst12565 (P2_U2996, P2_U4027, P2_U4028);
  nand ginst12566 (P2_U2997, P2_U4025, P2_U4026);
  nand ginst12567 (P2_U2998, P2_U4023, P2_U4024);
  nand ginst12568 (P2_U2999, P2_U4021, P2_U4022);
  nand ginst12569 (P2_U3000, P2_U4019, P2_U4020);
  nand ginst12570 (P2_U3001, P2_U4017, P2_U4018);
  nand ginst12571 (P2_U3002, P2_U4015, P2_U4016);
  nand ginst12572 (P2_U3003, P2_U4013, P2_U4014);
  nand ginst12573 (P2_U3004, P2_U4011, P2_U4012);
  nand ginst12574 (P2_U3005, P2_U4009, P2_U4010);
  nand ginst12575 (P2_U3006, P2_U4007, P2_U4008);
  nand ginst12576 (P2_U3007, P2_U4005, P2_U4006);
  nand ginst12577 (P2_U3008, P2_U4003, P2_U4004);
  nand ginst12578 (P2_U3009, P2_U4001, P2_U4002);
  nand ginst12579 (P2_U3010, P2_U3999, P2_U4000);
  nand ginst12580 (P2_U3011, P2_U3997, P2_U3998);
  nand ginst12581 (P2_U3012, P2_U3995, P2_U3996);
  nand ginst12582 (P2_U3013, P2_U3993, P2_U3994);
  nand ginst12583 (P2_U3014, P2_U3991, P2_U3992);
  nand ginst12584 (P2_U3015, P2_U3987, P2_U3988, P2_U5928, P2_U5932, P2_U5933);
  nand ginst12585 (P2_U3016, P2_U3985, P2_U3986, P2_U5920, P2_U5924, P2_U5925);
  nand ginst12586 (P2_U3017, P2_U3983, P2_U3984, P2_U5916, P2_U5917);
  nand ginst12587 (P2_U3018, P2_U3980, P2_U3981, P2_U3982, P2_U5908, P2_U5909);
  nand ginst12588 (P2_U3019, P2_U3977, P2_U3978, P2_U3979, P2_U5900, P2_U5901);
  nand ginst12589 (P2_U3020, P2_U3974, P2_U3975, P2_U3976, P2_U5892, P2_U5893);
  nand ginst12590 (P2_U3021, P2_U3971, P2_U3972, P2_U3973, P2_U5884, P2_U5885);
  nand ginst12591 (P2_U3022, P2_U3968, P2_U3969, P2_U3970, P2_U5876, P2_U5877);
  nand ginst12592 (P2_U3023, P2_U3965, P2_U3966, P2_U3967, P2_U5868, P2_U5869);
  nand ginst12593 (P2_U3024, P2_U3962, P2_U3963, P2_U3964, P2_U5860, P2_U5861);
  nand ginst12594 (P2_U3025, P2_U3959, P2_U3960, P2_U3961, P2_U5852, P2_U5853);
  nand ginst12595 (P2_U3026, P2_U3956, P2_U3957, P2_U3958, P2_U5844, P2_U5845);
  nand ginst12596 (P2_U3027, P2_U3953, P2_U3954, P2_U3955, P2_U5836, P2_U5837);
  nand ginst12597 (P2_U3028, P2_U3950, P2_U3951, P2_U3952, P2_U5828, P2_U5829);
  nand ginst12598 (P2_U3029, P2_U3947, P2_U3948, P2_U3949, P2_U5820, P2_U5821);
  nand ginst12599 (P2_U3030, P2_U3944, P2_U3945, P2_U3946, P2_U5812, P2_U5813);
  nand ginst12600 (P2_U3031, P2_U3941, P2_U3942, P2_U3943, P2_U5804, P2_U5805);
  nand ginst12601 (P2_U3032, P2_U3938, P2_U3939, P2_U3940, P2_U5796, P2_U5797);
  nand ginst12602 (P2_U3033, P2_U3935, P2_U3936, P2_U3937, P2_U5788, P2_U5789);
  nand ginst12603 (P2_U3034, P2_U3932, P2_U3933, P2_U3934, P2_U5780, P2_U5781);
  nand ginst12604 (P2_U3035, P2_U3929, P2_U3930, P2_U3931, P2_U5772, P2_U5773);
  nand ginst12605 (P2_U3036, P2_U3926, P2_U3927, P2_U3928, P2_U5764, P2_U5765);
  nand ginst12606 (P2_U3037, P2_U3923, P2_U3924, P2_U3925, P2_U5756, P2_U5757);
  nand ginst12607 (P2_U3038, P2_U3920, P2_U3921, P2_U3922, P2_U5748, P2_U5749);
  nand ginst12608 (P2_U3039, P2_U3917, P2_U3918, P2_U3919, P2_U5740, P2_U5741);
  nand ginst12609 (P2_U3040, P2_U3914, P2_U3915, P2_U3916, P2_U5732, P2_U5733);
  nand ginst12610 (P2_U3041, P2_U3911, P2_U3912, P2_U3913, P2_U5724, P2_U5725);
  nand ginst12611 (P2_U3042, P2_U3908, P2_U3909, P2_U3910, P2_U5716, P2_U5717);
  nand ginst12612 (P2_U3043, P2_U3905, P2_U3906, P2_U3907, P2_U5708, P2_U5709);
  nand ginst12613 (P2_U3044, P2_U3902, P2_U3903, P2_U3904, P2_U5700, P2_U5701);
  nand ginst12614 (P2_U3045, P2_U3899, P2_U3900, P2_U3901, P2_U5692, P2_U5693);
  nand ginst12615 (P2_U3046, P2_U3896, P2_U3897, P2_U3898, P2_U5684, P2_U5685);
  and ginst12616 (P2_U3047, P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN, P2_U5643);
  nand ginst12617 (P2_U3048, P2_U3865, P2_U5569, P2_U5570);
  nand ginst12618 (P2_U3049, P2_U3864, P2_U5564, P2_U5565);
  nand ginst12619 (P2_U3050, P2_U3863, P2_U5559, P2_U5560);
  nand ginst12620 (P2_U3051, P2_U3862, P2_U5554, P2_U5555);
  nand ginst12621 (P2_U3052, P2_U3861, P2_U5549, P2_U5550);
  nand ginst12622 (P2_U3053, P2_U3860, P2_U5544, P2_U5545);
  nand ginst12623 (P2_U3054, P2_U3859, P2_U5539, P2_U5540);
  nand ginst12624 (P2_U3055, P2_U3858, P2_U5534, P2_U5535);
  nand ginst12625 (P2_U3056, P2_U3856, P2_U5512, P2_U5513);
  nand ginst12626 (P2_U3057, P2_U3855, P2_U5507, P2_U5508);
  nand ginst12627 (P2_U3058, P2_U3854, P2_U5502, P2_U5503);
  nand ginst12628 (P2_U3059, P2_U3853, P2_U5497, P2_U5498);
  nand ginst12629 (P2_U3060, P2_U3852, P2_U5492, P2_U5493);
  nand ginst12630 (P2_U3061, P2_U3851, P2_U5487, P2_U5488);
  nand ginst12631 (P2_U3062, P2_U3850, P2_U5482, P2_U5483);
  nand ginst12632 (P2_U3063, P2_U3849, P2_U5477, P2_U5478);
  nand ginst12633 (P2_U3064, P2_U3847, P2_U5454, P2_U5455);
  nand ginst12634 (P2_U3065, P2_U3846, P2_U5449, P2_U5450);
  nand ginst12635 (P2_U3066, P2_U3845, P2_U5444, P2_U5445);
  nand ginst12636 (P2_U3067, P2_U3844, P2_U5439, P2_U5440);
  nand ginst12637 (P2_U3068, P2_U3843, P2_U5434, P2_U5435);
  nand ginst12638 (P2_U3069, P2_U3842, P2_U5429, P2_U5430);
  nand ginst12639 (P2_U3070, P2_U3841, P2_U5424, P2_U5425);
  nand ginst12640 (P2_U3071, P2_U3840, P2_U5419, P2_U5420);
  nand ginst12641 (P2_U3072, P2_U3838, P2_U5397, P2_U5398);
  nand ginst12642 (P2_U3073, P2_U3837, P2_U5392, P2_U5393);
  nand ginst12643 (P2_U3074, P2_U3836, P2_U5387, P2_U5388);
  nand ginst12644 (P2_U3075, P2_U3835, P2_U5382, P2_U5383);
  nand ginst12645 (P2_U3076, P2_U3834, P2_U5377, P2_U5378);
  nand ginst12646 (P2_U3077, P2_U3833, P2_U5372, P2_U5373);
  nand ginst12647 (P2_U3078, P2_U3832, P2_U5367, P2_U5368);
  nand ginst12648 (P2_U3079, P2_U3831, P2_U5362, P2_U5363);
  nand ginst12649 (P2_U3080, P2_U3829, P2_U5339, P2_U5340);
  nand ginst12650 (P2_U3081, P2_U3828, P2_U5334, P2_U5335);
  nand ginst12651 (P2_U3082, P2_U3827, P2_U5329, P2_U5330);
  nand ginst12652 (P2_U3083, P2_U3826, P2_U5324, P2_U5325);
  nand ginst12653 (P2_U3084, P2_U3825, P2_U5319, P2_U5320);
  nand ginst12654 (P2_U3085, P2_U3824, P2_U5314, P2_U5315);
  nand ginst12655 (P2_U3086, P2_U3823, P2_U5309, P2_U5310);
  nand ginst12656 (P2_U3087, P2_U3822, P2_U5304, P2_U5305);
  nand ginst12657 (P2_U3088, P2_U3820, P2_U5282, P2_U5283);
  nand ginst12658 (P2_U3089, P2_U3819, P2_U5277, P2_U5278);
  nand ginst12659 (P2_U3090, P2_U3818, P2_U5272, P2_U5273);
  nand ginst12660 (P2_U3091, P2_U3817, P2_U5267, P2_U5268);
  nand ginst12661 (P2_U3092, P2_U3816, P2_U5262, P2_U5263);
  nand ginst12662 (P2_U3093, P2_U3815, P2_U5257, P2_U5258);
  nand ginst12663 (P2_U3094, P2_U3814, P2_U5252, P2_U5253);
  nand ginst12664 (P2_U3095, P2_U3813, P2_U5247, P2_U5248);
  nand ginst12665 (P2_U3096, P2_U3811, P2_U5224, P2_U5225);
  nand ginst12666 (P2_U3097, P2_U3810, P2_U5219, P2_U5220);
  nand ginst12667 (P2_U3098, P2_U3809, P2_U5214, P2_U5215);
  nand ginst12668 (P2_U3099, P2_U3808, P2_U5209, P2_U5210);
  nand ginst12669 (P2_U3100, P2_U3807, P2_U5204, P2_U5205);
  nand ginst12670 (P2_U3101, P2_U3806, P2_U5199, P2_U5200);
  nand ginst12671 (P2_U3102, P2_U3805, P2_U5194, P2_U5195);
  nand ginst12672 (P2_U3103, P2_U3804, P2_U5189, P2_U5190);
  nand ginst12673 (P2_U3104, P2_U3802, P2_U5167, P2_U5168);
  nand ginst12674 (P2_U3105, P2_U3801, P2_U5162, P2_U5163);
  nand ginst12675 (P2_U3106, P2_U3800, P2_U5157, P2_U5158);
  nand ginst12676 (P2_U3107, P2_U3799, P2_U5152, P2_U5153);
  nand ginst12677 (P2_U3108, P2_U3798, P2_U5147, P2_U5148);
  nand ginst12678 (P2_U3109, P2_U3797, P2_U5142, P2_U5143);
  nand ginst12679 (P2_U3110, P2_U3796, P2_U5137, P2_U5138);
  nand ginst12680 (P2_U3111, P2_U3795, P2_U5132, P2_U5133);
  nand ginst12681 (P2_U3112, P2_U3793, P2_U5111, P2_U5112);
  nand ginst12682 (P2_U3113, P2_U3792, P2_U5106, P2_U5107);
  nand ginst12683 (P2_U3114, P2_U3791, P2_U5101, P2_U5102);
  nand ginst12684 (P2_U3115, P2_U3790, P2_U5096, P2_U5097);
  nand ginst12685 (P2_U3116, P2_U3789, P2_U5091, P2_U5092);
  nand ginst12686 (P2_U3117, P2_U3788, P2_U5086, P2_U5087);
  nand ginst12687 (P2_U3118, P2_U3787, P2_U5081, P2_U5082);
  nand ginst12688 (P2_U3119, P2_U3786, P2_U5076, P2_U5077);
  nand ginst12689 (P2_U3120, P2_U3784, P2_U5054, P2_U5055);
  nand ginst12690 (P2_U3121, P2_U3783, P2_U5049, P2_U5050);
  nand ginst12691 (P2_U3122, P2_U3782, P2_U5044, P2_U5045);
  nand ginst12692 (P2_U3123, P2_U3781, P2_U5039, P2_U5040);
  nand ginst12693 (P2_U3124, P2_U3780, P2_U5034, P2_U5035);
  nand ginst12694 (P2_U3125, P2_U3779, P2_U5029, P2_U5030);
  nand ginst12695 (P2_U3126, P2_U3778, P2_U5024, P2_U5025);
  nand ginst12696 (P2_U3127, P2_U3777, P2_U5019, P2_U5020);
  nand ginst12697 (P2_U3128, P2_U3775, P2_U4996, P2_U4997);
  nand ginst12698 (P2_U3129, P2_U3774, P2_U4991, P2_U4992);
  nand ginst12699 (P2_U3130, P2_U3773, P2_U4986, P2_U4987);
  nand ginst12700 (P2_U3131, P2_U3772, P2_U4981, P2_U4982);
  nand ginst12701 (P2_U3132, P2_U3771, P2_U4976, P2_U4977);
  nand ginst12702 (P2_U3133, P2_U3770, P2_U4971, P2_U4972);
  nand ginst12703 (P2_U3134, P2_U3769, P2_U4966, P2_U4967);
  nand ginst12704 (P2_U3135, P2_U3768, P2_U4961, P2_U4962);
  nand ginst12705 (P2_U3136, P2_U3766, P2_U4939, P2_U4940);
  nand ginst12706 (P2_U3137, P2_U3765, P2_U4934, P2_U4935);
  nand ginst12707 (P2_U3138, P2_U3764, P2_U4929, P2_U4930);
  nand ginst12708 (P2_U3139, P2_U3763, P2_U4924, P2_U4925);
  nand ginst12709 (P2_U3140, P2_U3762, P2_U4919, P2_U4920);
  nand ginst12710 (P2_U3141, P2_U3761, P2_U4914, P2_U4915);
  nand ginst12711 (P2_U3142, P2_U3760, P2_U4909, P2_U4910);
  nand ginst12712 (P2_U3143, P2_U3759, P2_U4904, P2_U4905);
  nand ginst12713 (P2_U3144, P2_U3757, P2_U4881, P2_U4882);
  nand ginst12714 (P2_U3145, P2_U3756, P2_U4876, P2_U4877);
  nand ginst12715 (P2_U3146, P2_U3755, P2_U4871, P2_U4872);
  nand ginst12716 (P2_U3147, P2_U3754, P2_U4866, P2_U4867);
  nand ginst12717 (P2_U3148, P2_U3753, P2_U4861, P2_U4862);
  nand ginst12718 (P2_U3149, P2_U3752, P2_U4856, P2_U4857);
  nand ginst12719 (P2_U3150, P2_U3751, P2_U4851, P2_U4852);
  nand ginst12720 (P2_U3151, P2_U3750, P2_U4846, P2_U4847);
  nand ginst12721 (P2_U3152, P2_U3748, P2_U4824, P2_U4825);
  nand ginst12722 (P2_U3153, P2_U3747, P2_U4819, P2_U4820);
  nand ginst12723 (P2_U3154, P2_U3746, P2_U4814, P2_U4815);
  nand ginst12724 (P2_U3155, P2_U3745, P2_U4809, P2_U4810);
  nand ginst12725 (P2_U3156, P2_U3744, P2_U4804, P2_U4805);
  nand ginst12726 (P2_U3157, P2_U3743, P2_U4799, P2_U4800);
  nand ginst12727 (P2_U3158, P2_U3742, P2_U4794, P2_U4795);
  nand ginst12728 (P2_U3159, P2_U3741, P2_U4789, P2_U4790);
  nand ginst12729 (P2_U3160, P2_U3739, P2_U4765, P2_U4766);
  nand ginst12730 (P2_U3161, P2_U3738, P2_U4760, P2_U4761);
  nand ginst12731 (P2_U3162, P2_U3737, P2_U4755, P2_U4756);
  nand ginst12732 (P2_U3163, P2_U3736, P2_U4750, P2_U4751);
  nand ginst12733 (P2_U3164, P2_U3735, P2_U4745, P2_U4746);
  nand ginst12734 (P2_U3165, P2_U3734, P2_U4740, P2_U4741);
  nand ginst12735 (P2_U3166, P2_U3733, P2_U4735, P2_U4736);
  nand ginst12736 (P2_U3167, P2_U3732, P2_U4730, P2_U4731);
  nand ginst12737 (P2_U3168, P2_U3730, P2_U4707, P2_U4708);
  nand ginst12738 (P2_U3169, P2_U3729, P2_U4702, P2_U4703);
  nand ginst12739 (P2_U3170, P2_U3728, P2_U4697, P2_U4698);
  nand ginst12740 (P2_U3171, P2_U3727, P2_U4692, P2_U4693);
  nand ginst12741 (P2_U3172, P2_U3726, P2_U4687, P2_U4688);
  nand ginst12742 (P2_U3173, P2_U3725, P2_U4682, P2_U4683);
  nand ginst12743 (P2_U3174, P2_U3724, P2_U4677, P2_U4678);
  nand ginst12744 (P2_U3175, P2_U3723, P2_U4672, P2_U4673);
  nand ginst12745 (P2_U3176, P2_U3721, P2_U8060, P2_U8061);
  nand ginst12746 (P2_U3177, P2_U4454, P2_U4627, P2_U4628, P2_U4629);
  nand ginst12747 (P2_U3178, P2_U3716, P2_U4625);
  and ginst12748 (P2_U3179, P2_DATAWIDTH_REG_31__SCAN_IN, P2_U7917);
  and ginst12749 (P2_U3180, P2_DATAWIDTH_REG_30__SCAN_IN, P2_U7917);
  and ginst12750 (P2_U3181, P2_DATAWIDTH_REG_29__SCAN_IN, P2_U7917);
  and ginst12751 (P2_U3182, P2_DATAWIDTH_REG_28__SCAN_IN, P2_U7917);
  and ginst12752 (P2_U3183, P2_DATAWIDTH_REG_27__SCAN_IN, P2_U7917);
  and ginst12753 (P2_U3184, P2_DATAWIDTH_REG_26__SCAN_IN, P2_U7917);
  and ginst12754 (P2_U3185, P2_DATAWIDTH_REG_25__SCAN_IN, P2_U7917);
  and ginst12755 (P2_U3186, P2_DATAWIDTH_REG_24__SCAN_IN, P2_U7917);
  and ginst12756 (P2_U3187, P2_DATAWIDTH_REG_23__SCAN_IN, P2_U7917);
  and ginst12757 (P2_U3188, P2_DATAWIDTH_REG_22__SCAN_IN, P2_U7917);
  and ginst12758 (P2_U3189, P2_DATAWIDTH_REG_21__SCAN_IN, P2_U7917);
  and ginst12759 (P2_U3190, P2_DATAWIDTH_REG_20__SCAN_IN, P2_U7917);
  and ginst12760 (P2_U3191, P2_DATAWIDTH_REG_19__SCAN_IN, P2_U7917);
  and ginst12761 (P2_U3192, P2_DATAWIDTH_REG_18__SCAN_IN, P2_U7917);
  and ginst12762 (P2_U3193, P2_DATAWIDTH_REG_17__SCAN_IN, P2_U7917);
  and ginst12763 (P2_U3194, P2_DATAWIDTH_REG_16__SCAN_IN, P2_U7917);
  and ginst12764 (P2_U3195, P2_DATAWIDTH_REG_15__SCAN_IN, P2_U7917);
  and ginst12765 (P2_U3196, P2_DATAWIDTH_REG_14__SCAN_IN, P2_U7917);
  and ginst12766 (P2_U3197, P2_DATAWIDTH_REG_13__SCAN_IN, P2_U7917);
  and ginst12767 (P2_U3198, P2_DATAWIDTH_REG_12__SCAN_IN, P2_U7917);
  and ginst12768 (P2_U3199, P2_DATAWIDTH_REG_11__SCAN_IN, P2_U7917);
  and ginst12769 (P2_U3200, P2_DATAWIDTH_REG_10__SCAN_IN, P2_U7917);
  and ginst12770 (P2_U3201, P2_DATAWIDTH_REG_9__SCAN_IN, P2_U7917);
  and ginst12771 (P2_U3202, P2_DATAWIDTH_REG_8__SCAN_IN, P2_U7917);
  and ginst12772 (P2_U3203, P2_DATAWIDTH_REG_7__SCAN_IN, P2_U7917);
  and ginst12773 (P2_U3204, P2_DATAWIDTH_REG_6__SCAN_IN, P2_U7917);
  and ginst12774 (P2_U3205, P2_DATAWIDTH_REG_5__SCAN_IN, P2_U7917);
  and ginst12775 (P2_U3206, P2_DATAWIDTH_REG_4__SCAN_IN, P2_U7917);
  and ginst12776 (P2_U3207, P2_DATAWIDTH_REG_3__SCAN_IN, P2_U7917);
  and ginst12777 (P2_U3208, P2_DATAWIDTH_REG_2__SCAN_IN, P2_U7917);
  nand ginst12778 (P2_U3209, P2_U4588, P2_U7913, P2_U7914);
  nand ginst12779 (P2_U3210, P2_U3691, P2_U7911, P2_U7912);
  nand ginst12780 (P2_U3211, P2_U3690, P2_U4579);
  nand ginst12781 (P2_U3212, P2_U4565, P2_U4566, P2_U4567);
  nand ginst12782 (P2_U3213, P2_U4562, P2_U4563, P2_U4564);
  nand ginst12783 (P2_U3214, P2_U4559, P2_U4560, P2_U4561);
  nand ginst12784 (P2_U3215, P2_U4556, P2_U4557, P2_U4558);
  nand ginst12785 (P2_U3216, P2_U4553, P2_U4554, P2_U4555);
  nand ginst12786 (P2_U3217, P2_U4550, P2_U4551, P2_U4552);
  nand ginst12787 (P2_U3218, P2_U4547, P2_U4548, P2_U4549);
  nand ginst12788 (P2_U3219, P2_U4544, P2_U4545, P2_U4546);
  nand ginst12789 (P2_U3220, P2_U4541, P2_U4542, P2_U4543);
  nand ginst12790 (P2_U3221, P2_U4538, P2_U4539, P2_U4540);
  nand ginst12791 (P2_U3222, P2_U4535, P2_U4536, P2_U4537);
  nand ginst12792 (P2_U3223, P2_U4532, P2_U4533, P2_U4534);
  nand ginst12793 (P2_U3224, P2_U4529, P2_U4530, P2_U4531);
  nand ginst12794 (P2_U3225, P2_U4526, P2_U4527, P2_U4528);
  nand ginst12795 (P2_U3226, P2_U4523, P2_U4524, P2_U4525);
  nand ginst12796 (P2_U3227, P2_U4520, P2_U4521, P2_U4522);
  nand ginst12797 (P2_U3228, P2_U4517, P2_U4518, P2_U4519);
  nand ginst12798 (P2_U3229, P2_U4514, P2_U4515, P2_U4516);
  nand ginst12799 (P2_U3230, P2_U4511, P2_U4512, P2_U4513);
  nand ginst12800 (P2_U3231, P2_U4508, P2_U4509, P2_U4510);
  nand ginst12801 (P2_U3232, P2_U4505, P2_U4506, P2_U4507);
  nand ginst12802 (P2_U3233, P2_U4502, P2_U4503, P2_U4504);
  nand ginst12803 (P2_U3234, P2_U4499, P2_U4500, P2_U4501);
  nand ginst12804 (P2_U3235, P2_U4496, P2_U4497, P2_U4498);
  nand ginst12805 (P2_U3236, P2_U4493, P2_U4494, P2_U4495);
  nand ginst12806 (P2_U3237, P2_U4490, P2_U4491, P2_U4492);
  nand ginst12807 (P2_U3238, P2_U4487, P2_U4488, P2_U4489);
  nand ginst12808 (P2_U3239, P2_U4484, P2_U4485, P2_U4486);
  nand ginst12809 (P2_U3240, P2_U4481, P2_U4482, P2_U4483);
  nand ginst12810 (P2_U3241, P2_U4478, P2_U4479, P2_U4480);
  nand ginst12811 (P2_U3242, P2_U4191, P2_U4192, P2_U4193, P2_U4194);
  nand ginst12812 (P2_U3243, P2_U3335, P2_U3349);
  not ginst12813 (P2_U3244, P2_STATE_REG_2__SCAN_IN);
  nand ginst12814 (P2_U3245, P2_U2440, P2_U3243);
  nand ginst12815 (P2_U3246, P2_U2440, P2_U4650);
  nand ginst12816 (P2_U3247, P2_U2442, P2_U3243);
  nand ginst12817 (P2_U3248, P2_U2442, P2_U4650);
  nand ginst12818 (P2_U3249, P2_U2441, P2_U3243);
  nand ginst12819 (P2_U3250, P2_U2441, P2_U4650);
  nand ginst12820 (P2_U3251, P2_U2443, P2_U3243);
  nand ginst12821 (P2_U3252, P2_U2443, P2_U4650);
  nand ginst12822 (P2_U3253, P2_U3707, P2_U3708);
  nand ginst12823 (P2_U3254, P2_U2590, P2_U4429);
  nand ginst12824 (P2_U3255, P2_U3695, P2_U3696);
  not ginst12825 (P2_U3256, P2_REQUESTPENDING_REG_SCAN_IN);
  nand ginst12826 (P2_U3257, P2_U4608, P2_U4609, P2_U8050, P2_U8051);
  not ginst12827 (P2_U3258, P2_STATE_REG_1__SCAN_IN);
  nand ginst12828 (P2_U3259, P2_STATE_REG_1__SCAN_IN, P2_U3266);
  nand ginst12829 (P2_U3260, P2_U3244, P2_U4439);
  nand ginst12830 (P2_U3261, P2_STATE_REG_2__SCAN_IN, P2_U4439);
  nand ginst12831 (P2_U3262, P2_STATE_REG_1__SCAN_IN, P2_U3244);
  or ginst12832 (P2_U3263, P2_STATE_REG_2__SCAN_IN, P2_STATE_REG_1__SCAN_IN);
  not ginst12833 (P2_U3264, HOLD);
  not ginst12834 (P2_U3265, U211);
  not ginst12835 (P2_U3266, P2_STATE_REG_0__SCAN_IN);
  nand ginst12836 (P2_U3267, P2_REQUESTPENDING_REG_SCAN_IN, P2_U3264);
  or ginst12837 (P2_U3268, HOLD, P2_REQUESTPENDING_REG_SCAN_IN);
  not ginst12838 (P2_U3269, P2_STATE2_REG_1__SCAN_IN);
  not ginst12839 (P2_U3270, P2_STATE2_REG_2__SCAN_IN);
  not ginst12840 (P2_U3271, P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN);
  not ginst12841 (P2_U3272, P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN);
  not ginst12842 (P2_U3273, P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN);
  nand ginst12843 (P2_U3274, P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN, P2_U3276);
  or ginst12844 (P2_U3275, P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN);
  not ginst12845 (P2_U3276, P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN);
  nand ginst12846 (P2_U3277, P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN);
  nand ginst12847 (P2_U3278, P2_U3699, P2_U3700);
  nand ginst12848 (P2_U3279, P2_U3701, P2_U3702);
  nand ginst12849 (P2_U3280, P2_U3703, P2_U3704);
  nand ginst12850 (P2_U3281, P2_U7859, P2_U7861, P2_U7863);
  nand ginst12851 (P2_U3282, P2_U2457, P2_U4476, P2_U7869);
  nand ginst12852 (P2_U3283, P2_U3253, P2_U7873);
  not ginst12853 (P2_U3284, P2_STATE2_REG_0__SCAN_IN);
  nand ginst12854 (P2_U3285, P2_U3709, P2_U4424);
  nand ginst12855 (P2_U3286, P2_U2616, P2_U3253);
  not ginst12856 (P2_U3287, P2_GTE_370_U6);
  nand ginst12857 (P2_U3288, P2_U2457, P2_U2458, P2_U7859);
  nand ginst12858 (P2_U3289, P2_U2616, P2_U7871);
  nand ginst12859 (P2_U3290, P2_U3266, P2_U4595);
  nand ginst12860 (P2_U3291, P2_U2459, P2_U3713);
  not ginst12861 (P2_U3292, P2_R2243_U8);
  nand ginst12862 (P2_U3293, P2_U2357, P2_U3280);
  nand ginst12863 (P2_U3294, P2_U7871, P2_U7873);
  nand ginst12864 (P2_U3295, P2_U2617, P2_U7861);
  nand ginst12865 (P2_U3296, P2_U2451, P2_U4428);
  not ginst12866 (P2_U3297, P2_R2167_U6);
  nand ginst12867 (P2_U3298, P2_LT_563_U6, P2_U4444, P2_U4610, P2_U4614, P2_U7894);
  nand ginst12868 (P2_U3299, P2_STATE2_REG_0__SCAN_IN, P2_U4619);
  not ginst12869 (P2_U3300, P2_STATE2_REG_3__SCAN_IN);
  nand ginst12870 (P2_U3301, P2_STATE2_REG_0__SCAN_IN, P2_U3270);
  not ginst12871 (P2_U3302, P2_STATEBS16_REG_SCAN_IN);
  or ginst12872 (P2_U3303, P2_STATE2_REG_3__SCAN_IN, P2_STATE2_REG_1__SCAN_IN);
  nand ginst12873 (P2_U3304, P2_STATE2_REG_2__SCAN_IN, P2_U3269);
  nand ginst12874 (P2_U3305, P2_STATE2_REG_3__SCAN_IN, P2_R2167_U6);
  nand ginst12875 (P2_U3306, P2_U3284, P2_U4656);
  not ginst12876 (P2_U3307, P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN);
  not ginst12877 (P2_U3308, P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN);
  not ginst12878 (P2_U3309, P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN);
  not ginst12879 (P2_U3310, P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN);
  nand ginst12880 (P2_U3311, P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN, P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN);
  nand ginst12881 (P2_U3312, P2_U2464, P2_U4642);
  or ginst12882 (P2_U3313, P2_STATE2_REG_3__SCAN_IN, P2_STATE2_REG_2__SCAN_IN);
  not ginst12883 (P2_U3314, P2_R2182_U69);
  not ginst12884 (P2_U3315, P2_R2182_U68);
  not ginst12885 (P2_U3316, P2_R2182_U40);
  not ginst12886 (P2_U3317, P2_R2182_U76);
  nand ginst12887 (P2_U3318, P2_R2182_U68, P2_R2182_U69);
  nand ginst12888 (P2_U3319, P2_U3314, P2_U3352);
  nand ginst12889 (P2_U3320, P2_U2461, P2_U4636);
  not ginst12890 (P2_U3321, P2_R2099_U95);
  not ginst12891 (P2_U3322, P2_R2099_U96);
  not ginst12892 (P2_U3323, P2_R2099_U94);
  not ginst12893 (P2_U3324, P2_R2099_U5);
  nand ginst12894 (P2_U3325, P2_U3312, P2_U4651);
  nand ginst12895 (P2_U3326, P2_U3312, P2_U3570);
  not ginst12896 (P2_U3327, P2_INSTQUEUE_REG_15__7__SCAN_IN);
  not ginst12897 (P2_U3328, P2_INSTQUEUE_REG_15__6__SCAN_IN);
  not ginst12898 (P2_U3329, P2_INSTQUEUE_REG_15__5__SCAN_IN);
  not ginst12899 (P2_U3330, P2_INSTQUEUE_REG_15__4__SCAN_IN);
  not ginst12900 (P2_U3331, P2_INSTQUEUE_REG_15__3__SCAN_IN);
  not ginst12901 (P2_U3332, P2_INSTQUEUE_REG_15__2__SCAN_IN);
  not ginst12902 (P2_U3333, P2_INSTQUEUE_REG_15__1__SCAN_IN);
  not ginst12903 (P2_U3334, P2_INSTQUEUE_REG_15__0__SCAN_IN);
  nand ginst12904 (P2_U3335, P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN, P2_U3307);
  nand ginst12905 (P2_U3336, P2_U2464, P2_U4649);
  nand ginst12906 (P2_U3337, P2_R2182_U68, P2_U3314);
  nand ginst12907 (P2_U3338, P2_R2182_U69, P2_U3352);
  nand ginst12908 (P2_U3339, P2_U2461, P2_U4709);
  nand ginst12909 (P2_U3340, P2_U3336, P2_U3569);
  not ginst12910 (P2_U3341, P2_INSTQUEUE_REG_14__7__SCAN_IN);
  not ginst12911 (P2_U3342, P2_INSTQUEUE_REG_14__6__SCAN_IN);
  not ginst12912 (P2_U3343, P2_INSTQUEUE_REG_14__5__SCAN_IN);
  not ginst12913 (P2_U3344, P2_INSTQUEUE_REG_14__4__SCAN_IN);
  not ginst12914 (P2_U3345, P2_INSTQUEUE_REG_14__3__SCAN_IN);
  not ginst12915 (P2_U3346, P2_INSTQUEUE_REG_14__2__SCAN_IN);
  not ginst12916 (P2_U3347, P2_INSTQUEUE_REG_14__1__SCAN_IN);
  not ginst12917 (P2_U3348, P2_INSTQUEUE_REG_14__0__SCAN_IN);
  nand ginst12918 (P2_U3349, P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P2_U3308);
  nand ginst12919 (P2_U3350, P2_U2464, P2_U4648);
  nand ginst12920 (P2_U3351, P2_R2182_U69, P2_U3315);
  nand ginst12921 (P2_U3352, P2_U3337, P2_U3351);
  nand ginst12922 (P2_U3353, P2_U3314, P2_U4635);
  nand ginst12923 (P2_U3354, P2_U2461, P2_U4767);
  nand ginst12924 (P2_U3355, P2_U3350, P2_U4770);
  nand ginst12925 (P2_U3356, P2_U3350, P2_U3568);
  not ginst12926 (P2_U3357, P2_INSTQUEUE_REG_13__7__SCAN_IN);
  not ginst12927 (P2_U3358, P2_INSTQUEUE_REG_13__6__SCAN_IN);
  not ginst12928 (P2_U3359, P2_INSTQUEUE_REG_13__5__SCAN_IN);
  not ginst12929 (P2_U3360, P2_INSTQUEUE_REG_13__4__SCAN_IN);
  not ginst12930 (P2_U3361, P2_INSTQUEUE_REG_13__3__SCAN_IN);
  not ginst12931 (P2_U3362, P2_INSTQUEUE_REG_13__2__SCAN_IN);
  not ginst12932 (P2_U3363, P2_INSTQUEUE_REG_13__1__SCAN_IN);
  not ginst12933 (P2_U3364, P2_INSTQUEUE_REG_13__0__SCAN_IN);
  nand ginst12934 (P2_U3365, P2_U2464, P2_U2478);
  nand ginst12935 (P2_U3366, P2_U2461, P2_U2475);
  nand ginst12936 (P2_U3367, P2_U3365, P2_U3567);
  not ginst12937 (P2_U3368, P2_INSTQUEUE_REG_12__7__SCAN_IN);
  not ginst12938 (P2_U3369, P2_INSTQUEUE_REG_12__6__SCAN_IN);
  not ginst12939 (P2_U3370, P2_INSTQUEUE_REG_12__5__SCAN_IN);
  not ginst12940 (P2_U3371, P2_INSTQUEUE_REG_12__4__SCAN_IN);
  not ginst12941 (P2_U3372, P2_INSTQUEUE_REG_12__3__SCAN_IN);
  not ginst12942 (P2_U3373, P2_INSTQUEUE_REG_12__2__SCAN_IN);
  not ginst12943 (P2_U3374, P2_INSTQUEUE_REG_12__1__SCAN_IN);
  not ginst12944 (P2_U3375, P2_INSTQUEUE_REG_12__0__SCAN_IN);
  nand ginst12945 (P2_U3376, P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN, P2_U3310);
  nand ginst12946 (P2_U3377, P2_U4642, P2_U4645);
  nand ginst12947 (P2_U3378, P2_R2182_U76, P2_U3316);
  nand ginst12948 (P2_U3379, P2_U2481, P2_U4636);
  nand ginst12949 (P2_U3380, P2_U3377, P2_U4885);
  nand ginst12950 (P2_U3381, P2_U3377, P2_U3566);
  not ginst12951 (P2_U3382, P2_INSTQUEUE_REG_11__7__SCAN_IN);
  not ginst12952 (P2_U3383, P2_INSTQUEUE_REG_11__6__SCAN_IN);
  not ginst12953 (P2_U3384, P2_INSTQUEUE_REG_11__5__SCAN_IN);
  not ginst12954 (P2_U3385, P2_INSTQUEUE_REG_11__4__SCAN_IN);
  not ginst12955 (P2_U3386, P2_INSTQUEUE_REG_11__3__SCAN_IN);
  not ginst12956 (P2_U3387, P2_INSTQUEUE_REG_11__2__SCAN_IN);
  not ginst12957 (P2_U3388, P2_INSTQUEUE_REG_11__1__SCAN_IN);
  not ginst12958 (P2_U3389, P2_INSTQUEUE_REG_11__0__SCAN_IN);
  nand ginst12959 (P2_U3390, P2_U4645, P2_U4649);
  nand ginst12960 (P2_U3391, P2_U2481, P2_U4709);
  nand ginst12961 (P2_U3392, P2_U3390, P2_U3565);
  not ginst12962 (P2_U3393, P2_INSTQUEUE_REG_10__7__SCAN_IN);
  not ginst12963 (P2_U3394, P2_INSTQUEUE_REG_10__6__SCAN_IN);
  not ginst12964 (P2_U3395, P2_INSTQUEUE_REG_10__5__SCAN_IN);
  not ginst12965 (P2_U3396, P2_INSTQUEUE_REG_10__4__SCAN_IN);
  not ginst12966 (P2_U3397, P2_INSTQUEUE_REG_10__3__SCAN_IN);
  not ginst12967 (P2_U3398, P2_INSTQUEUE_REG_10__2__SCAN_IN);
  not ginst12968 (P2_U3399, P2_INSTQUEUE_REG_10__1__SCAN_IN);
  not ginst12969 (P2_U3400, P2_INSTQUEUE_REG_10__0__SCAN_IN);
  nand ginst12970 (P2_U3401, P2_U4645, P2_U4648);
  nand ginst12971 (P2_U3402, P2_U2481, P2_U4767);
  nand ginst12972 (P2_U3403, P2_U3401, P2_U5000);
  nand ginst12973 (P2_U3404, P2_U3401, P2_U3564);
  not ginst12974 (P2_U3405, P2_INSTQUEUE_REG_9__7__SCAN_IN);
  not ginst12975 (P2_U3406, P2_INSTQUEUE_REG_9__6__SCAN_IN);
  not ginst12976 (P2_U3407, P2_INSTQUEUE_REG_9__5__SCAN_IN);
  not ginst12977 (P2_U3408, P2_INSTQUEUE_REG_9__4__SCAN_IN);
  not ginst12978 (P2_U3409, P2_INSTQUEUE_REG_9__3__SCAN_IN);
  not ginst12979 (P2_U3410, P2_INSTQUEUE_REG_9__2__SCAN_IN);
  not ginst12980 (P2_U3411, P2_INSTQUEUE_REG_9__1__SCAN_IN);
  not ginst12981 (P2_U3412, P2_INSTQUEUE_REG_9__0__SCAN_IN);
  nand ginst12982 (P2_U3413, P2_U2478, P2_U4645);
  nand ginst12983 (P2_U3414, P2_U2475, P2_U2481);
  nand ginst12984 (P2_U3415, P2_U3413, P2_U3563);
  not ginst12985 (P2_U3416, P2_INSTQUEUE_REG_8__7__SCAN_IN);
  not ginst12986 (P2_U3417, P2_INSTQUEUE_REG_8__6__SCAN_IN);
  not ginst12987 (P2_U3418, P2_INSTQUEUE_REG_8__5__SCAN_IN);
  not ginst12988 (P2_U3419, P2_INSTQUEUE_REG_8__4__SCAN_IN);
  not ginst12989 (P2_U3420, P2_INSTQUEUE_REG_8__3__SCAN_IN);
  not ginst12990 (P2_U3421, P2_INSTQUEUE_REG_8__2__SCAN_IN);
  not ginst12991 (P2_U3422, P2_INSTQUEUE_REG_8__1__SCAN_IN);
  not ginst12992 (P2_U3423, P2_INSTQUEUE_REG_8__0__SCAN_IN);
  nand ginst12993 (P2_U3424, P2_U2465, P2_U4642);
  nand ginst12994 (P2_U3425, P2_U2460, P2_U4637);
  nand ginst12995 (P2_U3426, P2_U3378, P2_U3425, P2_U4639);
  nand ginst12996 (P2_U3427, P2_U2491, P2_U4636);
  nand ginst12997 (P2_U3428, P2_U3376, P2_U3424, P2_U4646);
  nand ginst12998 (P2_U3429, P2_U3424, P2_U5114);
  nand ginst12999 (P2_U3430, P2_U3424, P2_U3562);
  not ginst13000 (P2_U3431, P2_INSTQUEUE_REG_7__7__SCAN_IN);
  not ginst13001 (P2_U3432, P2_INSTQUEUE_REG_7__6__SCAN_IN);
  not ginst13002 (P2_U3433, P2_INSTQUEUE_REG_7__5__SCAN_IN);
  not ginst13003 (P2_U3434, P2_INSTQUEUE_REG_7__4__SCAN_IN);
  not ginst13004 (P2_U3435, P2_INSTQUEUE_REG_7__3__SCAN_IN);
  not ginst13005 (P2_U3436, P2_INSTQUEUE_REG_7__2__SCAN_IN);
  not ginst13006 (P2_U3437, P2_INSTQUEUE_REG_7__1__SCAN_IN);
  not ginst13007 (P2_U3438, P2_INSTQUEUE_REG_7__0__SCAN_IN);
  nand ginst13008 (P2_U3439, P2_U2465, P2_U4649);
  nand ginst13009 (P2_U3440, P2_U2491, P2_U4709);
  nand ginst13010 (P2_U3441, P2_U3439, P2_U3561);
  not ginst13011 (P2_U3442, P2_INSTQUEUE_REG_6__7__SCAN_IN);
  not ginst13012 (P2_U3443, P2_INSTQUEUE_REG_6__6__SCAN_IN);
  not ginst13013 (P2_U3444, P2_INSTQUEUE_REG_6__5__SCAN_IN);
  not ginst13014 (P2_U3445, P2_INSTQUEUE_REG_6__4__SCAN_IN);
  not ginst13015 (P2_U3446, P2_INSTQUEUE_REG_6__3__SCAN_IN);
  not ginst13016 (P2_U3447, P2_INSTQUEUE_REG_6__2__SCAN_IN);
  not ginst13017 (P2_U3448, P2_INSTQUEUE_REG_6__1__SCAN_IN);
  not ginst13018 (P2_U3449, P2_INSTQUEUE_REG_6__0__SCAN_IN);
  nand ginst13019 (P2_U3450, P2_U2465, P2_U4648);
  nand ginst13020 (P2_U3451, P2_U2491, P2_U4767);
  nand ginst13021 (P2_U3452, P2_U3450, P2_U5228);
  nand ginst13022 (P2_U3453, P2_U3450, P2_U3560);
  not ginst13023 (P2_U3454, P2_INSTQUEUE_REG_5__7__SCAN_IN);
  not ginst13024 (P2_U3455, P2_INSTQUEUE_REG_5__6__SCAN_IN);
  not ginst13025 (P2_U3456, P2_INSTQUEUE_REG_5__5__SCAN_IN);
  not ginst13026 (P2_U3457, P2_INSTQUEUE_REG_5__4__SCAN_IN);
  not ginst13027 (P2_U3458, P2_INSTQUEUE_REG_5__3__SCAN_IN);
  not ginst13028 (P2_U3459, P2_INSTQUEUE_REG_5__2__SCAN_IN);
  not ginst13029 (P2_U3460, P2_INSTQUEUE_REG_5__1__SCAN_IN);
  not ginst13030 (P2_U3461, P2_INSTQUEUE_REG_5__0__SCAN_IN);
  nand ginst13031 (P2_U3462, P2_U2465, P2_U2478);
  nand ginst13032 (P2_U3463, P2_U2475, P2_U2491);
  nand ginst13033 (P2_U3464, P2_U3462, P2_U3559);
  not ginst13034 (P2_U3465, P2_INSTQUEUE_REG_4__7__SCAN_IN);
  not ginst13035 (P2_U3466, P2_INSTQUEUE_REG_4__6__SCAN_IN);
  not ginst13036 (P2_U3467, P2_INSTQUEUE_REG_4__5__SCAN_IN);
  not ginst13037 (P2_U3468, P2_INSTQUEUE_REG_4__4__SCAN_IN);
  not ginst13038 (P2_U3469, P2_INSTQUEUE_REG_4__3__SCAN_IN);
  not ginst13039 (P2_U3470, P2_INSTQUEUE_REG_4__2__SCAN_IN);
  not ginst13040 (P2_U3471, P2_INSTQUEUE_REG_4__1__SCAN_IN);
  not ginst13041 (P2_U3472, P2_INSTQUEUE_REG_4__0__SCAN_IN);
  nand ginst13042 (P2_U3473, P2_U2503, P2_U4642);
  nand ginst13043 (P2_U3474, P2_U2500, P2_U4636);
  nand ginst13044 (P2_U3475, P2_U3473, P2_U5343);
  nand ginst13045 (P2_U3476, P2_U3473, P2_U3558);
  not ginst13046 (P2_U3477, P2_INSTQUEUE_REG_3__7__SCAN_IN);
  not ginst13047 (P2_U3478, P2_INSTQUEUE_REG_3__6__SCAN_IN);
  not ginst13048 (P2_U3479, P2_INSTQUEUE_REG_3__5__SCAN_IN);
  not ginst13049 (P2_U3480, P2_INSTQUEUE_REG_3__4__SCAN_IN);
  not ginst13050 (P2_U3481, P2_INSTQUEUE_REG_3__3__SCAN_IN);
  not ginst13051 (P2_U3482, P2_INSTQUEUE_REG_3__2__SCAN_IN);
  not ginst13052 (P2_U3483, P2_INSTQUEUE_REG_3__1__SCAN_IN);
  not ginst13053 (P2_U3484, P2_INSTQUEUE_REG_3__0__SCAN_IN);
  nand ginst13054 (P2_U3485, P2_U2503, P2_U4649);
  nand ginst13055 (P2_U3486, P2_U2500, P2_U4709);
  nand ginst13056 (P2_U3487, P2_U3485, P2_U3557);
  not ginst13057 (P2_U3488, P2_INSTQUEUE_REG_2__7__SCAN_IN);
  not ginst13058 (P2_U3489, P2_INSTQUEUE_REG_2__6__SCAN_IN);
  not ginst13059 (P2_U3490, P2_INSTQUEUE_REG_2__5__SCAN_IN);
  not ginst13060 (P2_U3491, P2_INSTQUEUE_REG_2__4__SCAN_IN);
  not ginst13061 (P2_U3492, P2_INSTQUEUE_REG_2__3__SCAN_IN);
  not ginst13062 (P2_U3493, P2_INSTQUEUE_REG_2__2__SCAN_IN);
  not ginst13063 (P2_U3494, P2_INSTQUEUE_REG_2__1__SCAN_IN);
  not ginst13064 (P2_U3495, P2_INSTQUEUE_REG_2__0__SCAN_IN);
  nand ginst13065 (P2_U3496, P2_U2503, P2_U4648);
  nand ginst13066 (P2_U3497, P2_U2500, P2_U4767);
  nand ginst13067 (P2_U3498, P2_U3496, P2_U5458);
  nand ginst13068 (P2_U3499, P2_U3496, P2_U3556);
  not ginst13069 (P2_U3500, P2_INSTQUEUE_REG_1__7__SCAN_IN);
  not ginst13070 (P2_U3501, P2_INSTQUEUE_REG_1__6__SCAN_IN);
  not ginst13071 (P2_U3502, P2_INSTQUEUE_REG_1__5__SCAN_IN);
  not ginst13072 (P2_U3503, P2_INSTQUEUE_REG_1__4__SCAN_IN);
  not ginst13073 (P2_U3504, P2_INSTQUEUE_REG_1__3__SCAN_IN);
  not ginst13074 (P2_U3505, P2_INSTQUEUE_REG_1__2__SCAN_IN);
  not ginst13075 (P2_U3506, P2_INSTQUEUE_REG_1__1__SCAN_IN);
  not ginst13076 (P2_U3507, P2_INSTQUEUE_REG_1__0__SCAN_IN);
  nand ginst13077 (P2_U3508, P2_U2478, P2_U2503);
  nand ginst13078 (P2_U3509, P2_U2475, P2_U2500);
  nand ginst13079 (P2_U3510, P2_U3508, P2_U3555);
  not ginst13080 (P2_U3511, P2_INSTQUEUE_REG_0__7__SCAN_IN);
  not ginst13081 (P2_U3512, P2_INSTQUEUE_REG_0__6__SCAN_IN);
  not ginst13082 (P2_U3513, P2_INSTQUEUE_REG_0__5__SCAN_IN);
  not ginst13083 (P2_U3514, P2_INSTQUEUE_REG_0__4__SCAN_IN);
  not ginst13084 (P2_U3515, P2_INSTQUEUE_REG_0__3__SCAN_IN);
  not ginst13085 (P2_U3516, P2_INSTQUEUE_REG_0__2__SCAN_IN);
  not ginst13086 (P2_U3517, P2_INSTQUEUE_REG_0__1__SCAN_IN);
  not ginst13087 (P2_U3518, P2_INSTQUEUE_REG_0__0__SCAN_IN);
  not ginst13088 (P2_U3519, P2_FLUSH_REG_SCAN_IN);
  not ginst13089 (P2_U3520, P2_R2088_U6);
  nand ginst13090 (P2_U3521, P2_U3697, P2_U3698);
  nand ginst13091 (P2_U3522, P2_U2451, P2_U4429);
  nand ginst13092 (P2_U3523, P2_U4427, P2_U4475);
  nand ginst13093 (P2_U3524, P2_U4429, P2_U4475);
  nand ginst13094 (P2_U3525, P2_U3279, P2_U7863, P2_U7865, P2_U7869);
  not ginst13095 (P2_U3526, P2_R2147_U8);
  nand ginst13096 (P2_U3527, P2_U3283, P2_U3289);
  not ginst13097 (P2_U3528, P2_U3647);
  not ginst13098 (P2_U3529, P2_R2147_U9);
  nand ginst13099 (P2_U3530, P2_U3274, P2_U5615);
  not ginst13100 (P2_U3531, P2_R2147_U4);
  not ginst13101 (P2_U3532, P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN);
  nand ginst13102 (P2_U3533, P2_U3306, P2_U4455, P2_U5642);
  nand ginst13103 (P2_U3534, P2_U3269, P2_U4430);
  nand ginst13104 (P2_U3535, P2_U5671, P2_U5672);
  nand ginst13105 (P2_U3536, P2_STATE2_REG_0__SCAN_IN, P2_U7873);
  nand ginst13106 (P2_U3537, P2_U5936, P2_U5937);
  nand ginst13107 (P2_U3538, P2_U2446, P2_U4055);
  nand ginst13108 (P2_U3539, P2_U2357, P2_U4056);
  nand ginst13109 (P2_U3540, P2_STATE2_REG_2__SCAN_IN, P2_U3284);
  nand ginst13110 (P2_U3541, P2_U6230, P2_U6231);
  nand ginst13111 (P2_U3542, P2_U2374, P2_U6326);
  nand ginst13112 (P2_U3543, P2_U2374, P2_U6470);
  not ginst13113 (P2_U3544, P2_EBX_REG_31__SCAN_IN);
  or ginst13114 (P2_U3545, P2_STATEBS16_REG_SCAN_IN, U211);
  nand ginst13115 (P2_U3546, P2_U4069, P2_U4462);
  nand ginst13116 (P2_U3547, P2_U4171, P2_U4174, P2_U4177, P2_U4181);
  nand ginst13117 (P2_U3548, P2_REIP_REG_1__SCAN_IN, P2_U4438);
  nand ginst13118 (P2_U3549, P2_U2356, P2_U4420);
  nand ginst13119 (P2_U3550, P2_STATE2_REG_0__SCAN_IN, P2_U4427);
  not ginst13120 (P2_U3551, P2_CODEFETCH_REG_SCAN_IN);
  not ginst13121 (P2_U3552, P2_READREQUEST_REG_SCAN_IN);
  nand ginst13122 (P2_U3553, P2_U3275, P2_U4405);
  nand ginst13123 (P2_U3554, P2_U3576, P2_U4415);
  nand ginst13124 (P2_U3555, P2_U2479, P2_U2504);
  nand ginst13125 (P2_U3556, P2_U2473, P2_U2504);
  nand ginst13126 (P2_U3557, P2_U2470, P2_U2504);
  nand ginst13127 (P2_U3558, P2_U2467, P2_U2504);
  nand ginst13128 (P2_U3559, P2_U2479, P2_U2492);
  nand ginst13129 (P2_U3560, P2_U2473, P2_U2492);
  nand ginst13130 (P2_U3561, P2_U2470, P2_U2492);
  nand ginst13131 (P2_U3562, P2_U2467, P2_U2492);
  nand ginst13132 (P2_U3563, P2_U2479, P2_U2483);
  nand ginst13133 (P2_U3564, P2_U2473, P2_U2483);
  nand ginst13134 (P2_U3565, P2_U2470, P2_U2483);
  nand ginst13135 (P2_U3566, P2_U2467, P2_U2483);
  nand ginst13136 (P2_U3567, P2_U2466, P2_U2479);
  nand ginst13137 (P2_U3568, P2_U2466, P2_U2473);
  nand ginst13138 (P2_U3569, P2_U2466, P2_U2470);
  nand ginst13139 (P2_U3570, P2_U2466, P2_U2467);
  nand ginst13140 (P2_U3571, P2_U3300, P2_U7865);
  not ginst13141 (P2_U3572, P2_U3242);
  or ginst13142 (P2_U3573, P2_STATE2_REG_1__SCAN_IN, P2_STATE2_REG_0__SCAN_IN);
  nand ginst13143 (P2_U3574, P2_U3295, P2_U3521, P2_U5571);
  nand ginst13144 (P2_U3575, P2_U4419, P2_U7871);
  nand ginst13145 (P2_U3576, P2_U3279, P2_U4419);
  nand ginst13146 (P2_U3577, P2_U4424, P2_U6845);
  nand ginst13147 (P2_U3578, P2_U2590, P2_U4428);
  nand ginst13148 (P2_U3579, P2_U8062, P2_U8063);
  nand ginst13149 (P2_U3580, P2_U8065, P2_U8066);
  nand ginst13150 (P2_U3581, P2_U8080, P2_U8081);
  nand ginst13151 (P2_U3582, P2_U8098, P2_U8099);
  nand ginst13152 (P2_U3583, P2_U8147, P2_U8148);
  nand ginst13153 (P2_U3584, P2_U8150, P2_U8151);
  nand ginst13154 (P2_U3585, P2_U7899, P2_U7900);
  nand ginst13155 (P2_U3586, P2_U7901, P2_U7902);
  nand ginst13156 (P2_U3587, P2_U7903, P2_U7904);
  nand ginst13157 (P2_U3588, P2_U7905, P2_U7906);
  nand ginst13158 (P2_U3589, P2_U7915, P2_U7916);
  and ginst13159 (P2_U3590, P2_U3263, P2_U4401);
  nand ginst13160 (P2_U3591, P2_U7918, P2_U7919);
  nand ginst13161 (P2_U3592, P2_U7920, P2_U7921);
  nand ginst13162 (P2_U3593, P2_U8058, P2_U8059);
  and ginst13163 (P2_U3594, P2_U3866, P2_U4434);
  nand ginst13164 (P2_U3595, P2_U8072, P2_U8073);
  nand ginst13165 (P2_U3596, P2_U8083, P2_U8084);
  nand ginst13166 (P2_U3597, P2_U8085, P2_U8086);
  nand ginst13167 (P2_U3598, P2_U8088, P2_U8089);
  nand ginst13168 (P2_U3599, P2_U8093, P2_U8094);
  nand ginst13169 (P2_U3600, P2_U8101, P2_U8102);
  nand ginst13170 (P2_U3601, P2_U8103, P2_U8104);
  nand ginst13171 (P2_U3602, P2_U8105, P2_U8106);
  nand ginst13172 (P2_U3603, P2_U8110, P2_U8111);
  nand ginst13173 (P2_U3604, P2_U8112, P2_U8113);
  nand ginst13174 (P2_U3605, P2_U8114, P2_U8115);
  nor ginst13175 (P2_U3606, P2_DATAWIDTH_REG_1__SCAN_IN, P2_REIP_REG_1__SCAN_IN);
  and ginst13176 (P2_U3607, P2_U4183, P2_U7898);
  nand ginst13177 (P2_U3608, P2_U8129, P2_U8130);
  nand ginst13178 (P2_U3609, P2_U8133, P2_U8134);
  nand ginst13179 (P2_U3610, P2_U8137, P2_U8138);
  nand ginst13180 (P2_U3611, P2_U8141, P2_U8142);
  nand ginst13181 (P2_U3612, P2_U8143, P2_U8144);
  nand ginst13182 (P2_U3613, P2_U8281, P2_U8282);
  nand ginst13183 (P2_U3614, P2_U8283, P2_U8284);
  nand ginst13184 (P2_U3615, P2_U8285, P2_U8286);
  and ginst13185 (P2_U3616, P2_R2147_U7, P2_U4434);
  nand ginst13186 (P2_U3617, P2_U8287, P2_U8288);
  nand ginst13187 (P2_U3618, P2_U8289, P2_U8290);
  nand ginst13188 (P2_U3619, P2_U8291, P2_U8292);
  nand ginst13189 (P2_U3620, P2_U8293, P2_U8294);
  nand ginst13190 (P2_U3621, P2_U8295, P2_U8296);
  nand ginst13191 (P2_U3622, P2_U8297, P2_U8298);
  nand ginst13192 (P2_U3623, P2_U8299, P2_U8300);
  nand ginst13193 (P2_U3624, P2_U8301, P2_U8302);
  nand ginst13194 (P2_U3625, P2_U8303, P2_U8304);
  nand ginst13195 (P2_U3626, P2_U8305, P2_U8306);
  nand ginst13196 (P2_U3627, P2_U8307, P2_U8308);
  nand ginst13197 (P2_U3628, P2_U8309, P2_U8310);
  nand ginst13198 (P2_U3629, P2_U8311, P2_U8312);
  nand ginst13199 (P2_U3630, P2_U8313, P2_U8314);
  nand ginst13200 (P2_U3631, P2_U8315, P2_U8316);
  nand ginst13201 (P2_U3632, P2_U8317, P2_U8318);
  nand ginst13202 (P2_U3633, P2_U8319, P2_U8320);
  nand ginst13203 (P2_U3634, P2_U8321, P2_U8322);
  nand ginst13204 (P2_U3635, P2_U8323, P2_U8324);
  nand ginst13205 (P2_U3636, P2_U8325, P2_U8326);
  nand ginst13206 (P2_U3637, P2_U8327, P2_U8328);
  nand ginst13207 (P2_U3638, P2_U8329, P2_U8330);
  nand ginst13208 (P2_U3639, P2_U8331, P2_U8332);
  nand ginst13209 (P2_U3640, P2_U8333, P2_U8334);
  nand ginst13210 (P2_U3641, P2_U8335, P2_U8336);
  nand ginst13211 (P2_U3642, P2_U8337, P2_U8338);
  nand ginst13212 (P2_U3643, P2_U8339, P2_U8340);
  nand ginst13213 (P2_U3644, P2_U8341, P2_U8342);
  nand ginst13214 (P2_U3645, P2_U8343, P2_U8344);
  nand ginst13215 (P2_U3646, P2_U8345, P2_U8346);
  nand ginst13216 (P2_U3647, P2_U8349, P2_U8350);
  nand ginst13217 (P2_U3648, P2_U8351, P2_U8352);
  nand ginst13218 (P2_U3649, P2_U8353, P2_U8354);
  nand ginst13219 (P2_U3650, P2_U8355, P2_U8356);
  nand ginst13220 (P2_U3651, P2_U8357, P2_U8358);
  nand ginst13221 (P2_U3652, P2_U8359, P2_U8360);
  nand ginst13222 (P2_U3653, P2_U8361, P2_U8362);
  nand ginst13223 (P2_U3654, P2_U8363, P2_U8364);
  nand ginst13224 (P2_U3655, P2_U8365, P2_U8366);
  nand ginst13225 (P2_U3656, P2_U8367, P2_U8368);
  nand ginst13226 (P2_U3657, P2_U8369, P2_U8370);
  nand ginst13227 (P2_U3658, P2_U8371, P2_U8372);
  nand ginst13228 (P2_U3659, P2_U8373, P2_U8374);
  nand ginst13229 (P2_U3660, P2_U8375, P2_U8376);
  nand ginst13230 (P2_U3661, P2_U8377, P2_U8378);
  nand ginst13231 (P2_U3662, P2_U8379, P2_U8380);
  nand ginst13232 (P2_U3663, P2_U8381, P2_U8382);
  nand ginst13233 (P2_U3664, P2_U8383, P2_U8384);
  nand ginst13234 (P2_U3665, P2_U8385, P2_U8386);
  nand ginst13235 (P2_U3666, P2_U8387, P2_U8388);
  nand ginst13236 (P2_U3667, P2_U8389, P2_U8390);
  nand ginst13237 (P2_U3668, P2_U8391, P2_U8392);
  nand ginst13238 (P2_U3669, P2_U8393, P2_U8394);
  nand ginst13239 (P2_U3670, P2_U8395, P2_U8396);
  nand ginst13240 (P2_U3671, P2_U8397, P2_U8398);
  nand ginst13241 (P2_U3672, P2_U8399, P2_U8400);
  nand ginst13242 (P2_U3673, P2_U8401, P2_U8402);
  nand ginst13243 (P2_U3674, P2_U8403, P2_U8404);
  nand ginst13244 (P2_U3675, P2_U8405, P2_U8406);
  nand ginst13245 (P2_U3676, P2_U8407, P2_U8408);
  nand ginst13246 (P2_U3677, P2_U8409, P2_U8410);
  nand ginst13247 (P2_U3678, P2_U8411, P2_U8412);
  nand ginst13248 (P2_U3679, P2_U8413, P2_U8414);
  nand ginst13249 (P2_U3680, P2_U8415, P2_U8416);
  nand ginst13250 (P2_U3681, P2_U8417, P2_U8418);
  nand ginst13251 (P2_U3682, P2_U8419, P2_U8420);
  nand ginst13252 (P2_U3683, P2_U8421, P2_U8422);
  nand ginst13253 (P2_U3684, P2_U8423, P2_U8424);
  nand ginst13254 (P2_U3685, P2_U8425, P2_U8426);
  nand ginst13255 (P2_U3686, P2_U8427, P2_U8428);
  nand ginst13256 (P2_U3687, P2_U8429, P2_U8430);
  nand ginst13257 (P2_U3688, P2_U8431, P2_U8432);
  nand ginst13258 (P2_U3689, P2_U8433, P2_U8434);
  and ginst13259 (P2_U3690, P2_U3261, P2_U4578);
  and ginst13260 (P2_U3691, P2_U3260, P2_U4583);
  and ginst13261 (P2_U3692, P2_STATE_REG_0__SCAN_IN, P2_REQUESTPENDING_REG_SCAN_IN);
  and ginst13262 (P2_U3693, P2_U7751, P2_U7767, P2_U7783, P2_U7799);
  and ginst13263 (P2_U3694, P2_U7815, P2_U7831, P2_U7847, P2_U7868);
  and ginst13264 (P2_U3695, P2_U7750, P2_U7766, P2_U7782, P2_U7798);
  and ginst13265 (P2_U3696, P2_U7814, P2_U7830, P2_U7846, P2_U7866);
  and ginst13266 (P2_U3697, P2_U7749, P2_U7765, P2_U7781, P2_U7797);
  and ginst13267 (P2_U3698, P2_U7813, P2_U7829, P2_U7845, P2_U7864);
  and ginst13268 (P2_U3699, P2_U7748, P2_U7764, P2_U7780, P2_U7796);
  and ginst13269 (P2_U3700, P2_U7812, P2_U7828, P2_U7844, P2_U7862);
  and ginst13270 (P2_U3701, P2_U7747, P2_U7763, P2_U7779, P2_U7795);
  and ginst13271 (P2_U3702, P2_U7811, P2_U7827, P2_U7843, P2_U7860);
  and ginst13272 (P2_U3703, P2_U7746, P2_U7762, P2_U7778, P2_U7794);
  and ginst13273 (P2_U3704, P2_U7810, P2_U7826, P2_U7842, P2_U7858);
  and ginst13274 (P2_U3705, P2_U7753, P2_U7769, P2_U7785, P2_U7801);
  and ginst13275 (P2_U3706, P2_U7817, P2_U7833, P2_U7849, P2_U7872);
  and ginst13276 (P2_U3707, P2_U7752, P2_U7768, P2_U7784, P2_U7800);
  and ginst13277 (P2_U3708, P2_U7816, P2_U7832, P2_U7848, P2_U7870);
  and ginst13278 (P2_U3709, P2_U3710, P2_U4417);
  and ginst13279 (P2_U3710, P2_STATE2_REG_0__SCAN_IN, P2_U4595);
  and ginst13280 (P2_U3711, P2_U2360, P2_U3266);
  and ginst13281 (P2_U3712, P2_U3521, P2_U7867);
  and ginst13282 (P2_U3713, P2_U4598, P2_U4599);
  and ginst13283 (P2_U3714, P2_STATE2_REG_2__SCAN_IN, P2_U3573);
  and ginst13284 (P2_U3715, P2_U3714, P2_U4618);
  and ginst13285 (P2_U3716, P2_U3304, P2_U4624);
  and ginst13286 (P2_U3717, P2_U3265, P2_U4466);
  and ginst13287 (P2_U3718, P2_STATE2_REG_3__SCAN_IN, P2_U3269);
  nor ginst13288 (P2_U3719, P2_STATE2_REG_2__SCAN_IN, P2_STATE2_REG_1__SCAN_IN);
  and ginst13289 (P2_U3720, P2_U4453, P2_U4465);
  and ginst13290 (P2_U3721, P2_U3720, P2_U4632);
  and ginst13291 (P2_U3722, P2_U4443, P2_U4661, P2_U4662);
  and ginst13292 (P2_U3723, P2_U4669, P2_U4670, P2_U4671);
  and ginst13293 (P2_U3724, P2_U4674, P2_U4675, P2_U4676);
  and ginst13294 (P2_U3725, P2_U4679, P2_U4680, P2_U4681);
  and ginst13295 (P2_U3726, P2_U4684, P2_U4685, P2_U4686);
  and ginst13296 (P2_U3727, P2_U4689, P2_U4690, P2_U4691);
  and ginst13297 (P2_U3728, P2_U4694, P2_U4695, P2_U4696);
  and ginst13298 (P2_U3729, P2_U4699, P2_U4700, P2_U4701);
  and ginst13299 (P2_U3730, P2_U4704, P2_U4705, P2_U4706);
  and ginst13300 (P2_U3731, P2_U4443, P2_U4719, P2_U4720);
  and ginst13301 (P2_U3732, P2_U4727, P2_U4728, P2_U4729);
  and ginst13302 (P2_U3733, P2_U4732, P2_U4733, P2_U4734);
  and ginst13303 (P2_U3734, P2_U4737, P2_U4738, P2_U4739);
  and ginst13304 (P2_U3735, P2_U4742, P2_U4743, P2_U4744);
  and ginst13305 (P2_U3736, P2_U4747, P2_U4748, P2_U4749);
  and ginst13306 (P2_U3737, P2_U4752, P2_U4753, P2_U4754);
  and ginst13307 (P2_U3738, P2_U4757, P2_U4758, P2_U4759);
  and ginst13308 (P2_U3739, P2_U4762, P2_U4763, P2_U4764);
  and ginst13309 (P2_U3740, P2_U4443, P2_U4778, P2_U4779);
  and ginst13310 (P2_U3741, P2_U4786, P2_U4787, P2_U4788);
  and ginst13311 (P2_U3742, P2_U4791, P2_U4792, P2_U4793);
  and ginst13312 (P2_U3743, P2_U4796, P2_U4797, P2_U4798);
  and ginst13313 (P2_U3744, P2_U4801, P2_U4802, P2_U4803);
  and ginst13314 (P2_U3745, P2_U4806, P2_U4807, P2_U4808);
  and ginst13315 (P2_U3746, P2_U4811, P2_U4812, P2_U4813);
  and ginst13316 (P2_U3747, P2_U4816, P2_U4817, P2_U4818);
  and ginst13317 (P2_U3748, P2_U4821, P2_U4822, P2_U4823);
  and ginst13318 (P2_U3749, P2_U4443, P2_U4835, P2_U4836);
  and ginst13319 (P2_U3750, P2_U4843, P2_U4844, P2_U4845);
  and ginst13320 (P2_U3751, P2_U4848, P2_U4849, P2_U4850);
  and ginst13321 (P2_U3752, P2_U4853, P2_U4854, P2_U4855);
  and ginst13322 (P2_U3753, P2_U4858, P2_U4859, P2_U4860);
  and ginst13323 (P2_U3754, P2_U4863, P2_U4864, P2_U4865);
  and ginst13324 (P2_U3755, P2_U4868, P2_U4869, P2_U4870);
  and ginst13325 (P2_U3756, P2_U4873, P2_U4874, P2_U4875);
  and ginst13326 (P2_U3757, P2_U4878, P2_U4879, P2_U4880);
  and ginst13327 (P2_U3758, P2_U4443, P2_U4893, P2_U4894);
  and ginst13328 (P2_U3759, P2_U4901, P2_U4902, P2_U4903);
  and ginst13329 (P2_U3760, P2_U4906, P2_U4907, P2_U4908);
  and ginst13330 (P2_U3761, P2_U4911, P2_U4912, P2_U4913);
  and ginst13331 (P2_U3762, P2_U4916, P2_U4917, P2_U4918);
  and ginst13332 (P2_U3763, P2_U4921, P2_U4922, P2_U4923);
  and ginst13333 (P2_U3764, P2_U4926, P2_U4927, P2_U4928);
  and ginst13334 (P2_U3765, P2_U4931, P2_U4932, P2_U4933);
  and ginst13335 (P2_U3766, P2_U4936, P2_U4937, P2_U4938);
  and ginst13336 (P2_U3767, P2_U4443, P2_U4950, P2_U4951);
  and ginst13337 (P2_U3768, P2_U4958, P2_U4959, P2_U4960);
  and ginst13338 (P2_U3769, P2_U4963, P2_U4964, P2_U4965);
  and ginst13339 (P2_U3770, P2_U4968, P2_U4969, P2_U4970);
  and ginst13340 (P2_U3771, P2_U4973, P2_U4974, P2_U4975);
  and ginst13341 (P2_U3772, P2_U4978, P2_U4979, P2_U4980);
  and ginst13342 (P2_U3773, P2_U4983, P2_U4984, P2_U4985);
  and ginst13343 (P2_U3774, P2_U4988, P2_U4989, P2_U4990);
  and ginst13344 (P2_U3775, P2_U4993, P2_U4994, P2_U4995);
  and ginst13345 (P2_U3776, P2_U4443, P2_U5008, P2_U5009);
  and ginst13346 (P2_U3777, P2_U5016, P2_U5017, P2_U5018);
  and ginst13347 (P2_U3778, P2_U5021, P2_U5022, P2_U5023);
  and ginst13348 (P2_U3779, P2_U5026, P2_U5027, P2_U5028);
  and ginst13349 (P2_U3780, P2_U5031, P2_U5032, P2_U5033);
  and ginst13350 (P2_U3781, P2_U5036, P2_U5037, P2_U5038);
  and ginst13351 (P2_U3782, P2_U5041, P2_U5042, P2_U5043);
  and ginst13352 (P2_U3783, P2_U5046, P2_U5047, P2_U5048);
  and ginst13353 (P2_U3784, P2_U5051, P2_U5052, P2_U5053);
  and ginst13354 (P2_U3785, P2_U4443, P2_U5065, P2_U5066);
  and ginst13355 (P2_U3786, P2_U5073, P2_U5074, P2_U5075);
  and ginst13356 (P2_U3787, P2_U5078, P2_U5079, P2_U5080);
  and ginst13357 (P2_U3788, P2_U5083, P2_U5084, P2_U5085);
  and ginst13358 (P2_U3789, P2_U5088, P2_U5089, P2_U5090);
  and ginst13359 (P2_U3790, P2_U5093, P2_U5094, P2_U5095);
  and ginst13360 (P2_U3791, P2_U5098, P2_U5099, P2_U5100);
  and ginst13361 (P2_U3792, P2_U5103, P2_U5104, P2_U5105);
  and ginst13362 (P2_U3793, P2_U5108, P2_U5109, P2_U5110);
  and ginst13363 (P2_U3794, P2_U4443, P2_U5121, P2_U5122);
  and ginst13364 (P2_U3795, P2_U5129, P2_U5130, P2_U5131);
  and ginst13365 (P2_U3796, P2_U5134, P2_U5135, P2_U5136);
  and ginst13366 (P2_U3797, P2_U5139, P2_U5140, P2_U5141);
  and ginst13367 (P2_U3798, P2_U5144, P2_U5145, P2_U5146);
  and ginst13368 (P2_U3799, P2_U5149, P2_U5150, P2_U5151);
  and ginst13369 (P2_U3800, P2_U5154, P2_U5155, P2_U5156);
  and ginst13370 (P2_U3801, P2_U5159, P2_U5160, P2_U5161);
  and ginst13371 (P2_U3802, P2_U5164, P2_U5165, P2_U5166);
  and ginst13372 (P2_U3803, P2_U4443, P2_U5178, P2_U5179);
  and ginst13373 (P2_U3804, P2_U5186, P2_U5187, P2_U5188);
  and ginst13374 (P2_U3805, P2_U5191, P2_U5192, P2_U5193);
  and ginst13375 (P2_U3806, P2_U5196, P2_U5197, P2_U5198);
  and ginst13376 (P2_U3807, P2_U5201, P2_U5202, P2_U5203);
  and ginst13377 (P2_U3808, P2_U5206, P2_U5207, P2_U5208);
  and ginst13378 (P2_U3809, P2_U5211, P2_U5212, P2_U5213);
  and ginst13379 (P2_U3810, P2_U5216, P2_U5217, P2_U5218);
  and ginst13380 (P2_U3811, P2_U5221, P2_U5222, P2_U5223);
  and ginst13381 (P2_U3812, P2_U4443, P2_U5236, P2_U5237);
  and ginst13382 (P2_U3813, P2_U5244, P2_U5245, P2_U5246);
  and ginst13383 (P2_U3814, P2_U5249, P2_U5250, P2_U5251);
  and ginst13384 (P2_U3815, P2_U5254, P2_U5255, P2_U5256);
  and ginst13385 (P2_U3816, P2_U5259, P2_U5260, P2_U5261);
  and ginst13386 (P2_U3817, P2_U5264, P2_U5265, P2_U5266);
  and ginst13387 (P2_U3818, P2_U5269, P2_U5270, P2_U5271);
  and ginst13388 (P2_U3819, P2_U5274, P2_U5275, P2_U5276);
  and ginst13389 (P2_U3820, P2_U5279, P2_U5280, P2_U5281);
  and ginst13390 (P2_U3821, P2_U4443, P2_U5293, P2_U5294);
  and ginst13391 (P2_U3822, P2_U5301, P2_U5302, P2_U5303);
  and ginst13392 (P2_U3823, P2_U5306, P2_U5307, P2_U5308);
  and ginst13393 (P2_U3824, P2_U5311, P2_U5312, P2_U5313);
  and ginst13394 (P2_U3825, P2_U5316, P2_U5317, P2_U5318);
  and ginst13395 (P2_U3826, P2_U5321, P2_U5322, P2_U5323);
  and ginst13396 (P2_U3827, P2_U5326, P2_U5327, P2_U5328);
  and ginst13397 (P2_U3828, P2_U5331, P2_U5332, P2_U5333);
  and ginst13398 (P2_U3829, P2_U5336, P2_U5337, P2_U5338);
  and ginst13399 (P2_U3830, P2_U4443, P2_U5351, P2_U5352);
  and ginst13400 (P2_U3831, P2_U5359, P2_U5360, P2_U5361);
  and ginst13401 (P2_U3832, P2_U5364, P2_U5365, P2_U5366);
  and ginst13402 (P2_U3833, P2_U5369, P2_U5370, P2_U5371);
  and ginst13403 (P2_U3834, P2_U5374, P2_U5375, P2_U5376);
  and ginst13404 (P2_U3835, P2_U5379, P2_U5380, P2_U5381);
  and ginst13405 (P2_U3836, P2_U5384, P2_U5385, P2_U5386);
  and ginst13406 (P2_U3837, P2_U5389, P2_U5390, P2_U5391);
  and ginst13407 (P2_U3838, P2_U5394, P2_U5395, P2_U5396);
  and ginst13408 (P2_U3839, P2_U4443, P2_U5408, P2_U5409);
  and ginst13409 (P2_U3840, P2_U5416, P2_U5417, P2_U5418);
  and ginst13410 (P2_U3841, P2_U5421, P2_U5422, P2_U5423);
  and ginst13411 (P2_U3842, P2_U5426, P2_U5427, P2_U5428);
  and ginst13412 (P2_U3843, P2_U5431, P2_U5432, P2_U5433);
  and ginst13413 (P2_U3844, P2_U5436, P2_U5437, P2_U5438);
  and ginst13414 (P2_U3845, P2_U5441, P2_U5442, P2_U5443);
  and ginst13415 (P2_U3846, P2_U5446, P2_U5447, P2_U5448);
  and ginst13416 (P2_U3847, P2_U5451, P2_U5452, P2_U5453);
  and ginst13417 (P2_U3848, P2_U4443, P2_U5466, P2_U5467);
  and ginst13418 (P2_U3849, P2_U5474, P2_U5475, P2_U5476);
  and ginst13419 (P2_U3850, P2_U5479, P2_U5480, P2_U5481);
  and ginst13420 (P2_U3851, P2_U5484, P2_U5485, P2_U5486);
  and ginst13421 (P2_U3852, P2_U5489, P2_U5490, P2_U5491);
  and ginst13422 (P2_U3853, P2_U5494, P2_U5495, P2_U5496);
  and ginst13423 (P2_U3854, P2_U5499, P2_U5500, P2_U5501);
  and ginst13424 (P2_U3855, P2_U5504, P2_U5505, P2_U5506);
  and ginst13425 (P2_U3856, P2_U5509, P2_U5510, P2_U5511);
  and ginst13426 (P2_U3857, P2_U4443, P2_U5523, P2_U5524);
  and ginst13427 (P2_U3858, P2_U5531, P2_U5532, P2_U5533);
  and ginst13428 (P2_U3859, P2_U5536, P2_U5537, P2_U5538);
  and ginst13429 (P2_U3860, P2_U5541, P2_U5542, P2_U5543);
  and ginst13430 (P2_U3861, P2_U5546, P2_U5547, P2_U5548);
  and ginst13431 (P2_U3862, P2_U5551, P2_U5552, P2_U5553);
  and ginst13432 (P2_U3863, P2_U5556, P2_U5557, P2_U5558);
  and ginst13433 (P2_U3864, P2_U5561, P2_U5562, P2_U5563);
  and ginst13434 (P2_U3865, P2_U5566, P2_U5567, P2_U5568);
  and ginst13435 (P2_U3866, P2_R2147_U7, P2_U4466);
  and ginst13436 (P2_U3867, P2_STATE2_REG_0__SCAN_IN, P2_FLUSH_REG_SCAN_IN);
  and ginst13437 (P2_U3868, P2_U5571, P2_U5573);
  and ginst13438 (P2_U3869, P2_U3868, P2_U5576);
  and ginst13439 (P2_U3870, P2_U4456, P2_U4460);
  and ginst13440 (P2_U3871, P2_U2512, P2_U3870, P2_U8070, P2_U8071);
  and ginst13441 (P2_U3872, P2_U4455, P2_U5583);
  and ginst13442 (P2_U3873, P2_U3521, P2_U7869);
  and ginst13443 (P2_U3874, P2_U3278, P2_U7861);
  and ginst13444 (P2_U3875, P2_U3874, P2_U4429);
  and ginst13445 (P2_U3876, P2_U3279, P2_U4429);
  and ginst13446 (P2_U3877, P2_U5593, P2_U7859);
  and ginst13447 (P2_U3878, P2_U3521, P2_U7863);
  and ginst13448 (P2_U3879, P2_U3281, P2_U5587, P2_U5588);
  and ginst13449 (P2_U3880, P2_U3254, P2_U5599);
  and ginst13450 (P2_U3881, P2_U3880, P2_U5600, P2_U5601);
  and ginst13451 (P2_U3882, P2_U5602, P2_U7897);
  and ginst13452 (P2_U3883, P2_U5607, P2_U5608);
  and ginst13453 (P2_U3884, P2_U3883, P2_U5609);
  and ginst13454 (P2_U3885, P2_U4396, P2_U5617);
  and ginst13455 (P2_U3886, P2_U2449, P2_U4601);
  and ginst13456 (P2_U3887, P2_U3582, P2_U7859);
  and ginst13457 (P2_U3888, P2_U5626, P2_U5627);
  and ginst13458 (P2_U3889, P2_U3272, P2_U7859);
  and ginst13459 (P2_U3890, P2_U5634, P2_U5635);
  and ginst13460 (P2_U3891, P2_U5649, P2_U5650);
  and ginst13461 (P2_U3892, P2_U5653, P2_U5654);
  and ginst13462 (P2_U3893, P2_U5658, P2_U5659);
  and ginst13463 (P2_U3894, P2_U4456, P2_U4460, P2_U5668);
  and ginst13464 (P2_U3895, P2_U3578, P2_U5674);
  and ginst13465 (P2_U3896, P2_U5680, P2_U5681);
  and ginst13466 (P2_U3897, P2_U5682, P2_U5683);
  and ginst13467 (P2_U3898, P2_U5686, P2_U5687);
  and ginst13468 (P2_U3899, P2_U5688, P2_U5689);
  and ginst13469 (P2_U3900, P2_U5690, P2_U5691);
  and ginst13470 (P2_U3901, P2_U5694, P2_U5695);
  and ginst13471 (P2_U3902, P2_U5696, P2_U5697);
  and ginst13472 (P2_U3903, P2_U5698, P2_U5699);
  and ginst13473 (P2_U3904, P2_U5702, P2_U5703);
  and ginst13474 (P2_U3905, P2_U5704, P2_U5705);
  and ginst13475 (P2_U3906, P2_U5706, P2_U5707);
  and ginst13476 (P2_U3907, P2_U5710, P2_U5711);
  and ginst13477 (P2_U3908, P2_U5712, P2_U5713);
  and ginst13478 (P2_U3909, P2_U5714, P2_U5715);
  and ginst13479 (P2_U3910, P2_U5718, P2_U5719);
  and ginst13480 (P2_U3911, P2_U5720, P2_U5721);
  and ginst13481 (P2_U3912, P2_U5722, P2_U5723);
  and ginst13482 (P2_U3913, P2_U5726, P2_U5727);
  and ginst13483 (P2_U3914, P2_U5728, P2_U5729);
  and ginst13484 (P2_U3915, P2_U5730, P2_U5731);
  and ginst13485 (P2_U3916, P2_U5734, P2_U5735);
  and ginst13486 (P2_U3917, P2_U5736, P2_U5737);
  and ginst13487 (P2_U3918, P2_U5738, P2_U5739);
  and ginst13488 (P2_U3919, P2_U5742, P2_U5743);
  and ginst13489 (P2_U3920, P2_U5744, P2_U5745);
  and ginst13490 (P2_U3921, P2_U5746, P2_U5747);
  and ginst13491 (P2_U3922, P2_U5750, P2_U5751);
  and ginst13492 (P2_U3923, P2_U5752, P2_U5753);
  and ginst13493 (P2_U3924, P2_U5754, P2_U5755);
  and ginst13494 (P2_U3925, P2_U5758, P2_U5759);
  and ginst13495 (P2_U3926, P2_U5760, P2_U5761);
  and ginst13496 (P2_U3927, P2_U5762, P2_U5763);
  and ginst13497 (P2_U3928, P2_U5766, P2_U5767);
  and ginst13498 (P2_U3929, P2_U5768, P2_U5769);
  and ginst13499 (P2_U3930, P2_U5770, P2_U5771);
  and ginst13500 (P2_U3931, P2_U5774, P2_U5775);
  and ginst13501 (P2_U3932, P2_U5776, P2_U5777);
  and ginst13502 (P2_U3933, P2_U5778, P2_U5779);
  and ginst13503 (P2_U3934, P2_U5782, P2_U5783);
  and ginst13504 (P2_U3935, P2_U5784, P2_U5785);
  and ginst13505 (P2_U3936, P2_U5786, P2_U5787);
  and ginst13506 (P2_U3937, P2_U5790, P2_U5791);
  and ginst13507 (P2_U3938, P2_U5792, P2_U5793);
  and ginst13508 (P2_U3939, P2_U5794, P2_U5795);
  and ginst13509 (P2_U3940, P2_U5798, P2_U5799);
  and ginst13510 (P2_U3941, P2_U5800, P2_U5801);
  and ginst13511 (P2_U3942, P2_U5802, P2_U5803);
  and ginst13512 (P2_U3943, P2_U5806, P2_U5807);
  and ginst13513 (P2_U3944, P2_U5808, P2_U5809);
  and ginst13514 (P2_U3945, P2_U5810, P2_U5811);
  and ginst13515 (P2_U3946, P2_U5814, P2_U5815);
  and ginst13516 (P2_U3947, P2_U5816, P2_U5817);
  and ginst13517 (P2_U3948, P2_U5818, P2_U5819);
  and ginst13518 (P2_U3949, P2_U5822, P2_U5823);
  and ginst13519 (P2_U3950, P2_U5824, P2_U5825);
  and ginst13520 (P2_U3951, P2_U5826, P2_U5827);
  and ginst13521 (P2_U3952, P2_U5830, P2_U5831);
  and ginst13522 (P2_U3953, P2_U5832, P2_U5833);
  and ginst13523 (P2_U3954, P2_U5834, P2_U5835);
  and ginst13524 (P2_U3955, P2_U5838, P2_U5839);
  and ginst13525 (P2_U3956, P2_U5840, P2_U5841);
  and ginst13526 (P2_U3957, P2_U5842, P2_U5843);
  and ginst13527 (P2_U3958, P2_U5846, P2_U5847);
  and ginst13528 (P2_U3959, P2_U5848, P2_U5849);
  and ginst13529 (P2_U3960, P2_U5850, P2_U5851);
  and ginst13530 (P2_U3961, P2_U5854, P2_U5855);
  and ginst13531 (P2_U3962, P2_U5856, P2_U5857);
  and ginst13532 (P2_U3963, P2_U5858, P2_U5859);
  and ginst13533 (P2_U3964, P2_U5862, P2_U5863);
  and ginst13534 (P2_U3965, P2_U5864, P2_U5865);
  and ginst13535 (P2_U3966, P2_U5866, P2_U5867);
  and ginst13536 (P2_U3967, P2_U5870, P2_U5871);
  and ginst13537 (P2_U3968, P2_U5872, P2_U5873);
  and ginst13538 (P2_U3969, P2_U5874, P2_U5875);
  and ginst13539 (P2_U3970, P2_U5878, P2_U5879);
  and ginst13540 (P2_U3971, P2_U5880, P2_U5881);
  and ginst13541 (P2_U3972, P2_U5882, P2_U5883);
  and ginst13542 (P2_U3973, P2_U5886, P2_U5887);
  and ginst13543 (P2_U3974, P2_U5888, P2_U5889);
  and ginst13544 (P2_U3975, P2_U5890, P2_U5891);
  and ginst13545 (P2_U3976, P2_U5894, P2_U5895);
  and ginst13546 (P2_U3977, P2_U5896, P2_U5897);
  and ginst13547 (P2_U3978, P2_U5898, P2_U5899);
  and ginst13548 (P2_U3979, P2_U5902, P2_U5903);
  and ginst13549 (P2_U3980, P2_U5904, P2_U5905);
  and ginst13550 (P2_U3981, P2_U5906, P2_U5907);
  and ginst13551 (P2_U3982, P2_U5910, P2_U5911);
  and ginst13552 (P2_U3983, P2_U5912, P2_U5913, P2_U5914, P2_U5915);
  and ginst13553 (P2_U3984, P2_U5918, P2_U5919);
  and ginst13554 (P2_U3985, P2_U5921, P2_U5922, P2_U5923);
  and ginst13555 (P2_U3986, P2_U5926, P2_U5927);
  and ginst13556 (P2_U3987, P2_U5929, P2_U5930, P2_U5931);
  and ginst13557 (P2_U3988, P2_U5934, P2_U5935);
  and ginst13558 (P2_U3989, P2_STATE2_REG_1__SCAN_IN, P2_STATEBS16_REG_SCAN_IN);
  nor ginst13559 (P2_U3990, P2_STATE2_REG_2__SCAN_IN, P2_STATE2_REG_1__SCAN_IN);
  and ginst13560 (P2_U3991, P2_U5941, P2_U5942, P2_U5943);
  and ginst13561 (P2_U3992, P2_U5944, P2_U5945, P2_U5946);
  and ginst13562 (P2_U3993, P2_U5947, P2_U5948, P2_U5949);
  and ginst13563 (P2_U3994, P2_U5950, P2_U5951, P2_U5952);
  and ginst13564 (P2_U3995, P2_U5953, P2_U5954, P2_U5955);
  and ginst13565 (P2_U3996, P2_U5956, P2_U5957, P2_U5958);
  and ginst13566 (P2_U3997, P2_U5959, P2_U5960, P2_U5961);
  and ginst13567 (P2_U3998, P2_U5962, P2_U5963, P2_U5964);
  and ginst13568 (P2_U3999, P2_U5965, P2_U5966, P2_U5967);
  and ginst13569 (P2_U4000, P2_U5968, P2_U5969, P2_U5970);
  and ginst13570 (P2_U4001, P2_U5971, P2_U5972, P2_U5973);
  and ginst13571 (P2_U4002, P2_U5974, P2_U5975, P2_U5976);
  and ginst13572 (P2_U4003, P2_U5977, P2_U5978, P2_U5979);
  and ginst13573 (P2_U4004, P2_U5980, P2_U5981, P2_U5982);
  and ginst13574 (P2_U4005, P2_U5983, P2_U5984, P2_U5985);
  and ginst13575 (P2_U4006, P2_U5986, P2_U5987, P2_U5988);
  and ginst13576 (P2_U4007, P2_U5989, P2_U5990, P2_U5991);
  and ginst13577 (P2_U4008, P2_U5992, P2_U5993, P2_U5994);
  and ginst13578 (P2_U4009, P2_U5995, P2_U5996, P2_U5997);
  and ginst13579 (P2_U4010, P2_U5998, P2_U5999, P2_U6000);
  and ginst13580 (P2_U4011, P2_U6001, P2_U6002, P2_U6003);
  and ginst13581 (P2_U4012, P2_U6004, P2_U6005, P2_U6006);
  and ginst13582 (P2_U4013, P2_U6007, P2_U6008, P2_U6009);
  and ginst13583 (P2_U4014, P2_U6010, P2_U6011, P2_U6012);
  and ginst13584 (P2_U4015, P2_U6013, P2_U6014, P2_U6015);
  and ginst13585 (P2_U4016, P2_U6016, P2_U6017, P2_U6018);
  and ginst13586 (P2_U4017, P2_U6019, P2_U6020, P2_U6021);
  and ginst13587 (P2_U4018, P2_U6022, P2_U6023, P2_U6024);
  and ginst13588 (P2_U4019, P2_U6025, P2_U6026, P2_U6027);
  and ginst13589 (P2_U4020, P2_U6028, P2_U6029, P2_U6030);
  and ginst13590 (P2_U4021, P2_U6031, P2_U6032, P2_U6033);
  and ginst13591 (P2_U4022, P2_U6034, P2_U6035, P2_U6036);
  and ginst13592 (P2_U4023, P2_U6037, P2_U6038, P2_U6039);
  and ginst13593 (P2_U4024, P2_U6040, P2_U6041, P2_U6042);
  and ginst13594 (P2_U4025, P2_U6043, P2_U6044, P2_U6045);
  and ginst13595 (P2_U4026, P2_U6046, P2_U6047, P2_U6048);
  and ginst13596 (P2_U4027, P2_U6049, P2_U6050, P2_U6051);
  and ginst13597 (P2_U4028, P2_U6052, P2_U6053, P2_U6054);
  and ginst13598 (P2_U4029, P2_U6055, P2_U6056, P2_U6057);
  and ginst13599 (P2_U4030, P2_U6058, P2_U6059, P2_U6060);
  and ginst13600 (P2_U4031, P2_U6061, P2_U6062, P2_U6063);
  and ginst13601 (P2_U4032, P2_U6064, P2_U6065, P2_U6066);
  and ginst13602 (P2_U4033, P2_U6067, P2_U6068, P2_U6069);
  and ginst13603 (P2_U4034, P2_U6070, P2_U6071, P2_U6072);
  and ginst13604 (P2_U4035, P2_U6073, P2_U6074, P2_U6075);
  and ginst13605 (P2_U4036, P2_U6076, P2_U6077, P2_U6078);
  and ginst13606 (P2_U4037, P2_U6079, P2_U6080, P2_U6081);
  and ginst13607 (P2_U4038, P2_U6082, P2_U6083, P2_U6084);
  and ginst13608 (P2_U4039, P2_U6085, P2_U6086, P2_U6087);
  and ginst13609 (P2_U4040, P2_U6088, P2_U6089, P2_U6090);
  and ginst13610 (P2_U4041, P2_U6091, P2_U6092, P2_U6093);
  and ginst13611 (P2_U4042, P2_U6094, P2_U6095, P2_U6096);
  and ginst13612 (P2_U4043, P2_U6097, P2_U6098, P2_U6099);
  and ginst13613 (P2_U4044, P2_U6100, P2_U6101, P2_U6102);
  and ginst13614 (P2_U4045, P2_U6103, P2_U6104, P2_U6105);
  and ginst13615 (P2_U4046, P2_U6106, P2_U6107, P2_U6108);
  and ginst13616 (P2_U4047, P2_U6109, P2_U6110, P2_U6111);
  and ginst13617 (P2_U4048, P2_U6112, P2_U6113, P2_U6114);
  and ginst13618 (P2_U4049, P2_U6115, P2_U6116, P2_U6117);
  and ginst13619 (P2_U4050, P2_U6118, P2_U6119, P2_U6120);
  and ginst13620 (P2_U4051, P2_U6121, P2_U6122, P2_U6123);
  and ginst13621 (P2_U4052, P2_U6124, P2_U6125, P2_U6126);
  and ginst13622 (P2_U4053, P2_U6127, P2_U6128, P2_U6129);
  and ginst13623 (P2_U4054, P2_U6130, P2_U6131, P2_U6132);
  and ginst13624 (P2_U4055, P2_U2356, P2_U4468, P2_U6133);
  and ginst13625 (P2_U4056, P2_STATE2_REG_0__SCAN_IN, P2_U3280, P2_U7871);
  and ginst13626 (P2_U4057, P2_U2616, P2_U4468);
  and ginst13627 (P2_U4058, P2_U2374, P2_U4417);
  and ginst13628 (P2_U4059, P2_U6329, P2_U6330);
  and ginst13629 (P2_U4060, P2_U6333, P2_U6334);
  and ginst13630 (P2_U4061, P2_U6337, P2_U6338);
  and ginst13631 (P2_U4062, P2_U6341, P2_U6342);
  and ginst13632 (P2_U4063, P2_U6345, P2_U6346);
  and ginst13633 (P2_U4064, P2_U6349, P2_U6350);
  and ginst13634 (P2_U4065, P2_U6353, P2_U6354);
  and ginst13635 (P2_U4066, P2_U6357, P2_U6358);
  and ginst13636 (P2_U4067, P2_U6361, P2_U6362);
  and ginst13637 (P2_U4068, P2_U6365, P2_U6366);
  and ginst13638 (P2_U4069, P2_U4453, P2_U4454, P2_U6569);
  and ginst13639 (P2_U4070, P2_U4071, P2_U6573, P2_U6574);
  and ginst13640 (P2_U4071, P2_U6576, P2_U6577);
  and ginst13641 (P2_U4072, P2_U4073, P2_U6578);
  and ginst13642 (P2_U4073, P2_U6580, P2_U6581);
  and ginst13643 (P2_U4074, P2_U4075, P2_U6582, P2_U6583);
  and ginst13644 (P2_U4075, P2_U6585, P2_U6586);
  and ginst13645 (P2_U4076, P2_U4077, P2_U6587);
  and ginst13646 (P2_U4077, P2_U6589, P2_U6590);
  and ginst13647 (P2_U4078, P2_U4079, P2_U6591, P2_U6592);
  and ginst13648 (P2_U4079, P2_U6594, P2_U6595);
  and ginst13649 (P2_U4080, P2_U4081, P2_U6596);
  and ginst13650 (P2_U4081, P2_U6598, P2_U6599);
  and ginst13651 (P2_U4082, P2_U4083, P2_U6600, P2_U6601);
  and ginst13652 (P2_U4083, P2_U6603, P2_U6604);
  and ginst13653 (P2_U4084, P2_U4085, P2_U6605);
  and ginst13654 (P2_U4085, P2_U6607, P2_U6608);
  and ginst13655 (P2_U4086, P2_U4446, P2_U6609, P2_U6610);
  and ginst13656 (P2_U4087, P2_U4088, P2_U6615);
  and ginst13657 (P2_U4088, P2_U6616, P2_U6617);
  and ginst13658 (P2_U4089, P2_U4086, P2_U6611, P2_U6612, P2_U6613, P2_U6614);
  and ginst13659 (P2_U4090, P2_U4446, P2_U6618, P2_U6619);
  and ginst13660 (P2_U4091, P2_U4092, P2_U6624);
  and ginst13661 (P2_U4092, P2_U6625, P2_U6626);
  and ginst13662 (P2_U4093, P2_U4090, P2_U6620, P2_U6621, P2_U6622, P2_U6623);
  and ginst13663 (P2_U4094, P2_U4446, P2_U6627, P2_U6628);
  and ginst13664 (P2_U4095, P2_U4096, P2_U6631);
  and ginst13665 (P2_U4096, P2_U6633, P2_U6634);
  and ginst13666 (P2_U4097, P2_U4446, P2_U6635, P2_U6636);
  and ginst13667 (P2_U4098, P2_U4099, P2_U6639);
  and ginst13668 (P2_U4099, P2_U6641, P2_U6642);
  and ginst13669 (P2_U4100, P2_U4446, P2_U6643, P2_U6644);
  and ginst13670 (P2_U4101, P2_U4102, P2_U6647);
  and ginst13671 (P2_U4102, P2_U6649, P2_U6650);
  and ginst13672 (P2_U4103, P2_U4446, P2_U6651, P2_U6652);
  and ginst13673 (P2_U4104, P2_U4105, P2_U6655);
  and ginst13674 (P2_U4105, P2_U6657, P2_U6658);
  and ginst13675 (P2_U4106, P2_U4446, P2_U6659, P2_U6660);
  and ginst13676 (P2_U4107, P2_U4108, P2_U6663);
  and ginst13677 (P2_U4108, P2_U6665, P2_U6666);
  and ginst13678 (P2_U4109, P2_U4446, P2_U6667, P2_U6668);
  and ginst13679 (P2_U4110, P2_U4111, P2_U6671);
  and ginst13680 (P2_U4111, P2_U6673, P2_U6674);
  and ginst13681 (P2_U4112, P2_U4446, P2_U6675, P2_U6678);
  and ginst13682 (P2_U4113, P2_U4114, P2_U6679);
  and ginst13683 (P2_U4114, P2_U6681, P2_U6682);
  and ginst13684 (P2_U4115, P2_U4446, P2_U6683, P2_U6686);
  and ginst13685 (P2_U4116, P2_U4117, P2_U6687);
  and ginst13686 (P2_U4117, P2_U6689, P2_U6690);
  and ginst13687 (P2_U4118, P2_U4446, P2_U6691, P2_U6694);
  and ginst13688 (P2_U4119, P2_U4120, P2_U6695);
  and ginst13689 (P2_U4120, P2_U6697, P2_U6698);
  and ginst13690 (P2_U4121, P2_U4446, P2_U6699);
  and ginst13691 (P2_U4122, P2_U4123, P2_U6703);
  and ginst13692 (P2_U4123, P2_U6705, P2_U6706);
  and ginst13693 (P2_U4124, P2_U4121, P2_U6700, P2_U6701, P2_U6702, P2_U6704);
  and ginst13694 (P2_U4125, P2_U4446, P2_U6707);
  and ginst13695 (P2_U4126, P2_U4127, P2_U6711);
  and ginst13696 (P2_U4127, P2_U6713, P2_U6714);
  and ginst13697 (P2_U4128, P2_U4125, P2_U6708, P2_U6709, P2_U6710, P2_U6712);
  and ginst13698 (P2_U4129, P2_U4446, P2_U6715);
  and ginst13699 (P2_U4130, P2_U4131, P2_U6719);
  and ginst13700 (P2_U4131, P2_U6721, P2_U6722);
  and ginst13701 (P2_U4132, P2_U4129, P2_U6716, P2_U6717, P2_U6718, P2_U6720);
  and ginst13702 (P2_U4133, P2_U4446, P2_U6723);
  and ginst13703 (P2_U4134, P2_U4135, P2_U6727);
  and ginst13704 (P2_U4135, P2_U6729, P2_U6730);
  and ginst13705 (P2_U4136, P2_U4133, P2_U6724, P2_U6725, P2_U6726, P2_U6728);
  and ginst13706 (P2_U4137, P2_U4446, P2_U6731);
  and ginst13707 (P2_U4138, P2_U4139, P2_U6735);
  and ginst13708 (P2_U4139, P2_U6737, P2_U6738);
  and ginst13709 (P2_U4140, P2_U4137, P2_U6732, P2_U6733, P2_U6734, P2_U6736);
  and ginst13710 (P2_U4141, P2_U4142, P2_U6743);
  and ginst13711 (P2_U4142, P2_U6745, P2_U6746);
  and ginst13712 (P2_U4143, P2_U6739, P2_U6740, P2_U6741, P2_U6742, P2_U6744);
  and ginst13713 (P2_U4144, P2_U4145, P2_U6751);
  and ginst13714 (P2_U4145, P2_U6753, P2_U6754);
  and ginst13715 (P2_U4146, P2_U6747, P2_U6748, P2_U6749, P2_U6750, P2_U6752);
  and ginst13716 (P2_U4147, P2_U6761, P2_U6762);
  and ginst13717 (P2_U4148, P2_U4147, P2_U6759, P2_U6760);
  and ginst13718 (P2_U4149, P2_U4150, P2_U6763, P2_U6765, P2_U6766, P2_U6768);
  and ginst13719 (P2_U4150, P2_U4151, P2_U6767);
  and ginst13720 (P2_U4151, P2_U6769, P2_U6770);
  and ginst13721 (P2_U4152, P2_U4153, P2_U6771, P2_U6773, P2_U6774, P2_U6776);
  and ginst13722 (P2_U4153, P2_U4154, P2_U6775);
  and ginst13723 (P2_U4154, P2_U6777, P2_U6778);
  and ginst13724 (P2_U4155, P2_U6785, P2_U6786);
  and ginst13725 (P2_U4156, P2_U4155, P2_U6783, P2_U6784);
  and ginst13726 (P2_U4157, P2_U6793, P2_U6794);
  and ginst13727 (P2_U4158, P2_U4157, P2_U6791, P2_U6792);
  and ginst13728 (P2_U4159, P2_U6801, P2_U6802);
  and ginst13729 (P2_U4160, P2_U4159, P2_U6799, P2_U6800);
  and ginst13730 (P2_U4161, P2_U6809, P2_U6810);
  and ginst13731 (P2_U4162, P2_U4161, P2_U6807, P2_U6808);
  and ginst13732 (P2_U4163, P2_U6817, P2_U6818);
  and ginst13733 (P2_U4164, P2_U4163, P2_U6815, P2_U6816);
  and ginst13734 (P2_U4165, P2_U6825, P2_U6826);
  and ginst13735 (P2_U4166, P2_U4165, P2_U6823, P2_U6824);
  and ginst13736 (P2_U4167, P2_U6833, P2_U6834);
  and ginst13737 (P2_U4168, P2_U4167, P2_U6831, P2_U6832);
  nor ginst13738 (P2_U4169, P2_DATAWIDTH_REG_2__SCAN_IN, P2_DATAWIDTH_REG_3__SCAN_IN, P2_DATAWIDTH_REG_4__SCAN_IN, P2_DATAWIDTH_REG_5__SCAN_IN);
  nor ginst13739 (P2_U4170, P2_DATAWIDTH_REG_6__SCAN_IN, P2_DATAWIDTH_REG_7__SCAN_IN, P2_DATAWIDTH_REG_8__SCAN_IN, P2_DATAWIDTH_REG_9__SCAN_IN);
  and ginst13740 (P2_U4171, P2_U4169, P2_U4170);
  nor ginst13741 (P2_U4172, P2_DATAWIDTH_REG_10__SCAN_IN, P2_DATAWIDTH_REG_11__SCAN_IN, P2_DATAWIDTH_REG_12__SCAN_IN, P2_DATAWIDTH_REG_13__SCAN_IN);
  nor ginst13742 (P2_U4173, P2_DATAWIDTH_REG_14__SCAN_IN, P2_DATAWIDTH_REG_15__SCAN_IN, P2_DATAWIDTH_REG_16__SCAN_IN, P2_DATAWIDTH_REG_17__SCAN_IN);
  and ginst13743 (P2_U4174, P2_U4172, P2_U4173);
  nor ginst13744 (P2_U4175, P2_DATAWIDTH_REG_18__SCAN_IN, P2_DATAWIDTH_REG_19__SCAN_IN, P2_DATAWIDTH_REG_20__SCAN_IN, P2_DATAWIDTH_REG_21__SCAN_IN);
  nor ginst13745 (P2_U4176, P2_DATAWIDTH_REG_22__SCAN_IN, P2_DATAWIDTH_REG_23__SCAN_IN, P2_DATAWIDTH_REG_24__SCAN_IN, P2_DATAWIDTH_REG_25__SCAN_IN);
  and ginst13746 (P2_U4177, P2_U4175, P2_U4176);
  nor ginst13747 (P2_U4178, P2_DATAWIDTH_REG_26__SCAN_IN, P2_DATAWIDTH_REG_27__SCAN_IN);
  nor ginst13748 (P2_U4179, P2_DATAWIDTH_REG_28__SCAN_IN, P2_DATAWIDTH_REG_29__SCAN_IN);
  nor ginst13749 (P2_U4180, P2_DATAWIDTH_REG_30__SCAN_IN, P2_DATAWIDTH_REG_31__SCAN_IN);
  and ginst13750 (P2_U4181, P2_U4178, P2_U4179, P2_U4180, P2_U6835);
  nor ginst13751 (P2_U4182, P2_DATAWIDTH_REG_0__SCAN_IN, P2_DATAWIDTH_REG_1__SCAN_IN, P2_REIP_REG_0__SCAN_IN);
  nor ginst13752 (P2_U4183, P2_DATAWIDTH_REG_1__SCAN_IN, P2_REIP_REG_1__SCAN_IN);
  and ginst13753 (P2_U4184, P2_U6844, P2_U7873);
  and ginst13754 (P2_U4185, P2_U3301, P2_U6848);
  and ginst13755 (P2_U4186, P2_U4185, P2_U6849);
  and ginst13756 (P2_U4187, P2_STATE2_REG_1__SCAN_IN, P2_U3265);
  and ginst13757 (P2_U4188, P2_U3313, P2_U6841, P2_U6842);
  and ginst13758 (P2_U4189, P2_U2374, P2_U3253);
  and ginst13759 (P2_U4190, P2_U3534, P2_U6860);
  and ginst13760 (P2_U4191, P2_U6862, P2_U6863, P2_U6864, P2_U6865);
  and ginst13761 (P2_U4192, P2_U6866, P2_U6867, P2_U6868, P2_U6869);
  and ginst13762 (P2_U4193, P2_U6870, P2_U6871, P2_U6872, P2_U6873);
  and ginst13763 (P2_U4194, P2_U6874, P2_U6875, P2_U6876, P2_U6877);
  and ginst13764 (P2_U4195, P2_U6878, P2_U6879, P2_U6880, P2_U6881);
  and ginst13765 (P2_U4196, P2_U6882, P2_U6883, P2_U6884, P2_U6885);
  and ginst13766 (P2_U4197, P2_U6886, P2_U6887, P2_U6888, P2_U6889);
  and ginst13767 (P2_U4198, P2_U6890, P2_U6891, P2_U6892, P2_U6893);
  and ginst13768 (P2_U4199, P2_U6894, P2_U6895, P2_U6896, P2_U6897);
  and ginst13769 (P2_U4200, P2_U6898, P2_U6899, P2_U6900, P2_U6901);
  and ginst13770 (P2_U4201, P2_U6902, P2_U6903, P2_U6904, P2_U6905);
  and ginst13771 (P2_U4202, P2_U6906, P2_U6907, P2_U6908, P2_U6909);
  and ginst13772 (P2_U4203, P2_U6910, P2_U6911, P2_U6912, P2_U6913);
  and ginst13773 (P2_U4204, P2_U6914, P2_U6915, P2_U6916, P2_U6917);
  and ginst13774 (P2_U4205, P2_U6918, P2_U6919, P2_U6920, P2_U6921);
  and ginst13775 (P2_U4206, P2_U6922, P2_U6923, P2_U6924, P2_U6925);
  and ginst13776 (P2_U4207, P2_U6926, P2_U6927, P2_U6928, P2_U6929);
  and ginst13777 (P2_U4208, P2_U6930, P2_U6931, P2_U6932, P2_U6933);
  and ginst13778 (P2_U4209, P2_U6934, P2_U6935, P2_U6936, P2_U6937);
  and ginst13779 (P2_U4210, P2_U6938, P2_U6939, P2_U6940, P2_U6941);
  and ginst13780 (P2_U4211, P2_U6942, P2_U6943, P2_U6944, P2_U6945);
  and ginst13781 (P2_U4212, P2_U6946, P2_U6947, P2_U6948, P2_U6949);
  and ginst13782 (P2_U4213, P2_U6950, P2_U6951, P2_U6952, P2_U6953);
  and ginst13783 (P2_U4214, P2_U6954, P2_U6955, P2_U6956, P2_U6957);
  and ginst13784 (P2_U4215, P2_U6958, P2_U6959, P2_U6960, P2_U6961);
  and ginst13785 (P2_U4216, P2_U6962, P2_U6963, P2_U6964, P2_U6965);
  and ginst13786 (P2_U4217, P2_U6966, P2_U6967, P2_U6968, P2_U6969);
  and ginst13787 (P2_U4218, P2_U6970, P2_U6971, P2_U6972, P2_U6973);
  and ginst13788 (P2_U4219, P2_U6974, P2_U6975, P2_U6976, P2_U6977);
  and ginst13789 (P2_U4220, P2_U6978, P2_U6979, P2_U6980, P2_U6981);
  and ginst13790 (P2_U4221, P2_U6982, P2_U6983, P2_U6984, P2_U6985);
  and ginst13791 (P2_U4222, P2_U6986, P2_U6987, P2_U6988, P2_U6989);
  and ginst13792 (P2_U4223, P2_U6990, P2_U6991, P2_U6992, P2_U6993);
  and ginst13793 (P2_U4224, P2_U6994, P2_U6995, P2_U6996, P2_U6997);
  and ginst13794 (P2_U4225, P2_U6998, P2_U6999, P2_U7000, P2_U7001);
  and ginst13795 (P2_U4226, P2_U7002, P2_U7003, P2_U7004, P2_U7005);
  and ginst13796 (P2_U4227, P2_U7008, P2_U7009, P2_U7010, P2_U7011);
  and ginst13797 (P2_U4228, P2_U7012, P2_U7013, P2_U7014, P2_U7015);
  and ginst13798 (P2_U4229, P2_U7016, P2_U7017, P2_U7018, P2_U7019);
  and ginst13799 (P2_U4230, P2_U7020, P2_U7021, P2_U7022, P2_U7023);
  and ginst13800 (P2_U4231, P2_U7024, P2_U7025, P2_U7026, P2_U7027);
  and ginst13801 (P2_U4232, P2_U7028, P2_U7029, P2_U7030, P2_U7031);
  and ginst13802 (P2_U4233, P2_U7032, P2_U7033, P2_U7034, P2_U7035);
  and ginst13803 (P2_U4234, P2_U7036, P2_U7037, P2_U7038, P2_U7039);
  and ginst13804 (P2_U4235, P2_U7040, P2_U7041, P2_U7042, P2_U7043);
  and ginst13805 (P2_U4236, P2_U7044, P2_U7045, P2_U7046, P2_U7047);
  and ginst13806 (P2_U4237, P2_U7048, P2_U7049, P2_U7050, P2_U7051);
  and ginst13807 (P2_U4238, P2_U7052, P2_U7053, P2_U7054, P2_U7055);
  and ginst13808 (P2_U4239, P2_U7056, P2_U7057, P2_U7058, P2_U7059);
  and ginst13809 (P2_U4240, P2_U7060, P2_U7061, P2_U7062, P2_U7063);
  and ginst13810 (P2_U4241, P2_U7064, P2_U7065, P2_U7066, P2_U7067);
  and ginst13811 (P2_U4242, P2_U7068, P2_U7069, P2_U7070, P2_U7071);
  and ginst13812 (P2_U4243, P2_U7072, P2_U7073, P2_U7074, P2_U7075);
  and ginst13813 (P2_U4244, P2_U7076, P2_U7077, P2_U7078, P2_U7079);
  and ginst13814 (P2_U4245, P2_U7080, P2_U7081, P2_U7082, P2_U7083);
  and ginst13815 (P2_U4246, P2_U7084, P2_U7085, P2_U7086, P2_U7087);
  and ginst13816 (P2_U4247, P2_U7088, P2_U7089, P2_U7090, P2_U7091);
  and ginst13817 (P2_U4248, P2_U7092, P2_U7093, P2_U7094, P2_U7095);
  and ginst13818 (P2_U4249, P2_U7096, P2_U7097, P2_U7098, P2_U7099);
  and ginst13819 (P2_U4250, P2_U7100, P2_U7101, P2_U7102, P2_U7103);
  and ginst13820 (P2_U4251, P2_U7104, P2_U7105, P2_U7106, P2_U7107);
  and ginst13821 (P2_U4252, P2_U7108, P2_U7109, P2_U7110, P2_U7111);
  and ginst13822 (P2_U4253, P2_U7112, P2_U7113, P2_U7114, P2_U7115);
  and ginst13823 (P2_U4254, P2_U7116, P2_U7117, P2_U7118, P2_U7119);
  and ginst13824 (P2_U4255, P2_U7120, P2_U7121, P2_U7122, P2_U7123);
  and ginst13825 (P2_U4256, P2_U7124, P2_U7125, P2_U7126, P2_U7127);
  and ginst13826 (P2_U4257, P2_U7128, P2_U7129, P2_U7130, P2_U7131);
  and ginst13827 (P2_U4258, P2_U7132, P2_U7133, P2_U7134, P2_U7135);
  and ginst13828 (P2_U4259, P2_U7754, P2_U7770, P2_U7786, P2_U7802);
  and ginst13829 (P2_U4260, P2_U7818, P2_U7834, P2_U7850, P2_U7874);
  and ginst13830 (P2_U4261, P2_U7755, P2_U7771, P2_U7787, P2_U7803);
  and ginst13831 (P2_U4262, P2_U7819, P2_U7835, P2_U7851, P2_U7875);
  and ginst13832 (P2_U4263, P2_U7756, P2_U7772, P2_U7788, P2_U7804);
  and ginst13833 (P2_U4264, P2_U7820, P2_U7836, P2_U7852, P2_U7876);
  and ginst13834 (P2_U4265, P2_U7757, P2_U7773, P2_U7789, P2_U7805);
  and ginst13835 (P2_U4266, P2_U7821, P2_U7837, P2_U7853, P2_U7877);
  and ginst13836 (P2_U4267, P2_U7758, P2_U7774, P2_U7790, P2_U7806);
  and ginst13837 (P2_U4268, P2_U7822, P2_U7838, P2_U7854, P2_U7878);
  and ginst13838 (P2_U4269, P2_U7759, P2_U7775, P2_U7791, P2_U7807);
  and ginst13839 (P2_U4270, P2_U7823, P2_U7839, P2_U7855, P2_U7879);
  and ginst13840 (P2_U4271, P2_U7760, P2_U7776, P2_U7792, P2_U7808);
  and ginst13841 (P2_U4272, P2_U7824, P2_U7840, P2_U7856, P2_U7880);
  and ginst13842 (P2_U4273, P2_U7761, P2_U7777, P2_U7793, P2_U7809);
  and ginst13843 (P2_U4274, P2_U7825, P2_U7841, P2_U7857, P2_U7881);
  and ginst13844 (P2_U4275, P2_U4276, P2_U7861);
  and ginst13845 (P2_U4276, P2_STATE2_REG_2__SCAN_IN, P2_STATE2_REG_0__SCAN_IN, P2_U3300);
  and ginst13846 (P2_U4277, P2_U7167, P2_U7168, P2_U7169, P2_U7170);
  and ginst13847 (P2_U4278, P2_U7171, P2_U7172, P2_U7173, P2_U7174);
  and ginst13848 (P2_U4279, P2_U7175, P2_U7176, P2_U7177, P2_U7178);
  and ginst13849 (P2_U4280, P2_U7179, P2_U7180, P2_U7181, P2_U7182);
  and ginst13850 (P2_U4281, P2_U7184, P2_U7185, P2_U7186, P2_U7187);
  and ginst13851 (P2_U4282, P2_U7188, P2_U7189, P2_U7190, P2_U7191);
  and ginst13852 (P2_U4283, P2_U7192, P2_U7193, P2_U7194, P2_U7195);
  and ginst13853 (P2_U4284, P2_U7196, P2_U7197, P2_U7198, P2_U7199);
  and ginst13854 (P2_U4285, P2_U7201, P2_U7202, P2_U7203, P2_U7204);
  and ginst13855 (P2_U4286, P2_U7205, P2_U7206, P2_U7207, P2_U7208);
  and ginst13856 (P2_U4287, P2_U7209, P2_U7210, P2_U7211, P2_U7212);
  and ginst13857 (P2_U4288, P2_U7213, P2_U7214, P2_U7215, P2_U7216);
  and ginst13858 (P2_U4289, P2_U7218, P2_U7219, P2_U7220, P2_U7221);
  and ginst13859 (P2_U4290, P2_U7222, P2_U7223, P2_U7224, P2_U7225);
  and ginst13860 (P2_U4291, P2_U7226, P2_U7227, P2_U7228, P2_U7229);
  and ginst13861 (P2_U4292, P2_U7230, P2_U7231, P2_U7232, P2_U7233);
  and ginst13862 (P2_U4293, P2_U7235, P2_U7236, P2_U7237, P2_U7238);
  and ginst13863 (P2_U4294, P2_U7239, P2_U7240, P2_U7241, P2_U7242);
  and ginst13864 (P2_U4295, P2_U7243, P2_U7244, P2_U7245, P2_U7246);
  and ginst13865 (P2_U4296, P2_U7247, P2_U7248, P2_U7249, P2_U7250);
  and ginst13866 (P2_U4297, P2_U7252, P2_U7253, P2_U7254, P2_U7255);
  and ginst13867 (P2_U4298, P2_U7256, P2_U7257, P2_U7258, P2_U7259);
  and ginst13868 (P2_U4299, P2_U7260, P2_U7261, P2_U7262, P2_U7263);
  and ginst13869 (P2_U4300, P2_U7264, P2_U7265, P2_U7266, P2_U7267);
  and ginst13870 (P2_U4301, P2_U7269, P2_U7270, P2_U7271, P2_U7272);
  and ginst13871 (P2_U4302, P2_U7273, P2_U7274, P2_U7275, P2_U7276);
  and ginst13872 (P2_U4303, P2_U7277, P2_U7278, P2_U7279, P2_U7280);
  and ginst13873 (P2_U4304, P2_U7281, P2_U7282, P2_U7283, P2_U7284);
  and ginst13874 (P2_U4305, P2_U7286, P2_U7287, P2_U7288, P2_U7289);
  and ginst13875 (P2_U4306, P2_U7290, P2_U7291, P2_U7292, P2_U7293);
  and ginst13876 (P2_U4307, P2_U7294, P2_U7295, P2_U7296, P2_U7297);
  and ginst13877 (P2_U4308, P2_U7298, P2_U7299, P2_U7300, P2_U7301);
  and ginst13878 (P2_U4309, P2_U7303, P2_U7304, P2_U7305, P2_U7306);
  and ginst13879 (P2_U4310, P2_U7307, P2_U7308, P2_U7309, P2_U7310);
  and ginst13880 (P2_U4311, P2_U7311, P2_U7312, P2_U7313, P2_U7314);
  and ginst13881 (P2_U4312, P2_U7315, P2_U7316, P2_U7317, P2_U7318);
  and ginst13882 (P2_U4313, P2_U7320, P2_U7321, P2_U7322, P2_U7323);
  and ginst13883 (P2_U4314, P2_U7324, P2_U7325, P2_U7326, P2_U7327);
  and ginst13884 (P2_U4315, P2_U7328, P2_U7329, P2_U7330, P2_U7331);
  and ginst13885 (P2_U4316, P2_U7332, P2_U7333, P2_U7334, P2_U7335);
  and ginst13886 (P2_U4317, P2_U7337, P2_U7338, P2_U7339, P2_U7340);
  and ginst13887 (P2_U4318, P2_U7341, P2_U7342, P2_U7343, P2_U7344);
  and ginst13888 (P2_U4319, P2_U7345, P2_U7346, P2_U7347, P2_U7348);
  and ginst13889 (P2_U4320, P2_U7349, P2_U7350, P2_U7351, P2_U7352);
  and ginst13890 (P2_U4321, P2_U7354, P2_U7355, P2_U7356, P2_U7357);
  and ginst13891 (P2_U4322, P2_U7358, P2_U7359, P2_U7360, P2_U7361);
  and ginst13892 (P2_U4323, P2_U7362, P2_U7363, P2_U7364, P2_U7365);
  and ginst13893 (P2_U4324, P2_U7366, P2_U7367, P2_U7368, P2_U7369);
  and ginst13894 (P2_U4325, P2_U7371, P2_U7372, P2_U7373, P2_U7374);
  and ginst13895 (P2_U4326, P2_U7375, P2_U7376, P2_U7377, P2_U7378);
  and ginst13896 (P2_U4327, P2_U7379, P2_U7380, P2_U7381, P2_U7382);
  and ginst13897 (P2_U4328, P2_U7383, P2_U7384, P2_U7385, P2_U7386);
  and ginst13898 (P2_U4329, P2_U7388, P2_U7389, P2_U7390, P2_U7391);
  and ginst13899 (P2_U4330, P2_U7392, P2_U7393, P2_U7394, P2_U7395);
  and ginst13900 (P2_U4331, P2_U7396, P2_U7397, P2_U7398, P2_U7399);
  and ginst13901 (P2_U4332, P2_U7400, P2_U7401, P2_U7402, P2_U7403);
  and ginst13902 (P2_U4333, P2_U7405, P2_U7406, P2_U7407, P2_U7408);
  and ginst13903 (P2_U4334, P2_U7409, P2_U7410, P2_U7411, P2_U7412);
  and ginst13904 (P2_U4335, P2_U7413, P2_U7414, P2_U7415, P2_U7416);
  and ginst13905 (P2_U4336, P2_U7417, P2_U7418, P2_U7419, P2_U7420);
  and ginst13906 (P2_U4337, P2_U2616, P2_U3300);
  and ginst13907 (P2_U4338, P2_U4413, P2_U7425);
  and ginst13908 (P2_U4339, P2_U3300, P2_U4595);
  and ginst13909 (P2_U4340, P2_U4414, P2_U7426, P2_U7428);
  and ginst13910 (P2_U4341, P2_U3571, P2_U7430);
  and ginst13911 (P2_U4342, P2_U4341, P2_U4413);
  and ginst13912 (P2_U4343, P2_U7869, P2_U7873);
  and ginst13913 (P2_U4344, P2_U7435, P2_U7436);
  and ginst13914 (P2_U4345, P2_U7439, P2_U7440);
  and ginst13915 (P2_U4346, P2_U7442, P2_U7443);
  and ginst13916 (P2_U4347, P2_U7445, P2_U7446);
  and ginst13917 (P2_U4348, P2_U7448, P2_U7449);
  and ginst13918 (P2_U4349, P2_U7451, P2_U7452);
  and ginst13919 (P2_U4350, P2_U7454, P2_U7455);
  and ginst13920 (P2_U4351, P2_U7457, P2_U7458);
  and ginst13921 (P2_U4352, P2_U7460, P2_U7461);
  and ginst13922 (P2_U4353, P2_U7463, P2_U7464);
  and ginst13923 (P2_U4354, P2_U7466, P2_U7467);
  and ginst13924 (P2_U4355, P2_U7469, P2_U7470);
  and ginst13925 (P2_U4356, P2_U7472, P2_U7473);
  and ginst13926 (P2_U4357, P2_U7475, P2_U7476);
  and ginst13927 (P2_U4358, P2_U7478, P2_U7479);
  and ginst13928 (P2_U4359, P2_U7481, P2_U7482);
  and ginst13929 (P2_U4360, P2_U7484, P2_U7485);
  and ginst13930 (P2_U4361, P2_U7487, P2_U7488);
  and ginst13931 (P2_U4362, P2_U7490, P2_U7491);
  and ginst13932 (P2_U4363, P2_U7493, P2_U7494);
  and ginst13933 (P2_U4364, P2_U7496, P2_U7497);
  and ginst13934 (P2_U4365, P2_U7499, P2_U7500);
  and ginst13935 (P2_U4366, P2_U7502, P2_U7503);
  and ginst13936 (P2_U4367, P2_U7505, P2_U7506);
  and ginst13937 (P2_U4368, P2_U7509, P2_U7510);
  and ginst13938 (P2_U4369, P2_U7513, P2_U7514);
  and ginst13939 (P2_U4370, P2_U7517, P2_U7518);
  and ginst13940 (P2_U4371, P2_U7521, P2_U7522);
  and ginst13941 (P2_U4372, P2_U7525, P2_U7526);
  and ginst13942 (P2_U4373, P2_U7529, P2_U7530);
  and ginst13943 (P2_U4374, P2_U7532, P2_U7533);
  and ginst13944 (P2_U4375, P2_U7535, P2_U7536);
  and ginst13945 (P2_U4376, P2_U3255, P2_U6845);
  and ginst13946 (P2_U4377, P2_U3255, P2_U7863);
  and ginst13947 (P2_U4378, P2_U2356, P2_U7873);
  and ginst13948 (P2_U4379, P2_U7578, P2_U7579, P2_U7580);
  and ginst13949 (P2_U4380, P2_U3269, P2_U7585);
  and ginst13950 (P2_U4381, P2_U2356, P2_U4595);
  and ginst13951 (P2_U4382, P2_U3539, P2_U3577, P2_U4472, P2_U7586, P2_U7587);
  and ginst13952 (P2_U4383, P2_U4422, P2_U7579);
  and ginst13953 (P2_U4384, P2_U4383, P2_U7578);
  and ginst13954 (P2_U4385, P2_U4458, P2_U7580);
  and ginst13955 (P2_U4386, P2_U7589, P2_U7590);
  and ginst13956 (P2_U4387, P2_STATE2_REG_0__SCAN_IN, P2_U7736);
  and ginst13957 (P2_U4388, P2_U3549, P2_U3573, P2_U4457, P2_U4458);
  and ginst13958 (P2_U4389, P2_U7718, P2_U7719);
  and ginst13959 (P2_U4390, P2_U3536, P2_U7731);
  and ginst13960 (P2_U4391, P2_U3536, P2_U7735);
  and ginst13961 (P2_U4392, P2_U7907, P2_U7908);
  and ginst13962 (P2_U4393, P2_U8054, P2_U8055);
  nand ginst13963 (P2_U4394, P2_U3872, P2_U5582);
  and ginst13964 (P2_U4395, P2_U8078, P2_U8079);
  and ginst13965 (P2_U4396, P2_U8091, P2_U8092);
  and ginst13966 (P2_U4397, P2_U8119, P2_U8120);
  and ginst13967 (P2_U4398, P2_U8125, P2_U8126);
  and ginst13968 (P2_U4399, P2_U8131, P2_U8132);
  nand ginst13969 (P2_U4400, P2_U2374, P2_U3291);
  not ginst13970 (P2_U4401, BS16);
  nand ginst13971 (P2_U4402, P2_U4188, P2_U4462);
  nand ginst13972 (P2_U4403, P2_U3534, P2_U4462);
  and ginst13973 (P2_U4404, P2_U8145, P2_U8146);
  nand ginst13974 (P2_U4405, P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN, P2_U7006);
  nand ginst13975 (P2_U4406, P2_U2513, P2_U3871);
  not ginst13976 (P2_U4407, P2_R2219_U29);
  not ginst13977 (P2_U4408, P2_R2219_U8);
  not ginst13978 (P2_U4409, P2_U3553);
  nand ginst13979 (P2_U4410, HOLD, P2_U3265);
  not ginst13980 (P2_U4411, P2_U3290);
  not ginst13981 (P2_U4412, P2_U3571);
  nand ginst13982 (P2_U4413, P2_U4337, P2_U4601);
  nand ginst13983 (P2_U4414, P2_U2616, P2_U3300, P2_U7869);
  nand ginst13984 (P2_U4415, P2_U2447, P2_U3279);
  not ginst13985 (P2_U4416, P2_U3576);
  not ginst13986 (P2_U4417, P2_U3283);
  not ginst13987 (P2_U4418, P2_U3550);
  not ginst13988 (P2_U4419, P2_U3536);
  not ginst13989 (P2_U4420, P2_U3288);
  not ginst13990 (P2_U4421, P2_U3539);
  nand ginst13991 (P2_U4422, P2_U2376, P2_U2450, P2_U3278);
  not ginst13992 (P2_U4423, P2_U3577);
  not ginst13993 (P2_U4424, P2_U3282);
  not ginst13994 (P2_U4425, P2_U3285);
  not ginst13995 (P2_U4426, P2_U3549);
  not ginst13996 (P2_U4427, P2_U3289);
  not ginst13997 (P2_U4428, P2_U3286);
  not ginst13998 (P2_U4429, P2_U3294);
  not ginst13999 (P2_U4430, P2_U3313);
  not ginst14000 (P2_U4431, P2_U3578);
  not ginst14001 (P2_U4432, P2_U3254);
  not ginst14002 (P2_U4433, P2_U3523);
  not ginst14003 (P2_U4434, P2_U3524);
  not ginst14004 (P2_U4435, P2_U3296);
  not ginst14005 (P2_U4436, P2_U3522);
  nand ginst14006 (P2_U4437, P2_U2376, P2_U3875);
  not ginst14007 (P2_U4438, P2_U3547);
  not ginst14008 (P2_U4439, P2_U3259);
  not ginst14009 (P2_U4440, P2_U3543);
  not ginst14010 (P2_U4441, P2_U3542);
  not ginst14011 (P2_U4442, P2_U3538);
  not ginst14012 (P2_U4443, P2_U3306);
  not ginst14013 (P2_U4444, P2_LT_563_1260_U6);
  nand ginst14014 (P2_U4445, P2_U3302, P2_U4430);
  nand ginst14015 (P2_U4446, P2_U3546, P2_U4461);
  nand ginst14016 (P2_U4447, P2_R2219_U7, P2_U2617);
  nand ginst14017 (P2_U4448, P2_U2367, P2_U3290);
  not ginst14018 (P2_U4449, P2_U3261);
  not ginst14019 (P2_U4450, P2_U3260);
  not ginst14020 (P2_U4451, P2_U3425);
  nand ginst14021 (P2_U4452, P2_U4182, P2_U4438);
  nand ginst14022 (P2_U4453, P2_U3718, P2_U4474);
  nand ginst14023 (P2_U4454, P2_STATE2_REG_1__SCAN_IN, P2_U3270, P2_U3284, P2_U3302);
  nand ginst14024 (P2_U4455, P2_U2448, P2_U3867);
  nand ginst14025 (P2_U4456, P2_U2359, P2_U2446);
  nand ginst14026 (P2_U4457, P2_U2356, P2_U3280);
  nand ginst14027 (P2_U4458, P2_U4378, P2_U7577);
  not ginst14028 (P2_U4459, P2_U3575);
  nand ginst14029 (P2_U4460, P2_U2438, P2_U3295);
  not ginst14030 (P2_U4461, P2_U3534);
  nand ginst14031 (P2_U4462, P2_U2374, P2_U6568);
  nand ginst14032 (P2_U4463, P2_U3266, P2_U4574);
  nand ginst14033 (P2_U4464, P2_U2448, P2_U3292);
  nand ginst14034 (P2_U4465, P2_U4474, U211);
  not ginst14035 (P2_U4466, P2_U3303);
  not ginst14036 (P2_U4467, P2_U3540);
  not ginst14037 (P2_U4468, P2_U3304);
  not ginst14038 (P2_U4469, P2_U3305);
  nand ginst14039 (P2_U4470, P2_U2376, P2_U3876);
  not ginst14040 (P2_U4471, P2_U3573);
  nand ginst14041 (P2_U4472, P2_U2376, P2_U4416, P2_U7871);
  not ginst14042 (P2_U4473, P2_U3262);
  not ginst14043 (P2_U4474, P2_U3301);
  not ginst14044 (P2_U4475, P2_U3293);
  not ginst14045 (P2_U4476, P2_U3281);
  not ginst14046 (P2_U4477, P2_U3548);
  nand ginst14047 (P2_U4478, P2_REIP_REG_31__SCAN_IN, P2_U4450);
  nand ginst14048 (P2_U4479, P2_REIP_REG_30__SCAN_IN, P2_U4449);
  nand ginst14049 (P2_U4480, P2_ADDRESS_REG_29__SCAN_IN, P2_U3259);
  nand ginst14050 (P2_U4481, P2_REIP_REG_30__SCAN_IN, P2_U4450);
  nand ginst14051 (P2_U4482, P2_REIP_REG_29__SCAN_IN, P2_U4449);
  nand ginst14052 (P2_U4483, P2_ADDRESS_REG_28__SCAN_IN, P2_U3259);
  nand ginst14053 (P2_U4484, P2_REIP_REG_29__SCAN_IN, P2_U4450);
  nand ginst14054 (P2_U4485, P2_REIP_REG_28__SCAN_IN, P2_U4449);
  nand ginst14055 (P2_U4486, P2_ADDRESS_REG_27__SCAN_IN, P2_U3259);
  nand ginst14056 (P2_U4487, P2_REIP_REG_28__SCAN_IN, P2_U4450);
  nand ginst14057 (P2_U4488, P2_REIP_REG_27__SCAN_IN, P2_U4449);
  nand ginst14058 (P2_U4489, P2_ADDRESS_REG_26__SCAN_IN, P2_U3259);
  nand ginst14059 (P2_U4490, P2_REIP_REG_27__SCAN_IN, P2_U4450);
  nand ginst14060 (P2_U4491, P2_REIP_REG_26__SCAN_IN, P2_U4449);
  nand ginst14061 (P2_U4492, P2_ADDRESS_REG_25__SCAN_IN, P2_U3259);
  nand ginst14062 (P2_U4493, P2_REIP_REG_26__SCAN_IN, P2_U4450);
  nand ginst14063 (P2_U4494, P2_REIP_REG_25__SCAN_IN, P2_U4449);
  nand ginst14064 (P2_U4495, P2_ADDRESS_REG_24__SCAN_IN, P2_U3259);
  nand ginst14065 (P2_U4496, P2_REIP_REG_25__SCAN_IN, P2_U4450);
  nand ginst14066 (P2_U4497, P2_REIP_REG_24__SCAN_IN, P2_U4449);
  nand ginst14067 (P2_U4498, P2_ADDRESS_REG_23__SCAN_IN, P2_U3259);
  nand ginst14068 (P2_U4499, P2_REIP_REG_24__SCAN_IN, P2_U4450);
  nand ginst14069 (P2_U4500, P2_REIP_REG_23__SCAN_IN, P2_U4449);
  nand ginst14070 (P2_U4501, P2_ADDRESS_REG_22__SCAN_IN, P2_U3259);
  nand ginst14071 (P2_U4502, P2_REIP_REG_23__SCAN_IN, P2_U4450);
  nand ginst14072 (P2_U4503, P2_REIP_REG_22__SCAN_IN, P2_U4449);
  nand ginst14073 (P2_U4504, P2_ADDRESS_REG_21__SCAN_IN, P2_U3259);
  nand ginst14074 (P2_U4505, P2_REIP_REG_22__SCAN_IN, P2_U4450);
  nand ginst14075 (P2_U4506, P2_REIP_REG_21__SCAN_IN, P2_U4449);
  nand ginst14076 (P2_U4507, P2_ADDRESS_REG_20__SCAN_IN, P2_U3259);
  nand ginst14077 (P2_U4508, P2_REIP_REG_21__SCAN_IN, P2_U4450);
  nand ginst14078 (P2_U4509, P2_REIP_REG_20__SCAN_IN, P2_U4449);
  nand ginst14079 (P2_U4510, P2_ADDRESS_REG_19__SCAN_IN, P2_U3259);
  nand ginst14080 (P2_U4511, P2_REIP_REG_20__SCAN_IN, P2_U4450);
  nand ginst14081 (P2_U4512, P2_REIP_REG_19__SCAN_IN, P2_U4449);
  nand ginst14082 (P2_U4513, P2_ADDRESS_REG_18__SCAN_IN, P2_U3259);
  nand ginst14083 (P2_U4514, P2_REIP_REG_19__SCAN_IN, P2_U4450);
  nand ginst14084 (P2_U4515, P2_REIP_REG_18__SCAN_IN, P2_U4449);
  nand ginst14085 (P2_U4516, P2_ADDRESS_REG_17__SCAN_IN, P2_U3259);
  nand ginst14086 (P2_U4517, P2_REIP_REG_18__SCAN_IN, P2_U4450);
  nand ginst14087 (P2_U4518, P2_REIP_REG_17__SCAN_IN, P2_U4449);
  nand ginst14088 (P2_U4519, P2_ADDRESS_REG_16__SCAN_IN, P2_U3259);
  nand ginst14089 (P2_U4520, P2_REIP_REG_17__SCAN_IN, P2_U4450);
  nand ginst14090 (P2_U4521, P2_REIP_REG_16__SCAN_IN, P2_U4449);
  nand ginst14091 (P2_U4522, P2_ADDRESS_REG_15__SCAN_IN, P2_U3259);
  nand ginst14092 (P2_U4523, P2_REIP_REG_16__SCAN_IN, P2_U4450);
  nand ginst14093 (P2_U4524, P2_REIP_REG_15__SCAN_IN, P2_U4449);
  nand ginst14094 (P2_U4525, P2_ADDRESS_REG_14__SCAN_IN, P2_U3259);
  nand ginst14095 (P2_U4526, P2_REIP_REG_15__SCAN_IN, P2_U4450);
  nand ginst14096 (P2_U4527, P2_REIP_REG_14__SCAN_IN, P2_U4449);
  nand ginst14097 (P2_U4528, P2_ADDRESS_REG_13__SCAN_IN, P2_U3259);
  nand ginst14098 (P2_U4529, P2_REIP_REG_14__SCAN_IN, P2_U4450);
  nand ginst14099 (P2_U4530, P2_REIP_REG_13__SCAN_IN, P2_U4449);
  nand ginst14100 (P2_U4531, P2_ADDRESS_REG_12__SCAN_IN, P2_U3259);
  nand ginst14101 (P2_U4532, P2_REIP_REG_13__SCAN_IN, P2_U4450);
  nand ginst14102 (P2_U4533, P2_REIP_REG_12__SCAN_IN, P2_U4449);
  nand ginst14103 (P2_U4534, P2_ADDRESS_REG_11__SCAN_IN, P2_U3259);
  nand ginst14104 (P2_U4535, P2_REIP_REG_12__SCAN_IN, P2_U4450);
  nand ginst14105 (P2_U4536, P2_REIP_REG_11__SCAN_IN, P2_U4449);
  nand ginst14106 (P2_U4537, P2_ADDRESS_REG_10__SCAN_IN, P2_U3259);
  nand ginst14107 (P2_U4538, P2_REIP_REG_11__SCAN_IN, P2_U4450);
  nand ginst14108 (P2_U4539, P2_REIP_REG_10__SCAN_IN, P2_U4449);
  nand ginst14109 (P2_U4540, P2_ADDRESS_REG_9__SCAN_IN, P2_U3259);
  nand ginst14110 (P2_U4541, P2_REIP_REG_10__SCAN_IN, P2_U4450);
  nand ginst14111 (P2_U4542, P2_REIP_REG_9__SCAN_IN, P2_U4449);
  nand ginst14112 (P2_U4543, P2_ADDRESS_REG_8__SCAN_IN, P2_U3259);
  nand ginst14113 (P2_U4544, P2_REIP_REG_9__SCAN_IN, P2_U4450);
  nand ginst14114 (P2_U4545, P2_REIP_REG_8__SCAN_IN, P2_U4449);
  nand ginst14115 (P2_U4546, P2_ADDRESS_REG_7__SCAN_IN, P2_U3259);
  nand ginst14116 (P2_U4547, P2_REIP_REG_8__SCAN_IN, P2_U4450);
  nand ginst14117 (P2_U4548, P2_REIP_REG_7__SCAN_IN, P2_U4449);
  nand ginst14118 (P2_U4549, P2_ADDRESS_REG_6__SCAN_IN, P2_U3259);
  nand ginst14119 (P2_U4550, P2_REIP_REG_7__SCAN_IN, P2_U4450);
  nand ginst14120 (P2_U4551, P2_REIP_REG_6__SCAN_IN, P2_U4449);
  nand ginst14121 (P2_U4552, P2_ADDRESS_REG_5__SCAN_IN, P2_U3259);
  nand ginst14122 (P2_U4553, P2_REIP_REG_6__SCAN_IN, P2_U4450);
  nand ginst14123 (P2_U4554, P2_REIP_REG_5__SCAN_IN, P2_U4449);
  nand ginst14124 (P2_U4555, P2_ADDRESS_REG_4__SCAN_IN, P2_U3259);
  nand ginst14125 (P2_U4556, P2_REIP_REG_5__SCAN_IN, P2_U4450);
  nand ginst14126 (P2_U4557, P2_REIP_REG_4__SCAN_IN, P2_U4449);
  nand ginst14127 (P2_U4558, P2_ADDRESS_REG_3__SCAN_IN, P2_U3259);
  nand ginst14128 (P2_U4559, P2_REIP_REG_4__SCAN_IN, P2_U4450);
  nand ginst14129 (P2_U4560, P2_REIP_REG_3__SCAN_IN, P2_U4449);
  nand ginst14130 (P2_U4561, P2_ADDRESS_REG_2__SCAN_IN, P2_U3259);
  nand ginst14131 (P2_U4562, P2_REIP_REG_3__SCAN_IN, P2_U4450);
  nand ginst14132 (P2_U4563, P2_REIP_REG_2__SCAN_IN, P2_U4449);
  nand ginst14133 (P2_U4564, P2_ADDRESS_REG_1__SCAN_IN, P2_U3259);
  nand ginst14134 (P2_U4565, P2_REIP_REG_2__SCAN_IN, P2_U4450);
  nand ginst14135 (P2_U4566, P2_REIP_REG_1__SCAN_IN, P2_U4449);
  nand ginst14136 (P2_U4567, P2_ADDRESS_REG_0__SCAN_IN, P2_U3259);
  not ginst14137 (P2_U4568, P2_U3267);
  nand ginst14138 (P2_U4569, P2_U3265, P2_U4568);
  nand ginst14139 (P2_U4570, NA, P2_U4473);
  not ginst14140 (P2_U4571, P2_U3268);
  nand ginst14141 (P2_U4572, P2_U3265, P2_U4571);
  nand ginst14142 (P2_U4573, P2_U4392, P2_U7891);
  not ginst14143 (P2_U4574, P2_U3263);
  nand ginst14144 (P2_U4575, HOLD, P2_U3256, P2_U4574);
  nand ginst14145 (P2_U4576, P2_STATE_REG_1__SCAN_IN, P2_U3268, U211);
  nand ginst14146 (P2_U4577, P2_U4575, P2_U4576);
  nand ginst14147 (P2_U4578, P2_STATE_REG_0__SCAN_IN, P2_U4570, P2_U4577);
  nand ginst14148 (P2_U4579, P2_STATE_REG_2__SCAN_IN, P2_U4573);
  nand ginst14149 (P2_U4580, P2_STATE_REG_0__SCAN_IN, P2_U4410);
  nand ginst14150 (P2_U4581, P2_STATE_REG_2__SCAN_IN, P2_U4580);
  nand ginst14151 (P2_U4582, P2_U7892, P2_U7909, P2_U7910);
  nand ginst14152 (P2_U4583, P2_U4439, U211);
  nand ginst14153 (P2_U4584, P2_U3692, P2_U7893);
  nand ginst14154 (P2_U4585, P2_STATE_REG_2__SCAN_IN, P2_U3267);
  nand ginst14155 (P2_U4586, NA, P2_U3266);
  nand ginst14156 (P2_U4587, P2_U4585, P2_U4586);
  nand ginst14157 (P2_U4588, P2_U3258, P2_U4587);
  nand ginst14158 (P2_U4589, P2_U3263, P2_U4401);
  not ginst14159 (P2_U4590, P2_U3277);
  nand ginst14160 (P2_U4591, P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN);
  not ginst14161 (P2_U4592, P2_U3274);
  not ginst14162 (P2_U4593, P2_U3275);
  nand ginst14163 (P2_U4594, P2_STATE_REG_2__SCAN_IN, P2_U3258);
  nand ginst14164 (P2_U4595, P2_U3262, P2_U4594);
  not ginst14165 (P2_U4596, P2_U3527);
  nand ginst14166 (P2_U4597, P2_U3286, P2_U3294);
  nand ginst14167 (P2_U4598, P2_U3265, P2_U4597);
  nand ginst14168 (P2_U4599, P2_U2359, P2_U3527);
  not ginst14169 (P2_U4600, P2_U3291);
  not ginst14170 (P2_U4601, P2_U3295);
  nand ginst14171 (P2_U4602, P2_U3253, P2_U4424);
  nand ginst14172 (P2_U4603, P2_U3524, P2_U4602);
  nand ginst14173 (P2_U4604, P2_U3522, P2_U3523);
  nand ginst14174 (P2_U4605, P2_R2243_U8, P2_U4428);
  nand ginst14175 (P2_U4606, P2_U3287, P2_U4417);
  nand ginst14176 (P2_U4607, P2_U4605, P2_U4606);
  nand ginst14177 (P2_U4608, P2_U4420, P2_U4607);
  nand ginst14178 (P2_U4609, P2_U3520, P2_U4603);
  not ginst14179 (P2_U4610, P2_U3257);
  nand ginst14180 (P2_U4611, P2_U3292, P2_U4428);
  nand ginst14181 (P2_U4612, P2_GTE_370_U6, P2_U4417);
  nand ginst14182 (P2_U4613, P2_U4611, P2_U4612);
  nand ginst14183 (P2_U4614, P2_U4420, P2_U4613);
  or ginst14184 (P2_U4615, P2_FLUSH_REG_SCAN_IN, P2_MORE_REG_SCAN_IN);
  not ginst14185 (P2_U4616, P2_U3298);
  nand ginst14186 (P2_U4617, P2_U3269, P2_U4616);
  nand ginst14187 (P2_U4618, P2_U3711, P2_U4425);
  nand ginst14188 (P2_U4619, P2_U3715, P2_U8056, P2_U8057);
  not ginst14189 (P2_U4620, P2_U3299);
  nand ginst14190 (P2_U4621, P2_U3265, P2_U4474);
  nand ginst14191 (P2_U4622, P2_STATEBS16_REG_SCAN_IN, P2_U3284);
  nand ginst14192 (P2_U4623, P2_U4621, P2_U4622);
  nand ginst14193 (P2_U4624, P2_STATE2_REG_1__SCAN_IN, P2_U4623);
  nand ginst14194 (P2_U4625, P2_STATE2_REG_2__SCAN_IN, P2_U3299);
  nand ginst14195 (P2_U4626, P2_U4465, P2_U4619);
  nand ginst14196 (P2_U4627, P2_U3717, P2_U4620);
  nand ginst14197 (P2_U4628, P2_STATE2_REG_1__SCAN_IN, P2_U4626);
  nand ginst14198 (P2_U4629, P2_U2374, P2_U4619);
  nand ginst14199 (P2_U4630, P2_U3719, P2_U4469);
  nand ginst14200 (P2_U4631, P2_U4464, P2_U4619);
  nand ginst14201 (P2_U4632, P2_U2374, P2_U3298);
  not ginst14202 (P2_U4633, P2_U3337);
  not ginst14203 (P2_U4634, P2_U3351);
  not ginst14204 (P2_U4635, P2_U3352);
  not ginst14205 (P2_U4636, P2_U3319);
  not ginst14206 (P2_U4637, P2_U3318);
  not ginst14207 (P2_U4638, P2_U3378);
  nand ginst14208 (P2_U4639, P2_R2182_U76, P2_U3318);
  not ginst14209 (P2_U4640, P2_U3426);
  not ginst14210 (P2_U4641, P2_U3320);
  not ginst14211 (P2_U4642, P2_U3311);
  not ginst14212 (P2_U4643, P2_U3312);
  not ginst14213 (P2_U4644, P2_U3424);
  not ginst14214 (P2_U4645, P2_U3376);
  nand ginst14215 (P2_U4646, P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN, P2_U3311);
  not ginst14216 (P2_U4647, P2_U3428);
  not ginst14217 (P2_U4648, P2_U3349);
  not ginst14218 (P2_U4649, P2_U3335);
  not ginst14219 (P2_U4650, P2_U3243);
  nand ginst14220 (P2_U4651, P2_U2440, P2_U2444);
  not ginst14221 (P2_U4652, P2_U3325);
  not ginst14222 (P2_U4653, P2_U3570);
  not ginst14223 (P2_U4654, P2_U3326);
  nand ginst14224 (P2_U4655, P2_STATE2_REG_1__SCAN_IN, P2_U3270);
  nand ginst14225 (P2_U4656, P2_U3304, P2_U3305, P2_U4655);
  nand ginst14226 (P2_U4657, P2_U2462, P2_U4637);
  nand ginst14227 (P2_U4658, P2_U2362, P2_U2468);
  nand ginst14228 (P2_U4659, P2_U4445, P2_U4658);
  nand ginst14229 (P2_U4660, P2_U4652, P2_U4659);
  nand ginst14230 (P2_U4661, P2_STATE2_REG_2__SCAN_IN, P2_U4654);
  nand ginst14231 (P2_U4662, P2_STATE2_REG_3__SCAN_IN, P2_U3312);
  nand ginst14232 (P2_U4663, P2_U3722, P2_U4660);
  nand ginst14233 (P2_U4664, P2_U2398, P2_U2468);
  nand ginst14234 (P2_U4665, P2_U4445, P2_U4664);
  nand ginst14235 (P2_U4666, P2_U3325, P2_U4665);
  nand ginst14236 (P2_U4667, P2_STATE2_REG_2__SCAN_IN, P2_U3326);
  nand ginst14237 (P2_U4668, P2_U4666, P2_U4667);
  nand ginst14238 (P2_U4669, P2_U2425, P2_U4643);
  nand ginst14239 (P2_U4670, P2_U2422, P2_U2463);
  nand ginst14240 (P2_U4671, P2_U2421, P2_U4641);
  nand ginst14241 (P2_U4672, P2_U2406, P2_U4668);
  nand ginst14242 (P2_U4673, P2_INSTQUEUE_REG_15__7__SCAN_IN, P2_U4663);
  nand ginst14243 (P2_U4674, P2_U2426, P2_U4643);
  nand ginst14244 (P2_U4675, P2_U2420, P2_U2463);
  nand ginst14245 (P2_U4676, P2_U2419, P2_U4641);
  nand ginst14246 (P2_U4677, P2_U2405, P2_U4668);
  nand ginst14247 (P2_U4678, P2_INSTQUEUE_REG_15__6__SCAN_IN, P2_U4663);
  nand ginst14248 (P2_U4679, P2_U2429, P2_U4643);
  nand ginst14249 (P2_U4680, P2_U2418, P2_U2463);
  nand ginst14250 (P2_U4681, P2_U2417, P2_U4641);
  nand ginst14251 (P2_U4682, P2_U2404, P2_U4668);
  nand ginst14252 (P2_U4683, P2_INSTQUEUE_REG_15__5__SCAN_IN, P2_U4663);
  nand ginst14253 (P2_U4684, P2_U2424, P2_U4643);
  nand ginst14254 (P2_U4685, P2_U2416, P2_U2463);
  nand ginst14255 (P2_U4686, P2_U2415, P2_U4641);
  nand ginst14256 (P2_U4687, P2_U2403, P2_U4668);
  nand ginst14257 (P2_U4688, P2_INSTQUEUE_REG_15__4__SCAN_IN, P2_U4663);
  nand ginst14258 (P2_U4689, P2_U2423, P2_U4643);
  nand ginst14259 (P2_U4690, P2_U2414, P2_U2463);
  nand ginst14260 (P2_U4691, P2_U2413, P2_U4641);
  nand ginst14261 (P2_U4692, P2_U2402, P2_U4668);
  nand ginst14262 (P2_U4693, P2_INSTQUEUE_REG_15__3__SCAN_IN, P2_U4663);
  nand ginst14263 (P2_U4694, P2_U2432, P2_U4643);
  nand ginst14264 (P2_U4695, P2_U2412, P2_U2463);
  nand ginst14265 (P2_U4696, P2_U2411, P2_U4641);
  nand ginst14266 (P2_U4697, P2_U2401, P2_U4668);
  nand ginst14267 (P2_U4698, P2_INSTQUEUE_REG_15__2__SCAN_IN, P2_U4663);
  nand ginst14268 (P2_U4699, P2_U2428, P2_U4643);
  nand ginst14269 (P2_U4700, P2_U2410, P2_U2463);
  nand ginst14270 (P2_U4701, P2_U2409, P2_U4641);
  nand ginst14271 (P2_U4702, P2_U2400, P2_U4668);
  nand ginst14272 (P2_U4703, P2_INSTQUEUE_REG_15__1__SCAN_IN, P2_U4663);
  nand ginst14273 (P2_U4704, P2_U2431, P2_U4643);
  nand ginst14274 (P2_U4705, P2_U2408, P2_U2463);
  nand ginst14275 (P2_U4706, P2_U2407, P2_U4641);
  nand ginst14276 (P2_U4707, P2_U2399, P2_U4668);
  nand ginst14277 (P2_U4708, P2_INSTQUEUE_REG_15__0__SCAN_IN, P2_U4663);
  not ginst14278 (P2_U4709, P2_U3338);
  not ginst14279 (P2_U4710, P2_U3339);
  not ginst14280 (P2_U4711, P2_U3336);
  not ginst14281 (P2_U4712, P2_U3245);
  not ginst14282 (P2_U4713, P2_U3569);
  not ginst14283 (P2_U4714, P2_U3340);
  nand ginst14284 (P2_U4715, P2_U2462, P2_U4633);
  nand ginst14285 (P2_U4716, P2_U2362, P2_U2471);
  nand ginst14286 (P2_U4717, P2_U4445, P2_U4716);
  nand ginst14287 (P2_U4718, P2_U3245, P2_U4717);
  nand ginst14288 (P2_U4719, P2_STATE2_REG_2__SCAN_IN, P2_U4714);
  nand ginst14289 (P2_U4720, P2_STATE2_REG_3__SCAN_IN, P2_U3336);
  nand ginst14290 (P2_U4721, P2_U3731, P2_U4718);
  nand ginst14291 (P2_U4722, P2_U2398, P2_U2471);
  nand ginst14292 (P2_U4723, P2_U4445, P2_U4722);
  nand ginst14293 (P2_U4724, P2_U4712, P2_U4723);
  nand ginst14294 (P2_U4725, P2_STATE2_REG_2__SCAN_IN, P2_U3340);
  nand ginst14295 (P2_U4726, P2_U4724, P2_U4725);
  nand ginst14296 (P2_U4727, P2_U2425, P2_U4711);
  nand ginst14297 (P2_U4728, P2_U2422, P2_U2469);
  nand ginst14298 (P2_U4729, P2_U2421, P2_U4710);
  nand ginst14299 (P2_U4730, P2_U2406, P2_U4726);
  nand ginst14300 (P2_U4731, P2_INSTQUEUE_REG_14__7__SCAN_IN, P2_U4721);
  nand ginst14301 (P2_U4732, P2_U2426, P2_U4711);
  nand ginst14302 (P2_U4733, P2_U2420, P2_U2469);
  nand ginst14303 (P2_U4734, P2_U2419, P2_U4710);
  nand ginst14304 (P2_U4735, P2_U2405, P2_U4726);
  nand ginst14305 (P2_U4736, P2_INSTQUEUE_REG_14__6__SCAN_IN, P2_U4721);
  nand ginst14306 (P2_U4737, P2_U2429, P2_U4711);
  nand ginst14307 (P2_U4738, P2_U2418, P2_U2469);
  nand ginst14308 (P2_U4739, P2_U2417, P2_U4710);
  nand ginst14309 (P2_U4740, P2_U2404, P2_U4726);
  nand ginst14310 (P2_U4741, P2_INSTQUEUE_REG_14__5__SCAN_IN, P2_U4721);
  nand ginst14311 (P2_U4742, P2_U2424, P2_U4711);
  nand ginst14312 (P2_U4743, P2_U2416, P2_U2469);
  nand ginst14313 (P2_U4744, P2_U2415, P2_U4710);
  nand ginst14314 (P2_U4745, P2_U2403, P2_U4726);
  nand ginst14315 (P2_U4746, P2_INSTQUEUE_REG_14__4__SCAN_IN, P2_U4721);
  nand ginst14316 (P2_U4747, P2_U2423, P2_U4711);
  nand ginst14317 (P2_U4748, P2_U2414, P2_U2469);
  nand ginst14318 (P2_U4749, P2_U2413, P2_U4710);
  nand ginst14319 (P2_U4750, P2_U2402, P2_U4726);
  nand ginst14320 (P2_U4751, P2_INSTQUEUE_REG_14__3__SCAN_IN, P2_U4721);
  nand ginst14321 (P2_U4752, P2_U2432, P2_U4711);
  nand ginst14322 (P2_U4753, P2_U2412, P2_U2469);
  nand ginst14323 (P2_U4754, P2_U2411, P2_U4710);
  nand ginst14324 (P2_U4755, P2_U2401, P2_U4726);
  nand ginst14325 (P2_U4756, P2_INSTQUEUE_REG_14__2__SCAN_IN, P2_U4721);
  nand ginst14326 (P2_U4757, P2_U2428, P2_U4711);
  nand ginst14327 (P2_U4758, P2_U2410, P2_U2469);
  nand ginst14328 (P2_U4759, P2_U2409, P2_U4710);
  nand ginst14329 (P2_U4760, P2_U2400, P2_U4726);
  nand ginst14330 (P2_U4761, P2_INSTQUEUE_REG_14__1__SCAN_IN, P2_U4721);
  nand ginst14331 (P2_U4762, P2_U2431, P2_U4711);
  nand ginst14332 (P2_U4763, P2_U2408, P2_U2469);
  nand ginst14333 (P2_U4764, P2_U2407, P2_U4710);
  nand ginst14334 (P2_U4765, P2_U2399, P2_U4726);
  nand ginst14335 (P2_U4766, P2_INSTQUEUE_REG_14__0__SCAN_IN, P2_U4721);
  not ginst14336 (P2_U4767, P2_U3353);
  not ginst14337 (P2_U4768, P2_U3354);
  not ginst14338 (P2_U4769, P2_U3350);
  nand ginst14339 (P2_U4770, P2_U2440, P2_U2445);
  not ginst14340 (P2_U4771, P2_U3355);
  not ginst14341 (P2_U4772, P2_U3568);
  not ginst14342 (P2_U4773, P2_U3356);
  nand ginst14343 (P2_U4774, P2_U2462, P2_U4634);
  nand ginst14344 (P2_U4775, P2_U2362, P2_U2474);
  nand ginst14345 (P2_U4776, P2_U4445, P2_U4775);
  nand ginst14346 (P2_U4777, P2_U4771, P2_U4776);
  nand ginst14347 (P2_U4778, P2_STATE2_REG_2__SCAN_IN, P2_U4773);
  nand ginst14348 (P2_U4779, P2_STATE2_REG_3__SCAN_IN, P2_U3350);
  nand ginst14349 (P2_U4780, P2_U3740, P2_U4777);
  nand ginst14350 (P2_U4781, P2_U2398, P2_U2474);
  nand ginst14351 (P2_U4782, P2_U4445, P2_U4781);
  nand ginst14352 (P2_U4783, P2_U3355, P2_U4782);
  nand ginst14353 (P2_U4784, P2_STATE2_REG_2__SCAN_IN, P2_U3356);
  nand ginst14354 (P2_U4785, P2_U4783, P2_U4784);
  nand ginst14355 (P2_U4786, P2_U2425, P2_U4769);
  nand ginst14356 (P2_U4787, P2_U2422, P2_U2472);
  nand ginst14357 (P2_U4788, P2_U2421, P2_U4768);
  nand ginst14358 (P2_U4789, P2_U2406, P2_U4785);
  nand ginst14359 (P2_U4790, P2_INSTQUEUE_REG_13__7__SCAN_IN, P2_U4780);
  nand ginst14360 (P2_U4791, P2_U2426, P2_U4769);
  nand ginst14361 (P2_U4792, P2_U2420, P2_U2472);
  nand ginst14362 (P2_U4793, P2_U2419, P2_U4768);
  nand ginst14363 (P2_U4794, P2_U2405, P2_U4785);
  nand ginst14364 (P2_U4795, P2_INSTQUEUE_REG_13__6__SCAN_IN, P2_U4780);
  nand ginst14365 (P2_U4796, P2_U2429, P2_U4769);
  nand ginst14366 (P2_U4797, P2_U2418, P2_U2472);
  nand ginst14367 (P2_U4798, P2_U2417, P2_U4768);
  nand ginst14368 (P2_U4799, P2_U2404, P2_U4785);
  nand ginst14369 (P2_U4800, P2_INSTQUEUE_REG_13__5__SCAN_IN, P2_U4780);
  nand ginst14370 (P2_U4801, P2_U2424, P2_U4769);
  nand ginst14371 (P2_U4802, P2_U2416, P2_U2472);
  nand ginst14372 (P2_U4803, P2_U2415, P2_U4768);
  nand ginst14373 (P2_U4804, P2_U2403, P2_U4785);
  nand ginst14374 (P2_U4805, P2_INSTQUEUE_REG_13__4__SCAN_IN, P2_U4780);
  nand ginst14375 (P2_U4806, P2_U2423, P2_U4769);
  nand ginst14376 (P2_U4807, P2_U2414, P2_U2472);
  nand ginst14377 (P2_U4808, P2_U2413, P2_U4768);
  nand ginst14378 (P2_U4809, P2_U2402, P2_U4785);
  nand ginst14379 (P2_U4810, P2_INSTQUEUE_REG_13__3__SCAN_IN, P2_U4780);
  nand ginst14380 (P2_U4811, P2_U2432, P2_U4769);
  nand ginst14381 (P2_U4812, P2_U2412, P2_U2472);
  nand ginst14382 (P2_U4813, P2_U2411, P2_U4768);
  nand ginst14383 (P2_U4814, P2_U2401, P2_U4785);
  nand ginst14384 (P2_U4815, P2_INSTQUEUE_REG_13__2__SCAN_IN, P2_U4780);
  nand ginst14385 (P2_U4816, P2_U2428, P2_U4769);
  nand ginst14386 (P2_U4817, P2_U2410, P2_U2472);
  nand ginst14387 (P2_U4818, P2_U2409, P2_U4768);
  nand ginst14388 (P2_U4819, P2_U2400, P2_U4785);
  nand ginst14389 (P2_U4820, P2_INSTQUEUE_REG_13__1__SCAN_IN, P2_U4780);
  nand ginst14390 (P2_U4821, P2_U2431, P2_U4769);
  nand ginst14391 (P2_U4822, P2_U2408, P2_U2472);
  nand ginst14392 (P2_U4823, P2_U2407, P2_U4768);
  nand ginst14393 (P2_U4824, P2_U2399, P2_U4785);
  nand ginst14394 (P2_U4825, P2_INSTQUEUE_REG_13__0__SCAN_IN, P2_U4780);
  not ginst14395 (P2_U4826, P2_U3366);
  not ginst14396 (P2_U4827, P2_U3365);
  not ginst14397 (P2_U4828, P2_U3246);
  not ginst14398 (P2_U4829, P2_U3567);
  not ginst14399 (P2_U4830, P2_U3367);
  nand ginst14400 (P2_U4831, P2_U2462, P2_U2476);
  nand ginst14401 (P2_U4832, P2_U2362, P2_U2480);
  nand ginst14402 (P2_U4833, P2_U4445, P2_U4832);
  nand ginst14403 (P2_U4834, P2_U3246, P2_U4833);
  nand ginst14404 (P2_U4835, P2_STATE2_REG_2__SCAN_IN, P2_U4830);
  nand ginst14405 (P2_U4836, P2_STATE2_REG_3__SCAN_IN, P2_U3365);
  nand ginst14406 (P2_U4837, P2_U3749, P2_U4834);
  nand ginst14407 (P2_U4838, P2_U2398, P2_U2480);
  nand ginst14408 (P2_U4839, P2_U4445, P2_U4838);
  nand ginst14409 (P2_U4840, P2_U4828, P2_U4839);
  nand ginst14410 (P2_U4841, P2_STATE2_REG_2__SCAN_IN, P2_U3367);
  nand ginst14411 (P2_U4842, P2_U4840, P2_U4841);
  nand ginst14412 (P2_U4843, P2_U2425, P2_U4827);
  nand ginst14413 (P2_U4844, P2_U2422, P2_U2477);
  nand ginst14414 (P2_U4845, P2_U2421, P2_U4826);
  nand ginst14415 (P2_U4846, P2_U2406, P2_U4842);
  nand ginst14416 (P2_U4847, P2_INSTQUEUE_REG_12__7__SCAN_IN, P2_U4837);
  nand ginst14417 (P2_U4848, P2_U2426, P2_U4827);
  nand ginst14418 (P2_U4849, P2_U2420, P2_U2477);
  nand ginst14419 (P2_U4850, P2_U2419, P2_U4826);
  nand ginst14420 (P2_U4851, P2_U2405, P2_U4842);
  nand ginst14421 (P2_U4852, P2_INSTQUEUE_REG_12__6__SCAN_IN, P2_U4837);
  nand ginst14422 (P2_U4853, P2_U2429, P2_U4827);
  nand ginst14423 (P2_U4854, P2_U2418, P2_U2477);
  nand ginst14424 (P2_U4855, P2_U2417, P2_U4826);
  nand ginst14425 (P2_U4856, P2_U2404, P2_U4842);
  nand ginst14426 (P2_U4857, P2_INSTQUEUE_REG_12__5__SCAN_IN, P2_U4837);
  nand ginst14427 (P2_U4858, P2_U2424, P2_U4827);
  nand ginst14428 (P2_U4859, P2_U2416, P2_U2477);
  nand ginst14429 (P2_U4860, P2_U2415, P2_U4826);
  nand ginst14430 (P2_U4861, P2_U2403, P2_U4842);
  nand ginst14431 (P2_U4862, P2_INSTQUEUE_REG_12__4__SCAN_IN, P2_U4837);
  nand ginst14432 (P2_U4863, P2_U2423, P2_U4827);
  nand ginst14433 (P2_U4864, P2_U2414, P2_U2477);
  nand ginst14434 (P2_U4865, P2_U2413, P2_U4826);
  nand ginst14435 (P2_U4866, P2_U2402, P2_U4842);
  nand ginst14436 (P2_U4867, P2_INSTQUEUE_REG_12__3__SCAN_IN, P2_U4837);
  nand ginst14437 (P2_U4868, P2_U2432, P2_U4827);
  nand ginst14438 (P2_U4869, P2_U2412, P2_U2477);
  nand ginst14439 (P2_U4870, P2_U2411, P2_U4826);
  nand ginst14440 (P2_U4871, P2_U2401, P2_U4842);
  nand ginst14441 (P2_U4872, P2_INSTQUEUE_REG_12__2__SCAN_IN, P2_U4837);
  nand ginst14442 (P2_U4873, P2_U2428, P2_U4827);
  nand ginst14443 (P2_U4874, P2_U2410, P2_U2477);
  nand ginst14444 (P2_U4875, P2_U2409, P2_U4826);
  nand ginst14445 (P2_U4876, P2_U2400, P2_U4842);
  nand ginst14446 (P2_U4877, P2_INSTQUEUE_REG_12__1__SCAN_IN, P2_U4837);
  nand ginst14447 (P2_U4878, P2_U2431, P2_U4827);
  nand ginst14448 (P2_U4879, P2_U2408, P2_U2477);
  nand ginst14449 (P2_U4880, P2_U2407, P2_U4826);
  nand ginst14450 (P2_U4881, P2_U2399, P2_U4842);
  nand ginst14451 (P2_U4882, P2_INSTQUEUE_REG_12__0__SCAN_IN, P2_U4837);
  not ginst14452 (P2_U4883, P2_U3379);
  not ginst14453 (P2_U4884, P2_U3377);
  nand ginst14454 (P2_U4885, P2_U2442, P2_U2444);
  not ginst14455 (P2_U4886, P2_U3380);
  not ginst14456 (P2_U4887, P2_U3566);
  not ginst14457 (P2_U4888, P2_U3381);
  nand ginst14458 (P2_U4889, P2_U4637, P2_U4638);
  nand ginst14459 (P2_U4890, P2_U2362, P2_U2484);
  nand ginst14460 (P2_U4891, P2_U4445, P2_U4890);
  nand ginst14461 (P2_U4892, P2_U4886, P2_U4891);
  nand ginst14462 (P2_U4893, P2_STATE2_REG_2__SCAN_IN, P2_U4888);
  nand ginst14463 (P2_U4894, P2_STATE2_REG_3__SCAN_IN, P2_U3377);
  nand ginst14464 (P2_U4895, P2_U3758, P2_U4892);
  nand ginst14465 (P2_U4896, P2_U2398, P2_U2484);
  nand ginst14466 (P2_U4897, P2_U4445, P2_U4896);
  nand ginst14467 (P2_U4898, P2_U3380, P2_U4897);
  nand ginst14468 (P2_U4899, P2_STATE2_REG_2__SCAN_IN, P2_U3381);
  nand ginst14469 (P2_U4900, P2_U4898, P2_U4899);
  nand ginst14470 (P2_U4901, P2_U2425, P2_U4884);
  nand ginst14471 (P2_U4902, P2_U2422, P2_U2482);
  nand ginst14472 (P2_U4903, P2_U2421, P2_U4883);
  nand ginst14473 (P2_U4904, P2_U2406, P2_U4900);
  nand ginst14474 (P2_U4905, P2_INSTQUEUE_REG_11__7__SCAN_IN, P2_U4895);
  nand ginst14475 (P2_U4906, P2_U2426, P2_U4884);
  nand ginst14476 (P2_U4907, P2_U2420, P2_U2482);
  nand ginst14477 (P2_U4908, P2_U2419, P2_U4883);
  nand ginst14478 (P2_U4909, P2_U2405, P2_U4900);
  nand ginst14479 (P2_U4910, P2_INSTQUEUE_REG_11__6__SCAN_IN, P2_U4895);
  nand ginst14480 (P2_U4911, P2_U2429, P2_U4884);
  nand ginst14481 (P2_U4912, P2_U2418, P2_U2482);
  nand ginst14482 (P2_U4913, P2_U2417, P2_U4883);
  nand ginst14483 (P2_U4914, P2_U2404, P2_U4900);
  nand ginst14484 (P2_U4915, P2_INSTQUEUE_REG_11__5__SCAN_IN, P2_U4895);
  nand ginst14485 (P2_U4916, P2_U2424, P2_U4884);
  nand ginst14486 (P2_U4917, P2_U2416, P2_U2482);
  nand ginst14487 (P2_U4918, P2_U2415, P2_U4883);
  nand ginst14488 (P2_U4919, P2_U2403, P2_U4900);
  nand ginst14489 (P2_U4920, P2_INSTQUEUE_REG_11__4__SCAN_IN, P2_U4895);
  nand ginst14490 (P2_U4921, P2_U2423, P2_U4884);
  nand ginst14491 (P2_U4922, P2_U2414, P2_U2482);
  nand ginst14492 (P2_U4923, P2_U2413, P2_U4883);
  nand ginst14493 (P2_U4924, P2_U2402, P2_U4900);
  nand ginst14494 (P2_U4925, P2_INSTQUEUE_REG_11__3__SCAN_IN, P2_U4895);
  nand ginst14495 (P2_U4926, P2_U2432, P2_U4884);
  nand ginst14496 (P2_U4927, P2_U2412, P2_U2482);
  nand ginst14497 (P2_U4928, P2_U2411, P2_U4883);
  nand ginst14498 (P2_U4929, P2_U2401, P2_U4900);
  nand ginst14499 (P2_U4930, P2_INSTQUEUE_REG_11__2__SCAN_IN, P2_U4895);
  nand ginst14500 (P2_U4931, P2_U2428, P2_U4884);
  nand ginst14501 (P2_U4932, P2_U2410, P2_U2482);
  nand ginst14502 (P2_U4933, P2_U2409, P2_U4883);
  nand ginst14503 (P2_U4934, P2_U2400, P2_U4900);
  nand ginst14504 (P2_U4935, P2_INSTQUEUE_REG_11__1__SCAN_IN, P2_U4895);
  nand ginst14505 (P2_U4936, P2_U2431, P2_U4884);
  nand ginst14506 (P2_U4937, P2_U2408, P2_U2482);
  nand ginst14507 (P2_U4938, P2_U2407, P2_U4883);
  nand ginst14508 (P2_U4939, P2_U2399, P2_U4900);
  nand ginst14509 (P2_U4940, P2_INSTQUEUE_REG_11__0__SCAN_IN, P2_U4895);
  not ginst14510 (P2_U4941, P2_U3391);
  not ginst14511 (P2_U4942, P2_U3390);
  not ginst14512 (P2_U4943, P2_U3247);
  not ginst14513 (P2_U4944, P2_U3565);
  not ginst14514 (P2_U4945, P2_U3392);
  nand ginst14515 (P2_U4946, P2_U4633, P2_U4638);
  nand ginst14516 (P2_U4947, P2_U2362, P2_U2486);
  nand ginst14517 (P2_U4948, P2_U4445, P2_U4947);
  nand ginst14518 (P2_U4949, P2_U3247, P2_U4948);
  nand ginst14519 (P2_U4950, P2_STATE2_REG_2__SCAN_IN, P2_U4945);
  nand ginst14520 (P2_U4951, P2_STATE2_REG_3__SCAN_IN, P2_U3390);
  nand ginst14521 (P2_U4952, P2_U3767, P2_U4949);
  nand ginst14522 (P2_U4953, P2_U2398, P2_U2486);
  nand ginst14523 (P2_U4954, P2_U4445, P2_U4953);
  nand ginst14524 (P2_U4955, P2_U4943, P2_U4954);
  nand ginst14525 (P2_U4956, P2_STATE2_REG_2__SCAN_IN, P2_U3392);
  nand ginst14526 (P2_U4957, P2_U4955, P2_U4956);
  nand ginst14527 (P2_U4958, P2_U2425, P2_U4942);
  nand ginst14528 (P2_U4959, P2_U2422, P2_U2485);
  nand ginst14529 (P2_U4960, P2_U2421, P2_U4941);
  nand ginst14530 (P2_U4961, P2_U2406, P2_U4957);
  nand ginst14531 (P2_U4962, P2_INSTQUEUE_REG_10__7__SCAN_IN, P2_U4952);
  nand ginst14532 (P2_U4963, P2_U2426, P2_U4942);
  nand ginst14533 (P2_U4964, P2_U2420, P2_U2485);
  nand ginst14534 (P2_U4965, P2_U2419, P2_U4941);
  nand ginst14535 (P2_U4966, P2_U2405, P2_U4957);
  nand ginst14536 (P2_U4967, P2_INSTQUEUE_REG_10__6__SCAN_IN, P2_U4952);
  nand ginst14537 (P2_U4968, P2_U2429, P2_U4942);
  nand ginst14538 (P2_U4969, P2_U2418, P2_U2485);
  nand ginst14539 (P2_U4970, P2_U2417, P2_U4941);
  nand ginst14540 (P2_U4971, P2_U2404, P2_U4957);
  nand ginst14541 (P2_U4972, P2_INSTQUEUE_REG_10__5__SCAN_IN, P2_U4952);
  nand ginst14542 (P2_U4973, P2_U2424, P2_U4942);
  nand ginst14543 (P2_U4974, P2_U2416, P2_U2485);
  nand ginst14544 (P2_U4975, P2_U2415, P2_U4941);
  nand ginst14545 (P2_U4976, P2_U2403, P2_U4957);
  nand ginst14546 (P2_U4977, P2_INSTQUEUE_REG_10__4__SCAN_IN, P2_U4952);
  nand ginst14547 (P2_U4978, P2_U2423, P2_U4942);
  nand ginst14548 (P2_U4979, P2_U2414, P2_U2485);
  nand ginst14549 (P2_U4980, P2_U2413, P2_U4941);
  nand ginst14550 (P2_U4981, P2_U2402, P2_U4957);
  nand ginst14551 (P2_U4982, P2_INSTQUEUE_REG_10__3__SCAN_IN, P2_U4952);
  nand ginst14552 (P2_U4983, P2_U2432, P2_U4942);
  nand ginst14553 (P2_U4984, P2_U2412, P2_U2485);
  nand ginst14554 (P2_U4985, P2_U2411, P2_U4941);
  nand ginst14555 (P2_U4986, P2_U2401, P2_U4957);
  nand ginst14556 (P2_U4987, P2_INSTQUEUE_REG_10__2__SCAN_IN, P2_U4952);
  nand ginst14557 (P2_U4988, P2_U2428, P2_U4942);
  nand ginst14558 (P2_U4989, P2_U2410, P2_U2485);
  nand ginst14559 (P2_U4990, P2_U2409, P2_U4941);
  nand ginst14560 (P2_U4991, P2_U2400, P2_U4957);
  nand ginst14561 (P2_U4992, P2_INSTQUEUE_REG_10__1__SCAN_IN, P2_U4952);
  nand ginst14562 (P2_U4993, P2_U2431, P2_U4942);
  nand ginst14563 (P2_U4994, P2_U2408, P2_U2485);
  nand ginst14564 (P2_U4995, P2_U2407, P2_U4941);
  nand ginst14565 (P2_U4996, P2_U2399, P2_U4957);
  nand ginst14566 (P2_U4997, P2_INSTQUEUE_REG_10__0__SCAN_IN, P2_U4952);
  not ginst14567 (P2_U4998, P2_U3402);
  not ginst14568 (P2_U4999, P2_U3401);
  nand ginst14569 (P2_U5000, P2_U2442, P2_U2445);
  not ginst14570 (P2_U5001, P2_U3403);
  not ginst14571 (P2_U5002, P2_U3564);
  not ginst14572 (P2_U5003, P2_U3404);
  nand ginst14573 (P2_U5004, P2_U4634, P2_U4638);
  nand ginst14574 (P2_U5005, P2_U2362, P2_U2488);
  nand ginst14575 (P2_U5006, P2_U4445, P2_U5005);
  nand ginst14576 (P2_U5007, P2_U5001, P2_U5006);
  nand ginst14577 (P2_U5008, P2_STATE2_REG_2__SCAN_IN, P2_U5003);
  nand ginst14578 (P2_U5009, P2_STATE2_REG_3__SCAN_IN, P2_U3401);
  nand ginst14579 (P2_U5010, P2_U3776, P2_U5007);
  nand ginst14580 (P2_U5011, P2_U2398, P2_U2488);
  nand ginst14581 (P2_U5012, P2_U4445, P2_U5011);
  nand ginst14582 (P2_U5013, P2_U3403, P2_U5012);
  nand ginst14583 (P2_U5014, P2_STATE2_REG_2__SCAN_IN, P2_U3404);
  nand ginst14584 (P2_U5015, P2_U5013, P2_U5014);
  nand ginst14585 (P2_U5016, P2_U2425, P2_U4999);
  nand ginst14586 (P2_U5017, P2_U2422, P2_U2487);
  nand ginst14587 (P2_U5018, P2_U2421, P2_U4998);
  nand ginst14588 (P2_U5019, P2_U2406, P2_U5015);
  nand ginst14589 (P2_U5020, P2_INSTQUEUE_REG_9__7__SCAN_IN, P2_U5010);
  nand ginst14590 (P2_U5021, P2_U2426, P2_U4999);
  nand ginst14591 (P2_U5022, P2_U2420, P2_U2487);
  nand ginst14592 (P2_U5023, P2_U2419, P2_U4998);
  nand ginst14593 (P2_U5024, P2_U2405, P2_U5015);
  nand ginst14594 (P2_U5025, P2_INSTQUEUE_REG_9__6__SCAN_IN, P2_U5010);
  nand ginst14595 (P2_U5026, P2_U2429, P2_U4999);
  nand ginst14596 (P2_U5027, P2_U2418, P2_U2487);
  nand ginst14597 (P2_U5028, P2_U2417, P2_U4998);
  nand ginst14598 (P2_U5029, P2_U2404, P2_U5015);
  nand ginst14599 (P2_U5030, P2_INSTQUEUE_REG_9__5__SCAN_IN, P2_U5010);
  nand ginst14600 (P2_U5031, P2_U2424, P2_U4999);
  nand ginst14601 (P2_U5032, P2_U2416, P2_U2487);
  nand ginst14602 (P2_U5033, P2_U2415, P2_U4998);
  nand ginst14603 (P2_U5034, P2_U2403, P2_U5015);
  nand ginst14604 (P2_U5035, P2_INSTQUEUE_REG_9__4__SCAN_IN, P2_U5010);
  nand ginst14605 (P2_U5036, P2_U2423, P2_U4999);
  nand ginst14606 (P2_U5037, P2_U2414, P2_U2487);
  nand ginst14607 (P2_U5038, P2_U2413, P2_U4998);
  nand ginst14608 (P2_U5039, P2_U2402, P2_U5015);
  nand ginst14609 (P2_U5040, P2_INSTQUEUE_REG_9__3__SCAN_IN, P2_U5010);
  nand ginst14610 (P2_U5041, P2_U2432, P2_U4999);
  nand ginst14611 (P2_U5042, P2_U2412, P2_U2487);
  nand ginst14612 (P2_U5043, P2_U2411, P2_U4998);
  nand ginst14613 (P2_U5044, P2_U2401, P2_U5015);
  nand ginst14614 (P2_U5045, P2_INSTQUEUE_REG_9__2__SCAN_IN, P2_U5010);
  nand ginst14615 (P2_U5046, P2_U2428, P2_U4999);
  nand ginst14616 (P2_U5047, P2_U2410, P2_U2487);
  nand ginst14617 (P2_U5048, P2_U2409, P2_U4998);
  nand ginst14618 (P2_U5049, P2_U2400, P2_U5015);
  nand ginst14619 (P2_U5050, P2_INSTQUEUE_REG_9__1__SCAN_IN, P2_U5010);
  nand ginst14620 (P2_U5051, P2_U2431, P2_U4999);
  nand ginst14621 (P2_U5052, P2_U2408, P2_U2487);
  nand ginst14622 (P2_U5053, P2_U2407, P2_U4998);
  nand ginst14623 (P2_U5054, P2_U2399, P2_U5015);
  nand ginst14624 (P2_U5055, P2_INSTQUEUE_REG_9__0__SCAN_IN, P2_U5010);
  not ginst14625 (P2_U5056, P2_U3414);
  not ginst14626 (P2_U5057, P2_U3413);
  not ginst14627 (P2_U5058, P2_U3248);
  not ginst14628 (P2_U5059, P2_U3563);
  not ginst14629 (P2_U5060, P2_U3415);
  nand ginst14630 (P2_U5061, P2_U2476, P2_U4638);
  nand ginst14631 (P2_U5062, P2_U2362, P2_U2490);
  nand ginst14632 (P2_U5063, P2_U4445, P2_U5062);
  nand ginst14633 (P2_U5064, P2_U3248, P2_U5063);
  nand ginst14634 (P2_U5065, P2_STATE2_REG_2__SCAN_IN, P2_U5060);
  nand ginst14635 (P2_U5066, P2_STATE2_REG_3__SCAN_IN, P2_U3413);
  nand ginst14636 (P2_U5067, P2_U3785, P2_U5064);
  nand ginst14637 (P2_U5068, P2_U2398, P2_U2490);
  nand ginst14638 (P2_U5069, P2_U4445, P2_U5068);
  nand ginst14639 (P2_U5070, P2_U5058, P2_U5069);
  nand ginst14640 (P2_U5071, P2_STATE2_REG_2__SCAN_IN, P2_U3415);
  nand ginst14641 (P2_U5072, P2_U5070, P2_U5071);
  nand ginst14642 (P2_U5073, P2_U2425, P2_U5057);
  nand ginst14643 (P2_U5074, P2_U2422, P2_U2489);
  nand ginst14644 (P2_U5075, P2_U2421, P2_U5056);
  nand ginst14645 (P2_U5076, P2_U2406, P2_U5072);
  nand ginst14646 (P2_U5077, P2_INSTQUEUE_REG_8__7__SCAN_IN, P2_U5067);
  nand ginst14647 (P2_U5078, P2_U2426, P2_U5057);
  nand ginst14648 (P2_U5079, P2_U2420, P2_U2489);
  nand ginst14649 (P2_U5080, P2_U2419, P2_U5056);
  nand ginst14650 (P2_U5081, P2_U2405, P2_U5072);
  nand ginst14651 (P2_U5082, P2_INSTQUEUE_REG_8__6__SCAN_IN, P2_U5067);
  nand ginst14652 (P2_U5083, P2_U2429, P2_U5057);
  nand ginst14653 (P2_U5084, P2_U2418, P2_U2489);
  nand ginst14654 (P2_U5085, P2_U2417, P2_U5056);
  nand ginst14655 (P2_U5086, P2_U2404, P2_U5072);
  nand ginst14656 (P2_U5087, P2_INSTQUEUE_REG_8__5__SCAN_IN, P2_U5067);
  nand ginst14657 (P2_U5088, P2_U2424, P2_U5057);
  nand ginst14658 (P2_U5089, P2_U2416, P2_U2489);
  nand ginst14659 (P2_U5090, P2_U2415, P2_U5056);
  nand ginst14660 (P2_U5091, P2_U2403, P2_U5072);
  nand ginst14661 (P2_U5092, P2_INSTQUEUE_REG_8__4__SCAN_IN, P2_U5067);
  nand ginst14662 (P2_U5093, P2_U2423, P2_U5057);
  nand ginst14663 (P2_U5094, P2_U2414, P2_U2489);
  nand ginst14664 (P2_U5095, P2_U2413, P2_U5056);
  nand ginst14665 (P2_U5096, P2_U2402, P2_U5072);
  nand ginst14666 (P2_U5097, P2_INSTQUEUE_REG_8__3__SCAN_IN, P2_U5067);
  nand ginst14667 (P2_U5098, P2_U2432, P2_U5057);
  nand ginst14668 (P2_U5099, P2_U2412, P2_U2489);
  nand ginst14669 (P2_U5100, P2_U2411, P2_U5056);
  nand ginst14670 (P2_U5101, P2_U2401, P2_U5072);
  nand ginst14671 (P2_U5102, P2_INSTQUEUE_REG_8__2__SCAN_IN, P2_U5067);
  nand ginst14672 (P2_U5103, P2_U2428, P2_U5057);
  nand ginst14673 (P2_U5104, P2_U2410, P2_U2489);
  nand ginst14674 (P2_U5105, P2_U2409, P2_U5056);
  nand ginst14675 (P2_U5106, P2_U2400, P2_U5072);
  nand ginst14676 (P2_U5107, P2_INSTQUEUE_REG_8__1__SCAN_IN, P2_U5067);
  nand ginst14677 (P2_U5108, P2_U2431, P2_U5057);
  nand ginst14678 (P2_U5109, P2_U2408, P2_U2489);
  nand ginst14679 (P2_U5110, P2_U2407, P2_U5056);
  nand ginst14680 (P2_U5111, P2_U2399, P2_U5072);
  nand ginst14681 (P2_U5112, P2_INSTQUEUE_REG_8__0__SCAN_IN, P2_U5067);
  not ginst14682 (P2_U5113, P2_U3427);
  nand ginst14683 (P2_U5114, P2_U2441, P2_U2444);
  not ginst14684 (P2_U5115, P2_U3429);
  not ginst14685 (P2_U5116, P2_U3562);
  not ginst14686 (P2_U5117, P2_U3430);
  nand ginst14687 (P2_U5118, P2_U2362, P2_U2493);
  nand ginst14688 (P2_U5119, P2_U4445, P2_U5118);
  nand ginst14689 (P2_U5120, P2_U5115, P2_U5119);
  nand ginst14690 (P2_U5121, P2_STATE2_REG_2__SCAN_IN, P2_U5117);
  nand ginst14691 (P2_U5122, P2_STATE2_REG_3__SCAN_IN, P2_U3424);
  nand ginst14692 (P2_U5123, P2_U3794, P2_U5120);
  nand ginst14693 (P2_U5124, P2_U2398, P2_U2493);
  nand ginst14694 (P2_U5125, P2_U4445, P2_U5124);
  nand ginst14695 (P2_U5126, P2_U3429, P2_U5125);
  nand ginst14696 (P2_U5127, P2_STATE2_REG_2__SCAN_IN, P2_U3430);
  nand ginst14697 (P2_U5128, P2_U5126, P2_U5127);
  nand ginst14698 (P2_U5129, P2_U2425, P2_U4644);
  nand ginst14699 (P2_U5130, P2_U2422, P2_U4451);
  nand ginst14700 (P2_U5131, P2_U2421, P2_U5113);
  nand ginst14701 (P2_U5132, P2_U2406, P2_U5128);
  nand ginst14702 (P2_U5133, P2_INSTQUEUE_REG_7__7__SCAN_IN, P2_U5123);
  nand ginst14703 (P2_U5134, P2_U2426, P2_U4644);
  nand ginst14704 (P2_U5135, P2_U2420, P2_U4451);
  nand ginst14705 (P2_U5136, P2_U2419, P2_U5113);
  nand ginst14706 (P2_U5137, P2_U2405, P2_U5128);
  nand ginst14707 (P2_U5138, P2_INSTQUEUE_REG_7__6__SCAN_IN, P2_U5123);
  nand ginst14708 (P2_U5139, P2_U2429, P2_U4644);
  nand ginst14709 (P2_U5140, P2_U2418, P2_U4451);
  nand ginst14710 (P2_U5141, P2_U2417, P2_U5113);
  nand ginst14711 (P2_U5142, P2_U2404, P2_U5128);
  nand ginst14712 (P2_U5143, P2_INSTQUEUE_REG_7__5__SCAN_IN, P2_U5123);
  nand ginst14713 (P2_U5144, P2_U2424, P2_U4644);
  nand ginst14714 (P2_U5145, P2_U2416, P2_U4451);
  nand ginst14715 (P2_U5146, P2_U2415, P2_U5113);
  nand ginst14716 (P2_U5147, P2_U2403, P2_U5128);
  nand ginst14717 (P2_U5148, P2_INSTQUEUE_REG_7__4__SCAN_IN, P2_U5123);
  nand ginst14718 (P2_U5149, P2_U2423, P2_U4644);
  nand ginst14719 (P2_U5150, P2_U2414, P2_U4451);
  nand ginst14720 (P2_U5151, P2_U2413, P2_U5113);
  nand ginst14721 (P2_U5152, P2_U2402, P2_U5128);
  nand ginst14722 (P2_U5153, P2_INSTQUEUE_REG_7__3__SCAN_IN, P2_U5123);
  nand ginst14723 (P2_U5154, P2_U2432, P2_U4644);
  nand ginst14724 (P2_U5155, P2_U2412, P2_U4451);
  nand ginst14725 (P2_U5156, P2_U2411, P2_U5113);
  nand ginst14726 (P2_U5157, P2_U2401, P2_U5128);
  nand ginst14727 (P2_U5158, P2_INSTQUEUE_REG_7__2__SCAN_IN, P2_U5123);
  nand ginst14728 (P2_U5159, P2_U2428, P2_U4644);
  nand ginst14729 (P2_U5160, P2_U2410, P2_U4451);
  nand ginst14730 (P2_U5161, P2_U2409, P2_U5113);
  nand ginst14731 (P2_U5162, P2_U2400, P2_U5128);
  nand ginst14732 (P2_U5163, P2_INSTQUEUE_REG_7__1__SCAN_IN, P2_U5123);
  nand ginst14733 (P2_U5164, P2_U2431, P2_U4644);
  nand ginst14734 (P2_U5165, P2_U2408, P2_U4451);
  nand ginst14735 (P2_U5166, P2_U2407, P2_U5113);
  nand ginst14736 (P2_U5167, P2_U2399, P2_U5128);
  nand ginst14737 (P2_U5168, P2_INSTQUEUE_REG_7__0__SCAN_IN, P2_U5123);
  not ginst14738 (P2_U5169, P2_U3440);
  not ginst14739 (P2_U5170, P2_U3439);
  not ginst14740 (P2_U5171, P2_U3249);
  not ginst14741 (P2_U5172, P2_U3561);
  not ginst14742 (P2_U5173, P2_U3441);
  nand ginst14743 (P2_U5174, P2_U2460, P2_U4633);
  nand ginst14744 (P2_U5175, P2_U2362, P2_U2495);
  nand ginst14745 (P2_U5176, P2_U4445, P2_U5175);
  nand ginst14746 (P2_U5177, P2_U3249, P2_U5176);
  nand ginst14747 (P2_U5178, P2_STATE2_REG_2__SCAN_IN, P2_U5173);
  nand ginst14748 (P2_U5179, P2_STATE2_REG_3__SCAN_IN, P2_U3439);
  nand ginst14749 (P2_U5180, P2_U3803, P2_U5177);
  nand ginst14750 (P2_U5181, P2_U2398, P2_U2495);
  nand ginst14751 (P2_U5182, P2_U4445, P2_U5181);
  nand ginst14752 (P2_U5183, P2_U5171, P2_U5182);
  nand ginst14753 (P2_U5184, P2_STATE2_REG_2__SCAN_IN, P2_U3441);
  nand ginst14754 (P2_U5185, P2_U5183, P2_U5184);
  nand ginst14755 (P2_U5186, P2_U2425, P2_U5170);
  nand ginst14756 (P2_U5187, P2_U2422, P2_U2494);
  nand ginst14757 (P2_U5188, P2_U2421, P2_U5169);
  nand ginst14758 (P2_U5189, P2_U2406, P2_U5185);
  nand ginst14759 (P2_U5190, P2_INSTQUEUE_REG_6__7__SCAN_IN, P2_U5180);
  nand ginst14760 (P2_U5191, P2_U2426, P2_U5170);
  nand ginst14761 (P2_U5192, P2_U2420, P2_U2494);
  nand ginst14762 (P2_U5193, P2_U2419, P2_U5169);
  nand ginst14763 (P2_U5194, P2_U2405, P2_U5185);
  nand ginst14764 (P2_U5195, P2_INSTQUEUE_REG_6__6__SCAN_IN, P2_U5180);
  nand ginst14765 (P2_U5196, P2_U2429, P2_U5170);
  nand ginst14766 (P2_U5197, P2_U2418, P2_U2494);
  nand ginst14767 (P2_U5198, P2_U2417, P2_U5169);
  nand ginst14768 (P2_U5199, P2_U2404, P2_U5185);
  nand ginst14769 (P2_U5200, P2_INSTQUEUE_REG_6__5__SCAN_IN, P2_U5180);
  nand ginst14770 (P2_U5201, P2_U2424, P2_U5170);
  nand ginst14771 (P2_U5202, P2_U2416, P2_U2494);
  nand ginst14772 (P2_U5203, P2_U2415, P2_U5169);
  nand ginst14773 (P2_U5204, P2_U2403, P2_U5185);
  nand ginst14774 (P2_U5205, P2_INSTQUEUE_REG_6__4__SCAN_IN, P2_U5180);
  nand ginst14775 (P2_U5206, P2_U2423, P2_U5170);
  nand ginst14776 (P2_U5207, P2_U2414, P2_U2494);
  nand ginst14777 (P2_U5208, P2_U2413, P2_U5169);
  nand ginst14778 (P2_U5209, P2_U2402, P2_U5185);
  nand ginst14779 (P2_U5210, P2_INSTQUEUE_REG_6__3__SCAN_IN, P2_U5180);
  nand ginst14780 (P2_U5211, P2_U2432, P2_U5170);
  nand ginst14781 (P2_U5212, P2_U2412, P2_U2494);
  nand ginst14782 (P2_U5213, P2_U2411, P2_U5169);
  nand ginst14783 (P2_U5214, P2_U2401, P2_U5185);
  nand ginst14784 (P2_U5215, P2_INSTQUEUE_REG_6__2__SCAN_IN, P2_U5180);
  nand ginst14785 (P2_U5216, P2_U2428, P2_U5170);
  nand ginst14786 (P2_U5217, P2_U2410, P2_U2494);
  nand ginst14787 (P2_U5218, P2_U2409, P2_U5169);
  nand ginst14788 (P2_U5219, P2_U2400, P2_U5185);
  nand ginst14789 (P2_U5220, P2_INSTQUEUE_REG_6__1__SCAN_IN, P2_U5180);
  nand ginst14790 (P2_U5221, P2_U2431, P2_U5170);
  nand ginst14791 (P2_U5222, P2_U2408, P2_U2494);
  nand ginst14792 (P2_U5223, P2_U2407, P2_U5169);
  nand ginst14793 (P2_U5224, P2_U2399, P2_U5185);
  nand ginst14794 (P2_U5225, P2_INSTQUEUE_REG_6__0__SCAN_IN, P2_U5180);
  not ginst14795 (P2_U5226, P2_U3451);
  not ginst14796 (P2_U5227, P2_U3450);
  nand ginst14797 (P2_U5228, P2_U2441, P2_U2445);
  not ginst14798 (P2_U5229, P2_U3452);
  not ginst14799 (P2_U5230, P2_U3560);
  not ginst14800 (P2_U5231, P2_U3453);
  nand ginst14801 (P2_U5232, P2_U2460, P2_U4634);
  nand ginst14802 (P2_U5233, P2_U2362, P2_U2497);
  nand ginst14803 (P2_U5234, P2_U4445, P2_U5233);
  nand ginst14804 (P2_U5235, P2_U5229, P2_U5234);
  nand ginst14805 (P2_U5236, P2_STATE2_REG_2__SCAN_IN, P2_U5231);
  nand ginst14806 (P2_U5237, P2_STATE2_REG_3__SCAN_IN, P2_U3450);
  nand ginst14807 (P2_U5238, P2_U3812, P2_U5235);
  nand ginst14808 (P2_U5239, P2_U2398, P2_U2497);
  nand ginst14809 (P2_U5240, P2_U4445, P2_U5239);
  nand ginst14810 (P2_U5241, P2_U3452, P2_U5240);
  nand ginst14811 (P2_U5242, P2_STATE2_REG_2__SCAN_IN, P2_U3453);
  nand ginst14812 (P2_U5243, P2_U5241, P2_U5242);
  nand ginst14813 (P2_U5244, P2_U2425, P2_U5227);
  nand ginst14814 (P2_U5245, P2_U2422, P2_U2496);
  nand ginst14815 (P2_U5246, P2_U2421, P2_U5226);
  nand ginst14816 (P2_U5247, P2_U2406, P2_U5243);
  nand ginst14817 (P2_U5248, P2_INSTQUEUE_REG_5__7__SCAN_IN, P2_U5238);
  nand ginst14818 (P2_U5249, P2_U2426, P2_U5227);
  nand ginst14819 (P2_U5250, P2_U2420, P2_U2496);
  nand ginst14820 (P2_U5251, P2_U2419, P2_U5226);
  nand ginst14821 (P2_U5252, P2_U2405, P2_U5243);
  nand ginst14822 (P2_U5253, P2_INSTQUEUE_REG_5__6__SCAN_IN, P2_U5238);
  nand ginst14823 (P2_U5254, P2_U2429, P2_U5227);
  nand ginst14824 (P2_U5255, P2_U2418, P2_U2496);
  nand ginst14825 (P2_U5256, P2_U2417, P2_U5226);
  nand ginst14826 (P2_U5257, P2_U2404, P2_U5243);
  nand ginst14827 (P2_U5258, P2_INSTQUEUE_REG_5__5__SCAN_IN, P2_U5238);
  nand ginst14828 (P2_U5259, P2_U2424, P2_U5227);
  nand ginst14829 (P2_U5260, P2_U2416, P2_U2496);
  nand ginst14830 (P2_U5261, P2_U2415, P2_U5226);
  nand ginst14831 (P2_U5262, P2_U2403, P2_U5243);
  nand ginst14832 (P2_U5263, P2_INSTQUEUE_REG_5__4__SCAN_IN, P2_U5238);
  nand ginst14833 (P2_U5264, P2_U2423, P2_U5227);
  nand ginst14834 (P2_U5265, P2_U2414, P2_U2496);
  nand ginst14835 (P2_U5266, P2_U2413, P2_U5226);
  nand ginst14836 (P2_U5267, P2_U2402, P2_U5243);
  nand ginst14837 (P2_U5268, P2_INSTQUEUE_REG_5__3__SCAN_IN, P2_U5238);
  nand ginst14838 (P2_U5269, P2_U2432, P2_U5227);
  nand ginst14839 (P2_U5270, P2_U2412, P2_U2496);
  nand ginst14840 (P2_U5271, P2_U2411, P2_U5226);
  nand ginst14841 (P2_U5272, P2_U2401, P2_U5243);
  nand ginst14842 (P2_U5273, P2_INSTQUEUE_REG_5__2__SCAN_IN, P2_U5238);
  nand ginst14843 (P2_U5274, P2_U2428, P2_U5227);
  nand ginst14844 (P2_U5275, P2_U2410, P2_U2496);
  nand ginst14845 (P2_U5276, P2_U2409, P2_U5226);
  nand ginst14846 (P2_U5277, P2_U2400, P2_U5243);
  nand ginst14847 (P2_U5278, P2_INSTQUEUE_REG_5__1__SCAN_IN, P2_U5238);
  nand ginst14848 (P2_U5279, P2_U2431, P2_U5227);
  nand ginst14849 (P2_U5280, P2_U2408, P2_U2496);
  nand ginst14850 (P2_U5281, P2_U2407, P2_U5226);
  nand ginst14851 (P2_U5282, P2_U2399, P2_U5243);
  nand ginst14852 (P2_U5283, P2_INSTQUEUE_REG_5__0__SCAN_IN, P2_U5238);
  not ginst14853 (P2_U5284, P2_U3463);
  not ginst14854 (P2_U5285, P2_U3462);
  not ginst14855 (P2_U5286, P2_U3250);
  not ginst14856 (P2_U5287, P2_U3559);
  not ginst14857 (P2_U5288, P2_U3464);
  nand ginst14858 (P2_U5289, P2_U2460, P2_U2476);
  nand ginst14859 (P2_U5290, P2_U2362, P2_U2499);
  nand ginst14860 (P2_U5291, P2_U4445, P2_U5290);
  nand ginst14861 (P2_U5292, P2_U3250, P2_U5291);
  nand ginst14862 (P2_U5293, P2_STATE2_REG_2__SCAN_IN, P2_U5288);
  nand ginst14863 (P2_U5294, P2_STATE2_REG_3__SCAN_IN, P2_U3462);
  nand ginst14864 (P2_U5295, P2_U3821, P2_U5292);
  nand ginst14865 (P2_U5296, P2_U2398, P2_U2499);
  nand ginst14866 (P2_U5297, P2_U4445, P2_U5296);
  nand ginst14867 (P2_U5298, P2_U5286, P2_U5297);
  nand ginst14868 (P2_U5299, P2_STATE2_REG_2__SCAN_IN, P2_U3464);
  nand ginst14869 (P2_U5300, P2_U5298, P2_U5299);
  nand ginst14870 (P2_U5301, P2_U2425, P2_U5285);
  nand ginst14871 (P2_U5302, P2_U2422, P2_U2498);
  nand ginst14872 (P2_U5303, P2_U2421, P2_U5284);
  nand ginst14873 (P2_U5304, P2_U2406, P2_U5300);
  nand ginst14874 (P2_U5305, P2_INSTQUEUE_REG_4__7__SCAN_IN, P2_U5295);
  nand ginst14875 (P2_U5306, P2_U2426, P2_U5285);
  nand ginst14876 (P2_U5307, P2_U2420, P2_U2498);
  nand ginst14877 (P2_U5308, P2_U2419, P2_U5284);
  nand ginst14878 (P2_U5309, P2_U2405, P2_U5300);
  nand ginst14879 (P2_U5310, P2_INSTQUEUE_REG_4__6__SCAN_IN, P2_U5295);
  nand ginst14880 (P2_U5311, P2_U2429, P2_U5285);
  nand ginst14881 (P2_U5312, P2_U2418, P2_U2498);
  nand ginst14882 (P2_U5313, P2_U2417, P2_U5284);
  nand ginst14883 (P2_U5314, P2_U2404, P2_U5300);
  nand ginst14884 (P2_U5315, P2_INSTQUEUE_REG_4__5__SCAN_IN, P2_U5295);
  nand ginst14885 (P2_U5316, P2_U2424, P2_U5285);
  nand ginst14886 (P2_U5317, P2_U2416, P2_U2498);
  nand ginst14887 (P2_U5318, P2_U2415, P2_U5284);
  nand ginst14888 (P2_U5319, P2_U2403, P2_U5300);
  nand ginst14889 (P2_U5320, P2_INSTQUEUE_REG_4__4__SCAN_IN, P2_U5295);
  nand ginst14890 (P2_U5321, P2_U2423, P2_U5285);
  nand ginst14891 (P2_U5322, P2_U2414, P2_U2498);
  nand ginst14892 (P2_U5323, P2_U2413, P2_U5284);
  nand ginst14893 (P2_U5324, P2_U2402, P2_U5300);
  nand ginst14894 (P2_U5325, P2_INSTQUEUE_REG_4__3__SCAN_IN, P2_U5295);
  nand ginst14895 (P2_U5326, P2_U2432, P2_U5285);
  nand ginst14896 (P2_U5327, P2_U2412, P2_U2498);
  nand ginst14897 (P2_U5328, P2_U2411, P2_U5284);
  nand ginst14898 (P2_U5329, P2_U2401, P2_U5300);
  nand ginst14899 (P2_U5330, P2_INSTQUEUE_REG_4__2__SCAN_IN, P2_U5295);
  nand ginst14900 (P2_U5331, P2_U2428, P2_U5285);
  nand ginst14901 (P2_U5332, P2_U2410, P2_U2498);
  nand ginst14902 (P2_U5333, P2_U2409, P2_U5284);
  nand ginst14903 (P2_U5334, P2_U2400, P2_U5300);
  nand ginst14904 (P2_U5335, P2_INSTQUEUE_REG_4__1__SCAN_IN, P2_U5295);
  nand ginst14905 (P2_U5336, P2_U2431, P2_U5285);
  nand ginst14906 (P2_U5337, P2_U2408, P2_U2498);
  nand ginst14907 (P2_U5338, P2_U2407, P2_U5284);
  nand ginst14908 (P2_U5339, P2_U2399, P2_U5300);
  nand ginst14909 (P2_U5340, P2_INSTQUEUE_REG_4__0__SCAN_IN, P2_U5295);
  not ginst14910 (P2_U5341, P2_U3474);
  not ginst14911 (P2_U5342, P2_U3473);
  nand ginst14912 (P2_U5343, P2_U2443, P2_U2444);
  not ginst14913 (P2_U5344, P2_U3475);
  not ginst14914 (P2_U5345, P2_U3558);
  not ginst14915 (P2_U5346, P2_U3476);
  nand ginst14916 (P2_U5347, P2_U2501, P2_U4637);
  nand ginst14917 (P2_U5348, P2_U2362, P2_U2505);
  nand ginst14918 (P2_U5349, P2_U4445, P2_U5348);
  nand ginst14919 (P2_U5350, P2_U5344, P2_U5349);
  nand ginst14920 (P2_U5351, P2_STATE2_REG_2__SCAN_IN, P2_U5346);
  nand ginst14921 (P2_U5352, P2_STATE2_REG_3__SCAN_IN, P2_U3473);
  nand ginst14922 (P2_U5353, P2_U3830, P2_U5350);
  nand ginst14923 (P2_U5354, P2_U2398, P2_U2505);
  nand ginst14924 (P2_U5355, P2_U4445, P2_U5354);
  nand ginst14925 (P2_U5356, P2_U3475, P2_U5355);
  nand ginst14926 (P2_U5357, P2_STATE2_REG_2__SCAN_IN, P2_U3476);
  nand ginst14927 (P2_U5358, P2_U5356, P2_U5357);
  nand ginst14928 (P2_U5359, P2_U2425, P2_U5342);
  nand ginst14929 (P2_U5360, P2_U2422, P2_U2502);
  nand ginst14930 (P2_U5361, P2_U2421, P2_U5341);
  nand ginst14931 (P2_U5362, P2_U2406, P2_U5358);
  nand ginst14932 (P2_U5363, P2_INSTQUEUE_REG_3__7__SCAN_IN, P2_U5353);
  nand ginst14933 (P2_U5364, P2_U2426, P2_U5342);
  nand ginst14934 (P2_U5365, P2_U2420, P2_U2502);
  nand ginst14935 (P2_U5366, P2_U2419, P2_U5341);
  nand ginst14936 (P2_U5367, P2_U2405, P2_U5358);
  nand ginst14937 (P2_U5368, P2_INSTQUEUE_REG_3__6__SCAN_IN, P2_U5353);
  nand ginst14938 (P2_U5369, P2_U2429, P2_U5342);
  nand ginst14939 (P2_U5370, P2_U2418, P2_U2502);
  nand ginst14940 (P2_U5371, P2_U2417, P2_U5341);
  nand ginst14941 (P2_U5372, P2_U2404, P2_U5358);
  nand ginst14942 (P2_U5373, P2_INSTQUEUE_REG_3__5__SCAN_IN, P2_U5353);
  nand ginst14943 (P2_U5374, P2_U2424, P2_U5342);
  nand ginst14944 (P2_U5375, P2_U2416, P2_U2502);
  nand ginst14945 (P2_U5376, P2_U2415, P2_U5341);
  nand ginst14946 (P2_U5377, P2_U2403, P2_U5358);
  nand ginst14947 (P2_U5378, P2_INSTQUEUE_REG_3__4__SCAN_IN, P2_U5353);
  nand ginst14948 (P2_U5379, P2_U2423, P2_U5342);
  nand ginst14949 (P2_U5380, P2_U2414, P2_U2502);
  nand ginst14950 (P2_U5381, P2_U2413, P2_U5341);
  nand ginst14951 (P2_U5382, P2_U2402, P2_U5358);
  nand ginst14952 (P2_U5383, P2_INSTQUEUE_REG_3__3__SCAN_IN, P2_U5353);
  nand ginst14953 (P2_U5384, P2_U2432, P2_U5342);
  nand ginst14954 (P2_U5385, P2_U2412, P2_U2502);
  nand ginst14955 (P2_U5386, P2_U2411, P2_U5341);
  nand ginst14956 (P2_U5387, P2_U2401, P2_U5358);
  nand ginst14957 (P2_U5388, P2_INSTQUEUE_REG_3__2__SCAN_IN, P2_U5353);
  nand ginst14958 (P2_U5389, P2_U2428, P2_U5342);
  nand ginst14959 (P2_U5390, P2_U2410, P2_U2502);
  nand ginst14960 (P2_U5391, P2_U2409, P2_U5341);
  nand ginst14961 (P2_U5392, P2_U2400, P2_U5358);
  nand ginst14962 (P2_U5393, P2_INSTQUEUE_REG_3__1__SCAN_IN, P2_U5353);
  nand ginst14963 (P2_U5394, P2_U2431, P2_U5342);
  nand ginst14964 (P2_U5395, P2_U2408, P2_U2502);
  nand ginst14965 (P2_U5396, P2_U2407, P2_U5341);
  nand ginst14966 (P2_U5397, P2_U2399, P2_U5358);
  nand ginst14967 (P2_U5398, P2_INSTQUEUE_REG_3__0__SCAN_IN, P2_U5353);
  not ginst14968 (P2_U5399, P2_U3486);
  not ginst14969 (P2_U5400, P2_U3485);
  not ginst14970 (P2_U5401, P2_U3251);
  not ginst14971 (P2_U5402, P2_U3557);
  not ginst14972 (P2_U5403, P2_U3487);
  nand ginst14973 (P2_U5404, P2_U2501, P2_U4633);
  nand ginst14974 (P2_U5405, P2_U2362, P2_U2507);
  nand ginst14975 (P2_U5406, P2_U4445, P2_U5405);
  nand ginst14976 (P2_U5407, P2_U3251, P2_U5406);
  nand ginst14977 (P2_U5408, P2_STATE2_REG_2__SCAN_IN, P2_U5403);
  nand ginst14978 (P2_U5409, P2_STATE2_REG_3__SCAN_IN, P2_U3485);
  nand ginst14979 (P2_U5410, P2_U3839, P2_U5407);
  nand ginst14980 (P2_U5411, P2_U2398, P2_U2507);
  nand ginst14981 (P2_U5412, P2_U4445, P2_U5411);
  nand ginst14982 (P2_U5413, P2_U5401, P2_U5412);
  nand ginst14983 (P2_U5414, P2_STATE2_REG_2__SCAN_IN, P2_U3487);
  nand ginst14984 (P2_U5415, P2_U5413, P2_U5414);
  nand ginst14985 (P2_U5416, P2_U2425, P2_U5400);
  nand ginst14986 (P2_U5417, P2_U2422, P2_U2506);
  nand ginst14987 (P2_U5418, P2_U2421, P2_U5399);
  nand ginst14988 (P2_U5419, P2_U2406, P2_U5415);
  nand ginst14989 (P2_U5420, P2_INSTQUEUE_REG_2__7__SCAN_IN, P2_U5410);
  nand ginst14990 (P2_U5421, P2_U2426, P2_U5400);
  nand ginst14991 (P2_U5422, P2_U2420, P2_U2506);
  nand ginst14992 (P2_U5423, P2_U2419, P2_U5399);
  nand ginst14993 (P2_U5424, P2_U2405, P2_U5415);
  nand ginst14994 (P2_U5425, P2_INSTQUEUE_REG_2__6__SCAN_IN, P2_U5410);
  nand ginst14995 (P2_U5426, P2_U2429, P2_U5400);
  nand ginst14996 (P2_U5427, P2_U2418, P2_U2506);
  nand ginst14997 (P2_U5428, P2_U2417, P2_U5399);
  nand ginst14998 (P2_U5429, P2_U2404, P2_U5415);
  nand ginst14999 (P2_U5430, P2_INSTQUEUE_REG_2__5__SCAN_IN, P2_U5410);
  nand ginst15000 (P2_U5431, P2_U2424, P2_U5400);
  nand ginst15001 (P2_U5432, P2_U2416, P2_U2506);
  nand ginst15002 (P2_U5433, P2_U2415, P2_U5399);
  nand ginst15003 (P2_U5434, P2_U2403, P2_U5415);
  nand ginst15004 (P2_U5435, P2_INSTQUEUE_REG_2__4__SCAN_IN, P2_U5410);
  nand ginst15005 (P2_U5436, P2_U2423, P2_U5400);
  nand ginst15006 (P2_U5437, P2_U2414, P2_U2506);
  nand ginst15007 (P2_U5438, P2_U2413, P2_U5399);
  nand ginst15008 (P2_U5439, P2_U2402, P2_U5415);
  nand ginst15009 (P2_U5440, P2_INSTQUEUE_REG_2__3__SCAN_IN, P2_U5410);
  nand ginst15010 (P2_U5441, P2_U2432, P2_U5400);
  nand ginst15011 (P2_U5442, P2_U2412, P2_U2506);
  nand ginst15012 (P2_U5443, P2_U2411, P2_U5399);
  nand ginst15013 (P2_U5444, P2_U2401, P2_U5415);
  nand ginst15014 (P2_U5445, P2_INSTQUEUE_REG_2__2__SCAN_IN, P2_U5410);
  nand ginst15015 (P2_U5446, P2_U2428, P2_U5400);
  nand ginst15016 (P2_U5447, P2_U2410, P2_U2506);
  nand ginst15017 (P2_U5448, P2_U2409, P2_U5399);
  nand ginst15018 (P2_U5449, P2_U2400, P2_U5415);
  nand ginst15019 (P2_U5450, P2_INSTQUEUE_REG_2__1__SCAN_IN, P2_U5410);
  nand ginst15020 (P2_U5451, P2_U2431, P2_U5400);
  nand ginst15021 (P2_U5452, P2_U2408, P2_U2506);
  nand ginst15022 (P2_U5453, P2_U2407, P2_U5399);
  nand ginst15023 (P2_U5454, P2_U2399, P2_U5415);
  nand ginst15024 (P2_U5455, P2_INSTQUEUE_REG_2__0__SCAN_IN, P2_U5410);
  not ginst15025 (P2_U5456, P2_U3497);
  not ginst15026 (P2_U5457, P2_U3496);
  nand ginst15027 (P2_U5458, P2_U2443, P2_U2445);
  not ginst15028 (P2_U5459, P2_U3498);
  not ginst15029 (P2_U5460, P2_U3556);
  not ginst15030 (P2_U5461, P2_U3499);
  nand ginst15031 (P2_U5462, P2_U2501, P2_U4634);
  nand ginst15032 (P2_U5463, P2_U2362, P2_U2509);
  nand ginst15033 (P2_U5464, P2_U4445, P2_U5463);
  nand ginst15034 (P2_U5465, P2_U5459, P2_U5464);
  nand ginst15035 (P2_U5466, P2_STATE2_REG_2__SCAN_IN, P2_U5461);
  nand ginst15036 (P2_U5467, P2_STATE2_REG_3__SCAN_IN, P2_U3496);
  nand ginst15037 (P2_U5468, P2_U3848, P2_U5465);
  nand ginst15038 (P2_U5469, P2_U2398, P2_U2509);
  nand ginst15039 (P2_U5470, P2_U4445, P2_U5469);
  nand ginst15040 (P2_U5471, P2_U3498, P2_U5470);
  nand ginst15041 (P2_U5472, P2_STATE2_REG_2__SCAN_IN, P2_U3499);
  nand ginst15042 (P2_U5473, P2_U5471, P2_U5472);
  nand ginst15043 (P2_U5474, P2_U2425, P2_U5457);
  nand ginst15044 (P2_U5475, P2_U2422, P2_U2508);
  nand ginst15045 (P2_U5476, P2_U2421, P2_U5456);
  nand ginst15046 (P2_U5477, P2_U2406, P2_U5473);
  nand ginst15047 (P2_U5478, P2_INSTQUEUE_REG_1__7__SCAN_IN, P2_U5468);
  nand ginst15048 (P2_U5479, P2_U2426, P2_U5457);
  nand ginst15049 (P2_U5480, P2_U2420, P2_U2508);
  nand ginst15050 (P2_U5481, P2_U2419, P2_U5456);
  nand ginst15051 (P2_U5482, P2_U2405, P2_U5473);
  nand ginst15052 (P2_U5483, P2_INSTQUEUE_REG_1__6__SCAN_IN, P2_U5468);
  nand ginst15053 (P2_U5484, P2_U2429, P2_U5457);
  nand ginst15054 (P2_U5485, P2_U2418, P2_U2508);
  nand ginst15055 (P2_U5486, P2_U2417, P2_U5456);
  nand ginst15056 (P2_U5487, P2_U2404, P2_U5473);
  nand ginst15057 (P2_U5488, P2_INSTQUEUE_REG_1__5__SCAN_IN, P2_U5468);
  nand ginst15058 (P2_U5489, P2_U2424, P2_U5457);
  nand ginst15059 (P2_U5490, P2_U2416, P2_U2508);
  nand ginst15060 (P2_U5491, P2_U2415, P2_U5456);
  nand ginst15061 (P2_U5492, P2_U2403, P2_U5473);
  nand ginst15062 (P2_U5493, P2_INSTQUEUE_REG_1__4__SCAN_IN, P2_U5468);
  nand ginst15063 (P2_U5494, P2_U2423, P2_U5457);
  nand ginst15064 (P2_U5495, P2_U2414, P2_U2508);
  nand ginst15065 (P2_U5496, P2_U2413, P2_U5456);
  nand ginst15066 (P2_U5497, P2_U2402, P2_U5473);
  nand ginst15067 (P2_U5498, P2_INSTQUEUE_REG_1__3__SCAN_IN, P2_U5468);
  nand ginst15068 (P2_U5499, P2_U2432, P2_U5457);
  nand ginst15069 (P2_U5500, P2_U2412, P2_U2508);
  nand ginst15070 (P2_U5501, P2_U2411, P2_U5456);
  nand ginst15071 (P2_U5502, P2_U2401, P2_U5473);
  nand ginst15072 (P2_U5503, P2_INSTQUEUE_REG_1__2__SCAN_IN, P2_U5468);
  nand ginst15073 (P2_U5504, P2_U2428, P2_U5457);
  nand ginst15074 (P2_U5505, P2_U2410, P2_U2508);
  nand ginst15075 (P2_U5506, P2_U2409, P2_U5456);
  nand ginst15076 (P2_U5507, P2_U2400, P2_U5473);
  nand ginst15077 (P2_U5508, P2_INSTQUEUE_REG_1__1__SCAN_IN, P2_U5468);
  nand ginst15078 (P2_U5509, P2_U2431, P2_U5457);
  nand ginst15079 (P2_U5510, P2_U2408, P2_U2508);
  nand ginst15080 (P2_U5511, P2_U2407, P2_U5456);
  nand ginst15081 (P2_U5512, P2_U2399, P2_U5473);
  nand ginst15082 (P2_U5513, P2_INSTQUEUE_REG_1__0__SCAN_IN, P2_U5468);
  not ginst15083 (P2_U5514, P2_U3509);
  not ginst15084 (P2_U5515, P2_U3508);
  not ginst15085 (P2_U5516, P2_U3252);
  not ginst15086 (P2_U5517, P2_U3555);
  not ginst15087 (P2_U5518, P2_U3510);
  nand ginst15088 (P2_U5519, P2_U2476, P2_U2501);
  nand ginst15089 (P2_U5520, P2_U2362, P2_U2511);
  nand ginst15090 (P2_U5521, P2_U4445, P2_U5520);
  nand ginst15091 (P2_U5522, P2_U3252, P2_U5521);
  nand ginst15092 (P2_U5523, P2_STATE2_REG_2__SCAN_IN, P2_U5518);
  nand ginst15093 (P2_U5524, P2_STATE2_REG_3__SCAN_IN, P2_U3508);
  nand ginst15094 (P2_U5525, P2_U3857, P2_U5522);
  nand ginst15095 (P2_U5526, P2_U2398, P2_U2511);
  nand ginst15096 (P2_U5527, P2_U4445, P2_U5526);
  nand ginst15097 (P2_U5528, P2_U5516, P2_U5527);
  nand ginst15098 (P2_U5529, P2_STATE2_REG_2__SCAN_IN, P2_U3510);
  nand ginst15099 (P2_U5530, P2_U5528, P2_U5529);
  nand ginst15100 (P2_U5531, P2_U2425, P2_U5515);
  nand ginst15101 (P2_U5532, P2_U2422, P2_U2510);
  nand ginst15102 (P2_U5533, P2_U2421, P2_U5514);
  nand ginst15103 (P2_U5534, P2_U2406, P2_U5530);
  nand ginst15104 (P2_U5535, P2_INSTQUEUE_REG_0__7__SCAN_IN, P2_U5525);
  nand ginst15105 (P2_U5536, P2_U2426, P2_U5515);
  nand ginst15106 (P2_U5537, P2_U2420, P2_U2510);
  nand ginst15107 (P2_U5538, P2_U2419, P2_U5514);
  nand ginst15108 (P2_U5539, P2_U2405, P2_U5530);
  nand ginst15109 (P2_U5540, P2_INSTQUEUE_REG_0__6__SCAN_IN, P2_U5525);
  nand ginst15110 (P2_U5541, P2_U2429, P2_U5515);
  nand ginst15111 (P2_U5542, P2_U2418, P2_U2510);
  nand ginst15112 (P2_U5543, P2_U2417, P2_U5514);
  nand ginst15113 (P2_U5544, P2_U2404, P2_U5530);
  nand ginst15114 (P2_U5545, P2_INSTQUEUE_REG_0__5__SCAN_IN, P2_U5525);
  nand ginst15115 (P2_U5546, P2_U2424, P2_U5515);
  nand ginst15116 (P2_U5547, P2_U2416, P2_U2510);
  nand ginst15117 (P2_U5548, P2_U2415, P2_U5514);
  nand ginst15118 (P2_U5549, P2_U2403, P2_U5530);
  nand ginst15119 (P2_U5550, P2_INSTQUEUE_REG_0__4__SCAN_IN, P2_U5525);
  nand ginst15120 (P2_U5551, P2_U2423, P2_U5515);
  nand ginst15121 (P2_U5552, P2_U2414, P2_U2510);
  nand ginst15122 (P2_U5553, P2_U2413, P2_U5514);
  nand ginst15123 (P2_U5554, P2_U2402, P2_U5530);
  nand ginst15124 (P2_U5555, P2_INSTQUEUE_REG_0__3__SCAN_IN, P2_U5525);
  nand ginst15125 (P2_U5556, P2_U2432, P2_U5515);
  nand ginst15126 (P2_U5557, P2_U2412, P2_U2510);
  nand ginst15127 (P2_U5558, P2_U2411, P2_U5514);
  nand ginst15128 (P2_U5559, P2_U2401, P2_U5530);
  nand ginst15129 (P2_U5560, P2_INSTQUEUE_REG_0__2__SCAN_IN, P2_U5525);
  nand ginst15130 (P2_U5561, P2_U2428, P2_U5515);
  nand ginst15131 (P2_U5562, P2_U2410, P2_U2510);
  nand ginst15132 (P2_U5563, P2_U2409, P2_U5514);
  nand ginst15133 (P2_U5564, P2_U2400, P2_U5530);
  nand ginst15134 (P2_U5565, P2_INSTQUEUE_REG_0__1__SCAN_IN, P2_U5525);
  nand ginst15135 (P2_U5566, P2_U2431, P2_U5515);
  nand ginst15136 (P2_U5567, P2_U2408, P2_U2510);
  nand ginst15137 (P2_U5568, P2_U2407, P2_U5514);
  nand ginst15138 (P2_U5569, P2_U2399, P2_U5530);
  nand ginst15139 (P2_U5570, P2_INSTQUEUE_REG_0__0__SCAN_IN, P2_U5525);
  nand ginst15140 (P2_U5571, P2_U3279, P2_U7869);
  not ginst15141 (P2_U5572, P2_U3574);
  nand ginst15142 (P2_U5573, P2_U2617, P2_U7861, P2_U7863);
  nand ginst15143 (P2_U5574, P2_U3255, P2_U3289, P2_U3521, P2_U7895);
  nand ginst15144 (P2_U5575, P2_U2357, P2_U7871);
  nand ginst15145 (P2_U5576, P2_U3574, P2_U4417);
  nand ginst15146 (P2_U5577, P2_U4424, P2_U4428);
  nand ginst15147 (P2_U5578, P2_U3524, P2_U5577);
  nand ginst15148 (P2_U5579, P2_R2088_U6, P2_U3265, P2_U5578);
  nand ginst15149 (P2_U5580, P2_R2167_U6, P2_U4436);
  not ginst15150 (P2_U5581, P2_U4406);
  nand ginst15151 (P2_U5582, P2_U2374, P2_U4406);
  nand ginst15152 (P2_U5583, P2_STATE2_REG_3__SCAN_IN, P2_U3284);
  not ginst15153 (P2_U5584, P2_U4394);
  nand ginst15154 (P2_U5585, P2_U3276, P2_U4591);
  nand ginst15155 (P2_U5586, P2_U2617, P2_U3295, P2_U3878);
  nand ginst15156 (P2_U5587, P2_U3255, P2_U3295);
  nand ginst15157 (P2_U5588, P2_U3278, P2_U7865);
  nand ginst15158 (P2_U5589, P2_U3879, P2_U8074, P2_U8075);
  not ginst15159 (P2_U5590, P2_U3525);
  nand ginst15160 (P2_U5591, P2_U3278, P2_U7738);
  nand ginst15161 (P2_U5592, P2_U3521, P2_U5571, P2_U5573, P2_U5591);
  nand ginst15162 (P2_U5593, P2_U3574, P2_U4417);
  nand ginst15163 (P2_U5594, P2_U2616, P2_U5592);
  nand ginst15164 (P2_U5595, P2_U3877, P2_U5594);
  nand ginst15165 (P2_U5596, P2_U3295, P2_U7873);
  nand ginst15166 (P2_U5597, P2_U3279, P2_U7871);
  nand ginst15167 (P2_U5598, P2_U2617, P2_U3521);
  nand ginst15168 (P2_U5599, P2_U4427, P2_U5598);
  nand ginst15169 (P2_U5600, P2_U3280, P2_U5597);
  nand ginst15170 (P2_U5601, P2_U2436, P2_U7884);
  nand ginst15171 (P2_U5602, P2_U3278, P2_U3527);
  nand ginst15172 (P2_U5603, P2_U2514, P2_U3288);
  nand ginst15173 (P2_U5604, P2_U4470, P2_U8076, P2_U8077);
  nand ginst15174 (P2_U5605, P2_U3296, P2_U3522);
  nand ginst15175 (P2_U5606, P2_U3578, P2_U4437);
  nand ginst15176 (P2_U5607, P2_U4395, P2_U5605);
  nand ginst15177 (P2_U5608, P2_U3581, P2_U5606);
  nand ginst15178 (P2_U5609, P2_R2147_U8, P2_U5604);
  nand ginst15179 (P2_U5610, P2_R2099_U95, P2_U5603);
  nand ginst15180 (P2_U5611, P2_U3884, P2_U5610);
  nand ginst15181 (P2_U5612, P2_R2182_U76, P2_U4469);
  nand ginst15182 (P2_U5613, P2_U4466, P2_U5611);
  nand ginst15183 (P2_U5614, P2_U5612, P2_U5613);
  nand ginst15184 (P2_U5615, P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN, P2_U4591);
  not ginst15185 (P2_U5616, P2_U3530);
  nand ginst15186 (P2_U5617, P2_R2147_U9, P2_U5604);
  nand ginst15187 (P2_U5618, P2_R2099_U96, P2_U5603);
  nand ginst15188 (P2_U5619, P2_U3885, P2_U5618);
  nand ginst15189 (P2_U5620, P2_STATE2_REG_1__SCAN_IN, P2_U3597, P2_U3598);
  nand ginst15190 (P2_U5621, P2_R2182_U40, P2_U4469);
  nand ginst15191 (P2_U5622, P2_U4466, P2_U5619);
  nand ginst15192 (P2_U5623, P2_U5620, P2_U5621, P2_U5622);
  nand ginst15193 (P2_U5624, P2_U2449, P2_U4429, P2_U7861);
  nand ginst15194 (P2_U5625, P2_U5624, P2_U7882);
  nand ginst15195 (P2_U5626, P2_U3887, P2_U8097);
  nand ginst15196 (P2_U5627, P2_R2147_U4, P2_U5604);
  nand ginst15197 (P2_U5628, P2_R2099_U5, P2_U5603);
  nand ginst15198 (P2_U5629, P2_U3888, P2_U5628);
  nand ginst15199 (P2_U5630, P2_STATE2_REG_1__SCAN_IN, P2_U3597, P2_U8090);
  nand ginst15200 (P2_U5631, P2_R2182_U68, P2_U4469);
  nand ginst15201 (P2_U5632, P2_U4466, P2_U5629);
  nand ginst15202 (P2_U5633, P2_U5630, P2_U5631, P2_U5632);
  nand ginst15203 (P2_U5634, P2_U3889, P2_U8097);
  nand ginst15204 (P2_U5635, P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN, P2_U5604);
  nand ginst15205 (P2_U5636, P2_R2099_U94, P2_U5603);
  nand ginst15206 (P2_U5637, P2_U3890, P2_U5636);
  nand ginst15207 (P2_U5638, P2_R2182_U69, P2_U4469);
  nand ginst15208 (P2_U5639, P2_U4466, P2_U5637);
  nand ginst15209 (P2_U5640, P2_STATE2_REG_1__SCAN_IN, P2_U8087);
  nand ginst15210 (P2_U5641, P2_U5638, P2_U5639, P2_U5640);
  nand ginst15211 (P2_U5642, P2_STATE2_REG_0__SCAN_IN, P2_R2243_U8, P2_U2448);
  not ginst15212 (P2_U5643, P2_U3533);
  nand ginst15213 (P2_U5644, P2_U3303, P2_U4445);
  nand ginst15214 (P2_U5645, P2_U3579, P2_U4636);
  nand ginst15215 (P2_U5646, P2_U3426, P2_U5645);
  nand ginst15216 (P2_U5647, P2_U3427, P2_U5646);
  nand ginst15217 (P2_U5648, P2_U2398, P2_U5647);
  nand ginst15218 (P2_U5649, P2_R2182_U76, P2_U5644);
  nand ginst15219 (P2_U5650, P2_STATE2_REG_3__SCAN_IN, P2_R2096_U75);
  nand ginst15220 (P2_U5651, P2_U3891, P2_U5648);
  nand ginst15221 (P2_U5652, P2_U2398, P2_U8109);
  nand ginst15222 (P2_U5653, P2_R2182_U40, P2_U5644);
  nand ginst15223 (P2_U5654, P2_STATE2_REG_3__SCAN_IN, P2_R2096_U77);
  nand ginst15224 (P2_U5655, P2_U3892, P2_U5652);
  nand ginst15225 (P2_U5656, P2_U3338, P2_U3353);
  nand ginst15226 (P2_U5657, P2_U2398, P2_U5656);
  nand ginst15227 (P2_U5658, P2_R2182_U68, P2_U5644);
  nand ginst15228 (P2_U5659, P2_STATE2_REG_3__SCAN_IN, P2_R2096_U51);
  nand ginst15229 (P2_U5660, P2_U3893, P2_U5657);
  nand ginst15230 (P2_U5661, P2_U3303, P2_U3313);
  nand ginst15231 (P2_U5662, P2_R2182_U69, P2_U5661);
  nand ginst15232 (P2_U5663, P2_STATE2_REG_3__SCAN_IN, P2_R2096_U68);
  nand ginst15233 (P2_U5664, P2_U4464, P2_U5662, P2_U5663);
  nand ginst15234 (P2_U5665, P2_U2616, P2_U3292);
  nand ginst15235 (P2_U5666, P2_GTE_370_U6, P2_U4417);
  nand ginst15236 (P2_U5667, P2_U5665, P2_U5666);
  nand ginst15237 (P2_U5668, P2_R2088_U6, P2_U3265, P2_U8121, P2_U8122);
  nand ginst15238 (P2_U5669, P2_U4420, P2_U5667);
  nand ginst15239 (P2_U5670, P2_U2512, P2_U3894, P2_U4397, P2_U5669);
  nand ginst15240 (P2_U5671, P2_U2374, P2_U5670);
  nand ginst15241 (P2_U5672, P2_U3284, P2_U4461);
  not ginst15242 (P2_U5673, P2_U3535);
  nand ginst15243 (P2_U5674, P2_U4420, P2_U4427);
  nand ginst15244 (P2_U5675, P2_U2514, P2_U3895);
  nand ginst15245 (P2_U5676, P2_U4417, P2_U4424);
  nand ginst15246 (P2_U5677, P2_U3524, P2_U4437, P2_U4470, P2_U5676);
  nand ginst15247 (P2_U5678, P2_U4424, P2_U4428);
  nand ginst15248 (P2_U5679, P2_U3296, P2_U3523, P2_U5678);
  nand ginst15249 (P2_U5680, P2_R2096_U68, P2_U2390);
  nand ginst15250 (P2_U5681, P2_R2099_U94, P2_U2389);
  nand ginst15251 (P2_U5682, P2_R2027_U5, P2_U2388);
  nand ginst15252 (P2_U5683, P2_ADD_394_U4, P2_U2386);
  nand ginst15253 (P2_U5684, P2_R2278_U83, P2_U2385);
  nand ginst15254 (P2_U5685, P2_ADD_371_1212_U68, P2_U2384);
  nand ginst15255 (P2_U5686, P2_REIP_REG_0__SCAN_IN, P2_U2381);
  nand ginst15256 (P2_U5687, P2_INSTADDRPOINTER_REG_0__SCAN_IN, P2_U5673);
  nand ginst15257 (P2_U5688, P2_R2096_U51, P2_U2390);
  nand ginst15258 (P2_U5689, P2_R2099_U5, P2_U2389);
  nand ginst15259 (P2_U5690, P2_R2027_U85, P2_U2388);
  nand ginst15260 (P2_U5691, P2_ADD_394_U85, P2_U2386);
  nand ginst15261 (P2_U5692, P2_R2278_U6, P2_U2385);
  nand ginst15262 (P2_U5693, P2_ADD_371_1212_U25, P2_U2384);
  nand ginst15263 (P2_U5694, P2_REIP_REG_1__SCAN_IN, P2_U2381);
  nand ginst15264 (P2_U5695, P2_INSTADDRPOINTER_REG_1__SCAN_IN, P2_U5673);
  nand ginst15265 (P2_U5696, P2_R2096_U77, P2_U2390);
  nand ginst15266 (P2_U5697, P2_R2099_U96, P2_U2389);
  nand ginst15267 (P2_U5698, P2_R2027_U74, P2_U2388);
  nand ginst15268 (P2_U5699, P2_ADD_394_U5, P2_U2386);
  nand ginst15269 (P2_U5700, P2_R2278_U92, P2_U2385);
  nand ginst15270 (P2_U5701, P2_ADD_371_1212_U79, P2_U2384);
  nand ginst15271 (P2_U5702, P2_REIP_REG_2__SCAN_IN, P2_U2381);
  nand ginst15272 (P2_U5703, P2_INSTADDRPOINTER_REG_2__SCAN_IN, P2_U5673);
  nand ginst15273 (P2_U5704, P2_R2096_U75, P2_U2390);
  nand ginst15274 (P2_U5705, P2_R2099_U95, P2_U2389);
  nand ginst15275 (P2_U5706, P2_R2027_U71, P2_U2388);
  nand ginst15276 (P2_U5707, P2_ADD_394_U95, P2_U2386);
  nand ginst15277 (P2_U5708, P2_R2278_U90, P2_U2385);
  nand ginst15278 (P2_U5709, P2_ADD_371_1212_U84, P2_U2384);
  nand ginst15279 (P2_U5710, P2_REIP_REG_3__SCAN_IN, P2_U2381);
  nand ginst15280 (P2_U5711, P2_INSTADDRPOINTER_REG_3__SCAN_IN, P2_U5673);
  nand ginst15281 (P2_U5712, P2_R2096_U74, P2_U2390);
  nand ginst15282 (P2_U5713, P2_R2099_U98, P2_U2389);
  nand ginst15283 (P2_U5714, P2_R2027_U70, P2_U2388);
  nand ginst15284 (P2_U5715, P2_ADD_394_U76, P2_U2386);
  nand ginst15285 (P2_U5716, P2_R2278_U89, P2_U2385);
  nand ginst15286 (P2_U5717, P2_ADD_371_1212_U80, P2_U2384);
  nand ginst15287 (P2_U5718, P2_REIP_REG_4__SCAN_IN, P2_U2381);
  nand ginst15288 (P2_U5719, P2_INSTADDRPOINTER_REG_4__SCAN_IN, P2_U5673);
  nand ginst15289 (P2_U5720, P2_R2096_U73, P2_U2390);
  nand ginst15290 (P2_U5721, P2_R2099_U71, P2_U2389);
  nand ginst15291 (P2_U5722, P2_R2027_U69, P2_U2388);
  nand ginst15292 (P2_U5723, P2_ADD_394_U79, P2_U2386);
  nand ginst15293 (P2_U5724, P2_R2278_U88, P2_U2385);
  nand ginst15294 (P2_U5725, P2_ADD_371_1212_U81, P2_U2384);
  nand ginst15295 (P2_U5726, P2_REIP_REG_5__SCAN_IN, P2_U2381);
  nand ginst15296 (P2_U5727, P2_INSTADDRPOINTER_REG_5__SCAN_IN, P2_U5673);
  nand ginst15297 (P2_U5728, P2_R2096_U72, P2_U2390);
  nand ginst15298 (P2_U5729, P2_R2099_U70, P2_U2389);
  nand ginst15299 (P2_U5730, P2_R2027_U68, P2_U2388);
  nand ginst15300 (P2_U5731, P2_ADD_394_U63, P2_U2386);
  nand ginst15301 (P2_U5732, P2_R2278_U87, P2_U2385);
  nand ginst15302 (P2_U5733, P2_ADD_371_1212_U78, P2_U2384);
  nand ginst15303 (P2_U5734, P2_REIP_REG_6__SCAN_IN, P2_U2381);
  nand ginst15304 (P2_U5735, P2_INSTADDRPOINTER_REG_6__SCAN_IN, P2_U5673);
  nand ginst15305 (P2_U5736, P2_R2096_U71, P2_U2390);
  nand ginst15306 (P2_U5737, P2_R2099_U69, P2_U2389);
  nand ginst15307 (P2_U5738, P2_R2027_U67, P2_U2388);
  nand ginst15308 (P2_U5739, P2_ADD_394_U89, P2_U2386);
  nand ginst15309 (P2_U5740, P2_R2278_U86, P2_U2385);
  nand ginst15310 (P2_U5741, P2_ADD_371_1212_U85, P2_U2384);
  nand ginst15311 (P2_U5742, P2_REIP_REG_7__SCAN_IN, P2_U2381);
  nand ginst15312 (P2_U5743, P2_INSTADDRPOINTER_REG_7__SCAN_IN, P2_U5673);
  nand ginst15313 (P2_U5744, P2_R2096_U70, P2_U2390);
  nand ginst15314 (P2_U5745, P2_R2099_U68, P2_U2389);
  nand ginst15315 (P2_U5746, P2_R2027_U66, P2_U2388);
  nand ginst15316 (P2_U5747, P2_ADD_394_U80, P2_U2386);
  nand ginst15317 (P2_U5748, P2_R2278_U85, P2_U2385);
  nand ginst15318 (P2_U5749, P2_ADD_371_1212_U82, P2_U2384);
  nand ginst15319 (P2_U5750, P2_REIP_REG_8__SCAN_IN, P2_U2381);
  nand ginst15320 (P2_U5751, P2_INSTADDRPOINTER_REG_8__SCAN_IN, P2_U5673);
  nand ginst15321 (P2_U5752, P2_R2096_U69, P2_U2390);
  nand ginst15322 (P2_U5753, P2_R2099_U67, P2_U2389);
  nand ginst15323 (P2_U5754, P2_R2027_U65, P2_U2388);
  nand ginst15324 (P2_U5755, P2_ADD_394_U70, P2_U2386);
  nand ginst15325 (P2_U5756, P2_R2278_U84, P2_U2385);
  nand ginst15326 (P2_U5757, P2_ADD_371_1212_U118, P2_U2384);
  nand ginst15327 (P2_U5758, P2_REIP_REG_9__SCAN_IN, P2_U2381);
  nand ginst15328 (P2_U5759, P2_INSTADDRPOINTER_REG_9__SCAN_IN, P2_U5673);
  nand ginst15329 (P2_U5760, P2_R2096_U97, P2_U2390);
  nand ginst15330 (P2_U5761, P2_R2099_U93, P2_U2389);
  nand ginst15331 (P2_U5762, P2_R2027_U95, P2_U2388);
  nand ginst15332 (P2_U5763, P2_ADD_394_U83, P2_U2386);
  nand ginst15333 (P2_U5764, P2_R2278_U112, P2_U2385);
  nand ginst15334 (P2_U5765, P2_ADD_371_1212_U13, P2_U2384);
  nand ginst15335 (P2_U5766, P2_REIP_REG_10__SCAN_IN, P2_U2381);
  nand ginst15336 (P2_U5767, P2_INSTADDRPOINTER_REG_10__SCAN_IN, P2_U5673);
  nand ginst15337 (P2_U5768, P2_R2096_U96, P2_U2390);
  nand ginst15338 (P2_U5769, P2_R2099_U92, P2_U2389);
  nand ginst15339 (P2_U5770, P2_R2027_U94, P2_U2388);
  nand ginst15340 (P2_U5771, P2_ADD_394_U73, P2_U2386);
  nand ginst15341 (P2_U5772, P2_R2278_U111, P2_U2385);
  nand ginst15342 (P2_U5773, P2_ADD_371_1212_U14, P2_U2384);
  nand ginst15343 (P2_U5774, P2_REIP_REG_11__SCAN_IN, P2_U2381);
  nand ginst15344 (P2_U5775, P2_INSTADDRPOINTER_REG_11__SCAN_IN, P2_U5673);
  nand ginst15345 (P2_U5776, P2_R2096_U95, P2_U2390);
  nand ginst15346 (P2_U5777, P2_R2099_U91, P2_U2389);
  nand ginst15347 (P2_U5778, P2_R2027_U93, P2_U2388);
  nand ginst15348 (P2_U5779, P2_ADD_394_U88, P2_U2386);
  nand ginst15349 (P2_U5780, P2_R2278_U110, P2_U2385);
  nand ginst15350 (P2_U5781, P2_ADD_371_1212_U76, P2_U2384);
  nand ginst15351 (P2_U5782, P2_REIP_REG_12__SCAN_IN, P2_U2381);
  nand ginst15352 (P2_U5783, P2_INSTADDRPOINTER_REG_12__SCAN_IN, P2_U5673);
  nand ginst15353 (P2_U5784, P2_R2096_U94, P2_U2390);
  nand ginst15354 (P2_U5785, P2_R2099_U90, P2_U2389);
  nand ginst15355 (P2_U5786, P2_R2027_U92, P2_U2388);
  nand ginst15356 (P2_U5787, P2_ADD_394_U69, P2_U2386);
  nand ginst15357 (P2_U5788, P2_R2278_U109, P2_U2385);
  nand ginst15358 (P2_U5789, P2_ADD_371_1212_U15, P2_U2384);
  nand ginst15359 (P2_U5790, P2_REIP_REG_13__SCAN_IN, P2_U2381);
  nand ginst15360 (P2_U5791, P2_INSTADDRPOINTER_REG_13__SCAN_IN, P2_U5673);
  nand ginst15361 (P2_U5792, P2_R2096_U93, P2_U2390);
  nand ginst15362 (P2_U5793, P2_R2099_U89, P2_U2389);
  nand ginst15363 (P2_U5794, P2_R2027_U91, P2_U2388);
  nand ginst15364 (P2_U5795, P2_ADD_394_U78, P2_U2386);
  nand ginst15365 (P2_U5796, P2_R2278_U108, P2_U2385);
  nand ginst15366 (P2_U5797, P2_ADD_371_1212_U16, P2_U2384);
  nand ginst15367 (P2_U5798, P2_REIP_REG_14__SCAN_IN, P2_U2381);
  nand ginst15368 (P2_U5799, P2_INSTADDRPOINTER_REG_14__SCAN_IN, P2_U5673);
  nand ginst15369 (P2_U5800, P2_R2096_U92, P2_U2390);
  nand ginst15370 (P2_U5801, P2_R2099_U88, P2_U2389);
  nand ginst15371 (P2_U5802, P2_R2027_U90, P2_U2388);
  nand ginst15372 (P2_U5803, P2_ADD_394_U75, P2_U2386);
  nand ginst15373 (P2_U5804, P2_R2278_U107, P2_U2385);
  nand ginst15374 (P2_U5805, P2_ADD_371_1212_U73, P2_U2384);
  nand ginst15375 (P2_U5806, P2_REIP_REG_15__SCAN_IN, P2_U2381);
  nand ginst15376 (P2_U5807, P2_INSTADDRPOINTER_REG_15__SCAN_IN, P2_U5673);
  nand ginst15377 (P2_U5808, P2_R2096_U91, P2_U2390);
  nand ginst15378 (P2_U5809, P2_R2099_U87, P2_U2389);
  nand ginst15379 (P2_U5810, P2_R2027_U89, P2_U2388);
  nand ginst15380 (P2_U5811, P2_ADD_394_U91, P2_U2386);
  nand ginst15381 (P2_U5812, P2_R2278_U106, P2_U2385);
  nand ginst15382 (P2_U5813, P2_ADD_371_1212_U17, P2_U2384);
  nand ginst15383 (P2_U5814, P2_REIP_REG_16__SCAN_IN, P2_U2381);
  nand ginst15384 (P2_U5815, P2_INSTADDRPOINTER_REG_16__SCAN_IN, P2_U5673);
  nand ginst15385 (P2_U5816, P2_R2096_U90, P2_U2390);
  nand ginst15386 (P2_U5817, P2_R2099_U86, P2_U2389);
  nand ginst15387 (P2_U5818, P2_R2027_U88, P2_U2388);
  nand ginst15388 (P2_U5819, P2_ADD_394_U67, P2_U2386);
  nand ginst15389 (P2_U5820, P2_R2278_U105, P2_U2385);
  nand ginst15390 (P2_U5821, P2_ADD_371_1212_U71, P2_U2384);
  nand ginst15391 (P2_U5822, P2_REIP_REG_17__SCAN_IN, P2_U2381);
  nand ginst15392 (P2_U5823, P2_INSTADDRPOINTER_REG_17__SCAN_IN, P2_U5673);
  nand ginst15393 (P2_U5824, P2_R2096_U89, P2_U2390);
  nand ginst15394 (P2_U5825, P2_R2099_U85, P2_U2389);
  nand ginst15395 (P2_U5826, P2_R2027_U87, P2_U2388);
  nand ginst15396 (P2_U5827, P2_ADD_394_U72, P2_U2386);
  nand ginst15397 (P2_U5828, P2_R2278_U104, P2_U2385);
  nand ginst15398 (P2_U5829, P2_ADD_371_1212_U72, P2_U2384);
  nand ginst15399 (P2_U5830, P2_REIP_REG_18__SCAN_IN, P2_U2381);
  nand ginst15400 (P2_U5831, P2_INSTADDRPOINTER_REG_18__SCAN_IN, P2_U5673);
  nand ginst15401 (P2_U5832, P2_R2096_U88, P2_U2390);
  nand ginst15402 (P2_U5833, P2_R2099_U84, P2_U2389);
  nand ginst15403 (P2_U5834, P2_R2027_U86, P2_U2388);
  nand ginst15404 (P2_U5835, P2_ADD_394_U82, P2_U2386);
  nand ginst15405 (P2_U5836, P2_R2278_U103, P2_U2385);
  nand ginst15406 (P2_U5837, P2_ADD_371_1212_U18, P2_U2384);
  nand ginst15407 (P2_U5838, P2_REIP_REG_19__SCAN_IN, P2_U2381);
  nand ginst15408 (P2_U5839, P2_INSTADDRPOINTER_REG_19__SCAN_IN, P2_U5673);
  nand ginst15409 (P2_U5840, P2_R2096_U87, P2_U2390);
  nand ginst15410 (P2_U5841, P2_R2099_U83, P2_U2389);
  nand ginst15411 (P2_U5842, P2_R2027_U84, P2_U2388);
  nand ginst15412 (P2_U5843, P2_ADD_394_U68, P2_U2386);
  nand ginst15413 (P2_U5844, P2_R2278_U102, P2_U2385);
  nand ginst15414 (P2_U5845, P2_ADD_371_1212_U19, P2_U2384);
  nand ginst15415 (P2_U5846, P2_REIP_REG_20__SCAN_IN, P2_U2381);
  nand ginst15416 (P2_U5847, P2_INSTADDRPOINTER_REG_20__SCAN_IN, P2_U5673);
  nand ginst15417 (P2_U5848, P2_R2096_U86, P2_U2390);
  nand ginst15418 (P2_U5849, P2_R2099_U82, P2_U2389);
  nand ginst15419 (P2_U5850, P2_R2027_U83, P2_U2388);
  nand ginst15420 (P2_U5851, P2_ADD_394_U87, P2_U2386);
  nand ginst15421 (P2_U5852, P2_R2278_U101, P2_U2385);
  nand ginst15422 (P2_U5853, P2_ADD_371_1212_U75, P2_U2384);
  nand ginst15423 (P2_U5854, P2_REIP_REG_21__SCAN_IN, P2_U2381);
  nand ginst15424 (P2_U5855, P2_INSTADDRPOINTER_REG_21__SCAN_IN, P2_U5673);
  nand ginst15425 (P2_U5856, P2_R2096_U85, P2_U2390);
  nand ginst15426 (P2_U5857, P2_R2099_U81, P2_U2389);
  nand ginst15427 (P2_U5858, P2_R2027_U82, P2_U2388);
  nand ginst15428 (P2_U5859, P2_ADD_394_U71, P2_U2386);
  nand ginst15429 (P2_U5860, P2_R2278_U100, P2_U2385);
  nand ginst15430 (P2_U5861, P2_ADD_371_1212_U20, P2_U2384);
  nand ginst15431 (P2_U5862, P2_REIP_REG_22__SCAN_IN, P2_U2381);
  nand ginst15432 (P2_U5863, P2_INSTADDRPOINTER_REG_22__SCAN_IN, P2_U5673);
  nand ginst15433 (P2_U5864, P2_R2096_U84, P2_U2390);
  nand ginst15434 (P2_U5865, P2_R2099_U80, P2_U2389);
  nand ginst15435 (P2_U5866, P2_R2027_U81, P2_U2388);
  nand ginst15436 (P2_U5867, P2_ADD_394_U81, P2_U2386);
  nand ginst15437 (P2_U5868, P2_R2278_U99, P2_U2385);
  nand ginst15438 (P2_U5869, P2_ADD_371_1212_U21, P2_U2384);
  nand ginst15439 (P2_U5870, P2_REIP_REG_23__SCAN_IN, P2_U2381);
  nand ginst15440 (P2_U5871, P2_INSTADDRPOINTER_REG_23__SCAN_IN, P2_U5673);
  nand ginst15441 (P2_U5872, P2_R2096_U83, P2_U2390);
  nand ginst15442 (P2_U5873, P2_R2099_U79, P2_U2389);
  nand ginst15443 (P2_U5874, P2_R2027_U80, P2_U2388);
  nand ginst15444 (P2_U5875, P2_ADD_394_U66, P2_U2386);
  nand ginst15445 (P2_U5876, P2_R2278_U98, P2_U2385);
  nand ginst15446 (P2_U5877, P2_ADD_371_1212_U70, P2_U2384);
  nand ginst15447 (P2_U5878, P2_REIP_REG_24__SCAN_IN, P2_U2381);
  nand ginst15448 (P2_U5879, P2_INSTADDRPOINTER_REG_24__SCAN_IN, P2_U5673);
  nand ginst15449 (P2_U5880, P2_R2096_U82, P2_U2390);
  nand ginst15450 (P2_U5881, P2_R2099_U78, P2_U2389);
  nand ginst15451 (P2_U5882, P2_R2027_U79, P2_U2388);
  nand ginst15452 (P2_U5883, P2_ADD_394_U90, P2_U2386);
  nand ginst15453 (P2_U5884, P2_R2278_U97, P2_U2385);
  nand ginst15454 (P2_U5885, P2_ADD_371_1212_U77, P2_U2384);
  nand ginst15455 (P2_U5886, P2_REIP_REG_25__SCAN_IN, P2_U2381);
  nand ginst15456 (P2_U5887, P2_INSTADDRPOINTER_REG_25__SCAN_IN, P2_U5673);
  nand ginst15457 (P2_U5888, P2_R2096_U81, P2_U2390);
  nand ginst15458 (P2_U5889, P2_R2099_U77, P2_U2389);
  nand ginst15459 (P2_U5890, P2_R2027_U78, P2_U2388);
  nand ginst15460 (P2_U5891, P2_ADD_394_U74, P2_U2386);
  nand ginst15461 (P2_U5892, P2_R2278_U96, P2_U2385);
  nand ginst15462 (P2_U5893, P2_ADD_371_1212_U22, P2_U2384);
  nand ginst15463 (P2_U5894, P2_REIP_REG_26__SCAN_IN, P2_U2381);
  nand ginst15464 (P2_U5895, P2_INSTADDRPOINTER_REG_26__SCAN_IN, P2_U5673);
  nand ginst15465 (P2_U5896, P2_R2096_U80, P2_U2390);
  nand ginst15466 (P2_U5897, P2_R2099_U76, P2_U2389);
  nand ginst15467 (P2_U5898, P2_R2027_U77, P2_U2388);
  nand ginst15468 (P2_U5899, P2_ADD_394_U77, P2_U2386);
  nand ginst15469 (P2_U5900, P2_R2278_U95, P2_U2385);
  nand ginst15470 (P2_U5901, P2_ADD_371_1212_U74, P2_U2384);
  nand ginst15471 (P2_U5902, P2_REIP_REG_27__SCAN_IN, P2_U2381);
  nand ginst15472 (P2_U5903, P2_INSTADDRPOINTER_REG_27__SCAN_IN, P2_U5673);
  nand ginst15473 (P2_U5904, P2_R2096_U79, P2_U2390);
  nand ginst15474 (P2_U5905, P2_R2099_U75, P2_U2389);
  nand ginst15475 (P2_U5906, P2_R2027_U76, P2_U2388);
  nand ginst15476 (P2_U5907, P2_ADD_394_U86, P2_U2386);
  nand ginst15477 (P2_U5908, P2_R2278_U94, P2_U2385);
  nand ginst15478 (P2_U5909, P2_ADD_371_1212_U23, P2_U2384);
  nand ginst15479 (P2_U5910, P2_REIP_REG_28__SCAN_IN, P2_U2381);
  nand ginst15480 (P2_U5911, P2_INSTADDRPOINTER_REG_28__SCAN_IN, P2_U5673);
  nand ginst15481 (P2_U5912, P2_R2096_U78, P2_U2390);
  nand ginst15482 (P2_U5913, P2_R2099_U74, P2_U2389);
  nand ginst15483 (P2_U5914, P2_R2027_U75, P2_U2388);
  nand ginst15484 (P2_U5915, P2_ADD_394_U65, P2_U2386);
  nand ginst15485 (P2_U5916, P2_R2278_U93, P2_U2385);
  nand ginst15486 (P2_U5917, P2_ADD_371_1212_U24, P2_U2384);
  nand ginst15487 (P2_U5918, P2_REIP_REG_29__SCAN_IN, P2_U2381);
  nand ginst15488 (P2_U5919, P2_INSTADDRPOINTER_REG_29__SCAN_IN, P2_U5673);
  nand ginst15489 (P2_U5920, P2_R2096_U76, P2_U2390);
  nand ginst15490 (P2_U5921, P2_R2099_U73, P2_U2389);
  nand ginst15491 (P2_U5922, P2_R2027_U73, P2_U2388);
  nand ginst15492 (P2_U5923, P2_ADD_394_U64, P2_U2386);
  nand ginst15493 (P2_U5924, P2_R2278_U91, P2_U2385);
  nand ginst15494 (P2_U5925, P2_ADD_371_1212_U69, P2_U2384);
  nand ginst15495 (P2_U5926, P2_REIP_REG_30__SCAN_IN, P2_U2381);
  nand ginst15496 (P2_U5927, P2_INSTADDRPOINTER_REG_30__SCAN_IN, P2_U5673);
  nand ginst15497 (P2_U5928, P2_R2096_U50, P2_U2390);
  nand ginst15498 (P2_U5929, P2_R2099_U72, P2_U2389);
  nand ginst15499 (P2_U5930, P2_R2027_U72, P2_U2388);
  nand ginst15500 (P2_U5931, P2_ADD_394_U84, P2_U2386);
  nand ginst15501 (P2_U5932, P2_R2278_U5, P2_U2385);
  nand ginst15502 (P2_U5933, P2_ADD_371_1212_U83, P2_U2384);
  nand ginst15503 (P2_U5934, P2_REIP_REG_31__SCAN_IN, P2_U2381);
  nand ginst15504 (P2_U5935, P2_INSTADDRPOINTER_REG_31__SCAN_IN, P2_U5673);
  nand ginst15505 (P2_U5936, P2_U2374, P2_U4420, P2_U4613);
  nand ginst15506 (P2_U5937, P2_U3284, P2_U5661);
  not ginst15507 (P2_U5938, P2_U3537);
  nand ginst15508 (P2_U5939, P2_STATE2_REG_1__SCAN_IN, P2_U3302);
  nand ginst15509 (P2_U5940, P2_U3540, P2_U5939);
  nand ginst15510 (P2_U5941, P2_PHYADDRPOINTER_REG_0__SCAN_IN, P2_U2387);
  nand ginst15511 (P2_U5942, P2_ADD_371_1212_U68, P2_U2373);
  nand ginst15512 (P2_U5943, P2_R2099_U94, P2_U2372);
  nand ginst15513 (P2_U5944, P2_REIP_REG_0__SCAN_IN, P2_U2371);
  nand ginst15514 (P2_U5945, P2_R2278_U83, P2_U2370);
  nand ginst15515 (P2_U5946, P2_PHYADDRPOINTER_REG_0__SCAN_IN, P2_U5938);
  nand ginst15516 (P2_U5947, P2_R2337_U4, P2_U2387);
  nand ginst15517 (P2_U5948, P2_ADD_371_1212_U25, P2_U2373);
  nand ginst15518 (P2_U5949, P2_R2099_U5, P2_U2372);
  nand ginst15519 (P2_U5950, P2_REIP_REG_1__SCAN_IN, P2_U2371);
  nand ginst15520 (P2_U5951, P2_R2278_U6, P2_U2370);
  nand ginst15521 (P2_U5952, P2_PHYADDRPOINTER_REG_1__SCAN_IN, P2_U5938);
  nand ginst15522 (P2_U5953, P2_R2337_U70, P2_U2387);
  nand ginst15523 (P2_U5954, P2_ADD_371_1212_U79, P2_U2373);
  nand ginst15524 (P2_U5955, P2_R2099_U96, P2_U2372);
  nand ginst15525 (P2_U5956, P2_REIP_REG_2__SCAN_IN, P2_U2371);
  nand ginst15526 (P2_U5957, P2_R2278_U92, P2_U2370);
  nand ginst15527 (P2_U5958, P2_PHYADDRPOINTER_REG_2__SCAN_IN, P2_U5938);
  nand ginst15528 (P2_U5959, P2_R2337_U67, P2_U2387);
  nand ginst15529 (P2_U5960, P2_ADD_371_1212_U84, P2_U2373);
  nand ginst15530 (P2_U5961, P2_R2099_U95, P2_U2372);
  nand ginst15531 (P2_U5962, P2_REIP_REG_3__SCAN_IN, P2_U2371);
  nand ginst15532 (P2_U5963, P2_R2278_U90, P2_U2370);
  nand ginst15533 (P2_U5964, P2_PHYADDRPOINTER_REG_3__SCAN_IN, P2_U5938);
  nand ginst15534 (P2_U5965, P2_R2337_U66, P2_U2387);
  nand ginst15535 (P2_U5966, P2_ADD_371_1212_U80, P2_U2373);
  nand ginst15536 (P2_U5967, P2_R2099_U98, P2_U2372);
  nand ginst15537 (P2_U5968, P2_REIP_REG_4__SCAN_IN, P2_U2371);
  nand ginst15538 (P2_U5969, P2_R2278_U89, P2_U2370);
  nand ginst15539 (P2_U5970, P2_PHYADDRPOINTER_REG_4__SCAN_IN, P2_U5938);
  nand ginst15540 (P2_U5971, P2_R2337_U65, P2_U2387);
  nand ginst15541 (P2_U5972, P2_ADD_371_1212_U81, P2_U2373);
  nand ginst15542 (P2_U5973, P2_R2099_U71, P2_U2372);
  nand ginst15543 (P2_U5974, P2_REIP_REG_5__SCAN_IN, P2_U2371);
  nand ginst15544 (P2_U5975, P2_R2278_U88, P2_U2370);
  nand ginst15545 (P2_U5976, P2_PHYADDRPOINTER_REG_5__SCAN_IN, P2_U5938);
  nand ginst15546 (P2_U5977, P2_R2337_U64, P2_U2387);
  nand ginst15547 (P2_U5978, P2_ADD_371_1212_U78, P2_U2373);
  nand ginst15548 (P2_U5979, P2_R2099_U70, P2_U2372);
  nand ginst15549 (P2_U5980, P2_REIP_REG_6__SCAN_IN, P2_U2371);
  nand ginst15550 (P2_U5981, P2_R2278_U87, P2_U2370);
  nand ginst15551 (P2_U5982, P2_PHYADDRPOINTER_REG_6__SCAN_IN, P2_U5938);
  nand ginst15552 (P2_U5983, P2_R2337_U63, P2_U2387);
  nand ginst15553 (P2_U5984, P2_ADD_371_1212_U85, P2_U2373);
  nand ginst15554 (P2_U5985, P2_R2099_U69, P2_U2372);
  nand ginst15555 (P2_U5986, P2_REIP_REG_7__SCAN_IN, P2_U2371);
  nand ginst15556 (P2_U5987, P2_R2278_U86, P2_U2370);
  nand ginst15557 (P2_U5988, P2_PHYADDRPOINTER_REG_7__SCAN_IN, P2_U5938);
  nand ginst15558 (P2_U5989, P2_R2337_U62, P2_U2387);
  nand ginst15559 (P2_U5990, P2_ADD_371_1212_U82, P2_U2373);
  nand ginst15560 (P2_U5991, P2_R2099_U68, P2_U2372);
  nand ginst15561 (P2_U5992, P2_REIP_REG_8__SCAN_IN, P2_U2371);
  nand ginst15562 (P2_U5993, P2_R2278_U85, P2_U2370);
  nand ginst15563 (P2_U5994, P2_PHYADDRPOINTER_REG_8__SCAN_IN, P2_U5938);
  nand ginst15564 (P2_U5995, P2_R2337_U61, P2_U2387);
  nand ginst15565 (P2_U5996, P2_ADD_371_1212_U118, P2_U2373);
  nand ginst15566 (P2_U5997, P2_R2099_U67, P2_U2372);
  nand ginst15567 (P2_U5998, P2_REIP_REG_9__SCAN_IN, P2_U2371);
  nand ginst15568 (P2_U5999, P2_R2278_U84, P2_U2370);
  nand ginst15569 (P2_U6000, P2_PHYADDRPOINTER_REG_9__SCAN_IN, P2_U5938);
  nand ginst15570 (P2_U6001, P2_R2337_U90, P2_U2387);
  nand ginst15571 (P2_U6002, P2_ADD_371_1212_U13, P2_U2373);
  nand ginst15572 (P2_U6003, P2_R2099_U93, P2_U2372);
  nand ginst15573 (P2_U6004, P2_REIP_REG_10__SCAN_IN, P2_U2371);
  nand ginst15574 (P2_U6005, P2_R2278_U112, P2_U2370);
  nand ginst15575 (P2_U6006, P2_PHYADDRPOINTER_REG_10__SCAN_IN, P2_U5938);
  nand ginst15576 (P2_U6007, P2_R2337_U89, P2_U2387);
  nand ginst15577 (P2_U6008, P2_ADD_371_1212_U14, P2_U2373);
  nand ginst15578 (P2_U6009, P2_R2099_U92, P2_U2372);
  nand ginst15579 (P2_U6010, P2_REIP_REG_11__SCAN_IN, P2_U2371);
  nand ginst15580 (P2_U6011, P2_R2278_U111, P2_U2370);
  nand ginst15581 (P2_U6012, P2_PHYADDRPOINTER_REG_11__SCAN_IN, P2_U5938);
  nand ginst15582 (P2_U6013, P2_R2337_U88, P2_U2387);
  nand ginst15583 (P2_U6014, P2_ADD_371_1212_U76, P2_U2373);
  nand ginst15584 (P2_U6015, P2_R2099_U91, P2_U2372);
  nand ginst15585 (P2_U6016, P2_REIP_REG_12__SCAN_IN, P2_U2371);
  nand ginst15586 (P2_U6017, P2_R2278_U110, P2_U2370);
  nand ginst15587 (P2_U6018, P2_PHYADDRPOINTER_REG_12__SCAN_IN, P2_U5938);
  nand ginst15588 (P2_U6019, P2_R2337_U87, P2_U2387);
  nand ginst15589 (P2_U6020, P2_ADD_371_1212_U15, P2_U2373);
  nand ginst15590 (P2_U6021, P2_R2099_U90, P2_U2372);
  nand ginst15591 (P2_U6022, P2_REIP_REG_13__SCAN_IN, P2_U2371);
  nand ginst15592 (P2_U6023, P2_R2278_U109, P2_U2370);
  nand ginst15593 (P2_U6024, P2_PHYADDRPOINTER_REG_13__SCAN_IN, P2_U5938);
  nand ginst15594 (P2_U6025, P2_R2337_U86, P2_U2387);
  nand ginst15595 (P2_U6026, P2_ADD_371_1212_U16, P2_U2373);
  nand ginst15596 (P2_U6027, P2_R2099_U89, P2_U2372);
  nand ginst15597 (P2_U6028, P2_REIP_REG_14__SCAN_IN, P2_U2371);
  nand ginst15598 (P2_U6029, P2_R2278_U108, P2_U2370);
  nand ginst15599 (P2_U6030, P2_PHYADDRPOINTER_REG_14__SCAN_IN, P2_U5938);
  nand ginst15600 (P2_U6031, P2_R2337_U85, P2_U2387);
  nand ginst15601 (P2_U6032, P2_ADD_371_1212_U73, P2_U2373);
  nand ginst15602 (P2_U6033, P2_R2099_U88, P2_U2372);
  nand ginst15603 (P2_U6034, P2_REIP_REG_15__SCAN_IN, P2_U2371);
  nand ginst15604 (P2_U6035, P2_R2278_U107, P2_U2370);
  nand ginst15605 (P2_U6036, P2_PHYADDRPOINTER_REG_15__SCAN_IN, P2_U5938);
  nand ginst15606 (P2_U6037, P2_R2337_U84, P2_U2387);
  nand ginst15607 (P2_U6038, P2_ADD_371_1212_U17, P2_U2373);
  nand ginst15608 (P2_U6039, P2_R2099_U87, P2_U2372);
  nand ginst15609 (P2_U6040, P2_REIP_REG_16__SCAN_IN, P2_U2371);
  nand ginst15610 (P2_U6041, P2_R2278_U106, P2_U2370);
  nand ginst15611 (P2_U6042, P2_PHYADDRPOINTER_REG_16__SCAN_IN, P2_U5938);
  nand ginst15612 (P2_U6043, P2_R2337_U83, P2_U2387);
  nand ginst15613 (P2_U6044, P2_ADD_371_1212_U71, P2_U2373);
  nand ginst15614 (P2_U6045, P2_R2099_U86, P2_U2372);
  nand ginst15615 (P2_U6046, P2_REIP_REG_17__SCAN_IN, P2_U2371);
  nand ginst15616 (P2_U6047, P2_R2278_U105, P2_U2370);
  nand ginst15617 (P2_U6048, P2_PHYADDRPOINTER_REG_17__SCAN_IN, P2_U5938);
  nand ginst15618 (P2_U6049, P2_R2337_U82, P2_U2387);
  nand ginst15619 (P2_U6050, P2_ADD_371_1212_U72, P2_U2373);
  nand ginst15620 (P2_U6051, P2_R2099_U85, P2_U2372);
  nand ginst15621 (P2_U6052, P2_REIP_REG_18__SCAN_IN, P2_U2371);
  nand ginst15622 (P2_U6053, P2_R2278_U104, P2_U2370);
  nand ginst15623 (P2_U6054, P2_PHYADDRPOINTER_REG_18__SCAN_IN, P2_U5938);
  nand ginst15624 (P2_U6055, P2_R2337_U81, P2_U2387);
  nand ginst15625 (P2_U6056, P2_ADD_371_1212_U18, P2_U2373);
  nand ginst15626 (P2_U6057, P2_R2099_U84, P2_U2372);
  nand ginst15627 (P2_U6058, P2_REIP_REG_19__SCAN_IN, P2_U2371);
  nand ginst15628 (P2_U6059, P2_R2278_U103, P2_U2370);
  nand ginst15629 (P2_U6060, P2_PHYADDRPOINTER_REG_19__SCAN_IN, P2_U5938);
  nand ginst15630 (P2_U6061, P2_R2337_U80, P2_U2387);
  nand ginst15631 (P2_U6062, P2_ADD_371_1212_U19, P2_U2373);
  nand ginst15632 (P2_U6063, P2_R2099_U83, P2_U2372);
  nand ginst15633 (P2_U6064, P2_REIP_REG_20__SCAN_IN, P2_U2371);
  nand ginst15634 (P2_U6065, P2_R2278_U102, P2_U2370);
  nand ginst15635 (P2_U6066, P2_PHYADDRPOINTER_REG_20__SCAN_IN, P2_U5938);
  nand ginst15636 (P2_U6067, P2_R2337_U79, P2_U2387);
  nand ginst15637 (P2_U6068, P2_ADD_371_1212_U75, P2_U2373);
  nand ginst15638 (P2_U6069, P2_R2099_U82, P2_U2372);
  nand ginst15639 (P2_U6070, P2_REIP_REG_21__SCAN_IN, P2_U2371);
  nand ginst15640 (P2_U6071, P2_R2278_U101, P2_U2370);
  nand ginst15641 (P2_U6072, P2_PHYADDRPOINTER_REG_21__SCAN_IN, P2_U5938);
  nand ginst15642 (P2_U6073, P2_R2337_U78, P2_U2387);
  nand ginst15643 (P2_U6074, P2_ADD_371_1212_U20, P2_U2373);
  nand ginst15644 (P2_U6075, P2_R2099_U81, P2_U2372);
  nand ginst15645 (P2_U6076, P2_REIP_REG_22__SCAN_IN, P2_U2371);
  nand ginst15646 (P2_U6077, P2_R2278_U100, P2_U2370);
  nand ginst15647 (P2_U6078, P2_PHYADDRPOINTER_REG_22__SCAN_IN, P2_U5938);
  nand ginst15648 (P2_U6079, P2_R2337_U77, P2_U2387);
  nand ginst15649 (P2_U6080, P2_ADD_371_1212_U21, P2_U2373);
  nand ginst15650 (P2_U6081, P2_R2099_U80, P2_U2372);
  nand ginst15651 (P2_U6082, P2_REIP_REG_23__SCAN_IN, P2_U2371);
  nand ginst15652 (P2_U6083, P2_R2278_U99, P2_U2370);
  nand ginst15653 (P2_U6084, P2_PHYADDRPOINTER_REG_23__SCAN_IN, P2_U5938);
  nand ginst15654 (P2_U6085, P2_R2337_U76, P2_U2387);
  nand ginst15655 (P2_U6086, P2_ADD_371_1212_U70, P2_U2373);
  nand ginst15656 (P2_U6087, P2_R2099_U79, P2_U2372);
  nand ginst15657 (P2_U6088, P2_REIP_REG_24__SCAN_IN, P2_U2371);
  nand ginst15658 (P2_U6089, P2_R2278_U98, P2_U2370);
  nand ginst15659 (P2_U6090, P2_PHYADDRPOINTER_REG_24__SCAN_IN, P2_U5938);
  nand ginst15660 (P2_U6091, P2_R2337_U75, P2_U2387);
  nand ginst15661 (P2_U6092, P2_ADD_371_1212_U77, P2_U2373);
  nand ginst15662 (P2_U6093, P2_R2099_U78, P2_U2372);
  nand ginst15663 (P2_U6094, P2_REIP_REG_25__SCAN_IN, P2_U2371);
  nand ginst15664 (P2_U6095, P2_R2278_U97, P2_U2370);
  nand ginst15665 (P2_U6096, P2_PHYADDRPOINTER_REG_25__SCAN_IN, P2_U5938);
  nand ginst15666 (P2_U6097, P2_R2337_U74, P2_U2387);
  nand ginst15667 (P2_U6098, P2_ADD_371_1212_U22, P2_U2373);
  nand ginst15668 (P2_U6099, P2_R2099_U77, P2_U2372);
  nand ginst15669 (P2_U6100, P2_REIP_REG_26__SCAN_IN, P2_U2371);
  nand ginst15670 (P2_U6101, P2_R2278_U96, P2_U2370);
  nand ginst15671 (P2_U6102, P2_PHYADDRPOINTER_REG_26__SCAN_IN, P2_U5938);
  nand ginst15672 (P2_U6103, P2_R2337_U73, P2_U2387);
  nand ginst15673 (P2_U6104, P2_ADD_371_1212_U74, P2_U2373);
  nand ginst15674 (P2_U6105, P2_R2099_U76, P2_U2372);
  nand ginst15675 (P2_U6106, P2_REIP_REG_27__SCAN_IN, P2_U2371);
  nand ginst15676 (P2_U6107, P2_R2278_U95, P2_U2370);
  nand ginst15677 (P2_U6108, P2_PHYADDRPOINTER_REG_27__SCAN_IN, P2_U5938);
  nand ginst15678 (P2_U6109, P2_R2337_U72, P2_U2387);
  nand ginst15679 (P2_U6110, P2_ADD_371_1212_U23, P2_U2373);
  nand ginst15680 (P2_U6111, P2_R2099_U75, P2_U2372);
  nand ginst15681 (P2_U6112, P2_REIP_REG_28__SCAN_IN, P2_U2371);
  nand ginst15682 (P2_U6113, P2_R2278_U94, P2_U2370);
  nand ginst15683 (P2_U6114, P2_PHYADDRPOINTER_REG_28__SCAN_IN, P2_U5938);
  nand ginst15684 (P2_U6115, P2_R2337_U71, P2_U2387);
  nand ginst15685 (P2_U6116, P2_ADD_371_1212_U24, P2_U2373);
  nand ginst15686 (P2_U6117, P2_R2099_U74, P2_U2372);
  nand ginst15687 (P2_U6118, P2_REIP_REG_29__SCAN_IN, P2_U2371);
  nand ginst15688 (P2_U6119, P2_R2278_U93, P2_U2370);
  nand ginst15689 (P2_U6120, P2_PHYADDRPOINTER_REG_29__SCAN_IN, P2_U5938);
  nand ginst15690 (P2_U6121, P2_R2337_U69, P2_U2387);
  nand ginst15691 (P2_U6122, P2_ADD_371_1212_U69, P2_U2373);
  nand ginst15692 (P2_U6123, P2_R2099_U73, P2_U2372);
  nand ginst15693 (P2_U6124, P2_REIP_REG_30__SCAN_IN, P2_U2371);
  nand ginst15694 (P2_U6125, P2_R2278_U91, P2_U2370);
  nand ginst15695 (P2_U6126, P2_PHYADDRPOINTER_REG_30__SCAN_IN, P2_U5938);
  nand ginst15696 (P2_U6127, P2_R2337_U68, P2_U2387);
  nand ginst15697 (P2_U6128, P2_ADD_371_1212_U83, P2_U2373);
  nand ginst15698 (P2_U6129, P2_R2099_U72, P2_U2372);
  nand ginst15699 (P2_U6130, P2_REIP_REG_31__SCAN_IN, P2_U2371);
  nand ginst15700 (P2_U6131, P2_R2278_U5, P2_U2370);
  nand ginst15701 (P2_U6132, P2_PHYADDRPOINTER_REG_31__SCAN_IN, P2_U5938);
  nand ginst15702 (P2_U6133, P2_U2616, U211);
  nand ginst15703 (P2_U6134, P2_EAX_REG_15__SCAN_IN, P2_U2395);
  nand ginst15704 (P2_U6135, P2_U2394, U308);
  nand ginst15705 (P2_U6136, P2_LWORD_REG_15__SCAN_IN, P2_U3538);
  nand ginst15706 (P2_U6137, P2_EAX_REG_14__SCAN_IN, P2_U2395);
  nand ginst15707 (P2_U6138, P2_U2394, U309);
  nand ginst15708 (P2_U6139, P2_LWORD_REG_14__SCAN_IN, P2_U3538);
  nand ginst15709 (P2_U6140, P2_EAX_REG_13__SCAN_IN, P2_U2395);
  nand ginst15710 (P2_U6141, P2_U2394, U310);
  nand ginst15711 (P2_U6142, P2_LWORD_REG_13__SCAN_IN, P2_U3538);
  nand ginst15712 (P2_U6143, P2_EAX_REG_12__SCAN_IN, P2_U2395);
  nand ginst15713 (P2_U6144, P2_U2394, U311);
  nand ginst15714 (P2_U6145, P2_LWORD_REG_12__SCAN_IN, P2_U3538);
  nand ginst15715 (P2_U6146, P2_EAX_REG_11__SCAN_IN, P2_U2395);
  nand ginst15716 (P2_U6147, P2_U2394, U312);
  nand ginst15717 (P2_U6148, P2_LWORD_REG_11__SCAN_IN, P2_U3538);
  nand ginst15718 (P2_U6149, P2_EAX_REG_10__SCAN_IN, P2_U2395);
  nand ginst15719 (P2_U6150, P2_U2394, U313);
  nand ginst15720 (P2_U6151, P2_LWORD_REG_10__SCAN_IN, P2_U3538);
  nand ginst15721 (P2_U6152, P2_EAX_REG_9__SCAN_IN, P2_U2395);
  nand ginst15722 (P2_U6153, P2_U2394, U283);
  nand ginst15723 (P2_U6154, P2_LWORD_REG_9__SCAN_IN, P2_U3538);
  nand ginst15724 (P2_U6155, P2_EAX_REG_8__SCAN_IN, P2_U2395);
  nand ginst15725 (P2_U6156, P2_U2394, U284);
  nand ginst15726 (P2_U6157, P2_LWORD_REG_8__SCAN_IN, P2_U3538);
  nand ginst15727 (P2_U6158, P2_EAX_REG_7__SCAN_IN, P2_U2395);
  nand ginst15728 (P2_U6159, P2_U2394, U285);
  nand ginst15729 (P2_U6160, P2_LWORD_REG_7__SCAN_IN, P2_U3538);
  nand ginst15730 (P2_U6161, P2_EAX_REG_6__SCAN_IN, P2_U2395);
  nand ginst15731 (P2_U6162, P2_U2394, U286);
  nand ginst15732 (P2_U6163, P2_LWORD_REG_6__SCAN_IN, P2_U3538);
  nand ginst15733 (P2_U6164, P2_EAX_REG_5__SCAN_IN, P2_U2395);
  nand ginst15734 (P2_U6165, P2_U2394, U287);
  nand ginst15735 (P2_U6166, P2_LWORD_REG_5__SCAN_IN, P2_U3538);
  nand ginst15736 (P2_U6167, P2_EAX_REG_4__SCAN_IN, P2_U2395);
  nand ginst15737 (P2_U6168, P2_U2394, U288);
  nand ginst15738 (P2_U6169, P2_LWORD_REG_4__SCAN_IN, P2_U3538);
  nand ginst15739 (P2_U6170, P2_EAX_REG_3__SCAN_IN, P2_U2395);
  nand ginst15740 (P2_U6171, P2_U2394, U289);
  nand ginst15741 (P2_U6172, P2_LWORD_REG_3__SCAN_IN, P2_U3538);
  nand ginst15742 (P2_U6173, P2_EAX_REG_2__SCAN_IN, P2_U2395);
  nand ginst15743 (P2_U6174, P2_U2394, U292);
  nand ginst15744 (P2_U6175, P2_LWORD_REG_2__SCAN_IN, P2_U3538);
  nand ginst15745 (P2_U6176, P2_EAX_REG_1__SCAN_IN, P2_U2395);
  nand ginst15746 (P2_U6177, P2_U2394, U303);
  nand ginst15747 (P2_U6178, P2_LWORD_REG_1__SCAN_IN, P2_U3538);
  nand ginst15748 (P2_U6179, P2_EAX_REG_0__SCAN_IN, P2_U2395);
  nand ginst15749 (P2_U6180, P2_U2394, U314);
  nand ginst15750 (P2_U6181, P2_LWORD_REG_0__SCAN_IN, P2_U3538);
  nand ginst15751 (P2_U6182, P2_EAX_REG_30__SCAN_IN, P2_U2395);
  nand ginst15752 (P2_U6183, P2_U2394, U309);
  nand ginst15753 (P2_U6184, P2_UWORD_REG_14__SCAN_IN, P2_U3538);
  nand ginst15754 (P2_U6185, P2_EAX_REG_29__SCAN_IN, P2_U2395);
  nand ginst15755 (P2_U6186, P2_U2394, U310);
  nand ginst15756 (P2_U6187, P2_UWORD_REG_13__SCAN_IN, P2_U3538);
  nand ginst15757 (P2_U6188, P2_EAX_REG_28__SCAN_IN, P2_U2395);
  nand ginst15758 (P2_U6189, P2_U2394, U311);
  nand ginst15759 (P2_U6190, P2_UWORD_REG_12__SCAN_IN, P2_U3538);
  nand ginst15760 (P2_U6191, P2_EAX_REG_27__SCAN_IN, P2_U2395);
  nand ginst15761 (P2_U6192, P2_U2394, U312);
  nand ginst15762 (P2_U6193, P2_UWORD_REG_11__SCAN_IN, P2_U3538);
  nand ginst15763 (P2_U6194, P2_EAX_REG_26__SCAN_IN, P2_U2395);
  nand ginst15764 (P2_U6195, P2_U2394, U313);
  nand ginst15765 (P2_U6196, P2_UWORD_REG_10__SCAN_IN, P2_U3538);
  nand ginst15766 (P2_U6197, P2_EAX_REG_25__SCAN_IN, P2_U2395);
  nand ginst15767 (P2_U6198, P2_U2394, U283);
  nand ginst15768 (P2_U6199, P2_UWORD_REG_9__SCAN_IN, P2_U3538);
  nand ginst15769 (P2_U6200, P2_EAX_REG_24__SCAN_IN, P2_U2395);
  nand ginst15770 (P2_U6201, P2_U2394, U284);
  nand ginst15771 (P2_U6202, P2_UWORD_REG_8__SCAN_IN, P2_U3538);
  nand ginst15772 (P2_U6203, P2_EAX_REG_23__SCAN_IN, P2_U2395);
  nand ginst15773 (P2_U6204, P2_U2394, U285);
  nand ginst15774 (P2_U6205, P2_UWORD_REG_7__SCAN_IN, P2_U3538);
  nand ginst15775 (P2_U6206, P2_EAX_REG_22__SCAN_IN, P2_U2395);
  nand ginst15776 (P2_U6207, P2_U2394, U286);
  nand ginst15777 (P2_U6208, P2_UWORD_REG_6__SCAN_IN, P2_U3538);
  nand ginst15778 (P2_U6209, P2_EAX_REG_21__SCAN_IN, P2_U2395);
  nand ginst15779 (P2_U6210, P2_U2394, U287);
  nand ginst15780 (P2_U6211, P2_UWORD_REG_5__SCAN_IN, P2_U3538);
  nand ginst15781 (P2_U6212, P2_EAX_REG_20__SCAN_IN, P2_U2395);
  nand ginst15782 (P2_U6213, P2_U2394, U288);
  nand ginst15783 (P2_U6214, P2_UWORD_REG_4__SCAN_IN, P2_U3538);
  nand ginst15784 (P2_U6215, P2_EAX_REG_19__SCAN_IN, P2_U2395);
  nand ginst15785 (P2_U6216, P2_U2394, U289);
  nand ginst15786 (P2_U6217, P2_UWORD_REG_3__SCAN_IN, P2_U3538);
  nand ginst15787 (P2_U6218, P2_EAX_REG_18__SCAN_IN, P2_U2395);
  nand ginst15788 (P2_U6219, P2_U2394, U292);
  nand ginst15789 (P2_U6220, P2_UWORD_REG_2__SCAN_IN, P2_U3538);
  nand ginst15790 (P2_U6221, P2_EAX_REG_17__SCAN_IN, P2_U2395);
  nand ginst15791 (P2_U6222, P2_U2394, U303);
  nand ginst15792 (P2_U6223, P2_UWORD_REG_1__SCAN_IN, P2_U3538);
  nand ginst15793 (P2_U6224, P2_EAX_REG_16__SCAN_IN, P2_U2395);
  nand ginst15794 (P2_U6225, P2_U2394, U314);
  nand ginst15795 (P2_U6226, P2_UWORD_REG_0__SCAN_IN, P2_U3538);
  nand ginst15796 (P2_U6227, P2_R2167_U6, P2_U4057, P2_U4421);
  nand ginst15797 (P2_U6228, P2_U2446, P2_U4058);
  nand ginst15798 (P2_U6229, P2_U6227, P2_U6228);
  nand ginst15799 (P2_U6230, P2_U4411, P2_U6229);
  nand ginst15800 (P2_U6231, P2_STATE2_REG_1__SCAN_IN, P2_U4467);
  not ginst15801 (P2_U6232, P2_U3541);
  nand ginst15802 (P2_U6233, P2_EAX_REG_0__SCAN_IN, P2_U2430);
  nand ginst15803 (P2_U6234, P2_LWORD_REG_0__SCAN_IN, P2_U2396);
  nand ginst15804 (P2_U6235, P2_DATAO_REG_0__SCAN_IN, P2_U6232);
  nand ginst15805 (P2_U6236, P2_EAX_REG_1__SCAN_IN, P2_U2430);
  nand ginst15806 (P2_U6237, P2_LWORD_REG_1__SCAN_IN, P2_U2396);
  nand ginst15807 (P2_U6238, P2_DATAO_REG_1__SCAN_IN, P2_U6232);
  nand ginst15808 (P2_U6239, P2_EAX_REG_2__SCAN_IN, P2_U2430);
  nand ginst15809 (P2_U6240, P2_LWORD_REG_2__SCAN_IN, P2_U2396);
  nand ginst15810 (P2_U6241, P2_DATAO_REG_2__SCAN_IN, P2_U6232);
  nand ginst15811 (P2_U6242, P2_EAX_REG_3__SCAN_IN, P2_U2430);
  nand ginst15812 (P2_U6243, P2_LWORD_REG_3__SCAN_IN, P2_U2396);
  nand ginst15813 (P2_U6244, P2_DATAO_REG_3__SCAN_IN, P2_U6232);
  nand ginst15814 (P2_U6245, P2_EAX_REG_4__SCAN_IN, P2_U2430);
  nand ginst15815 (P2_U6246, P2_LWORD_REG_4__SCAN_IN, P2_U2396);
  nand ginst15816 (P2_U6247, P2_DATAO_REG_4__SCAN_IN, P2_U6232);
  nand ginst15817 (P2_U6248, P2_EAX_REG_5__SCAN_IN, P2_U2430);
  nand ginst15818 (P2_U6249, P2_LWORD_REG_5__SCAN_IN, P2_U2396);
  nand ginst15819 (P2_U6250, P2_DATAO_REG_5__SCAN_IN, P2_U6232);
  nand ginst15820 (P2_U6251, P2_EAX_REG_6__SCAN_IN, P2_U2430);
  nand ginst15821 (P2_U6252, P2_LWORD_REG_6__SCAN_IN, P2_U2396);
  nand ginst15822 (P2_U6253, P2_DATAO_REG_6__SCAN_IN, P2_U6232);
  nand ginst15823 (P2_U6254, P2_EAX_REG_7__SCAN_IN, P2_U2430);
  nand ginst15824 (P2_U6255, P2_LWORD_REG_7__SCAN_IN, P2_U2396);
  nand ginst15825 (P2_U6256, P2_DATAO_REG_7__SCAN_IN, P2_U6232);
  nand ginst15826 (P2_U6257, P2_EAX_REG_8__SCAN_IN, P2_U2430);
  nand ginst15827 (P2_U6258, P2_LWORD_REG_8__SCAN_IN, P2_U2396);
  nand ginst15828 (P2_U6259, P2_DATAO_REG_8__SCAN_IN, P2_U6232);
  nand ginst15829 (P2_U6260, P2_EAX_REG_9__SCAN_IN, P2_U2430);
  nand ginst15830 (P2_U6261, P2_LWORD_REG_9__SCAN_IN, P2_U2396);
  nand ginst15831 (P2_U6262, P2_DATAO_REG_9__SCAN_IN, P2_U6232);
  nand ginst15832 (P2_U6263, P2_EAX_REG_10__SCAN_IN, P2_U2430);
  nand ginst15833 (P2_U6264, P2_LWORD_REG_10__SCAN_IN, P2_U2396);
  nand ginst15834 (P2_U6265, P2_DATAO_REG_10__SCAN_IN, P2_U6232);
  nand ginst15835 (P2_U6266, P2_EAX_REG_11__SCAN_IN, P2_U2430);
  nand ginst15836 (P2_U6267, P2_LWORD_REG_11__SCAN_IN, P2_U2396);
  nand ginst15837 (P2_U6268, P2_DATAO_REG_11__SCAN_IN, P2_U6232);
  nand ginst15838 (P2_U6269, P2_EAX_REG_12__SCAN_IN, P2_U2430);
  nand ginst15839 (P2_U6270, P2_LWORD_REG_12__SCAN_IN, P2_U2396);
  nand ginst15840 (P2_U6271, P2_DATAO_REG_12__SCAN_IN, P2_U6232);
  nand ginst15841 (P2_U6272, P2_EAX_REG_13__SCAN_IN, P2_U2430);
  nand ginst15842 (P2_U6273, P2_LWORD_REG_13__SCAN_IN, P2_U2396);
  nand ginst15843 (P2_U6274, P2_DATAO_REG_13__SCAN_IN, P2_U6232);
  nand ginst15844 (P2_U6275, P2_EAX_REG_14__SCAN_IN, P2_U2430);
  nand ginst15845 (P2_U6276, P2_LWORD_REG_14__SCAN_IN, P2_U2396);
  nand ginst15846 (P2_U6277, P2_DATAO_REG_14__SCAN_IN, P2_U6232);
  nand ginst15847 (P2_U6278, P2_EAX_REG_15__SCAN_IN, P2_U2430);
  nand ginst15848 (P2_U6279, P2_LWORD_REG_15__SCAN_IN, P2_U2396);
  nand ginst15849 (P2_U6280, P2_DATAO_REG_15__SCAN_IN, P2_U6232);
  nand ginst15850 (P2_U6281, P2_EAX_REG_16__SCAN_IN, P2_U2435);
  nand ginst15851 (P2_U6282, P2_UWORD_REG_0__SCAN_IN, P2_U2396);
  nand ginst15852 (P2_U6283, P2_DATAO_REG_16__SCAN_IN, P2_U6232);
  nand ginst15853 (P2_U6284, P2_EAX_REG_17__SCAN_IN, P2_U2435);
  nand ginst15854 (P2_U6285, P2_UWORD_REG_1__SCAN_IN, P2_U2396);
  nand ginst15855 (P2_U6286, P2_DATAO_REG_17__SCAN_IN, P2_U6232);
  nand ginst15856 (P2_U6287, P2_EAX_REG_18__SCAN_IN, P2_U2435);
  nand ginst15857 (P2_U6288, P2_UWORD_REG_2__SCAN_IN, P2_U2396);
  nand ginst15858 (P2_U6289, P2_DATAO_REG_18__SCAN_IN, P2_U6232);
  nand ginst15859 (P2_U6290, P2_EAX_REG_19__SCAN_IN, P2_U2435);
  nand ginst15860 (P2_U6291, P2_UWORD_REG_3__SCAN_IN, P2_U2396);
  nand ginst15861 (P2_U6292, P2_DATAO_REG_19__SCAN_IN, P2_U6232);
  nand ginst15862 (P2_U6293, P2_EAX_REG_20__SCAN_IN, P2_U2435);
  nand ginst15863 (P2_U6294, P2_UWORD_REG_4__SCAN_IN, P2_U2396);
  nand ginst15864 (P2_U6295, P2_DATAO_REG_20__SCAN_IN, P2_U6232);
  nand ginst15865 (P2_U6296, P2_EAX_REG_21__SCAN_IN, P2_U2435);
  nand ginst15866 (P2_U6297, P2_UWORD_REG_5__SCAN_IN, P2_U2396);
  nand ginst15867 (P2_U6298, P2_DATAO_REG_21__SCAN_IN, P2_U6232);
  nand ginst15868 (P2_U6299, P2_EAX_REG_22__SCAN_IN, P2_U2435);
  nand ginst15869 (P2_U6300, P2_UWORD_REG_6__SCAN_IN, P2_U2396);
  nand ginst15870 (P2_U6301, P2_DATAO_REG_22__SCAN_IN, P2_U6232);
  nand ginst15871 (P2_U6302, P2_EAX_REG_23__SCAN_IN, P2_U2435);
  nand ginst15872 (P2_U6303, P2_UWORD_REG_7__SCAN_IN, P2_U2396);
  nand ginst15873 (P2_U6304, P2_DATAO_REG_23__SCAN_IN, P2_U6232);
  nand ginst15874 (P2_U6305, P2_EAX_REG_24__SCAN_IN, P2_U2435);
  nand ginst15875 (P2_U6306, P2_UWORD_REG_8__SCAN_IN, P2_U2396);
  nand ginst15876 (P2_U6307, P2_DATAO_REG_24__SCAN_IN, P2_U6232);
  nand ginst15877 (P2_U6308, P2_EAX_REG_25__SCAN_IN, P2_U2435);
  nand ginst15878 (P2_U6309, P2_UWORD_REG_9__SCAN_IN, P2_U2396);
  nand ginst15879 (P2_U6310, P2_DATAO_REG_25__SCAN_IN, P2_U6232);
  nand ginst15880 (P2_U6311, P2_EAX_REG_26__SCAN_IN, P2_U2435);
  nand ginst15881 (P2_U6312, P2_UWORD_REG_10__SCAN_IN, P2_U2396);
  nand ginst15882 (P2_U6313, P2_DATAO_REG_26__SCAN_IN, P2_U6232);
  nand ginst15883 (P2_U6314, P2_EAX_REG_27__SCAN_IN, P2_U2435);
  nand ginst15884 (P2_U6315, P2_UWORD_REG_11__SCAN_IN, P2_U2396);
  nand ginst15885 (P2_U6316, P2_DATAO_REG_27__SCAN_IN, P2_U6232);
  nand ginst15886 (P2_U6317, P2_EAX_REG_28__SCAN_IN, P2_U2435);
  nand ginst15887 (P2_U6318, P2_UWORD_REG_12__SCAN_IN, P2_U2396);
  nand ginst15888 (P2_U6319, P2_DATAO_REG_28__SCAN_IN, P2_U6232);
  nand ginst15889 (P2_U6320, P2_EAX_REG_29__SCAN_IN, P2_U2435);
  nand ginst15890 (P2_U6321, P2_UWORD_REG_13__SCAN_IN, P2_U2396);
  nand ginst15891 (P2_U6322, P2_DATAO_REG_29__SCAN_IN, P2_U6232);
  nand ginst15892 (P2_U6323, P2_EAX_REG_30__SCAN_IN, P2_U2435);
  nand ginst15893 (P2_U6324, P2_UWORD_REG_14__SCAN_IN, P2_U2396);
  nand ginst15894 (P2_U6325, P2_DATAO_REG_30__SCAN_IN, P2_U6232);
  nand ginst15895 (P2_U6326, P2_U2513, P2_U3254);
  nand ginst15896 (P2_U6327, P2_U2433, U314);
  nand ginst15897 (P2_U6328, P2_ADD_391_1196_U87, P2_U2397);
  nand ginst15898 (P2_U6329, P2_R2096_U68, P2_U2380);
  nand ginst15899 (P2_U6330, P2_EAX_REG_0__SCAN_IN, P2_U3542);
  nand ginst15900 (P2_U6331, P2_U2433, U303);
  nand ginst15901 (P2_U6332, P2_ADD_391_1196_U12, P2_U2397);
  nand ginst15902 (P2_U6333, P2_R2096_U51, P2_U2380);
  nand ginst15903 (P2_U6334, P2_EAX_REG_1__SCAN_IN, P2_U3542);
  nand ginst15904 (P2_U6335, P2_U2433, U292);
  nand ginst15905 (P2_U6336, P2_ADD_391_1196_U92, P2_U2397);
  nand ginst15906 (P2_U6337, P2_R2096_U77, P2_U2380);
  nand ginst15907 (P2_U6338, P2_EAX_REG_2__SCAN_IN, P2_U3542);
  nand ginst15908 (P2_U6339, P2_U2433, U289);
  nand ginst15909 (P2_U6340, P2_ADD_391_1196_U91, P2_U2397);
  nand ginst15910 (P2_U6341, P2_R2096_U75, P2_U2380);
  nand ginst15911 (P2_U6342, P2_EAX_REG_3__SCAN_IN, P2_U3542);
  nand ginst15912 (P2_U6343, P2_U2433, U288);
  nand ginst15913 (P2_U6344, P2_ADD_391_1196_U90, P2_U2397);
  nand ginst15914 (P2_U6345, P2_R2096_U74, P2_U2380);
  nand ginst15915 (P2_U6346, P2_EAX_REG_4__SCAN_IN, P2_U3542);
  nand ginst15916 (P2_U6347, P2_U2433, U287);
  nand ginst15917 (P2_U6348, P2_ADD_391_1196_U9, P2_U2397);
  nand ginst15918 (P2_U6349, P2_R2096_U73, P2_U2380);
  nand ginst15919 (P2_U6350, P2_EAX_REG_5__SCAN_IN, P2_U3542);
  nand ginst15920 (P2_U6351, P2_U2433, U286);
  nand ginst15921 (P2_U6352, P2_ADD_391_1196_U89, P2_U2397);
  nand ginst15922 (P2_U6353, P2_R2096_U72, P2_U2380);
  nand ginst15923 (P2_U6354, P2_EAX_REG_6__SCAN_IN, P2_U3542);
  nand ginst15924 (P2_U6355, P2_U2433, U285);
  nand ginst15925 (P2_U6356, P2_ADD_391_1196_U10, P2_U2397);
  nand ginst15926 (P2_U6357, P2_R2096_U71, P2_U2380);
  nand ginst15927 (P2_U6358, P2_EAX_REG_7__SCAN_IN, P2_U3542);
  nand ginst15928 (P2_U6359, P2_U2433, U284);
  nand ginst15929 (P2_U6360, P2_ADD_391_1196_U88, P2_U2397);
  nand ginst15930 (P2_U6361, P2_R2096_U70, P2_U2380);
  nand ginst15931 (P2_U6362, P2_EAX_REG_8__SCAN_IN, P2_U3542);
  nand ginst15932 (P2_U6363, P2_U2433, U283);
  nand ginst15933 (P2_U6364, P2_ADD_391_1196_U11, P2_U2397);
  nand ginst15934 (P2_U6365, P2_R2096_U69, P2_U2380);
  nand ginst15935 (P2_U6366, P2_EAX_REG_9__SCAN_IN, P2_U3542);
  nand ginst15936 (P2_U6367, P2_U2433, U313);
  nand ginst15937 (P2_U6368, P2_ADD_391_1196_U109, P2_U2397);
  nand ginst15938 (P2_U6369, P2_R2096_U97, P2_U2380);
  nand ginst15939 (P2_U6370, P2_EAX_REG_10__SCAN_IN, P2_U3542);
  nand ginst15940 (P2_U6371, P2_U2433, U312);
  nand ginst15941 (P2_U6372, P2_ADD_391_1196_U5, P2_U2397);
  nand ginst15942 (P2_U6373, P2_R2096_U96, P2_U2380);
  nand ginst15943 (P2_U6374, P2_EAX_REG_11__SCAN_IN, P2_U3542);
  nand ginst15944 (P2_U6375, P2_U2433, U311);
  nand ginst15945 (P2_U6376, P2_ADD_391_1196_U108, P2_U2397);
  nand ginst15946 (P2_U6377, P2_R2096_U95, P2_U2380);
  nand ginst15947 (P2_U6378, P2_EAX_REG_12__SCAN_IN, P2_U3542);
  nand ginst15948 (P2_U6379, P2_U2433, U310);
  nand ginst15949 (P2_U6380, P2_ADD_391_1196_U6, P2_U2397);
  nand ginst15950 (P2_U6381, P2_R2096_U94, P2_U2380);
  nand ginst15951 (P2_U6382, P2_EAX_REG_13__SCAN_IN, P2_U3542);
  nand ginst15952 (P2_U6383, P2_U2433, U309);
  nand ginst15953 (P2_U6384, P2_ADD_391_1196_U107, P2_U2397);
  nand ginst15954 (P2_U6385, P2_R2096_U93, P2_U2380);
  nand ginst15955 (P2_U6386, P2_EAX_REG_14__SCAN_IN, P2_U3542);
  nand ginst15956 (P2_U6387, P2_U2433, U308);
  nand ginst15957 (P2_U6388, P2_ADD_391_1196_U7, P2_U2397);
  nand ginst15958 (P2_U6389, P2_R2096_U92, P2_U2380);
  nand ginst15959 (P2_U6390, P2_EAX_REG_15__SCAN_IN, P2_U3542);
  nand ginst15960 (P2_U6391, P2_U2434, U314);
  nand ginst15961 (P2_U6392, P2_U2427, U307);
  nand ginst15962 (P2_U6393, P2_ADD_391_1196_U106, P2_U2397);
  nand ginst15963 (P2_U6394, P2_R2096_U91, P2_U2380);
  nand ginst15964 (P2_U6395, P2_EAX_REG_16__SCAN_IN, P2_U3542);
  nand ginst15965 (P2_U6396, P2_U2434, U303);
  nand ginst15966 (P2_U6397, P2_U2427, U306);
  nand ginst15967 (P2_U6398, P2_ADD_391_1196_U105, P2_U2397);
  nand ginst15968 (P2_U6399, P2_R2096_U90, P2_U2380);
  nand ginst15969 (P2_U6400, P2_EAX_REG_17__SCAN_IN, P2_U3542);
  nand ginst15970 (P2_U6401, P2_U2434, U292);
  nand ginst15971 (P2_U6402, P2_U2427, U305);
  nand ginst15972 (P2_U6403, P2_ADD_391_1196_U104, P2_U2397);
  nand ginst15973 (P2_U6404, P2_R2096_U89, P2_U2380);
  nand ginst15974 (P2_U6405, P2_EAX_REG_18__SCAN_IN, P2_U3542);
  nand ginst15975 (P2_U6406, P2_U2434, U289);
  nand ginst15976 (P2_U6407, P2_U2427, U304);
  nand ginst15977 (P2_U6408, P2_ADD_391_1196_U103, P2_U2397);
  nand ginst15978 (P2_U6409, P2_R2096_U88, P2_U2380);
  nand ginst15979 (P2_U6410, P2_EAX_REG_19__SCAN_IN, P2_U3542);
  nand ginst15980 (P2_U6411, P2_U2434, U288);
  nand ginst15981 (P2_U6412, P2_U2427, U302);
  nand ginst15982 (P2_U6413, P2_ADD_391_1196_U102, P2_U2397);
  nand ginst15983 (P2_U6414, P2_R2096_U87, P2_U2380);
  nand ginst15984 (P2_U6415, P2_EAX_REG_20__SCAN_IN, P2_U3542);
  nand ginst15985 (P2_U6416, P2_U2434, U287);
  nand ginst15986 (P2_U6417, P2_U2427, U301);
  nand ginst15987 (P2_U6418, P2_ADD_391_1196_U101, P2_U2397);
  nand ginst15988 (P2_U6419, P2_R2096_U86, P2_U2380);
  nand ginst15989 (P2_U6420, P2_EAX_REG_21__SCAN_IN, P2_U3542);
  nand ginst15990 (P2_U6421, P2_U2434, U286);
  nand ginst15991 (P2_U6422, P2_U2427, U300);
  nand ginst15992 (P2_U6423, P2_ADD_391_1196_U100, P2_U2397);
  nand ginst15993 (P2_U6424, P2_R2096_U85, P2_U2380);
  nand ginst15994 (P2_U6425, P2_EAX_REG_22__SCAN_IN, P2_U3542);
  nand ginst15995 (P2_U6426, P2_U2434, U285);
  nand ginst15996 (P2_U6427, P2_U2427, U299);
  nand ginst15997 (P2_U6428, P2_ADD_391_1196_U99, P2_U2397);
  nand ginst15998 (P2_U6429, P2_R2096_U84, P2_U2380);
  nand ginst15999 (P2_U6430, P2_EAX_REG_23__SCAN_IN, P2_U3542);
  nand ginst16000 (P2_U6431, P2_U2434, U284);
  nand ginst16001 (P2_U6432, P2_U2427, U298);
  nand ginst16002 (P2_U6433, P2_ADD_391_1196_U98, P2_U2397);
  nand ginst16003 (P2_U6434, P2_R2096_U83, P2_U2380);
  nand ginst16004 (P2_U6435, P2_EAX_REG_24__SCAN_IN, P2_U3542);
  nand ginst16005 (P2_U6436, P2_U2434, U283);
  nand ginst16006 (P2_U6437, P2_U2427, U297);
  nand ginst16007 (P2_U6438, P2_ADD_391_1196_U97, P2_U2397);
  nand ginst16008 (P2_U6439, P2_R2096_U82, P2_U2380);
  nand ginst16009 (P2_U6440, P2_EAX_REG_25__SCAN_IN, P2_U3542);
  nand ginst16010 (P2_U6441, P2_U2434, U313);
  nand ginst16011 (P2_U6442, P2_U2427, U296);
  nand ginst16012 (P2_U6443, P2_ADD_391_1196_U96, P2_U2397);
  nand ginst16013 (P2_U6444, P2_R2096_U81, P2_U2380);
  nand ginst16014 (P2_U6445, P2_EAX_REG_26__SCAN_IN, P2_U3542);
  nand ginst16015 (P2_U6446, P2_U2434, U312);
  nand ginst16016 (P2_U6447, P2_U2427, U295);
  nand ginst16017 (P2_U6448, P2_ADD_391_1196_U95, P2_U2397);
  nand ginst16018 (P2_U6449, P2_R2096_U80, P2_U2380);
  nand ginst16019 (P2_U6450, P2_EAX_REG_27__SCAN_IN, P2_U3542);
  nand ginst16020 (P2_U6451, P2_U2434, U311);
  nand ginst16021 (P2_U6452, P2_U2427, U294);
  nand ginst16022 (P2_U6453, P2_ADD_391_1196_U94, P2_U2397);
  nand ginst16023 (P2_U6454, P2_R2096_U79, P2_U2380);
  nand ginst16024 (P2_U6455, P2_EAX_REG_28__SCAN_IN, P2_U3542);
  nand ginst16025 (P2_U6456, P2_U2434, U310);
  nand ginst16026 (P2_U6457, P2_U2427, U293);
  nand ginst16027 (P2_U6458, P2_ADD_391_1196_U93, P2_U2397);
  nand ginst16028 (P2_U6459, P2_R2096_U78, P2_U2380);
  nand ginst16029 (P2_U6460, P2_EAX_REG_29__SCAN_IN, P2_U3542);
  nand ginst16030 (P2_U6461, P2_U2434, U309);
  nand ginst16031 (P2_U6462, P2_U2427, U291);
  nand ginst16032 (P2_U6463, P2_ADD_391_1196_U8, P2_U2397);
  nand ginst16033 (P2_U6464, P2_R2096_U76, P2_U2380);
  nand ginst16034 (P2_U6465, P2_EAX_REG_30__SCAN_IN, P2_U3542);
  nand ginst16035 (P2_U6466, P2_U2427, U290);
  nand ginst16036 (P2_U6467, P2_R2096_U50, P2_U2380);
  nand ginst16037 (P2_U6468, P2_EAX_REG_31__SCAN_IN, P2_U3542);
  nand ginst16038 (P2_U6469, P2_U3297, P2_U4435);
  nand ginst16039 (P2_U6470, P2_U3578, P2_U6469);
  nand ginst16040 (P2_U6471, P2_R2182_U69, P2_U2393);
  nand ginst16041 (P2_U6472, P2_R2099_U94, P2_U2379);
  nand ginst16042 (P2_U6473, P2_EBX_REG_0__SCAN_IN, P2_U3543);
  nand ginst16043 (P2_U6474, P2_R2182_U68, P2_U2393);
  nand ginst16044 (P2_U6475, P2_R2099_U5, P2_U2379);
  nand ginst16045 (P2_U6476, P2_EBX_REG_1__SCAN_IN, P2_U3543);
  nand ginst16046 (P2_U6477, P2_R2182_U40, P2_U2393);
  nand ginst16047 (P2_U6478, P2_R2099_U96, P2_U2379);
  nand ginst16048 (P2_U6479, P2_EBX_REG_2__SCAN_IN, P2_U3543);
  nand ginst16049 (P2_U6480, P2_R2182_U76, P2_U2393);
  nand ginst16050 (P2_U6481, P2_R2099_U95, P2_U2379);
  nand ginst16051 (P2_U6482, P2_EBX_REG_3__SCAN_IN, P2_U3543);
  nand ginst16052 (P2_U6483, P2_R2182_U75, P2_U2393);
  nand ginst16053 (P2_U6484, P2_R2099_U98, P2_U2379);
  nand ginst16054 (P2_U6485, P2_EBX_REG_4__SCAN_IN, P2_U3543);
  nand ginst16055 (P2_U6486, P2_R2182_U74, P2_U2393);
  nand ginst16056 (P2_U6487, P2_R2099_U71, P2_U2379);
  nand ginst16057 (P2_U6488, P2_EBX_REG_5__SCAN_IN, P2_U3543);
  nand ginst16058 (P2_U6489, P2_R2182_U73, P2_U2393);
  nand ginst16059 (P2_U6490, P2_R2099_U70, P2_U2379);
  nand ginst16060 (P2_U6491, P2_EBX_REG_6__SCAN_IN, P2_U3543);
  nand ginst16061 (P2_U6492, P2_R2182_U72, P2_U2393);
  nand ginst16062 (P2_U6493, P2_R2099_U69, P2_U2379);
  nand ginst16063 (P2_U6494, P2_EBX_REG_7__SCAN_IN, P2_U3543);
  nand ginst16064 (P2_U6495, P2_R2182_U71, P2_U2393);
  nand ginst16065 (P2_U6496, P2_R2099_U68, P2_U2379);
  nand ginst16066 (P2_U6497, P2_EBX_REG_8__SCAN_IN, P2_U3543);
  nand ginst16067 (P2_U6498, P2_R2182_U70, P2_U2393);
  nand ginst16068 (P2_U6499, P2_R2099_U67, P2_U2379);
  nand ginst16069 (P2_U6500, P2_EBX_REG_9__SCAN_IN, P2_U3543);
  nand ginst16070 (P2_U6501, P2_R2182_U96, P2_U2393);
  nand ginst16071 (P2_U6502, P2_R2099_U93, P2_U2379);
  nand ginst16072 (P2_U6503, P2_EBX_REG_10__SCAN_IN, P2_U3543);
  nand ginst16073 (P2_U6504, P2_R2182_U95, P2_U2393);
  nand ginst16074 (P2_U6505, P2_R2099_U92, P2_U2379);
  nand ginst16075 (P2_U6506, P2_EBX_REG_11__SCAN_IN, P2_U3543);
  nand ginst16076 (P2_U6507, P2_R2182_U94, P2_U2393);
  nand ginst16077 (P2_U6508, P2_R2099_U91, P2_U2379);
  nand ginst16078 (P2_U6509, P2_EBX_REG_12__SCAN_IN, P2_U3543);
  nand ginst16079 (P2_U6510, P2_R2182_U93, P2_U2393);
  nand ginst16080 (P2_U6511, P2_R2099_U90, P2_U2379);
  nand ginst16081 (P2_U6512, P2_EBX_REG_13__SCAN_IN, P2_U3543);
  nand ginst16082 (P2_U6513, P2_R2182_U92, P2_U2393);
  nand ginst16083 (P2_U6514, P2_R2099_U89, P2_U2379);
  nand ginst16084 (P2_U6515, P2_EBX_REG_14__SCAN_IN, P2_U3543);
  nand ginst16085 (P2_U6516, P2_R2182_U91, P2_U2393);
  nand ginst16086 (P2_U6517, P2_R2099_U88, P2_U2379);
  nand ginst16087 (P2_U6518, P2_EBX_REG_15__SCAN_IN, P2_U3543);
  nand ginst16088 (P2_U6519, P2_R2182_U90, P2_U2393);
  nand ginst16089 (P2_U6520, P2_R2099_U87, P2_U2379);
  nand ginst16090 (P2_U6521, P2_EBX_REG_16__SCAN_IN, P2_U3543);
  nand ginst16091 (P2_U6522, P2_R2182_U89, P2_U2393);
  nand ginst16092 (P2_U6523, P2_R2099_U86, P2_U2379);
  nand ginst16093 (P2_U6524, P2_EBX_REG_17__SCAN_IN, P2_U3543);
  nand ginst16094 (P2_U6525, P2_R2182_U88, P2_U2393);
  nand ginst16095 (P2_U6526, P2_R2099_U85, P2_U2379);
  nand ginst16096 (P2_U6527, P2_EBX_REG_18__SCAN_IN, P2_U3543);
  nand ginst16097 (P2_U6528, P2_R2182_U87, P2_U2393);
  nand ginst16098 (P2_U6529, P2_R2099_U84, P2_U2379);
  nand ginst16099 (P2_U6530, P2_EBX_REG_19__SCAN_IN, P2_U3543);
  nand ginst16100 (P2_U6531, P2_R2182_U86, P2_U2393);
  nand ginst16101 (P2_U6532, P2_R2099_U83, P2_U2379);
  nand ginst16102 (P2_U6533, P2_EBX_REG_20__SCAN_IN, P2_U3543);
  nand ginst16103 (P2_U6534, P2_R2182_U85, P2_U2393);
  nand ginst16104 (P2_U6535, P2_R2099_U82, P2_U2379);
  nand ginst16105 (P2_U6536, P2_EBX_REG_21__SCAN_IN, P2_U3543);
  nand ginst16106 (P2_U6537, P2_R2182_U84, P2_U2393);
  nand ginst16107 (P2_U6538, P2_R2099_U81, P2_U2379);
  nand ginst16108 (P2_U6539, P2_EBX_REG_22__SCAN_IN, P2_U3543);
  nand ginst16109 (P2_U6540, P2_R2182_U83, P2_U2393);
  nand ginst16110 (P2_U6541, P2_R2099_U80, P2_U2379);
  nand ginst16111 (P2_U6542, P2_EBX_REG_23__SCAN_IN, P2_U3543);
  nand ginst16112 (P2_U6543, P2_R2182_U82, P2_U2393);
  nand ginst16113 (P2_U6544, P2_R2099_U79, P2_U2379);
  nand ginst16114 (P2_U6545, P2_EBX_REG_24__SCAN_IN, P2_U3543);
  nand ginst16115 (P2_U6546, P2_R2182_U81, P2_U2393);
  nand ginst16116 (P2_U6547, P2_R2099_U78, P2_U2379);
  nand ginst16117 (P2_U6548, P2_EBX_REG_25__SCAN_IN, P2_U3543);
  nand ginst16118 (P2_U6549, P2_R2182_U80, P2_U2393);
  nand ginst16119 (P2_U6550, P2_R2099_U77, P2_U2379);
  nand ginst16120 (P2_U6551, P2_EBX_REG_26__SCAN_IN, P2_U3543);
  nand ginst16121 (P2_U6552, P2_R2182_U79, P2_U2393);
  nand ginst16122 (P2_U6553, P2_R2099_U76, P2_U2379);
  nand ginst16123 (P2_U6554, P2_EBX_REG_27__SCAN_IN, P2_U3543);
  nand ginst16124 (P2_U6555, P2_R2182_U78, P2_U2393);
  nand ginst16125 (P2_U6556, P2_R2099_U75, P2_U2379);
  nand ginst16126 (P2_U6557, P2_EBX_REG_28__SCAN_IN, P2_U3543);
  nand ginst16127 (P2_U6558, P2_R2182_U77, P2_U2393);
  nand ginst16128 (P2_U6559, P2_R2099_U74, P2_U2379);
  nand ginst16129 (P2_U6560, P2_EBX_REG_29__SCAN_IN, P2_U3543);
  nand ginst16130 (P2_U6561, P2_R2182_U41, P2_U2393);
  nand ginst16131 (P2_U6562, P2_R2099_U73, P2_U2379);
  nand ginst16132 (P2_U6563, P2_EBX_REG_30__SCAN_IN, P2_U3543);
  nand ginst16133 (P2_U6564, P2_R2099_U72, P2_U2379);
  nand ginst16134 (P2_U6565, P2_EBX_REG_31__SCAN_IN, P2_U3543);
  nand ginst16135 (P2_U6566, P2_R2088_U6, P2_U4603);
  nand ginst16136 (P2_U6567, P2_R2167_U6, P2_U4433);
  nand ginst16137 (P2_U6568, P2_U6566, P2_U6567);
  nand ginst16138 (P2_U6569, P2_U3284, P2_U4461);
  not ginst16139 (P2_U6570, P2_U3546);
  not ginst16140 (P2_U6571, P2_U3545);
  or ginst16141 (P2_U6572, P2_STATEBS16_REG_SCAN_IN, U211);
  nand ginst16142 (P2_U6573, P2_R2267_U21, P2_U2587);
  nand ginst16143 (P2_U6574, P2_R2096_U68, P2_U2588);
  nand ginst16144 (P2_U6575, P2_EBX_REG_0__SCAN_IN, P2_U7743);
  nand ginst16145 (P2_U6576, P2_R2182_U69, P2_U2437);
  nand ginst16146 (P2_U6577, P2_R2099_U94, P2_U2392);
  nand ginst16147 (P2_U6578, P2_PHYADDRPOINTER_REG_0__SCAN_IN, P2_U2383);
  nand ginst16148 (P2_U6579, P2_U2382, P2_U3683);
  nand ginst16149 (P2_U6580, P2_PHYADDRPOINTER_REG_0__SCAN_IN, P2_U2378);
  nand ginst16150 (P2_U6581, P2_REIP_REG_0__SCAN_IN, P2_U6570);
  nand ginst16151 (P2_U6582, P2_R2267_U43, P2_U2587);
  nand ginst16152 (P2_U6583, P2_R2096_U51, P2_U2588);
  nand ginst16153 (P2_U6584, P2_EBX_REG_1__SCAN_IN, P2_U7743);
  nand ginst16154 (P2_U6585, P2_R2182_U68, P2_U2437);
  nand ginst16155 (P2_U6586, P2_R2099_U5, P2_U2392);
  nand ginst16156 (P2_U6587, P2_R2337_U4, P2_U2383);
  nand ginst16157 (P2_U6588, P2_R1957_U49, P2_U2382);
  nand ginst16158 (P2_U6589, P2_PHYADDRPOINTER_REG_1__SCAN_IN, P2_U2378);
  nand ginst16159 (P2_U6590, P2_REIP_REG_1__SCAN_IN, P2_U6570);
  nand ginst16160 (P2_U6591, P2_R2267_U65, P2_U2587);
  nand ginst16161 (P2_U6592, P2_R2096_U77, P2_U2588);
  nand ginst16162 (P2_U6593, P2_EBX_REG_2__SCAN_IN, P2_U7743);
  nand ginst16163 (P2_U6594, P2_R2182_U40, P2_U2437);
  nand ginst16164 (P2_U6595, P2_R2099_U96, P2_U2392);
  nand ginst16165 (P2_U6596, P2_R2337_U70, P2_U2383);
  nand ginst16166 (P2_U6597, P2_R1957_U17, P2_U2382);
  nand ginst16167 (P2_U6598, P2_PHYADDRPOINTER_REG_2__SCAN_IN, P2_U2378);
  nand ginst16168 (P2_U6599, P2_REIP_REG_2__SCAN_IN, P2_U6570);
  nand ginst16169 (P2_U6600, P2_R2267_U17, P2_U2587);
  nand ginst16170 (P2_U6601, P2_R2096_U75, P2_U2588);
  nand ginst16171 (P2_U6602, P2_EBX_REG_3__SCAN_IN, P2_U7743);
  nand ginst16172 (P2_U6603, P2_R2182_U76, P2_U2437);
  nand ginst16173 (P2_U6604, P2_R2099_U95, P2_U2392);
  nand ginst16174 (P2_U6605, P2_R2337_U67, P2_U2383);
  nand ginst16175 (P2_U6606, P2_R1957_U59, P2_U2382);
  nand ginst16176 (P2_U6607, P2_PHYADDRPOINTER_REG_3__SCAN_IN, P2_U2378);
  nand ginst16177 (P2_U6608, P2_REIP_REG_3__SCAN_IN, P2_U6570);
  nand ginst16178 (P2_U6609, P2_R2267_U60, P2_U2587);
  nand ginst16179 (P2_U6610, P2_R2096_U74, P2_U2588);
  nand ginst16180 (P2_U6611, P2_EBX_REG_4__SCAN_IN, P2_U7743);
  nand ginst16181 (P2_U6612, P2_R2182_U75, P2_U2437);
  nand ginst16182 (P2_U6613, P2_R2099_U98, P2_U2392);
  nand ginst16183 (P2_U6614, P2_R2337_U66, P2_U2383);
  nand ginst16184 (P2_U6615, P2_R1957_U18, P2_U2382);
  nand ginst16185 (P2_U6616, P2_PHYADDRPOINTER_REG_4__SCAN_IN, P2_U2378);
  nand ginst16186 (P2_U6617, P2_REIP_REG_4__SCAN_IN, P2_U6570);
  nand ginst16187 (P2_U6618, P2_R2267_U18, P2_U2587);
  nand ginst16188 (P2_U6619, P2_R2096_U73, P2_U2588);
  nand ginst16189 (P2_U6620, P2_EBX_REG_5__SCAN_IN, P2_U7743);
  nand ginst16190 (P2_U6621, P2_R2182_U74, P2_U2437);
  nand ginst16191 (P2_U6622, P2_R2099_U71, P2_U2392);
  nand ginst16192 (P2_U6623, P2_R2337_U65, P2_U2383);
  nand ginst16193 (P2_U6624, P2_R1957_U57, P2_U2382);
  nand ginst16194 (P2_U6625, P2_PHYADDRPOINTER_REG_5__SCAN_IN, P2_U2378);
  nand ginst16195 (P2_U6626, P2_REIP_REG_5__SCAN_IN, P2_U6570);
  nand ginst16196 (P2_U6627, P2_R2267_U58, P2_U2587);
  nand ginst16197 (P2_U6628, P2_R2096_U72, P2_U2588);
  nand ginst16198 (P2_U6629, P2_EBX_REG_6__SCAN_IN, P2_U7743);
  nand ginst16199 (P2_U6630, P2_R2099_U70, P2_U2392);
  nand ginst16200 (P2_U6631, P2_R2337_U64, P2_U2383);
  nand ginst16201 (P2_U6632, P2_R1957_U19, P2_U2382);
  nand ginst16202 (P2_U6633, P2_PHYADDRPOINTER_REG_6__SCAN_IN, P2_U2378);
  nand ginst16203 (P2_U6634, P2_REIP_REG_6__SCAN_IN, P2_U6570);
  nand ginst16204 (P2_U6635, P2_R2267_U19, P2_U2587);
  nand ginst16205 (P2_U6636, P2_R2096_U71, P2_U2588);
  nand ginst16206 (P2_U6637, P2_EBX_REG_7__SCAN_IN, P2_U7743);
  nand ginst16207 (P2_U6638, P2_R2099_U69, P2_U2392);
  nand ginst16208 (P2_U6639, P2_R2337_U63, P2_U2383);
  nand ginst16209 (P2_U6640, P2_R1957_U55, P2_U2382);
  nand ginst16210 (P2_U6641, P2_PHYADDRPOINTER_REG_7__SCAN_IN, P2_U2378);
  nand ginst16211 (P2_U6642, P2_REIP_REG_7__SCAN_IN, P2_U6570);
  nand ginst16212 (P2_U6643, P2_R2267_U56, P2_U2587);
  nand ginst16213 (P2_U6644, P2_R2096_U70, P2_U2588);
  nand ginst16214 (P2_U6645, P2_EBX_REG_8__SCAN_IN, P2_U7743);
  nand ginst16215 (P2_U6646, P2_R2099_U68, P2_U2392);
  nand ginst16216 (P2_U6647, P2_R2337_U62, P2_U2383);
  nand ginst16217 (P2_U6648, P2_R1957_U20, P2_U2382);
  nand ginst16218 (P2_U6649, P2_PHYADDRPOINTER_REG_8__SCAN_IN, P2_U2378);
  nand ginst16219 (P2_U6650, P2_REIP_REG_8__SCAN_IN, P2_U6570);
  nand ginst16220 (P2_U6651, P2_R2267_U20, P2_U2587);
  nand ginst16221 (P2_U6652, P2_R2096_U69, P2_U2588);
  nand ginst16222 (P2_U6653, P2_EBX_REG_9__SCAN_IN, P2_U7743);
  nand ginst16223 (P2_U6654, P2_R2099_U67, P2_U2392);
  nand ginst16224 (P2_U6655, P2_R2337_U61, P2_U2383);
  nand ginst16225 (P2_U6656, P2_R1957_U53, P2_U2382);
  nand ginst16226 (P2_U6657, P2_PHYADDRPOINTER_REG_9__SCAN_IN, P2_U2378);
  nand ginst16227 (P2_U6658, P2_REIP_REG_9__SCAN_IN, P2_U6570);
  nand ginst16228 (P2_U6659, P2_R2267_U87, P2_U2587);
  nand ginst16229 (P2_U6660, P2_R2096_U97, P2_U2588);
  nand ginst16230 (P2_U6661, P2_EBX_REG_10__SCAN_IN, P2_U7743);
  nand ginst16231 (P2_U6662, P2_R2099_U93, P2_U2392);
  nand ginst16232 (P2_U6663, P2_R2337_U90, P2_U2383);
  nand ginst16233 (P2_U6664, P2_R1957_U6, P2_U2382);
  nand ginst16234 (P2_U6665, P2_PHYADDRPOINTER_REG_10__SCAN_IN, P2_U2378);
  nand ginst16235 (P2_U6666, P2_REIP_REG_10__SCAN_IN, P2_U6570);
  nand ginst16236 (P2_U6667, P2_R2267_U6, P2_U2587);
  nand ginst16237 (P2_U6668, P2_R2096_U96, P2_U2588);
  nand ginst16238 (P2_U6669, P2_EBX_REG_11__SCAN_IN, P2_U7743);
  nand ginst16239 (P2_U6670, P2_R2099_U92, P2_U2392);
  nand ginst16240 (P2_U6671, P2_R2337_U89, P2_U2383);
  nand ginst16241 (P2_U6672, P2_R1957_U82, P2_U2382);
  nand ginst16242 (P2_U6673, P2_PHYADDRPOINTER_REG_11__SCAN_IN, P2_U2378);
  nand ginst16243 (P2_U6674, P2_REIP_REG_11__SCAN_IN, P2_U6570);
  nand ginst16244 (P2_U6675, P2_R2267_U85, P2_U2587);
  nand ginst16245 (P2_U6676, P2_R2096_U95, P2_U2588);
  nand ginst16246 (P2_U6677, P2_EBX_REG_12__SCAN_IN, P2_U7743);
  nand ginst16247 (P2_U6678, P2_R2099_U91, P2_U2392);
  nand ginst16248 (P2_U6679, P2_R2337_U88, P2_U2383);
  nand ginst16249 (P2_U6680, P2_R1957_U7, P2_U2382);
  nand ginst16250 (P2_U6681, P2_PHYADDRPOINTER_REG_12__SCAN_IN, P2_U2378);
  nand ginst16251 (P2_U6682, P2_REIP_REG_12__SCAN_IN, P2_U6570);
  nand ginst16252 (P2_U6683, P2_R2267_U7, P2_U2587);
  nand ginst16253 (P2_U6684, P2_R2096_U94, P2_U2588);
  nand ginst16254 (P2_U6685, P2_EBX_REG_13__SCAN_IN, P2_U7743);
  nand ginst16255 (P2_U6686, P2_R2099_U90, P2_U2392);
  nand ginst16256 (P2_U6687, P2_R2337_U87, P2_U2383);
  nand ginst16257 (P2_U6688, P2_R1957_U80, P2_U2382);
  nand ginst16258 (P2_U6689, P2_PHYADDRPOINTER_REG_13__SCAN_IN, P2_U2378);
  nand ginst16259 (P2_U6690, P2_REIP_REG_13__SCAN_IN, P2_U6570);
  nand ginst16260 (P2_U6691, P2_R2267_U83, P2_U2587);
  nand ginst16261 (P2_U6692, P2_R2096_U93, P2_U2588);
  nand ginst16262 (P2_U6693, P2_EBX_REG_14__SCAN_IN, P2_U7743);
  nand ginst16263 (P2_U6694, P2_R2099_U89, P2_U2392);
  nand ginst16264 (P2_U6695, P2_R2337_U86, P2_U2383);
  nand ginst16265 (P2_U6696, P2_R1957_U8, P2_U2382);
  nand ginst16266 (P2_U6697, P2_PHYADDRPOINTER_REG_14__SCAN_IN, P2_U2378);
  nand ginst16267 (P2_U6698, P2_REIP_REG_14__SCAN_IN, P2_U6570);
  nand ginst16268 (P2_U6699, P2_R2267_U8, P2_U2587);
  nand ginst16269 (P2_U6700, P2_R2096_U92, P2_U2588);
  nand ginst16270 (P2_U6701, P2_EBX_REG_15__SCAN_IN, P2_U7743);
  nand ginst16271 (P2_U6702, P2_R2099_U88, P2_U2392);
  nand ginst16272 (P2_U6703, P2_R2337_U85, P2_U2383);
  nand ginst16273 (P2_U6704, P2_R1957_U78, P2_U2382);
  nand ginst16274 (P2_U6705, P2_PHYADDRPOINTER_REG_15__SCAN_IN, P2_U2378);
  nand ginst16275 (P2_U6706, P2_REIP_REG_15__SCAN_IN, P2_U6570);
  nand ginst16276 (P2_U6707, P2_R2267_U81, P2_U2587);
  nand ginst16277 (P2_U6708, P2_R2096_U91, P2_U2588);
  nand ginst16278 (P2_U6709, P2_EBX_REG_16__SCAN_IN, P2_U7743);
  nand ginst16279 (P2_U6710, P2_R2099_U87, P2_U2392);
  nand ginst16280 (P2_U6711, P2_R2337_U84, P2_U2383);
  nand ginst16281 (P2_U6712, P2_R1957_U9, P2_U2382);
  nand ginst16282 (P2_U6713, P2_PHYADDRPOINTER_REG_16__SCAN_IN, P2_U2378);
  nand ginst16283 (P2_U6714, P2_REIP_REG_16__SCAN_IN, P2_U6570);
  nand ginst16284 (P2_U6715, P2_R2267_U9, P2_U2587);
  nand ginst16285 (P2_U6716, P2_R2096_U90, P2_U2588);
  nand ginst16286 (P2_U6717, P2_EBX_REG_17__SCAN_IN, P2_U7743);
  nand ginst16287 (P2_U6718, P2_R2099_U86, P2_U2392);
  nand ginst16288 (P2_U6719, P2_R2337_U83, P2_U2383);
  nand ginst16289 (P2_U6720, P2_R1957_U76, P2_U2382);
  nand ginst16290 (P2_U6721, P2_PHYADDRPOINTER_REG_17__SCAN_IN, P2_U2378);
  nand ginst16291 (P2_U6722, P2_REIP_REG_17__SCAN_IN, P2_U6570);
  nand ginst16292 (P2_U6723, P2_R2267_U79, P2_U2587);
  nand ginst16293 (P2_U6724, P2_R2096_U89, P2_U2588);
  nand ginst16294 (P2_U6725, P2_EBX_REG_18__SCAN_IN, P2_U7743);
  nand ginst16295 (P2_U6726, P2_R2099_U85, P2_U2392);
  nand ginst16296 (P2_U6727, P2_R2337_U82, P2_U2383);
  nand ginst16297 (P2_U6728, P2_R1957_U10, P2_U2382);
  nand ginst16298 (P2_U6729, P2_PHYADDRPOINTER_REG_18__SCAN_IN, P2_U2378);
  nand ginst16299 (P2_U6730, P2_REIP_REG_18__SCAN_IN, P2_U6570);
  nand ginst16300 (P2_U6731, P2_R2267_U10, P2_U2587);
  nand ginst16301 (P2_U6732, P2_R2096_U88, P2_U2588);
  nand ginst16302 (P2_U6733, P2_EBX_REG_19__SCAN_IN, P2_U7743);
  nand ginst16303 (P2_U6734, P2_R2099_U84, P2_U2392);
  nand ginst16304 (P2_U6735, P2_R2337_U81, P2_U2383);
  nand ginst16305 (P2_U6736, P2_R1957_U74, P2_U2382);
  nand ginst16306 (P2_U6737, P2_PHYADDRPOINTER_REG_19__SCAN_IN, P2_U2378);
  nand ginst16307 (P2_U6738, P2_REIP_REG_19__SCAN_IN, P2_U6570);
  nand ginst16308 (P2_U6739, P2_R2267_U75, P2_U2587);
  nand ginst16309 (P2_U6740, P2_R2096_U87, P2_U2588);
  nand ginst16310 (P2_U6741, P2_EBX_REG_20__SCAN_IN, P2_U7743);
  nand ginst16311 (P2_U6742, P2_R2099_U83, P2_U2392);
  nand ginst16312 (P2_U6743, P2_R2337_U80, P2_U2383);
  nand ginst16313 (P2_U6744, P2_R1957_U11, P2_U2382);
  nand ginst16314 (P2_U6745, P2_PHYADDRPOINTER_REG_20__SCAN_IN, P2_U2378);
  nand ginst16315 (P2_U6746, P2_REIP_REG_20__SCAN_IN, P2_U6570);
  nand ginst16316 (P2_U6747, P2_R2267_U11, P2_U2587);
  nand ginst16317 (P2_U6748, P2_R2096_U86, P2_U2588);
  nand ginst16318 (P2_U6749, P2_EBX_REG_21__SCAN_IN, P2_U7743);
  nand ginst16319 (P2_U6750, P2_R2099_U82, P2_U2392);
  nand ginst16320 (P2_U6751, P2_R2337_U79, P2_U2383);
  nand ginst16321 (P2_U6752, P2_R1957_U70, P2_U2382);
  nand ginst16322 (P2_U6753, P2_PHYADDRPOINTER_REG_21__SCAN_IN, P2_U2378);
  nand ginst16323 (P2_U6754, P2_REIP_REG_21__SCAN_IN, P2_U6570);
  nand ginst16324 (P2_U6755, P2_R2267_U73, P2_U2587);
  nand ginst16325 (P2_U6756, P2_R2096_U85, P2_U2588);
  nand ginst16326 (P2_U6757, P2_EBX_REG_22__SCAN_IN, P2_U7743);
  nand ginst16327 (P2_U6758, P2_R2099_U81, P2_U2392);
  nand ginst16328 (P2_U6759, P2_R2337_U78, P2_U2383);
  nand ginst16329 (P2_U6760, P2_R1957_U12, P2_U2382);
  nand ginst16330 (P2_U6761, P2_PHYADDRPOINTER_REG_22__SCAN_IN, P2_U2378);
  nand ginst16331 (P2_U6762, P2_REIP_REG_22__SCAN_IN, P2_U6570);
  nand ginst16332 (P2_U6763, P2_R2267_U12, P2_U2587);
  nand ginst16333 (P2_U6764, P2_R2096_U84, P2_U2588);
  nand ginst16334 (P2_U6765, P2_EBX_REG_23__SCAN_IN, P2_U7743);
  nand ginst16335 (P2_U6766, P2_R2099_U80, P2_U2392);
  nand ginst16336 (P2_U6767, P2_R2337_U77, P2_U2383);
  nand ginst16337 (P2_U6768, P2_R1957_U68, P2_U2382);
  nand ginst16338 (P2_U6769, P2_PHYADDRPOINTER_REG_23__SCAN_IN, P2_U2378);
  nand ginst16339 (P2_U6770, P2_REIP_REG_23__SCAN_IN, P2_U6570);
  nand ginst16340 (P2_U6771, P2_R2267_U71, P2_U2587);
  nand ginst16341 (P2_U6772, P2_R2096_U83, P2_U2588);
  nand ginst16342 (P2_U6773, P2_EBX_REG_24__SCAN_IN, P2_U7743);
  nand ginst16343 (P2_U6774, P2_R2099_U79, P2_U2392);
  nand ginst16344 (P2_U6775, P2_R2337_U76, P2_U2383);
  nand ginst16345 (P2_U6776, P2_R1957_U13, P2_U2382);
  nand ginst16346 (P2_U6777, P2_PHYADDRPOINTER_REG_24__SCAN_IN, P2_U2378);
  nand ginst16347 (P2_U6778, P2_REIP_REG_24__SCAN_IN, P2_U6570);
  nand ginst16348 (P2_U6779, P2_R2267_U13, P2_U2587);
  nand ginst16349 (P2_U6780, P2_R2096_U82, P2_U2588);
  nand ginst16350 (P2_U6781, P2_EBX_REG_25__SCAN_IN, P2_U7743);
  nand ginst16351 (P2_U6782, P2_R2099_U78, P2_U2392);
  nand ginst16352 (P2_U6783, P2_R2337_U75, P2_U2383);
  nand ginst16353 (P2_U6784, P2_R1957_U66, P2_U2382);
  nand ginst16354 (P2_U6785, P2_PHYADDRPOINTER_REG_25__SCAN_IN, P2_U2378);
  nand ginst16355 (P2_U6786, P2_REIP_REG_25__SCAN_IN, P2_U6570);
  nand ginst16356 (P2_U6787, P2_R2267_U69, P2_U2587);
  nand ginst16357 (P2_U6788, P2_R2096_U81, P2_U2588);
  nand ginst16358 (P2_U6789, P2_EBX_REG_26__SCAN_IN, P2_U7743);
  nand ginst16359 (P2_U6790, P2_R2099_U77, P2_U2392);
  nand ginst16360 (P2_U6791, P2_R2337_U74, P2_U2383);
  nand ginst16361 (P2_U6792, P2_R1957_U14, P2_U2382);
  nand ginst16362 (P2_U6793, P2_PHYADDRPOINTER_REG_26__SCAN_IN, P2_U2378);
  nand ginst16363 (P2_U6794, P2_REIP_REG_26__SCAN_IN, P2_U6570);
  nand ginst16364 (P2_U6795, P2_R2267_U14, P2_U2587);
  nand ginst16365 (P2_U6796, P2_R2096_U80, P2_U2588);
  nand ginst16366 (P2_U6797, P2_EBX_REG_27__SCAN_IN, P2_U7743);
  nand ginst16367 (P2_U6798, P2_R2099_U76, P2_U2392);
  nand ginst16368 (P2_U6799, P2_R2337_U73, P2_U2383);
  nand ginst16369 (P2_U6800, P2_R1957_U64, P2_U2382);
  nand ginst16370 (P2_U6801, P2_PHYADDRPOINTER_REG_27__SCAN_IN, P2_U2378);
  nand ginst16371 (P2_U6802, P2_REIP_REG_27__SCAN_IN, P2_U6570);
  nand ginst16372 (P2_U6803, P2_R2267_U67, P2_U2587);
  nand ginst16373 (P2_U6804, P2_R2096_U79, P2_U2588);
  nand ginst16374 (P2_U6805, P2_EBX_REG_28__SCAN_IN, P2_U7743);
  nand ginst16375 (P2_U6806, P2_R2099_U75, P2_U2392);
  nand ginst16376 (P2_U6807, P2_R2337_U72, P2_U2383);
  nand ginst16377 (P2_U6808, P2_R1957_U15, P2_U2382);
  nand ginst16378 (P2_U6809, P2_PHYADDRPOINTER_REG_28__SCAN_IN, P2_U2378);
  nand ginst16379 (P2_U6810, P2_REIP_REG_28__SCAN_IN, P2_U6570);
  nand ginst16380 (P2_U6811, P2_R2267_U15, P2_U2587);
  nand ginst16381 (P2_U6812, P2_R2096_U78, P2_U2588);
  nand ginst16382 (P2_U6813, P2_EBX_REG_29__SCAN_IN, P2_U7743);
  nand ginst16383 (P2_U6814, P2_R2099_U74, P2_U2392);
  nand ginst16384 (P2_U6815, P2_R2337_U71, P2_U2383);
  nand ginst16385 (P2_U6816, P2_R1957_U16, P2_U2382);
  nand ginst16386 (P2_U6817, P2_PHYADDRPOINTER_REG_29__SCAN_IN, P2_U2378);
  nand ginst16387 (P2_U6818, P2_REIP_REG_29__SCAN_IN, P2_U6570);
  nand ginst16388 (P2_U6819, P2_R2267_U16, P2_U2587);
  nand ginst16389 (P2_U6820, P2_R2096_U76, P2_U2588);
  nand ginst16390 (P2_U6821, P2_EBX_REG_30__SCAN_IN, P2_U7743);
  nand ginst16391 (P2_U6822, P2_R2099_U73, P2_U2392);
  nand ginst16392 (P2_U6823, P2_R2337_U69, P2_U2383);
  nand ginst16393 (P2_U6824, P2_R1957_U62, P2_U2382);
  nand ginst16394 (P2_U6825, P2_PHYADDRPOINTER_REG_30__SCAN_IN, P2_U2378);
  nand ginst16395 (P2_U6826, P2_REIP_REG_30__SCAN_IN, P2_U6570);
  nand ginst16396 (P2_U6827, P2_R2267_U63, P2_U2587);
  nand ginst16397 (P2_U6828, P2_R2096_U50, P2_U2588);
  nand ginst16398 (P2_U6829, P2_EBX_REG_31__SCAN_IN, P2_U7743);
  nand ginst16399 (P2_U6830, P2_R2099_U72, P2_U2392);
  nand ginst16400 (P2_U6831, P2_R2337_U68, P2_U2383);
  nand ginst16401 (P2_U6832, P2_R1957_U50, P2_U2382);
  nand ginst16402 (P2_U6833, P2_PHYADDRPOINTER_REG_31__SCAN_IN, P2_U2378);
  nand ginst16403 (P2_U6834, P2_REIP_REG_31__SCAN_IN, P2_U6570);
  nand ginst16404 (P2_U6835, P2_DATAWIDTH_REG_0__SCAN_IN, P2_DATAWIDTH_REG_1__SCAN_IN);
  nand ginst16405 (P2_U6836, P2_REIP_REG_0__SCAN_IN, P2_U4477);
  nand ginst16406 (P2_U6837, P2_BYTEENABLE_REG_1__SCAN_IN, P2_U3547);
  not ginst16407 (P2_U6838, P2_U4400);
  nand ginst16408 (P2_U6839, P2_U4399, P2_U4426, P2_U4468);
  nand ginst16409 (P2_U6840, P2_FLUSH_REG_SCAN_IN, P2_U4400);
  nand ginst16410 (P2_U6841, P2_U4187, P2_U4467);
  nand ginst16411 (P2_U6842, P2_U3284, P2_U4466);
  not ginst16412 (P2_U6843, P2_U4402);
  nand ginst16413 (P2_U6844, P2_STATEBS16_REG_SCAN_IN, P2_U4411);
  not ginst16414 (P2_U6845, P2_U2715);
  nand ginst16415 (P2_U6846, P2_U2715, P2_U3536);
  nand ginst16416 (P2_U6847, P2_U3265, P2_U4411);
  nand ginst16417 (P2_U6848, P2_U2356, P2_U4184);
  nand ginst16418 (P2_U6849, P2_U4418, P2_U6847);
  nand ginst16419 (P2_U6850, P2_U6846, U211);
  or ginst16420 (P2_U6851, P2_STATE2_REG_2__SCAN_IN, P2_STATE2_REG_1__SCAN_IN);
  nand ginst16421 (P2_U6852, P2_U4186, P2_U6850, P2_U6851);
  nand ginst16422 (P2_U6853, P2_U2374, P2_U2459);
  nand ginst16423 (P2_U6854, P2_CODEFETCH_REG_SCAN_IN, P2_U6853);
  nand ginst16424 (P2_U6855, P2_STATE2_REG_0__SCAN_IN, P2_U4461);
  nand ginst16425 (P2_U6856, P2_STATE_REG_0__SCAN_IN, P2_ADS_N_REG_SCAN_IN);
  not ginst16426 (P2_U6857, P2_U4403);
  nand ginst16427 (P2_U6858, P2_STATE2_REG_2__SCAN_IN, P2_U3286, P2_U3294);
  nand ginst16428 (P2_U6859, P2_U4404, P2_U4421, P2_U4468);
  nand ginst16429 (P2_U6860, P2_U2446, P2_U4189);
  nand ginst16430 (P2_U6861, P2_MEMORYFETCH_REG_SCAN_IN, P2_U6859);
  nand ginst16431 (P2_U6862, P2_INSTQUEUE_REG_8__7__SCAN_IN, P2_U2538);
  nand ginst16432 (P2_U6863, P2_INSTQUEUE_REG_9__7__SCAN_IN, P2_U2537);
  nand ginst16433 (P2_U6864, P2_INSTQUEUE_REG_10__7__SCAN_IN, P2_U2536);
  nand ginst16434 (P2_U6865, P2_INSTQUEUE_REG_11__7__SCAN_IN, P2_U2535);
  nand ginst16435 (P2_U6866, P2_INSTQUEUE_REG_12__7__SCAN_IN, P2_U2534);
  nand ginst16436 (P2_U6867, P2_INSTQUEUE_REG_13__7__SCAN_IN, P2_U2533);
  nand ginst16437 (P2_U6868, P2_INSTQUEUE_REG_14__7__SCAN_IN, P2_U2531);
  nand ginst16438 (P2_U6869, P2_INSTQUEUE_REG_15__7__SCAN_IN, P2_U2530);
  nand ginst16439 (P2_U6870, P2_INSTQUEUE_REG_7__7__SCAN_IN, P2_U2528);
  nand ginst16440 (P2_U6871, P2_INSTQUEUE_REG_6__7__SCAN_IN, P2_U2527);
  nand ginst16441 (P2_U6872, P2_INSTQUEUE_REG_5__7__SCAN_IN, P2_U2526);
  nand ginst16442 (P2_U6873, P2_INSTQUEUE_REG_4__7__SCAN_IN, P2_U2524);
  nand ginst16443 (P2_U6874, P2_INSTQUEUE_REG_3__7__SCAN_IN, P2_U2522);
  nand ginst16444 (P2_U6875, P2_INSTQUEUE_REG_2__7__SCAN_IN, P2_U2521);
  nand ginst16445 (P2_U6876, P2_INSTQUEUE_REG_1__7__SCAN_IN, P2_U2519);
  nand ginst16446 (P2_U6877, P2_INSTQUEUE_REG_0__7__SCAN_IN, P2_U2517);
  nand ginst16447 (P2_U6878, P2_INSTQUEUE_REG_15__7__SCAN_IN, P2_U2562);
  nand ginst16448 (P2_U6879, P2_INSTQUEUE_REG_14__7__SCAN_IN, P2_U2561);
  nand ginst16449 (P2_U6880, P2_INSTQUEUE_REG_13__7__SCAN_IN, P2_U2560);
  nand ginst16450 (P2_U6881, P2_INSTQUEUE_REG_12__7__SCAN_IN, P2_U2559);
  nand ginst16451 (P2_U6882, P2_INSTQUEUE_REG_11__7__SCAN_IN, P2_U2558);
  nand ginst16452 (P2_U6883, P2_INSTQUEUE_REG_10__7__SCAN_IN, P2_U2557);
  nand ginst16453 (P2_U6884, P2_INSTQUEUE_REG_9__7__SCAN_IN, P2_U2555);
  nand ginst16454 (P2_U6885, P2_INSTQUEUE_REG_8__7__SCAN_IN, P2_U2554);
  nand ginst16455 (P2_U6886, P2_INSTQUEUE_REG_7__7__SCAN_IN, P2_U2552);
  nand ginst16456 (P2_U6887, P2_INSTQUEUE_REG_6__7__SCAN_IN, P2_U2551);
  nand ginst16457 (P2_U6888, P2_INSTQUEUE_REG_5__7__SCAN_IN, P2_U2550);
  nand ginst16458 (P2_U6889, P2_INSTQUEUE_REG_4__7__SCAN_IN, P2_U2548);
  nand ginst16459 (P2_U6890, P2_INSTQUEUE_REG_3__7__SCAN_IN, P2_U2546);
  nand ginst16460 (P2_U6891, P2_INSTQUEUE_REG_2__7__SCAN_IN, P2_U2545);
  nand ginst16461 (P2_U6892, P2_INSTQUEUE_REG_1__7__SCAN_IN, P2_U2543);
  nand ginst16462 (P2_U6893, P2_INSTQUEUE_REG_0__7__SCAN_IN, P2_U2541);
  nand ginst16463 (P2_U6894, P2_INSTQUEUE_REG_15__6__SCAN_IN, P2_U2562);
  nand ginst16464 (P2_U6895, P2_INSTQUEUE_REG_14__6__SCAN_IN, P2_U2561);
  nand ginst16465 (P2_U6896, P2_INSTQUEUE_REG_13__6__SCAN_IN, P2_U2560);
  nand ginst16466 (P2_U6897, P2_INSTQUEUE_REG_12__6__SCAN_IN, P2_U2559);
  nand ginst16467 (P2_U6898, P2_INSTQUEUE_REG_11__6__SCAN_IN, P2_U2558);
  nand ginst16468 (P2_U6899, P2_INSTQUEUE_REG_10__6__SCAN_IN, P2_U2557);
  nand ginst16469 (P2_U6900, P2_INSTQUEUE_REG_9__6__SCAN_IN, P2_U2555);
  nand ginst16470 (P2_U6901, P2_INSTQUEUE_REG_8__6__SCAN_IN, P2_U2554);
  nand ginst16471 (P2_U6902, P2_INSTQUEUE_REG_7__6__SCAN_IN, P2_U2552);
  nand ginst16472 (P2_U6903, P2_INSTQUEUE_REG_6__6__SCAN_IN, P2_U2551);
  nand ginst16473 (P2_U6904, P2_INSTQUEUE_REG_5__6__SCAN_IN, P2_U2550);
  nand ginst16474 (P2_U6905, P2_INSTQUEUE_REG_4__6__SCAN_IN, P2_U2548);
  nand ginst16475 (P2_U6906, P2_INSTQUEUE_REG_3__6__SCAN_IN, P2_U2546);
  nand ginst16476 (P2_U6907, P2_INSTQUEUE_REG_2__6__SCAN_IN, P2_U2545);
  nand ginst16477 (P2_U6908, P2_INSTQUEUE_REG_1__6__SCAN_IN, P2_U2543);
  nand ginst16478 (P2_U6909, P2_INSTQUEUE_REG_0__6__SCAN_IN, P2_U2541);
  nand ginst16479 (P2_U6910, P2_INSTQUEUE_REG_15__5__SCAN_IN, P2_U2562);
  nand ginst16480 (P2_U6911, P2_INSTQUEUE_REG_14__5__SCAN_IN, P2_U2561);
  nand ginst16481 (P2_U6912, P2_INSTQUEUE_REG_13__5__SCAN_IN, P2_U2560);
  nand ginst16482 (P2_U6913, P2_INSTQUEUE_REG_12__5__SCAN_IN, P2_U2559);
  nand ginst16483 (P2_U6914, P2_INSTQUEUE_REG_11__5__SCAN_IN, P2_U2558);
  nand ginst16484 (P2_U6915, P2_INSTQUEUE_REG_10__5__SCAN_IN, P2_U2557);
  nand ginst16485 (P2_U6916, P2_INSTQUEUE_REG_9__5__SCAN_IN, P2_U2555);
  nand ginst16486 (P2_U6917, P2_INSTQUEUE_REG_8__5__SCAN_IN, P2_U2554);
  nand ginst16487 (P2_U6918, P2_INSTQUEUE_REG_7__5__SCAN_IN, P2_U2552);
  nand ginst16488 (P2_U6919, P2_INSTQUEUE_REG_6__5__SCAN_IN, P2_U2551);
  nand ginst16489 (P2_U6920, P2_INSTQUEUE_REG_5__5__SCAN_IN, P2_U2550);
  nand ginst16490 (P2_U6921, P2_INSTQUEUE_REG_4__5__SCAN_IN, P2_U2548);
  nand ginst16491 (P2_U6922, P2_INSTQUEUE_REG_3__5__SCAN_IN, P2_U2546);
  nand ginst16492 (P2_U6923, P2_INSTQUEUE_REG_2__5__SCAN_IN, P2_U2545);
  nand ginst16493 (P2_U6924, P2_INSTQUEUE_REG_1__5__SCAN_IN, P2_U2543);
  nand ginst16494 (P2_U6925, P2_INSTQUEUE_REG_0__5__SCAN_IN, P2_U2541);
  nand ginst16495 (P2_U6926, P2_INSTQUEUE_REG_15__4__SCAN_IN, P2_U2562);
  nand ginst16496 (P2_U6927, P2_INSTQUEUE_REG_14__4__SCAN_IN, P2_U2561);
  nand ginst16497 (P2_U6928, P2_INSTQUEUE_REG_13__4__SCAN_IN, P2_U2560);
  nand ginst16498 (P2_U6929, P2_INSTQUEUE_REG_12__4__SCAN_IN, P2_U2559);
  nand ginst16499 (P2_U6930, P2_INSTQUEUE_REG_11__4__SCAN_IN, P2_U2558);
  nand ginst16500 (P2_U6931, P2_INSTQUEUE_REG_10__4__SCAN_IN, P2_U2557);
  nand ginst16501 (P2_U6932, P2_INSTQUEUE_REG_9__4__SCAN_IN, P2_U2555);
  nand ginst16502 (P2_U6933, P2_INSTQUEUE_REG_8__4__SCAN_IN, P2_U2554);
  nand ginst16503 (P2_U6934, P2_INSTQUEUE_REG_7__4__SCAN_IN, P2_U2552);
  nand ginst16504 (P2_U6935, P2_INSTQUEUE_REG_6__4__SCAN_IN, P2_U2551);
  nand ginst16505 (P2_U6936, P2_INSTQUEUE_REG_5__4__SCAN_IN, P2_U2550);
  nand ginst16506 (P2_U6937, P2_INSTQUEUE_REG_4__4__SCAN_IN, P2_U2548);
  nand ginst16507 (P2_U6938, P2_INSTQUEUE_REG_3__4__SCAN_IN, P2_U2546);
  nand ginst16508 (P2_U6939, P2_INSTQUEUE_REG_2__4__SCAN_IN, P2_U2545);
  nand ginst16509 (P2_U6940, P2_INSTQUEUE_REG_1__4__SCAN_IN, P2_U2543);
  nand ginst16510 (P2_U6941, P2_INSTQUEUE_REG_0__4__SCAN_IN, P2_U2541);
  nand ginst16511 (P2_U6942, P2_INSTQUEUE_REG_15__3__SCAN_IN, P2_U2562);
  nand ginst16512 (P2_U6943, P2_INSTQUEUE_REG_14__3__SCAN_IN, P2_U2561);
  nand ginst16513 (P2_U6944, P2_INSTQUEUE_REG_13__3__SCAN_IN, P2_U2560);
  nand ginst16514 (P2_U6945, P2_INSTQUEUE_REG_12__3__SCAN_IN, P2_U2559);
  nand ginst16515 (P2_U6946, P2_INSTQUEUE_REG_11__3__SCAN_IN, P2_U2558);
  nand ginst16516 (P2_U6947, P2_INSTQUEUE_REG_10__3__SCAN_IN, P2_U2557);
  nand ginst16517 (P2_U6948, P2_INSTQUEUE_REG_9__3__SCAN_IN, P2_U2555);
  nand ginst16518 (P2_U6949, P2_INSTQUEUE_REG_8__3__SCAN_IN, P2_U2554);
  nand ginst16519 (P2_U6950, P2_INSTQUEUE_REG_7__3__SCAN_IN, P2_U2552);
  nand ginst16520 (P2_U6951, P2_INSTQUEUE_REG_6__3__SCAN_IN, P2_U2551);
  nand ginst16521 (P2_U6952, P2_INSTQUEUE_REG_5__3__SCAN_IN, P2_U2550);
  nand ginst16522 (P2_U6953, P2_INSTQUEUE_REG_4__3__SCAN_IN, P2_U2548);
  nand ginst16523 (P2_U6954, P2_INSTQUEUE_REG_3__3__SCAN_IN, P2_U2546);
  nand ginst16524 (P2_U6955, P2_INSTQUEUE_REG_2__3__SCAN_IN, P2_U2545);
  nand ginst16525 (P2_U6956, P2_INSTQUEUE_REG_1__3__SCAN_IN, P2_U2543);
  nand ginst16526 (P2_U6957, P2_INSTQUEUE_REG_0__3__SCAN_IN, P2_U2541);
  nand ginst16527 (P2_U6958, P2_INSTQUEUE_REG_15__2__SCAN_IN, P2_U2562);
  nand ginst16528 (P2_U6959, P2_INSTQUEUE_REG_14__2__SCAN_IN, P2_U2561);
  nand ginst16529 (P2_U6960, P2_INSTQUEUE_REG_13__2__SCAN_IN, P2_U2560);
  nand ginst16530 (P2_U6961, P2_INSTQUEUE_REG_12__2__SCAN_IN, P2_U2559);
  nand ginst16531 (P2_U6962, P2_INSTQUEUE_REG_11__2__SCAN_IN, P2_U2558);
  nand ginst16532 (P2_U6963, P2_INSTQUEUE_REG_10__2__SCAN_IN, P2_U2557);
  nand ginst16533 (P2_U6964, P2_INSTQUEUE_REG_9__2__SCAN_IN, P2_U2555);
  nand ginst16534 (P2_U6965, P2_INSTQUEUE_REG_8__2__SCAN_IN, P2_U2554);
  nand ginst16535 (P2_U6966, P2_INSTQUEUE_REG_7__2__SCAN_IN, P2_U2552);
  nand ginst16536 (P2_U6967, P2_INSTQUEUE_REG_6__2__SCAN_IN, P2_U2551);
  nand ginst16537 (P2_U6968, P2_INSTQUEUE_REG_5__2__SCAN_IN, P2_U2550);
  nand ginst16538 (P2_U6969, P2_INSTQUEUE_REG_4__2__SCAN_IN, P2_U2548);
  nand ginst16539 (P2_U6970, P2_INSTQUEUE_REG_3__2__SCAN_IN, P2_U2546);
  nand ginst16540 (P2_U6971, P2_INSTQUEUE_REG_2__2__SCAN_IN, P2_U2545);
  nand ginst16541 (P2_U6972, P2_INSTQUEUE_REG_1__2__SCAN_IN, P2_U2543);
  nand ginst16542 (P2_U6973, P2_INSTQUEUE_REG_0__2__SCAN_IN, P2_U2541);
  nand ginst16543 (P2_U6974, P2_INSTQUEUE_REG_15__1__SCAN_IN, P2_U2562);
  nand ginst16544 (P2_U6975, P2_INSTQUEUE_REG_14__1__SCAN_IN, P2_U2561);
  nand ginst16545 (P2_U6976, P2_INSTQUEUE_REG_13__1__SCAN_IN, P2_U2560);
  nand ginst16546 (P2_U6977, P2_INSTQUEUE_REG_12__1__SCAN_IN, P2_U2559);
  nand ginst16547 (P2_U6978, P2_INSTQUEUE_REG_11__1__SCAN_IN, P2_U2558);
  nand ginst16548 (P2_U6979, P2_INSTQUEUE_REG_10__1__SCAN_IN, P2_U2557);
  nand ginst16549 (P2_U6980, P2_INSTQUEUE_REG_9__1__SCAN_IN, P2_U2555);
  nand ginst16550 (P2_U6981, P2_INSTQUEUE_REG_8__1__SCAN_IN, P2_U2554);
  nand ginst16551 (P2_U6982, P2_INSTQUEUE_REG_7__1__SCAN_IN, P2_U2552);
  nand ginst16552 (P2_U6983, P2_INSTQUEUE_REG_6__1__SCAN_IN, P2_U2551);
  nand ginst16553 (P2_U6984, P2_INSTQUEUE_REG_5__1__SCAN_IN, P2_U2550);
  nand ginst16554 (P2_U6985, P2_INSTQUEUE_REG_4__1__SCAN_IN, P2_U2548);
  nand ginst16555 (P2_U6986, P2_INSTQUEUE_REG_3__1__SCAN_IN, P2_U2546);
  nand ginst16556 (P2_U6987, P2_INSTQUEUE_REG_2__1__SCAN_IN, P2_U2545);
  nand ginst16557 (P2_U6988, P2_INSTQUEUE_REG_1__1__SCAN_IN, P2_U2543);
  nand ginst16558 (P2_U6989, P2_INSTQUEUE_REG_0__1__SCAN_IN, P2_U2541);
  nand ginst16559 (P2_U6990, P2_INSTQUEUE_REG_15__0__SCAN_IN, P2_U2562);
  nand ginst16560 (P2_U6991, P2_INSTQUEUE_REG_14__0__SCAN_IN, P2_U2561);
  nand ginst16561 (P2_U6992, P2_INSTQUEUE_REG_13__0__SCAN_IN, P2_U2560);
  nand ginst16562 (P2_U6993, P2_INSTQUEUE_REG_12__0__SCAN_IN, P2_U2559);
  nand ginst16563 (P2_U6994, P2_INSTQUEUE_REG_11__0__SCAN_IN, P2_U2558);
  nand ginst16564 (P2_U6995, P2_INSTQUEUE_REG_10__0__SCAN_IN, P2_U2557);
  nand ginst16565 (P2_U6996, P2_INSTQUEUE_REG_9__0__SCAN_IN, P2_U2555);
  nand ginst16566 (P2_U6997, P2_INSTQUEUE_REG_8__0__SCAN_IN, P2_U2554);
  nand ginst16567 (P2_U6998, P2_INSTQUEUE_REG_7__0__SCAN_IN, P2_U2552);
  nand ginst16568 (P2_U6999, P2_INSTQUEUE_REG_6__0__SCAN_IN, P2_U2551);
  nand ginst16569 (P2_U7000, P2_INSTQUEUE_REG_5__0__SCAN_IN, P2_U2550);
  nand ginst16570 (P2_U7001, P2_INSTQUEUE_REG_4__0__SCAN_IN, P2_U2548);
  nand ginst16571 (P2_U7002, P2_INSTQUEUE_REG_3__0__SCAN_IN, P2_U2546);
  nand ginst16572 (P2_U7003, P2_INSTQUEUE_REG_2__0__SCAN_IN, P2_U2545);
  nand ginst16573 (P2_U7004, P2_INSTQUEUE_REG_1__0__SCAN_IN, P2_U2543);
  nand ginst16574 (P2_U7005, P2_INSTQUEUE_REG_0__0__SCAN_IN, P2_U2541);
  or ginst16575 (P2_U7006, P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN);
  not ginst16576 (P2_U7007, P2_U4405);
  nand ginst16577 (P2_U7008, P2_INSTQUEUE_REG_0__7__SCAN_IN, P2_U2586);
  nand ginst16578 (P2_U7009, P2_INSTQUEUE_REG_1__7__SCAN_IN, P2_U2585);
  nand ginst16579 (P2_U7010, P2_INSTQUEUE_REG_2__7__SCAN_IN, P2_U2584);
  nand ginst16580 (P2_U7011, P2_INSTQUEUE_REG_3__7__SCAN_IN, P2_U2583);
  nand ginst16581 (P2_U7012, P2_INSTQUEUE_REG_4__7__SCAN_IN, P2_U2581);
  nand ginst16582 (P2_U7013, P2_INSTQUEUE_REG_5__7__SCAN_IN, P2_U2580);
  nand ginst16583 (P2_U7014, P2_INSTQUEUE_REG_6__7__SCAN_IN, P2_U2579);
  nand ginst16584 (P2_U7015, P2_INSTQUEUE_REG_7__7__SCAN_IN, P2_U2578);
  nand ginst16585 (P2_U7016, P2_INSTQUEUE_REG_8__7__SCAN_IN, P2_U2576);
  nand ginst16586 (P2_U7017, P2_INSTQUEUE_REG_9__7__SCAN_IN, P2_U2575);
  nand ginst16587 (P2_U7018, P2_INSTQUEUE_REG_10__7__SCAN_IN, P2_U2574);
  nand ginst16588 (P2_U7019, P2_INSTQUEUE_REG_11__7__SCAN_IN, P2_U2573);
  nand ginst16589 (P2_U7020, P2_INSTQUEUE_REG_12__7__SCAN_IN, P2_U2571);
  nand ginst16590 (P2_U7021, P2_INSTQUEUE_REG_13__7__SCAN_IN, P2_U2569);
  nand ginst16591 (P2_U7022, P2_INSTQUEUE_REG_14__7__SCAN_IN, P2_U2567);
  nand ginst16592 (P2_U7023, P2_INSTQUEUE_REG_15__7__SCAN_IN, P2_U2565);
  nand ginst16593 (P2_U7024, P2_INSTQUEUE_REG_0__6__SCAN_IN, P2_U2586);
  nand ginst16594 (P2_U7025, P2_INSTQUEUE_REG_1__6__SCAN_IN, P2_U2585);
  nand ginst16595 (P2_U7026, P2_INSTQUEUE_REG_2__6__SCAN_IN, P2_U2584);
  nand ginst16596 (P2_U7027, P2_INSTQUEUE_REG_3__6__SCAN_IN, P2_U2583);
  nand ginst16597 (P2_U7028, P2_INSTQUEUE_REG_4__6__SCAN_IN, P2_U2581);
  nand ginst16598 (P2_U7029, P2_INSTQUEUE_REG_5__6__SCAN_IN, P2_U2580);
  nand ginst16599 (P2_U7030, P2_INSTQUEUE_REG_6__6__SCAN_IN, P2_U2579);
  nand ginst16600 (P2_U7031, P2_INSTQUEUE_REG_7__6__SCAN_IN, P2_U2578);
  nand ginst16601 (P2_U7032, P2_INSTQUEUE_REG_8__6__SCAN_IN, P2_U2576);
  nand ginst16602 (P2_U7033, P2_INSTQUEUE_REG_9__6__SCAN_IN, P2_U2575);
  nand ginst16603 (P2_U7034, P2_INSTQUEUE_REG_10__6__SCAN_IN, P2_U2574);
  nand ginst16604 (P2_U7035, P2_INSTQUEUE_REG_11__6__SCAN_IN, P2_U2573);
  nand ginst16605 (P2_U7036, P2_INSTQUEUE_REG_12__6__SCAN_IN, P2_U2571);
  nand ginst16606 (P2_U7037, P2_INSTQUEUE_REG_13__6__SCAN_IN, P2_U2569);
  nand ginst16607 (P2_U7038, P2_INSTQUEUE_REG_14__6__SCAN_IN, P2_U2567);
  nand ginst16608 (P2_U7039, P2_INSTQUEUE_REG_15__6__SCAN_IN, P2_U2565);
  nand ginst16609 (P2_U7040, P2_INSTQUEUE_REG_0__5__SCAN_IN, P2_U2586);
  nand ginst16610 (P2_U7041, P2_INSTQUEUE_REG_1__5__SCAN_IN, P2_U2585);
  nand ginst16611 (P2_U7042, P2_INSTQUEUE_REG_2__5__SCAN_IN, P2_U2584);
  nand ginst16612 (P2_U7043, P2_INSTQUEUE_REG_3__5__SCAN_IN, P2_U2583);
  nand ginst16613 (P2_U7044, P2_INSTQUEUE_REG_4__5__SCAN_IN, P2_U2581);
  nand ginst16614 (P2_U7045, P2_INSTQUEUE_REG_5__5__SCAN_IN, P2_U2580);
  nand ginst16615 (P2_U7046, P2_INSTQUEUE_REG_6__5__SCAN_IN, P2_U2579);
  nand ginst16616 (P2_U7047, P2_INSTQUEUE_REG_7__5__SCAN_IN, P2_U2578);
  nand ginst16617 (P2_U7048, P2_INSTQUEUE_REG_8__5__SCAN_IN, P2_U2576);
  nand ginst16618 (P2_U7049, P2_INSTQUEUE_REG_9__5__SCAN_IN, P2_U2575);
  nand ginst16619 (P2_U7050, P2_INSTQUEUE_REG_10__5__SCAN_IN, P2_U2574);
  nand ginst16620 (P2_U7051, P2_INSTQUEUE_REG_11__5__SCAN_IN, P2_U2573);
  nand ginst16621 (P2_U7052, P2_INSTQUEUE_REG_12__5__SCAN_IN, P2_U2571);
  nand ginst16622 (P2_U7053, P2_INSTQUEUE_REG_13__5__SCAN_IN, P2_U2569);
  nand ginst16623 (P2_U7054, P2_INSTQUEUE_REG_14__5__SCAN_IN, P2_U2567);
  nand ginst16624 (P2_U7055, P2_INSTQUEUE_REG_15__5__SCAN_IN, P2_U2565);
  nand ginst16625 (P2_U7056, P2_INSTQUEUE_REG_0__4__SCAN_IN, P2_U2586);
  nand ginst16626 (P2_U7057, P2_INSTQUEUE_REG_1__4__SCAN_IN, P2_U2585);
  nand ginst16627 (P2_U7058, P2_INSTQUEUE_REG_2__4__SCAN_IN, P2_U2584);
  nand ginst16628 (P2_U7059, P2_INSTQUEUE_REG_3__4__SCAN_IN, P2_U2583);
  nand ginst16629 (P2_U7060, P2_INSTQUEUE_REG_4__4__SCAN_IN, P2_U2581);
  nand ginst16630 (P2_U7061, P2_INSTQUEUE_REG_5__4__SCAN_IN, P2_U2580);
  nand ginst16631 (P2_U7062, P2_INSTQUEUE_REG_6__4__SCAN_IN, P2_U2579);
  nand ginst16632 (P2_U7063, P2_INSTQUEUE_REG_7__4__SCAN_IN, P2_U2578);
  nand ginst16633 (P2_U7064, P2_INSTQUEUE_REG_8__4__SCAN_IN, P2_U2576);
  nand ginst16634 (P2_U7065, P2_INSTQUEUE_REG_9__4__SCAN_IN, P2_U2575);
  nand ginst16635 (P2_U7066, P2_INSTQUEUE_REG_10__4__SCAN_IN, P2_U2574);
  nand ginst16636 (P2_U7067, P2_INSTQUEUE_REG_11__4__SCAN_IN, P2_U2573);
  nand ginst16637 (P2_U7068, P2_INSTQUEUE_REG_12__4__SCAN_IN, P2_U2571);
  nand ginst16638 (P2_U7069, P2_INSTQUEUE_REG_13__4__SCAN_IN, P2_U2569);
  nand ginst16639 (P2_U7070, P2_INSTQUEUE_REG_14__4__SCAN_IN, P2_U2567);
  nand ginst16640 (P2_U7071, P2_INSTQUEUE_REG_15__4__SCAN_IN, P2_U2565);
  nand ginst16641 (P2_U7072, P2_INSTQUEUE_REG_0__3__SCAN_IN, P2_U2586);
  nand ginst16642 (P2_U7073, P2_INSTQUEUE_REG_1__3__SCAN_IN, P2_U2585);
  nand ginst16643 (P2_U7074, P2_INSTQUEUE_REG_2__3__SCAN_IN, P2_U2584);
  nand ginst16644 (P2_U7075, P2_INSTQUEUE_REG_3__3__SCAN_IN, P2_U2583);
  nand ginst16645 (P2_U7076, P2_INSTQUEUE_REG_4__3__SCAN_IN, P2_U2581);
  nand ginst16646 (P2_U7077, P2_INSTQUEUE_REG_5__3__SCAN_IN, P2_U2580);
  nand ginst16647 (P2_U7078, P2_INSTQUEUE_REG_6__3__SCAN_IN, P2_U2579);
  nand ginst16648 (P2_U7079, P2_INSTQUEUE_REG_7__3__SCAN_IN, P2_U2578);
  nand ginst16649 (P2_U7080, P2_INSTQUEUE_REG_8__3__SCAN_IN, P2_U2576);
  nand ginst16650 (P2_U7081, P2_INSTQUEUE_REG_9__3__SCAN_IN, P2_U2575);
  nand ginst16651 (P2_U7082, P2_INSTQUEUE_REG_10__3__SCAN_IN, P2_U2574);
  nand ginst16652 (P2_U7083, P2_INSTQUEUE_REG_11__3__SCAN_IN, P2_U2573);
  nand ginst16653 (P2_U7084, P2_INSTQUEUE_REG_12__3__SCAN_IN, P2_U2571);
  nand ginst16654 (P2_U7085, P2_INSTQUEUE_REG_13__3__SCAN_IN, P2_U2569);
  nand ginst16655 (P2_U7086, P2_INSTQUEUE_REG_14__3__SCAN_IN, P2_U2567);
  nand ginst16656 (P2_U7087, P2_INSTQUEUE_REG_15__3__SCAN_IN, P2_U2565);
  nand ginst16657 (P2_U7088, P2_INSTQUEUE_REG_0__2__SCAN_IN, P2_U2586);
  nand ginst16658 (P2_U7089, P2_INSTQUEUE_REG_1__2__SCAN_IN, P2_U2585);
  nand ginst16659 (P2_U7090, P2_INSTQUEUE_REG_2__2__SCAN_IN, P2_U2584);
  nand ginst16660 (P2_U7091, P2_INSTQUEUE_REG_3__2__SCAN_IN, P2_U2583);
  nand ginst16661 (P2_U7092, P2_INSTQUEUE_REG_4__2__SCAN_IN, P2_U2581);
  nand ginst16662 (P2_U7093, P2_INSTQUEUE_REG_5__2__SCAN_IN, P2_U2580);
  nand ginst16663 (P2_U7094, P2_INSTQUEUE_REG_6__2__SCAN_IN, P2_U2579);
  nand ginst16664 (P2_U7095, P2_INSTQUEUE_REG_7__2__SCAN_IN, P2_U2578);
  nand ginst16665 (P2_U7096, P2_INSTQUEUE_REG_8__2__SCAN_IN, P2_U2576);
  nand ginst16666 (P2_U7097, P2_INSTQUEUE_REG_9__2__SCAN_IN, P2_U2575);
  nand ginst16667 (P2_U7098, P2_INSTQUEUE_REG_10__2__SCAN_IN, P2_U2574);
  nand ginst16668 (P2_U7099, P2_INSTQUEUE_REG_11__2__SCAN_IN, P2_U2573);
  nand ginst16669 (P2_U7100, P2_INSTQUEUE_REG_12__2__SCAN_IN, P2_U2571);
  nand ginst16670 (P2_U7101, P2_INSTQUEUE_REG_13__2__SCAN_IN, P2_U2569);
  nand ginst16671 (P2_U7102, P2_INSTQUEUE_REG_14__2__SCAN_IN, P2_U2567);
  nand ginst16672 (P2_U7103, P2_INSTQUEUE_REG_15__2__SCAN_IN, P2_U2565);
  nand ginst16673 (P2_U7104, P2_INSTQUEUE_REG_0__1__SCAN_IN, P2_U2586);
  nand ginst16674 (P2_U7105, P2_INSTQUEUE_REG_1__1__SCAN_IN, P2_U2585);
  nand ginst16675 (P2_U7106, P2_INSTQUEUE_REG_2__1__SCAN_IN, P2_U2584);
  nand ginst16676 (P2_U7107, P2_INSTQUEUE_REG_3__1__SCAN_IN, P2_U2583);
  nand ginst16677 (P2_U7108, P2_INSTQUEUE_REG_4__1__SCAN_IN, P2_U2581);
  nand ginst16678 (P2_U7109, P2_INSTQUEUE_REG_5__1__SCAN_IN, P2_U2580);
  nand ginst16679 (P2_U7110, P2_INSTQUEUE_REG_6__1__SCAN_IN, P2_U2579);
  nand ginst16680 (P2_U7111, P2_INSTQUEUE_REG_7__1__SCAN_IN, P2_U2578);
  nand ginst16681 (P2_U7112, P2_INSTQUEUE_REG_8__1__SCAN_IN, P2_U2576);
  nand ginst16682 (P2_U7113, P2_INSTQUEUE_REG_9__1__SCAN_IN, P2_U2575);
  nand ginst16683 (P2_U7114, P2_INSTQUEUE_REG_10__1__SCAN_IN, P2_U2574);
  nand ginst16684 (P2_U7115, P2_INSTQUEUE_REG_11__1__SCAN_IN, P2_U2573);
  nand ginst16685 (P2_U7116, P2_INSTQUEUE_REG_12__1__SCAN_IN, P2_U2571);
  nand ginst16686 (P2_U7117, P2_INSTQUEUE_REG_13__1__SCAN_IN, P2_U2569);
  nand ginst16687 (P2_U7118, P2_INSTQUEUE_REG_14__1__SCAN_IN, P2_U2567);
  nand ginst16688 (P2_U7119, P2_INSTQUEUE_REG_15__1__SCAN_IN, P2_U2565);
  nand ginst16689 (P2_U7120, P2_INSTQUEUE_REG_0__0__SCAN_IN, P2_U2586);
  nand ginst16690 (P2_U7121, P2_INSTQUEUE_REG_1__0__SCAN_IN, P2_U2585);
  nand ginst16691 (P2_U7122, P2_INSTQUEUE_REG_2__0__SCAN_IN, P2_U2584);
  nand ginst16692 (P2_U7123, P2_INSTQUEUE_REG_3__0__SCAN_IN, P2_U2583);
  nand ginst16693 (P2_U7124, P2_INSTQUEUE_REG_4__0__SCAN_IN, P2_U2581);
  nand ginst16694 (P2_U7125, P2_INSTQUEUE_REG_5__0__SCAN_IN, P2_U2580);
  nand ginst16695 (P2_U7126, P2_INSTQUEUE_REG_6__0__SCAN_IN, P2_U2579);
  nand ginst16696 (P2_U7127, P2_INSTQUEUE_REG_7__0__SCAN_IN, P2_U2578);
  nand ginst16697 (P2_U7128, P2_INSTQUEUE_REG_8__0__SCAN_IN, P2_U2576);
  nand ginst16698 (P2_U7129, P2_INSTQUEUE_REG_9__0__SCAN_IN, P2_U2575);
  nand ginst16699 (P2_U7130, P2_INSTQUEUE_REG_10__0__SCAN_IN, P2_U2574);
  nand ginst16700 (P2_U7131, P2_INSTQUEUE_REG_11__0__SCAN_IN, P2_U2573);
  nand ginst16701 (P2_U7132, P2_INSTQUEUE_REG_12__0__SCAN_IN, P2_U2571);
  nand ginst16702 (P2_U7133, P2_INSTQUEUE_REG_13__0__SCAN_IN, P2_U2569);
  nand ginst16703 (P2_U7134, P2_INSTQUEUE_REG_14__0__SCAN_IN, P2_U2567);
  nand ginst16704 (P2_U7135, P2_INSTQUEUE_REG_15__0__SCAN_IN, P2_U2565);
  not ginst16705 (P2_U7136, P2_U3554);
  nand ginst16706 (P2_U7137, P2_U3300, P2_U7136);
  nand ginst16707 (P2_U7138, P2_R2099_U95, P2_U4467);
  nand ginst16708 (P2_U7139, P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P2_U7137);
  nand ginst16709 (P2_U7140, P2_U3428, P2_U4430);
  nand ginst16710 (P2_U7141, P2_ADD_402_1132_U23, P2_U2355);
  nand ginst16711 (P2_U7142, P2_U2354, P2_U2606);
  nand ginst16712 (P2_U7143, P2_U2355, P2_U2605);
  nand ginst16713 (P2_U7144, P2_U2354, P2_U2605);
  nand ginst16714 (P2_U7145, P2_U2355, P2_U2604);
  nand ginst16715 (P2_U7146, P2_U2354, P2_U2604);
  nand ginst16716 (P2_U7147, P2_U2355, P2_U2603);
  nand ginst16717 (P2_U7148, P2_U2354, P2_U2603);
  nand ginst16718 (P2_U7149, P2_R2099_U96, P2_U4467);
  nand ginst16719 (P2_U7150, P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN, P2_U7137);
  nand ginst16720 (P2_U7151, P2_U3580, P2_U4430);
  nand ginst16721 (P2_U7152, P2_U2355, P2_U2602);
  nand ginst16722 (P2_U7153, P2_U2354, P2_U2602);
  nand ginst16723 (P2_U7154, P2_U2355, P2_U2601);
  nand ginst16724 (P2_U7155, P2_U2354, P2_U2601);
  nand ginst16725 (P2_U7156, P2_U2355, P2_U2600);
  nand ginst16726 (P2_U7157, P2_U2354, P2_U2600);
  nand ginst16727 (P2_U7158, P2_U2355, P2_U2599);
  nand ginst16728 (P2_U7159, P2_U2354, P2_U2599);
  nand ginst16729 (P2_U7160, P2_R2099_U5, P2_U4467);
  nand ginst16730 (P2_U7161, P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P2_U7137);
  nand ginst16731 (P2_U7162, P2_U3243, P2_U4430);
  nand ginst16732 (P2_U7163, P2_R2099_U94, P2_U4467);
  nand ginst16733 (P2_U7164, P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN, P2_U7137);
  nand ginst16734 (P2_U7165, P2_U3307, P2_U4430);
  nand ginst16735 (P2_U7166, P2_INSTQUEUE_REG_0__0__SCAN_IN, P2_U2355);
  nand ginst16736 (P2_U7167, P2_INSTQUEUE_REG_0__7__SCAN_IN, P2_U5517);
  nand ginst16737 (P2_U7168, P2_INSTQUEUE_REG_1__7__SCAN_IN, P2_U5460);
  nand ginst16738 (P2_U7169, P2_INSTQUEUE_REG_2__7__SCAN_IN, P2_U5402);
  nand ginst16739 (P2_U7170, P2_INSTQUEUE_REG_3__7__SCAN_IN, P2_U5345);
  nand ginst16740 (P2_U7171, P2_INSTQUEUE_REG_4__7__SCAN_IN, P2_U5287);
  nand ginst16741 (P2_U7172, P2_INSTQUEUE_REG_5__7__SCAN_IN, P2_U5230);
  nand ginst16742 (P2_U7173, P2_INSTQUEUE_REG_6__7__SCAN_IN, P2_U5172);
  nand ginst16743 (P2_U7174, P2_INSTQUEUE_REG_7__7__SCAN_IN, P2_U5116);
  nand ginst16744 (P2_U7175, P2_INSTQUEUE_REG_8__7__SCAN_IN, P2_U5059);
  nand ginst16745 (P2_U7176, P2_INSTQUEUE_REG_9__7__SCAN_IN, P2_U5002);
  nand ginst16746 (P2_U7177, P2_INSTQUEUE_REG_10__7__SCAN_IN, P2_U4944);
  nand ginst16747 (P2_U7178, P2_INSTQUEUE_REG_11__7__SCAN_IN, P2_U4887);
  nand ginst16748 (P2_U7179, P2_INSTQUEUE_REG_12__7__SCAN_IN, P2_U4829);
  nand ginst16749 (P2_U7180, P2_INSTQUEUE_REG_13__7__SCAN_IN, P2_U4772);
  nand ginst16750 (P2_U7181, P2_INSTQUEUE_REG_14__7__SCAN_IN, P2_U4713);
  nand ginst16751 (P2_U7182, P2_INSTQUEUE_REG_15__7__SCAN_IN, P2_U4653);
  nand ginst16752 (P2_U7183, P2_U4277, P2_U4278, P2_U4279, P2_U4280);
  nand ginst16753 (P2_U7184, P2_INSTQUEUE_REG_0__6__SCAN_IN, P2_U5517);
  nand ginst16754 (P2_U7185, P2_INSTQUEUE_REG_1__6__SCAN_IN, P2_U5460);
  nand ginst16755 (P2_U7186, P2_INSTQUEUE_REG_2__6__SCAN_IN, P2_U5402);
  nand ginst16756 (P2_U7187, P2_INSTQUEUE_REG_3__6__SCAN_IN, P2_U5345);
  nand ginst16757 (P2_U7188, P2_INSTQUEUE_REG_4__6__SCAN_IN, P2_U5287);
  nand ginst16758 (P2_U7189, P2_INSTQUEUE_REG_5__6__SCAN_IN, P2_U5230);
  nand ginst16759 (P2_U7190, P2_INSTQUEUE_REG_6__6__SCAN_IN, P2_U5172);
  nand ginst16760 (P2_U7191, P2_INSTQUEUE_REG_7__6__SCAN_IN, P2_U5116);
  nand ginst16761 (P2_U7192, P2_INSTQUEUE_REG_8__6__SCAN_IN, P2_U5059);
  nand ginst16762 (P2_U7193, P2_INSTQUEUE_REG_9__6__SCAN_IN, P2_U5002);
  nand ginst16763 (P2_U7194, P2_INSTQUEUE_REG_10__6__SCAN_IN, P2_U4944);
  nand ginst16764 (P2_U7195, P2_INSTQUEUE_REG_11__6__SCAN_IN, P2_U4887);
  nand ginst16765 (P2_U7196, P2_INSTQUEUE_REG_12__6__SCAN_IN, P2_U4829);
  nand ginst16766 (P2_U7197, P2_INSTQUEUE_REG_13__6__SCAN_IN, P2_U4772);
  nand ginst16767 (P2_U7198, P2_INSTQUEUE_REG_14__6__SCAN_IN, P2_U4713);
  nand ginst16768 (P2_U7199, P2_INSTQUEUE_REG_15__6__SCAN_IN, P2_U4653);
  nand ginst16769 (P2_U7200, P2_U4281, P2_U4282, P2_U4283, P2_U4284);
  nand ginst16770 (P2_U7201, P2_INSTQUEUE_REG_8__6__SCAN_IN, P2_U2538);
  nand ginst16771 (P2_U7202, P2_INSTQUEUE_REG_9__6__SCAN_IN, P2_U2537);
  nand ginst16772 (P2_U7203, P2_INSTQUEUE_REG_10__6__SCAN_IN, P2_U2536);
  nand ginst16773 (P2_U7204, P2_INSTQUEUE_REG_11__6__SCAN_IN, P2_U2535);
  nand ginst16774 (P2_U7205, P2_INSTQUEUE_REG_12__6__SCAN_IN, P2_U2534);
  nand ginst16775 (P2_U7206, P2_INSTQUEUE_REG_13__6__SCAN_IN, P2_U2533);
  nand ginst16776 (P2_U7207, P2_INSTQUEUE_REG_14__6__SCAN_IN, P2_U2531);
  nand ginst16777 (P2_U7208, P2_INSTQUEUE_REG_15__6__SCAN_IN, P2_U2530);
  nand ginst16778 (P2_U7209, P2_INSTQUEUE_REG_7__6__SCAN_IN, P2_U2528);
  nand ginst16779 (P2_U7210, P2_INSTQUEUE_REG_6__6__SCAN_IN, P2_U2527);
  nand ginst16780 (P2_U7211, P2_INSTQUEUE_REG_5__6__SCAN_IN, P2_U2526);
  nand ginst16781 (P2_U7212, P2_INSTQUEUE_REG_4__6__SCAN_IN, P2_U2524);
  nand ginst16782 (P2_U7213, P2_INSTQUEUE_REG_3__6__SCAN_IN, P2_U2522);
  nand ginst16783 (P2_U7214, P2_INSTQUEUE_REG_2__6__SCAN_IN, P2_U2521);
  nand ginst16784 (P2_U7215, P2_INSTQUEUE_REG_1__6__SCAN_IN, P2_U2519);
  nand ginst16785 (P2_U7216, P2_INSTQUEUE_REG_0__6__SCAN_IN, P2_U2517);
  nand ginst16786 (P2_U7217, P2_U4285, P2_U4286, P2_U4287, P2_U4288);
  nand ginst16787 (P2_U7218, P2_INSTQUEUE_REG_0__5__SCAN_IN, P2_U5517);
  nand ginst16788 (P2_U7219, P2_INSTQUEUE_REG_1__5__SCAN_IN, P2_U5460);
  nand ginst16789 (P2_U7220, P2_INSTQUEUE_REG_2__5__SCAN_IN, P2_U5402);
  nand ginst16790 (P2_U7221, P2_INSTQUEUE_REG_3__5__SCAN_IN, P2_U5345);
  nand ginst16791 (P2_U7222, P2_INSTQUEUE_REG_4__5__SCAN_IN, P2_U5287);
  nand ginst16792 (P2_U7223, P2_INSTQUEUE_REG_5__5__SCAN_IN, P2_U5230);
  nand ginst16793 (P2_U7224, P2_INSTQUEUE_REG_6__5__SCAN_IN, P2_U5172);
  nand ginst16794 (P2_U7225, P2_INSTQUEUE_REG_7__5__SCAN_IN, P2_U5116);
  nand ginst16795 (P2_U7226, P2_INSTQUEUE_REG_8__5__SCAN_IN, P2_U5059);
  nand ginst16796 (P2_U7227, P2_INSTQUEUE_REG_9__5__SCAN_IN, P2_U5002);
  nand ginst16797 (P2_U7228, P2_INSTQUEUE_REG_10__5__SCAN_IN, P2_U4944);
  nand ginst16798 (P2_U7229, P2_INSTQUEUE_REG_11__5__SCAN_IN, P2_U4887);
  nand ginst16799 (P2_U7230, P2_INSTQUEUE_REG_12__5__SCAN_IN, P2_U4829);
  nand ginst16800 (P2_U7231, P2_INSTQUEUE_REG_13__5__SCAN_IN, P2_U4772);
  nand ginst16801 (P2_U7232, P2_INSTQUEUE_REG_14__5__SCAN_IN, P2_U4713);
  nand ginst16802 (P2_U7233, P2_INSTQUEUE_REG_15__5__SCAN_IN, P2_U4653);
  nand ginst16803 (P2_U7234, P2_U4289, P2_U4290, P2_U4291, P2_U4292);
  nand ginst16804 (P2_U7235, P2_INSTQUEUE_REG_8__5__SCAN_IN, P2_U2538);
  nand ginst16805 (P2_U7236, P2_INSTQUEUE_REG_9__5__SCAN_IN, P2_U2537);
  nand ginst16806 (P2_U7237, P2_INSTQUEUE_REG_10__5__SCAN_IN, P2_U2536);
  nand ginst16807 (P2_U7238, P2_INSTQUEUE_REG_11__5__SCAN_IN, P2_U2535);
  nand ginst16808 (P2_U7239, P2_INSTQUEUE_REG_12__5__SCAN_IN, P2_U2534);
  nand ginst16809 (P2_U7240, P2_INSTQUEUE_REG_13__5__SCAN_IN, P2_U2533);
  nand ginst16810 (P2_U7241, P2_INSTQUEUE_REG_14__5__SCAN_IN, P2_U2531);
  nand ginst16811 (P2_U7242, P2_INSTQUEUE_REG_15__5__SCAN_IN, P2_U2530);
  nand ginst16812 (P2_U7243, P2_INSTQUEUE_REG_7__5__SCAN_IN, P2_U2528);
  nand ginst16813 (P2_U7244, P2_INSTQUEUE_REG_6__5__SCAN_IN, P2_U2527);
  nand ginst16814 (P2_U7245, P2_INSTQUEUE_REG_5__5__SCAN_IN, P2_U2526);
  nand ginst16815 (P2_U7246, P2_INSTQUEUE_REG_4__5__SCAN_IN, P2_U2524);
  nand ginst16816 (P2_U7247, P2_INSTQUEUE_REG_3__5__SCAN_IN, P2_U2522);
  nand ginst16817 (P2_U7248, P2_INSTQUEUE_REG_2__5__SCAN_IN, P2_U2521);
  nand ginst16818 (P2_U7249, P2_INSTQUEUE_REG_1__5__SCAN_IN, P2_U2519);
  nand ginst16819 (P2_U7250, P2_INSTQUEUE_REG_0__5__SCAN_IN, P2_U2517);
  nand ginst16820 (P2_U7251, P2_U4293, P2_U4294, P2_U4295, P2_U4296);
  nand ginst16821 (P2_U7252, P2_INSTQUEUE_REG_0__4__SCAN_IN, P2_U5517);
  nand ginst16822 (P2_U7253, P2_INSTQUEUE_REG_1__4__SCAN_IN, P2_U5460);
  nand ginst16823 (P2_U7254, P2_INSTQUEUE_REG_2__4__SCAN_IN, P2_U5402);
  nand ginst16824 (P2_U7255, P2_INSTQUEUE_REG_3__4__SCAN_IN, P2_U5345);
  nand ginst16825 (P2_U7256, P2_INSTQUEUE_REG_4__4__SCAN_IN, P2_U5287);
  nand ginst16826 (P2_U7257, P2_INSTQUEUE_REG_5__4__SCAN_IN, P2_U5230);
  nand ginst16827 (P2_U7258, P2_INSTQUEUE_REG_6__4__SCAN_IN, P2_U5172);
  nand ginst16828 (P2_U7259, P2_INSTQUEUE_REG_7__4__SCAN_IN, P2_U5116);
  nand ginst16829 (P2_U7260, P2_INSTQUEUE_REG_8__4__SCAN_IN, P2_U5059);
  nand ginst16830 (P2_U7261, P2_INSTQUEUE_REG_9__4__SCAN_IN, P2_U5002);
  nand ginst16831 (P2_U7262, P2_INSTQUEUE_REG_10__4__SCAN_IN, P2_U4944);
  nand ginst16832 (P2_U7263, P2_INSTQUEUE_REG_11__4__SCAN_IN, P2_U4887);
  nand ginst16833 (P2_U7264, P2_INSTQUEUE_REG_12__4__SCAN_IN, P2_U4829);
  nand ginst16834 (P2_U7265, P2_INSTQUEUE_REG_13__4__SCAN_IN, P2_U4772);
  nand ginst16835 (P2_U7266, P2_INSTQUEUE_REG_14__4__SCAN_IN, P2_U4713);
  nand ginst16836 (P2_U7267, P2_INSTQUEUE_REG_15__4__SCAN_IN, P2_U4653);
  nand ginst16837 (P2_U7268, P2_U4297, P2_U4298, P2_U4299, P2_U4300);
  nand ginst16838 (P2_U7269, P2_INSTQUEUE_REG_8__4__SCAN_IN, P2_U2538);
  nand ginst16839 (P2_U7270, P2_INSTQUEUE_REG_9__4__SCAN_IN, P2_U2537);
  nand ginst16840 (P2_U7271, P2_INSTQUEUE_REG_10__4__SCAN_IN, P2_U2536);
  nand ginst16841 (P2_U7272, P2_INSTQUEUE_REG_11__4__SCAN_IN, P2_U2535);
  nand ginst16842 (P2_U7273, P2_INSTQUEUE_REG_12__4__SCAN_IN, P2_U2534);
  nand ginst16843 (P2_U7274, P2_INSTQUEUE_REG_13__4__SCAN_IN, P2_U2533);
  nand ginst16844 (P2_U7275, P2_INSTQUEUE_REG_14__4__SCAN_IN, P2_U2531);
  nand ginst16845 (P2_U7276, P2_INSTQUEUE_REG_15__4__SCAN_IN, P2_U2530);
  nand ginst16846 (P2_U7277, P2_INSTQUEUE_REG_7__4__SCAN_IN, P2_U2528);
  nand ginst16847 (P2_U7278, P2_INSTQUEUE_REG_6__4__SCAN_IN, P2_U2527);
  nand ginst16848 (P2_U7279, P2_INSTQUEUE_REG_5__4__SCAN_IN, P2_U2526);
  nand ginst16849 (P2_U7280, P2_INSTQUEUE_REG_4__4__SCAN_IN, P2_U2524);
  nand ginst16850 (P2_U7281, P2_INSTQUEUE_REG_3__4__SCAN_IN, P2_U2522);
  nand ginst16851 (P2_U7282, P2_INSTQUEUE_REG_2__4__SCAN_IN, P2_U2521);
  nand ginst16852 (P2_U7283, P2_INSTQUEUE_REG_1__4__SCAN_IN, P2_U2519);
  nand ginst16853 (P2_U7284, P2_INSTQUEUE_REG_0__4__SCAN_IN, P2_U2517);
  nand ginst16854 (P2_U7285, P2_U4301, P2_U4302, P2_U4303, P2_U4304);
  nand ginst16855 (P2_U7286, P2_INSTQUEUE_REG_0__3__SCAN_IN, P2_U5517);
  nand ginst16856 (P2_U7287, P2_INSTQUEUE_REG_1__3__SCAN_IN, P2_U5460);
  nand ginst16857 (P2_U7288, P2_INSTQUEUE_REG_2__3__SCAN_IN, P2_U5402);
  nand ginst16858 (P2_U7289, P2_INSTQUEUE_REG_3__3__SCAN_IN, P2_U5345);
  nand ginst16859 (P2_U7290, P2_INSTQUEUE_REG_4__3__SCAN_IN, P2_U5287);
  nand ginst16860 (P2_U7291, P2_INSTQUEUE_REG_5__3__SCAN_IN, P2_U5230);
  nand ginst16861 (P2_U7292, P2_INSTQUEUE_REG_6__3__SCAN_IN, P2_U5172);
  nand ginst16862 (P2_U7293, P2_INSTQUEUE_REG_7__3__SCAN_IN, P2_U5116);
  nand ginst16863 (P2_U7294, P2_INSTQUEUE_REG_8__3__SCAN_IN, P2_U5059);
  nand ginst16864 (P2_U7295, P2_INSTQUEUE_REG_9__3__SCAN_IN, P2_U5002);
  nand ginst16865 (P2_U7296, P2_INSTQUEUE_REG_10__3__SCAN_IN, P2_U4944);
  nand ginst16866 (P2_U7297, P2_INSTQUEUE_REG_11__3__SCAN_IN, P2_U4887);
  nand ginst16867 (P2_U7298, P2_INSTQUEUE_REG_12__3__SCAN_IN, P2_U4829);
  nand ginst16868 (P2_U7299, P2_INSTQUEUE_REG_13__3__SCAN_IN, P2_U4772);
  nand ginst16869 (P2_U7300, P2_INSTQUEUE_REG_14__3__SCAN_IN, P2_U4713);
  nand ginst16870 (P2_U7301, P2_INSTQUEUE_REG_15__3__SCAN_IN, P2_U4653);
  nand ginst16871 (P2_U7302, P2_U4305, P2_U4306, P2_U4307, P2_U4308);
  nand ginst16872 (P2_U7303, P2_INSTQUEUE_REG_8__3__SCAN_IN, P2_U2538);
  nand ginst16873 (P2_U7304, P2_INSTQUEUE_REG_9__3__SCAN_IN, P2_U2537);
  nand ginst16874 (P2_U7305, P2_INSTQUEUE_REG_10__3__SCAN_IN, P2_U2536);
  nand ginst16875 (P2_U7306, P2_INSTQUEUE_REG_11__3__SCAN_IN, P2_U2535);
  nand ginst16876 (P2_U7307, P2_INSTQUEUE_REG_12__3__SCAN_IN, P2_U2534);
  nand ginst16877 (P2_U7308, P2_INSTQUEUE_REG_13__3__SCAN_IN, P2_U2533);
  nand ginst16878 (P2_U7309, P2_INSTQUEUE_REG_14__3__SCAN_IN, P2_U2531);
  nand ginst16879 (P2_U7310, P2_INSTQUEUE_REG_15__3__SCAN_IN, P2_U2530);
  nand ginst16880 (P2_U7311, P2_INSTQUEUE_REG_7__3__SCAN_IN, P2_U2528);
  nand ginst16881 (P2_U7312, P2_INSTQUEUE_REG_6__3__SCAN_IN, P2_U2527);
  nand ginst16882 (P2_U7313, P2_INSTQUEUE_REG_5__3__SCAN_IN, P2_U2526);
  nand ginst16883 (P2_U7314, P2_INSTQUEUE_REG_4__3__SCAN_IN, P2_U2524);
  nand ginst16884 (P2_U7315, P2_INSTQUEUE_REG_3__3__SCAN_IN, P2_U2522);
  nand ginst16885 (P2_U7316, P2_INSTQUEUE_REG_2__3__SCAN_IN, P2_U2521);
  nand ginst16886 (P2_U7317, P2_INSTQUEUE_REG_1__3__SCAN_IN, P2_U2519);
  nand ginst16887 (P2_U7318, P2_INSTQUEUE_REG_0__3__SCAN_IN, P2_U2517);
  nand ginst16888 (P2_U7319, P2_U4309, P2_U4310, P2_U4311, P2_U4312);
  nand ginst16889 (P2_U7320, P2_INSTQUEUE_REG_0__2__SCAN_IN, P2_U5517);
  nand ginst16890 (P2_U7321, P2_INSTQUEUE_REG_1__2__SCAN_IN, P2_U5460);
  nand ginst16891 (P2_U7322, P2_INSTQUEUE_REG_2__2__SCAN_IN, P2_U5402);
  nand ginst16892 (P2_U7323, P2_INSTQUEUE_REG_3__2__SCAN_IN, P2_U5345);
  nand ginst16893 (P2_U7324, P2_INSTQUEUE_REG_4__2__SCAN_IN, P2_U5287);
  nand ginst16894 (P2_U7325, P2_INSTQUEUE_REG_5__2__SCAN_IN, P2_U5230);
  nand ginst16895 (P2_U7326, P2_INSTQUEUE_REG_6__2__SCAN_IN, P2_U5172);
  nand ginst16896 (P2_U7327, P2_INSTQUEUE_REG_7__2__SCAN_IN, P2_U5116);
  nand ginst16897 (P2_U7328, P2_INSTQUEUE_REG_8__2__SCAN_IN, P2_U5059);
  nand ginst16898 (P2_U7329, P2_INSTQUEUE_REG_9__2__SCAN_IN, P2_U5002);
  nand ginst16899 (P2_U7330, P2_INSTQUEUE_REG_10__2__SCAN_IN, P2_U4944);
  nand ginst16900 (P2_U7331, P2_INSTQUEUE_REG_11__2__SCAN_IN, P2_U4887);
  nand ginst16901 (P2_U7332, P2_INSTQUEUE_REG_12__2__SCAN_IN, P2_U4829);
  nand ginst16902 (P2_U7333, P2_INSTQUEUE_REG_13__2__SCAN_IN, P2_U4772);
  nand ginst16903 (P2_U7334, P2_INSTQUEUE_REG_14__2__SCAN_IN, P2_U4713);
  nand ginst16904 (P2_U7335, P2_INSTQUEUE_REG_15__2__SCAN_IN, P2_U4653);
  nand ginst16905 (P2_U7336, P2_U4313, P2_U4314, P2_U4315, P2_U4316);
  nand ginst16906 (P2_U7337, P2_INSTQUEUE_REG_8__2__SCAN_IN, P2_U2538);
  nand ginst16907 (P2_U7338, P2_INSTQUEUE_REG_9__2__SCAN_IN, P2_U2537);
  nand ginst16908 (P2_U7339, P2_INSTQUEUE_REG_10__2__SCAN_IN, P2_U2536);
  nand ginst16909 (P2_U7340, P2_INSTQUEUE_REG_11__2__SCAN_IN, P2_U2535);
  nand ginst16910 (P2_U7341, P2_INSTQUEUE_REG_12__2__SCAN_IN, P2_U2534);
  nand ginst16911 (P2_U7342, P2_INSTQUEUE_REG_13__2__SCAN_IN, P2_U2533);
  nand ginst16912 (P2_U7343, P2_INSTQUEUE_REG_14__2__SCAN_IN, P2_U2531);
  nand ginst16913 (P2_U7344, P2_INSTQUEUE_REG_15__2__SCAN_IN, P2_U2530);
  nand ginst16914 (P2_U7345, P2_INSTQUEUE_REG_7__2__SCAN_IN, P2_U2528);
  nand ginst16915 (P2_U7346, P2_INSTQUEUE_REG_6__2__SCAN_IN, P2_U2527);
  nand ginst16916 (P2_U7347, P2_INSTQUEUE_REG_5__2__SCAN_IN, P2_U2526);
  nand ginst16917 (P2_U7348, P2_INSTQUEUE_REG_4__2__SCAN_IN, P2_U2524);
  nand ginst16918 (P2_U7349, P2_INSTQUEUE_REG_3__2__SCAN_IN, P2_U2522);
  nand ginst16919 (P2_U7350, P2_INSTQUEUE_REG_2__2__SCAN_IN, P2_U2521);
  nand ginst16920 (P2_U7351, P2_INSTQUEUE_REG_1__2__SCAN_IN, P2_U2519);
  nand ginst16921 (P2_U7352, P2_INSTQUEUE_REG_0__2__SCAN_IN, P2_U2517);
  nand ginst16922 (P2_U7353, P2_U4317, P2_U4318, P2_U4319, P2_U4320);
  nand ginst16923 (P2_U7354, P2_INSTQUEUE_REG_0__1__SCAN_IN, P2_U5517);
  nand ginst16924 (P2_U7355, P2_INSTQUEUE_REG_1__1__SCAN_IN, P2_U5460);
  nand ginst16925 (P2_U7356, P2_INSTQUEUE_REG_2__1__SCAN_IN, P2_U5402);
  nand ginst16926 (P2_U7357, P2_INSTQUEUE_REG_3__1__SCAN_IN, P2_U5345);
  nand ginst16927 (P2_U7358, P2_INSTQUEUE_REG_4__1__SCAN_IN, P2_U5287);
  nand ginst16928 (P2_U7359, P2_INSTQUEUE_REG_5__1__SCAN_IN, P2_U5230);
  nand ginst16929 (P2_U7360, P2_INSTQUEUE_REG_6__1__SCAN_IN, P2_U5172);
  nand ginst16930 (P2_U7361, P2_INSTQUEUE_REG_7__1__SCAN_IN, P2_U5116);
  nand ginst16931 (P2_U7362, P2_INSTQUEUE_REG_8__1__SCAN_IN, P2_U5059);
  nand ginst16932 (P2_U7363, P2_INSTQUEUE_REG_9__1__SCAN_IN, P2_U5002);
  nand ginst16933 (P2_U7364, P2_INSTQUEUE_REG_10__1__SCAN_IN, P2_U4944);
  nand ginst16934 (P2_U7365, P2_INSTQUEUE_REG_11__1__SCAN_IN, P2_U4887);
  nand ginst16935 (P2_U7366, P2_INSTQUEUE_REG_12__1__SCAN_IN, P2_U4829);
  nand ginst16936 (P2_U7367, P2_INSTQUEUE_REG_13__1__SCAN_IN, P2_U4772);
  nand ginst16937 (P2_U7368, P2_INSTQUEUE_REG_14__1__SCAN_IN, P2_U4713);
  nand ginst16938 (P2_U7369, P2_INSTQUEUE_REG_15__1__SCAN_IN, P2_U4653);
  nand ginst16939 (P2_U7370, P2_U4321, P2_U4322, P2_U4323, P2_U4324);
  nand ginst16940 (P2_U7371, P2_INSTQUEUE_REG_8__1__SCAN_IN, P2_U2538);
  nand ginst16941 (P2_U7372, P2_INSTQUEUE_REG_9__1__SCAN_IN, P2_U2537);
  nand ginst16942 (P2_U7373, P2_INSTQUEUE_REG_10__1__SCAN_IN, P2_U2536);
  nand ginst16943 (P2_U7374, P2_INSTQUEUE_REG_11__1__SCAN_IN, P2_U2535);
  nand ginst16944 (P2_U7375, P2_INSTQUEUE_REG_12__1__SCAN_IN, P2_U2534);
  nand ginst16945 (P2_U7376, P2_INSTQUEUE_REG_13__1__SCAN_IN, P2_U2533);
  nand ginst16946 (P2_U7377, P2_INSTQUEUE_REG_14__1__SCAN_IN, P2_U2531);
  nand ginst16947 (P2_U7378, P2_INSTQUEUE_REG_15__1__SCAN_IN, P2_U2530);
  nand ginst16948 (P2_U7379, P2_INSTQUEUE_REG_7__1__SCAN_IN, P2_U2528);
  nand ginst16949 (P2_U7380, P2_INSTQUEUE_REG_6__1__SCAN_IN, P2_U2527);
  nand ginst16950 (P2_U7381, P2_INSTQUEUE_REG_5__1__SCAN_IN, P2_U2526);
  nand ginst16951 (P2_U7382, P2_INSTQUEUE_REG_4__1__SCAN_IN, P2_U2524);
  nand ginst16952 (P2_U7383, P2_INSTQUEUE_REG_3__1__SCAN_IN, P2_U2522);
  nand ginst16953 (P2_U7384, P2_INSTQUEUE_REG_2__1__SCAN_IN, P2_U2521);
  nand ginst16954 (P2_U7385, P2_INSTQUEUE_REG_1__1__SCAN_IN, P2_U2519);
  nand ginst16955 (P2_U7386, P2_INSTQUEUE_REG_0__1__SCAN_IN, P2_U2517);
  nand ginst16956 (P2_U7387, P2_U4325, P2_U4326, P2_U4327, P2_U4328);
  nand ginst16957 (P2_U7388, P2_INSTQUEUE_REG_0__0__SCAN_IN, P2_U5517);
  nand ginst16958 (P2_U7389, P2_INSTQUEUE_REG_1__0__SCAN_IN, P2_U5460);
  nand ginst16959 (P2_U7390, P2_INSTQUEUE_REG_2__0__SCAN_IN, P2_U5402);
  nand ginst16960 (P2_U7391, P2_INSTQUEUE_REG_3__0__SCAN_IN, P2_U5345);
  nand ginst16961 (P2_U7392, P2_INSTQUEUE_REG_4__0__SCAN_IN, P2_U5287);
  nand ginst16962 (P2_U7393, P2_INSTQUEUE_REG_5__0__SCAN_IN, P2_U5230);
  nand ginst16963 (P2_U7394, P2_INSTQUEUE_REG_6__0__SCAN_IN, P2_U5172);
  nand ginst16964 (P2_U7395, P2_INSTQUEUE_REG_7__0__SCAN_IN, P2_U5116);
  nand ginst16965 (P2_U7396, P2_INSTQUEUE_REG_8__0__SCAN_IN, P2_U5059);
  nand ginst16966 (P2_U7397, P2_INSTQUEUE_REG_9__0__SCAN_IN, P2_U5002);
  nand ginst16967 (P2_U7398, P2_INSTQUEUE_REG_10__0__SCAN_IN, P2_U4944);
  nand ginst16968 (P2_U7399, P2_INSTQUEUE_REG_11__0__SCAN_IN, P2_U4887);
  nand ginst16969 (P2_U7400, P2_INSTQUEUE_REG_12__0__SCAN_IN, P2_U4829);
  nand ginst16970 (P2_U7401, P2_INSTQUEUE_REG_13__0__SCAN_IN, P2_U4772);
  nand ginst16971 (P2_U7402, P2_INSTQUEUE_REG_14__0__SCAN_IN, P2_U4713);
  nand ginst16972 (P2_U7403, P2_INSTQUEUE_REG_15__0__SCAN_IN, P2_U4653);
  nand ginst16973 (P2_U7404, P2_U4329, P2_U4330, P2_U4331, P2_U4332);
  nand ginst16974 (P2_U7405, P2_INSTQUEUE_REG_8__0__SCAN_IN, P2_U2538);
  nand ginst16975 (P2_U7406, P2_INSTQUEUE_REG_9__0__SCAN_IN, P2_U2537);
  nand ginst16976 (P2_U7407, P2_INSTQUEUE_REG_10__0__SCAN_IN, P2_U2536);
  nand ginst16977 (P2_U7408, P2_INSTQUEUE_REG_11__0__SCAN_IN, P2_U2535);
  nand ginst16978 (P2_U7409, P2_INSTQUEUE_REG_12__0__SCAN_IN, P2_U2534);
  nand ginst16979 (P2_U7410, P2_INSTQUEUE_REG_13__0__SCAN_IN, P2_U2533);
  nand ginst16980 (P2_U7411, P2_INSTQUEUE_REG_14__0__SCAN_IN, P2_U2531);
  nand ginst16981 (P2_U7412, P2_INSTQUEUE_REG_15__0__SCAN_IN, P2_U2530);
  nand ginst16982 (P2_U7413, P2_INSTQUEUE_REG_7__0__SCAN_IN, P2_U2528);
  nand ginst16983 (P2_U7414, P2_INSTQUEUE_REG_6__0__SCAN_IN, P2_U2527);
  nand ginst16984 (P2_U7415, P2_INSTQUEUE_REG_5__0__SCAN_IN, P2_U2526);
  nand ginst16985 (P2_U7416, P2_INSTQUEUE_REG_4__0__SCAN_IN, P2_U2524);
  nand ginst16986 (P2_U7417, P2_INSTQUEUE_REG_3__0__SCAN_IN, P2_U2522);
  nand ginst16987 (P2_U7418, P2_INSTQUEUE_REG_2__0__SCAN_IN, P2_U2521);
  nand ginst16988 (P2_U7419, P2_INSTQUEUE_REG_1__0__SCAN_IN, P2_U2519);
  nand ginst16989 (P2_U7420, P2_INSTQUEUE_REG_0__0__SCAN_IN, P2_U2517);
  nand ginst16990 (P2_U7421, P2_U4333, P2_U4334, P2_U4335, P2_U4336);
  nand ginst16991 (P2_U7422, P2_U2352, P2_U7319);
  nand ginst16992 (P2_U7423, P2_STATE2_REG_3__SCAN_IN, P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN);
  nand ginst16993 (P2_U7424, P2_U2352, P2_U7353);
  nand ginst16994 (P2_U7425, P2_STATE2_REG_3__SCAN_IN, P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN);
  nand ginst16995 (P2_U7426, P2_U2439, P2_U3295);
  nand ginst16996 (P2_U7427, P2_U2352, P2_U7387);
  nand ginst16997 (P2_U7428, P2_STATE2_REG_3__SCAN_IN, P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN);
  nand ginst16998 (P2_U7429, P2_U2352, P2_U7421);
  nand ginst16999 (P2_U7430, P2_STATE2_REG_3__SCAN_IN, P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN);
  nand ginst17000 (P2_U7431, P2_U2439, P2_U3279);
  nand ginst17001 (P2_U7432, P2_U4413, P2_U4414, P2_U7431);
  nand ginst17002 (P2_U7433, P2_INSTADDRPOINTER_REG_9__SCAN_IN, P2_U7432);
  nand ginst17003 (P2_U7434, P2_REIP_REG_9__SCAN_IN, P2_U2353);
  nand ginst17004 (P2_U7435, P2_EAX_REG_9__SCAN_IN, P2_U4412);
  nand ginst17005 (P2_U7436, P2_U2352, P2_U2608);
  nand ginst17006 (P2_U7437, P2_INSTADDRPOINTER_REG_8__SCAN_IN, P2_U7432);
  nand ginst17007 (P2_U7438, P2_REIP_REG_8__SCAN_IN, P2_U2353);
  nand ginst17008 (P2_U7439, P2_EAX_REG_8__SCAN_IN, P2_U4412);
  nand ginst17009 (P2_U7440, P2_U2352, P2_U2607);
  nand ginst17010 (P2_U7441, P2_INSTADDRPOINTER_REG_7__SCAN_IN, P2_U7432);
  nand ginst17011 (P2_U7442, P2_REIP_REG_7__SCAN_IN, P2_U2353);
  nand ginst17012 (P2_U7443, P2_EAX_REG_7__SCAN_IN, P2_U4412);
  nand ginst17013 (P2_U7444, P2_INSTADDRPOINTER_REG_6__SCAN_IN, P2_U7432);
  nand ginst17014 (P2_U7445, P2_REIP_REG_6__SCAN_IN, P2_U2353);
  nand ginst17015 (P2_U7446, P2_EAX_REG_6__SCAN_IN, P2_U4412);
  nand ginst17016 (P2_U7447, P2_INSTADDRPOINTER_REG_5__SCAN_IN, P2_U7432);
  nand ginst17017 (P2_U7448, P2_REIP_REG_5__SCAN_IN, P2_U2353);
  nand ginst17018 (P2_U7449, P2_EAX_REG_5__SCAN_IN, P2_U4412);
  nand ginst17019 (P2_U7450, P2_INSTADDRPOINTER_REG_4__SCAN_IN, P2_U7432);
  nand ginst17020 (P2_U7451, P2_REIP_REG_4__SCAN_IN, P2_U2353);
  nand ginst17021 (P2_U7452, P2_EAX_REG_4__SCAN_IN, P2_U4412);
  nand ginst17022 (P2_U7453, P2_INSTADDRPOINTER_REG_31__SCAN_IN, P2_U7432);
  nand ginst17023 (P2_U7454, P2_REIP_REG_31__SCAN_IN, P2_U2353);
  nand ginst17024 (P2_U7455, P2_EAX_REG_31__SCAN_IN, P2_U4412);
  nand ginst17025 (P2_U7456, P2_INSTADDRPOINTER_REG_30__SCAN_IN, P2_U7432);
  nand ginst17026 (P2_U7457, P2_REIP_REG_30__SCAN_IN, P2_U2353);
  nand ginst17027 (P2_U7458, P2_EAX_REG_30__SCAN_IN, P2_U4412);
  nand ginst17028 (P2_U7459, P2_INSTADDRPOINTER_REG_3__SCAN_IN, P2_U7432);
  nand ginst17029 (P2_U7460, P2_REIP_REG_3__SCAN_IN, P2_U2353);
  nand ginst17030 (P2_U7461, P2_EAX_REG_3__SCAN_IN, P2_U4412);
  nand ginst17031 (P2_U7462, P2_INSTADDRPOINTER_REG_29__SCAN_IN, P2_U7432);
  nand ginst17032 (P2_U7463, P2_REIP_REG_29__SCAN_IN, P2_U2353);
  nand ginst17033 (P2_U7464, P2_EAX_REG_29__SCAN_IN, P2_U4412);
  nand ginst17034 (P2_U7465, P2_INSTADDRPOINTER_REG_28__SCAN_IN, P2_U7432);
  nand ginst17035 (P2_U7466, P2_REIP_REG_28__SCAN_IN, P2_U2353);
  nand ginst17036 (P2_U7467, P2_EAX_REG_28__SCAN_IN, P2_U4412);
  nand ginst17037 (P2_U7468, P2_INSTADDRPOINTER_REG_27__SCAN_IN, P2_U7432);
  nand ginst17038 (P2_U7469, P2_REIP_REG_27__SCAN_IN, P2_U2353);
  nand ginst17039 (P2_U7470, P2_EAX_REG_27__SCAN_IN, P2_U4412);
  nand ginst17040 (P2_U7471, P2_INSTADDRPOINTER_REG_26__SCAN_IN, P2_U7432);
  nand ginst17041 (P2_U7472, P2_REIP_REG_26__SCAN_IN, P2_U2353);
  nand ginst17042 (P2_U7473, P2_EAX_REG_26__SCAN_IN, P2_U4412);
  nand ginst17043 (P2_U7474, P2_INSTADDRPOINTER_REG_25__SCAN_IN, P2_U7432);
  nand ginst17044 (P2_U7475, P2_REIP_REG_25__SCAN_IN, P2_U2353);
  nand ginst17045 (P2_U7476, P2_EAX_REG_25__SCAN_IN, P2_U4412);
  nand ginst17046 (P2_U7477, P2_INSTADDRPOINTER_REG_24__SCAN_IN, P2_U7432);
  nand ginst17047 (P2_U7478, P2_REIP_REG_24__SCAN_IN, P2_U2353);
  nand ginst17048 (P2_U7479, P2_EAX_REG_24__SCAN_IN, P2_U4412);
  nand ginst17049 (P2_U7480, P2_INSTADDRPOINTER_REG_23__SCAN_IN, P2_U7432);
  nand ginst17050 (P2_U7481, P2_REIP_REG_23__SCAN_IN, P2_U2353);
  nand ginst17051 (P2_U7482, P2_EAX_REG_23__SCAN_IN, P2_U4412);
  nand ginst17052 (P2_U7483, P2_INSTADDRPOINTER_REG_22__SCAN_IN, P2_U7432);
  nand ginst17053 (P2_U7484, P2_REIP_REG_22__SCAN_IN, P2_U2353);
  nand ginst17054 (P2_U7485, P2_EAX_REG_22__SCAN_IN, P2_U4412);
  nand ginst17055 (P2_U7486, P2_INSTADDRPOINTER_REG_21__SCAN_IN, P2_U7432);
  nand ginst17056 (P2_U7487, P2_REIP_REG_21__SCAN_IN, P2_U2353);
  nand ginst17057 (P2_U7488, P2_EAX_REG_21__SCAN_IN, P2_U4412);
  nand ginst17058 (P2_U7489, P2_INSTADDRPOINTER_REG_20__SCAN_IN, P2_U7432);
  nand ginst17059 (P2_U7490, P2_REIP_REG_20__SCAN_IN, P2_U2353);
  nand ginst17060 (P2_U7491, P2_EAX_REG_20__SCAN_IN, P2_U4412);
  nand ginst17061 (P2_U7492, P2_INSTADDRPOINTER_REG_2__SCAN_IN, P2_U7432);
  nand ginst17062 (P2_U7493, P2_REIP_REG_2__SCAN_IN, P2_U2353);
  nand ginst17063 (P2_U7494, P2_EAX_REG_2__SCAN_IN, P2_U4412);
  nand ginst17064 (P2_U7495, P2_INSTADDRPOINTER_REG_19__SCAN_IN, P2_U7432);
  nand ginst17065 (P2_U7496, P2_REIP_REG_19__SCAN_IN, P2_U2353);
  nand ginst17066 (P2_U7497, P2_EAX_REG_19__SCAN_IN, P2_U4412);
  nand ginst17067 (P2_U7498, P2_INSTADDRPOINTER_REG_18__SCAN_IN, P2_U7432);
  nand ginst17068 (P2_U7499, P2_REIP_REG_18__SCAN_IN, P2_U2353);
  nand ginst17069 (P2_U7500, P2_EAX_REG_18__SCAN_IN, P2_U4412);
  nand ginst17070 (P2_U7501, P2_INSTADDRPOINTER_REG_17__SCAN_IN, P2_U7432);
  nand ginst17071 (P2_U7502, P2_REIP_REG_17__SCAN_IN, P2_U2353);
  nand ginst17072 (P2_U7503, P2_EAX_REG_17__SCAN_IN, P2_U4412);
  nand ginst17073 (P2_U7504, P2_INSTADDRPOINTER_REG_16__SCAN_IN, P2_U7432);
  nand ginst17074 (P2_U7505, P2_REIP_REG_16__SCAN_IN, P2_U2353);
  nand ginst17075 (P2_U7506, P2_EAX_REG_16__SCAN_IN, P2_U4412);
  nand ginst17076 (P2_U7507, P2_INSTADDRPOINTER_REG_15__SCAN_IN, P2_U7432);
  nand ginst17077 (P2_U7508, P2_REIP_REG_15__SCAN_IN, P2_U2353);
  nand ginst17078 (P2_U7509, P2_EAX_REG_15__SCAN_IN, P2_U4412);
  nand ginst17079 (P2_U7510, P2_U2352, P2_U2614);
  nand ginst17080 (P2_U7511, P2_INSTADDRPOINTER_REG_14__SCAN_IN, P2_U7432);
  nand ginst17081 (P2_U7512, P2_REIP_REG_14__SCAN_IN, P2_U2353);
  nand ginst17082 (P2_U7513, P2_EAX_REG_14__SCAN_IN, P2_U4412);
  nand ginst17083 (P2_U7514, P2_U2352, P2_U2613);
  nand ginst17084 (P2_U7515, P2_INSTADDRPOINTER_REG_13__SCAN_IN, P2_U7432);
  nand ginst17085 (P2_U7516, P2_REIP_REG_13__SCAN_IN, P2_U2353);
  nand ginst17086 (P2_U7517, P2_EAX_REG_13__SCAN_IN, P2_U4412);
  nand ginst17087 (P2_U7518, P2_U2352, P2_U2612);
  nand ginst17088 (P2_U7519, P2_INSTADDRPOINTER_REG_12__SCAN_IN, P2_U7432);
  nand ginst17089 (P2_U7520, P2_REIP_REG_12__SCAN_IN, P2_U2353);
  nand ginst17090 (P2_U7521, P2_EAX_REG_12__SCAN_IN, P2_U4412);
  nand ginst17091 (P2_U7522, P2_U2352, P2_U2611);
  nand ginst17092 (P2_U7523, P2_INSTADDRPOINTER_REG_11__SCAN_IN, P2_U7432);
  nand ginst17093 (P2_U7524, P2_REIP_REG_11__SCAN_IN, P2_U2353);
  nand ginst17094 (P2_U7525, P2_EAX_REG_11__SCAN_IN, P2_U4412);
  nand ginst17095 (P2_U7526, P2_U2352, P2_U2610);
  nand ginst17096 (P2_U7527, P2_INSTADDRPOINTER_REG_10__SCAN_IN, P2_U7432);
  nand ginst17097 (P2_U7528, P2_REIP_REG_10__SCAN_IN, P2_U2353);
  nand ginst17098 (P2_U7529, P2_EAX_REG_10__SCAN_IN, P2_U4412);
  nand ginst17099 (P2_U7530, P2_U2352, P2_U2609);
  nand ginst17100 (P2_U7531, P2_INSTADDRPOINTER_REG_1__SCAN_IN, P2_U7432);
  nand ginst17101 (P2_U7532, P2_REIP_REG_1__SCAN_IN, P2_U2353);
  nand ginst17102 (P2_U7533, P2_EAX_REG_1__SCAN_IN, P2_U4412);
  nand ginst17103 (P2_U7534, P2_INSTADDRPOINTER_REG_0__SCAN_IN, P2_U7432);
  nand ginst17104 (P2_U7535, P2_REIP_REG_0__SCAN_IN, P2_U2353);
  nand ginst17105 (P2_U7536, P2_EAX_REG_0__SCAN_IN, P2_U4412);
  nand ginst17106 (P2_U7537, P2_EBX_REG_9__SCAN_IN, P2_U7869);
  nand ginst17107 (P2_U7538, P2_EBX_REG_8__SCAN_IN, P2_U7869);
  nand ginst17108 (P2_U7539, P2_EBX_REG_31__SCAN_IN, P2_U7869);
  nand ginst17109 (P2_U7540, P2_EBX_REG_30__SCAN_IN, P2_U7869);
  nand ginst17110 (P2_U7541, P2_EBX_REG_29__SCAN_IN, P2_U7869);
  nand ginst17111 (P2_U7542, P2_EBX_REG_28__SCAN_IN, P2_U7869);
  nand ginst17112 (P2_U7543, P2_EBX_REG_27__SCAN_IN, P2_U7869);
  nand ginst17113 (P2_U7544, P2_EBX_REG_26__SCAN_IN, P2_U7869);
  nand ginst17114 (P2_U7545, P2_EBX_REG_25__SCAN_IN, P2_U7869);
  nand ginst17115 (P2_U7546, P2_EBX_REG_24__SCAN_IN, P2_U7869);
  nand ginst17116 (P2_U7547, P2_EBX_REG_23__SCAN_IN, P2_U7869);
  nand ginst17117 (P2_U7548, P2_EBX_REG_22__SCAN_IN, P2_U7869);
  nand ginst17118 (P2_U7549, P2_EBX_REG_21__SCAN_IN, P2_U7869);
  nand ginst17119 (P2_U7550, P2_EBX_REG_20__SCAN_IN, P2_U7869);
  nand ginst17120 (P2_U7551, P2_EBX_REG_19__SCAN_IN, P2_U7869);
  nand ginst17121 (P2_U7552, P2_EBX_REG_18__SCAN_IN, P2_U7869);
  nand ginst17122 (P2_U7553, P2_EBX_REG_17__SCAN_IN, P2_U7869);
  nand ginst17123 (P2_U7554, P2_EBX_REG_16__SCAN_IN, P2_U7869);
  nand ginst17124 (P2_U7555, P2_EBX_REG_15__SCAN_IN, P2_U7869);
  nand ginst17125 (P2_U7556, P2_EBX_REG_14__SCAN_IN, P2_U7869);
  nand ginst17126 (P2_U7557, P2_EBX_REG_13__SCAN_IN, P2_U7869);
  nand ginst17127 (P2_U7558, P2_EBX_REG_12__SCAN_IN, P2_U7869);
  nand ginst17128 (P2_U7559, P2_EBX_REG_11__SCAN_IN, P2_U7869);
  nand ginst17129 (P2_U7560, P2_EBX_REG_10__SCAN_IN, P2_U7869);
  nand ginst17130 (P2_U7561, P2_U3294, P2_U4596);
  nand ginst17131 (P2_U7562, P2_U4428, P2_U7285);
  nand ginst17132 (P2_U7563, P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN, P2_U7561);
  nand ginst17133 (P2_U7564, P2_U4428, P2_U7319);
  nand ginst17134 (P2_U7565, P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P2_U7561);
  nand ginst17135 (P2_U7566, P2_U4428, P2_U7353);
  nand ginst17136 (P2_U7567, P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN, P2_U7561);
  nand ginst17137 (P2_U7568, P2_U4428, P2_U7387);
  nand ginst17138 (P2_U7569, P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P2_U7561);
  nand ginst17139 (P2_U7570, P2_U4428, P2_U7421);
  nand ginst17140 (P2_U7571, P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN, P2_U7561);
  nand ginst17141 (P2_U7572, P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN, P2_U7561);
  nand ginst17142 (P2_U7573, P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN, P2_U7561);
  nand ginst17143 (P2_U7574, P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN, P2_U7561);
  nand ginst17144 (P2_U7575, P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN, P2_U7561);
  nand ginst17145 (P2_U7576, P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P2_U7561);
  nand ginst17146 (P2_U7577, P2_U4377, P2_U5572);
  nand ginst17147 (P2_U7578, P2_STATE2_REG_0__SCAN_IN, P2_U4432);
  nand ginst17148 (P2_U7579, P2_U2450, P2_U2617);
  nand ginst17149 (P2_U7580, P2_U4376, P2_U5592);
  nand ginst17150 (P2_U7581, P2_U3525, P2_U6845, P2_U7867);
  nand ginst17151 (P2_U7582, P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN, P2_U4471);
  nand ginst17152 (P2_U7583, P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P2_U7890);
  nand ginst17153 (P2_U7584, P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN, P2_U7890);
  nand ginst17154 (P2_U7585, P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN, P2_U3284);
  nand ginst17155 (P2_U7586, P2_U4381, P2_U4424);
  nand ginst17156 (P2_U7587, P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN, P2_U4471);
  nand ginst17157 (P2_U7588, P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P2_U7890);
  nand ginst17158 (P2_U7589, P2_U2590, P2_U6845);
  nand ginst17159 (P2_U7590, P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P2_U4471);
  nand ginst17160 (P2_U7591, P2_U2376, P2_U4416, P2_U7871);
  nand ginst17161 (P2_U7592, P2_U3285, P2_U3539, P2_U4422, P2_U7591);
  nand ginst17162 (P2_U7593, P2_INSTADDRPOINTER_REG_9__SCAN_IN, P2_U7592);
  nand ginst17163 (P2_U7594, P2_STATE2_REG_1__SCAN_IN, P2_PHYADDRPOINTER_REG_9__SCAN_IN);
  nand ginst17164 (P2_U7595, P2_REIP_REG_9__SCAN_IN, P2_U4423);
  nand ginst17165 (P2_U7596, P2_EBX_REG_9__SCAN_IN, P2_U2358);
  nand ginst17166 (P2_U7597, P2_INSTADDRPOINTER_REG_8__SCAN_IN, P2_U7592);
  nand ginst17167 (P2_U7598, P2_STATE2_REG_1__SCAN_IN, P2_PHYADDRPOINTER_REG_8__SCAN_IN);
  nand ginst17168 (P2_U7599, P2_REIP_REG_8__SCAN_IN, P2_U4423);
  nand ginst17169 (P2_U7600, P2_EBX_REG_8__SCAN_IN, P2_U2358);
  nand ginst17170 (P2_U7601, P2_INSTADDRPOINTER_REG_7__SCAN_IN, P2_U7592);
  nand ginst17171 (P2_U7602, P2_STATE2_REG_1__SCAN_IN, P2_PHYADDRPOINTER_REG_7__SCAN_IN);
  nand ginst17172 (P2_U7603, P2_REIP_REG_7__SCAN_IN, P2_U4423);
  nand ginst17173 (P2_U7604, P2_EBX_REG_7__SCAN_IN, P2_U2358);
  nand ginst17174 (P2_U7605, P2_INSTADDRPOINTER_REG_6__SCAN_IN, P2_U7592);
  nand ginst17175 (P2_U7606, P2_STATE2_REG_1__SCAN_IN, P2_PHYADDRPOINTER_REG_6__SCAN_IN);
  nand ginst17176 (P2_U7607, P2_REIP_REG_6__SCAN_IN, P2_U4423);
  nand ginst17177 (P2_U7608, P2_EBX_REG_6__SCAN_IN, P2_U2358);
  nand ginst17178 (P2_U7609, P2_INSTADDRPOINTER_REG_5__SCAN_IN, P2_U7592);
  nand ginst17179 (P2_U7610, P2_STATE2_REG_1__SCAN_IN, P2_PHYADDRPOINTER_REG_5__SCAN_IN);
  nand ginst17180 (P2_U7611, P2_REIP_REG_5__SCAN_IN, P2_U4423);
  nand ginst17181 (P2_U7612, P2_EBX_REG_5__SCAN_IN, P2_U2358);
  nand ginst17182 (P2_U7613, P2_INSTADDRPOINTER_REG_4__SCAN_IN, P2_U7592);
  nand ginst17183 (P2_U7614, P2_STATE2_REG_1__SCAN_IN, P2_PHYADDRPOINTER_REG_4__SCAN_IN);
  nand ginst17184 (P2_U7615, P2_REIP_REG_4__SCAN_IN, P2_U4423);
  nand ginst17185 (P2_U7616, P2_EBX_REG_4__SCAN_IN, P2_U2358);
  nand ginst17186 (P2_U7617, P2_INSTADDRPOINTER_REG_31__SCAN_IN, P2_U7592);
  nand ginst17187 (P2_U7618, P2_STATE2_REG_1__SCAN_IN, P2_PHYADDRPOINTER_REG_31__SCAN_IN);
  nand ginst17188 (P2_U7619, P2_REIP_REG_31__SCAN_IN, P2_U4423);
  nand ginst17189 (P2_U7620, P2_EBX_REG_31__SCAN_IN, P2_U2358);
  nand ginst17190 (P2_U7621, P2_INSTADDRPOINTER_REG_30__SCAN_IN, P2_U7592);
  nand ginst17191 (P2_U7622, P2_STATE2_REG_1__SCAN_IN, P2_PHYADDRPOINTER_REG_30__SCAN_IN);
  nand ginst17192 (P2_U7623, P2_REIP_REG_30__SCAN_IN, P2_U4423);
  nand ginst17193 (P2_U7624, P2_EBX_REG_30__SCAN_IN, P2_U2358);
  nand ginst17194 (P2_U7625, P2_INSTADDRPOINTER_REG_3__SCAN_IN, P2_U7592);
  nand ginst17195 (P2_U7626, P2_STATE2_REG_1__SCAN_IN, P2_PHYADDRPOINTER_REG_3__SCAN_IN);
  nand ginst17196 (P2_U7627, P2_REIP_REG_3__SCAN_IN, P2_U4423);
  nand ginst17197 (P2_U7628, P2_EBX_REG_3__SCAN_IN, P2_U2358);
  nand ginst17198 (P2_U7629, P2_INSTADDRPOINTER_REG_29__SCAN_IN, P2_U7592);
  nand ginst17199 (P2_U7630, P2_STATE2_REG_1__SCAN_IN, P2_PHYADDRPOINTER_REG_29__SCAN_IN);
  nand ginst17200 (P2_U7631, P2_REIP_REG_29__SCAN_IN, P2_U4423);
  nand ginst17201 (P2_U7632, P2_EBX_REG_29__SCAN_IN, P2_U2358);
  nand ginst17202 (P2_U7633, P2_INSTADDRPOINTER_REG_28__SCAN_IN, P2_U7592);
  nand ginst17203 (P2_U7634, P2_STATE2_REG_1__SCAN_IN, P2_PHYADDRPOINTER_REG_28__SCAN_IN);
  nand ginst17204 (P2_U7635, P2_REIP_REG_28__SCAN_IN, P2_U4423);
  nand ginst17205 (P2_U7636, P2_EBX_REG_28__SCAN_IN, P2_U2358);
  nand ginst17206 (P2_U7637, P2_INSTADDRPOINTER_REG_27__SCAN_IN, P2_U7592);
  nand ginst17207 (P2_U7638, P2_STATE2_REG_1__SCAN_IN, P2_PHYADDRPOINTER_REG_27__SCAN_IN);
  nand ginst17208 (P2_U7639, P2_REIP_REG_27__SCAN_IN, P2_U4423);
  nand ginst17209 (P2_U7640, P2_EBX_REG_27__SCAN_IN, P2_U2358);
  nand ginst17210 (P2_U7641, P2_INSTADDRPOINTER_REG_26__SCAN_IN, P2_U7592);
  nand ginst17211 (P2_U7642, P2_STATE2_REG_1__SCAN_IN, P2_PHYADDRPOINTER_REG_26__SCAN_IN);
  nand ginst17212 (P2_U7643, P2_REIP_REG_26__SCAN_IN, P2_U4423);
  nand ginst17213 (P2_U7644, P2_EBX_REG_26__SCAN_IN, P2_U2358);
  nand ginst17214 (P2_U7645, P2_INSTADDRPOINTER_REG_25__SCAN_IN, P2_U7592);
  nand ginst17215 (P2_U7646, P2_STATE2_REG_1__SCAN_IN, P2_PHYADDRPOINTER_REG_25__SCAN_IN);
  nand ginst17216 (P2_U7647, P2_REIP_REG_25__SCAN_IN, P2_U4423);
  nand ginst17217 (P2_U7648, P2_EBX_REG_25__SCAN_IN, P2_U2358);
  nand ginst17218 (P2_U7649, P2_INSTADDRPOINTER_REG_24__SCAN_IN, P2_U7592);
  nand ginst17219 (P2_U7650, P2_STATE2_REG_1__SCAN_IN, P2_PHYADDRPOINTER_REG_24__SCAN_IN);
  nand ginst17220 (P2_U7651, P2_REIP_REG_24__SCAN_IN, P2_U4423);
  nand ginst17221 (P2_U7652, P2_EBX_REG_24__SCAN_IN, P2_U2358);
  nand ginst17222 (P2_U7653, P2_INSTADDRPOINTER_REG_23__SCAN_IN, P2_U7592);
  nand ginst17223 (P2_U7654, P2_STATE2_REG_1__SCAN_IN, P2_PHYADDRPOINTER_REG_23__SCAN_IN);
  nand ginst17224 (P2_U7655, P2_REIP_REG_23__SCAN_IN, P2_U4423);
  nand ginst17225 (P2_U7656, P2_EBX_REG_23__SCAN_IN, P2_U2358);
  nand ginst17226 (P2_U7657, P2_INSTADDRPOINTER_REG_22__SCAN_IN, P2_U7592);
  nand ginst17227 (P2_U7658, P2_STATE2_REG_1__SCAN_IN, P2_PHYADDRPOINTER_REG_22__SCAN_IN);
  nand ginst17228 (P2_U7659, P2_REIP_REG_22__SCAN_IN, P2_U4423);
  nand ginst17229 (P2_U7660, P2_EBX_REG_22__SCAN_IN, P2_U2358);
  nand ginst17230 (P2_U7661, P2_INSTADDRPOINTER_REG_21__SCAN_IN, P2_U7592);
  nand ginst17231 (P2_U7662, P2_STATE2_REG_1__SCAN_IN, P2_PHYADDRPOINTER_REG_21__SCAN_IN);
  nand ginst17232 (P2_U7663, P2_REIP_REG_21__SCAN_IN, P2_U4423);
  nand ginst17233 (P2_U7664, P2_EBX_REG_21__SCAN_IN, P2_U2358);
  nand ginst17234 (P2_U7665, P2_INSTADDRPOINTER_REG_20__SCAN_IN, P2_U7592);
  nand ginst17235 (P2_U7666, P2_STATE2_REG_1__SCAN_IN, P2_PHYADDRPOINTER_REG_20__SCAN_IN);
  nand ginst17236 (P2_U7667, P2_REIP_REG_20__SCAN_IN, P2_U4423);
  nand ginst17237 (P2_U7668, P2_EBX_REG_20__SCAN_IN, P2_U2358);
  nand ginst17238 (P2_U7669, P2_INSTADDRPOINTER_REG_2__SCAN_IN, P2_U7592);
  nand ginst17239 (P2_U7670, P2_STATE2_REG_1__SCAN_IN, P2_PHYADDRPOINTER_REG_2__SCAN_IN);
  nand ginst17240 (P2_U7671, P2_REIP_REG_2__SCAN_IN, P2_U4423);
  nand ginst17241 (P2_U7672, P2_EBX_REG_2__SCAN_IN, P2_U2358);
  nand ginst17242 (P2_U7673, P2_INSTADDRPOINTER_REG_19__SCAN_IN, P2_U7592);
  nand ginst17243 (P2_U7674, P2_STATE2_REG_1__SCAN_IN, P2_PHYADDRPOINTER_REG_19__SCAN_IN);
  nand ginst17244 (P2_U7675, P2_REIP_REG_19__SCAN_IN, P2_U4423);
  nand ginst17245 (P2_U7676, P2_EBX_REG_19__SCAN_IN, P2_U2358);
  nand ginst17246 (P2_U7677, P2_INSTADDRPOINTER_REG_18__SCAN_IN, P2_U7592);
  nand ginst17247 (P2_U7678, P2_STATE2_REG_1__SCAN_IN, P2_PHYADDRPOINTER_REG_18__SCAN_IN);
  nand ginst17248 (P2_U7679, P2_REIP_REG_18__SCAN_IN, P2_U4423);
  nand ginst17249 (P2_U7680, P2_EBX_REG_18__SCAN_IN, P2_U2358);
  nand ginst17250 (P2_U7681, P2_INSTADDRPOINTER_REG_17__SCAN_IN, P2_U7592);
  nand ginst17251 (P2_U7682, P2_STATE2_REG_1__SCAN_IN, P2_PHYADDRPOINTER_REG_17__SCAN_IN);
  nand ginst17252 (P2_U7683, P2_REIP_REG_17__SCAN_IN, P2_U4423);
  nand ginst17253 (P2_U7684, P2_EBX_REG_17__SCAN_IN, P2_U2358);
  nand ginst17254 (P2_U7685, P2_INSTADDRPOINTER_REG_16__SCAN_IN, P2_U7592);
  nand ginst17255 (P2_U7686, P2_STATE2_REG_1__SCAN_IN, P2_PHYADDRPOINTER_REG_16__SCAN_IN);
  nand ginst17256 (P2_U7687, P2_REIP_REG_16__SCAN_IN, P2_U4423);
  nand ginst17257 (P2_U7688, P2_EBX_REG_16__SCAN_IN, P2_U2358);
  nand ginst17258 (P2_U7689, P2_INSTADDRPOINTER_REG_15__SCAN_IN, P2_U7592);
  nand ginst17259 (P2_U7690, P2_STATE2_REG_1__SCAN_IN, P2_PHYADDRPOINTER_REG_15__SCAN_IN);
  nand ginst17260 (P2_U7691, P2_REIP_REG_15__SCAN_IN, P2_U4423);
  nand ginst17261 (P2_U7692, P2_EBX_REG_15__SCAN_IN, P2_U2358);
  nand ginst17262 (P2_U7693, P2_INSTADDRPOINTER_REG_14__SCAN_IN, P2_U7592);
  nand ginst17263 (P2_U7694, P2_STATE2_REG_1__SCAN_IN, P2_PHYADDRPOINTER_REG_14__SCAN_IN);
  nand ginst17264 (P2_U7695, P2_REIP_REG_14__SCAN_IN, P2_U4423);
  nand ginst17265 (P2_U7696, P2_EBX_REG_14__SCAN_IN, P2_U2358);
  nand ginst17266 (P2_U7697, P2_INSTADDRPOINTER_REG_13__SCAN_IN, P2_U7592);
  nand ginst17267 (P2_U7698, P2_STATE2_REG_1__SCAN_IN, P2_PHYADDRPOINTER_REG_13__SCAN_IN);
  nand ginst17268 (P2_U7699, P2_REIP_REG_13__SCAN_IN, P2_U4423);
  nand ginst17269 (P2_U7700, P2_EBX_REG_13__SCAN_IN, P2_U2358);
  nand ginst17270 (P2_U7701, P2_INSTADDRPOINTER_REG_12__SCAN_IN, P2_U7592);
  nand ginst17271 (P2_U7702, P2_STATE2_REG_1__SCAN_IN, P2_PHYADDRPOINTER_REG_12__SCAN_IN);
  nand ginst17272 (P2_U7703, P2_REIP_REG_12__SCAN_IN, P2_U4423);
  nand ginst17273 (P2_U7704, P2_EBX_REG_12__SCAN_IN, P2_U2358);
  nand ginst17274 (P2_U7705, P2_INSTADDRPOINTER_REG_11__SCAN_IN, P2_U7592);
  nand ginst17275 (P2_U7706, P2_STATE2_REG_1__SCAN_IN, P2_PHYADDRPOINTER_REG_11__SCAN_IN);
  nand ginst17276 (P2_U7707, P2_REIP_REG_11__SCAN_IN, P2_U4423);
  nand ginst17277 (P2_U7708, P2_EBX_REG_11__SCAN_IN, P2_U2358);
  nand ginst17278 (P2_U7709, P2_INSTADDRPOINTER_REG_10__SCAN_IN, P2_U7592);
  nand ginst17279 (P2_U7710, P2_STATE2_REG_1__SCAN_IN, P2_PHYADDRPOINTER_REG_10__SCAN_IN);
  nand ginst17280 (P2_U7711, P2_REIP_REG_10__SCAN_IN, P2_U4423);
  nand ginst17281 (P2_U7712, P2_EBX_REG_10__SCAN_IN, P2_U2358);
  nand ginst17282 (P2_U7713, P2_INSTADDRPOINTER_REG_1__SCAN_IN, P2_U7592);
  nand ginst17283 (P2_U7714, P2_STATE2_REG_1__SCAN_IN, P2_PHYADDRPOINTER_REG_1__SCAN_IN);
  nand ginst17284 (P2_U7715, P2_REIP_REG_1__SCAN_IN, P2_U4423);
  nand ginst17285 (P2_U7716, P2_EBX_REG_1__SCAN_IN, P2_U2358);
  nand ginst17286 (P2_U7717, P2_U4387, P2_U7885);
  nand ginst17287 (P2_U7718, P2_INSTADDRPOINTER_REG_0__SCAN_IN, P2_U7739);
  nand ginst17288 (P2_U7719, P2_STATE2_REG_1__SCAN_IN, P2_PHYADDRPOINTER_REG_0__SCAN_IN);
  nand ginst17289 (P2_U7720, P2_REIP_REG_0__SCAN_IN, P2_U4423);
  nand ginst17290 (P2_U7721, P2_EBX_REG_0__SCAN_IN, P2_U2358);
  nand ginst17291 (P2_U7722, P2_U3575, P2_U7720);
  nand ginst17292 (P2_U7723, P2_U3536, P2_U3550);
  nand ginst17293 (P2_U7724, P2_R2219_U28, P2_U7723);
  nand ginst17294 (P2_U7725, P2_R2219_U30, P2_U7723);
  nand ginst17295 (P2_U7726, P2_R2238_U19, P2_U2356);
  nand ginst17296 (P2_U7727, P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN, P2_U3284);
  nand ginst17297 (P2_U7728, P2_R2238_U20, P2_U2356);
  nand ginst17298 (P2_U7729, P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P2_U3284);
  nand ginst17299 (P2_U7730, P2_R2238_U21, P2_U2356);
  nand ginst17300 (P2_U7731, P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN, P2_U3284);
  nand ginst17301 (P2_U7732, P2_R2238_U22, P2_U2356);
  nand ginst17302 (P2_U7733, P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P2_U3284);
  nand ginst17303 (P2_U7734, P2_R2238_U7, P2_U2356);
  nand ginst17304 (P2_U7735, P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN, P2_U3284);
  nand ginst17305 (P2_U7736, P2_U3295, P2_U3525, P2_U7873);
  nand ginst17306 (P2_U7737, P2_U3272, P2_U4422, P2_U7589, P2_U7590);
  nand ginst17307 (P2_U7738, P2_U2617, P2_U7861);
  nand ginst17308 (P2_U7739, P2_U3285, P2_U3539, P2_U4422, P2_U7591);
  nand ginst17309 (P2_U7740, P2_U3521, P2_U5571, P2_U5573, P2_U7744);
  nand ginst17310 (P2_U7741, P2_U2391, P2_U3544);
  nand ginst17311 (P2_U7742, P2_U2377, P2_U6572);
  nand ginst17312 (P2_U7743, P2_U4448, P2_U7741, P2_U7742);
  nand ginst17313 (P2_U7744, P2_U3278, P2_U7745);
  nand ginst17314 (P2_U7745, P2_U2617, P2_U7861);
  nand ginst17315 (P2_U7746, P2_U4592, P2_U8002, P2_U8003);
  nand ginst17316 (P2_U7747, P2_U4592, P2_U7970, P2_U7971);
  nand ginst17317 (P2_U7748, P2_U4592, P2_U7954, P2_U7955);
  nand ginst17318 (P2_U7749, P2_U4592, P2_U8034, P2_U8035);
  nand ginst17319 (P2_U7750, P2_U4592, P2_U8018, P2_U8019);
  nand ginst17320 (P2_U7751, P2_U4592, P2_U7986, P2_U7987);
  nand ginst17321 (P2_U7752, P2_U4592, P2_U7938, P2_U7939);
  nand ginst17322 (P2_U7753, P2_U4592, P2_U7922, P2_U7923);
  nand ginst17323 (P2_U7754, P2_U4592, P2_U8153, P2_U8154);
  nand ginst17324 (P2_U7755, P2_U4592, P2_U8169, P2_U8170);
  nand ginst17325 (P2_U7756, P2_U4592, P2_U8185, P2_U8186);
  nand ginst17326 (P2_U7757, P2_U4592, P2_U8201, P2_U8202);
  nand ginst17327 (P2_U7758, P2_U4592, P2_U8217, P2_U8218);
  nand ginst17328 (P2_U7759, P2_U4592, P2_U8233, P2_U8234);
  nand ginst17329 (P2_U7760, P2_U4592, P2_U8249, P2_U8250);
  nand ginst17330 (P2_U7761, P2_U4592, P2_U8265, P2_U8266);
  nand ginst17331 (P2_U7762, P2_U4593, P2_U8004, P2_U8005);
  nand ginst17332 (P2_U7763, P2_U4593, P2_U7972, P2_U7973);
  nand ginst17333 (P2_U7764, P2_U4593, P2_U7956, P2_U7957);
  nand ginst17334 (P2_U7765, P2_U4593, P2_U8036, P2_U8037);
  nand ginst17335 (P2_U7766, P2_U4593, P2_U8020, P2_U8021);
  nand ginst17336 (P2_U7767, P2_U4593, P2_U7988, P2_U7989);
  nand ginst17337 (P2_U7768, P2_U4593, P2_U7940, P2_U7941);
  nand ginst17338 (P2_U7769, P2_U4593, P2_U7924, P2_U7925);
  nand ginst17339 (P2_U7770, P2_U4593, P2_U8155, P2_U8156);
  nand ginst17340 (P2_U7771, P2_U4593, P2_U8171, P2_U8172);
  nand ginst17341 (P2_U7772, P2_U4593, P2_U8187, P2_U8188);
  nand ginst17342 (P2_U7773, P2_U4593, P2_U8203, P2_U8204);
  nand ginst17343 (P2_U7774, P2_U4593, P2_U8219, P2_U8220);
  nand ginst17344 (P2_U7775, P2_U4593, P2_U8235, P2_U8236);
  nand ginst17345 (P2_U7776, P2_U4593, P2_U8251, P2_U8252);
  nand ginst17346 (P2_U7777, P2_U4593, P2_U8267, P2_U8268);
  nand ginst17347 (P2_U7778, P2_U2456, P2_U8006, P2_U8007);
  nand ginst17348 (P2_U7779, P2_U2456, P2_U7974, P2_U7975);
  nand ginst17349 (P2_U7780, P2_U2456, P2_U7958, P2_U7959);
  nand ginst17350 (P2_U7781, P2_U2456, P2_U8038, P2_U8039);
  nand ginst17351 (P2_U7782, P2_U2456, P2_U8022, P2_U8023);
  nand ginst17352 (P2_U7783, P2_U2456, P2_U7990, P2_U7991);
  nand ginst17353 (P2_U7784, P2_U2456, P2_U7942, P2_U7943);
  nand ginst17354 (P2_U7785, P2_U2456, P2_U7926, P2_U7927);
  nand ginst17355 (P2_U7786, P2_U2456, P2_U8157, P2_U8158);
  nand ginst17356 (P2_U7787, P2_U2456, P2_U8173, P2_U8174);
  nand ginst17357 (P2_U7788, P2_U2456, P2_U8189, P2_U8190);
  nand ginst17358 (P2_U7789, P2_U2456, P2_U8205, P2_U8206);
  nand ginst17359 (P2_U7790, P2_U2456, P2_U8221, P2_U8222);
  nand ginst17360 (P2_U7791, P2_U2456, P2_U8237, P2_U8238);
  nand ginst17361 (P2_U7792, P2_U2456, P2_U8253, P2_U8254);
  nand ginst17362 (P2_U7793, P2_U2456, P2_U8269, P2_U8270);
  nand ginst17363 (P2_U7794, P2_U2454, P2_U8008, P2_U8009);
  nand ginst17364 (P2_U7795, P2_U2454, P2_U7976, P2_U7977);
  nand ginst17365 (P2_U7796, P2_U2454, P2_U7960, P2_U7961);
  nand ginst17366 (P2_U7797, P2_U2454, P2_U8040, P2_U8041);
  nand ginst17367 (P2_U7798, P2_U2454, P2_U8024, P2_U8025);
  nand ginst17368 (P2_U7799, P2_U2454, P2_U7992, P2_U7993);
  nand ginst17369 (P2_U7800, P2_U2454, P2_U7944, P2_U7945);
  nand ginst17370 (P2_U7801, P2_U2454, P2_U7928, P2_U7929);
  nand ginst17371 (P2_U7802, P2_U2454, P2_U8159, P2_U8160);
  nand ginst17372 (P2_U7803, P2_U2454, P2_U8175, P2_U8176);
  nand ginst17373 (P2_U7804, P2_U2454, P2_U8191, P2_U8192);
  nand ginst17374 (P2_U7805, P2_U2454, P2_U8207, P2_U8208);
  nand ginst17375 (P2_U7806, P2_U2454, P2_U8223, P2_U8224);
  nand ginst17376 (P2_U7807, P2_U2454, P2_U8239, P2_U8240);
  nand ginst17377 (P2_U7808, P2_U2454, P2_U8255, P2_U8256);
  nand ginst17378 (P2_U7809, P2_U2454, P2_U8271, P2_U8272);
  nand ginst17379 (P2_U7810, P2_U4590, P2_U8010, P2_U8011);
  nand ginst17380 (P2_U7811, P2_U4590, P2_U7978, P2_U7979);
  nand ginst17381 (P2_U7812, P2_U4590, P2_U7962, P2_U7963);
  nand ginst17382 (P2_U7813, P2_U4590, P2_U8042, P2_U8043);
  nand ginst17383 (P2_U7814, P2_U4590, P2_U8026, P2_U8027);
  nand ginst17384 (P2_U7815, P2_U4590, P2_U7994, P2_U7995);
  nand ginst17385 (P2_U7816, P2_U4590, P2_U7946, P2_U7947);
  nand ginst17386 (P2_U7817, P2_U4590, P2_U7930, P2_U7931);
  nand ginst17387 (P2_U7818, P2_U4590, P2_U8161, P2_U8162);
  nand ginst17388 (P2_U7819, P2_U4590, P2_U8177, P2_U8178);
  nand ginst17389 (P2_U7820, P2_U4590, P2_U8193, P2_U8194);
  nand ginst17390 (P2_U7821, P2_U4590, P2_U8209, P2_U8210);
  nand ginst17391 (P2_U7822, P2_U4590, P2_U8225, P2_U8226);
  nand ginst17392 (P2_U7823, P2_U4590, P2_U8241, P2_U8242);
  nand ginst17393 (P2_U7824, P2_U4590, P2_U8257, P2_U8258);
  nand ginst17394 (P2_U7825, P2_U4590, P2_U8273, P2_U8274);
  nand ginst17395 (P2_U7826, P2_U2453, P2_U8012, P2_U8013);
  nand ginst17396 (P2_U7827, P2_U2453, P2_U7980, P2_U7981);
  nand ginst17397 (P2_U7828, P2_U2453, P2_U7964, P2_U7965);
  nand ginst17398 (P2_U7829, P2_U2453, P2_U8044, P2_U8045);
  nand ginst17399 (P2_U7830, P2_U2453, P2_U8028, P2_U8029);
  nand ginst17400 (P2_U7831, P2_U2453, P2_U7996, P2_U7997);
  nand ginst17401 (P2_U7832, P2_U2453, P2_U7948, P2_U7949);
  nand ginst17402 (P2_U7833, P2_U2453, P2_U7932, P2_U7933);
  nand ginst17403 (P2_U7834, P2_U2453, P2_U8163, P2_U8164);
  nand ginst17404 (P2_U7835, P2_U2453, P2_U8179, P2_U8180);
  nand ginst17405 (P2_U7836, P2_U2453, P2_U8195, P2_U8196);
  nand ginst17406 (P2_U7837, P2_U2453, P2_U8211, P2_U8212);
  nand ginst17407 (P2_U7838, P2_U2453, P2_U8227, P2_U8228);
  nand ginst17408 (P2_U7839, P2_U2453, P2_U8243, P2_U8244);
  nand ginst17409 (P2_U7840, P2_U2453, P2_U8259, P2_U8260);
  nand ginst17410 (P2_U7841, P2_U2453, P2_U8275, P2_U8276);
  nand ginst17411 (P2_U7842, P2_U2452, P2_U8014, P2_U8015);
  nand ginst17412 (P2_U7843, P2_U2452, P2_U7982, P2_U7983);
  nand ginst17413 (P2_U7844, P2_U2452, P2_U7966, P2_U7967);
  nand ginst17414 (P2_U7845, P2_U2452, P2_U8046, P2_U8047);
  nand ginst17415 (P2_U7846, P2_U2452, P2_U8030, P2_U8031);
  nand ginst17416 (P2_U7847, P2_U2452, P2_U7998, P2_U7999);
  nand ginst17417 (P2_U7848, P2_U2452, P2_U7950, P2_U7951);
  nand ginst17418 (P2_U7849, P2_U2452, P2_U7934, P2_U7935);
  nand ginst17419 (P2_U7850, P2_U2452, P2_U8165, P2_U8166);
  nand ginst17420 (P2_U7851, P2_U2452, P2_U8181, P2_U8182);
  nand ginst17421 (P2_U7852, P2_U2452, P2_U8197, P2_U8198);
  nand ginst17422 (P2_U7853, P2_U2452, P2_U8213, P2_U8214);
  nand ginst17423 (P2_U7854, P2_U2452, P2_U8229, P2_U8230);
  nand ginst17424 (P2_U7855, P2_U2452, P2_U8245, P2_U8246);
  nand ginst17425 (P2_U7856, P2_U2452, P2_U8261, P2_U8262);
  nand ginst17426 (P2_U7857, P2_U2452, P2_U8277, P2_U8278);
  nand ginst17427 (P2_U7858, P2_U2455, P2_U8016, P2_U8017);
  not ginst17428 (P2_U7859, P2_U3280);
  nand ginst17429 (P2_U7860, P2_U2455, P2_U7984, P2_U7985);
  not ginst17430 (P2_U7861, P2_U3279);
  nand ginst17431 (P2_U7862, P2_U2455, P2_U7968, P2_U7969);
  not ginst17432 (P2_U7863, P2_U3278);
  nand ginst17433 (P2_U7864, P2_U2455, P2_U8048, P2_U8049);
  not ginst17434 (P2_U7865, P2_U3521);
  nand ginst17435 (P2_U7866, P2_U2455, P2_U8032, P2_U8033);
  not ginst17436 (P2_U7867, P2_U3255);
  nand ginst17437 (P2_U7868, P2_U2455, P2_U8000, P2_U8001);
  not ginst17438 (P2_U7869, P2_U2617);
  nand ginst17439 (P2_U7870, P2_U2455, P2_U7952, P2_U7953);
  not ginst17440 (P2_U7871, P2_U3253);
  nand ginst17441 (P2_U7872, P2_U2455, P2_U7936, P2_U7937);
  not ginst17442 (P2_U7873, P2_U2616);
  nand ginst17443 (P2_U7874, P2_U2455, P2_U8167, P2_U8168);
  nand ginst17444 (P2_U7875, P2_U2455, P2_U8183, P2_U8184);
  nand ginst17445 (P2_U7876, P2_U2455, P2_U8199, P2_U8200);
  nand ginst17446 (P2_U7877, P2_U2455, P2_U8215, P2_U8216);
  nand ginst17447 (P2_U7878, P2_U2455, P2_U8231, P2_U8232);
  nand ginst17448 (P2_U7879, P2_U2455, P2_U8247, P2_U8248);
  nand ginst17449 (P2_U7880, P2_U2455, P2_U8263, P2_U8264);
  nand ginst17450 (P2_U7881, P2_U2455, P2_U8279, P2_U8280);
  nand ginst17451 (P2_U7882, P2_U4428, P2_U5590);
  nand ginst17452 (P2_U7883, P2_U3525, P2_U5596);
  nand ginst17453 (P2_U7884, P2_U4596, P2_U7883);
  nand ginst17454 (P2_U7885, P2_U3253, P2_U8347, P2_U8348);
  nand ginst17455 (P2_U7886, P2_U5589, P2_U7722);
  nand ginst17456 (P2_U7887, P2_U4459, P2_U5589);
  nand ginst17457 (P2_U7888, P2_U2589, P2_U4384, P2_U4385, P2_U4386, P2_U7887);
  nand ginst17458 (P2_U7889, P2_U4459, P2_U5589);
  nand ginst17459 (P2_U7890, P2_U2589, P2_U4379, P2_U4458, P2_U7889);
  nand ginst17460 (P2_U7891, P2_STATE_REG_1__SCAN_IN, P2_U4569, P2_U4572);
  nand ginst17461 (P2_U7892, P2_STATE_REG_0__SCAN_IN, P2_REQUESTPENDING_REG_SCAN_IN, P2_U3244);
  nand ginst17462 (P2_U7893, P2_STATE_REG_1__SCAN_IN, P2_U4569);
  nand ginst17463 (P2_U7894, P2_U4600, P2_U4615);
  nand ginst17464 (P2_U7895, P2_U7863, P2_U7871);
  nand ginst17465 (P2_U7896, P2_U3255, P2_U5595);
  nand ginst17466 (P2_U7897, P2_U4429, P2_U5589);
  nand ginst17467 (P2_U7898, P2_DATAWIDTH_REG_0__SCAN_IN, P2_REIP_REG_0__SCAN_IN);
  nand ginst17468 (P2_U7899, P2_BE_N_REG_3__SCAN_IN, P2_U3259);
  nand ginst17469 (P2_U7900, P2_BYTEENABLE_REG_3__SCAN_IN, P2_U4439);
  nand ginst17470 (P2_U7901, P2_BE_N_REG_2__SCAN_IN, P2_U3259);
  nand ginst17471 (P2_U7902, P2_BYTEENABLE_REG_2__SCAN_IN, P2_U4439);
  nand ginst17472 (P2_U7903, P2_BE_N_REG_1__SCAN_IN, P2_U3259);
  nand ginst17473 (P2_U7904, P2_BYTEENABLE_REG_1__SCAN_IN, P2_U4439);
  nand ginst17474 (P2_U7905, P2_BE_N_REG_0__SCAN_IN, P2_U3259);
  nand ginst17475 (P2_U7906, P2_BYTEENABLE_REG_0__SCAN_IN, P2_U4439);
  nand ginst17476 (P2_U7907, P2_STATE_REG_0__SCAN_IN, P2_U3267, P2_U3268);
  or ginst17477 (P2_U7908, NA, P2_STATE_REG_0__SCAN_IN);
  nand ginst17478 (P2_U7909, P2_STATE_REG_2__SCAN_IN, P2_U3266);
  nand ginst17479 (P2_U7910, P2_STATE_REG_0__SCAN_IN, P2_U4568);
  nand ginst17480 (P2_U7911, P2_STATE_REG_1__SCAN_IN, P2_U4572, P2_U4581);
  nand ginst17481 (P2_U7912, P2_U3258, P2_U4582);
  nand ginst17482 (P2_U7913, P2_STATE_REG_2__SCAN_IN, P2_STATE_REG_0__SCAN_IN, P2_U3267);
  nand ginst17483 (P2_U7914, P2_U3244, P2_U4584);
  or ginst17484 (P2_U7915, P2_STATE_REG_1__SCAN_IN, P2_STATE_REG_0__SCAN_IN);
  nand ginst17485 (P2_U7916, P2_STATE_REG_0__SCAN_IN, P2_U4473);
  not ginst17486 (P2_U7917, P2_U3589);
  nand ginst17487 (P2_U7918, P2_DATAWIDTH_REG_0__SCAN_IN, P2_U7917);
  nand ginst17488 (P2_U7919, P2_U3589, P2_U3590);
  nand ginst17489 (P2_U7920, P2_U3589, P2_U4589);
  nand ginst17490 (P2_U7921, P2_DATAWIDTH_REG_1__SCAN_IN, P2_U7917);
  nand ginst17491 (P2_U7922, P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P2_U3388);
  or ginst17492 (P2_U7923, P2_INSTQUEUE_REG_3__1__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN);
  or ginst17493 (P2_U7924, P2_INSTQUEUE_REG_0__1__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN);
  nand ginst17494 (P2_U7925, P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P2_U3422);
  or ginst17495 (P2_U7926, P2_INSTQUEUE_REG_1__1__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN);
  nand ginst17496 (P2_U7927, P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P2_U3411);
  nand ginst17497 (P2_U7928, P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P2_U3374);
  or ginst17498 (P2_U7929, P2_INSTQUEUE_REG_4__1__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN);
  nand ginst17499 (P2_U7930, P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P2_U3333);
  or ginst17500 (P2_U7931, P2_INSTQUEUE_REG_7__1__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN);
  nand ginst17501 (P2_U7932, P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P2_U3363);
  or ginst17502 (P2_U7933, P2_INSTQUEUE_REG_5__1__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN);
  nand ginst17503 (P2_U7934, P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P2_U3347);
  or ginst17504 (P2_U7935, P2_INSTQUEUE_REG_6__1__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN);
  nand ginst17505 (P2_U7936, P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P2_U3399);
  or ginst17506 (P2_U7937, P2_INSTQUEUE_REG_2__1__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN);
  nand ginst17507 (P2_U7938, P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P2_U3389);
  or ginst17508 (P2_U7939, P2_INSTQUEUE_REG_3__0__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN);
  or ginst17509 (P2_U7940, P2_INSTQUEUE_REG_0__0__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN);
  nand ginst17510 (P2_U7941, P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P2_U3423);
  or ginst17511 (P2_U7942, P2_INSTQUEUE_REG_1__0__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN);
  nand ginst17512 (P2_U7943, P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P2_U3412);
  nand ginst17513 (P2_U7944, P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P2_U3375);
  or ginst17514 (P2_U7945, P2_INSTQUEUE_REG_4__0__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN);
  nand ginst17515 (P2_U7946, P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P2_U3334);
  or ginst17516 (P2_U7947, P2_INSTQUEUE_REG_7__0__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN);
  nand ginst17517 (P2_U7948, P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P2_U3364);
  or ginst17518 (P2_U7949, P2_INSTQUEUE_REG_5__0__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN);
  nand ginst17519 (P2_U7950, P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P2_U3348);
  or ginst17520 (P2_U7951, P2_INSTQUEUE_REG_6__0__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN);
  nand ginst17521 (P2_U7952, P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P2_U3400);
  or ginst17522 (P2_U7953, P2_INSTQUEUE_REG_2__0__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN);
  nand ginst17523 (P2_U7954, P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P2_U3385);
  or ginst17524 (P2_U7955, P2_INSTQUEUE_REG_3__4__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN);
  or ginst17525 (P2_U7956, P2_INSTQUEUE_REG_0__4__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN);
  nand ginst17526 (P2_U7957, P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P2_U3419);
  or ginst17527 (P2_U7958, P2_INSTQUEUE_REG_1__4__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN);
  nand ginst17528 (P2_U7959, P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P2_U3408);
  nand ginst17529 (P2_U7960, P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P2_U3371);
  or ginst17530 (P2_U7961, P2_INSTQUEUE_REG_4__4__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN);
  nand ginst17531 (P2_U7962, P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P2_U3330);
  or ginst17532 (P2_U7963, P2_INSTQUEUE_REG_7__4__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN);
  nand ginst17533 (P2_U7964, P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P2_U3360);
  or ginst17534 (P2_U7965, P2_INSTQUEUE_REG_5__4__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN);
  nand ginst17535 (P2_U7966, P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P2_U3344);
  or ginst17536 (P2_U7967, P2_INSTQUEUE_REG_6__4__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN);
  nand ginst17537 (P2_U7968, P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P2_U3396);
  or ginst17538 (P2_U7969, P2_INSTQUEUE_REG_2__4__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN);
  nand ginst17539 (P2_U7970, P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P2_U3383);
  or ginst17540 (P2_U7971, P2_INSTQUEUE_REG_3__6__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN);
  or ginst17541 (P2_U7972, P2_INSTQUEUE_REG_0__6__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN);
  nand ginst17542 (P2_U7973, P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P2_U3417);
  or ginst17543 (P2_U7974, P2_INSTQUEUE_REG_1__6__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN);
  nand ginst17544 (P2_U7975, P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P2_U3406);
  nand ginst17545 (P2_U7976, P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P2_U3369);
  or ginst17546 (P2_U7977, P2_INSTQUEUE_REG_4__6__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN);
  nand ginst17547 (P2_U7978, P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P2_U3328);
  or ginst17548 (P2_U7979, P2_INSTQUEUE_REG_7__6__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN);
  nand ginst17549 (P2_U7980, P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P2_U3358);
  or ginst17550 (P2_U7981, P2_INSTQUEUE_REG_5__6__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN);
  nand ginst17551 (P2_U7982, P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P2_U3342);
  or ginst17552 (P2_U7983, P2_INSTQUEUE_REG_6__6__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN);
  nand ginst17553 (P2_U7984, P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P2_U3394);
  or ginst17554 (P2_U7985, P2_INSTQUEUE_REG_2__6__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN);
  nand ginst17555 (P2_U7986, P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P2_U3384);
  or ginst17556 (P2_U7987, P2_INSTQUEUE_REG_3__5__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN);
  or ginst17557 (P2_U7988, P2_INSTQUEUE_REG_0__5__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN);
  nand ginst17558 (P2_U7989, P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P2_U3418);
  or ginst17559 (P2_U7990, P2_INSTQUEUE_REG_1__5__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN);
  nand ginst17560 (P2_U7991, P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P2_U3407);
  nand ginst17561 (P2_U7992, P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P2_U3370);
  or ginst17562 (P2_U7993, P2_INSTQUEUE_REG_4__5__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN);
  nand ginst17563 (P2_U7994, P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P2_U3329);
  or ginst17564 (P2_U7995, P2_INSTQUEUE_REG_7__5__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN);
  nand ginst17565 (P2_U7996, P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P2_U3359);
  or ginst17566 (P2_U7997, P2_INSTQUEUE_REG_5__5__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN);
  nand ginst17567 (P2_U7998, P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P2_U3343);
  or ginst17568 (P2_U7999, P2_INSTQUEUE_REG_6__5__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN);
  nand ginst17569 (P2_U8000, P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P2_U3395);
  or ginst17570 (P2_U8001, P2_INSTQUEUE_REG_2__5__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN);
  nand ginst17571 (P2_U8002, P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P2_U3387);
  or ginst17572 (P2_U8003, P2_INSTQUEUE_REG_3__2__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN);
  or ginst17573 (P2_U8004, P2_INSTQUEUE_REG_0__2__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN);
  nand ginst17574 (P2_U8005, P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P2_U3421);
  or ginst17575 (P2_U8006, P2_INSTQUEUE_REG_1__2__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN);
  nand ginst17576 (P2_U8007, P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P2_U3410);
  nand ginst17577 (P2_U8008, P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P2_U3373);
  or ginst17578 (P2_U8009, P2_INSTQUEUE_REG_4__2__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN);
  nand ginst17579 (P2_U8010, P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P2_U3332);
  or ginst17580 (P2_U8011, P2_INSTQUEUE_REG_7__2__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN);
  nand ginst17581 (P2_U8012, P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P2_U3362);
  or ginst17582 (P2_U8013, P2_INSTQUEUE_REG_5__2__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN);
  nand ginst17583 (P2_U8014, P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P2_U3346);
  or ginst17584 (P2_U8015, P2_INSTQUEUE_REG_6__2__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN);
  nand ginst17585 (P2_U8016, P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P2_U3398);
  or ginst17586 (P2_U8017, P2_INSTQUEUE_REG_2__2__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN);
  nand ginst17587 (P2_U8018, P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P2_U3386);
  or ginst17588 (P2_U8019, P2_INSTQUEUE_REG_3__3__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN);
  or ginst17589 (P2_U8020, P2_INSTQUEUE_REG_0__3__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN);
  nand ginst17590 (P2_U8021, P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P2_U3420);
  or ginst17591 (P2_U8022, P2_INSTQUEUE_REG_1__3__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN);
  nand ginst17592 (P2_U8023, P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P2_U3409);
  nand ginst17593 (P2_U8024, P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P2_U3372);
  or ginst17594 (P2_U8025, P2_INSTQUEUE_REG_4__3__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN);
  nand ginst17595 (P2_U8026, P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P2_U3331);
  or ginst17596 (P2_U8027, P2_INSTQUEUE_REG_7__3__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN);
  nand ginst17597 (P2_U8028, P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P2_U3361);
  or ginst17598 (P2_U8029, P2_INSTQUEUE_REG_5__3__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN);
  nand ginst17599 (P2_U8030, P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P2_U3345);
  or ginst17600 (P2_U8031, P2_INSTQUEUE_REG_6__3__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN);
  nand ginst17601 (P2_U8032, P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P2_U3397);
  or ginst17602 (P2_U8033, P2_INSTQUEUE_REG_2__3__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN);
  nand ginst17603 (P2_U8034, P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P2_U3382);
  or ginst17604 (P2_U8035, P2_INSTQUEUE_REG_3__7__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN);
  or ginst17605 (P2_U8036, P2_INSTQUEUE_REG_0__7__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN);
  nand ginst17606 (P2_U8037, P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P2_U3416);
  or ginst17607 (P2_U8038, P2_INSTQUEUE_REG_1__7__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN);
  nand ginst17608 (P2_U8039, P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P2_U3405);
  nand ginst17609 (P2_U8040, P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P2_U3368);
  or ginst17610 (P2_U8041, P2_INSTQUEUE_REG_4__7__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN);
  nand ginst17611 (P2_U8042, P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P2_U3327);
  or ginst17612 (P2_U8043, P2_INSTQUEUE_REG_7__7__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN);
  nand ginst17613 (P2_U8044, P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P2_U3357);
  or ginst17614 (P2_U8045, P2_INSTQUEUE_REG_5__7__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN);
  nand ginst17615 (P2_U8046, P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P2_U3341);
  or ginst17616 (P2_U8047, P2_INSTQUEUE_REG_6__7__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN);
  nand ginst17617 (P2_U8048, P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P2_U3393);
  or ginst17618 (P2_U8049, P2_INSTQUEUE_REG_2__7__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN);
  nand ginst17619 (P2_U8050, P2_R2167_U6, P2_U4435);
  nand ginst17620 (P2_U8051, P2_U3297, P2_U4604);
  nand ginst17621 (P2_U8052, P2_U3293, P2_U7871);
  nand ginst17622 (P2_U8053, P2_U3253, P2_U3282);
  nand ginst17623 (P2_U8054, P2_U3297, P2_U4427);
  nand ginst17624 (P2_U8055, P2_U3289, P2_U3520);
  or ginst17625 (P2_U8056, P2_STATE2_REG_0__SCAN_IN, U211);
  nand ginst17626 (P2_U8057, P2_STATE2_REG_0__SCAN_IN, P2_U4617);
  nand ginst17627 (P2_U8058, P2_STATE2_REG_3__SCAN_IN, P2_U3299);
  nand ginst17628 (P2_U8059, P2_U2448, P2_U4620);
  nand ginst17629 (P2_U8060, P2_STATE2_REG_0__SCAN_IN, P2_U4631);
  nand ginst17630 (P2_U8061, P2_U3284, P2_U4619, P2_U4630);
  nand ginst17631 (P2_U8062, P2_R2182_U40, P2_U3318);
  nand ginst17632 (P2_U8063, P2_U3316, P2_U4637);
  not ginst17633 (P2_U8064, P2_U3579);
  nand ginst17634 (P2_U8065, P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN, P2_U3311);
  nand ginst17635 (P2_U8066, P2_U3310, P2_U4642);
  not ginst17636 (P2_U8067, P2_U3580);
  nand ginst17637 (P2_U8068, P2_U5574, P2_U7859);
  nand ginst17638 (P2_U8069, P2_U3280, P2_U5575);
  nand ginst17639 (P2_U8070, P2_U3297, P2_U4435);
  nand ginst17640 (P2_U8071, P2_R2167_U6, P2_U2359, P2_U4433);
  nand ginst17641 (P2_U8072, P2_U3594, P2_U4394);
  nand ginst17642 (P2_U8073, P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN, P2_U5584);
  nand ginst17643 (P2_U8074, P2_U3280, P2_U5586);
  nand ginst17644 (P2_U8075, P2_U2617, P2_U3279, P2_U7859);
  nand ginst17645 (P2_U8076, P2_U3253, P2_U4424);
  nand ginst17646 (P2_U8077, P2_U4475, P2_U7871);
  nand ginst17647 (P2_U8078, P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P2_U5585);
  nand ginst17648 (P2_U8079, P2_U3273, P2_U3276, P2_U4591);
  nand ginst17649 (P2_U8080, P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P2_U3277);
  nand ginst17650 (P2_U8081, P2_U3273, P2_U4590);
  not ginst17651 (P2_U8082, P2_U3581);
  nand ginst17652 (P2_U8083, P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P2_U5584);
  nand ginst17653 (P2_U8084, P2_U4394, P2_U5614);
  nand ginst17654 (P2_U8085, P2_INSTADDRPOINTER_REG_0__SCAN_IN, P2_U3528);
  nand ginst17655 (P2_U8086, P2_U3647, P2_U3683);
  not ginst17656 (P2_U8087, P2_U3597);
  nand ginst17657 (P2_U8088, P2_INSTADDRPOINTER_REG_1__SCAN_IN, P2_U3528);
  nand ginst17658 (P2_U8089, P2_R1957_U49, P2_U3647);
  not ginst17659 (P2_U8090, P2_U3598);
  nand ginst17660 (P2_U8091, P2_U5605, P2_U5616);
  nand ginst17661 (P2_U8092, P2_U3530, P2_U5606);
  nand ginst17662 (P2_U8093, P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN, P2_U5584);
  nand ginst17663 (P2_U8094, P2_U4394, P2_U5623);
  nand ginst17664 (P2_U8095, P2_U3255, P2_U3886, P2_U4597);
  nand ginst17665 (P2_U8096, P2_U5625, P2_U7867, P2_U7869);
  nand ginst17666 (P2_U8097, P2_U8095, P2_U8096);
  nand ginst17667 (P2_U8098, P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN, P2_U3271);
  nand ginst17668 (P2_U8099, P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P2_U3272);
  not ginst17669 (P2_U8100, P2_U3582);
  nand ginst17670 (P2_U8101, P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P2_U5584);
  nand ginst17671 (P2_U8102, P2_U4394, P2_U5633);
  nand ginst17672 (P2_U8103, P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN, P2_U5584);
  nand ginst17673 (P2_U8104, P2_U4394, P2_U5641);
  nand ginst17674 (P2_U8105, P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN, P2_U5643);
  nand ginst17675 (P2_U8106, P2_U3533, P2_U5651);
  nand ginst17676 (P2_U8107, P2_U4636, P2_U8064);
  nand ginst17677 (P2_U8108, P2_U3319, P2_U3579);
  nand ginst17678 (P2_U8109, P2_U8107, P2_U8108);
  nand ginst17679 (P2_U8110, P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN, P2_U5643);
  nand ginst17680 (P2_U8111, P2_U3533, P2_U5655);
  nand ginst17681 (P2_U8112, P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN, P2_U5643);
  nand ginst17682 (P2_U8113, P2_U3533, P2_U5660);
  nand ginst17683 (P2_U8114, P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P2_U5643);
  nand ginst17684 (P2_U8115, P2_U3533, P2_U5664);
  nand ginst17685 (P2_U8116, P2_U2359, P2_U2616, P2_U3280);
  nand ginst17686 (P2_U8117, P2_U2438, P2_U7873);
  nand ginst17687 (P2_U8118, P2_U8116, P2_U8117);
  nand ginst17688 (P2_U8119, P2_U3253, P2_U3278, P2_U3297);
  nand ginst17689 (P2_U8120, P2_R2167_U6, P2_U8118);
  nand ginst17690 (P2_U8121, P2_U7859, P2_U7873);
  nand ginst17691 (P2_U8122, P2_U2616, P2_U3282);
  nand ginst17692 (P2_U8123, P2_BYTEENABLE_REG_3__SCAN_IN, P2_U3547);
  nand ginst17693 (P2_U8124, P2_U3606, P2_U4438);
  nand ginst17694 (P2_U8125, P2_BYTEENABLE_REG_2__SCAN_IN, P2_U3547);
  nand ginst17695 (P2_U8126, P2_U3607, P2_U4438);
  nand ginst17696 (P2_U8127, P2_BYTEENABLE_REG_0__SCAN_IN, P2_U3547);
  nand ginst17697 (P2_U8128, P2_REIP_REG_0__SCAN_IN, P2_U4438);
  nand ginst17698 (P2_U8129, P2_U3552, P2_U4439);
  nand ginst17699 (P2_U8130, P2_W_R_N_REG_SCAN_IN, P2_U3259);
  nand ginst17700 (P2_U8131, P2_U3287, P2_U7873);
  nand ginst17701 (P2_U8132, P2_R2243_U8, P2_U2616);
  nand ginst17702 (P2_U8133, P2_U3257, P2_U6838);
  nand ginst17703 (P2_U8134, P2_MORE_REG_SCAN_IN, P2_U4400);
  nand ginst17704 (P2_U8135, P2_STATEBS16_REG_SCAN_IN, P2_U7917);
  nand ginst17705 (P2_U8136, BS16, P2_U3589);
  nand ginst17706 (P2_U8137, P2_REQUESTPENDING_REG_SCAN_IN, P2_U6843);
  nand ginst17707 (P2_U8138, P2_U4402, P2_U6852);
  nand ginst17708 (P2_U8139, P2_U3551, P2_U4439);
  nand ginst17709 (P2_U8140, P2_D_C_N_REG_SCAN_IN, P2_U3259);
  nand ginst17710 (P2_U8141, P2_M_IO_N_REG_SCAN_IN, P2_U3259);
  nand ginst17711 (P2_U8142, P2_MEMORYFETCH_REG_SCAN_IN, P2_U4439);
  nand ginst17712 (P2_U8143, P2_READREQUEST_REG_SCAN_IN, P2_U6857);
  nand ginst17713 (P2_U8144, P2_U4403, P2_U6858);
  nand ginst17714 (P2_U8145, P2_U3520, P2_U7873);
  nand ginst17715 (P2_U8146, P2_U2616, P2_U3297);
  nand ginst17716 (P2_U8147, P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P2_U4405);
  nand ginst17717 (P2_U8148, P2_U3273, P2_U7007);
  not ginst17718 (P2_U8149, P2_U3583);
  nand ginst17719 (P2_U8150, P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN, P2_U3273);
  nand ginst17720 (P2_U8151, P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P2_U3276);
  not ginst17721 (P2_U8152, P2_U3584);
  nand ginst17722 (P2_U8153, P2_U3327, P2_U3584);
  nand ginst17723 (P2_U8154, P2_U3431, P2_U8152);
  nand ginst17724 (P2_U8155, P2_U3368, P2_U3584);
  nand ginst17725 (P2_U8156, P2_U3465, P2_U8152);
  nand ginst17726 (P2_U8157, P2_U3357, P2_U3584);
  nand ginst17727 (P2_U8158, P2_U3454, P2_U8152);
  nand ginst17728 (P2_U8159, P2_U3416, P2_U3584);
  nand ginst17729 (P2_U8160, P2_U3511, P2_U8152);
  nand ginst17730 (P2_U8161, P2_U3382, P2_U3584);
  nand ginst17731 (P2_U8162, P2_U3477, P2_U8152);
  nand ginst17732 (P2_U8163, P2_U3405, P2_U3584);
  nand ginst17733 (P2_U8164, P2_U3500, P2_U8152);
  nand ginst17734 (P2_U8165, P2_U3393, P2_U3584);
  nand ginst17735 (P2_U8166, P2_U3488, P2_U8152);
  nand ginst17736 (P2_U8167, P2_U3341, P2_U3584);
  nand ginst17737 (P2_U8168, P2_U3442, P2_U8152);
  nand ginst17738 (P2_U8169, P2_U3328, P2_U3584);
  nand ginst17739 (P2_U8170, P2_U3432, P2_U8152);
  nand ginst17740 (P2_U8171, P2_U3369, P2_U3584);
  nand ginst17741 (P2_U8172, P2_U3466, P2_U8152);
  nand ginst17742 (P2_U8173, P2_U3358, P2_U3584);
  nand ginst17743 (P2_U8174, P2_U3455, P2_U8152);
  nand ginst17744 (P2_U8175, P2_U3417, P2_U3584);
  nand ginst17745 (P2_U8176, P2_U3512, P2_U8152);
  nand ginst17746 (P2_U8177, P2_U3383, P2_U3584);
  nand ginst17747 (P2_U8178, P2_U3478, P2_U8152);
  nand ginst17748 (P2_U8179, P2_U3406, P2_U3584);
  nand ginst17749 (P2_U8180, P2_U3501, P2_U8152);
  nand ginst17750 (P2_U8181, P2_U3394, P2_U3584);
  nand ginst17751 (P2_U8182, P2_U3489, P2_U8152);
  nand ginst17752 (P2_U8183, P2_U3342, P2_U3584);
  nand ginst17753 (P2_U8184, P2_U3443, P2_U8152);
  nand ginst17754 (P2_U8185, P2_U3329, P2_U3584);
  nand ginst17755 (P2_U8186, P2_U3433, P2_U8152);
  nand ginst17756 (P2_U8187, P2_U3370, P2_U3584);
  nand ginst17757 (P2_U8188, P2_U3467, P2_U8152);
  nand ginst17758 (P2_U8189, P2_U3359, P2_U3584);
  nand ginst17759 (P2_U8190, P2_U3456, P2_U8152);
  nand ginst17760 (P2_U8191, P2_U3418, P2_U3584);
  nand ginst17761 (P2_U8192, P2_U3513, P2_U8152);
  nand ginst17762 (P2_U8193, P2_U3384, P2_U3584);
  nand ginst17763 (P2_U8194, P2_U3479, P2_U8152);
  nand ginst17764 (P2_U8195, P2_U3407, P2_U3584);
  nand ginst17765 (P2_U8196, P2_U3502, P2_U8152);
  nand ginst17766 (P2_U8197, P2_U3395, P2_U3584);
  nand ginst17767 (P2_U8198, P2_U3490, P2_U8152);
  nand ginst17768 (P2_U8199, P2_U3343, P2_U3584);
  nand ginst17769 (P2_U8200, P2_U3444, P2_U8152);
  nand ginst17770 (P2_U8201, P2_U3330, P2_U3584);
  nand ginst17771 (P2_U8202, P2_U3434, P2_U8152);
  nand ginst17772 (P2_U8203, P2_U3371, P2_U3584);
  nand ginst17773 (P2_U8204, P2_U3468, P2_U8152);
  nand ginst17774 (P2_U8205, P2_U3360, P2_U3584);
  nand ginst17775 (P2_U8206, P2_U3457, P2_U8152);
  nand ginst17776 (P2_U8207, P2_U3419, P2_U3584);
  nand ginst17777 (P2_U8208, P2_U3514, P2_U8152);
  nand ginst17778 (P2_U8209, P2_U3385, P2_U3584);
  nand ginst17779 (P2_U8210, P2_U3480, P2_U8152);
  nand ginst17780 (P2_U8211, P2_U3408, P2_U3584);
  nand ginst17781 (P2_U8212, P2_U3503, P2_U8152);
  nand ginst17782 (P2_U8213, P2_U3396, P2_U3584);
  nand ginst17783 (P2_U8214, P2_U3491, P2_U8152);
  nand ginst17784 (P2_U8215, P2_U3344, P2_U3584);
  nand ginst17785 (P2_U8216, P2_U3445, P2_U8152);
  nand ginst17786 (P2_U8217, P2_U3331, P2_U3584);
  nand ginst17787 (P2_U8218, P2_U3435, P2_U8152);
  nand ginst17788 (P2_U8219, P2_U3372, P2_U3584);
  nand ginst17789 (P2_U8220, P2_U3469, P2_U8152);
  nand ginst17790 (P2_U8221, P2_U3361, P2_U3584);
  nand ginst17791 (P2_U8222, P2_U3458, P2_U8152);
  nand ginst17792 (P2_U8223, P2_U3420, P2_U3584);
  nand ginst17793 (P2_U8224, P2_U3515, P2_U8152);
  nand ginst17794 (P2_U8225, P2_U3386, P2_U3584);
  nand ginst17795 (P2_U8226, P2_U3481, P2_U8152);
  nand ginst17796 (P2_U8227, P2_U3409, P2_U3584);
  nand ginst17797 (P2_U8228, P2_U3504, P2_U8152);
  nand ginst17798 (P2_U8229, P2_U3397, P2_U3584);
  nand ginst17799 (P2_U8230, P2_U3492, P2_U8152);
  nand ginst17800 (P2_U8231, P2_U3345, P2_U3584);
  nand ginst17801 (P2_U8232, P2_U3446, P2_U8152);
  nand ginst17802 (P2_U8233, P2_U3332, P2_U3584);
  nand ginst17803 (P2_U8234, P2_U3436, P2_U8152);
  nand ginst17804 (P2_U8235, P2_U3373, P2_U3584);
  nand ginst17805 (P2_U8236, P2_U3470, P2_U8152);
  nand ginst17806 (P2_U8237, P2_U3362, P2_U3584);
  nand ginst17807 (P2_U8238, P2_U3459, P2_U8152);
  nand ginst17808 (P2_U8239, P2_U3421, P2_U3584);
  nand ginst17809 (P2_U8240, P2_U3516, P2_U8152);
  nand ginst17810 (P2_U8241, P2_U3387, P2_U3584);
  nand ginst17811 (P2_U8242, P2_U3482, P2_U8152);
  nand ginst17812 (P2_U8243, P2_U3410, P2_U3584);
  nand ginst17813 (P2_U8244, P2_U3505, P2_U8152);
  nand ginst17814 (P2_U8245, P2_U3398, P2_U3584);
  nand ginst17815 (P2_U8246, P2_U3493, P2_U8152);
  nand ginst17816 (P2_U8247, P2_U3346, P2_U3584);
  nand ginst17817 (P2_U8248, P2_U3447, P2_U8152);
  nand ginst17818 (P2_U8249, P2_U3333, P2_U3584);
  nand ginst17819 (P2_U8250, P2_U3437, P2_U8152);
  nand ginst17820 (P2_U8251, P2_U3374, P2_U3584);
  nand ginst17821 (P2_U8252, P2_U3471, P2_U8152);
  nand ginst17822 (P2_U8253, P2_U3363, P2_U3584);
  nand ginst17823 (P2_U8254, P2_U3460, P2_U8152);
  nand ginst17824 (P2_U8255, P2_U3422, P2_U3584);
  nand ginst17825 (P2_U8256, P2_U3517, P2_U8152);
  nand ginst17826 (P2_U8257, P2_U3388, P2_U3584);
  nand ginst17827 (P2_U8258, P2_U3483, P2_U8152);
  nand ginst17828 (P2_U8259, P2_U3411, P2_U3584);
  nand ginst17829 (P2_U8260, P2_U3506, P2_U8152);
  nand ginst17830 (P2_U8261, P2_U3399, P2_U3584);
  nand ginst17831 (P2_U8262, P2_U3494, P2_U8152);
  nand ginst17832 (P2_U8263, P2_U3347, P2_U3584);
  nand ginst17833 (P2_U8264, P2_U3448, P2_U8152);
  nand ginst17834 (P2_U8265, P2_U3334, P2_U3584);
  nand ginst17835 (P2_U8266, P2_U3438, P2_U8152);
  nand ginst17836 (P2_U8267, P2_U3375, P2_U3584);
  nand ginst17837 (P2_U8268, P2_U3472, P2_U8152);
  nand ginst17838 (P2_U8269, P2_U3364, P2_U3584);
  nand ginst17839 (P2_U8270, P2_U3461, P2_U8152);
  nand ginst17840 (P2_U8271, P2_U3423, P2_U3584);
  nand ginst17841 (P2_U8272, P2_U3518, P2_U8152);
  nand ginst17842 (P2_U8273, P2_U3389, P2_U3584);
  nand ginst17843 (P2_U8274, P2_U3484, P2_U8152);
  nand ginst17844 (P2_U8275, P2_U3412, P2_U3584);
  nand ginst17845 (P2_U8276, P2_U3507, P2_U8152);
  nand ginst17846 (P2_U8277, P2_U3400, P2_U3584);
  nand ginst17847 (P2_U8278, P2_U3495, P2_U8152);
  nand ginst17848 (P2_U8279, P2_U3348, P2_U3584);
  nand ginst17849 (P2_U8280, P2_U3449, P2_U8152);
  nand ginst17850 (P2_U8281, P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN, P2_U3519);
  nand ginst17851 (P2_U8282, P2_FLUSH_REG_SCAN_IN, P2_U3597, P2_U3598);
  nand ginst17852 (P2_U8283, P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P2_U3519);
  nand ginst17853 (P2_U8284, P2_FLUSH_REG_SCAN_IN, P2_U3597, P2_U8090);
  nand ginst17854 (P2_U8285, P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN, P2_U3519);
  nand ginst17855 (P2_U8286, P2_FLUSH_REG_SCAN_IN, P2_U8087);
  nand ginst17856 (P2_U8287, P2_U3616, P2_U4406);
  nand ginst17857 (P2_U8288, P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN, P2_U5581);
  nand ginst17858 (P2_U8289, P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P2_U5581);
  nand ginst17859 (P2_U8290, P2_U4406, P2_U5611);
  nand ginst17860 (P2_U8291, P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN, P2_U5581);
  nand ginst17861 (P2_U8292, P2_U4406, P2_U5619);
  nand ginst17862 (P2_U8293, P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P2_U5581);
  nand ginst17863 (P2_U8294, P2_U4406, P2_U5629);
  nand ginst17864 (P2_U8295, P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN, P2_U5581);
  nand ginst17865 (P2_U8296, P2_U4406, P2_U5637);
  nand ginst17866 (P2_U8297, P2_U3242, P2_U7873);
  nand ginst17867 (P2_U8298, P2_U2616, P2_U7183);
  nand ginst17868 (P2_U8299, P2_U7217, P2_U7873);
  nand ginst17869 (P2_U8300, P2_U2616, P2_U7200);
  nand ginst17870 (P2_U8301, P2_U7251, P2_U7873);
  nand ginst17871 (P2_U8302, P2_U2616, P2_U7234);
  nand ginst17872 (P2_U8303, P2_U7285, P2_U7873);
  nand ginst17873 (P2_U8304, P2_U2616, P2_U7268);
  nand ginst17874 (P2_U8305, P2_U7319, P2_U7873);
  nand ginst17875 (P2_U8306, P2_U2616, P2_U7302);
  nand ginst17876 (P2_U8307, P2_U7353, P2_U7873);
  nand ginst17877 (P2_U8308, P2_U2616, P2_U7336);
  nand ginst17878 (P2_U8309, P2_U7387, P2_U7873);
  nand ginst17879 (P2_U8310, P2_U2616, P2_U7370);
  nand ginst17880 (P2_U8311, P2_U7421, P2_U7873);
  nand ginst17881 (P2_U8312, P2_U2616, P2_U7404);
  nand ginst17882 (P2_U8313, P2_R2256_U5, P2_U3572);
  nand ginst17883 (P2_U8314, P2_R2267_U56, P2_U3242);
  nand ginst17884 (P2_U8315, P2_R2256_U17, P2_U3572);
  nand ginst17885 (P2_U8316, P2_R2267_U19, P2_U3242);
  nand ginst17886 (P2_U8317, P2_R2256_U18, P2_U3572);
  nand ginst17887 (P2_U8318, P2_R2267_U58, P2_U3242);
  nand ginst17888 (P2_U8319, P2_R2256_U19, P2_U3572);
  nand ginst17889 (P2_U8320, P2_R2267_U18, P2_U3242);
  nand ginst17890 (P2_U8321, P2_R2256_U20, P2_U3572);
  nand ginst17891 (P2_U8322, P2_R2267_U60, P2_U3242);
  nand ginst17892 (P2_U8323, P2_R2256_U26, P2_U3572);
  nand ginst17893 (P2_U8324, P2_R2267_U17, P2_U3242);
  nand ginst17894 (P2_U8325, P2_R2256_U22, P2_U3572);
  nand ginst17895 (P2_U8326, P2_R2267_U65, P2_U3242);
  nand ginst17896 (P2_U8327, P2_R2256_U4, P2_U3572);
  nand ginst17897 (P2_U8328, P2_R2267_U43, P2_U3242);
  nand ginst17898 (P2_U8329, P2_R2256_U21, P2_U3572);
  nand ginst17899 (P2_U8330, P2_R2267_U21, P2_U3242);
  nand ginst17900 (P2_U8331, P2_R2219_U24, P2_U2617);
  nand ginst17901 (P2_U8332, P2_EBX_REG_7__SCAN_IN, P2_U7869);
  nand ginst17902 (P2_U8333, P2_R2219_U25, P2_U2617);
  nand ginst17903 (P2_U8334, P2_EBX_REG_6__SCAN_IN, P2_U7869);
  nand ginst17904 (P2_U8335, P2_R2219_U26, P2_U2617);
  nand ginst17905 (P2_U8336, P2_EBX_REG_5__SCAN_IN, P2_U7869);
  nand ginst17906 (P2_U8337, P2_R2219_U27, P2_U2617);
  nand ginst17907 (P2_U8338, P2_EBX_REG_4__SCAN_IN, P2_U7869);
  nand ginst17908 (P2_U8339, P2_R2219_U28, P2_U2617);
  nand ginst17909 (P2_U8340, P2_EBX_REG_3__SCAN_IN, P2_U7869);
  nand ginst17910 (P2_U8341, P2_R2219_U29, P2_U2617);
  nand ginst17911 (P2_U8342, P2_EBX_REG_2__SCAN_IN, P2_U7869);
  nand ginst17912 (P2_U8343, P2_R2219_U30, P2_U2617);
  nand ginst17913 (P2_U8344, P2_EBX_REG_1__SCAN_IN, P2_U7869);
  nand ginst17914 (P2_U8345, P2_R2219_U8, P2_U2617);
  nand ginst17915 (P2_U8346, P2_EBX_REG_0__SCAN_IN, P2_U7869);
  nand ginst17916 (P2_U8347, P2_U3255, P2_U7740);
  nand ginst17917 (P2_U8348, P2_U3525, P2_U7867);
  nand ginst17918 (P2_U8349, P2_R2337_U68, P2_U3284);
  nand ginst17919 (P2_U8350, P2_STATE2_REG_0__SCAN_IN, P2_INSTADDRPOINTER_REG_31__SCAN_IN);
  nand ginst17920 (P2_U8351, P2_R2238_U6, P2_U3283);
  nand ginst17921 (P2_U8352, P2_SUB_450_U6, P2_U4417);
  nand ginst17922 (P2_U8353, P2_R2238_U19, P2_U3283);
  nand ginst17923 (P2_U8354, P2_SUB_450_U17, P2_U4417);
  nand ginst17924 (P2_U8355, P2_R2238_U20, P2_U3283);
  nand ginst17925 (P2_U8356, P2_SUB_450_U18, P2_U4417);
  nand ginst17926 (P2_U8357, P2_R2238_U21, P2_U3283);
  nand ginst17927 (P2_U8358, P2_SUB_450_U19, P2_U4417);
  nand ginst17928 (P2_U8359, P2_R2238_U22, P2_U3283);
  nand ginst17929 (P2_U8360, P2_SUB_450_U20, P2_U4417);
  nand ginst17930 (P2_U8361, P2_R2337_U61, P2_U3284);
  nand ginst17931 (P2_U8362, P2_STATE2_REG_0__SCAN_IN, P2_INSTADDRPOINTER_REG_9__SCAN_IN);
  nand ginst17932 (P2_U8363, P2_R2337_U62, P2_U3284);
  nand ginst17933 (P2_U8364, P2_STATE2_REG_0__SCAN_IN, P2_INSTADDRPOINTER_REG_8__SCAN_IN);
  nand ginst17934 (P2_U8365, P2_R2337_U63, P2_U3284);
  nand ginst17935 (P2_U8366, P2_STATE2_REG_0__SCAN_IN, P2_INSTADDRPOINTER_REG_7__SCAN_IN);
  nand ginst17936 (P2_U8367, P2_R2337_U64, P2_U3284);
  nand ginst17937 (P2_U8368, P2_STATE2_REG_0__SCAN_IN, P2_INSTADDRPOINTER_REG_6__SCAN_IN);
  nand ginst17938 (P2_U8369, P2_R2337_U65, P2_U3284);
  nand ginst17939 (P2_U8370, P2_STATE2_REG_0__SCAN_IN, P2_INSTADDRPOINTER_REG_5__SCAN_IN);
  nand ginst17940 (P2_U8371, P2_R2337_U66, P2_U3284);
  nand ginst17941 (P2_U8372, P2_STATE2_REG_0__SCAN_IN, P2_INSTADDRPOINTER_REG_4__SCAN_IN);
  nand ginst17942 (P2_U8373, P2_R2337_U69, P2_U3284);
  nand ginst17943 (P2_U8374, P2_STATE2_REG_0__SCAN_IN, P2_INSTADDRPOINTER_REG_30__SCAN_IN);
  nand ginst17944 (P2_U8375, P2_R2337_U67, P2_U3284);
  nand ginst17945 (P2_U8376, P2_STATE2_REG_0__SCAN_IN, P2_INSTADDRPOINTER_REG_3__SCAN_IN);
  nand ginst17946 (P2_U8377, P2_R2337_U71, P2_U3284);
  nand ginst17947 (P2_U8378, P2_STATE2_REG_0__SCAN_IN, P2_INSTADDRPOINTER_REG_29__SCAN_IN);
  nand ginst17948 (P2_U8379, P2_R2337_U72, P2_U3284);
  nand ginst17949 (P2_U8380, P2_STATE2_REG_0__SCAN_IN, P2_INSTADDRPOINTER_REG_28__SCAN_IN);
  nand ginst17950 (P2_U8381, P2_R2337_U73, P2_U3284);
  nand ginst17951 (P2_U8382, P2_STATE2_REG_0__SCAN_IN, P2_INSTADDRPOINTER_REG_27__SCAN_IN);
  nand ginst17952 (P2_U8383, P2_R2337_U74, P2_U3284);
  nand ginst17953 (P2_U8384, P2_STATE2_REG_0__SCAN_IN, P2_INSTADDRPOINTER_REG_26__SCAN_IN);
  nand ginst17954 (P2_U8385, P2_R2337_U75, P2_U3284);
  nand ginst17955 (P2_U8386, P2_STATE2_REG_0__SCAN_IN, P2_INSTADDRPOINTER_REG_25__SCAN_IN);
  nand ginst17956 (P2_U8387, P2_R2337_U76, P2_U3284);
  nand ginst17957 (P2_U8388, P2_STATE2_REG_0__SCAN_IN, P2_INSTADDRPOINTER_REG_24__SCAN_IN);
  nand ginst17958 (P2_U8389, P2_R2337_U77, P2_U3284);
  nand ginst17959 (P2_U8390, P2_STATE2_REG_0__SCAN_IN, P2_INSTADDRPOINTER_REG_23__SCAN_IN);
  nand ginst17960 (P2_U8391, P2_R2337_U78, P2_U3284);
  nand ginst17961 (P2_U8392, P2_STATE2_REG_0__SCAN_IN, P2_INSTADDRPOINTER_REG_22__SCAN_IN);
  nand ginst17962 (P2_U8393, P2_R2337_U79, P2_U3284);
  nand ginst17963 (P2_U8394, P2_STATE2_REG_0__SCAN_IN, P2_INSTADDRPOINTER_REG_21__SCAN_IN);
  nand ginst17964 (P2_U8395, P2_R2337_U80, P2_U3284);
  nand ginst17965 (P2_U8396, P2_STATE2_REG_0__SCAN_IN, P2_INSTADDRPOINTER_REG_20__SCAN_IN);
  nand ginst17966 (P2_U8397, P2_R2337_U70, P2_U3284);
  nand ginst17967 (P2_U8398, P2_STATE2_REG_0__SCAN_IN, P2_INSTADDRPOINTER_REG_2__SCAN_IN);
  nand ginst17968 (P2_U8399, P2_R2337_U81, P2_U3284);
  nand ginst17969 (P2_U8400, P2_STATE2_REG_0__SCAN_IN, P2_INSTADDRPOINTER_REG_19__SCAN_IN);
  nand ginst17970 (P2_U8401, P2_R2337_U82, P2_U3284);
  nand ginst17971 (P2_U8402, P2_STATE2_REG_0__SCAN_IN, P2_INSTADDRPOINTER_REG_18__SCAN_IN);
  nand ginst17972 (P2_U8403, P2_R2337_U83, P2_U3284);
  nand ginst17973 (P2_U8404, P2_STATE2_REG_0__SCAN_IN, P2_INSTADDRPOINTER_REG_17__SCAN_IN);
  nand ginst17974 (P2_U8405, P2_R2337_U84, P2_U3284);
  nand ginst17975 (P2_U8406, P2_STATE2_REG_0__SCAN_IN, P2_INSTADDRPOINTER_REG_16__SCAN_IN);
  nand ginst17976 (P2_U8407, P2_R2337_U85, P2_U3284);
  nand ginst17977 (P2_U8408, P2_STATE2_REG_0__SCAN_IN, P2_INSTADDRPOINTER_REG_15__SCAN_IN);
  nand ginst17978 (P2_U8409, P2_R2337_U86, P2_U3284);
  nand ginst17979 (P2_U8410, P2_STATE2_REG_0__SCAN_IN, P2_INSTADDRPOINTER_REG_14__SCAN_IN);
  nand ginst17980 (P2_U8411, P2_R2337_U87, P2_U3284);
  nand ginst17981 (P2_U8412, P2_STATE2_REG_0__SCAN_IN, P2_INSTADDRPOINTER_REG_13__SCAN_IN);
  nand ginst17982 (P2_U8413, P2_R2337_U88, P2_U3284);
  nand ginst17983 (P2_U8414, P2_STATE2_REG_0__SCAN_IN, P2_INSTADDRPOINTER_REG_12__SCAN_IN);
  nand ginst17984 (P2_U8415, P2_R2337_U89, P2_U3284);
  nand ginst17985 (P2_U8416, P2_STATE2_REG_0__SCAN_IN, P2_INSTADDRPOINTER_REG_11__SCAN_IN);
  nand ginst17986 (P2_U8417, P2_R2337_U90, P2_U3284);
  nand ginst17987 (P2_U8418, P2_STATE2_REG_0__SCAN_IN, P2_INSTADDRPOINTER_REG_10__SCAN_IN);
  nand ginst17988 (P2_U8419, P2_R2337_U4, P2_U3284);
  nand ginst17989 (P2_U8420, P2_STATE2_REG_0__SCAN_IN, P2_INSTADDRPOINTER_REG_1__SCAN_IN);
  nand ginst17990 (P2_U8421, P2_PHYADDRPOINTER_REG_0__SCAN_IN, P2_U3284);
  nand ginst17991 (P2_U8422, P2_STATE2_REG_0__SCAN_IN, P2_INSTADDRPOINTER_REG_0__SCAN_IN);
  nand ginst17992 (P2_U8423, P2_R2238_U6, P2_U3269);
  nand ginst17993 (P2_U8424, P2_STATE2_REG_1__SCAN_IN, P2_U2615);
  nand ginst17994 (P2_U8425, P2_R2238_U19, P2_U3269);
  nand ginst17995 (P2_U8426, P2_STATE2_REG_1__SCAN_IN, P2_U2615);
  nand ginst17996 (P2_U8427, P2_R2238_U20, P2_U3269);
  nand ginst17997 (P2_U8428, P2_STATE2_REG_1__SCAN_IN, P2_SUB_589_U8);
  nand ginst17998 (P2_U8429, P2_R2238_U21, P2_U3269);
  nand ginst17999 (P2_U8430, P2_STATE2_REG_1__SCAN_IN, P2_SUB_589_U9);
  nand ginst18000 (P2_U8431, P2_R2238_U22, P2_U3269);
  nand ginst18001 (P2_U8432, P2_STATE2_REG_1__SCAN_IN, P2_SUB_589_U6);
  nand ginst18002 (P2_U8433, P2_R2238_U7, P2_U3269);
  nand ginst18003 (P2_U8434, P2_STATE2_REG_1__SCAN_IN, P2_SUB_589_U7);
  nand ginst18004 (P3_ADD_315_U10, P3_PHYADDRPOINTER_REG_5__SCAN_IN, P3_ADD_315_U92);
  not ginst18005 (P3_ADD_315_U100, P3_ADD_315_U24);
  not ginst18006 (P3_ADD_315_U101, P3_ADD_315_U26);
  not ginst18007 (P3_ADD_315_U102, P3_ADD_315_U28);
  not ginst18008 (P3_ADD_315_U103, P3_ADD_315_U30);
  not ginst18009 (P3_ADD_315_U104, P3_ADD_315_U32);
  not ginst18010 (P3_ADD_315_U105, P3_ADD_315_U34);
  not ginst18011 (P3_ADD_315_U106, P3_ADD_315_U36);
  not ginst18012 (P3_ADD_315_U107, P3_ADD_315_U38);
  not ginst18013 (P3_ADD_315_U108, P3_ADD_315_U40);
  not ginst18014 (P3_ADD_315_U109, P3_ADD_315_U42);
  not ginst18015 (P3_ADD_315_U11, P3_PHYADDRPOINTER_REG_6__SCAN_IN);
  not ginst18016 (P3_ADD_315_U110, P3_ADD_315_U44);
  not ginst18017 (P3_ADD_315_U111, P3_ADD_315_U46);
  not ginst18018 (P3_ADD_315_U112, P3_ADD_315_U48);
  not ginst18019 (P3_ADD_315_U113, P3_ADD_315_U50);
  not ginst18020 (P3_ADD_315_U114, P3_ADD_315_U52);
  not ginst18021 (P3_ADD_315_U115, P3_ADD_315_U54);
  not ginst18022 (P3_ADD_315_U116, P3_ADD_315_U56);
  not ginst18023 (P3_ADD_315_U117, P3_ADD_315_U58);
  not ginst18024 (P3_ADD_315_U118, P3_ADD_315_U90);
  nand ginst18025 (P3_ADD_315_U119, P3_PHYADDRPOINTER_REG_9__SCAN_IN, P3_ADD_315_U17);
  nand ginst18026 (P3_ADD_315_U12, P3_PHYADDRPOINTER_REG_6__SCAN_IN, P3_ADD_315_U93);
  nand ginst18027 (P3_ADD_315_U120, P3_ADD_315_U16, P3_ADD_315_U96);
  nand ginst18028 (P3_ADD_315_U121, P3_PHYADDRPOINTER_REG_8__SCAN_IN, P3_ADD_315_U14);
  nand ginst18029 (P3_ADD_315_U122, P3_ADD_315_U15, P3_ADD_315_U95);
  nand ginst18030 (P3_ADD_315_U123, P3_PHYADDRPOINTER_REG_7__SCAN_IN, P3_ADD_315_U12);
  nand ginst18031 (P3_ADD_315_U124, P3_ADD_315_U13, P3_ADD_315_U94);
  nand ginst18032 (P3_ADD_315_U125, P3_PHYADDRPOINTER_REG_6__SCAN_IN, P3_ADD_315_U10);
  nand ginst18033 (P3_ADD_315_U126, P3_ADD_315_U11, P3_ADD_315_U93);
  nand ginst18034 (P3_ADD_315_U127, P3_PHYADDRPOINTER_REG_5__SCAN_IN, P3_ADD_315_U8);
  nand ginst18035 (P3_ADD_315_U128, P3_ADD_315_U9, P3_ADD_315_U92);
  nand ginst18036 (P3_ADD_315_U129, P3_PHYADDRPOINTER_REG_4__SCAN_IN, P3_ADD_315_U6);
  not ginst18037 (P3_ADD_315_U13, P3_PHYADDRPOINTER_REG_7__SCAN_IN);
  nand ginst18038 (P3_ADD_315_U130, P3_ADD_315_U7, P3_ADD_315_U91);
  nand ginst18039 (P3_ADD_315_U131, P3_PHYADDRPOINTER_REG_3__SCAN_IN, P3_ADD_315_U4);
  nand ginst18040 (P3_ADD_315_U132, P3_PHYADDRPOINTER_REG_2__SCAN_IN, P3_ADD_315_U5);
  nand ginst18041 (P3_ADD_315_U133, P3_PHYADDRPOINTER_REG_31__SCAN_IN, P3_ADD_315_U90);
  nand ginst18042 (P3_ADD_315_U134, P3_ADD_315_U118, P3_ADD_315_U89);
  nand ginst18043 (P3_ADD_315_U135, P3_PHYADDRPOINTER_REG_30__SCAN_IN, P3_ADD_315_U58);
  nand ginst18044 (P3_ADD_315_U136, P3_ADD_315_U117, P3_ADD_315_U59);
  nand ginst18045 (P3_ADD_315_U137, P3_PHYADDRPOINTER_REG_29__SCAN_IN, P3_ADD_315_U56);
  nand ginst18046 (P3_ADD_315_U138, P3_ADD_315_U116, P3_ADD_315_U57);
  nand ginst18047 (P3_ADD_315_U139, P3_PHYADDRPOINTER_REG_28__SCAN_IN, P3_ADD_315_U54);
  nand ginst18048 (P3_ADD_315_U14, P3_PHYADDRPOINTER_REG_7__SCAN_IN, P3_ADD_315_U94);
  nand ginst18049 (P3_ADD_315_U140, P3_ADD_315_U115, P3_ADD_315_U55);
  nand ginst18050 (P3_ADD_315_U141, P3_PHYADDRPOINTER_REG_27__SCAN_IN, P3_ADD_315_U52);
  nand ginst18051 (P3_ADD_315_U142, P3_ADD_315_U114, P3_ADD_315_U53);
  nand ginst18052 (P3_ADD_315_U143, P3_PHYADDRPOINTER_REG_26__SCAN_IN, P3_ADD_315_U50);
  nand ginst18053 (P3_ADD_315_U144, P3_ADD_315_U113, P3_ADD_315_U51);
  nand ginst18054 (P3_ADD_315_U145, P3_PHYADDRPOINTER_REG_25__SCAN_IN, P3_ADD_315_U48);
  nand ginst18055 (P3_ADD_315_U146, P3_ADD_315_U112, P3_ADD_315_U49);
  nand ginst18056 (P3_ADD_315_U147, P3_PHYADDRPOINTER_REG_24__SCAN_IN, P3_ADD_315_U46);
  nand ginst18057 (P3_ADD_315_U148, P3_ADD_315_U111, P3_ADD_315_U47);
  nand ginst18058 (P3_ADD_315_U149, P3_PHYADDRPOINTER_REG_23__SCAN_IN, P3_ADD_315_U44);
  not ginst18059 (P3_ADD_315_U15, P3_PHYADDRPOINTER_REG_8__SCAN_IN);
  nand ginst18060 (P3_ADD_315_U150, P3_ADD_315_U110, P3_ADD_315_U45);
  nand ginst18061 (P3_ADD_315_U151, P3_PHYADDRPOINTER_REG_22__SCAN_IN, P3_ADD_315_U42);
  nand ginst18062 (P3_ADD_315_U152, P3_ADD_315_U109, P3_ADD_315_U43);
  nand ginst18063 (P3_ADD_315_U153, P3_PHYADDRPOINTER_REG_21__SCAN_IN, P3_ADD_315_U40);
  nand ginst18064 (P3_ADD_315_U154, P3_ADD_315_U108, P3_ADD_315_U41);
  nand ginst18065 (P3_ADD_315_U155, P3_PHYADDRPOINTER_REG_20__SCAN_IN, P3_ADD_315_U38);
  nand ginst18066 (P3_ADD_315_U156, P3_ADD_315_U107, P3_ADD_315_U39);
  nand ginst18067 (P3_ADD_315_U157, P3_PHYADDRPOINTER_REG_19__SCAN_IN, P3_ADD_315_U36);
  nand ginst18068 (P3_ADD_315_U158, P3_ADD_315_U106, P3_ADD_315_U37);
  nand ginst18069 (P3_ADD_315_U159, P3_PHYADDRPOINTER_REG_18__SCAN_IN, P3_ADD_315_U34);
  not ginst18070 (P3_ADD_315_U16, P3_PHYADDRPOINTER_REG_9__SCAN_IN);
  nand ginst18071 (P3_ADD_315_U160, P3_ADD_315_U105, P3_ADD_315_U35);
  nand ginst18072 (P3_ADD_315_U161, P3_PHYADDRPOINTER_REG_17__SCAN_IN, P3_ADD_315_U32);
  nand ginst18073 (P3_ADD_315_U162, P3_ADD_315_U104, P3_ADD_315_U33);
  nand ginst18074 (P3_ADD_315_U163, P3_PHYADDRPOINTER_REG_16__SCAN_IN, P3_ADD_315_U30);
  nand ginst18075 (P3_ADD_315_U164, P3_ADD_315_U103, P3_ADD_315_U31);
  nand ginst18076 (P3_ADD_315_U165, P3_PHYADDRPOINTER_REG_15__SCAN_IN, P3_ADD_315_U28);
  nand ginst18077 (P3_ADD_315_U166, P3_ADD_315_U102, P3_ADD_315_U29);
  nand ginst18078 (P3_ADD_315_U167, P3_PHYADDRPOINTER_REG_14__SCAN_IN, P3_ADD_315_U26);
  nand ginst18079 (P3_ADD_315_U168, P3_ADD_315_U101, P3_ADD_315_U27);
  nand ginst18080 (P3_ADD_315_U169, P3_PHYADDRPOINTER_REG_13__SCAN_IN, P3_ADD_315_U24);
  nand ginst18081 (P3_ADD_315_U17, P3_PHYADDRPOINTER_REG_8__SCAN_IN, P3_ADD_315_U95);
  nand ginst18082 (P3_ADD_315_U170, P3_ADD_315_U100, P3_ADD_315_U25);
  nand ginst18083 (P3_ADD_315_U171, P3_PHYADDRPOINTER_REG_12__SCAN_IN, P3_ADD_315_U22);
  nand ginst18084 (P3_ADD_315_U172, P3_ADD_315_U23, P3_ADD_315_U99);
  nand ginst18085 (P3_ADD_315_U173, P3_PHYADDRPOINTER_REG_11__SCAN_IN, P3_ADD_315_U20);
  nand ginst18086 (P3_ADD_315_U174, P3_ADD_315_U21, P3_ADD_315_U98);
  nand ginst18087 (P3_ADD_315_U175, P3_PHYADDRPOINTER_REG_10__SCAN_IN, P3_ADD_315_U18);
  nand ginst18088 (P3_ADD_315_U176, P3_ADD_315_U19, P3_ADD_315_U97);
  nand ginst18089 (P3_ADD_315_U18, P3_PHYADDRPOINTER_REG_9__SCAN_IN, P3_ADD_315_U96);
  not ginst18090 (P3_ADD_315_U19, P3_PHYADDRPOINTER_REG_10__SCAN_IN);
  nand ginst18091 (P3_ADD_315_U20, P3_PHYADDRPOINTER_REG_10__SCAN_IN, P3_ADD_315_U97);
  not ginst18092 (P3_ADD_315_U21, P3_PHYADDRPOINTER_REG_11__SCAN_IN);
  nand ginst18093 (P3_ADD_315_U22, P3_PHYADDRPOINTER_REG_11__SCAN_IN, P3_ADD_315_U98);
  not ginst18094 (P3_ADD_315_U23, P3_PHYADDRPOINTER_REG_12__SCAN_IN);
  nand ginst18095 (P3_ADD_315_U24, P3_PHYADDRPOINTER_REG_12__SCAN_IN, P3_ADD_315_U99);
  not ginst18096 (P3_ADD_315_U25, P3_PHYADDRPOINTER_REG_13__SCAN_IN);
  nand ginst18097 (P3_ADD_315_U26, P3_PHYADDRPOINTER_REG_13__SCAN_IN, P3_ADD_315_U100);
  not ginst18098 (P3_ADD_315_U27, P3_PHYADDRPOINTER_REG_14__SCAN_IN);
  nand ginst18099 (P3_ADD_315_U28, P3_PHYADDRPOINTER_REG_14__SCAN_IN, P3_ADD_315_U101);
  not ginst18100 (P3_ADD_315_U29, P3_PHYADDRPOINTER_REG_15__SCAN_IN);
  nand ginst18101 (P3_ADD_315_U30, P3_PHYADDRPOINTER_REG_15__SCAN_IN, P3_ADD_315_U102);
  not ginst18102 (P3_ADD_315_U31, P3_PHYADDRPOINTER_REG_16__SCAN_IN);
  nand ginst18103 (P3_ADD_315_U32, P3_PHYADDRPOINTER_REG_16__SCAN_IN, P3_ADD_315_U103);
  not ginst18104 (P3_ADD_315_U33, P3_PHYADDRPOINTER_REG_17__SCAN_IN);
  nand ginst18105 (P3_ADD_315_U34, P3_PHYADDRPOINTER_REG_17__SCAN_IN, P3_ADD_315_U104);
  not ginst18106 (P3_ADD_315_U35, P3_PHYADDRPOINTER_REG_18__SCAN_IN);
  nand ginst18107 (P3_ADD_315_U36, P3_PHYADDRPOINTER_REG_18__SCAN_IN, P3_ADD_315_U105);
  not ginst18108 (P3_ADD_315_U37, P3_PHYADDRPOINTER_REG_19__SCAN_IN);
  nand ginst18109 (P3_ADD_315_U38, P3_PHYADDRPOINTER_REG_19__SCAN_IN, P3_ADD_315_U106);
  not ginst18110 (P3_ADD_315_U39, P3_PHYADDRPOINTER_REG_20__SCAN_IN);
  not ginst18111 (P3_ADD_315_U4, P3_PHYADDRPOINTER_REG_2__SCAN_IN);
  nand ginst18112 (P3_ADD_315_U40, P3_PHYADDRPOINTER_REG_20__SCAN_IN, P3_ADD_315_U107);
  not ginst18113 (P3_ADD_315_U41, P3_PHYADDRPOINTER_REG_21__SCAN_IN);
  nand ginst18114 (P3_ADD_315_U42, P3_PHYADDRPOINTER_REG_21__SCAN_IN, P3_ADD_315_U108);
  not ginst18115 (P3_ADD_315_U43, P3_PHYADDRPOINTER_REG_22__SCAN_IN);
  nand ginst18116 (P3_ADD_315_U44, P3_PHYADDRPOINTER_REG_22__SCAN_IN, P3_ADD_315_U109);
  not ginst18117 (P3_ADD_315_U45, P3_PHYADDRPOINTER_REG_23__SCAN_IN);
  nand ginst18118 (P3_ADD_315_U46, P3_PHYADDRPOINTER_REG_23__SCAN_IN, P3_ADD_315_U110);
  not ginst18119 (P3_ADD_315_U47, P3_PHYADDRPOINTER_REG_24__SCAN_IN);
  nand ginst18120 (P3_ADD_315_U48, P3_PHYADDRPOINTER_REG_24__SCAN_IN, P3_ADD_315_U111);
  not ginst18121 (P3_ADD_315_U49, P3_PHYADDRPOINTER_REG_25__SCAN_IN);
  not ginst18122 (P3_ADD_315_U5, P3_PHYADDRPOINTER_REG_3__SCAN_IN);
  nand ginst18123 (P3_ADD_315_U50, P3_PHYADDRPOINTER_REG_25__SCAN_IN, P3_ADD_315_U112);
  not ginst18124 (P3_ADD_315_U51, P3_PHYADDRPOINTER_REG_26__SCAN_IN);
  nand ginst18125 (P3_ADD_315_U52, P3_PHYADDRPOINTER_REG_26__SCAN_IN, P3_ADD_315_U113);
  not ginst18126 (P3_ADD_315_U53, P3_PHYADDRPOINTER_REG_27__SCAN_IN);
  nand ginst18127 (P3_ADD_315_U54, P3_PHYADDRPOINTER_REG_27__SCAN_IN, P3_ADD_315_U114);
  not ginst18128 (P3_ADD_315_U55, P3_PHYADDRPOINTER_REG_28__SCAN_IN);
  nand ginst18129 (P3_ADD_315_U56, P3_PHYADDRPOINTER_REG_28__SCAN_IN, P3_ADD_315_U115);
  not ginst18130 (P3_ADD_315_U57, P3_PHYADDRPOINTER_REG_29__SCAN_IN);
  nand ginst18131 (P3_ADD_315_U58, P3_PHYADDRPOINTER_REG_29__SCAN_IN, P3_ADD_315_U116);
  not ginst18132 (P3_ADD_315_U59, P3_PHYADDRPOINTER_REG_30__SCAN_IN);
  nand ginst18133 (P3_ADD_315_U6, P3_PHYADDRPOINTER_REG_2__SCAN_IN, P3_PHYADDRPOINTER_REG_3__SCAN_IN);
  nand ginst18134 (P3_ADD_315_U60, P3_ADD_315_U119, P3_ADD_315_U120);
  nand ginst18135 (P3_ADD_315_U61, P3_ADD_315_U121, P3_ADD_315_U122);
  nand ginst18136 (P3_ADD_315_U62, P3_ADD_315_U123, P3_ADD_315_U124);
  nand ginst18137 (P3_ADD_315_U63, P3_ADD_315_U125, P3_ADD_315_U126);
  nand ginst18138 (P3_ADD_315_U64, P3_ADD_315_U127, P3_ADD_315_U128);
  nand ginst18139 (P3_ADD_315_U65, P3_ADD_315_U129, P3_ADD_315_U130);
  nand ginst18140 (P3_ADD_315_U66, P3_ADD_315_U131, P3_ADD_315_U132);
  nand ginst18141 (P3_ADD_315_U67, P3_ADD_315_U133, P3_ADD_315_U134);
  nand ginst18142 (P3_ADD_315_U68, P3_ADD_315_U135, P3_ADD_315_U136);
  nand ginst18143 (P3_ADD_315_U69, P3_ADD_315_U137, P3_ADD_315_U138);
  not ginst18144 (P3_ADD_315_U7, P3_PHYADDRPOINTER_REG_4__SCAN_IN);
  nand ginst18145 (P3_ADD_315_U70, P3_ADD_315_U139, P3_ADD_315_U140);
  nand ginst18146 (P3_ADD_315_U71, P3_ADD_315_U141, P3_ADD_315_U142);
  nand ginst18147 (P3_ADD_315_U72, P3_ADD_315_U143, P3_ADD_315_U144);
  nand ginst18148 (P3_ADD_315_U73, P3_ADD_315_U145, P3_ADD_315_U146);
  nand ginst18149 (P3_ADD_315_U74, P3_ADD_315_U147, P3_ADD_315_U148);
  nand ginst18150 (P3_ADD_315_U75, P3_ADD_315_U149, P3_ADD_315_U150);
  nand ginst18151 (P3_ADD_315_U76, P3_ADD_315_U151, P3_ADD_315_U152);
  nand ginst18152 (P3_ADD_315_U77, P3_ADD_315_U153, P3_ADD_315_U154);
  nand ginst18153 (P3_ADD_315_U78, P3_ADD_315_U155, P3_ADD_315_U156);
  nand ginst18154 (P3_ADD_315_U79, P3_ADD_315_U157, P3_ADD_315_U158);
  nand ginst18155 (P3_ADD_315_U8, P3_PHYADDRPOINTER_REG_4__SCAN_IN, P3_ADD_315_U91);
  nand ginst18156 (P3_ADD_315_U80, P3_ADD_315_U159, P3_ADD_315_U160);
  nand ginst18157 (P3_ADD_315_U81, P3_ADD_315_U161, P3_ADD_315_U162);
  nand ginst18158 (P3_ADD_315_U82, P3_ADD_315_U163, P3_ADD_315_U164);
  nand ginst18159 (P3_ADD_315_U83, P3_ADD_315_U165, P3_ADD_315_U166);
  nand ginst18160 (P3_ADD_315_U84, P3_ADD_315_U167, P3_ADD_315_U168);
  nand ginst18161 (P3_ADD_315_U85, P3_ADD_315_U169, P3_ADD_315_U170);
  nand ginst18162 (P3_ADD_315_U86, P3_ADD_315_U171, P3_ADD_315_U172);
  nand ginst18163 (P3_ADD_315_U87, P3_ADD_315_U173, P3_ADD_315_U174);
  nand ginst18164 (P3_ADD_315_U88, P3_ADD_315_U175, P3_ADD_315_U176);
  not ginst18165 (P3_ADD_315_U89, P3_PHYADDRPOINTER_REG_31__SCAN_IN);
  not ginst18166 (P3_ADD_315_U9, P3_PHYADDRPOINTER_REG_5__SCAN_IN);
  nand ginst18167 (P3_ADD_315_U90, P3_PHYADDRPOINTER_REG_30__SCAN_IN, P3_ADD_315_U117);
  not ginst18168 (P3_ADD_315_U91, P3_ADD_315_U6);
  not ginst18169 (P3_ADD_315_U92, P3_ADD_315_U8);
  not ginst18170 (P3_ADD_315_U93, P3_ADD_315_U10);
  not ginst18171 (P3_ADD_315_U94, P3_ADD_315_U12);
  not ginst18172 (P3_ADD_315_U95, P3_ADD_315_U14);
  not ginst18173 (P3_ADD_315_U96, P3_ADD_315_U17);
  not ginst18174 (P3_ADD_315_U97, P3_ADD_315_U18);
  not ginst18175 (P3_ADD_315_U98, P3_ADD_315_U20);
  not ginst18176 (P3_ADD_315_U99, P3_ADD_315_U22);
  nand ginst18177 (P3_ADD_318_U10, P3_PHYADDRPOINTER_REG_4__SCAN_IN, P3_ADD_318_U95);
  not ginst18178 (P3_ADD_318_U100, P3_ADD_318_U19);
  not ginst18179 (P3_ADD_318_U101, P3_ADD_318_U20);
  not ginst18180 (P3_ADD_318_U102, P3_ADD_318_U22);
  not ginst18181 (P3_ADD_318_U103, P3_ADD_318_U24);
  not ginst18182 (P3_ADD_318_U104, P3_ADD_318_U26);
  not ginst18183 (P3_ADD_318_U105, P3_ADD_318_U28);
  not ginst18184 (P3_ADD_318_U106, P3_ADD_318_U30);
  not ginst18185 (P3_ADD_318_U107, P3_ADD_318_U32);
  not ginst18186 (P3_ADD_318_U108, P3_ADD_318_U34);
  not ginst18187 (P3_ADD_318_U109, P3_ADD_318_U36);
  not ginst18188 (P3_ADD_318_U11, P3_PHYADDRPOINTER_REG_5__SCAN_IN);
  not ginst18189 (P3_ADD_318_U110, P3_ADD_318_U38);
  not ginst18190 (P3_ADD_318_U111, P3_ADD_318_U40);
  not ginst18191 (P3_ADD_318_U112, P3_ADD_318_U42);
  not ginst18192 (P3_ADD_318_U113, P3_ADD_318_U44);
  not ginst18193 (P3_ADD_318_U114, P3_ADD_318_U46);
  not ginst18194 (P3_ADD_318_U115, P3_ADD_318_U48);
  not ginst18195 (P3_ADD_318_U116, P3_ADD_318_U50);
  not ginst18196 (P3_ADD_318_U117, P3_ADD_318_U52);
  not ginst18197 (P3_ADD_318_U118, P3_ADD_318_U54);
  not ginst18198 (P3_ADD_318_U119, P3_ADD_318_U56);
  nand ginst18199 (P3_ADD_318_U12, P3_PHYADDRPOINTER_REG_5__SCAN_IN, P3_ADD_318_U96);
  not ginst18200 (P3_ADD_318_U120, P3_ADD_318_U58);
  not ginst18201 (P3_ADD_318_U121, P3_ADD_318_U60);
  not ginst18202 (P3_ADD_318_U122, P3_ADD_318_U93);
  nand ginst18203 (P3_ADD_318_U123, P3_PHYADDRPOINTER_REG_9__SCAN_IN, P3_ADD_318_U19);
  nand ginst18204 (P3_ADD_318_U124, P3_ADD_318_U100, P3_ADD_318_U18);
  nand ginst18205 (P3_ADD_318_U125, P3_PHYADDRPOINTER_REG_8__SCAN_IN, P3_ADD_318_U16);
  nand ginst18206 (P3_ADD_318_U126, P3_ADD_318_U17, P3_ADD_318_U99);
  nand ginst18207 (P3_ADD_318_U127, P3_PHYADDRPOINTER_REG_7__SCAN_IN, P3_ADD_318_U14);
  nand ginst18208 (P3_ADD_318_U128, P3_ADD_318_U15, P3_ADD_318_U98);
  nand ginst18209 (P3_ADD_318_U129, P3_PHYADDRPOINTER_REG_6__SCAN_IN, P3_ADD_318_U12);
  not ginst18210 (P3_ADD_318_U13, P3_PHYADDRPOINTER_REG_6__SCAN_IN);
  nand ginst18211 (P3_ADD_318_U130, P3_ADD_318_U13, P3_ADD_318_U97);
  nand ginst18212 (P3_ADD_318_U131, P3_PHYADDRPOINTER_REG_5__SCAN_IN, P3_ADD_318_U10);
  nand ginst18213 (P3_ADD_318_U132, P3_ADD_318_U11, P3_ADD_318_U96);
  nand ginst18214 (P3_ADD_318_U133, P3_PHYADDRPOINTER_REG_4__SCAN_IN, P3_ADD_318_U8);
  nand ginst18215 (P3_ADD_318_U134, P3_ADD_318_U9, P3_ADD_318_U95);
  nand ginst18216 (P3_ADD_318_U135, P3_PHYADDRPOINTER_REG_3__SCAN_IN, P3_ADD_318_U6);
  nand ginst18217 (P3_ADD_318_U136, P3_ADD_318_U7, P3_ADD_318_U94);
  nand ginst18218 (P3_ADD_318_U137, P3_PHYADDRPOINTER_REG_31__SCAN_IN, P3_ADD_318_U93);
  nand ginst18219 (P3_ADD_318_U138, P3_ADD_318_U122, P3_ADD_318_U92);
  nand ginst18220 (P3_ADD_318_U139, P3_PHYADDRPOINTER_REG_30__SCAN_IN, P3_ADD_318_U60);
  nand ginst18221 (P3_ADD_318_U14, P3_PHYADDRPOINTER_REG_6__SCAN_IN, P3_ADD_318_U97);
  nand ginst18222 (P3_ADD_318_U140, P3_ADD_318_U121, P3_ADD_318_U61);
  nand ginst18223 (P3_ADD_318_U141, P3_PHYADDRPOINTER_REG_2__SCAN_IN, P3_ADD_318_U4);
  nand ginst18224 (P3_ADD_318_U142, P3_PHYADDRPOINTER_REG_1__SCAN_IN, P3_ADD_318_U5);
  nand ginst18225 (P3_ADD_318_U143, P3_PHYADDRPOINTER_REG_29__SCAN_IN, P3_ADD_318_U58);
  nand ginst18226 (P3_ADD_318_U144, P3_ADD_318_U120, P3_ADD_318_U59);
  nand ginst18227 (P3_ADD_318_U145, P3_PHYADDRPOINTER_REG_28__SCAN_IN, P3_ADD_318_U56);
  nand ginst18228 (P3_ADD_318_U146, P3_ADD_318_U119, P3_ADD_318_U57);
  nand ginst18229 (P3_ADD_318_U147, P3_PHYADDRPOINTER_REG_27__SCAN_IN, P3_ADD_318_U54);
  nand ginst18230 (P3_ADD_318_U148, P3_ADD_318_U118, P3_ADD_318_U55);
  nand ginst18231 (P3_ADD_318_U149, P3_PHYADDRPOINTER_REG_26__SCAN_IN, P3_ADD_318_U52);
  not ginst18232 (P3_ADD_318_U15, P3_PHYADDRPOINTER_REG_7__SCAN_IN);
  nand ginst18233 (P3_ADD_318_U150, P3_ADD_318_U117, P3_ADD_318_U53);
  nand ginst18234 (P3_ADD_318_U151, P3_PHYADDRPOINTER_REG_25__SCAN_IN, P3_ADD_318_U50);
  nand ginst18235 (P3_ADD_318_U152, P3_ADD_318_U116, P3_ADD_318_U51);
  nand ginst18236 (P3_ADD_318_U153, P3_PHYADDRPOINTER_REG_24__SCAN_IN, P3_ADD_318_U48);
  nand ginst18237 (P3_ADD_318_U154, P3_ADD_318_U115, P3_ADD_318_U49);
  nand ginst18238 (P3_ADD_318_U155, P3_PHYADDRPOINTER_REG_23__SCAN_IN, P3_ADD_318_U46);
  nand ginst18239 (P3_ADD_318_U156, P3_ADD_318_U114, P3_ADD_318_U47);
  nand ginst18240 (P3_ADD_318_U157, P3_PHYADDRPOINTER_REG_22__SCAN_IN, P3_ADD_318_U44);
  nand ginst18241 (P3_ADD_318_U158, P3_ADD_318_U113, P3_ADD_318_U45);
  nand ginst18242 (P3_ADD_318_U159, P3_PHYADDRPOINTER_REG_21__SCAN_IN, P3_ADD_318_U42);
  nand ginst18243 (P3_ADD_318_U16, P3_PHYADDRPOINTER_REG_7__SCAN_IN, P3_ADD_318_U98);
  nand ginst18244 (P3_ADD_318_U160, P3_ADD_318_U112, P3_ADD_318_U43);
  nand ginst18245 (P3_ADD_318_U161, P3_PHYADDRPOINTER_REG_20__SCAN_IN, P3_ADD_318_U40);
  nand ginst18246 (P3_ADD_318_U162, P3_ADD_318_U111, P3_ADD_318_U41);
  nand ginst18247 (P3_ADD_318_U163, P3_PHYADDRPOINTER_REG_19__SCAN_IN, P3_ADD_318_U38);
  nand ginst18248 (P3_ADD_318_U164, P3_ADD_318_U110, P3_ADD_318_U39);
  nand ginst18249 (P3_ADD_318_U165, P3_PHYADDRPOINTER_REG_18__SCAN_IN, P3_ADD_318_U36);
  nand ginst18250 (P3_ADD_318_U166, P3_ADD_318_U109, P3_ADD_318_U37);
  nand ginst18251 (P3_ADD_318_U167, P3_PHYADDRPOINTER_REG_17__SCAN_IN, P3_ADD_318_U34);
  nand ginst18252 (P3_ADD_318_U168, P3_ADD_318_U108, P3_ADD_318_U35);
  nand ginst18253 (P3_ADD_318_U169, P3_PHYADDRPOINTER_REG_16__SCAN_IN, P3_ADD_318_U32);
  not ginst18254 (P3_ADD_318_U17, P3_PHYADDRPOINTER_REG_8__SCAN_IN);
  nand ginst18255 (P3_ADD_318_U170, P3_ADD_318_U107, P3_ADD_318_U33);
  nand ginst18256 (P3_ADD_318_U171, P3_PHYADDRPOINTER_REG_15__SCAN_IN, P3_ADD_318_U30);
  nand ginst18257 (P3_ADD_318_U172, P3_ADD_318_U106, P3_ADD_318_U31);
  nand ginst18258 (P3_ADD_318_U173, P3_PHYADDRPOINTER_REG_14__SCAN_IN, P3_ADD_318_U28);
  nand ginst18259 (P3_ADD_318_U174, P3_ADD_318_U105, P3_ADD_318_U29);
  nand ginst18260 (P3_ADD_318_U175, P3_PHYADDRPOINTER_REG_13__SCAN_IN, P3_ADD_318_U26);
  nand ginst18261 (P3_ADD_318_U176, P3_ADD_318_U104, P3_ADD_318_U27);
  nand ginst18262 (P3_ADD_318_U177, P3_PHYADDRPOINTER_REG_12__SCAN_IN, P3_ADD_318_U24);
  nand ginst18263 (P3_ADD_318_U178, P3_ADD_318_U103, P3_ADD_318_U25);
  nand ginst18264 (P3_ADD_318_U179, P3_PHYADDRPOINTER_REG_11__SCAN_IN, P3_ADD_318_U22);
  not ginst18265 (P3_ADD_318_U18, P3_PHYADDRPOINTER_REG_9__SCAN_IN);
  nand ginst18266 (P3_ADD_318_U180, P3_ADD_318_U102, P3_ADD_318_U23);
  nand ginst18267 (P3_ADD_318_U181, P3_PHYADDRPOINTER_REG_10__SCAN_IN, P3_ADD_318_U20);
  nand ginst18268 (P3_ADD_318_U182, P3_ADD_318_U101, P3_ADD_318_U21);
  nand ginst18269 (P3_ADD_318_U19, P3_PHYADDRPOINTER_REG_8__SCAN_IN, P3_ADD_318_U99);
  nand ginst18270 (P3_ADD_318_U20, P3_PHYADDRPOINTER_REG_9__SCAN_IN, P3_ADD_318_U100);
  not ginst18271 (P3_ADD_318_U21, P3_PHYADDRPOINTER_REG_10__SCAN_IN);
  nand ginst18272 (P3_ADD_318_U22, P3_PHYADDRPOINTER_REG_10__SCAN_IN, P3_ADD_318_U101);
  not ginst18273 (P3_ADD_318_U23, P3_PHYADDRPOINTER_REG_11__SCAN_IN);
  nand ginst18274 (P3_ADD_318_U24, P3_PHYADDRPOINTER_REG_11__SCAN_IN, P3_ADD_318_U102);
  not ginst18275 (P3_ADD_318_U25, P3_PHYADDRPOINTER_REG_12__SCAN_IN);
  nand ginst18276 (P3_ADD_318_U26, P3_PHYADDRPOINTER_REG_12__SCAN_IN, P3_ADD_318_U103);
  not ginst18277 (P3_ADD_318_U27, P3_PHYADDRPOINTER_REG_13__SCAN_IN);
  nand ginst18278 (P3_ADD_318_U28, P3_PHYADDRPOINTER_REG_13__SCAN_IN, P3_ADD_318_U104);
  not ginst18279 (P3_ADD_318_U29, P3_PHYADDRPOINTER_REG_14__SCAN_IN);
  nand ginst18280 (P3_ADD_318_U30, P3_PHYADDRPOINTER_REG_14__SCAN_IN, P3_ADD_318_U105);
  not ginst18281 (P3_ADD_318_U31, P3_PHYADDRPOINTER_REG_15__SCAN_IN);
  nand ginst18282 (P3_ADD_318_U32, P3_PHYADDRPOINTER_REG_15__SCAN_IN, P3_ADD_318_U106);
  not ginst18283 (P3_ADD_318_U33, P3_PHYADDRPOINTER_REG_16__SCAN_IN);
  nand ginst18284 (P3_ADD_318_U34, P3_PHYADDRPOINTER_REG_16__SCAN_IN, P3_ADD_318_U107);
  not ginst18285 (P3_ADD_318_U35, P3_PHYADDRPOINTER_REG_17__SCAN_IN);
  nand ginst18286 (P3_ADD_318_U36, P3_PHYADDRPOINTER_REG_17__SCAN_IN, P3_ADD_318_U108);
  not ginst18287 (P3_ADD_318_U37, P3_PHYADDRPOINTER_REG_18__SCAN_IN);
  nand ginst18288 (P3_ADD_318_U38, P3_PHYADDRPOINTER_REG_18__SCAN_IN, P3_ADD_318_U109);
  not ginst18289 (P3_ADD_318_U39, P3_PHYADDRPOINTER_REG_19__SCAN_IN);
  not ginst18290 (P3_ADD_318_U4, P3_PHYADDRPOINTER_REG_1__SCAN_IN);
  nand ginst18291 (P3_ADD_318_U40, P3_PHYADDRPOINTER_REG_19__SCAN_IN, P3_ADD_318_U110);
  not ginst18292 (P3_ADD_318_U41, P3_PHYADDRPOINTER_REG_20__SCAN_IN);
  nand ginst18293 (P3_ADD_318_U42, P3_PHYADDRPOINTER_REG_20__SCAN_IN, P3_ADD_318_U111);
  not ginst18294 (P3_ADD_318_U43, P3_PHYADDRPOINTER_REG_21__SCAN_IN);
  nand ginst18295 (P3_ADD_318_U44, P3_PHYADDRPOINTER_REG_21__SCAN_IN, P3_ADD_318_U112);
  not ginst18296 (P3_ADD_318_U45, P3_PHYADDRPOINTER_REG_22__SCAN_IN);
  nand ginst18297 (P3_ADD_318_U46, P3_PHYADDRPOINTER_REG_22__SCAN_IN, P3_ADD_318_U113);
  not ginst18298 (P3_ADD_318_U47, P3_PHYADDRPOINTER_REG_23__SCAN_IN);
  nand ginst18299 (P3_ADD_318_U48, P3_PHYADDRPOINTER_REG_23__SCAN_IN, P3_ADD_318_U114);
  not ginst18300 (P3_ADD_318_U49, P3_PHYADDRPOINTER_REG_24__SCAN_IN);
  not ginst18301 (P3_ADD_318_U5, P3_PHYADDRPOINTER_REG_2__SCAN_IN);
  nand ginst18302 (P3_ADD_318_U50, P3_PHYADDRPOINTER_REG_24__SCAN_IN, P3_ADD_318_U115);
  not ginst18303 (P3_ADD_318_U51, P3_PHYADDRPOINTER_REG_25__SCAN_IN);
  nand ginst18304 (P3_ADD_318_U52, P3_PHYADDRPOINTER_REG_25__SCAN_IN, P3_ADD_318_U116);
  not ginst18305 (P3_ADD_318_U53, P3_PHYADDRPOINTER_REG_26__SCAN_IN);
  nand ginst18306 (P3_ADD_318_U54, P3_PHYADDRPOINTER_REG_26__SCAN_IN, P3_ADD_318_U117);
  not ginst18307 (P3_ADD_318_U55, P3_PHYADDRPOINTER_REG_27__SCAN_IN);
  nand ginst18308 (P3_ADD_318_U56, P3_PHYADDRPOINTER_REG_27__SCAN_IN, P3_ADD_318_U118);
  not ginst18309 (P3_ADD_318_U57, P3_PHYADDRPOINTER_REG_28__SCAN_IN);
  nand ginst18310 (P3_ADD_318_U58, P3_PHYADDRPOINTER_REG_28__SCAN_IN, P3_ADD_318_U119);
  not ginst18311 (P3_ADD_318_U59, P3_PHYADDRPOINTER_REG_29__SCAN_IN);
  nand ginst18312 (P3_ADD_318_U6, P3_PHYADDRPOINTER_REG_1__SCAN_IN, P3_PHYADDRPOINTER_REG_2__SCAN_IN);
  nand ginst18313 (P3_ADD_318_U60, P3_PHYADDRPOINTER_REG_29__SCAN_IN, P3_ADD_318_U120);
  not ginst18314 (P3_ADD_318_U61, P3_PHYADDRPOINTER_REG_30__SCAN_IN);
  nand ginst18315 (P3_ADD_318_U62, P3_ADD_318_U123, P3_ADD_318_U124);
  nand ginst18316 (P3_ADD_318_U63, P3_ADD_318_U125, P3_ADD_318_U126);
  nand ginst18317 (P3_ADD_318_U64, P3_ADD_318_U127, P3_ADD_318_U128);
  nand ginst18318 (P3_ADD_318_U65, P3_ADD_318_U129, P3_ADD_318_U130);
  nand ginst18319 (P3_ADD_318_U66, P3_ADD_318_U131, P3_ADD_318_U132);
  nand ginst18320 (P3_ADD_318_U67, P3_ADD_318_U133, P3_ADD_318_U134);
  nand ginst18321 (P3_ADD_318_U68, P3_ADD_318_U135, P3_ADD_318_U136);
  nand ginst18322 (P3_ADD_318_U69, P3_ADD_318_U137, P3_ADD_318_U138);
  not ginst18323 (P3_ADD_318_U7, P3_PHYADDRPOINTER_REG_3__SCAN_IN);
  nand ginst18324 (P3_ADD_318_U70, P3_ADD_318_U139, P3_ADD_318_U140);
  nand ginst18325 (P3_ADD_318_U71, P3_ADD_318_U141, P3_ADD_318_U142);
  nand ginst18326 (P3_ADD_318_U72, P3_ADD_318_U143, P3_ADD_318_U144);
  nand ginst18327 (P3_ADD_318_U73, P3_ADD_318_U145, P3_ADD_318_U146);
  nand ginst18328 (P3_ADD_318_U74, P3_ADD_318_U147, P3_ADD_318_U148);
  nand ginst18329 (P3_ADD_318_U75, P3_ADD_318_U149, P3_ADD_318_U150);
  nand ginst18330 (P3_ADD_318_U76, P3_ADD_318_U151, P3_ADD_318_U152);
  nand ginst18331 (P3_ADD_318_U77, P3_ADD_318_U153, P3_ADD_318_U154);
  nand ginst18332 (P3_ADD_318_U78, P3_ADD_318_U155, P3_ADD_318_U156);
  nand ginst18333 (P3_ADD_318_U79, P3_ADD_318_U157, P3_ADD_318_U158);
  nand ginst18334 (P3_ADD_318_U8, P3_PHYADDRPOINTER_REG_3__SCAN_IN, P3_ADD_318_U94);
  nand ginst18335 (P3_ADD_318_U80, P3_ADD_318_U159, P3_ADD_318_U160);
  nand ginst18336 (P3_ADD_318_U81, P3_ADD_318_U161, P3_ADD_318_U162);
  nand ginst18337 (P3_ADD_318_U82, P3_ADD_318_U163, P3_ADD_318_U164);
  nand ginst18338 (P3_ADD_318_U83, P3_ADD_318_U165, P3_ADD_318_U166);
  nand ginst18339 (P3_ADD_318_U84, P3_ADD_318_U167, P3_ADD_318_U168);
  nand ginst18340 (P3_ADD_318_U85, P3_ADD_318_U169, P3_ADD_318_U170);
  nand ginst18341 (P3_ADD_318_U86, P3_ADD_318_U171, P3_ADD_318_U172);
  nand ginst18342 (P3_ADD_318_U87, P3_ADD_318_U173, P3_ADD_318_U174);
  nand ginst18343 (P3_ADD_318_U88, P3_ADD_318_U175, P3_ADD_318_U176);
  nand ginst18344 (P3_ADD_318_U89, P3_ADD_318_U177, P3_ADD_318_U178);
  not ginst18345 (P3_ADD_318_U9, P3_PHYADDRPOINTER_REG_4__SCAN_IN);
  nand ginst18346 (P3_ADD_318_U90, P3_ADD_318_U179, P3_ADD_318_U180);
  nand ginst18347 (P3_ADD_318_U91, P3_ADD_318_U181, P3_ADD_318_U182);
  not ginst18348 (P3_ADD_318_U92, P3_PHYADDRPOINTER_REG_31__SCAN_IN);
  nand ginst18349 (P3_ADD_318_U93, P3_PHYADDRPOINTER_REG_30__SCAN_IN, P3_ADD_318_U121);
  not ginst18350 (P3_ADD_318_U94, P3_ADD_318_U6);
  not ginst18351 (P3_ADD_318_U95, P3_ADD_318_U8);
  not ginst18352 (P3_ADD_318_U96, P3_ADD_318_U10);
  not ginst18353 (P3_ADD_318_U97, P3_ADD_318_U12);
  not ginst18354 (P3_ADD_318_U98, P3_ADD_318_U14);
  not ginst18355 (P3_ADD_318_U99, P3_ADD_318_U16);
  nand ginst18356 (P3_ADD_339_U10, P3_PHYADDRPOINTER_REG_4__SCAN_IN, P3_ADD_339_U95);
  not ginst18357 (P3_ADD_339_U100, P3_ADD_339_U19);
  not ginst18358 (P3_ADD_339_U101, P3_ADD_339_U20);
  not ginst18359 (P3_ADD_339_U102, P3_ADD_339_U22);
  not ginst18360 (P3_ADD_339_U103, P3_ADD_339_U24);
  not ginst18361 (P3_ADD_339_U104, P3_ADD_339_U26);
  not ginst18362 (P3_ADD_339_U105, P3_ADD_339_U28);
  not ginst18363 (P3_ADD_339_U106, P3_ADD_339_U30);
  not ginst18364 (P3_ADD_339_U107, P3_ADD_339_U32);
  not ginst18365 (P3_ADD_339_U108, P3_ADD_339_U34);
  not ginst18366 (P3_ADD_339_U109, P3_ADD_339_U36);
  not ginst18367 (P3_ADD_339_U11, P3_PHYADDRPOINTER_REG_5__SCAN_IN);
  not ginst18368 (P3_ADD_339_U110, P3_ADD_339_U38);
  not ginst18369 (P3_ADD_339_U111, P3_ADD_339_U40);
  not ginst18370 (P3_ADD_339_U112, P3_ADD_339_U42);
  not ginst18371 (P3_ADD_339_U113, P3_ADD_339_U44);
  not ginst18372 (P3_ADD_339_U114, P3_ADD_339_U46);
  not ginst18373 (P3_ADD_339_U115, P3_ADD_339_U48);
  not ginst18374 (P3_ADD_339_U116, P3_ADD_339_U50);
  not ginst18375 (P3_ADD_339_U117, P3_ADD_339_U52);
  not ginst18376 (P3_ADD_339_U118, P3_ADD_339_U54);
  not ginst18377 (P3_ADD_339_U119, P3_ADD_339_U56);
  nand ginst18378 (P3_ADD_339_U12, P3_PHYADDRPOINTER_REG_5__SCAN_IN, P3_ADD_339_U96);
  not ginst18379 (P3_ADD_339_U120, P3_ADD_339_U58);
  not ginst18380 (P3_ADD_339_U121, P3_ADD_339_U60);
  not ginst18381 (P3_ADD_339_U122, P3_ADD_339_U93);
  nand ginst18382 (P3_ADD_339_U123, P3_PHYADDRPOINTER_REG_9__SCAN_IN, P3_ADD_339_U19);
  nand ginst18383 (P3_ADD_339_U124, P3_ADD_339_U100, P3_ADD_339_U18);
  nand ginst18384 (P3_ADD_339_U125, P3_PHYADDRPOINTER_REG_8__SCAN_IN, P3_ADD_339_U16);
  nand ginst18385 (P3_ADD_339_U126, P3_ADD_339_U17, P3_ADD_339_U99);
  nand ginst18386 (P3_ADD_339_U127, P3_PHYADDRPOINTER_REG_7__SCAN_IN, P3_ADD_339_U14);
  nand ginst18387 (P3_ADD_339_U128, P3_ADD_339_U15, P3_ADD_339_U98);
  nand ginst18388 (P3_ADD_339_U129, P3_PHYADDRPOINTER_REG_6__SCAN_IN, P3_ADD_339_U12);
  not ginst18389 (P3_ADD_339_U13, P3_PHYADDRPOINTER_REG_6__SCAN_IN);
  nand ginst18390 (P3_ADD_339_U130, P3_ADD_339_U13, P3_ADD_339_U97);
  nand ginst18391 (P3_ADD_339_U131, P3_PHYADDRPOINTER_REG_5__SCAN_IN, P3_ADD_339_U10);
  nand ginst18392 (P3_ADD_339_U132, P3_ADD_339_U11, P3_ADD_339_U96);
  nand ginst18393 (P3_ADD_339_U133, P3_PHYADDRPOINTER_REG_4__SCAN_IN, P3_ADD_339_U8);
  nand ginst18394 (P3_ADD_339_U134, P3_ADD_339_U9, P3_ADD_339_U95);
  nand ginst18395 (P3_ADD_339_U135, P3_PHYADDRPOINTER_REG_3__SCAN_IN, P3_ADD_339_U6);
  nand ginst18396 (P3_ADD_339_U136, P3_ADD_339_U7, P3_ADD_339_U94);
  nand ginst18397 (P3_ADD_339_U137, P3_PHYADDRPOINTER_REG_31__SCAN_IN, P3_ADD_339_U93);
  nand ginst18398 (P3_ADD_339_U138, P3_ADD_339_U122, P3_ADD_339_U92);
  nand ginst18399 (P3_ADD_339_U139, P3_PHYADDRPOINTER_REG_30__SCAN_IN, P3_ADD_339_U60);
  nand ginst18400 (P3_ADD_339_U14, P3_PHYADDRPOINTER_REG_6__SCAN_IN, P3_ADD_339_U97);
  nand ginst18401 (P3_ADD_339_U140, P3_ADD_339_U121, P3_ADD_339_U61);
  nand ginst18402 (P3_ADD_339_U141, P3_PHYADDRPOINTER_REG_2__SCAN_IN, P3_ADD_339_U4);
  nand ginst18403 (P3_ADD_339_U142, P3_PHYADDRPOINTER_REG_1__SCAN_IN, P3_ADD_339_U5);
  nand ginst18404 (P3_ADD_339_U143, P3_PHYADDRPOINTER_REG_29__SCAN_IN, P3_ADD_339_U58);
  nand ginst18405 (P3_ADD_339_U144, P3_ADD_339_U120, P3_ADD_339_U59);
  nand ginst18406 (P3_ADD_339_U145, P3_PHYADDRPOINTER_REG_28__SCAN_IN, P3_ADD_339_U56);
  nand ginst18407 (P3_ADD_339_U146, P3_ADD_339_U119, P3_ADD_339_U57);
  nand ginst18408 (P3_ADD_339_U147, P3_PHYADDRPOINTER_REG_27__SCAN_IN, P3_ADD_339_U54);
  nand ginst18409 (P3_ADD_339_U148, P3_ADD_339_U118, P3_ADD_339_U55);
  nand ginst18410 (P3_ADD_339_U149, P3_PHYADDRPOINTER_REG_26__SCAN_IN, P3_ADD_339_U52);
  not ginst18411 (P3_ADD_339_U15, P3_PHYADDRPOINTER_REG_7__SCAN_IN);
  nand ginst18412 (P3_ADD_339_U150, P3_ADD_339_U117, P3_ADD_339_U53);
  nand ginst18413 (P3_ADD_339_U151, P3_PHYADDRPOINTER_REG_25__SCAN_IN, P3_ADD_339_U50);
  nand ginst18414 (P3_ADD_339_U152, P3_ADD_339_U116, P3_ADD_339_U51);
  nand ginst18415 (P3_ADD_339_U153, P3_PHYADDRPOINTER_REG_24__SCAN_IN, P3_ADD_339_U48);
  nand ginst18416 (P3_ADD_339_U154, P3_ADD_339_U115, P3_ADD_339_U49);
  nand ginst18417 (P3_ADD_339_U155, P3_PHYADDRPOINTER_REG_23__SCAN_IN, P3_ADD_339_U46);
  nand ginst18418 (P3_ADD_339_U156, P3_ADD_339_U114, P3_ADD_339_U47);
  nand ginst18419 (P3_ADD_339_U157, P3_PHYADDRPOINTER_REG_22__SCAN_IN, P3_ADD_339_U44);
  nand ginst18420 (P3_ADD_339_U158, P3_ADD_339_U113, P3_ADD_339_U45);
  nand ginst18421 (P3_ADD_339_U159, P3_PHYADDRPOINTER_REG_21__SCAN_IN, P3_ADD_339_U42);
  nand ginst18422 (P3_ADD_339_U16, P3_PHYADDRPOINTER_REG_7__SCAN_IN, P3_ADD_339_U98);
  nand ginst18423 (P3_ADD_339_U160, P3_ADD_339_U112, P3_ADD_339_U43);
  nand ginst18424 (P3_ADD_339_U161, P3_PHYADDRPOINTER_REG_20__SCAN_IN, P3_ADD_339_U40);
  nand ginst18425 (P3_ADD_339_U162, P3_ADD_339_U111, P3_ADD_339_U41);
  nand ginst18426 (P3_ADD_339_U163, P3_PHYADDRPOINTER_REG_19__SCAN_IN, P3_ADD_339_U38);
  nand ginst18427 (P3_ADD_339_U164, P3_ADD_339_U110, P3_ADD_339_U39);
  nand ginst18428 (P3_ADD_339_U165, P3_PHYADDRPOINTER_REG_18__SCAN_IN, P3_ADD_339_U36);
  nand ginst18429 (P3_ADD_339_U166, P3_ADD_339_U109, P3_ADD_339_U37);
  nand ginst18430 (P3_ADD_339_U167, P3_PHYADDRPOINTER_REG_17__SCAN_IN, P3_ADD_339_U34);
  nand ginst18431 (P3_ADD_339_U168, P3_ADD_339_U108, P3_ADD_339_U35);
  nand ginst18432 (P3_ADD_339_U169, P3_PHYADDRPOINTER_REG_16__SCAN_IN, P3_ADD_339_U32);
  not ginst18433 (P3_ADD_339_U17, P3_PHYADDRPOINTER_REG_8__SCAN_IN);
  nand ginst18434 (P3_ADD_339_U170, P3_ADD_339_U107, P3_ADD_339_U33);
  nand ginst18435 (P3_ADD_339_U171, P3_PHYADDRPOINTER_REG_15__SCAN_IN, P3_ADD_339_U30);
  nand ginst18436 (P3_ADD_339_U172, P3_ADD_339_U106, P3_ADD_339_U31);
  nand ginst18437 (P3_ADD_339_U173, P3_PHYADDRPOINTER_REG_14__SCAN_IN, P3_ADD_339_U28);
  nand ginst18438 (P3_ADD_339_U174, P3_ADD_339_U105, P3_ADD_339_U29);
  nand ginst18439 (P3_ADD_339_U175, P3_PHYADDRPOINTER_REG_13__SCAN_IN, P3_ADD_339_U26);
  nand ginst18440 (P3_ADD_339_U176, P3_ADD_339_U104, P3_ADD_339_U27);
  nand ginst18441 (P3_ADD_339_U177, P3_PHYADDRPOINTER_REG_12__SCAN_IN, P3_ADD_339_U24);
  nand ginst18442 (P3_ADD_339_U178, P3_ADD_339_U103, P3_ADD_339_U25);
  nand ginst18443 (P3_ADD_339_U179, P3_PHYADDRPOINTER_REG_11__SCAN_IN, P3_ADD_339_U22);
  not ginst18444 (P3_ADD_339_U18, P3_PHYADDRPOINTER_REG_9__SCAN_IN);
  nand ginst18445 (P3_ADD_339_U180, P3_ADD_339_U102, P3_ADD_339_U23);
  nand ginst18446 (P3_ADD_339_U181, P3_PHYADDRPOINTER_REG_10__SCAN_IN, P3_ADD_339_U20);
  nand ginst18447 (P3_ADD_339_U182, P3_ADD_339_U101, P3_ADD_339_U21);
  nand ginst18448 (P3_ADD_339_U19, P3_PHYADDRPOINTER_REG_8__SCAN_IN, P3_ADD_339_U99);
  nand ginst18449 (P3_ADD_339_U20, P3_PHYADDRPOINTER_REG_9__SCAN_IN, P3_ADD_339_U100);
  not ginst18450 (P3_ADD_339_U21, P3_PHYADDRPOINTER_REG_10__SCAN_IN);
  nand ginst18451 (P3_ADD_339_U22, P3_PHYADDRPOINTER_REG_10__SCAN_IN, P3_ADD_339_U101);
  not ginst18452 (P3_ADD_339_U23, P3_PHYADDRPOINTER_REG_11__SCAN_IN);
  nand ginst18453 (P3_ADD_339_U24, P3_PHYADDRPOINTER_REG_11__SCAN_IN, P3_ADD_339_U102);
  not ginst18454 (P3_ADD_339_U25, P3_PHYADDRPOINTER_REG_12__SCAN_IN);
  nand ginst18455 (P3_ADD_339_U26, P3_PHYADDRPOINTER_REG_12__SCAN_IN, P3_ADD_339_U103);
  not ginst18456 (P3_ADD_339_U27, P3_PHYADDRPOINTER_REG_13__SCAN_IN);
  nand ginst18457 (P3_ADD_339_U28, P3_PHYADDRPOINTER_REG_13__SCAN_IN, P3_ADD_339_U104);
  not ginst18458 (P3_ADD_339_U29, P3_PHYADDRPOINTER_REG_14__SCAN_IN);
  nand ginst18459 (P3_ADD_339_U30, P3_PHYADDRPOINTER_REG_14__SCAN_IN, P3_ADD_339_U105);
  not ginst18460 (P3_ADD_339_U31, P3_PHYADDRPOINTER_REG_15__SCAN_IN);
  nand ginst18461 (P3_ADD_339_U32, P3_PHYADDRPOINTER_REG_15__SCAN_IN, P3_ADD_339_U106);
  not ginst18462 (P3_ADD_339_U33, P3_PHYADDRPOINTER_REG_16__SCAN_IN);
  nand ginst18463 (P3_ADD_339_U34, P3_PHYADDRPOINTER_REG_16__SCAN_IN, P3_ADD_339_U107);
  not ginst18464 (P3_ADD_339_U35, P3_PHYADDRPOINTER_REG_17__SCAN_IN);
  nand ginst18465 (P3_ADD_339_U36, P3_PHYADDRPOINTER_REG_17__SCAN_IN, P3_ADD_339_U108);
  not ginst18466 (P3_ADD_339_U37, P3_PHYADDRPOINTER_REG_18__SCAN_IN);
  nand ginst18467 (P3_ADD_339_U38, P3_PHYADDRPOINTER_REG_18__SCAN_IN, P3_ADD_339_U109);
  not ginst18468 (P3_ADD_339_U39, P3_PHYADDRPOINTER_REG_19__SCAN_IN);
  not ginst18469 (P3_ADD_339_U4, P3_PHYADDRPOINTER_REG_1__SCAN_IN);
  nand ginst18470 (P3_ADD_339_U40, P3_PHYADDRPOINTER_REG_19__SCAN_IN, P3_ADD_339_U110);
  not ginst18471 (P3_ADD_339_U41, P3_PHYADDRPOINTER_REG_20__SCAN_IN);
  nand ginst18472 (P3_ADD_339_U42, P3_PHYADDRPOINTER_REG_20__SCAN_IN, P3_ADD_339_U111);
  not ginst18473 (P3_ADD_339_U43, P3_PHYADDRPOINTER_REG_21__SCAN_IN);
  nand ginst18474 (P3_ADD_339_U44, P3_PHYADDRPOINTER_REG_21__SCAN_IN, P3_ADD_339_U112);
  not ginst18475 (P3_ADD_339_U45, P3_PHYADDRPOINTER_REG_22__SCAN_IN);
  nand ginst18476 (P3_ADD_339_U46, P3_PHYADDRPOINTER_REG_22__SCAN_IN, P3_ADD_339_U113);
  not ginst18477 (P3_ADD_339_U47, P3_PHYADDRPOINTER_REG_23__SCAN_IN);
  nand ginst18478 (P3_ADD_339_U48, P3_PHYADDRPOINTER_REG_23__SCAN_IN, P3_ADD_339_U114);
  not ginst18479 (P3_ADD_339_U49, P3_PHYADDRPOINTER_REG_24__SCAN_IN);
  not ginst18480 (P3_ADD_339_U5, P3_PHYADDRPOINTER_REG_2__SCAN_IN);
  nand ginst18481 (P3_ADD_339_U50, P3_PHYADDRPOINTER_REG_24__SCAN_IN, P3_ADD_339_U115);
  not ginst18482 (P3_ADD_339_U51, P3_PHYADDRPOINTER_REG_25__SCAN_IN);
  nand ginst18483 (P3_ADD_339_U52, P3_PHYADDRPOINTER_REG_25__SCAN_IN, P3_ADD_339_U116);
  not ginst18484 (P3_ADD_339_U53, P3_PHYADDRPOINTER_REG_26__SCAN_IN);
  nand ginst18485 (P3_ADD_339_U54, P3_PHYADDRPOINTER_REG_26__SCAN_IN, P3_ADD_339_U117);
  not ginst18486 (P3_ADD_339_U55, P3_PHYADDRPOINTER_REG_27__SCAN_IN);
  nand ginst18487 (P3_ADD_339_U56, P3_PHYADDRPOINTER_REG_27__SCAN_IN, P3_ADD_339_U118);
  not ginst18488 (P3_ADD_339_U57, P3_PHYADDRPOINTER_REG_28__SCAN_IN);
  nand ginst18489 (P3_ADD_339_U58, P3_PHYADDRPOINTER_REG_28__SCAN_IN, P3_ADD_339_U119);
  not ginst18490 (P3_ADD_339_U59, P3_PHYADDRPOINTER_REG_29__SCAN_IN);
  nand ginst18491 (P3_ADD_339_U6, P3_PHYADDRPOINTER_REG_1__SCAN_IN, P3_PHYADDRPOINTER_REG_2__SCAN_IN);
  nand ginst18492 (P3_ADD_339_U60, P3_PHYADDRPOINTER_REG_29__SCAN_IN, P3_ADD_339_U120);
  not ginst18493 (P3_ADD_339_U61, P3_PHYADDRPOINTER_REG_30__SCAN_IN);
  nand ginst18494 (P3_ADD_339_U62, P3_ADD_339_U123, P3_ADD_339_U124);
  nand ginst18495 (P3_ADD_339_U63, P3_ADD_339_U125, P3_ADD_339_U126);
  nand ginst18496 (P3_ADD_339_U64, P3_ADD_339_U127, P3_ADD_339_U128);
  nand ginst18497 (P3_ADD_339_U65, P3_ADD_339_U129, P3_ADD_339_U130);
  nand ginst18498 (P3_ADD_339_U66, P3_ADD_339_U131, P3_ADD_339_U132);
  nand ginst18499 (P3_ADD_339_U67, P3_ADD_339_U133, P3_ADD_339_U134);
  nand ginst18500 (P3_ADD_339_U68, P3_ADD_339_U135, P3_ADD_339_U136);
  nand ginst18501 (P3_ADD_339_U69, P3_ADD_339_U137, P3_ADD_339_U138);
  not ginst18502 (P3_ADD_339_U7, P3_PHYADDRPOINTER_REG_3__SCAN_IN);
  nand ginst18503 (P3_ADD_339_U70, P3_ADD_339_U139, P3_ADD_339_U140);
  nand ginst18504 (P3_ADD_339_U71, P3_ADD_339_U141, P3_ADD_339_U142);
  nand ginst18505 (P3_ADD_339_U72, P3_ADD_339_U143, P3_ADD_339_U144);
  nand ginst18506 (P3_ADD_339_U73, P3_ADD_339_U145, P3_ADD_339_U146);
  nand ginst18507 (P3_ADD_339_U74, P3_ADD_339_U147, P3_ADD_339_U148);
  nand ginst18508 (P3_ADD_339_U75, P3_ADD_339_U149, P3_ADD_339_U150);
  nand ginst18509 (P3_ADD_339_U76, P3_ADD_339_U151, P3_ADD_339_U152);
  nand ginst18510 (P3_ADD_339_U77, P3_ADD_339_U153, P3_ADD_339_U154);
  nand ginst18511 (P3_ADD_339_U78, P3_ADD_339_U155, P3_ADD_339_U156);
  nand ginst18512 (P3_ADD_339_U79, P3_ADD_339_U157, P3_ADD_339_U158);
  nand ginst18513 (P3_ADD_339_U8, P3_PHYADDRPOINTER_REG_3__SCAN_IN, P3_ADD_339_U94);
  nand ginst18514 (P3_ADD_339_U80, P3_ADD_339_U159, P3_ADD_339_U160);
  nand ginst18515 (P3_ADD_339_U81, P3_ADD_339_U161, P3_ADD_339_U162);
  nand ginst18516 (P3_ADD_339_U82, P3_ADD_339_U163, P3_ADD_339_U164);
  nand ginst18517 (P3_ADD_339_U83, P3_ADD_339_U165, P3_ADD_339_U166);
  nand ginst18518 (P3_ADD_339_U84, P3_ADD_339_U167, P3_ADD_339_U168);
  nand ginst18519 (P3_ADD_339_U85, P3_ADD_339_U169, P3_ADD_339_U170);
  nand ginst18520 (P3_ADD_339_U86, P3_ADD_339_U171, P3_ADD_339_U172);
  nand ginst18521 (P3_ADD_339_U87, P3_ADD_339_U173, P3_ADD_339_U174);
  nand ginst18522 (P3_ADD_339_U88, P3_ADD_339_U175, P3_ADD_339_U176);
  nand ginst18523 (P3_ADD_339_U89, P3_ADD_339_U177, P3_ADD_339_U178);
  not ginst18524 (P3_ADD_339_U9, P3_PHYADDRPOINTER_REG_4__SCAN_IN);
  nand ginst18525 (P3_ADD_339_U90, P3_ADD_339_U179, P3_ADD_339_U180);
  nand ginst18526 (P3_ADD_339_U91, P3_ADD_339_U181, P3_ADD_339_U182);
  not ginst18527 (P3_ADD_339_U92, P3_PHYADDRPOINTER_REG_31__SCAN_IN);
  nand ginst18528 (P3_ADD_339_U93, P3_PHYADDRPOINTER_REG_30__SCAN_IN, P3_ADD_339_U121);
  not ginst18529 (P3_ADD_339_U94, P3_ADD_339_U6);
  not ginst18530 (P3_ADD_339_U95, P3_ADD_339_U8);
  not ginst18531 (P3_ADD_339_U96, P3_ADD_339_U10);
  not ginst18532 (P3_ADD_339_U97, P3_ADD_339_U12);
  not ginst18533 (P3_ADD_339_U98, P3_ADD_339_U14);
  not ginst18534 (P3_ADD_339_U99, P3_ADD_339_U16);
  not ginst18535 (P3_ADD_344_U10, P3_INSTADDRPOINTER_REG_3__SCAN_IN);
  not ginst18536 (P3_ADD_344_U100, P3_ADD_344_U11);
  not ginst18537 (P3_ADD_344_U101, P3_ADD_344_U13);
  not ginst18538 (P3_ADD_344_U102, P3_ADD_344_U15);
  not ginst18539 (P3_ADD_344_U103, P3_ADD_344_U17);
  not ginst18540 (P3_ADD_344_U104, P3_ADD_344_U19);
  not ginst18541 (P3_ADD_344_U105, P3_ADD_344_U22);
  not ginst18542 (P3_ADD_344_U106, P3_ADD_344_U23);
  not ginst18543 (P3_ADD_344_U107, P3_ADD_344_U25);
  not ginst18544 (P3_ADD_344_U108, P3_ADD_344_U27);
  not ginst18545 (P3_ADD_344_U109, P3_ADD_344_U29);
  nand ginst18546 (P3_ADD_344_U11, P3_INSTADDRPOINTER_REG_3__SCAN_IN, P3_ADD_344_U99);
  not ginst18547 (P3_ADD_344_U110, P3_ADD_344_U31);
  not ginst18548 (P3_ADD_344_U111, P3_ADD_344_U33);
  not ginst18549 (P3_ADD_344_U112, P3_ADD_344_U35);
  not ginst18550 (P3_ADD_344_U113, P3_ADD_344_U37);
  not ginst18551 (P3_ADD_344_U114, P3_ADD_344_U39);
  not ginst18552 (P3_ADD_344_U115, P3_ADD_344_U41);
  not ginst18553 (P3_ADD_344_U116, P3_ADD_344_U43);
  not ginst18554 (P3_ADD_344_U117, P3_ADD_344_U45);
  not ginst18555 (P3_ADD_344_U118, P3_ADD_344_U47);
  not ginst18556 (P3_ADD_344_U119, P3_ADD_344_U49);
  not ginst18557 (P3_ADD_344_U12, P3_INSTADDRPOINTER_REG_4__SCAN_IN);
  not ginst18558 (P3_ADD_344_U120, P3_ADD_344_U51);
  not ginst18559 (P3_ADD_344_U121, P3_ADD_344_U53);
  not ginst18560 (P3_ADD_344_U122, P3_ADD_344_U55);
  not ginst18561 (P3_ADD_344_U123, P3_ADD_344_U57);
  not ginst18562 (P3_ADD_344_U124, P3_ADD_344_U59);
  not ginst18563 (P3_ADD_344_U125, P3_ADD_344_U61);
  not ginst18564 (P3_ADD_344_U126, P3_ADD_344_U63);
  not ginst18565 (P3_ADD_344_U127, P3_ADD_344_U97);
  nand ginst18566 (P3_ADD_344_U128, P3_INSTADDRPOINTER_REG_9__SCAN_IN, P3_ADD_344_U22);
  nand ginst18567 (P3_ADD_344_U129, P3_ADD_344_U105, P3_ADD_344_U21);
  nand ginst18568 (P3_ADD_344_U13, P3_INSTADDRPOINTER_REG_4__SCAN_IN, P3_ADD_344_U100);
  nand ginst18569 (P3_ADD_344_U130, P3_INSTADDRPOINTER_REG_8__SCAN_IN, P3_ADD_344_U19);
  nand ginst18570 (P3_ADD_344_U131, P3_ADD_344_U104, P3_ADD_344_U20);
  nand ginst18571 (P3_ADD_344_U132, P3_INSTADDRPOINTER_REG_7__SCAN_IN, P3_ADD_344_U17);
  nand ginst18572 (P3_ADD_344_U133, P3_ADD_344_U103, P3_ADD_344_U18);
  nand ginst18573 (P3_ADD_344_U134, P3_INSTADDRPOINTER_REG_6__SCAN_IN, P3_ADD_344_U15);
  nand ginst18574 (P3_ADD_344_U135, P3_ADD_344_U102, P3_ADD_344_U16);
  nand ginst18575 (P3_ADD_344_U136, P3_INSTADDRPOINTER_REG_5__SCAN_IN, P3_ADD_344_U13);
  nand ginst18576 (P3_ADD_344_U137, P3_ADD_344_U101, P3_ADD_344_U14);
  nand ginst18577 (P3_ADD_344_U138, P3_INSTADDRPOINTER_REG_4__SCAN_IN, P3_ADD_344_U11);
  nand ginst18578 (P3_ADD_344_U139, P3_ADD_344_U100, P3_ADD_344_U12);
  not ginst18579 (P3_ADD_344_U14, P3_INSTADDRPOINTER_REG_5__SCAN_IN);
  nand ginst18580 (P3_ADD_344_U140, P3_INSTADDRPOINTER_REG_3__SCAN_IN, P3_ADD_344_U9);
  nand ginst18581 (P3_ADD_344_U141, P3_ADD_344_U10, P3_ADD_344_U99);
  nand ginst18582 (P3_ADD_344_U142, P3_INSTADDRPOINTER_REG_31__SCAN_IN, P3_ADD_344_U97);
  nand ginst18583 (P3_ADD_344_U143, P3_ADD_344_U127, P3_ADD_344_U96);
  nand ginst18584 (P3_ADD_344_U144, P3_INSTADDRPOINTER_REG_30__SCAN_IN, P3_ADD_344_U63);
  nand ginst18585 (P3_ADD_344_U145, P3_ADD_344_U126, P3_ADD_344_U64);
  nand ginst18586 (P3_ADD_344_U146, P3_INSTADDRPOINTER_REG_2__SCAN_IN, P3_ADD_344_U7);
  nand ginst18587 (P3_ADD_344_U147, P3_ADD_344_U8, P3_ADD_344_U98);
  nand ginst18588 (P3_ADD_344_U148, P3_INSTADDRPOINTER_REG_29__SCAN_IN, P3_ADD_344_U61);
  nand ginst18589 (P3_ADD_344_U149, P3_ADD_344_U125, P3_ADD_344_U62);
  nand ginst18590 (P3_ADD_344_U15, P3_INSTADDRPOINTER_REG_5__SCAN_IN, P3_ADD_344_U101);
  nand ginst18591 (P3_ADD_344_U150, P3_INSTADDRPOINTER_REG_28__SCAN_IN, P3_ADD_344_U59);
  nand ginst18592 (P3_ADD_344_U151, P3_ADD_344_U124, P3_ADD_344_U60);
  nand ginst18593 (P3_ADD_344_U152, P3_INSTADDRPOINTER_REG_27__SCAN_IN, P3_ADD_344_U57);
  nand ginst18594 (P3_ADD_344_U153, P3_ADD_344_U123, P3_ADD_344_U58);
  nand ginst18595 (P3_ADD_344_U154, P3_INSTADDRPOINTER_REG_26__SCAN_IN, P3_ADD_344_U55);
  nand ginst18596 (P3_ADD_344_U155, P3_ADD_344_U122, P3_ADD_344_U56);
  nand ginst18597 (P3_ADD_344_U156, P3_INSTADDRPOINTER_REG_25__SCAN_IN, P3_ADD_344_U53);
  nand ginst18598 (P3_ADD_344_U157, P3_ADD_344_U121, P3_ADD_344_U54);
  nand ginst18599 (P3_ADD_344_U158, P3_INSTADDRPOINTER_REG_24__SCAN_IN, P3_ADD_344_U51);
  nand ginst18600 (P3_ADD_344_U159, P3_ADD_344_U120, P3_ADD_344_U52);
  not ginst18601 (P3_ADD_344_U16, P3_INSTADDRPOINTER_REG_6__SCAN_IN);
  nand ginst18602 (P3_ADD_344_U160, P3_INSTADDRPOINTER_REG_23__SCAN_IN, P3_ADD_344_U49);
  nand ginst18603 (P3_ADD_344_U161, P3_ADD_344_U119, P3_ADD_344_U50);
  nand ginst18604 (P3_ADD_344_U162, P3_INSTADDRPOINTER_REG_22__SCAN_IN, P3_ADD_344_U47);
  nand ginst18605 (P3_ADD_344_U163, P3_ADD_344_U118, P3_ADD_344_U48);
  nand ginst18606 (P3_ADD_344_U164, P3_INSTADDRPOINTER_REG_21__SCAN_IN, P3_ADD_344_U45);
  nand ginst18607 (P3_ADD_344_U165, P3_ADD_344_U117, P3_ADD_344_U46);
  nand ginst18608 (P3_ADD_344_U166, P3_INSTADDRPOINTER_REG_20__SCAN_IN, P3_ADD_344_U43);
  nand ginst18609 (P3_ADD_344_U167, P3_ADD_344_U116, P3_ADD_344_U44);
  nand ginst18610 (P3_ADD_344_U168, P3_INSTADDRPOINTER_REG_1__SCAN_IN, P3_ADD_344_U5);
  nand ginst18611 (P3_ADD_344_U169, P3_INSTADDRPOINTER_REG_0__SCAN_IN, P3_ADD_344_U6);
  nand ginst18612 (P3_ADD_344_U17, P3_INSTADDRPOINTER_REG_6__SCAN_IN, P3_ADD_344_U102);
  nand ginst18613 (P3_ADD_344_U170, P3_INSTADDRPOINTER_REG_19__SCAN_IN, P3_ADD_344_U41);
  nand ginst18614 (P3_ADD_344_U171, P3_ADD_344_U115, P3_ADD_344_U42);
  nand ginst18615 (P3_ADD_344_U172, P3_INSTADDRPOINTER_REG_18__SCAN_IN, P3_ADD_344_U39);
  nand ginst18616 (P3_ADD_344_U173, P3_ADD_344_U114, P3_ADD_344_U40);
  nand ginst18617 (P3_ADD_344_U174, P3_INSTADDRPOINTER_REG_17__SCAN_IN, P3_ADD_344_U37);
  nand ginst18618 (P3_ADD_344_U175, P3_ADD_344_U113, P3_ADD_344_U38);
  nand ginst18619 (P3_ADD_344_U176, P3_INSTADDRPOINTER_REG_16__SCAN_IN, P3_ADD_344_U35);
  nand ginst18620 (P3_ADD_344_U177, P3_ADD_344_U112, P3_ADD_344_U36);
  nand ginst18621 (P3_ADD_344_U178, P3_INSTADDRPOINTER_REG_15__SCAN_IN, P3_ADD_344_U33);
  nand ginst18622 (P3_ADD_344_U179, P3_ADD_344_U111, P3_ADD_344_U34);
  not ginst18623 (P3_ADD_344_U18, P3_INSTADDRPOINTER_REG_7__SCAN_IN);
  nand ginst18624 (P3_ADD_344_U180, P3_INSTADDRPOINTER_REG_14__SCAN_IN, P3_ADD_344_U31);
  nand ginst18625 (P3_ADD_344_U181, P3_ADD_344_U110, P3_ADD_344_U32);
  nand ginst18626 (P3_ADD_344_U182, P3_INSTADDRPOINTER_REG_13__SCAN_IN, P3_ADD_344_U29);
  nand ginst18627 (P3_ADD_344_U183, P3_ADD_344_U109, P3_ADD_344_U30);
  nand ginst18628 (P3_ADD_344_U184, P3_INSTADDRPOINTER_REG_12__SCAN_IN, P3_ADD_344_U27);
  nand ginst18629 (P3_ADD_344_U185, P3_ADD_344_U108, P3_ADD_344_U28);
  nand ginst18630 (P3_ADD_344_U186, P3_INSTADDRPOINTER_REG_11__SCAN_IN, P3_ADD_344_U25);
  nand ginst18631 (P3_ADD_344_U187, P3_ADD_344_U107, P3_ADD_344_U26);
  nand ginst18632 (P3_ADD_344_U188, P3_INSTADDRPOINTER_REG_10__SCAN_IN, P3_ADD_344_U23);
  nand ginst18633 (P3_ADD_344_U189, P3_ADD_344_U106, P3_ADD_344_U24);
  nand ginst18634 (P3_ADD_344_U19, P3_INSTADDRPOINTER_REG_7__SCAN_IN, P3_ADD_344_U103);
  not ginst18635 (P3_ADD_344_U20, P3_INSTADDRPOINTER_REG_8__SCAN_IN);
  not ginst18636 (P3_ADD_344_U21, P3_INSTADDRPOINTER_REG_9__SCAN_IN);
  nand ginst18637 (P3_ADD_344_U22, P3_INSTADDRPOINTER_REG_8__SCAN_IN, P3_ADD_344_U104);
  nand ginst18638 (P3_ADD_344_U23, P3_INSTADDRPOINTER_REG_9__SCAN_IN, P3_ADD_344_U105);
  not ginst18639 (P3_ADD_344_U24, P3_INSTADDRPOINTER_REG_10__SCAN_IN);
  nand ginst18640 (P3_ADD_344_U25, P3_INSTADDRPOINTER_REG_10__SCAN_IN, P3_ADD_344_U106);
  not ginst18641 (P3_ADD_344_U26, P3_INSTADDRPOINTER_REG_11__SCAN_IN);
  nand ginst18642 (P3_ADD_344_U27, P3_INSTADDRPOINTER_REG_11__SCAN_IN, P3_ADD_344_U107);
  not ginst18643 (P3_ADD_344_U28, P3_INSTADDRPOINTER_REG_12__SCAN_IN);
  nand ginst18644 (P3_ADD_344_U29, P3_INSTADDRPOINTER_REG_12__SCAN_IN, P3_ADD_344_U108);
  not ginst18645 (P3_ADD_344_U30, P3_INSTADDRPOINTER_REG_13__SCAN_IN);
  nand ginst18646 (P3_ADD_344_U31, P3_INSTADDRPOINTER_REG_13__SCAN_IN, P3_ADD_344_U109);
  not ginst18647 (P3_ADD_344_U32, P3_INSTADDRPOINTER_REG_14__SCAN_IN);
  nand ginst18648 (P3_ADD_344_U33, P3_INSTADDRPOINTER_REG_14__SCAN_IN, P3_ADD_344_U110);
  not ginst18649 (P3_ADD_344_U34, P3_INSTADDRPOINTER_REG_15__SCAN_IN);
  nand ginst18650 (P3_ADD_344_U35, P3_INSTADDRPOINTER_REG_15__SCAN_IN, P3_ADD_344_U111);
  not ginst18651 (P3_ADD_344_U36, P3_INSTADDRPOINTER_REG_16__SCAN_IN);
  nand ginst18652 (P3_ADD_344_U37, P3_INSTADDRPOINTER_REG_16__SCAN_IN, P3_ADD_344_U112);
  not ginst18653 (P3_ADD_344_U38, P3_INSTADDRPOINTER_REG_17__SCAN_IN);
  nand ginst18654 (P3_ADD_344_U39, P3_INSTADDRPOINTER_REG_17__SCAN_IN, P3_ADD_344_U113);
  not ginst18655 (P3_ADD_344_U40, P3_INSTADDRPOINTER_REG_18__SCAN_IN);
  nand ginst18656 (P3_ADD_344_U41, P3_INSTADDRPOINTER_REG_18__SCAN_IN, P3_ADD_344_U114);
  not ginst18657 (P3_ADD_344_U42, P3_INSTADDRPOINTER_REG_19__SCAN_IN);
  nand ginst18658 (P3_ADD_344_U43, P3_INSTADDRPOINTER_REG_19__SCAN_IN, P3_ADD_344_U115);
  not ginst18659 (P3_ADD_344_U44, P3_INSTADDRPOINTER_REG_20__SCAN_IN);
  nand ginst18660 (P3_ADD_344_U45, P3_INSTADDRPOINTER_REG_20__SCAN_IN, P3_ADD_344_U116);
  not ginst18661 (P3_ADD_344_U46, P3_INSTADDRPOINTER_REG_21__SCAN_IN);
  nand ginst18662 (P3_ADD_344_U47, P3_INSTADDRPOINTER_REG_21__SCAN_IN, P3_ADD_344_U117);
  not ginst18663 (P3_ADD_344_U48, P3_INSTADDRPOINTER_REG_22__SCAN_IN);
  nand ginst18664 (P3_ADD_344_U49, P3_INSTADDRPOINTER_REG_22__SCAN_IN, P3_ADD_344_U118);
  not ginst18665 (P3_ADD_344_U5, P3_INSTADDRPOINTER_REG_0__SCAN_IN);
  not ginst18666 (P3_ADD_344_U50, P3_INSTADDRPOINTER_REG_23__SCAN_IN);
  nand ginst18667 (P3_ADD_344_U51, P3_INSTADDRPOINTER_REG_23__SCAN_IN, P3_ADD_344_U119);
  not ginst18668 (P3_ADD_344_U52, P3_INSTADDRPOINTER_REG_24__SCAN_IN);
  nand ginst18669 (P3_ADD_344_U53, P3_INSTADDRPOINTER_REG_24__SCAN_IN, P3_ADD_344_U120);
  not ginst18670 (P3_ADD_344_U54, P3_INSTADDRPOINTER_REG_25__SCAN_IN);
  nand ginst18671 (P3_ADD_344_U55, P3_INSTADDRPOINTER_REG_25__SCAN_IN, P3_ADD_344_U121);
  not ginst18672 (P3_ADD_344_U56, P3_INSTADDRPOINTER_REG_26__SCAN_IN);
  nand ginst18673 (P3_ADD_344_U57, P3_INSTADDRPOINTER_REG_26__SCAN_IN, P3_ADD_344_U122);
  not ginst18674 (P3_ADD_344_U58, P3_INSTADDRPOINTER_REG_27__SCAN_IN);
  nand ginst18675 (P3_ADD_344_U59, P3_INSTADDRPOINTER_REG_27__SCAN_IN, P3_ADD_344_U123);
  not ginst18676 (P3_ADD_344_U6, P3_INSTADDRPOINTER_REG_1__SCAN_IN);
  not ginst18677 (P3_ADD_344_U60, P3_INSTADDRPOINTER_REG_28__SCAN_IN);
  nand ginst18678 (P3_ADD_344_U61, P3_INSTADDRPOINTER_REG_28__SCAN_IN, P3_ADD_344_U124);
  not ginst18679 (P3_ADD_344_U62, P3_INSTADDRPOINTER_REG_29__SCAN_IN);
  nand ginst18680 (P3_ADD_344_U63, P3_INSTADDRPOINTER_REG_29__SCAN_IN, P3_ADD_344_U125);
  not ginst18681 (P3_ADD_344_U64, P3_INSTADDRPOINTER_REG_30__SCAN_IN);
  nand ginst18682 (P3_ADD_344_U65, P3_ADD_344_U128, P3_ADD_344_U129);
  nand ginst18683 (P3_ADD_344_U66, P3_ADD_344_U130, P3_ADD_344_U131);
  nand ginst18684 (P3_ADD_344_U67, P3_ADD_344_U132, P3_ADD_344_U133);
  nand ginst18685 (P3_ADD_344_U68, P3_ADD_344_U134, P3_ADD_344_U135);
  nand ginst18686 (P3_ADD_344_U69, P3_ADD_344_U136, P3_ADD_344_U137);
  nand ginst18687 (P3_ADD_344_U7, P3_INSTADDRPOINTER_REG_0__SCAN_IN, P3_INSTADDRPOINTER_REG_1__SCAN_IN);
  nand ginst18688 (P3_ADD_344_U70, P3_ADD_344_U138, P3_ADD_344_U139);
  nand ginst18689 (P3_ADD_344_U71, P3_ADD_344_U140, P3_ADD_344_U141);
  nand ginst18690 (P3_ADD_344_U72, P3_ADD_344_U142, P3_ADD_344_U143);
  nand ginst18691 (P3_ADD_344_U73, P3_ADD_344_U144, P3_ADD_344_U145);
  nand ginst18692 (P3_ADD_344_U74, P3_ADD_344_U146, P3_ADD_344_U147);
  nand ginst18693 (P3_ADD_344_U75, P3_ADD_344_U148, P3_ADD_344_U149);
  nand ginst18694 (P3_ADD_344_U76, P3_ADD_344_U150, P3_ADD_344_U151);
  nand ginst18695 (P3_ADD_344_U77, P3_ADD_344_U152, P3_ADD_344_U153);
  nand ginst18696 (P3_ADD_344_U78, P3_ADD_344_U154, P3_ADD_344_U155);
  nand ginst18697 (P3_ADD_344_U79, P3_ADD_344_U156, P3_ADD_344_U157);
  not ginst18698 (P3_ADD_344_U8, P3_INSTADDRPOINTER_REG_2__SCAN_IN);
  nand ginst18699 (P3_ADD_344_U80, P3_ADD_344_U158, P3_ADD_344_U159);
  nand ginst18700 (P3_ADD_344_U81, P3_ADD_344_U160, P3_ADD_344_U161);
  nand ginst18701 (P3_ADD_344_U82, P3_ADD_344_U162, P3_ADD_344_U163);
  nand ginst18702 (P3_ADD_344_U83, P3_ADD_344_U164, P3_ADD_344_U165);
  nand ginst18703 (P3_ADD_344_U84, P3_ADD_344_U166, P3_ADD_344_U167);
  nand ginst18704 (P3_ADD_344_U85, P3_ADD_344_U168, P3_ADD_344_U169);
  nand ginst18705 (P3_ADD_344_U86, P3_ADD_344_U170, P3_ADD_344_U171);
  nand ginst18706 (P3_ADD_344_U87, P3_ADD_344_U172, P3_ADD_344_U173);
  nand ginst18707 (P3_ADD_344_U88, P3_ADD_344_U174, P3_ADD_344_U175);
  nand ginst18708 (P3_ADD_344_U89, P3_ADD_344_U176, P3_ADD_344_U177);
  nand ginst18709 (P3_ADD_344_U9, P3_INSTADDRPOINTER_REG_2__SCAN_IN, P3_ADD_344_U98);
  nand ginst18710 (P3_ADD_344_U90, P3_ADD_344_U178, P3_ADD_344_U179);
  nand ginst18711 (P3_ADD_344_U91, P3_ADD_344_U180, P3_ADD_344_U181);
  nand ginst18712 (P3_ADD_344_U92, P3_ADD_344_U182, P3_ADD_344_U183);
  nand ginst18713 (P3_ADD_344_U93, P3_ADD_344_U184, P3_ADD_344_U185);
  nand ginst18714 (P3_ADD_344_U94, P3_ADD_344_U186, P3_ADD_344_U187);
  nand ginst18715 (P3_ADD_344_U95, P3_ADD_344_U188, P3_ADD_344_U189);
  not ginst18716 (P3_ADD_344_U96, P3_INSTADDRPOINTER_REG_31__SCAN_IN);
  nand ginst18717 (P3_ADD_344_U97, P3_INSTADDRPOINTER_REG_30__SCAN_IN, P3_ADD_344_U126);
  not ginst18718 (P3_ADD_344_U98, P3_ADD_344_U7);
  not ginst18719 (P3_ADD_344_U99, P3_ADD_344_U9);
  not ginst18720 (P3_ADD_349_U10, P3_INSTADDRPOINTER_REG_3__SCAN_IN);
  not ginst18721 (P3_ADD_349_U100, P3_ADD_349_U11);
  not ginst18722 (P3_ADD_349_U101, P3_ADD_349_U13);
  not ginst18723 (P3_ADD_349_U102, P3_ADD_349_U15);
  not ginst18724 (P3_ADD_349_U103, P3_ADD_349_U17);
  not ginst18725 (P3_ADD_349_U104, P3_ADD_349_U19);
  not ginst18726 (P3_ADD_349_U105, P3_ADD_349_U22);
  not ginst18727 (P3_ADD_349_U106, P3_ADD_349_U23);
  not ginst18728 (P3_ADD_349_U107, P3_ADD_349_U25);
  not ginst18729 (P3_ADD_349_U108, P3_ADD_349_U27);
  not ginst18730 (P3_ADD_349_U109, P3_ADD_349_U29);
  nand ginst18731 (P3_ADD_349_U11, P3_INSTADDRPOINTER_REG_3__SCAN_IN, P3_ADD_349_U99);
  not ginst18732 (P3_ADD_349_U110, P3_ADD_349_U31);
  not ginst18733 (P3_ADD_349_U111, P3_ADD_349_U33);
  not ginst18734 (P3_ADD_349_U112, P3_ADD_349_U35);
  not ginst18735 (P3_ADD_349_U113, P3_ADD_349_U37);
  not ginst18736 (P3_ADD_349_U114, P3_ADD_349_U39);
  not ginst18737 (P3_ADD_349_U115, P3_ADD_349_U41);
  not ginst18738 (P3_ADD_349_U116, P3_ADD_349_U43);
  not ginst18739 (P3_ADD_349_U117, P3_ADD_349_U45);
  not ginst18740 (P3_ADD_349_U118, P3_ADD_349_U47);
  not ginst18741 (P3_ADD_349_U119, P3_ADD_349_U49);
  not ginst18742 (P3_ADD_349_U12, P3_INSTADDRPOINTER_REG_4__SCAN_IN);
  not ginst18743 (P3_ADD_349_U120, P3_ADD_349_U51);
  not ginst18744 (P3_ADD_349_U121, P3_ADD_349_U53);
  not ginst18745 (P3_ADD_349_U122, P3_ADD_349_U55);
  not ginst18746 (P3_ADD_349_U123, P3_ADD_349_U57);
  not ginst18747 (P3_ADD_349_U124, P3_ADD_349_U59);
  not ginst18748 (P3_ADD_349_U125, P3_ADD_349_U61);
  not ginst18749 (P3_ADD_349_U126, P3_ADD_349_U63);
  not ginst18750 (P3_ADD_349_U127, P3_ADD_349_U97);
  nand ginst18751 (P3_ADD_349_U128, P3_INSTADDRPOINTER_REG_9__SCAN_IN, P3_ADD_349_U22);
  nand ginst18752 (P3_ADD_349_U129, P3_ADD_349_U105, P3_ADD_349_U21);
  nand ginst18753 (P3_ADD_349_U13, P3_INSTADDRPOINTER_REG_4__SCAN_IN, P3_ADD_349_U100);
  nand ginst18754 (P3_ADD_349_U130, P3_INSTADDRPOINTER_REG_8__SCAN_IN, P3_ADD_349_U19);
  nand ginst18755 (P3_ADD_349_U131, P3_ADD_349_U104, P3_ADD_349_U20);
  nand ginst18756 (P3_ADD_349_U132, P3_INSTADDRPOINTER_REG_7__SCAN_IN, P3_ADD_349_U17);
  nand ginst18757 (P3_ADD_349_U133, P3_ADD_349_U103, P3_ADD_349_U18);
  nand ginst18758 (P3_ADD_349_U134, P3_INSTADDRPOINTER_REG_6__SCAN_IN, P3_ADD_349_U15);
  nand ginst18759 (P3_ADD_349_U135, P3_ADD_349_U102, P3_ADD_349_U16);
  nand ginst18760 (P3_ADD_349_U136, P3_INSTADDRPOINTER_REG_5__SCAN_IN, P3_ADD_349_U13);
  nand ginst18761 (P3_ADD_349_U137, P3_ADD_349_U101, P3_ADD_349_U14);
  nand ginst18762 (P3_ADD_349_U138, P3_INSTADDRPOINTER_REG_4__SCAN_IN, P3_ADD_349_U11);
  nand ginst18763 (P3_ADD_349_U139, P3_ADD_349_U100, P3_ADD_349_U12);
  not ginst18764 (P3_ADD_349_U14, P3_INSTADDRPOINTER_REG_5__SCAN_IN);
  nand ginst18765 (P3_ADD_349_U140, P3_INSTADDRPOINTER_REG_3__SCAN_IN, P3_ADD_349_U9);
  nand ginst18766 (P3_ADD_349_U141, P3_ADD_349_U10, P3_ADD_349_U99);
  nand ginst18767 (P3_ADD_349_U142, P3_INSTADDRPOINTER_REG_31__SCAN_IN, P3_ADD_349_U97);
  nand ginst18768 (P3_ADD_349_U143, P3_ADD_349_U127, P3_ADD_349_U96);
  nand ginst18769 (P3_ADD_349_U144, P3_INSTADDRPOINTER_REG_30__SCAN_IN, P3_ADD_349_U63);
  nand ginst18770 (P3_ADD_349_U145, P3_ADD_349_U126, P3_ADD_349_U64);
  nand ginst18771 (P3_ADD_349_U146, P3_INSTADDRPOINTER_REG_2__SCAN_IN, P3_ADD_349_U7);
  nand ginst18772 (P3_ADD_349_U147, P3_ADD_349_U8, P3_ADD_349_U98);
  nand ginst18773 (P3_ADD_349_U148, P3_INSTADDRPOINTER_REG_29__SCAN_IN, P3_ADD_349_U61);
  nand ginst18774 (P3_ADD_349_U149, P3_ADD_349_U125, P3_ADD_349_U62);
  nand ginst18775 (P3_ADD_349_U15, P3_INSTADDRPOINTER_REG_5__SCAN_IN, P3_ADD_349_U101);
  nand ginst18776 (P3_ADD_349_U150, P3_INSTADDRPOINTER_REG_28__SCAN_IN, P3_ADD_349_U59);
  nand ginst18777 (P3_ADD_349_U151, P3_ADD_349_U124, P3_ADD_349_U60);
  nand ginst18778 (P3_ADD_349_U152, P3_INSTADDRPOINTER_REG_27__SCAN_IN, P3_ADD_349_U57);
  nand ginst18779 (P3_ADD_349_U153, P3_ADD_349_U123, P3_ADD_349_U58);
  nand ginst18780 (P3_ADD_349_U154, P3_INSTADDRPOINTER_REG_26__SCAN_IN, P3_ADD_349_U55);
  nand ginst18781 (P3_ADD_349_U155, P3_ADD_349_U122, P3_ADD_349_U56);
  nand ginst18782 (P3_ADD_349_U156, P3_INSTADDRPOINTER_REG_25__SCAN_IN, P3_ADD_349_U53);
  nand ginst18783 (P3_ADD_349_U157, P3_ADD_349_U121, P3_ADD_349_U54);
  nand ginst18784 (P3_ADD_349_U158, P3_INSTADDRPOINTER_REG_24__SCAN_IN, P3_ADD_349_U51);
  nand ginst18785 (P3_ADD_349_U159, P3_ADD_349_U120, P3_ADD_349_U52);
  not ginst18786 (P3_ADD_349_U16, P3_INSTADDRPOINTER_REG_6__SCAN_IN);
  nand ginst18787 (P3_ADD_349_U160, P3_INSTADDRPOINTER_REG_23__SCAN_IN, P3_ADD_349_U49);
  nand ginst18788 (P3_ADD_349_U161, P3_ADD_349_U119, P3_ADD_349_U50);
  nand ginst18789 (P3_ADD_349_U162, P3_INSTADDRPOINTER_REG_22__SCAN_IN, P3_ADD_349_U47);
  nand ginst18790 (P3_ADD_349_U163, P3_ADD_349_U118, P3_ADD_349_U48);
  nand ginst18791 (P3_ADD_349_U164, P3_INSTADDRPOINTER_REG_21__SCAN_IN, P3_ADD_349_U45);
  nand ginst18792 (P3_ADD_349_U165, P3_ADD_349_U117, P3_ADD_349_U46);
  nand ginst18793 (P3_ADD_349_U166, P3_INSTADDRPOINTER_REG_20__SCAN_IN, P3_ADD_349_U43);
  nand ginst18794 (P3_ADD_349_U167, P3_ADD_349_U116, P3_ADD_349_U44);
  nand ginst18795 (P3_ADD_349_U168, P3_INSTADDRPOINTER_REG_1__SCAN_IN, P3_ADD_349_U5);
  nand ginst18796 (P3_ADD_349_U169, P3_INSTADDRPOINTER_REG_0__SCAN_IN, P3_ADD_349_U6);
  nand ginst18797 (P3_ADD_349_U17, P3_INSTADDRPOINTER_REG_6__SCAN_IN, P3_ADD_349_U102);
  nand ginst18798 (P3_ADD_349_U170, P3_INSTADDRPOINTER_REG_19__SCAN_IN, P3_ADD_349_U41);
  nand ginst18799 (P3_ADD_349_U171, P3_ADD_349_U115, P3_ADD_349_U42);
  nand ginst18800 (P3_ADD_349_U172, P3_INSTADDRPOINTER_REG_18__SCAN_IN, P3_ADD_349_U39);
  nand ginst18801 (P3_ADD_349_U173, P3_ADD_349_U114, P3_ADD_349_U40);
  nand ginst18802 (P3_ADD_349_U174, P3_INSTADDRPOINTER_REG_17__SCAN_IN, P3_ADD_349_U37);
  nand ginst18803 (P3_ADD_349_U175, P3_ADD_349_U113, P3_ADD_349_U38);
  nand ginst18804 (P3_ADD_349_U176, P3_INSTADDRPOINTER_REG_16__SCAN_IN, P3_ADD_349_U35);
  nand ginst18805 (P3_ADD_349_U177, P3_ADD_349_U112, P3_ADD_349_U36);
  nand ginst18806 (P3_ADD_349_U178, P3_INSTADDRPOINTER_REG_15__SCAN_IN, P3_ADD_349_U33);
  nand ginst18807 (P3_ADD_349_U179, P3_ADD_349_U111, P3_ADD_349_U34);
  not ginst18808 (P3_ADD_349_U18, P3_INSTADDRPOINTER_REG_7__SCAN_IN);
  nand ginst18809 (P3_ADD_349_U180, P3_INSTADDRPOINTER_REG_14__SCAN_IN, P3_ADD_349_U31);
  nand ginst18810 (P3_ADD_349_U181, P3_ADD_349_U110, P3_ADD_349_U32);
  nand ginst18811 (P3_ADD_349_U182, P3_INSTADDRPOINTER_REG_13__SCAN_IN, P3_ADD_349_U29);
  nand ginst18812 (P3_ADD_349_U183, P3_ADD_349_U109, P3_ADD_349_U30);
  nand ginst18813 (P3_ADD_349_U184, P3_INSTADDRPOINTER_REG_12__SCAN_IN, P3_ADD_349_U27);
  nand ginst18814 (P3_ADD_349_U185, P3_ADD_349_U108, P3_ADD_349_U28);
  nand ginst18815 (P3_ADD_349_U186, P3_INSTADDRPOINTER_REG_11__SCAN_IN, P3_ADD_349_U25);
  nand ginst18816 (P3_ADD_349_U187, P3_ADD_349_U107, P3_ADD_349_U26);
  nand ginst18817 (P3_ADD_349_U188, P3_INSTADDRPOINTER_REG_10__SCAN_IN, P3_ADD_349_U23);
  nand ginst18818 (P3_ADD_349_U189, P3_ADD_349_U106, P3_ADD_349_U24);
  nand ginst18819 (P3_ADD_349_U19, P3_INSTADDRPOINTER_REG_7__SCAN_IN, P3_ADD_349_U103);
  not ginst18820 (P3_ADD_349_U20, P3_INSTADDRPOINTER_REG_8__SCAN_IN);
  not ginst18821 (P3_ADD_349_U21, P3_INSTADDRPOINTER_REG_9__SCAN_IN);
  nand ginst18822 (P3_ADD_349_U22, P3_INSTADDRPOINTER_REG_8__SCAN_IN, P3_ADD_349_U104);
  nand ginst18823 (P3_ADD_349_U23, P3_INSTADDRPOINTER_REG_9__SCAN_IN, P3_ADD_349_U105);
  not ginst18824 (P3_ADD_349_U24, P3_INSTADDRPOINTER_REG_10__SCAN_IN);
  nand ginst18825 (P3_ADD_349_U25, P3_INSTADDRPOINTER_REG_10__SCAN_IN, P3_ADD_349_U106);
  not ginst18826 (P3_ADD_349_U26, P3_INSTADDRPOINTER_REG_11__SCAN_IN);
  nand ginst18827 (P3_ADD_349_U27, P3_INSTADDRPOINTER_REG_11__SCAN_IN, P3_ADD_349_U107);
  not ginst18828 (P3_ADD_349_U28, P3_INSTADDRPOINTER_REG_12__SCAN_IN);
  nand ginst18829 (P3_ADD_349_U29, P3_INSTADDRPOINTER_REG_12__SCAN_IN, P3_ADD_349_U108);
  not ginst18830 (P3_ADD_349_U30, P3_INSTADDRPOINTER_REG_13__SCAN_IN);
  nand ginst18831 (P3_ADD_349_U31, P3_INSTADDRPOINTER_REG_13__SCAN_IN, P3_ADD_349_U109);
  not ginst18832 (P3_ADD_349_U32, P3_INSTADDRPOINTER_REG_14__SCAN_IN);
  nand ginst18833 (P3_ADD_349_U33, P3_INSTADDRPOINTER_REG_14__SCAN_IN, P3_ADD_349_U110);
  not ginst18834 (P3_ADD_349_U34, P3_INSTADDRPOINTER_REG_15__SCAN_IN);
  nand ginst18835 (P3_ADD_349_U35, P3_INSTADDRPOINTER_REG_15__SCAN_IN, P3_ADD_349_U111);
  not ginst18836 (P3_ADD_349_U36, P3_INSTADDRPOINTER_REG_16__SCAN_IN);
  nand ginst18837 (P3_ADD_349_U37, P3_INSTADDRPOINTER_REG_16__SCAN_IN, P3_ADD_349_U112);
  not ginst18838 (P3_ADD_349_U38, P3_INSTADDRPOINTER_REG_17__SCAN_IN);
  nand ginst18839 (P3_ADD_349_U39, P3_INSTADDRPOINTER_REG_17__SCAN_IN, P3_ADD_349_U113);
  not ginst18840 (P3_ADD_349_U40, P3_INSTADDRPOINTER_REG_18__SCAN_IN);
  nand ginst18841 (P3_ADD_349_U41, P3_INSTADDRPOINTER_REG_18__SCAN_IN, P3_ADD_349_U114);
  not ginst18842 (P3_ADD_349_U42, P3_INSTADDRPOINTER_REG_19__SCAN_IN);
  nand ginst18843 (P3_ADD_349_U43, P3_INSTADDRPOINTER_REG_19__SCAN_IN, P3_ADD_349_U115);
  not ginst18844 (P3_ADD_349_U44, P3_INSTADDRPOINTER_REG_20__SCAN_IN);
  nand ginst18845 (P3_ADD_349_U45, P3_INSTADDRPOINTER_REG_20__SCAN_IN, P3_ADD_349_U116);
  not ginst18846 (P3_ADD_349_U46, P3_INSTADDRPOINTER_REG_21__SCAN_IN);
  nand ginst18847 (P3_ADD_349_U47, P3_INSTADDRPOINTER_REG_21__SCAN_IN, P3_ADD_349_U117);
  not ginst18848 (P3_ADD_349_U48, P3_INSTADDRPOINTER_REG_22__SCAN_IN);
  nand ginst18849 (P3_ADD_349_U49, P3_INSTADDRPOINTER_REG_22__SCAN_IN, P3_ADD_349_U118);
  not ginst18850 (P3_ADD_349_U5, P3_INSTADDRPOINTER_REG_0__SCAN_IN);
  not ginst18851 (P3_ADD_349_U50, P3_INSTADDRPOINTER_REG_23__SCAN_IN);
  nand ginst18852 (P3_ADD_349_U51, P3_INSTADDRPOINTER_REG_23__SCAN_IN, P3_ADD_349_U119);
  not ginst18853 (P3_ADD_349_U52, P3_INSTADDRPOINTER_REG_24__SCAN_IN);
  nand ginst18854 (P3_ADD_349_U53, P3_INSTADDRPOINTER_REG_24__SCAN_IN, P3_ADD_349_U120);
  not ginst18855 (P3_ADD_349_U54, P3_INSTADDRPOINTER_REG_25__SCAN_IN);
  nand ginst18856 (P3_ADD_349_U55, P3_INSTADDRPOINTER_REG_25__SCAN_IN, P3_ADD_349_U121);
  not ginst18857 (P3_ADD_349_U56, P3_INSTADDRPOINTER_REG_26__SCAN_IN);
  nand ginst18858 (P3_ADD_349_U57, P3_INSTADDRPOINTER_REG_26__SCAN_IN, P3_ADD_349_U122);
  not ginst18859 (P3_ADD_349_U58, P3_INSTADDRPOINTER_REG_27__SCAN_IN);
  nand ginst18860 (P3_ADD_349_U59, P3_INSTADDRPOINTER_REG_27__SCAN_IN, P3_ADD_349_U123);
  not ginst18861 (P3_ADD_349_U6, P3_INSTADDRPOINTER_REG_1__SCAN_IN);
  not ginst18862 (P3_ADD_349_U60, P3_INSTADDRPOINTER_REG_28__SCAN_IN);
  nand ginst18863 (P3_ADD_349_U61, P3_INSTADDRPOINTER_REG_28__SCAN_IN, P3_ADD_349_U124);
  not ginst18864 (P3_ADD_349_U62, P3_INSTADDRPOINTER_REG_29__SCAN_IN);
  nand ginst18865 (P3_ADD_349_U63, P3_INSTADDRPOINTER_REG_29__SCAN_IN, P3_ADD_349_U125);
  not ginst18866 (P3_ADD_349_U64, P3_INSTADDRPOINTER_REG_30__SCAN_IN);
  nand ginst18867 (P3_ADD_349_U65, P3_ADD_349_U128, P3_ADD_349_U129);
  nand ginst18868 (P3_ADD_349_U66, P3_ADD_349_U130, P3_ADD_349_U131);
  nand ginst18869 (P3_ADD_349_U67, P3_ADD_349_U132, P3_ADD_349_U133);
  nand ginst18870 (P3_ADD_349_U68, P3_ADD_349_U134, P3_ADD_349_U135);
  nand ginst18871 (P3_ADD_349_U69, P3_ADD_349_U136, P3_ADD_349_U137);
  nand ginst18872 (P3_ADD_349_U7, P3_INSTADDRPOINTER_REG_0__SCAN_IN, P3_INSTADDRPOINTER_REG_1__SCAN_IN);
  nand ginst18873 (P3_ADD_349_U70, P3_ADD_349_U138, P3_ADD_349_U139);
  nand ginst18874 (P3_ADD_349_U71, P3_ADD_349_U140, P3_ADD_349_U141);
  nand ginst18875 (P3_ADD_349_U72, P3_ADD_349_U142, P3_ADD_349_U143);
  nand ginst18876 (P3_ADD_349_U73, P3_ADD_349_U144, P3_ADD_349_U145);
  nand ginst18877 (P3_ADD_349_U74, P3_ADD_349_U146, P3_ADD_349_U147);
  nand ginst18878 (P3_ADD_349_U75, P3_ADD_349_U148, P3_ADD_349_U149);
  nand ginst18879 (P3_ADD_349_U76, P3_ADD_349_U150, P3_ADD_349_U151);
  nand ginst18880 (P3_ADD_349_U77, P3_ADD_349_U152, P3_ADD_349_U153);
  nand ginst18881 (P3_ADD_349_U78, P3_ADD_349_U154, P3_ADD_349_U155);
  nand ginst18882 (P3_ADD_349_U79, P3_ADD_349_U156, P3_ADD_349_U157);
  not ginst18883 (P3_ADD_349_U8, P3_INSTADDRPOINTER_REG_2__SCAN_IN);
  nand ginst18884 (P3_ADD_349_U80, P3_ADD_349_U158, P3_ADD_349_U159);
  nand ginst18885 (P3_ADD_349_U81, P3_ADD_349_U160, P3_ADD_349_U161);
  nand ginst18886 (P3_ADD_349_U82, P3_ADD_349_U162, P3_ADD_349_U163);
  nand ginst18887 (P3_ADD_349_U83, P3_ADD_349_U164, P3_ADD_349_U165);
  nand ginst18888 (P3_ADD_349_U84, P3_ADD_349_U166, P3_ADD_349_U167);
  nand ginst18889 (P3_ADD_349_U85, P3_ADD_349_U168, P3_ADD_349_U169);
  nand ginst18890 (P3_ADD_349_U86, P3_ADD_349_U170, P3_ADD_349_U171);
  nand ginst18891 (P3_ADD_349_U87, P3_ADD_349_U172, P3_ADD_349_U173);
  nand ginst18892 (P3_ADD_349_U88, P3_ADD_349_U174, P3_ADD_349_U175);
  nand ginst18893 (P3_ADD_349_U89, P3_ADD_349_U176, P3_ADD_349_U177);
  nand ginst18894 (P3_ADD_349_U9, P3_INSTADDRPOINTER_REG_2__SCAN_IN, P3_ADD_349_U98);
  nand ginst18895 (P3_ADD_349_U90, P3_ADD_349_U178, P3_ADD_349_U179);
  nand ginst18896 (P3_ADD_349_U91, P3_ADD_349_U180, P3_ADD_349_U181);
  nand ginst18897 (P3_ADD_349_U92, P3_ADD_349_U182, P3_ADD_349_U183);
  nand ginst18898 (P3_ADD_349_U93, P3_ADD_349_U184, P3_ADD_349_U185);
  nand ginst18899 (P3_ADD_349_U94, P3_ADD_349_U186, P3_ADD_349_U187);
  nand ginst18900 (P3_ADD_349_U95, P3_ADD_349_U188, P3_ADD_349_U189);
  not ginst18901 (P3_ADD_349_U96, P3_INSTADDRPOINTER_REG_31__SCAN_IN);
  nand ginst18902 (P3_ADD_349_U97, P3_INSTADDRPOINTER_REG_30__SCAN_IN, P3_ADD_349_U126);
  not ginst18903 (P3_ADD_349_U98, P3_ADD_349_U7);
  not ginst18904 (P3_ADD_349_U99, P3_ADD_349_U9);
  not ginst18905 (P3_ADD_357_U10, P3_SUB_357_U10);
  or ginst18906 (P3_ADD_357_U11, P3_SUB_357_U11, P3_SUB_357_U12, P3_SUB_357_U7);
  nand ginst18907 (P3_ADD_357_U12, P3_ADD_357_U14, P3_ADD_357_U22);
  nand ginst18908 (P3_ADD_357_U13, P3_ADD_357_U34, P3_ADD_357_U35);
  nor ginst18909 (P3_ADD_357_U14, P3_SUB_357_U13, P3_SUB_357_U9);
  nor ginst18910 (P3_ADD_357_U15, P3_SUB_357_U6, P3_SUB_357_U8);
  not ginst18911 (P3_ADD_357_U16, P3_SUB_357_U6);
  and ginst18912 (P3_ADD_357_U17, P3_ADD_357_U30, P3_ADD_357_U31);
  not ginst18913 (P3_ADD_357_U18, P3_SUB_357_U13);
  and ginst18914 (P3_ADD_357_U19, P3_ADD_357_U32, P3_ADD_357_U33);
  not ginst18915 (P3_ADD_357_U20, P3_SUB_357_U7);
  not ginst18916 (P3_ADD_357_U21, P3_SUB_357_U12);
  not ginst18917 (P3_ADD_357_U22, P3_ADD_357_U11);
  not ginst18918 (P3_ADD_357_U23, P3_ADD_357_U12);
  nand ginst18919 (P3_ADD_357_U24, P3_ADD_357_U16, P3_ADD_357_U23);
  nand ginst18920 (P3_ADD_357_U25, P3_ADD_357_U24, P3_SUB_357_U8);
  nand ginst18921 (P3_ADD_357_U26, P3_ADD_357_U18, P3_ADD_357_U22);
  nand ginst18922 (P3_ADD_357_U27, P3_ADD_357_U26, P3_SUB_357_U9);
  or ginst18923 (P3_ADD_357_U28, P3_SUB_357_U12, P3_SUB_357_U7);
  nand ginst18924 (P3_ADD_357_U29, P3_ADD_357_U28, P3_SUB_357_U11);
  nand ginst18925 (P3_ADD_357_U30, P3_ADD_357_U12, P3_SUB_357_U6);
  nand ginst18926 (P3_ADD_357_U31, P3_ADD_357_U16, P3_ADD_357_U23);
  nand ginst18927 (P3_ADD_357_U32, P3_ADD_357_U11, P3_SUB_357_U13);
  nand ginst18928 (P3_ADD_357_U33, P3_ADD_357_U18, P3_ADD_357_U22);
  nand ginst18929 (P3_ADD_357_U34, P3_ADD_357_U21, P3_SUB_357_U7);
  nand ginst18930 (P3_ADD_357_U35, P3_ADD_357_U20, P3_SUB_357_U12);
  nand ginst18931 (P3_ADD_357_U6, P3_ADD_357_U15, P3_ADD_357_U23);
  and ginst18932 (P3_ADD_357_U7, P3_ADD_357_U11, P3_ADD_357_U29);
  and ginst18933 (P3_ADD_357_U8, P3_ADD_357_U12, P3_ADD_357_U27);
  and ginst18934 (P3_ADD_357_U9, P3_ADD_357_U25, P3_ADD_357_U6);
  and ginst18935 (P3_ADD_360_1242_U10, P3_ADD_360_1242_U175, P3_ADD_360_1242_U58);
  and ginst18936 (P3_ADD_360_1242_U100, P3_INSTADDRPOINTER_REG_16__SCAN_IN, P3_INSTADDRPOINTER_REG_17__SCAN_IN);
  and ginst18937 (P3_ADD_360_1242_U101, P3_INSTADDRPOINTER_REG_18__SCAN_IN, P3_INSTADDRPOINTER_REG_19__SCAN_IN);
  and ginst18938 (P3_ADD_360_1242_U102, P3_INSTADDRPOINTER_REG_22__SCAN_IN, P3_INSTADDRPOINTER_REG_23__SCAN_IN);
  and ginst18939 (P3_ADD_360_1242_U103, P3_INSTADDRPOINTER_REG_24__SCAN_IN, P3_INSTADDRPOINTER_REG_25__SCAN_IN);
  and ginst18940 (P3_ADD_360_1242_U104, P3_INSTADDRPOINTER_REG_27__SCAN_IN, P3_INSTADDRPOINTER_REG_28__SCAN_IN);
  nand ginst18941 (P3_ADD_360_1242_U105, P3_ADD_360_1242_U146, P3_ADD_360_1242_U147);
  and ginst18942 (P3_ADD_360_1242_U106, P3_ADD_360_1242_U193, P3_ADD_360_1242_U194);
  and ginst18943 (P3_ADD_360_1242_U107, P3_ADD_360_1242_U195, P3_ADD_360_1242_U196);
  nand ginst18944 (P3_ADD_360_1242_U108, P3_ADD_360_1242_U120, P3_ADD_360_1242_U143, P3_ADD_360_1242_U189);
  and ginst18945 (P3_ADD_360_1242_U109, P3_ADD_360_1242_U202, P3_ADD_360_1242_U203);
  and ginst18946 (P3_ADD_360_1242_U11, P3_ADD_360_1242_U174, P3_ADD_360_1242_U60);
  nand ginst18947 (P3_ADD_360_1242_U110, P3_ADD_360_1242_U140, P3_ADD_360_1242_U141);
  and ginst18948 (P3_ADD_360_1242_U111, P3_ADD_360_1242_U209, P3_ADD_360_1242_U210);
  nand ginst18949 (P3_ADD_360_1242_U112, P3_ADD_360_1242_U121, P3_ADD_360_1242_U137, P3_ADD_360_1242_U188);
  and ginst18950 (P3_ADD_360_1242_U113, P3_ADD_360_1242_U216, P3_ADD_360_1242_U217);
  nand ginst18951 (P3_ADD_360_1242_U114, P3_ADD_360_1242_U191, P3_ADD_360_1242_U94);
  and ginst18952 (P3_ADD_360_1242_U115, P3_ADD_360_1242_U225, P3_ADD_360_1242_U226);
  not ginst18953 (P3_ADD_360_1242_U116, P3_INSTADDRPOINTER_REG_31__SCAN_IN);
  and ginst18954 (P3_ADD_360_1242_U117, P3_ADD_360_1242_U231, P3_ADD_360_1242_U232);
  nand ginst18955 (P3_ADD_360_1242_U118, P3_ADD_360_1242_U127, P3_ADD_360_1242_U75);
  not ginst18956 (P3_ADD_360_1242_U119, P3_ADD_360_1242_U45);
  and ginst18957 (P3_ADD_360_1242_U12, P3_ADD_360_1242_U173, P3_ADD_360_1242_U63);
  nand ginst18958 (P3_ADD_360_1242_U120, P3_INSTADDRPOINTER_REG_7__SCAN_IN, P3_ADD_360_1242_U110);
  nand ginst18959 (P3_ADD_360_1242_U121, P3_INSTADDRPOINTER_REG_5__SCAN_IN, P3_ADD_360_1242_U114);
  not ginst18960 (P3_ADD_360_1242_U122, P3_ADD_360_1242_U75);
  or ginst18961 (P3_ADD_360_1242_U123, P3_INSTADDRPOINTER_REG_4__SCAN_IN, P3_ADD_360_U19);
  not ginst18962 (P3_ADD_360_1242_U124, P3_ADD_360_1242_U27);
  nand ginst18963 (P3_ADD_360_1242_U125, P3_INSTADDRPOINTER_REG_4__SCAN_IN, P3_ADD_360_U19);
  nand ginst18964 (P3_ADD_360_1242_U126, P3_ADD_360_1242_U27, P3_ADD_360_1242_U28);
  nand ginst18965 (P3_ADD_360_1242_U127, P3_INSTADDRPOINTER_REG_1__SCAN_IN, P3_ADD_360_1242_U126);
  not ginst18966 (P3_ADD_360_1242_U128, P3_ADD_360_1242_U118);
  or ginst18967 (P3_ADD_360_1242_U129, P3_INSTADDRPOINTER_REG_2__SCAN_IN, P3_ADD_360_U21);
  and ginst18968 (P3_ADD_360_1242_U13, P3_ADD_360_1242_U171, P3_ADD_360_1242_U66);
  nand ginst18969 (P3_ADD_360_1242_U130, P3_ADD_360_1242_U118, P3_ADD_360_1242_U129);
  nand ginst18970 (P3_ADD_360_1242_U131, P3_INSTADDRPOINTER_REG_2__SCAN_IN, P3_ADD_360_U21);
  not ginst18971 (P3_ADD_360_1242_U132, P3_ADD_360_1242_U40);
  or ginst18972 (P3_ADD_360_1242_U133, P3_INSTADDRPOINTER_REG_3__SCAN_IN, P3_ADD_360_U20);
  not ginst18973 (P3_ADD_360_1242_U134, P3_ADD_360_1242_U41);
  nand ginst18974 (P3_ADD_360_1242_U135, P3_INSTADDRPOINTER_REG_3__SCAN_IN, P3_ADD_360_U20);
  not ginst18975 (P3_ADD_360_1242_U136, P3_ADD_360_1242_U114);
  nand ginst18976 (P3_ADD_360_1242_U137, P3_ADD_360_1242_U114, P3_ADD_360_U18);
  not ginst18977 (P3_ADD_360_1242_U138, P3_ADD_360_1242_U112);
  or ginst18978 (P3_ADD_360_1242_U139, P3_INSTADDRPOINTER_REG_6__SCAN_IN, P3_ADD_360_U17);
  and ginst18979 (P3_ADD_360_1242_U14, P3_ADD_360_1242_U169, P3_ADD_360_1242_U68);
  nand ginst18980 (P3_ADD_360_1242_U140, P3_ADD_360_1242_U112, P3_ADD_360_1242_U139);
  nand ginst18981 (P3_ADD_360_1242_U141, P3_INSTADDRPOINTER_REG_6__SCAN_IN, P3_ADD_360_U17);
  not ginst18982 (P3_ADD_360_1242_U142, P3_ADD_360_1242_U110);
  nand ginst18983 (P3_ADD_360_1242_U143, P3_ADD_360_1242_U110, P3_ADD_360_U16);
  not ginst18984 (P3_ADD_360_1242_U144, P3_ADD_360_1242_U108);
  or ginst18985 (P3_ADD_360_1242_U145, P3_INSTADDRPOINTER_REG_8__SCAN_IN, P3_ADD_360_U5);
  nand ginst18986 (P3_ADD_360_1242_U146, P3_ADD_360_1242_U108, P3_ADD_360_1242_U145);
  nand ginst18987 (P3_ADD_360_1242_U147, P3_INSTADDRPOINTER_REG_8__SCAN_IN, P3_ADD_360_U5);
  not ginst18988 (P3_ADD_360_1242_U148, P3_ADD_360_1242_U105);
  nand ginst18989 (P3_ADD_360_1242_U149, P3_ADD_360_1242_U41, P3_ADD_360_1242_U95);
  and ginst18990 (P3_ADD_360_1242_U15, P3_ADD_360_1242_U168, P3_ADD_360_1242_U71);
  nand ginst18991 (P3_ADD_360_1242_U150, P3_ADD_360_1242_U135, P3_ADD_360_1242_U41);
  nand ginst18992 (P3_ADD_360_1242_U151, P3_ADD_360_1242_U150, P3_ADD_360_1242_U96);
  nand ginst18993 (P3_ADD_360_1242_U152, P3_ADD_360_1242_U115, P3_ADD_360_1242_U132);
  nand ginst18994 (P3_ADD_360_1242_U153, P3_ADD_360_1242_U134, P3_ADD_360_1242_U135);
  not ginst18995 (P3_ADD_360_1242_U154, P3_ADD_360_1242_U46);
  not ginst18996 (P3_ADD_360_1242_U155, P3_ADD_360_1242_U76);
  not ginst18997 (P3_ADD_360_1242_U156, P3_ADD_360_1242_U50);
  not ginst18998 (P3_ADD_360_1242_U157, P3_ADD_360_1242_U53);
  not ginst18999 (P3_ADD_360_1242_U158, P3_ADD_360_1242_U56);
  not ginst19000 (P3_ADD_360_1242_U159, P3_ADD_360_1242_U58);
  and ginst19001 (P3_ADD_360_1242_U16, P3_ADD_360_1242_U166, P3_ADD_360_1242_U73);
  not ginst19002 (P3_ADD_360_1242_U160, P3_ADD_360_1242_U60);
  not ginst19003 (P3_ADD_360_1242_U161, P3_ADD_360_1242_U63);
  not ginst19004 (P3_ADD_360_1242_U162, P3_ADD_360_1242_U66);
  not ginst19005 (P3_ADD_360_1242_U163, P3_ADD_360_1242_U68);
  not ginst19006 (P3_ADD_360_1242_U164, P3_ADD_360_1242_U71);
  not ginst19007 (P3_ADD_360_1242_U165, P3_ADD_360_1242_U73);
  nand ginst19008 (P3_ADD_360_1242_U166, P3_ADD_360_1242_U71, P3_ADD_360_1242_U72);
  nand ginst19009 (P3_ADD_360_1242_U167, P3_INSTADDRPOINTER_REG_27__SCAN_IN, P3_ADD_360_1242_U163);
  nand ginst19010 (P3_ADD_360_1242_U168, P3_ADD_360_1242_U167, P3_ADD_360_1242_U69);
  nand ginst19011 (P3_ADD_360_1242_U169, P3_ADD_360_1242_U66, P3_ADD_360_1242_U67);
  and ginst19012 (P3_ADD_360_1242_U17, P3_ADD_360_1242_U152, P3_ADD_360_1242_U153);
  nand ginst19013 (P3_ADD_360_1242_U170, P3_INSTADDRPOINTER_REG_24__SCAN_IN, P3_ADD_360_1242_U161);
  nand ginst19014 (P3_ADD_360_1242_U171, P3_ADD_360_1242_U170, P3_ADD_360_1242_U64);
  nand ginst19015 (P3_ADD_360_1242_U172, P3_INSTADDRPOINTER_REG_22__SCAN_IN, P3_ADD_360_1242_U160);
  nand ginst19016 (P3_ADD_360_1242_U173, P3_ADD_360_1242_U172, P3_ADD_360_1242_U61);
  nand ginst19017 (P3_ADD_360_1242_U174, P3_ADD_360_1242_U58, P3_ADD_360_1242_U59);
  nand ginst19018 (P3_ADD_360_1242_U175, P3_ADD_360_1242_U56, P3_ADD_360_1242_U57);
  nand ginst19019 (P3_ADD_360_1242_U176, P3_INSTADDRPOINTER_REG_18__SCAN_IN, P3_ADD_360_1242_U157);
  nand ginst19020 (P3_ADD_360_1242_U177, P3_ADD_360_1242_U176, P3_ADD_360_1242_U55);
  nand ginst19021 (P3_ADD_360_1242_U178, P3_INSTADDRPOINTER_REG_16__SCAN_IN, P3_ADD_360_1242_U156);
  nand ginst19022 (P3_ADD_360_1242_U179, P3_ADD_360_1242_U178, P3_ADD_360_1242_U51);
  and ginst19023 (P3_ADD_360_1242_U18, P3_ADD_360_1242_U149, P3_ADD_360_1242_U151);
  nand ginst19024 (P3_ADD_360_1242_U180, P3_INSTADDRPOINTER_REG_14__SCAN_IN, P3_ADD_360_1242_U155);
  nand ginst19025 (P3_ADD_360_1242_U181, P3_ADD_360_1242_U180, P3_ADD_360_1242_U48);
  nand ginst19026 (P3_ADD_360_1242_U182, P3_ADD_360_1242_U46, P3_ADD_360_1242_U47);
  nand ginst19027 (P3_ADD_360_1242_U183, P3_INSTADDRPOINTER_REG_11__SCAN_IN, P3_ADD_360_1242_U119);
  nand ginst19028 (P3_ADD_360_1242_U184, P3_ADD_360_1242_U183, P3_ADD_360_1242_U44);
  nand ginst19029 (P3_ADD_360_1242_U185, P3_INSTADDRPOINTER_REG_9__SCAN_IN, P3_ADD_360_1242_U105);
  nand ginst19030 (P3_ADD_360_1242_U186, P3_ADD_360_1242_U185, P3_ADD_360_1242_U42);
  nand ginst19031 (P3_ADD_360_1242_U187, P3_INSTADDRPOINTER_REG_30__SCAN_IN, P3_ADD_360_1242_U165);
  nand ginst19032 (P3_ADD_360_1242_U188, P3_INSTADDRPOINTER_REG_5__SCAN_IN, P3_ADD_360_U18);
  nand ginst19033 (P3_ADD_360_1242_U189, P3_INSTADDRPOINTER_REG_7__SCAN_IN, P3_ADD_360_U16);
  nand ginst19034 (P3_ADD_360_1242_U19, P3_ADD_360_1242_U192, P3_ADD_360_1242_U247, P3_ADD_360_1242_U248);
  nand ginst19035 (P3_ADD_360_1242_U190, P3_ADD_360_1242_U123, P3_ADD_360_1242_U92);
  nand ginst19036 (P3_ADD_360_1242_U191, P3_ADD_360_1242_U40, P3_ADD_360_1242_U93);
  nand ginst19037 (P3_ADD_360_1242_U192, P3_INSTADDRPOINTER_REG_1__SCAN_IN, P3_ADD_360_1242_U122);
  nand ginst19038 (P3_ADD_360_1242_U193, P3_INSTADDRPOINTER_REG_9__SCAN_IN, P3_ADD_360_1242_U105);
  nand ginst19039 (P3_ADD_360_1242_U194, P3_ADD_360_1242_U148, P3_ADD_360_1242_U39);
  nand ginst19040 (P3_ADD_360_1242_U195, P3_INSTADDRPOINTER_REG_8__SCAN_IN, P3_ADD_360_1242_U37);
  nand ginst19041 (P3_ADD_360_1242_U196, P3_ADD_360_1242_U38, P3_ADD_360_U5);
  nand ginst19042 (P3_ADD_360_1242_U197, P3_INSTADDRPOINTER_REG_8__SCAN_IN, P3_ADD_360_1242_U37);
  nand ginst19043 (P3_ADD_360_1242_U198, P3_ADD_360_1242_U38, P3_ADD_360_U5);
  nand ginst19044 (P3_ADD_360_1242_U199, P3_ADD_360_1242_U197, P3_ADD_360_1242_U198);
  not ginst19045 (P3_ADD_360_1242_U20, P3_ADD_360_U19);
  nand ginst19046 (P3_ADD_360_1242_U200, P3_ADD_360_1242_U107, P3_ADD_360_1242_U108);
  nand ginst19047 (P3_ADD_360_1242_U201, P3_ADD_360_1242_U144, P3_ADD_360_1242_U199);
  nand ginst19048 (P3_ADD_360_1242_U202, P3_INSTADDRPOINTER_REG_7__SCAN_IN, P3_ADD_360_1242_U36);
  nand ginst19049 (P3_ADD_360_1242_U203, P3_ADD_360_1242_U35, P3_ADD_360_U16);
  nand ginst19050 (P3_ADD_360_1242_U204, P3_INSTADDRPOINTER_REG_7__SCAN_IN, P3_ADD_360_1242_U36);
  nand ginst19051 (P3_ADD_360_1242_U205, P3_ADD_360_1242_U35, P3_ADD_360_U16);
  nand ginst19052 (P3_ADD_360_1242_U206, P3_ADD_360_1242_U204, P3_ADD_360_1242_U205);
  nand ginst19053 (P3_ADD_360_1242_U207, P3_ADD_360_1242_U109, P3_ADD_360_1242_U110);
  nand ginst19054 (P3_ADD_360_1242_U208, P3_ADD_360_1242_U142, P3_ADD_360_1242_U206);
  nand ginst19055 (P3_ADD_360_1242_U209, P3_INSTADDRPOINTER_REG_6__SCAN_IN, P3_ADD_360_1242_U33);
  not ginst19056 (P3_ADD_360_1242_U21, P3_INSTADDRPOINTER_REG_4__SCAN_IN);
  nand ginst19057 (P3_ADD_360_1242_U210, P3_ADD_360_1242_U34, P3_ADD_360_U17);
  nand ginst19058 (P3_ADD_360_1242_U211, P3_INSTADDRPOINTER_REG_6__SCAN_IN, P3_ADD_360_1242_U33);
  nand ginst19059 (P3_ADD_360_1242_U212, P3_ADD_360_1242_U34, P3_ADD_360_U17);
  nand ginst19060 (P3_ADD_360_1242_U213, P3_ADD_360_1242_U211, P3_ADD_360_1242_U212);
  nand ginst19061 (P3_ADD_360_1242_U214, P3_ADD_360_1242_U111, P3_ADD_360_1242_U112);
  nand ginst19062 (P3_ADD_360_1242_U215, P3_ADD_360_1242_U138, P3_ADD_360_1242_U213);
  nand ginst19063 (P3_ADD_360_1242_U216, P3_INSTADDRPOINTER_REG_5__SCAN_IN, P3_ADD_360_1242_U32);
  nand ginst19064 (P3_ADD_360_1242_U217, P3_ADD_360_1242_U31, P3_ADD_360_U18);
  nand ginst19065 (P3_ADD_360_1242_U218, P3_INSTADDRPOINTER_REG_5__SCAN_IN, P3_ADD_360_1242_U32);
  nand ginst19066 (P3_ADD_360_1242_U219, P3_ADD_360_1242_U31, P3_ADD_360_U18);
  not ginst19067 (P3_ADD_360_1242_U22, P3_ADD_360_U20);
  nand ginst19068 (P3_ADD_360_1242_U220, P3_ADD_360_1242_U218, P3_ADD_360_1242_U219);
  nand ginst19069 (P3_ADD_360_1242_U221, P3_ADD_360_1242_U113, P3_ADD_360_1242_U114);
  nand ginst19070 (P3_ADD_360_1242_U222, P3_ADD_360_1242_U136, P3_ADD_360_1242_U220);
  nand ginst19071 (P3_ADD_360_1242_U223, P3_INSTADDRPOINTER_REG_4__SCAN_IN, P3_ADD_360_1242_U20);
  nand ginst19072 (P3_ADD_360_1242_U224, P3_ADD_360_1242_U21, P3_ADD_360_U19);
  nand ginst19073 (P3_ADD_360_1242_U225, P3_INSTADDRPOINTER_REG_3__SCAN_IN, P3_ADD_360_1242_U22);
  nand ginst19074 (P3_ADD_360_1242_U226, P3_ADD_360_1242_U23, P3_ADD_360_U20);
  nand ginst19075 (P3_ADD_360_1242_U227, P3_INSTADDRPOINTER_REG_31__SCAN_IN, P3_ADD_360_1242_U187);
  nand ginst19076 (P3_ADD_360_1242_U228, P3_INSTADDRPOINTER_REG_30__SCAN_IN, P3_ADD_360_1242_U116, P3_ADD_360_1242_U165);
  nand ginst19077 (P3_ADD_360_1242_U229, P3_INSTADDRPOINTER_REG_30__SCAN_IN, P3_ADD_360_1242_U73);
  not ginst19078 (P3_ADD_360_1242_U23, P3_INSTADDRPOINTER_REG_3__SCAN_IN);
  nand ginst19079 (P3_ADD_360_1242_U230, P3_ADD_360_1242_U165, P3_ADD_360_1242_U74);
  nand ginst19080 (P3_ADD_360_1242_U231, P3_INSTADDRPOINTER_REG_2__SCAN_IN, P3_ADD_360_1242_U29);
  nand ginst19081 (P3_ADD_360_1242_U232, P3_ADD_360_1242_U30, P3_ADD_360_U21);
  nand ginst19082 (P3_ADD_360_1242_U233, P3_INSTADDRPOINTER_REG_2__SCAN_IN, P3_ADD_360_1242_U29);
  nand ginst19083 (P3_ADD_360_1242_U234, P3_ADD_360_1242_U30, P3_ADD_360_U21);
  nand ginst19084 (P3_ADD_360_1242_U235, P3_ADD_360_1242_U233, P3_ADD_360_1242_U234);
  nand ginst19085 (P3_ADD_360_1242_U236, P3_ADD_360_1242_U117, P3_ADD_360_1242_U118);
  nand ginst19086 (P3_ADD_360_1242_U237, P3_ADD_360_1242_U128, P3_ADD_360_1242_U235);
  nand ginst19087 (P3_ADD_360_1242_U238, P3_INSTADDRPOINTER_REG_27__SCAN_IN, P3_ADD_360_1242_U68);
  nand ginst19088 (P3_ADD_360_1242_U239, P3_ADD_360_1242_U163, P3_ADD_360_1242_U70);
  not ginst19089 (P3_ADD_360_1242_U24, P3_U2621);
  nand ginst19090 (P3_ADD_360_1242_U240, P3_INSTADDRPOINTER_REG_24__SCAN_IN, P3_ADD_360_1242_U63);
  nand ginst19091 (P3_ADD_360_1242_U241, P3_ADD_360_1242_U161, P3_ADD_360_1242_U65);
  nand ginst19092 (P3_ADD_360_1242_U242, P3_INSTADDRPOINTER_REG_22__SCAN_IN, P3_ADD_360_1242_U60);
  nand ginst19093 (P3_ADD_360_1242_U243, P3_ADD_360_1242_U160, P3_ADD_360_1242_U62);
  nand ginst19094 (P3_ADD_360_1242_U244, P3_INSTADDRPOINTER_REG_1__SCAN_IN, P3_ADD_360_1242_U27);
  nand ginst19095 (P3_ADD_360_1242_U245, P3_ADD_360_1242_U124, P3_ADD_360_1242_U26);
  nand ginst19096 (P3_ADD_360_1242_U246, P3_ADD_360_1242_U244, P3_ADD_360_1242_U245);
  nand ginst19097 (P3_ADD_360_1242_U247, P3_ADD_360_1242_U26, P3_ADD_360_1242_U27, P3_ADD_360_U4);
  nand ginst19098 (P3_ADD_360_1242_U248, P3_ADD_360_1242_U246, P3_ADD_360_1242_U28);
  nand ginst19099 (P3_ADD_360_1242_U249, P3_INSTADDRPOINTER_REG_18__SCAN_IN, P3_ADD_360_1242_U53);
  not ginst19100 (P3_ADD_360_1242_U25, P3_INSTADDRPOINTER_REG_0__SCAN_IN);
  nand ginst19101 (P3_ADD_360_1242_U250, P3_ADD_360_1242_U157, P3_ADD_360_1242_U54);
  nand ginst19102 (P3_ADD_360_1242_U251, P3_INSTADDRPOINTER_REG_16__SCAN_IN, P3_ADD_360_1242_U50);
  nand ginst19103 (P3_ADD_360_1242_U252, P3_ADD_360_1242_U156, P3_ADD_360_1242_U52);
  nand ginst19104 (P3_ADD_360_1242_U253, P3_INSTADDRPOINTER_REG_14__SCAN_IN, P3_ADD_360_1242_U76);
  nand ginst19105 (P3_ADD_360_1242_U254, P3_ADD_360_1242_U155, P3_ADD_360_1242_U49);
  nand ginst19106 (P3_ADD_360_1242_U255, P3_ADD_360_1242_U119, P3_ADD_360_1242_U43);
  nand ginst19107 (P3_ADD_360_1242_U256, P3_INSTADDRPOINTER_REG_11__SCAN_IN, P3_ADD_360_1242_U45);
  nand ginst19108 (P3_ADD_360_1242_U257, P3_INSTADDRPOINTER_REG_0__SCAN_IN, P3_ADD_360_1242_U24);
  nand ginst19109 (P3_ADD_360_1242_U258, P3_ADD_360_1242_U25, P3_U2621);
  not ginst19110 (P3_ADD_360_1242_U26, P3_INSTADDRPOINTER_REG_1__SCAN_IN);
  nand ginst19111 (P3_ADD_360_1242_U27, P3_INSTADDRPOINTER_REG_0__SCAN_IN, P3_U2621);
  not ginst19112 (P3_ADD_360_1242_U28, P3_ADD_360_U4);
  not ginst19113 (P3_ADD_360_1242_U29, P3_ADD_360_U21);
  not ginst19114 (P3_ADD_360_1242_U30, P3_INSTADDRPOINTER_REG_2__SCAN_IN);
  not ginst19115 (P3_ADD_360_1242_U31, P3_INSTADDRPOINTER_REG_5__SCAN_IN);
  not ginst19116 (P3_ADD_360_1242_U32, P3_ADD_360_U18);
  not ginst19117 (P3_ADD_360_1242_U33, P3_ADD_360_U17);
  not ginst19118 (P3_ADD_360_1242_U34, P3_INSTADDRPOINTER_REG_6__SCAN_IN);
  not ginst19119 (P3_ADD_360_1242_U35, P3_INSTADDRPOINTER_REG_7__SCAN_IN);
  not ginst19120 (P3_ADD_360_1242_U36, P3_ADD_360_U16);
  not ginst19121 (P3_ADD_360_1242_U37, P3_ADD_360_U5);
  not ginst19122 (P3_ADD_360_1242_U38, P3_INSTADDRPOINTER_REG_8__SCAN_IN);
  not ginst19123 (P3_ADD_360_1242_U39, P3_INSTADDRPOINTER_REG_9__SCAN_IN);
  and ginst19124 (P3_ADD_360_1242_U4, P3_ADD_360_1242_U186, P3_ADD_360_1242_U45);
  nand ginst19125 (P3_ADD_360_1242_U40, P3_ADD_360_1242_U130, P3_ADD_360_1242_U131);
  nand ginst19126 (P3_ADD_360_1242_U41, P3_ADD_360_1242_U133, P3_ADD_360_1242_U40);
  not ginst19127 (P3_ADD_360_1242_U42, P3_INSTADDRPOINTER_REG_10__SCAN_IN);
  not ginst19128 (P3_ADD_360_1242_U43, P3_INSTADDRPOINTER_REG_11__SCAN_IN);
  not ginst19129 (P3_ADD_360_1242_U44, P3_INSTADDRPOINTER_REG_12__SCAN_IN);
  nand ginst19130 (P3_ADD_360_1242_U45, P3_ADD_360_1242_U105, P3_ADD_360_1242_U97);
  nand ginst19131 (P3_ADD_360_1242_U46, P3_ADD_360_1242_U119, P3_ADD_360_1242_U98);
  not ginst19132 (P3_ADD_360_1242_U47, P3_INSTADDRPOINTER_REG_13__SCAN_IN);
  not ginst19133 (P3_ADD_360_1242_U48, P3_INSTADDRPOINTER_REG_15__SCAN_IN);
  not ginst19134 (P3_ADD_360_1242_U49, P3_INSTADDRPOINTER_REG_14__SCAN_IN);
  and ginst19135 (P3_ADD_360_1242_U5, P3_ADD_360_1242_U184, P3_ADD_360_1242_U46);
  nand ginst19136 (P3_ADD_360_1242_U50, P3_ADD_360_1242_U154, P3_ADD_360_1242_U99);
  not ginst19137 (P3_ADD_360_1242_U51, P3_INSTADDRPOINTER_REG_17__SCAN_IN);
  not ginst19138 (P3_ADD_360_1242_U52, P3_INSTADDRPOINTER_REG_16__SCAN_IN);
  nand ginst19139 (P3_ADD_360_1242_U53, P3_ADD_360_1242_U100, P3_ADD_360_1242_U156);
  not ginst19140 (P3_ADD_360_1242_U54, P3_INSTADDRPOINTER_REG_18__SCAN_IN);
  not ginst19141 (P3_ADD_360_1242_U55, P3_INSTADDRPOINTER_REG_19__SCAN_IN);
  nand ginst19142 (P3_ADD_360_1242_U56, P3_ADD_360_1242_U101, P3_ADD_360_1242_U157);
  not ginst19143 (P3_ADD_360_1242_U57, P3_INSTADDRPOINTER_REG_20__SCAN_IN);
  nand ginst19144 (P3_ADD_360_1242_U58, P3_INSTADDRPOINTER_REG_20__SCAN_IN, P3_ADD_360_1242_U158);
  not ginst19145 (P3_ADD_360_1242_U59, P3_INSTADDRPOINTER_REG_21__SCAN_IN);
  and ginst19146 (P3_ADD_360_1242_U6, P3_ADD_360_1242_U182, P3_ADD_360_1242_U76);
  nand ginst19147 (P3_ADD_360_1242_U60, P3_INSTADDRPOINTER_REG_21__SCAN_IN, P3_ADD_360_1242_U159);
  not ginst19148 (P3_ADD_360_1242_U61, P3_INSTADDRPOINTER_REG_23__SCAN_IN);
  not ginst19149 (P3_ADD_360_1242_U62, P3_INSTADDRPOINTER_REG_22__SCAN_IN);
  nand ginst19150 (P3_ADD_360_1242_U63, P3_ADD_360_1242_U102, P3_ADD_360_1242_U160);
  not ginst19151 (P3_ADD_360_1242_U64, P3_INSTADDRPOINTER_REG_25__SCAN_IN);
  not ginst19152 (P3_ADD_360_1242_U65, P3_INSTADDRPOINTER_REG_24__SCAN_IN);
  nand ginst19153 (P3_ADD_360_1242_U66, P3_ADD_360_1242_U103, P3_ADD_360_1242_U161);
  not ginst19154 (P3_ADD_360_1242_U67, P3_INSTADDRPOINTER_REG_26__SCAN_IN);
  nand ginst19155 (P3_ADD_360_1242_U68, P3_INSTADDRPOINTER_REG_26__SCAN_IN, P3_ADD_360_1242_U162);
  not ginst19156 (P3_ADD_360_1242_U69, P3_INSTADDRPOINTER_REG_28__SCAN_IN);
  and ginst19157 (P3_ADD_360_1242_U7, P3_ADD_360_1242_U181, P3_ADD_360_1242_U50);
  not ginst19158 (P3_ADD_360_1242_U70, P3_INSTADDRPOINTER_REG_27__SCAN_IN);
  nand ginst19159 (P3_ADD_360_1242_U71, P3_ADD_360_1242_U104, P3_ADD_360_1242_U163);
  not ginst19160 (P3_ADD_360_1242_U72, P3_INSTADDRPOINTER_REG_29__SCAN_IN);
  nand ginst19161 (P3_ADD_360_1242_U73, P3_INSTADDRPOINTER_REG_29__SCAN_IN, P3_ADD_360_1242_U164);
  not ginst19162 (P3_ADD_360_1242_U74, P3_INSTADDRPOINTER_REG_30__SCAN_IN);
  nand ginst19163 (P3_ADD_360_1242_U75, P3_ADD_360_1242_U124, P3_ADD_360_U4);
  nand ginst19164 (P3_ADD_360_1242_U76, P3_INSTADDRPOINTER_REG_13__SCAN_IN, P3_ADD_360_1242_U154);
  nand ginst19165 (P3_ADD_360_1242_U77, P3_ADD_360_1242_U229, P3_ADD_360_1242_U230);
  nand ginst19166 (P3_ADD_360_1242_U78, P3_ADD_360_1242_U238, P3_ADD_360_1242_U239);
  nand ginst19167 (P3_ADD_360_1242_U79, P3_ADD_360_1242_U240, P3_ADD_360_1242_U241);
  and ginst19168 (P3_ADD_360_1242_U8, P3_ADD_360_1242_U179, P3_ADD_360_1242_U53);
  nand ginst19169 (P3_ADD_360_1242_U80, P3_ADD_360_1242_U242, P3_ADD_360_1242_U243);
  nand ginst19170 (P3_ADD_360_1242_U81, P3_ADD_360_1242_U249, P3_ADD_360_1242_U250);
  nand ginst19171 (P3_ADD_360_1242_U82, P3_ADD_360_1242_U251, P3_ADD_360_1242_U252);
  nand ginst19172 (P3_ADD_360_1242_U83, P3_ADD_360_1242_U253, P3_ADD_360_1242_U254);
  nand ginst19173 (P3_ADD_360_1242_U84, P3_ADD_360_1242_U255, P3_ADD_360_1242_U256);
  nand ginst19174 (P3_ADD_360_1242_U85, P3_ADD_360_1242_U257, P3_ADD_360_1242_U258);
  nand ginst19175 (P3_ADD_360_1242_U86, P3_ADD_360_1242_U200, P3_ADD_360_1242_U201);
  nand ginst19176 (P3_ADD_360_1242_U87, P3_ADD_360_1242_U207, P3_ADD_360_1242_U208);
  nand ginst19177 (P3_ADD_360_1242_U88, P3_ADD_360_1242_U214, P3_ADD_360_1242_U215);
  nand ginst19178 (P3_ADD_360_1242_U89, P3_ADD_360_1242_U221, P3_ADD_360_1242_U222);
  and ginst19179 (P3_ADD_360_1242_U9, P3_ADD_360_1242_U177, P3_ADD_360_1242_U56);
  nand ginst19180 (P3_ADD_360_1242_U90, P3_ADD_360_1242_U227, P3_ADD_360_1242_U228);
  nand ginst19181 (P3_ADD_360_1242_U91, P3_ADD_360_1242_U236, P3_ADD_360_1242_U237);
  and ginst19182 (P3_ADD_360_1242_U92, P3_INSTADDRPOINTER_REG_3__SCAN_IN, P3_ADD_360_U20);
  and ginst19183 (P3_ADD_360_1242_U93, P3_ADD_360_1242_U123, P3_ADD_360_1242_U133);
  and ginst19184 (P3_ADD_360_1242_U94, P3_ADD_360_1242_U125, P3_ADD_360_1242_U190);
  and ginst19185 (P3_ADD_360_1242_U95, P3_ADD_360_1242_U135, P3_ADD_360_1242_U223, P3_ADD_360_1242_U224);
  and ginst19186 (P3_ADD_360_1242_U96, P3_ADD_360_1242_U123, P3_ADD_360_1242_U125);
  and ginst19187 (P3_ADD_360_1242_U97, P3_INSTADDRPOINTER_REG_9__SCAN_IN, P3_INSTADDRPOINTER_REG_10__SCAN_IN);
  and ginst19188 (P3_ADD_360_1242_U98, P3_INSTADDRPOINTER_REG_11__SCAN_IN, P3_INSTADDRPOINTER_REG_12__SCAN_IN);
  and ginst19189 (P3_ADD_360_1242_U99, P3_INSTADDRPOINTER_REG_13__SCAN_IN, P3_INSTADDRPOINTER_REG_14__SCAN_IN, P3_INSTADDRPOINTER_REG_15__SCAN_IN);
  not ginst19190 (P3_ADD_360_U10, P3_U2625);
  nand ginst19191 (P3_ADD_360_U11, P3_ADD_360_U25, P3_U2625);
  not ginst19192 (P3_ADD_360_U12, P3_U2626);
  nand ginst19193 (P3_ADD_360_U13, P3_ADD_360_U26, P3_U2626);
  not ginst19194 (P3_ADD_360_U14, P3_U2628);
  not ginst19195 (P3_ADD_360_U15, P3_U2627);
  nand ginst19196 (P3_ADD_360_U16, P3_ADD_360_U29, P3_ADD_360_U30);
  nand ginst19197 (P3_ADD_360_U17, P3_ADD_360_U31, P3_ADD_360_U32);
  nand ginst19198 (P3_ADD_360_U18, P3_ADD_360_U33, P3_ADD_360_U34);
  nand ginst19199 (P3_ADD_360_U19, P3_ADD_360_U35, P3_ADD_360_U36);
  nand ginst19200 (P3_ADD_360_U20, P3_ADD_360_U37, P3_ADD_360_U38);
  nand ginst19201 (P3_ADD_360_U21, P3_ADD_360_U39, P3_ADD_360_U40);
  and ginst19202 (P3_ADD_360_U22, P3_U2627, P3_U2628);
  nand ginst19203 (P3_ADD_360_U23, P3_ADD_360_U27, P3_U2627);
  not ginst19204 (P3_ADD_360_U24, P3_ADD_360_U7);
  not ginst19205 (P3_ADD_360_U25, P3_ADD_360_U9);
  not ginst19206 (P3_ADD_360_U26, P3_ADD_360_U11);
  not ginst19207 (P3_ADD_360_U27, P3_ADD_360_U13);
  not ginst19208 (P3_ADD_360_U28, P3_ADD_360_U23);
  nand ginst19209 (P3_ADD_360_U29, P3_ADD_360_U23, P3_U2628);
  nand ginst19210 (P3_ADD_360_U30, P3_ADD_360_U14, P3_ADD_360_U28);
  nand ginst19211 (P3_ADD_360_U31, P3_ADD_360_U13, P3_U2627);
  nand ginst19212 (P3_ADD_360_U32, P3_ADD_360_U15, P3_ADD_360_U27);
  nand ginst19213 (P3_ADD_360_U33, P3_ADD_360_U11, P3_U2626);
  nand ginst19214 (P3_ADD_360_U34, P3_ADD_360_U12, P3_ADD_360_U26);
  nand ginst19215 (P3_ADD_360_U35, P3_ADD_360_U9, P3_U2625);
  nand ginst19216 (P3_ADD_360_U36, P3_ADD_360_U10, P3_ADD_360_U25);
  nand ginst19217 (P3_ADD_360_U37, P3_ADD_360_U7, P3_U2624);
  nand ginst19218 (P3_ADD_360_U38, P3_ADD_360_U24, P3_ADD_360_U8);
  nand ginst19219 (P3_ADD_360_U39, P3_ADD_360_U4, P3_U2623);
  not ginst19220 (P3_ADD_360_U4, P3_U2622);
  nand ginst19221 (P3_ADD_360_U40, P3_ADD_360_U6, P3_U2622);
  and ginst19222 (P3_ADD_360_U5, P3_ADD_360_U22, P3_ADD_360_U27);
  not ginst19223 (P3_ADD_360_U6, P3_U2623);
  nand ginst19224 (P3_ADD_360_U7, P3_U2622, P3_U2623);
  not ginst19225 (P3_ADD_360_U8, P3_U2624);
  nand ginst19226 (P3_ADD_360_U9, P3_ADD_360_U24, P3_U2624);
  and ginst19227 (P3_ADD_371_1212_U10, P3_ADD_371_1212_U187, P3_ADD_371_1212_U59);
  and ginst19228 (P3_ADD_371_1212_U100, P3_INSTADDRPOINTER_REG_11__SCAN_IN, P3_INSTADDRPOINTER_REG_12__SCAN_IN);
  and ginst19229 (P3_ADD_371_1212_U101, P3_INSTADDRPOINTER_REG_13__SCAN_IN, P3_INSTADDRPOINTER_REG_14__SCAN_IN, P3_INSTADDRPOINTER_REG_15__SCAN_IN);
  and ginst19230 (P3_ADD_371_1212_U102, P3_INSTADDRPOINTER_REG_16__SCAN_IN, P3_INSTADDRPOINTER_REG_17__SCAN_IN);
  and ginst19231 (P3_ADD_371_1212_U103, P3_INSTADDRPOINTER_REG_18__SCAN_IN, P3_INSTADDRPOINTER_REG_19__SCAN_IN);
  and ginst19232 (P3_ADD_371_1212_U104, P3_INSTADDRPOINTER_REG_20__SCAN_IN, P3_INSTADDRPOINTER_REG_21__SCAN_IN);
  and ginst19233 (P3_ADD_371_1212_U105, P3_INSTADDRPOINTER_REG_22__SCAN_IN, P3_INSTADDRPOINTER_REG_23__SCAN_IN);
  and ginst19234 (P3_ADD_371_1212_U106, P3_INSTADDRPOINTER_REG_24__SCAN_IN, P3_INSTADDRPOINTER_REG_25__SCAN_IN);
  and ginst19235 (P3_ADD_371_1212_U107, P3_INSTADDRPOINTER_REG_27__SCAN_IN, P3_INSTADDRPOINTER_REG_28__SCAN_IN);
  nand ginst19236 (P3_ADD_371_1212_U108, P3_ADD_371_1212_U147, P3_ADD_371_1212_U148);
  and ginst19237 (P3_ADD_371_1212_U109, P3_ADD_371_1212_U204, P3_ADD_371_1212_U205);
  and ginst19238 (P3_ADD_371_1212_U11, P3_ADD_371_1212_U168, P3_ADD_371_1212_U185);
  and ginst19239 (P3_ADD_371_1212_U110, P3_ADD_371_1212_U206, P3_ADD_371_1212_U207);
  nand ginst19240 (P3_ADD_371_1212_U111, P3_ADD_371_1212_U118, P3_ADD_371_1212_U144, P3_ADD_371_1212_U200);
  and ginst19241 (P3_ADD_371_1212_U112, P3_ADD_371_1212_U213, P3_ADD_371_1212_U214);
  nand ginst19242 (P3_ADD_371_1212_U113, P3_ADD_371_1212_U141, P3_ADD_371_1212_U142);
  and ginst19243 (P3_ADD_371_1212_U114, P3_ADD_371_1212_U220, P3_ADD_371_1212_U221);
  nand ginst19244 (P3_ADD_371_1212_U115, P3_ADD_371_1212_U138, P3_ADD_371_1212_U95);
  not ginst19245 (P3_ADD_371_1212_U116, P3_INSTADDRPOINTER_REG_31__SCAN_IN);
  not ginst19246 (P3_ADD_371_1212_U117, P3_ADD_371_1212_U48);
  nand ginst19247 (P3_ADD_371_1212_U118, P3_INSTADDRPOINTER_REG_7__SCAN_IN, P3_ADD_371_1212_U113);
  nand ginst19248 (P3_ADD_371_1212_U119, P3_ADD_371_1212_U201, P3_ADD_371_1212_U202);
  and ginst19249 (P3_ADD_371_1212_U12, P3_ADD_371_1212_U184, P3_ADD_371_1212_U62);
  not ginst19250 (P3_ADD_371_1212_U120, P3_ADD_371_1212_U77);
  not ginst19251 (P3_ADD_371_1212_U121, P3_ADD_371_1212_U34);
  nand ginst19252 (P3_ADD_371_1212_U122, P3_ADD_371_1212_U34, P3_ADD_371_1212_U35);
  nand ginst19253 (P3_ADD_371_1212_U123, P3_INSTADDRPOINTER_REG_1__SCAN_IN, P3_ADD_371_1212_U122);
  not ginst19254 (P3_ADD_371_1212_U124, P3_ADD_371_1212_U44);
  or ginst19255 (P3_ADD_371_1212_U125, P3_INSTADDRPOINTER_REG_2__SCAN_IN, P3_ADD_371_U5);
  not ginst19256 (P3_ADD_371_1212_U126, P3_ADD_371_1212_U29);
  nand ginst19257 (P3_ADD_371_1212_U127, P3_ADD_371_1212_U29, P3_ADD_371_1212_U30);
  nand ginst19258 (P3_ADD_371_1212_U128, P3_INSTADDRPOINTER_REG_3__SCAN_IN, P3_ADD_371_1212_U127);
  nand ginst19259 (P3_ADD_371_1212_U129, P3_ADD_371_1212_U126, P3_ADD_371_U25);
  and ginst19260 (P3_ADD_371_1212_U13, P3_ADD_371_1212_U183, P3_ADD_371_1212_U65);
  nand ginst19261 (P3_ADD_371_1212_U130, P3_ADD_371_1212_U119, P3_ADD_371_1212_U44);
  not ginst19262 (P3_ADD_371_1212_U131, P3_ADD_371_1212_U43);
  or ginst19263 (P3_ADD_371_1212_U132, P3_INSTADDRPOINTER_REG_5__SCAN_IN, P3_ADD_371_U19);
  or ginst19264 (P3_ADD_371_1212_U133, P3_INSTADDRPOINTER_REG_4__SCAN_IN, P3_ADD_371_U20);
  not ginst19265 (P3_ADD_371_1212_U134, P3_ADD_371_1212_U24);
  nand ginst19266 (P3_ADD_371_1212_U135, P3_ADD_371_1212_U24, P3_ADD_371_1212_U25);
  nand ginst19267 (P3_ADD_371_1212_U136, P3_INSTADDRPOINTER_REG_5__SCAN_IN, P3_ADD_371_1212_U135);
  nand ginst19268 (P3_ADD_371_1212_U137, P3_ADD_371_1212_U134, P3_ADD_371_U19);
  nand ginst19269 (P3_ADD_371_1212_U138, P3_ADD_371_1212_U4, P3_ADD_371_1212_U43);
  not ginst19270 (P3_ADD_371_1212_U139, P3_ADD_371_1212_U115);
  and ginst19271 (P3_ADD_371_1212_U14, P3_ADD_371_1212_U181, P3_ADD_371_1212_U68);
  or ginst19272 (P3_ADD_371_1212_U140, P3_INSTADDRPOINTER_REG_6__SCAN_IN, P3_ADD_371_U18);
  nand ginst19273 (P3_ADD_371_1212_U141, P3_ADD_371_1212_U115, P3_ADD_371_1212_U140);
  nand ginst19274 (P3_ADD_371_1212_U142, P3_INSTADDRPOINTER_REG_6__SCAN_IN, P3_ADD_371_U18);
  not ginst19275 (P3_ADD_371_1212_U143, P3_ADD_371_1212_U113);
  nand ginst19276 (P3_ADD_371_1212_U144, P3_ADD_371_1212_U113, P3_ADD_371_U17);
  not ginst19277 (P3_ADD_371_1212_U145, P3_ADD_371_1212_U111);
  or ginst19278 (P3_ADD_371_1212_U146, P3_INSTADDRPOINTER_REG_8__SCAN_IN, P3_ADD_371_U6);
  nand ginst19279 (P3_ADD_371_1212_U147, P3_ADD_371_1212_U111, P3_ADD_371_1212_U146);
  nand ginst19280 (P3_ADD_371_1212_U148, P3_INSTADDRPOINTER_REG_8__SCAN_IN, P3_ADD_371_U6);
  not ginst19281 (P3_ADD_371_1212_U149, P3_ADD_371_1212_U108);
  and ginst19282 (P3_ADD_371_1212_U15, P3_ADD_371_1212_U179, P3_ADD_371_1212_U70);
  or ginst19283 (P3_ADD_371_1212_U150, P3_INSTADDRPOINTER_REG_4__SCAN_IN, P3_ADD_371_U20);
  nand ginst19284 (P3_ADD_371_1212_U151, P3_ADD_371_1212_U150, P3_ADD_371_1212_U43);
  nand ginst19285 (P3_ADD_371_1212_U152, P3_ADD_371_1212_U151, P3_ADD_371_1212_U96);
  nand ginst19286 (P3_ADD_371_1212_U153, P3_ADD_371_1212_U131, P3_ADD_371_1212_U24);
  nand ginst19287 (P3_ADD_371_1212_U154, P3_INSTADDRPOINTER_REG_5__SCAN_IN, P3_ADD_371_U19);
  nand ginst19288 (P3_ADD_371_1212_U155, P3_ADD_371_1212_U153, P3_ADD_371_1212_U97);
  or ginst19289 (P3_ADD_371_1212_U156, P3_INSTADDRPOINTER_REG_4__SCAN_IN, P3_ADD_371_U20);
  or ginst19290 (P3_ADD_371_1212_U157, P3_INSTADDRPOINTER_REG_2__SCAN_IN, P3_ADD_371_U5);
  nand ginst19291 (P3_ADD_371_1212_U158, P3_ADD_371_1212_U157, P3_ADD_371_1212_U44);
  nand ginst19292 (P3_ADD_371_1212_U159, P3_ADD_371_1212_U158, P3_ADD_371_1212_U98);
  and ginst19293 (P3_ADD_371_1212_U16, P3_ADD_371_1212_U178, P3_ADD_371_1212_U73);
  nand ginst19294 (P3_ADD_371_1212_U160, P3_ADD_371_1212_U124, P3_ADD_371_1212_U29);
  nand ginst19295 (P3_ADD_371_1212_U161, P3_INSTADDRPOINTER_REG_3__SCAN_IN, P3_ADD_371_U25);
  nand ginst19296 (P3_ADD_371_1212_U162, P3_ADD_371_1212_U119, P3_ADD_371_1212_U160, P3_ADD_371_1212_U161);
  not ginst19297 (P3_ADD_371_1212_U163, P3_ADD_371_1212_U49);
  not ginst19298 (P3_ADD_371_1212_U164, P3_ADD_371_1212_U78);
  not ginst19299 (P3_ADD_371_1212_U165, P3_ADD_371_1212_U53);
  not ginst19300 (P3_ADD_371_1212_U166, P3_ADD_371_1212_U56);
  not ginst19301 (P3_ADD_371_1212_U167, P3_ADD_371_1212_U59);
  nand ginst19302 (P3_ADD_371_1212_U168, P3_INSTADDRPOINTER_REG_20__SCAN_IN, P3_ADD_371_1212_U167);
  not ginst19303 (P3_ADD_371_1212_U169, P3_ADD_371_1212_U62);
  and ginst19304 (P3_ADD_371_1212_U17, P3_ADD_371_1212_U176, P3_ADD_371_1212_U75);
  not ginst19305 (P3_ADD_371_1212_U170, P3_ADD_371_1212_U65);
  not ginst19306 (P3_ADD_371_1212_U171, P3_ADD_371_1212_U68);
  not ginst19307 (P3_ADD_371_1212_U172, P3_ADD_371_1212_U70);
  not ginst19308 (P3_ADD_371_1212_U173, P3_ADD_371_1212_U73);
  not ginst19309 (P3_ADD_371_1212_U174, P3_ADD_371_1212_U75);
  or ginst19310 (P3_ADD_371_1212_U175, P3_INSTADDRPOINTER_REG_2__SCAN_IN, P3_ADD_371_U5);
  nand ginst19311 (P3_ADD_371_1212_U176, P3_ADD_371_1212_U73, P3_ADD_371_1212_U74);
  nand ginst19312 (P3_ADD_371_1212_U177, P3_INSTADDRPOINTER_REG_27__SCAN_IN, P3_ADD_371_1212_U172);
  nand ginst19313 (P3_ADD_371_1212_U178, P3_ADD_371_1212_U177, P3_ADD_371_1212_U71);
  nand ginst19314 (P3_ADD_371_1212_U179, P3_ADD_371_1212_U68, P3_ADD_371_1212_U69);
  and ginst19315 (P3_ADD_371_1212_U18, P3_ADD_371_1212_U159, P3_ADD_371_1212_U162);
  nand ginst19316 (P3_ADD_371_1212_U180, P3_INSTADDRPOINTER_REG_24__SCAN_IN, P3_ADD_371_1212_U170);
  nand ginst19317 (P3_ADD_371_1212_U181, P3_ADD_371_1212_U180, P3_ADD_371_1212_U66);
  nand ginst19318 (P3_ADD_371_1212_U182, P3_INSTADDRPOINTER_REG_22__SCAN_IN, P3_ADD_371_1212_U169);
  nand ginst19319 (P3_ADD_371_1212_U183, P3_ADD_371_1212_U182, P3_ADD_371_1212_U63);
  nand ginst19320 (P3_ADD_371_1212_U184, P3_ADD_371_1212_U168, P3_ADD_371_1212_U61);
  nand ginst19321 (P3_ADD_371_1212_U185, P3_ADD_371_1212_U59, P3_ADD_371_1212_U60);
  nand ginst19322 (P3_ADD_371_1212_U186, P3_INSTADDRPOINTER_REG_18__SCAN_IN, P3_ADD_371_1212_U166);
  nand ginst19323 (P3_ADD_371_1212_U187, P3_ADD_371_1212_U186, P3_ADD_371_1212_U58);
  nand ginst19324 (P3_ADD_371_1212_U188, P3_INSTADDRPOINTER_REG_16__SCAN_IN, P3_ADD_371_1212_U165);
  nand ginst19325 (P3_ADD_371_1212_U189, P3_ADD_371_1212_U188, P3_ADD_371_1212_U54);
  and ginst19326 (P3_ADD_371_1212_U19, P3_ADD_371_1212_U152, P3_ADD_371_1212_U155);
  nand ginst19327 (P3_ADD_371_1212_U190, P3_INSTADDRPOINTER_REG_14__SCAN_IN, P3_ADD_371_1212_U164);
  nand ginst19328 (P3_ADD_371_1212_U191, P3_ADD_371_1212_U190, P3_ADD_371_1212_U51);
  nand ginst19329 (P3_ADD_371_1212_U192, P3_ADD_371_1212_U49, P3_ADD_371_1212_U50);
  nand ginst19330 (P3_ADD_371_1212_U193, P3_INSTADDRPOINTER_REG_11__SCAN_IN, P3_ADD_371_1212_U117);
  nand ginst19331 (P3_ADD_371_1212_U194, P3_ADD_371_1212_U193, P3_ADD_371_1212_U47);
  nand ginst19332 (P3_ADD_371_1212_U195, P3_INSTADDRPOINTER_REG_9__SCAN_IN, P3_ADD_371_1212_U108);
  nand ginst19333 (P3_ADD_371_1212_U196, P3_ADD_371_1212_U195, P3_ADD_371_1212_U45);
  nand ginst19334 (P3_ADD_371_1212_U197, P3_ADD_371_1212_U156, P3_ADD_371_1212_U24);
  nand ginst19335 (P3_ADD_371_1212_U198, P3_INSTADDRPOINTER_REG_30__SCAN_IN, P3_ADD_371_1212_U174);
  nand ginst19336 (P3_ADD_371_1212_U199, P3_ADD_371_1212_U175, P3_ADD_371_1212_U29);
  nand ginst19337 (P3_ADD_371_1212_U20, P3_ADD_371_1212_U203, P3_ADD_371_1212_U254, P3_ADD_371_1212_U255);
  nand ginst19338 (P3_ADD_371_1212_U200, P3_INSTADDRPOINTER_REG_7__SCAN_IN, P3_ADD_371_U17);
  nand ginst19339 (P3_ADD_371_1212_U201, P3_INSTADDRPOINTER_REG_3__SCAN_IN, P3_ADD_371_1212_U125);
  nand ginst19340 (P3_ADD_371_1212_U202, P3_ADD_371_1212_U125, P3_ADD_371_U25);
  nand ginst19341 (P3_ADD_371_1212_U203, P3_INSTADDRPOINTER_REG_1__SCAN_IN, P3_ADD_371_1212_U120);
  nand ginst19342 (P3_ADD_371_1212_U204, P3_INSTADDRPOINTER_REG_9__SCAN_IN, P3_ADD_371_1212_U108);
  nand ginst19343 (P3_ADD_371_1212_U205, P3_ADD_371_1212_U149, P3_ADD_371_1212_U42);
  nand ginst19344 (P3_ADD_371_1212_U206, P3_INSTADDRPOINTER_REG_8__SCAN_IN, P3_ADD_371_1212_U40);
  nand ginst19345 (P3_ADD_371_1212_U207, P3_ADD_371_1212_U41, P3_ADD_371_U6);
  nand ginst19346 (P3_ADD_371_1212_U208, P3_INSTADDRPOINTER_REG_8__SCAN_IN, P3_ADD_371_1212_U40);
  nand ginst19347 (P3_ADD_371_1212_U209, P3_ADD_371_1212_U41, P3_ADD_371_U6);
  not ginst19348 (P3_ADD_371_1212_U21, P3_ADD_371_U20);
  nand ginst19349 (P3_ADD_371_1212_U210, P3_ADD_371_1212_U208, P3_ADD_371_1212_U209);
  nand ginst19350 (P3_ADD_371_1212_U211, P3_ADD_371_1212_U110, P3_ADD_371_1212_U111);
  nand ginst19351 (P3_ADD_371_1212_U212, P3_ADD_371_1212_U145, P3_ADD_371_1212_U210);
  nand ginst19352 (P3_ADD_371_1212_U213, P3_INSTADDRPOINTER_REG_7__SCAN_IN, P3_ADD_371_1212_U39);
  nand ginst19353 (P3_ADD_371_1212_U214, P3_ADD_371_1212_U38, P3_ADD_371_U17);
  nand ginst19354 (P3_ADD_371_1212_U215, P3_INSTADDRPOINTER_REG_7__SCAN_IN, P3_ADD_371_1212_U39);
  nand ginst19355 (P3_ADD_371_1212_U216, P3_ADD_371_1212_U38, P3_ADD_371_U17);
  nand ginst19356 (P3_ADD_371_1212_U217, P3_ADD_371_1212_U215, P3_ADD_371_1212_U216);
  nand ginst19357 (P3_ADD_371_1212_U218, P3_ADD_371_1212_U112, P3_ADD_371_1212_U113);
  nand ginst19358 (P3_ADD_371_1212_U219, P3_ADD_371_1212_U143, P3_ADD_371_1212_U217);
  not ginst19359 (P3_ADD_371_1212_U22, P3_INSTADDRPOINTER_REG_4__SCAN_IN);
  nand ginst19360 (P3_ADD_371_1212_U220, P3_INSTADDRPOINTER_REG_6__SCAN_IN, P3_ADD_371_1212_U36);
  nand ginst19361 (P3_ADD_371_1212_U221, P3_ADD_371_1212_U37, P3_ADD_371_U18);
  nand ginst19362 (P3_ADD_371_1212_U222, P3_INSTADDRPOINTER_REG_6__SCAN_IN, P3_ADD_371_1212_U36);
  nand ginst19363 (P3_ADD_371_1212_U223, P3_ADD_371_1212_U37, P3_ADD_371_U18);
  nand ginst19364 (P3_ADD_371_1212_U224, P3_ADD_371_1212_U222, P3_ADD_371_1212_U223);
  nand ginst19365 (P3_ADD_371_1212_U225, P3_ADD_371_1212_U114, P3_ADD_371_1212_U115);
  nand ginst19366 (P3_ADD_371_1212_U226, P3_ADD_371_1212_U139, P3_ADD_371_1212_U224);
  nand ginst19367 (P3_ADD_371_1212_U227, P3_INSTADDRPOINTER_REG_5__SCAN_IN, P3_ADD_371_1212_U25);
  nand ginst19368 (P3_ADD_371_1212_U228, P3_ADD_371_1212_U23, P3_ADD_371_U19);
  nand ginst19369 (P3_ADD_371_1212_U229, P3_INSTADDRPOINTER_REG_4__SCAN_IN, P3_ADD_371_1212_U21);
  not ginst19370 (P3_ADD_371_1212_U23, P3_INSTADDRPOINTER_REG_5__SCAN_IN);
  nand ginst19371 (P3_ADD_371_1212_U230, P3_ADD_371_1212_U22, P3_ADD_371_U20);
  nand ginst19372 (P3_ADD_371_1212_U231, P3_ADD_371_1212_U229, P3_ADD_371_1212_U230);
  nand ginst19373 (P3_ADD_371_1212_U232, P3_ADD_371_1212_U197, P3_ADD_371_1212_U43);
  nand ginst19374 (P3_ADD_371_1212_U233, P3_ADD_371_1212_U131, P3_ADD_371_1212_U231);
  nand ginst19375 (P3_ADD_371_1212_U234, P3_INSTADDRPOINTER_REG_3__SCAN_IN, P3_ADD_371_1212_U30);
  nand ginst19376 (P3_ADD_371_1212_U235, P3_ADD_371_1212_U28, P3_ADD_371_U25);
  nand ginst19377 (P3_ADD_371_1212_U236, P3_INSTADDRPOINTER_REG_31__SCAN_IN, P3_ADD_371_1212_U198);
  nand ginst19378 (P3_ADD_371_1212_U237, P3_INSTADDRPOINTER_REG_30__SCAN_IN, P3_ADD_371_1212_U116, P3_ADD_371_1212_U174);
  nand ginst19379 (P3_ADD_371_1212_U238, P3_INSTADDRPOINTER_REG_30__SCAN_IN, P3_ADD_371_1212_U75);
  nand ginst19380 (P3_ADD_371_1212_U239, P3_ADD_371_1212_U174, P3_ADD_371_1212_U76);
  nand ginst19381 (P3_ADD_371_1212_U24, P3_INSTADDRPOINTER_REG_4__SCAN_IN, P3_ADD_371_U20);
  nand ginst19382 (P3_ADD_371_1212_U240, P3_INSTADDRPOINTER_REG_2__SCAN_IN, P3_ADD_371_1212_U26);
  nand ginst19383 (P3_ADD_371_1212_U241, P3_ADD_371_1212_U27, P3_ADD_371_U5);
  nand ginst19384 (P3_ADD_371_1212_U242, P3_ADD_371_1212_U240, P3_ADD_371_1212_U241);
  nand ginst19385 (P3_ADD_371_1212_U243, P3_ADD_371_1212_U199, P3_ADD_371_1212_U44);
  nand ginst19386 (P3_ADD_371_1212_U244, P3_ADD_371_1212_U124, P3_ADD_371_1212_U242);
  nand ginst19387 (P3_ADD_371_1212_U245, P3_INSTADDRPOINTER_REG_27__SCAN_IN, P3_ADD_371_1212_U70);
  nand ginst19388 (P3_ADD_371_1212_U246, P3_ADD_371_1212_U172, P3_ADD_371_1212_U72);
  nand ginst19389 (P3_ADD_371_1212_U247, P3_INSTADDRPOINTER_REG_24__SCAN_IN, P3_ADD_371_1212_U65);
  nand ginst19390 (P3_ADD_371_1212_U248, P3_ADD_371_1212_U170, P3_ADD_371_1212_U67);
  nand ginst19391 (P3_ADD_371_1212_U249, P3_INSTADDRPOINTER_REG_22__SCAN_IN, P3_ADD_371_1212_U62);
  not ginst19392 (P3_ADD_371_1212_U25, P3_ADD_371_U19);
  nand ginst19393 (P3_ADD_371_1212_U250, P3_ADD_371_1212_U169, P3_ADD_371_1212_U64);
  nand ginst19394 (P3_ADD_371_1212_U251, P3_INSTADDRPOINTER_REG_1__SCAN_IN, P3_ADD_371_1212_U34);
  nand ginst19395 (P3_ADD_371_1212_U252, P3_ADD_371_1212_U121, P3_ADD_371_1212_U33);
  nand ginst19396 (P3_ADD_371_1212_U253, P3_ADD_371_1212_U251, P3_ADD_371_1212_U252);
  nand ginst19397 (P3_ADD_371_1212_U254, P3_ADD_371_1212_U33, P3_ADD_371_1212_U34, P3_ADD_371_U21);
  nand ginst19398 (P3_ADD_371_1212_U255, P3_ADD_371_1212_U253, P3_ADD_371_1212_U35);
  nand ginst19399 (P3_ADD_371_1212_U256, P3_INSTADDRPOINTER_REG_18__SCAN_IN, P3_ADD_371_1212_U56);
  nand ginst19400 (P3_ADD_371_1212_U257, P3_ADD_371_1212_U166, P3_ADD_371_1212_U57);
  nand ginst19401 (P3_ADD_371_1212_U258, P3_INSTADDRPOINTER_REG_16__SCAN_IN, P3_ADD_371_1212_U53);
  nand ginst19402 (P3_ADD_371_1212_U259, P3_ADD_371_1212_U165, P3_ADD_371_1212_U55);
  not ginst19403 (P3_ADD_371_1212_U26, P3_ADD_371_U5);
  nand ginst19404 (P3_ADD_371_1212_U260, P3_INSTADDRPOINTER_REG_14__SCAN_IN, P3_ADD_371_1212_U78);
  nand ginst19405 (P3_ADD_371_1212_U261, P3_ADD_371_1212_U164, P3_ADD_371_1212_U52);
  nand ginst19406 (P3_ADD_371_1212_U262, P3_ADD_371_1212_U117, P3_ADD_371_1212_U46);
  nand ginst19407 (P3_ADD_371_1212_U263, P3_INSTADDRPOINTER_REG_11__SCAN_IN, P3_ADD_371_1212_U48);
  nand ginst19408 (P3_ADD_371_1212_U264, P3_INSTADDRPOINTER_REG_0__SCAN_IN, P3_ADD_371_1212_U31);
  nand ginst19409 (P3_ADD_371_1212_U265, P3_ADD_371_1212_U32, P3_ADD_371_U4);
  not ginst19410 (P3_ADD_371_1212_U27, P3_INSTADDRPOINTER_REG_2__SCAN_IN);
  not ginst19411 (P3_ADD_371_1212_U28, P3_INSTADDRPOINTER_REG_3__SCAN_IN);
  nand ginst19412 (P3_ADD_371_1212_U29, P3_INSTADDRPOINTER_REG_2__SCAN_IN, P3_ADD_371_U5);
  not ginst19413 (P3_ADD_371_1212_U30, P3_ADD_371_U25);
  not ginst19414 (P3_ADD_371_1212_U31, P3_ADD_371_U4);
  not ginst19415 (P3_ADD_371_1212_U32, P3_INSTADDRPOINTER_REG_0__SCAN_IN);
  not ginst19416 (P3_ADD_371_1212_U33, P3_INSTADDRPOINTER_REG_1__SCAN_IN);
  nand ginst19417 (P3_ADD_371_1212_U34, P3_INSTADDRPOINTER_REG_0__SCAN_IN, P3_ADD_371_U4);
  not ginst19418 (P3_ADD_371_1212_U35, P3_ADD_371_U21);
  not ginst19419 (P3_ADD_371_1212_U36, P3_ADD_371_U18);
  not ginst19420 (P3_ADD_371_1212_U37, P3_INSTADDRPOINTER_REG_6__SCAN_IN);
  not ginst19421 (P3_ADD_371_1212_U38, P3_INSTADDRPOINTER_REG_7__SCAN_IN);
  not ginst19422 (P3_ADD_371_1212_U39, P3_ADD_371_U17);
  and ginst19423 (P3_ADD_371_1212_U4, P3_ADD_371_1212_U132, P3_ADD_371_1212_U133);
  not ginst19424 (P3_ADD_371_1212_U40, P3_ADD_371_U6);
  not ginst19425 (P3_ADD_371_1212_U41, P3_INSTADDRPOINTER_REG_8__SCAN_IN);
  not ginst19426 (P3_ADD_371_1212_U42, P3_INSTADDRPOINTER_REG_9__SCAN_IN);
  nand ginst19427 (P3_ADD_371_1212_U43, P3_ADD_371_1212_U130, P3_ADD_371_1212_U94);
  nand ginst19428 (P3_ADD_371_1212_U44, P3_ADD_371_1212_U123, P3_ADD_371_1212_U77);
  not ginst19429 (P3_ADD_371_1212_U45, P3_INSTADDRPOINTER_REG_10__SCAN_IN);
  not ginst19430 (P3_ADD_371_1212_U46, P3_INSTADDRPOINTER_REG_11__SCAN_IN);
  not ginst19431 (P3_ADD_371_1212_U47, P3_INSTADDRPOINTER_REG_12__SCAN_IN);
  nand ginst19432 (P3_ADD_371_1212_U48, P3_ADD_371_1212_U108, P3_ADD_371_1212_U99);
  nand ginst19433 (P3_ADD_371_1212_U49, P3_ADD_371_1212_U100, P3_ADD_371_1212_U117);
  and ginst19434 (P3_ADD_371_1212_U5, P3_ADD_371_1212_U196, P3_ADD_371_1212_U48);
  not ginst19435 (P3_ADD_371_1212_U50, P3_INSTADDRPOINTER_REG_13__SCAN_IN);
  not ginst19436 (P3_ADD_371_1212_U51, P3_INSTADDRPOINTER_REG_15__SCAN_IN);
  not ginst19437 (P3_ADD_371_1212_U52, P3_INSTADDRPOINTER_REG_14__SCAN_IN);
  nand ginst19438 (P3_ADD_371_1212_U53, P3_ADD_371_1212_U101, P3_ADD_371_1212_U163);
  not ginst19439 (P3_ADD_371_1212_U54, P3_INSTADDRPOINTER_REG_17__SCAN_IN);
  not ginst19440 (P3_ADD_371_1212_U55, P3_INSTADDRPOINTER_REG_16__SCAN_IN);
  nand ginst19441 (P3_ADD_371_1212_U56, P3_ADD_371_1212_U102, P3_ADD_371_1212_U165);
  not ginst19442 (P3_ADD_371_1212_U57, P3_INSTADDRPOINTER_REG_18__SCAN_IN);
  not ginst19443 (P3_ADD_371_1212_U58, P3_INSTADDRPOINTER_REG_19__SCAN_IN);
  nand ginst19444 (P3_ADD_371_1212_U59, P3_ADD_371_1212_U103, P3_ADD_371_1212_U166);
  and ginst19445 (P3_ADD_371_1212_U6, P3_ADD_371_1212_U194, P3_ADD_371_1212_U49);
  not ginst19446 (P3_ADD_371_1212_U60, P3_INSTADDRPOINTER_REG_20__SCAN_IN);
  not ginst19447 (P3_ADD_371_1212_U61, P3_INSTADDRPOINTER_REG_21__SCAN_IN);
  nand ginst19448 (P3_ADD_371_1212_U62, P3_ADD_371_1212_U104, P3_ADD_371_1212_U167);
  not ginst19449 (P3_ADD_371_1212_U63, P3_INSTADDRPOINTER_REG_23__SCAN_IN);
  not ginst19450 (P3_ADD_371_1212_U64, P3_INSTADDRPOINTER_REG_22__SCAN_IN);
  nand ginst19451 (P3_ADD_371_1212_U65, P3_ADD_371_1212_U105, P3_ADD_371_1212_U169);
  not ginst19452 (P3_ADD_371_1212_U66, P3_INSTADDRPOINTER_REG_25__SCAN_IN);
  not ginst19453 (P3_ADD_371_1212_U67, P3_INSTADDRPOINTER_REG_24__SCAN_IN);
  nand ginst19454 (P3_ADD_371_1212_U68, P3_ADD_371_1212_U106, P3_ADD_371_1212_U170);
  not ginst19455 (P3_ADD_371_1212_U69, P3_INSTADDRPOINTER_REG_26__SCAN_IN);
  and ginst19456 (P3_ADD_371_1212_U7, P3_ADD_371_1212_U192, P3_ADD_371_1212_U78);
  nand ginst19457 (P3_ADD_371_1212_U70, P3_INSTADDRPOINTER_REG_26__SCAN_IN, P3_ADD_371_1212_U171);
  not ginst19458 (P3_ADD_371_1212_U71, P3_INSTADDRPOINTER_REG_28__SCAN_IN);
  not ginst19459 (P3_ADD_371_1212_U72, P3_INSTADDRPOINTER_REG_27__SCAN_IN);
  nand ginst19460 (P3_ADD_371_1212_U73, P3_ADD_371_1212_U107, P3_ADD_371_1212_U172);
  not ginst19461 (P3_ADD_371_1212_U74, P3_INSTADDRPOINTER_REG_29__SCAN_IN);
  nand ginst19462 (P3_ADD_371_1212_U75, P3_INSTADDRPOINTER_REG_29__SCAN_IN, P3_ADD_371_1212_U173);
  not ginst19463 (P3_ADD_371_1212_U76, P3_INSTADDRPOINTER_REG_30__SCAN_IN);
  nand ginst19464 (P3_ADD_371_1212_U77, P3_ADD_371_1212_U121, P3_ADD_371_U21);
  nand ginst19465 (P3_ADD_371_1212_U78, P3_INSTADDRPOINTER_REG_13__SCAN_IN, P3_ADD_371_1212_U163);
  nand ginst19466 (P3_ADD_371_1212_U79, P3_ADD_371_1212_U238, P3_ADD_371_1212_U239);
  and ginst19467 (P3_ADD_371_1212_U8, P3_ADD_371_1212_U191, P3_ADD_371_1212_U53);
  nand ginst19468 (P3_ADD_371_1212_U80, P3_ADD_371_1212_U245, P3_ADD_371_1212_U246);
  nand ginst19469 (P3_ADD_371_1212_U81, P3_ADD_371_1212_U247, P3_ADD_371_1212_U248);
  nand ginst19470 (P3_ADD_371_1212_U82, P3_ADD_371_1212_U249, P3_ADD_371_1212_U250);
  nand ginst19471 (P3_ADD_371_1212_U83, P3_ADD_371_1212_U256, P3_ADD_371_1212_U257);
  nand ginst19472 (P3_ADD_371_1212_U84, P3_ADD_371_1212_U258, P3_ADD_371_1212_U259);
  nand ginst19473 (P3_ADD_371_1212_U85, P3_ADD_371_1212_U260, P3_ADD_371_1212_U261);
  nand ginst19474 (P3_ADD_371_1212_U86, P3_ADD_371_1212_U262, P3_ADD_371_1212_U263);
  nand ginst19475 (P3_ADD_371_1212_U87, P3_ADD_371_1212_U264, P3_ADD_371_1212_U265);
  nand ginst19476 (P3_ADD_371_1212_U88, P3_ADD_371_1212_U211, P3_ADD_371_1212_U212);
  nand ginst19477 (P3_ADD_371_1212_U89, P3_ADD_371_1212_U218, P3_ADD_371_1212_U219);
  and ginst19478 (P3_ADD_371_1212_U9, P3_ADD_371_1212_U189, P3_ADD_371_1212_U56);
  nand ginst19479 (P3_ADD_371_1212_U90, P3_ADD_371_1212_U225, P3_ADD_371_1212_U226);
  nand ginst19480 (P3_ADD_371_1212_U91, P3_ADD_371_1212_U232, P3_ADD_371_1212_U233);
  nand ginst19481 (P3_ADD_371_1212_U92, P3_ADD_371_1212_U236, P3_ADD_371_1212_U237);
  nand ginst19482 (P3_ADD_371_1212_U93, P3_ADD_371_1212_U243, P3_ADD_371_1212_U244);
  and ginst19483 (P3_ADD_371_1212_U94, P3_ADD_371_1212_U128, P3_ADD_371_1212_U129);
  and ginst19484 (P3_ADD_371_1212_U95, P3_ADD_371_1212_U136, P3_ADD_371_1212_U137);
  and ginst19485 (P3_ADD_371_1212_U96, P3_ADD_371_1212_U227, P3_ADD_371_1212_U228, P3_ADD_371_1212_U24);
  and ginst19486 (P3_ADD_371_1212_U97, P3_ADD_371_1212_U154, P3_ADD_371_1212_U4);
  and ginst19487 (P3_ADD_371_1212_U98, P3_ADD_371_1212_U234, P3_ADD_371_1212_U235, P3_ADD_371_1212_U29);
  and ginst19488 (P3_ADD_371_1212_U99, P3_INSTADDRPOINTER_REG_9__SCAN_IN, P3_INSTADDRPOINTER_REG_10__SCAN_IN);
  not ginst19489 (P3_ADD_371_U10, P3_U2625);
  nand ginst19490 (P3_ADD_371_U11, P3_ADD_371_U28, P3_U2625);
  not ginst19491 (P3_ADD_371_U12, P3_U2626);
  nand ginst19492 (P3_ADD_371_U13, P3_ADD_371_U29, P3_U2626);
  not ginst19493 (P3_ADD_371_U14, P3_U2628);
  not ginst19494 (P3_ADD_371_U15, P3_U2627);
  not ginst19495 (P3_ADD_371_U16, P3_U2623);
  nand ginst19496 (P3_ADD_371_U17, P3_ADD_371_U33, P3_ADD_371_U34);
  nand ginst19497 (P3_ADD_371_U18, P3_ADD_371_U35, P3_ADD_371_U36);
  nand ginst19498 (P3_ADD_371_U19, P3_ADD_371_U37, P3_ADD_371_U38);
  nand ginst19499 (P3_ADD_371_U20, P3_ADD_371_U39, P3_ADD_371_U40);
  nand ginst19500 (P3_ADD_371_U21, P3_ADD_371_U43, P3_ADD_371_U44);
  and ginst19501 (P3_ADD_371_U22, P3_U2627, P3_U2628);
  nand ginst19502 (P3_ADD_371_U23, P3_ADD_371_U30, P3_U2627);
  nand ginst19503 (P3_ADD_371_U24, P3_ADD_371_U16, P3_ADD_371_U26);
  and ginst19504 (P3_ADD_371_U25, P3_ADD_371_U41, P3_ADD_371_U42);
  nand ginst19505 (P3_ADD_371_U26, P3_U2621, P3_U2622);
  not ginst19506 (P3_ADD_371_U27, P3_ADD_371_U24);
  not ginst19507 (P3_ADD_371_U28, P3_ADD_371_U9);
  not ginst19508 (P3_ADD_371_U29, P3_ADD_371_U11);
  not ginst19509 (P3_ADD_371_U30, P3_ADD_371_U13);
  not ginst19510 (P3_ADD_371_U31, P3_ADD_371_U23);
  nand ginst19511 (P3_ADD_371_U32, P3_U2621, P3_U2622, P3_U2623);
  nand ginst19512 (P3_ADD_371_U33, P3_ADD_371_U23, P3_U2628);
  nand ginst19513 (P3_ADD_371_U34, P3_ADD_371_U14, P3_ADD_371_U31);
  nand ginst19514 (P3_ADD_371_U35, P3_ADD_371_U13, P3_U2627);
  nand ginst19515 (P3_ADD_371_U36, P3_ADD_371_U15, P3_ADD_371_U30);
  nand ginst19516 (P3_ADD_371_U37, P3_ADD_371_U11, P3_U2626);
  nand ginst19517 (P3_ADD_371_U38, P3_ADD_371_U12, P3_ADD_371_U29);
  nand ginst19518 (P3_ADD_371_U39, P3_ADD_371_U9, P3_U2625);
  not ginst19519 (P3_ADD_371_U4, P3_U2621);
  nand ginst19520 (P3_ADD_371_U40, P3_ADD_371_U10, P3_ADD_371_U28);
  nand ginst19521 (P3_ADD_371_U41, P3_ADD_371_U24, P3_U2624);
  nand ginst19522 (P3_ADD_371_U42, P3_ADD_371_U27, P3_ADD_371_U8);
  nand ginst19523 (P3_ADD_371_U43, P3_ADD_371_U4, P3_U2622);
  nand ginst19524 (P3_ADD_371_U44, P3_ADD_371_U7, P3_U2621);
  nand ginst19525 (P3_ADD_371_U5, P3_ADD_371_U24, P3_ADD_371_U32);
  and ginst19526 (P3_ADD_371_U6, P3_ADD_371_U22, P3_ADD_371_U30);
  not ginst19527 (P3_ADD_371_U7, P3_U2622);
  not ginst19528 (P3_ADD_371_U8, P3_U2624);
  nand ginst19529 (P3_ADD_371_U9, P3_ADD_371_U24, P3_U2624);
  not ginst19530 (P3_ADD_380_U10, P3_INSTADDRPOINTER_REG_3__SCAN_IN);
  not ginst19531 (P3_ADD_380_U100, P3_ADD_380_U11);
  not ginst19532 (P3_ADD_380_U101, P3_ADD_380_U13);
  not ginst19533 (P3_ADD_380_U102, P3_ADD_380_U15);
  not ginst19534 (P3_ADD_380_U103, P3_ADD_380_U17);
  not ginst19535 (P3_ADD_380_U104, P3_ADD_380_U19);
  not ginst19536 (P3_ADD_380_U105, P3_ADD_380_U22);
  not ginst19537 (P3_ADD_380_U106, P3_ADD_380_U23);
  not ginst19538 (P3_ADD_380_U107, P3_ADD_380_U25);
  not ginst19539 (P3_ADD_380_U108, P3_ADD_380_U27);
  not ginst19540 (P3_ADD_380_U109, P3_ADD_380_U29);
  nand ginst19541 (P3_ADD_380_U11, P3_INSTADDRPOINTER_REG_3__SCAN_IN, P3_ADD_380_U99);
  not ginst19542 (P3_ADD_380_U110, P3_ADD_380_U31);
  not ginst19543 (P3_ADD_380_U111, P3_ADD_380_U33);
  not ginst19544 (P3_ADD_380_U112, P3_ADD_380_U35);
  not ginst19545 (P3_ADD_380_U113, P3_ADD_380_U37);
  not ginst19546 (P3_ADD_380_U114, P3_ADD_380_U39);
  not ginst19547 (P3_ADD_380_U115, P3_ADD_380_U41);
  not ginst19548 (P3_ADD_380_U116, P3_ADD_380_U43);
  not ginst19549 (P3_ADD_380_U117, P3_ADD_380_U45);
  not ginst19550 (P3_ADD_380_U118, P3_ADD_380_U47);
  not ginst19551 (P3_ADD_380_U119, P3_ADD_380_U49);
  not ginst19552 (P3_ADD_380_U12, P3_INSTADDRPOINTER_REG_4__SCAN_IN);
  not ginst19553 (P3_ADD_380_U120, P3_ADD_380_U51);
  not ginst19554 (P3_ADD_380_U121, P3_ADD_380_U53);
  not ginst19555 (P3_ADD_380_U122, P3_ADD_380_U55);
  not ginst19556 (P3_ADD_380_U123, P3_ADD_380_U57);
  not ginst19557 (P3_ADD_380_U124, P3_ADD_380_U59);
  not ginst19558 (P3_ADD_380_U125, P3_ADD_380_U61);
  not ginst19559 (P3_ADD_380_U126, P3_ADD_380_U63);
  not ginst19560 (P3_ADD_380_U127, P3_ADD_380_U97);
  nand ginst19561 (P3_ADD_380_U128, P3_INSTADDRPOINTER_REG_9__SCAN_IN, P3_ADD_380_U22);
  nand ginst19562 (P3_ADD_380_U129, P3_ADD_380_U105, P3_ADD_380_U21);
  nand ginst19563 (P3_ADD_380_U13, P3_INSTADDRPOINTER_REG_4__SCAN_IN, P3_ADD_380_U100);
  nand ginst19564 (P3_ADD_380_U130, P3_INSTADDRPOINTER_REG_8__SCAN_IN, P3_ADD_380_U19);
  nand ginst19565 (P3_ADD_380_U131, P3_ADD_380_U104, P3_ADD_380_U20);
  nand ginst19566 (P3_ADD_380_U132, P3_INSTADDRPOINTER_REG_7__SCAN_IN, P3_ADD_380_U17);
  nand ginst19567 (P3_ADD_380_U133, P3_ADD_380_U103, P3_ADD_380_U18);
  nand ginst19568 (P3_ADD_380_U134, P3_INSTADDRPOINTER_REG_6__SCAN_IN, P3_ADD_380_U15);
  nand ginst19569 (P3_ADD_380_U135, P3_ADD_380_U102, P3_ADD_380_U16);
  nand ginst19570 (P3_ADD_380_U136, P3_INSTADDRPOINTER_REG_5__SCAN_IN, P3_ADD_380_U13);
  nand ginst19571 (P3_ADD_380_U137, P3_ADD_380_U101, P3_ADD_380_U14);
  nand ginst19572 (P3_ADD_380_U138, P3_INSTADDRPOINTER_REG_4__SCAN_IN, P3_ADD_380_U11);
  nand ginst19573 (P3_ADD_380_U139, P3_ADD_380_U100, P3_ADD_380_U12);
  not ginst19574 (P3_ADD_380_U14, P3_INSTADDRPOINTER_REG_5__SCAN_IN);
  nand ginst19575 (P3_ADD_380_U140, P3_INSTADDRPOINTER_REG_3__SCAN_IN, P3_ADD_380_U9);
  nand ginst19576 (P3_ADD_380_U141, P3_ADD_380_U10, P3_ADD_380_U99);
  nand ginst19577 (P3_ADD_380_U142, P3_INSTADDRPOINTER_REG_31__SCAN_IN, P3_ADD_380_U97);
  nand ginst19578 (P3_ADD_380_U143, P3_ADD_380_U127, P3_ADD_380_U96);
  nand ginst19579 (P3_ADD_380_U144, P3_INSTADDRPOINTER_REG_30__SCAN_IN, P3_ADD_380_U63);
  nand ginst19580 (P3_ADD_380_U145, P3_ADD_380_U126, P3_ADD_380_U64);
  nand ginst19581 (P3_ADD_380_U146, P3_INSTADDRPOINTER_REG_2__SCAN_IN, P3_ADD_380_U7);
  nand ginst19582 (P3_ADD_380_U147, P3_ADD_380_U8, P3_ADD_380_U98);
  nand ginst19583 (P3_ADD_380_U148, P3_INSTADDRPOINTER_REG_29__SCAN_IN, P3_ADD_380_U61);
  nand ginst19584 (P3_ADD_380_U149, P3_ADD_380_U125, P3_ADD_380_U62);
  nand ginst19585 (P3_ADD_380_U15, P3_INSTADDRPOINTER_REG_5__SCAN_IN, P3_ADD_380_U101);
  nand ginst19586 (P3_ADD_380_U150, P3_INSTADDRPOINTER_REG_28__SCAN_IN, P3_ADD_380_U59);
  nand ginst19587 (P3_ADD_380_U151, P3_ADD_380_U124, P3_ADD_380_U60);
  nand ginst19588 (P3_ADD_380_U152, P3_INSTADDRPOINTER_REG_27__SCAN_IN, P3_ADD_380_U57);
  nand ginst19589 (P3_ADD_380_U153, P3_ADD_380_U123, P3_ADD_380_U58);
  nand ginst19590 (P3_ADD_380_U154, P3_INSTADDRPOINTER_REG_26__SCAN_IN, P3_ADD_380_U55);
  nand ginst19591 (P3_ADD_380_U155, P3_ADD_380_U122, P3_ADD_380_U56);
  nand ginst19592 (P3_ADD_380_U156, P3_INSTADDRPOINTER_REG_25__SCAN_IN, P3_ADD_380_U53);
  nand ginst19593 (P3_ADD_380_U157, P3_ADD_380_U121, P3_ADD_380_U54);
  nand ginst19594 (P3_ADD_380_U158, P3_INSTADDRPOINTER_REG_24__SCAN_IN, P3_ADD_380_U51);
  nand ginst19595 (P3_ADD_380_U159, P3_ADD_380_U120, P3_ADD_380_U52);
  not ginst19596 (P3_ADD_380_U16, P3_INSTADDRPOINTER_REG_6__SCAN_IN);
  nand ginst19597 (P3_ADD_380_U160, P3_INSTADDRPOINTER_REG_23__SCAN_IN, P3_ADD_380_U49);
  nand ginst19598 (P3_ADD_380_U161, P3_ADD_380_U119, P3_ADD_380_U50);
  nand ginst19599 (P3_ADD_380_U162, P3_INSTADDRPOINTER_REG_22__SCAN_IN, P3_ADD_380_U47);
  nand ginst19600 (P3_ADD_380_U163, P3_ADD_380_U118, P3_ADD_380_U48);
  nand ginst19601 (P3_ADD_380_U164, P3_INSTADDRPOINTER_REG_21__SCAN_IN, P3_ADD_380_U45);
  nand ginst19602 (P3_ADD_380_U165, P3_ADD_380_U117, P3_ADD_380_U46);
  nand ginst19603 (P3_ADD_380_U166, P3_INSTADDRPOINTER_REG_20__SCAN_IN, P3_ADD_380_U43);
  nand ginst19604 (P3_ADD_380_U167, P3_ADD_380_U116, P3_ADD_380_U44);
  nand ginst19605 (P3_ADD_380_U168, P3_INSTADDRPOINTER_REG_1__SCAN_IN, P3_ADD_380_U5);
  nand ginst19606 (P3_ADD_380_U169, P3_INSTADDRPOINTER_REG_0__SCAN_IN, P3_ADD_380_U6);
  nand ginst19607 (P3_ADD_380_U17, P3_INSTADDRPOINTER_REG_6__SCAN_IN, P3_ADD_380_U102);
  nand ginst19608 (P3_ADD_380_U170, P3_INSTADDRPOINTER_REG_19__SCAN_IN, P3_ADD_380_U41);
  nand ginst19609 (P3_ADD_380_U171, P3_ADD_380_U115, P3_ADD_380_U42);
  nand ginst19610 (P3_ADD_380_U172, P3_INSTADDRPOINTER_REG_18__SCAN_IN, P3_ADD_380_U39);
  nand ginst19611 (P3_ADD_380_U173, P3_ADD_380_U114, P3_ADD_380_U40);
  nand ginst19612 (P3_ADD_380_U174, P3_INSTADDRPOINTER_REG_17__SCAN_IN, P3_ADD_380_U37);
  nand ginst19613 (P3_ADD_380_U175, P3_ADD_380_U113, P3_ADD_380_U38);
  nand ginst19614 (P3_ADD_380_U176, P3_INSTADDRPOINTER_REG_16__SCAN_IN, P3_ADD_380_U35);
  nand ginst19615 (P3_ADD_380_U177, P3_ADD_380_U112, P3_ADD_380_U36);
  nand ginst19616 (P3_ADD_380_U178, P3_INSTADDRPOINTER_REG_15__SCAN_IN, P3_ADD_380_U33);
  nand ginst19617 (P3_ADD_380_U179, P3_ADD_380_U111, P3_ADD_380_U34);
  not ginst19618 (P3_ADD_380_U18, P3_INSTADDRPOINTER_REG_7__SCAN_IN);
  nand ginst19619 (P3_ADD_380_U180, P3_INSTADDRPOINTER_REG_14__SCAN_IN, P3_ADD_380_U31);
  nand ginst19620 (P3_ADD_380_U181, P3_ADD_380_U110, P3_ADD_380_U32);
  nand ginst19621 (P3_ADD_380_U182, P3_INSTADDRPOINTER_REG_13__SCAN_IN, P3_ADD_380_U29);
  nand ginst19622 (P3_ADD_380_U183, P3_ADD_380_U109, P3_ADD_380_U30);
  nand ginst19623 (P3_ADD_380_U184, P3_INSTADDRPOINTER_REG_12__SCAN_IN, P3_ADD_380_U27);
  nand ginst19624 (P3_ADD_380_U185, P3_ADD_380_U108, P3_ADD_380_U28);
  nand ginst19625 (P3_ADD_380_U186, P3_INSTADDRPOINTER_REG_11__SCAN_IN, P3_ADD_380_U25);
  nand ginst19626 (P3_ADD_380_U187, P3_ADD_380_U107, P3_ADD_380_U26);
  nand ginst19627 (P3_ADD_380_U188, P3_INSTADDRPOINTER_REG_10__SCAN_IN, P3_ADD_380_U23);
  nand ginst19628 (P3_ADD_380_U189, P3_ADD_380_U106, P3_ADD_380_U24);
  nand ginst19629 (P3_ADD_380_U19, P3_INSTADDRPOINTER_REG_7__SCAN_IN, P3_ADD_380_U103);
  not ginst19630 (P3_ADD_380_U20, P3_INSTADDRPOINTER_REG_8__SCAN_IN);
  not ginst19631 (P3_ADD_380_U21, P3_INSTADDRPOINTER_REG_9__SCAN_IN);
  nand ginst19632 (P3_ADD_380_U22, P3_INSTADDRPOINTER_REG_8__SCAN_IN, P3_ADD_380_U104);
  nand ginst19633 (P3_ADD_380_U23, P3_INSTADDRPOINTER_REG_9__SCAN_IN, P3_ADD_380_U105);
  not ginst19634 (P3_ADD_380_U24, P3_INSTADDRPOINTER_REG_10__SCAN_IN);
  nand ginst19635 (P3_ADD_380_U25, P3_INSTADDRPOINTER_REG_10__SCAN_IN, P3_ADD_380_U106);
  not ginst19636 (P3_ADD_380_U26, P3_INSTADDRPOINTER_REG_11__SCAN_IN);
  nand ginst19637 (P3_ADD_380_U27, P3_INSTADDRPOINTER_REG_11__SCAN_IN, P3_ADD_380_U107);
  not ginst19638 (P3_ADD_380_U28, P3_INSTADDRPOINTER_REG_12__SCAN_IN);
  nand ginst19639 (P3_ADD_380_U29, P3_INSTADDRPOINTER_REG_12__SCAN_IN, P3_ADD_380_U108);
  not ginst19640 (P3_ADD_380_U30, P3_INSTADDRPOINTER_REG_13__SCAN_IN);
  nand ginst19641 (P3_ADD_380_U31, P3_INSTADDRPOINTER_REG_13__SCAN_IN, P3_ADD_380_U109);
  not ginst19642 (P3_ADD_380_U32, P3_INSTADDRPOINTER_REG_14__SCAN_IN);
  nand ginst19643 (P3_ADD_380_U33, P3_INSTADDRPOINTER_REG_14__SCAN_IN, P3_ADD_380_U110);
  not ginst19644 (P3_ADD_380_U34, P3_INSTADDRPOINTER_REG_15__SCAN_IN);
  nand ginst19645 (P3_ADD_380_U35, P3_INSTADDRPOINTER_REG_15__SCAN_IN, P3_ADD_380_U111);
  not ginst19646 (P3_ADD_380_U36, P3_INSTADDRPOINTER_REG_16__SCAN_IN);
  nand ginst19647 (P3_ADD_380_U37, P3_INSTADDRPOINTER_REG_16__SCAN_IN, P3_ADD_380_U112);
  not ginst19648 (P3_ADD_380_U38, P3_INSTADDRPOINTER_REG_17__SCAN_IN);
  nand ginst19649 (P3_ADD_380_U39, P3_INSTADDRPOINTER_REG_17__SCAN_IN, P3_ADD_380_U113);
  not ginst19650 (P3_ADD_380_U40, P3_INSTADDRPOINTER_REG_18__SCAN_IN);
  nand ginst19651 (P3_ADD_380_U41, P3_INSTADDRPOINTER_REG_18__SCAN_IN, P3_ADD_380_U114);
  not ginst19652 (P3_ADD_380_U42, P3_INSTADDRPOINTER_REG_19__SCAN_IN);
  nand ginst19653 (P3_ADD_380_U43, P3_INSTADDRPOINTER_REG_19__SCAN_IN, P3_ADD_380_U115);
  not ginst19654 (P3_ADD_380_U44, P3_INSTADDRPOINTER_REG_20__SCAN_IN);
  nand ginst19655 (P3_ADD_380_U45, P3_INSTADDRPOINTER_REG_20__SCAN_IN, P3_ADD_380_U116);
  not ginst19656 (P3_ADD_380_U46, P3_INSTADDRPOINTER_REG_21__SCAN_IN);
  nand ginst19657 (P3_ADD_380_U47, P3_INSTADDRPOINTER_REG_21__SCAN_IN, P3_ADD_380_U117);
  not ginst19658 (P3_ADD_380_U48, P3_INSTADDRPOINTER_REG_22__SCAN_IN);
  nand ginst19659 (P3_ADD_380_U49, P3_INSTADDRPOINTER_REG_22__SCAN_IN, P3_ADD_380_U118);
  not ginst19660 (P3_ADD_380_U5, P3_INSTADDRPOINTER_REG_0__SCAN_IN);
  not ginst19661 (P3_ADD_380_U50, P3_INSTADDRPOINTER_REG_23__SCAN_IN);
  nand ginst19662 (P3_ADD_380_U51, P3_INSTADDRPOINTER_REG_23__SCAN_IN, P3_ADD_380_U119);
  not ginst19663 (P3_ADD_380_U52, P3_INSTADDRPOINTER_REG_24__SCAN_IN);
  nand ginst19664 (P3_ADD_380_U53, P3_INSTADDRPOINTER_REG_24__SCAN_IN, P3_ADD_380_U120);
  not ginst19665 (P3_ADD_380_U54, P3_INSTADDRPOINTER_REG_25__SCAN_IN);
  nand ginst19666 (P3_ADD_380_U55, P3_INSTADDRPOINTER_REG_25__SCAN_IN, P3_ADD_380_U121);
  not ginst19667 (P3_ADD_380_U56, P3_INSTADDRPOINTER_REG_26__SCAN_IN);
  nand ginst19668 (P3_ADD_380_U57, P3_INSTADDRPOINTER_REG_26__SCAN_IN, P3_ADD_380_U122);
  not ginst19669 (P3_ADD_380_U58, P3_INSTADDRPOINTER_REG_27__SCAN_IN);
  nand ginst19670 (P3_ADD_380_U59, P3_INSTADDRPOINTER_REG_27__SCAN_IN, P3_ADD_380_U123);
  not ginst19671 (P3_ADD_380_U6, P3_INSTADDRPOINTER_REG_1__SCAN_IN);
  not ginst19672 (P3_ADD_380_U60, P3_INSTADDRPOINTER_REG_28__SCAN_IN);
  nand ginst19673 (P3_ADD_380_U61, P3_INSTADDRPOINTER_REG_28__SCAN_IN, P3_ADD_380_U124);
  not ginst19674 (P3_ADD_380_U62, P3_INSTADDRPOINTER_REG_29__SCAN_IN);
  nand ginst19675 (P3_ADD_380_U63, P3_INSTADDRPOINTER_REG_29__SCAN_IN, P3_ADD_380_U125);
  not ginst19676 (P3_ADD_380_U64, P3_INSTADDRPOINTER_REG_30__SCAN_IN);
  nand ginst19677 (P3_ADD_380_U65, P3_ADD_380_U128, P3_ADD_380_U129);
  nand ginst19678 (P3_ADD_380_U66, P3_ADD_380_U130, P3_ADD_380_U131);
  nand ginst19679 (P3_ADD_380_U67, P3_ADD_380_U132, P3_ADD_380_U133);
  nand ginst19680 (P3_ADD_380_U68, P3_ADD_380_U134, P3_ADD_380_U135);
  nand ginst19681 (P3_ADD_380_U69, P3_ADD_380_U136, P3_ADD_380_U137);
  nand ginst19682 (P3_ADD_380_U7, P3_INSTADDRPOINTER_REG_0__SCAN_IN, P3_INSTADDRPOINTER_REG_1__SCAN_IN);
  nand ginst19683 (P3_ADD_380_U70, P3_ADD_380_U138, P3_ADD_380_U139);
  nand ginst19684 (P3_ADD_380_U71, P3_ADD_380_U140, P3_ADD_380_U141);
  nand ginst19685 (P3_ADD_380_U72, P3_ADD_380_U142, P3_ADD_380_U143);
  nand ginst19686 (P3_ADD_380_U73, P3_ADD_380_U144, P3_ADD_380_U145);
  nand ginst19687 (P3_ADD_380_U74, P3_ADD_380_U146, P3_ADD_380_U147);
  nand ginst19688 (P3_ADD_380_U75, P3_ADD_380_U148, P3_ADD_380_U149);
  nand ginst19689 (P3_ADD_380_U76, P3_ADD_380_U150, P3_ADD_380_U151);
  nand ginst19690 (P3_ADD_380_U77, P3_ADD_380_U152, P3_ADD_380_U153);
  nand ginst19691 (P3_ADD_380_U78, P3_ADD_380_U154, P3_ADD_380_U155);
  nand ginst19692 (P3_ADD_380_U79, P3_ADD_380_U156, P3_ADD_380_U157);
  not ginst19693 (P3_ADD_380_U8, P3_INSTADDRPOINTER_REG_2__SCAN_IN);
  nand ginst19694 (P3_ADD_380_U80, P3_ADD_380_U158, P3_ADD_380_U159);
  nand ginst19695 (P3_ADD_380_U81, P3_ADD_380_U160, P3_ADD_380_U161);
  nand ginst19696 (P3_ADD_380_U82, P3_ADD_380_U162, P3_ADD_380_U163);
  nand ginst19697 (P3_ADD_380_U83, P3_ADD_380_U164, P3_ADD_380_U165);
  nand ginst19698 (P3_ADD_380_U84, P3_ADD_380_U166, P3_ADD_380_U167);
  nand ginst19699 (P3_ADD_380_U85, P3_ADD_380_U168, P3_ADD_380_U169);
  nand ginst19700 (P3_ADD_380_U86, P3_ADD_380_U170, P3_ADD_380_U171);
  nand ginst19701 (P3_ADD_380_U87, P3_ADD_380_U172, P3_ADD_380_U173);
  nand ginst19702 (P3_ADD_380_U88, P3_ADD_380_U174, P3_ADD_380_U175);
  nand ginst19703 (P3_ADD_380_U89, P3_ADD_380_U176, P3_ADD_380_U177);
  nand ginst19704 (P3_ADD_380_U9, P3_INSTADDRPOINTER_REG_2__SCAN_IN, P3_ADD_380_U98);
  nand ginst19705 (P3_ADD_380_U90, P3_ADD_380_U178, P3_ADD_380_U179);
  nand ginst19706 (P3_ADD_380_U91, P3_ADD_380_U180, P3_ADD_380_U181);
  nand ginst19707 (P3_ADD_380_U92, P3_ADD_380_U182, P3_ADD_380_U183);
  nand ginst19708 (P3_ADD_380_U93, P3_ADD_380_U184, P3_ADD_380_U185);
  nand ginst19709 (P3_ADD_380_U94, P3_ADD_380_U186, P3_ADD_380_U187);
  nand ginst19710 (P3_ADD_380_U95, P3_ADD_380_U188, P3_ADD_380_U189);
  not ginst19711 (P3_ADD_380_U96, P3_INSTADDRPOINTER_REG_31__SCAN_IN);
  nand ginst19712 (P3_ADD_380_U97, P3_INSTADDRPOINTER_REG_30__SCAN_IN, P3_ADD_380_U126);
  not ginst19713 (P3_ADD_380_U98, P3_ADD_380_U7);
  not ginst19714 (P3_ADD_380_U99, P3_ADD_380_U9);
  not ginst19715 (P3_ADD_385_U10, P3_INSTADDRPOINTER_REG_3__SCAN_IN);
  not ginst19716 (P3_ADD_385_U100, P3_ADD_385_U11);
  not ginst19717 (P3_ADD_385_U101, P3_ADD_385_U13);
  not ginst19718 (P3_ADD_385_U102, P3_ADD_385_U15);
  not ginst19719 (P3_ADD_385_U103, P3_ADD_385_U17);
  not ginst19720 (P3_ADD_385_U104, P3_ADD_385_U19);
  not ginst19721 (P3_ADD_385_U105, P3_ADD_385_U22);
  not ginst19722 (P3_ADD_385_U106, P3_ADD_385_U23);
  not ginst19723 (P3_ADD_385_U107, P3_ADD_385_U25);
  not ginst19724 (P3_ADD_385_U108, P3_ADD_385_U27);
  not ginst19725 (P3_ADD_385_U109, P3_ADD_385_U29);
  nand ginst19726 (P3_ADD_385_U11, P3_INSTADDRPOINTER_REG_3__SCAN_IN, P3_ADD_385_U99);
  not ginst19727 (P3_ADD_385_U110, P3_ADD_385_U31);
  not ginst19728 (P3_ADD_385_U111, P3_ADD_385_U33);
  not ginst19729 (P3_ADD_385_U112, P3_ADD_385_U35);
  not ginst19730 (P3_ADD_385_U113, P3_ADD_385_U37);
  not ginst19731 (P3_ADD_385_U114, P3_ADD_385_U39);
  not ginst19732 (P3_ADD_385_U115, P3_ADD_385_U41);
  not ginst19733 (P3_ADD_385_U116, P3_ADD_385_U43);
  not ginst19734 (P3_ADD_385_U117, P3_ADD_385_U45);
  not ginst19735 (P3_ADD_385_U118, P3_ADD_385_U47);
  not ginst19736 (P3_ADD_385_U119, P3_ADD_385_U49);
  not ginst19737 (P3_ADD_385_U12, P3_INSTADDRPOINTER_REG_4__SCAN_IN);
  not ginst19738 (P3_ADD_385_U120, P3_ADD_385_U51);
  not ginst19739 (P3_ADD_385_U121, P3_ADD_385_U53);
  not ginst19740 (P3_ADD_385_U122, P3_ADD_385_U55);
  not ginst19741 (P3_ADD_385_U123, P3_ADD_385_U57);
  not ginst19742 (P3_ADD_385_U124, P3_ADD_385_U59);
  not ginst19743 (P3_ADD_385_U125, P3_ADD_385_U61);
  not ginst19744 (P3_ADD_385_U126, P3_ADD_385_U63);
  not ginst19745 (P3_ADD_385_U127, P3_ADD_385_U97);
  nand ginst19746 (P3_ADD_385_U128, P3_INSTADDRPOINTER_REG_9__SCAN_IN, P3_ADD_385_U22);
  nand ginst19747 (P3_ADD_385_U129, P3_ADD_385_U105, P3_ADD_385_U21);
  nand ginst19748 (P3_ADD_385_U13, P3_INSTADDRPOINTER_REG_4__SCAN_IN, P3_ADD_385_U100);
  nand ginst19749 (P3_ADD_385_U130, P3_INSTADDRPOINTER_REG_8__SCAN_IN, P3_ADD_385_U19);
  nand ginst19750 (P3_ADD_385_U131, P3_ADD_385_U104, P3_ADD_385_U20);
  nand ginst19751 (P3_ADD_385_U132, P3_INSTADDRPOINTER_REG_7__SCAN_IN, P3_ADD_385_U17);
  nand ginst19752 (P3_ADD_385_U133, P3_ADD_385_U103, P3_ADD_385_U18);
  nand ginst19753 (P3_ADD_385_U134, P3_INSTADDRPOINTER_REG_6__SCAN_IN, P3_ADD_385_U15);
  nand ginst19754 (P3_ADD_385_U135, P3_ADD_385_U102, P3_ADD_385_U16);
  nand ginst19755 (P3_ADD_385_U136, P3_INSTADDRPOINTER_REG_5__SCAN_IN, P3_ADD_385_U13);
  nand ginst19756 (P3_ADD_385_U137, P3_ADD_385_U101, P3_ADD_385_U14);
  nand ginst19757 (P3_ADD_385_U138, P3_INSTADDRPOINTER_REG_4__SCAN_IN, P3_ADD_385_U11);
  nand ginst19758 (P3_ADD_385_U139, P3_ADD_385_U100, P3_ADD_385_U12);
  not ginst19759 (P3_ADD_385_U14, P3_INSTADDRPOINTER_REG_5__SCAN_IN);
  nand ginst19760 (P3_ADD_385_U140, P3_INSTADDRPOINTER_REG_3__SCAN_IN, P3_ADD_385_U9);
  nand ginst19761 (P3_ADD_385_U141, P3_ADD_385_U10, P3_ADD_385_U99);
  nand ginst19762 (P3_ADD_385_U142, P3_INSTADDRPOINTER_REG_31__SCAN_IN, P3_ADD_385_U97);
  nand ginst19763 (P3_ADD_385_U143, P3_ADD_385_U127, P3_ADD_385_U96);
  nand ginst19764 (P3_ADD_385_U144, P3_INSTADDRPOINTER_REG_30__SCAN_IN, P3_ADD_385_U63);
  nand ginst19765 (P3_ADD_385_U145, P3_ADD_385_U126, P3_ADD_385_U64);
  nand ginst19766 (P3_ADD_385_U146, P3_INSTADDRPOINTER_REG_2__SCAN_IN, P3_ADD_385_U7);
  nand ginst19767 (P3_ADD_385_U147, P3_ADD_385_U8, P3_ADD_385_U98);
  nand ginst19768 (P3_ADD_385_U148, P3_INSTADDRPOINTER_REG_29__SCAN_IN, P3_ADD_385_U61);
  nand ginst19769 (P3_ADD_385_U149, P3_ADD_385_U125, P3_ADD_385_U62);
  nand ginst19770 (P3_ADD_385_U15, P3_INSTADDRPOINTER_REG_5__SCAN_IN, P3_ADD_385_U101);
  nand ginst19771 (P3_ADD_385_U150, P3_INSTADDRPOINTER_REG_28__SCAN_IN, P3_ADD_385_U59);
  nand ginst19772 (P3_ADD_385_U151, P3_ADD_385_U124, P3_ADD_385_U60);
  nand ginst19773 (P3_ADD_385_U152, P3_INSTADDRPOINTER_REG_27__SCAN_IN, P3_ADD_385_U57);
  nand ginst19774 (P3_ADD_385_U153, P3_ADD_385_U123, P3_ADD_385_U58);
  nand ginst19775 (P3_ADD_385_U154, P3_INSTADDRPOINTER_REG_26__SCAN_IN, P3_ADD_385_U55);
  nand ginst19776 (P3_ADD_385_U155, P3_ADD_385_U122, P3_ADD_385_U56);
  nand ginst19777 (P3_ADD_385_U156, P3_INSTADDRPOINTER_REG_25__SCAN_IN, P3_ADD_385_U53);
  nand ginst19778 (P3_ADD_385_U157, P3_ADD_385_U121, P3_ADD_385_U54);
  nand ginst19779 (P3_ADD_385_U158, P3_INSTADDRPOINTER_REG_24__SCAN_IN, P3_ADD_385_U51);
  nand ginst19780 (P3_ADD_385_U159, P3_ADD_385_U120, P3_ADD_385_U52);
  not ginst19781 (P3_ADD_385_U16, P3_INSTADDRPOINTER_REG_6__SCAN_IN);
  nand ginst19782 (P3_ADD_385_U160, P3_INSTADDRPOINTER_REG_23__SCAN_IN, P3_ADD_385_U49);
  nand ginst19783 (P3_ADD_385_U161, P3_ADD_385_U119, P3_ADD_385_U50);
  nand ginst19784 (P3_ADD_385_U162, P3_INSTADDRPOINTER_REG_22__SCAN_IN, P3_ADD_385_U47);
  nand ginst19785 (P3_ADD_385_U163, P3_ADD_385_U118, P3_ADD_385_U48);
  nand ginst19786 (P3_ADD_385_U164, P3_INSTADDRPOINTER_REG_21__SCAN_IN, P3_ADD_385_U45);
  nand ginst19787 (P3_ADD_385_U165, P3_ADD_385_U117, P3_ADD_385_U46);
  nand ginst19788 (P3_ADD_385_U166, P3_INSTADDRPOINTER_REG_20__SCAN_IN, P3_ADD_385_U43);
  nand ginst19789 (P3_ADD_385_U167, P3_ADD_385_U116, P3_ADD_385_U44);
  nand ginst19790 (P3_ADD_385_U168, P3_INSTADDRPOINTER_REG_1__SCAN_IN, P3_ADD_385_U5);
  nand ginst19791 (P3_ADD_385_U169, P3_INSTADDRPOINTER_REG_0__SCAN_IN, P3_ADD_385_U6);
  nand ginst19792 (P3_ADD_385_U17, P3_INSTADDRPOINTER_REG_6__SCAN_IN, P3_ADD_385_U102);
  nand ginst19793 (P3_ADD_385_U170, P3_INSTADDRPOINTER_REG_19__SCAN_IN, P3_ADD_385_U41);
  nand ginst19794 (P3_ADD_385_U171, P3_ADD_385_U115, P3_ADD_385_U42);
  nand ginst19795 (P3_ADD_385_U172, P3_INSTADDRPOINTER_REG_18__SCAN_IN, P3_ADD_385_U39);
  nand ginst19796 (P3_ADD_385_U173, P3_ADD_385_U114, P3_ADD_385_U40);
  nand ginst19797 (P3_ADD_385_U174, P3_INSTADDRPOINTER_REG_17__SCAN_IN, P3_ADD_385_U37);
  nand ginst19798 (P3_ADD_385_U175, P3_ADD_385_U113, P3_ADD_385_U38);
  nand ginst19799 (P3_ADD_385_U176, P3_INSTADDRPOINTER_REG_16__SCAN_IN, P3_ADD_385_U35);
  nand ginst19800 (P3_ADD_385_U177, P3_ADD_385_U112, P3_ADD_385_U36);
  nand ginst19801 (P3_ADD_385_U178, P3_INSTADDRPOINTER_REG_15__SCAN_IN, P3_ADD_385_U33);
  nand ginst19802 (P3_ADD_385_U179, P3_ADD_385_U111, P3_ADD_385_U34);
  not ginst19803 (P3_ADD_385_U18, P3_INSTADDRPOINTER_REG_7__SCAN_IN);
  nand ginst19804 (P3_ADD_385_U180, P3_INSTADDRPOINTER_REG_14__SCAN_IN, P3_ADD_385_U31);
  nand ginst19805 (P3_ADD_385_U181, P3_ADD_385_U110, P3_ADD_385_U32);
  nand ginst19806 (P3_ADD_385_U182, P3_INSTADDRPOINTER_REG_13__SCAN_IN, P3_ADD_385_U29);
  nand ginst19807 (P3_ADD_385_U183, P3_ADD_385_U109, P3_ADD_385_U30);
  nand ginst19808 (P3_ADD_385_U184, P3_INSTADDRPOINTER_REG_12__SCAN_IN, P3_ADD_385_U27);
  nand ginst19809 (P3_ADD_385_U185, P3_ADD_385_U108, P3_ADD_385_U28);
  nand ginst19810 (P3_ADD_385_U186, P3_INSTADDRPOINTER_REG_11__SCAN_IN, P3_ADD_385_U25);
  nand ginst19811 (P3_ADD_385_U187, P3_ADD_385_U107, P3_ADD_385_U26);
  nand ginst19812 (P3_ADD_385_U188, P3_INSTADDRPOINTER_REG_10__SCAN_IN, P3_ADD_385_U23);
  nand ginst19813 (P3_ADD_385_U189, P3_ADD_385_U106, P3_ADD_385_U24);
  nand ginst19814 (P3_ADD_385_U19, P3_INSTADDRPOINTER_REG_7__SCAN_IN, P3_ADD_385_U103);
  not ginst19815 (P3_ADD_385_U20, P3_INSTADDRPOINTER_REG_8__SCAN_IN);
  not ginst19816 (P3_ADD_385_U21, P3_INSTADDRPOINTER_REG_9__SCAN_IN);
  nand ginst19817 (P3_ADD_385_U22, P3_INSTADDRPOINTER_REG_8__SCAN_IN, P3_ADD_385_U104);
  nand ginst19818 (P3_ADD_385_U23, P3_INSTADDRPOINTER_REG_9__SCAN_IN, P3_ADD_385_U105);
  not ginst19819 (P3_ADD_385_U24, P3_INSTADDRPOINTER_REG_10__SCAN_IN);
  nand ginst19820 (P3_ADD_385_U25, P3_INSTADDRPOINTER_REG_10__SCAN_IN, P3_ADD_385_U106);
  not ginst19821 (P3_ADD_385_U26, P3_INSTADDRPOINTER_REG_11__SCAN_IN);
  nand ginst19822 (P3_ADD_385_U27, P3_INSTADDRPOINTER_REG_11__SCAN_IN, P3_ADD_385_U107);
  not ginst19823 (P3_ADD_385_U28, P3_INSTADDRPOINTER_REG_12__SCAN_IN);
  nand ginst19824 (P3_ADD_385_U29, P3_INSTADDRPOINTER_REG_12__SCAN_IN, P3_ADD_385_U108);
  not ginst19825 (P3_ADD_385_U30, P3_INSTADDRPOINTER_REG_13__SCAN_IN);
  nand ginst19826 (P3_ADD_385_U31, P3_INSTADDRPOINTER_REG_13__SCAN_IN, P3_ADD_385_U109);
  not ginst19827 (P3_ADD_385_U32, P3_INSTADDRPOINTER_REG_14__SCAN_IN);
  nand ginst19828 (P3_ADD_385_U33, P3_INSTADDRPOINTER_REG_14__SCAN_IN, P3_ADD_385_U110);
  not ginst19829 (P3_ADD_385_U34, P3_INSTADDRPOINTER_REG_15__SCAN_IN);
  nand ginst19830 (P3_ADD_385_U35, P3_INSTADDRPOINTER_REG_15__SCAN_IN, P3_ADD_385_U111);
  not ginst19831 (P3_ADD_385_U36, P3_INSTADDRPOINTER_REG_16__SCAN_IN);
  nand ginst19832 (P3_ADD_385_U37, P3_INSTADDRPOINTER_REG_16__SCAN_IN, P3_ADD_385_U112);
  not ginst19833 (P3_ADD_385_U38, P3_INSTADDRPOINTER_REG_17__SCAN_IN);
  nand ginst19834 (P3_ADD_385_U39, P3_INSTADDRPOINTER_REG_17__SCAN_IN, P3_ADD_385_U113);
  not ginst19835 (P3_ADD_385_U40, P3_INSTADDRPOINTER_REG_18__SCAN_IN);
  nand ginst19836 (P3_ADD_385_U41, P3_INSTADDRPOINTER_REG_18__SCAN_IN, P3_ADD_385_U114);
  not ginst19837 (P3_ADD_385_U42, P3_INSTADDRPOINTER_REG_19__SCAN_IN);
  nand ginst19838 (P3_ADD_385_U43, P3_INSTADDRPOINTER_REG_19__SCAN_IN, P3_ADD_385_U115);
  not ginst19839 (P3_ADD_385_U44, P3_INSTADDRPOINTER_REG_20__SCAN_IN);
  nand ginst19840 (P3_ADD_385_U45, P3_INSTADDRPOINTER_REG_20__SCAN_IN, P3_ADD_385_U116);
  not ginst19841 (P3_ADD_385_U46, P3_INSTADDRPOINTER_REG_21__SCAN_IN);
  nand ginst19842 (P3_ADD_385_U47, P3_INSTADDRPOINTER_REG_21__SCAN_IN, P3_ADD_385_U117);
  not ginst19843 (P3_ADD_385_U48, P3_INSTADDRPOINTER_REG_22__SCAN_IN);
  nand ginst19844 (P3_ADD_385_U49, P3_INSTADDRPOINTER_REG_22__SCAN_IN, P3_ADD_385_U118);
  not ginst19845 (P3_ADD_385_U5, P3_INSTADDRPOINTER_REG_0__SCAN_IN);
  not ginst19846 (P3_ADD_385_U50, P3_INSTADDRPOINTER_REG_23__SCAN_IN);
  nand ginst19847 (P3_ADD_385_U51, P3_INSTADDRPOINTER_REG_23__SCAN_IN, P3_ADD_385_U119);
  not ginst19848 (P3_ADD_385_U52, P3_INSTADDRPOINTER_REG_24__SCAN_IN);
  nand ginst19849 (P3_ADD_385_U53, P3_INSTADDRPOINTER_REG_24__SCAN_IN, P3_ADD_385_U120);
  not ginst19850 (P3_ADD_385_U54, P3_INSTADDRPOINTER_REG_25__SCAN_IN);
  nand ginst19851 (P3_ADD_385_U55, P3_INSTADDRPOINTER_REG_25__SCAN_IN, P3_ADD_385_U121);
  not ginst19852 (P3_ADD_385_U56, P3_INSTADDRPOINTER_REG_26__SCAN_IN);
  nand ginst19853 (P3_ADD_385_U57, P3_INSTADDRPOINTER_REG_26__SCAN_IN, P3_ADD_385_U122);
  not ginst19854 (P3_ADD_385_U58, P3_INSTADDRPOINTER_REG_27__SCAN_IN);
  nand ginst19855 (P3_ADD_385_U59, P3_INSTADDRPOINTER_REG_27__SCAN_IN, P3_ADD_385_U123);
  not ginst19856 (P3_ADD_385_U6, P3_INSTADDRPOINTER_REG_1__SCAN_IN);
  not ginst19857 (P3_ADD_385_U60, P3_INSTADDRPOINTER_REG_28__SCAN_IN);
  nand ginst19858 (P3_ADD_385_U61, P3_INSTADDRPOINTER_REG_28__SCAN_IN, P3_ADD_385_U124);
  not ginst19859 (P3_ADD_385_U62, P3_INSTADDRPOINTER_REG_29__SCAN_IN);
  nand ginst19860 (P3_ADD_385_U63, P3_INSTADDRPOINTER_REG_29__SCAN_IN, P3_ADD_385_U125);
  not ginst19861 (P3_ADD_385_U64, P3_INSTADDRPOINTER_REG_30__SCAN_IN);
  nand ginst19862 (P3_ADD_385_U65, P3_ADD_385_U128, P3_ADD_385_U129);
  nand ginst19863 (P3_ADD_385_U66, P3_ADD_385_U130, P3_ADD_385_U131);
  nand ginst19864 (P3_ADD_385_U67, P3_ADD_385_U132, P3_ADD_385_U133);
  nand ginst19865 (P3_ADD_385_U68, P3_ADD_385_U134, P3_ADD_385_U135);
  nand ginst19866 (P3_ADD_385_U69, P3_ADD_385_U136, P3_ADD_385_U137);
  nand ginst19867 (P3_ADD_385_U7, P3_INSTADDRPOINTER_REG_0__SCAN_IN, P3_INSTADDRPOINTER_REG_1__SCAN_IN);
  nand ginst19868 (P3_ADD_385_U70, P3_ADD_385_U138, P3_ADD_385_U139);
  nand ginst19869 (P3_ADD_385_U71, P3_ADD_385_U140, P3_ADD_385_U141);
  nand ginst19870 (P3_ADD_385_U72, P3_ADD_385_U142, P3_ADD_385_U143);
  nand ginst19871 (P3_ADD_385_U73, P3_ADD_385_U144, P3_ADD_385_U145);
  nand ginst19872 (P3_ADD_385_U74, P3_ADD_385_U146, P3_ADD_385_U147);
  nand ginst19873 (P3_ADD_385_U75, P3_ADD_385_U148, P3_ADD_385_U149);
  nand ginst19874 (P3_ADD_385_U76, P3_ADD_385_U150, P3_ADD_385_U151);
  nand ginst19875 (P3_ADD_385_U77, P3_ADD_385_U152, P3_ADD_385_U153);
  nand ginst19876 (P3_ADD_385_U78, P3_ADD_385_U154, P3_ADD_385_U155);
  nand ginst19877 (P3_ADD_385_U79, P3_ADD_385_U156, P3_ADD_385_U157);
  not ginst19878 (P3_ADD_385_U8, P3_INSTADDRPOINTER_REG_2__SCAN_IN);
  nand ginst19879 (P3_ADD_385_U80, P3_ADD_385_U158, P3_ADD_385_U159);
  nand ginst19880 (P3_ADD_385_U81, P3_ADD_385_U160, P3_ADD_385_U161);
  nand ginst19881 (P3_ADD_385_U82, P3_ADD_385_U162, P3_ADD_385_U163);
  nand ginst19882 (P3_ADD_385_U83, P3_ADD_385_U164, P3_ADD_385_U165);
  nand ginst19883 (P3_ADD_385_U84, P3_ADD_385_U166, P3_ADD_385_U167);
  nand ginst19884 (P3_ADD_385_U85, P3_ADD_385_U168, P3_ADD_385_U169);
  nand ginst19885 (P3_ADD_385_U86, P3_ADD_385_U170, P3_ADD_385_U171);
  nand ginst19886 (P3_ADD_385_U87, P3_ADD_385_U172, P3_ADD_385_U173);
  nand ginst19887 (P3_ADD_385_U88, P3_ADD_385_U174, P3_ADD_385_U175);
  nand ginst19888 (P3_ADD_385_U89, P3_ADD_385_U176, P3_ADD_385_U177);
  nand ginst19889 (P3_ADD_385_U9, P3_INSTADDRPOINTER_REG_2__SCAN_IN, P3_ADD_385_U98);
  nand ginst19890 (P3_ADD_385_U90, P3_ADD_385_U178, P3_ADD_385_U179);
  nand ginst19891 (P3_ADD_385_U91, P3_ADD_385_U180, P3_ADD_385_U181);
  nand ginst19892 (P3_ADD_385_U92, P3_ADD_385_U182, P3_ADD_385_U183);
  nand ginst19893 (P3_ADD_385_U93, P3_ADD_385_U184, P3_ADD_385_U185);
  nand ginst19894 (P3_ADD_385_U94, P3_ADD_385_U186, P3_ADD_385_U187);
  nand ginst19895 (P3_ADD_385_U95, P3_ADD_385_U188, P3_ADD_385_U189);
  not ginst19896 (P3_ADD_385_U96, P3_INSTADDRPOINTER_REG_31__SCAN_IN);
  nand ginst19897 (P3_ADD_385_U97, P3_INSTADDRPOINTER_REG_30__SCAN_IN, P3_ADD_385_U126);
  not ginst19898 (P3_ADD_385_U98, P3_ADD_385_U7);
  not ginst19899 (P3_ADD_385_U99, P3_ADD_385_U9);
  nand ginst19900 (P3_ADD_391_1180_U10, P3_ADD_391_1180_U29, P3_U2615);
  not ginst19901 (P3_ADD_391_1180_U11, P3_U2616);
  nand ginst19902 (P3_ADD_391_1180_U12, P3_ADD_391_1180_U30, P3_U2616);
  not ginst19903 (P3_ADD_391_1180_U13, P3_U2617);
  nand ginst19904 (P3_ADD_391_1180_U14, P3_ADD_391_1180_U31, P3_U2617);
  not ginst19905 (P3_ADD_391_1180_U15, P3_U2618);
  nand ginst19906 (P3_ADD_391_1180_U16, P3_ADD_391_1180_U32, P3_U2618);
  not ginst19907 (P3_ADD_391_1180_U17, P3_U2619);
  nand ginst19908 (P3_ADD_391_1180_U18, P3_ADD_391_1180_U35, P3_ADD_391_1180_U36);
  nand ginst19909 (P3_ADD_391_1180_U19, P3_ADD_391_1180_U37, P3_ADD_391_1180_U38);
  nand ginst19910 (P3_ADD_391_1180_U20, P3_ADD_391_1180_U39, P3_ADD_391_1180_U40);
  nand ginst19911 (P3_ADD_391_1180_U21, P3_ADD_391_1180_U41, P3_ADD_391_1180_U42);
  nand ginst19912 (P3_ADD_391_1180_U22, P3_ADD_391_1180_U43, P3_ADD_391_1180_U44);
  nand ginst19913 (P3_ADD_391_1180_U23, P3_ADD_391_1180_U45, P3_ADD_391_1180_U46);
  nand ginst19914 (P3_ADD_391_1180_U24, P3_ADD_391_1180_U47, P3_ADD_391_1180_U48);
  nand ginst19915 (P3_ADD_391_1180_U25, P3_ADD_391_1180_U49, P3_ADD_391_1180_U50);
  not ginst19916 (P3_ADD_391_1180_U26, P3_U2620);
  nand ginst19917 (P3_ADD_391_1180_U27, P3_ADD_391_1180_U33, P3_U2619);
  not ginst19918 (P3_ADD_391_1180_U28, P3_ADD_391_1180_U6);
  not ginst19919 (P3_ADD_391_1180_U29, P3_ADD_391_1180_U8);
  not ginst19920 (P3_ADD_391_1180_U30, P3_ADD_391_1180_U10);
  not ginst19921 (P3_ADD_391_1180_U31, P3_ADD_391_1180_U12);
  not ginst19922 (P3_ADD_391_1180_U32, P3_ADD_391_1180_U14);
  not ginst19923 (P3_ADD_391_1180_U33, P3_ADD_391_1180_U16);
  not ginst19924 (P3_ADD_391_1180_U34, P3_ADD_391_1180_U27);
  nand ginst19925 (P3_ADD_391_1180_U35, P3_ADD_391_1180_U27, P3_U2620);
  nand ginst19926 (P3_ADD_391_1180_U36, P3_ADD_391_1180_U26, P3_ADD_391_1180_U34);
  nand ginst19927 (P3_ADD_391_1180_U37, P3_ADD_391_1180_U16, P3_U2619);
  nand ginst19928 (P3_ADD_391_1180_U38, P3_ADD_391_1180_U17, P3_ADD_391_1180_U33);
  nand ginst19929 (P3_ADD_391_1180_U39, P3_ADD_391_1180_U14, P3_U2618);
  not ginst19930 (P3_ADD_391_1180_U4, P3_U2613);
  nand ginst19931 (P3_ADD_391_1180_U40, P3_ADD_391_1180_U15, P3_ADD_391_1180_U32);
  nand ginst19932 (P3_ADD_391_1180_U41, P3_ADD_391_1180_U12, P3_U2617);
  nand ginst19933 (P3_ADD_391_1180_U42, P3_ADD_391_1180_U13, P3_ADD_391_1180_U31);
  nand ginst19934 (P3_ADD_391_1180_U43, P3_ADD_391_1180_U10, P3_U2616);
  nand ginst19935 (P3_ADD_391_1180_U44, P3_ADD_391_1180_U11, P3_ADD_391_1180_U30);
  nand ginst19936 (P3_ADD_391_1180_U45, P3_ADD_391_1180_U8, P3_U2615);
  nand ginst19937 (P3_ADD_391_1180_U46, P3_ADD_391_1180_U29, P3_ADD_391_1180_U9);
  nand ginst19938 (P3_ADD_391_1180_U47, P3_ADD_391_1180_U6, P3_U2614);
  nand ginst19939 (P3_ADD_391_1180_U48, P3_ADD_391_1180_U28, P3_ADD_391_1180_U7);
  nand ginst19940 (P3_ADD_391_1180_U49, P3_ADD_391_1180_U4, P3_U3069);
  not ginst19941 (P3_ADD_391_1180_U5, P3_U3069);
  nand ginst19942 (P3_ADD_391_1180_U50, P3_ADD_391_1180_U5, P3_U2613);
  nand ginst19943 (P3_ADD_391_1180_U6, P3_U2613, P3_U3069);
  not ginst19944 (P3_ADD_391_1180_U7, P3_U2614);
  nand ginst19945 (P3_ADD_391_1180_U8, P3_ADD_391_1180_U28, P3_U2614);
  not ginst19946 (P3_ADD_391_1180_U9, P3_U2615);
  nand ginst19947 (P3_ADD_394_U10, P3_INSTADDRPOINTER_REG_4__SCAN_IN, P3_ADD_394_U98);
  not ginst19948 (P3_ADD_394_U100, P3_ADD_394_U12);
  not ginst19949 (P3_ADD_394_U101, P3_ADD_394_U14);
  not ginst19950 (P3_ADD_394_U102, P3_ADD_394_U16);
  not ginst19951 (P3_ADD_394_U103, P3_ADD_394_U19);
  not ginst19952 (P3_ADD_394_U104, P3_ADD_394_U20);
  not ginst19953 (P3_ADD_394_U105, P3_ADD_394_U22);
  not ginst19954 (P3_ADD_394_U106, P3_ADD_394_U24);
  not ginst19955 (P3_ADD_394_U107, P3_ADD_394_U26);
  not ginst19956 (P3_ADD_394_U108, P3_ADD_394_U28);
  not ginst19957 (P3_ADD_394_U109, P3_ADD_394_U30);
  not ginst19958 (P3_ADD_394_U11, P3_INSTADDRPOINTER_REG_5__SCAN_IN);
  not ginst19959 (P3_ADD_394_U110, P3_ADD_394_U32);
  not ginst19960 (P3_ADD_394_U111, P3_ADD_394_U34);
  not ginst19961 (P3_ADD_394_U112, P3_ADD_394_U36);
  not ginst19962 (P3_ADD_394_U113, P3_ADD_394_U38);
  not ginst19963 (P3_ADD_394_U114, P3_ADD_394_U40);
  not ginst19964 (P3_ADD_394_U115, P3_ADD_394_U42);
  not ginst19965 (P3_ADD_394_U116, P3_ADD_394_U44);
  not ginst19966 (P3_ADD_394_U117, P3_ADD_394_U46);
  not ginst19967 (P3_ADD_394_U118, P3_ADD_394_U48);
  not ginst19968 (P3_ADD_394_U119, P3_ADD_394_U50);
  nand ginst19969 (P3_ADD_394_U12, P3_INSTADDRPOINTER_REG_5__SCAN_IN, P3_ADD_394_U99);
  not ginst19970 (P3_ADD_394_U120, P3_ADD_394_U52);
  not ginst19971 (P3_ADD_394_U121, P3_ADD_394_U54);
  not ginst19972 (P3_ADD_394_U122, P3_ADD_394_U56);
  not ginst19973 (P3_ADD_394_U123, P3_ADD_394_U58);
  not ginst19974 (P3_ADD_394_U124, P3_ADD_394_U60);
  not ginst19975 (P3_ADD_394_U125, P3_ADD_394_U95);
  nand ginst19976 (P3_ADD_394_U126, P3_INSTADDRPOINTER_REG_0__SCAN_IN, P3_INSTADDRPOINTER_REG_1__SCAN_IN, P3_INSTADDRPOINTER_REG_2__SCAN_IN);
  nand ginst19977 (P3_ADD_394_U127, P3_INSTADDRPOINTER_REG_9__SCAN_IN, P3_ADD_394_U19);
  nand ginst19978 (P3_ADD_394_U128, P3_ADD_394_U103, P3_ADD_394_U18);
  nand ginst19979 (P3_ADD_394_U129, P3_INSTADDRPOINTER_REG_8__SCAN_IN, P3_ADD_394_U16);
  not ginst19980 (P3_ADD_394_U13, P3_INSTADDRPOINTER_REG_6__SCAN_IN);
  nand ginst19981 (P3_ADD_394_U130, P3_ADD_394_U102, P3_ADD_394_U17);
  nand ginst19982 (P3_ADD_394_U131, P3_INSTADDRPOINTER_REG_7__SCAN_IN, P3_ADD_394_U14);
  nand ginst19983 (P3_ADD_394_U132, P3_ADD_394_U101, P3_ADD_394_U15);
  nand ginst19984 (P3_ADD_394_U133, P3_INSTADDRPOINTER_REG_6__SCAN_IN, P3_ADD_394_U12);
  nand ginst19985 (P3_ADD_394_U134, P3_ADD_394_U100, P3_ADD_394_U13);
  nand ginst19986 (P3_ADD_394_U135, P3_INSTADDRPOINTER_REG_5__SCAN_IN, P3_ADD_394_U10);
  nand ginst19987 (P3_ADD_394_U136, P3_ADD_394_U11, P3_ADD_394_U99);
  nand ginst19988 (P3_ADD_394_U137, P3_INSTADDRPOINTER_REG_4__SCAN_IN, P3_ADD_394_U8);
  nand ginst19989 (P3_ADD_394_U138, P3_ADD_394_U9, P3_ADD_394_U98);
  nand ginst19990 (P3_ADD_394_U139, P3_INSTADDRPOINTER_REG_3__SCAN_IN, P3_ADD_394_U92);
  nand ginst19991 (P3_ADD_394_U14, P3_INSTADDRPOINTER_REG_6__SCAN_IN, P3_ADD_394_U100);
  nand ginst19992 (P3_ADD_394_U140, P3_ADD_394_U7, P3_ADD_394_U97);
  nand ginst19993 (P3_ADD_394_U141, P3_INSTADDRPOINTER_REG_31__SCAN_IN, P3_ADD_394_U95);
  nand ginst19994 (P3_ADD_394_U142, P3_ADD_394_U125, P3_ADD_394_U94);
  nand ginst19995 (P3_ADD_394_U143, P3_INSTADDRPOINTER_REG_30__SCAN_IN, P3_ADD_394_U60);
  nand ginst19996 (P3_ADD_394_U144, P3_ADD_394_U124, P3_ADD_394_U61);
  nand ginst19997 (P3_ADD_394_U145, P3_INSTADDRPOINTER_REG_29__SCAN_IN, P3_ADD_394_U58);
  nand ginst19998 (P3_ADD_394_U146, P3_ADD_394_U123, P3_ADD_394_U59);
  nand ginst19999 (P3_ADD_394_U147, P3_INSTADDRPOINTER_REG_28__SCAN_IN, P3_ADD_394_U56);
  nand ginst20000 (P3_ADD_394_U148, P3_ADD_394_U122, P3_ADD_394_U57);
  nand ginst20001 (P3_ADD_394_U149, P3_INSTADDRPOINTER_REG_27__SCAN_IN, P3_ADD_394_U54);
  not ginst20002 (P3_ADD_394_U15, P3_INSTADDRPOINTER_REG_7__SCAN_IN);
  nand ginst20003 (P3_ADD_394_U150, P3_ADD_394_U121, P3_ADD_394_U55);
  nand ginst20004 (P3_ADD_394_U151, P3_INSTADDRPOINTER_REG_26__SCAN_IN, P3_ADD_394_U52);
  nand ginst20005 (P3_ADD_394_U152, P3_ADD_394_U120, P3_ADD_394_U53);
  nand ginst20006 (P3_ADD_394_U153, P3_INSTADDRPOINTER_REG_25__SCAN_IN, P3_ADD_394_U50);
  nand ginst20007 (P3_ADD_394_U154, P3_ADD_394_U119, P3_ADD_394_U51);
  nand ginst20008 (P3_ADD_394_U155, P3_INSTADDRPOINTER_REG_24__SCAN_IN, P3_ADD_394_U48);
  nand ginst20009 (P3_ADD_394_U156, P3_ADD_394_U118, P3_ADD_394_U49);
  nand ginst20010 (P3_ADD_394_U157, P3_INSTADDRPOINTER_REG_23__SCAN_IN, P3_ADD_394_U46);
  nand ginst20011 (P3_ADD_394_U158, P3_ADD_394_U117, P3_ADD_394_U47);
  nand ginst20012 (P3_ADD_394_U159, P3_INSTADDRPOINTER_REG_22__SCAN_IN, P3_ADD_394_U44);
  nand ginst20013 (P3_ADD_394_U16, P3_INSTADDRPOINTER_REG_7__SCAN_IN, P3_ADD_394_U101);
  nand ginst20014 (P3_ADD_394_U160, P3_ADD_394_U116, P3_ADD_394_U45);
  nand ginst20015 (P3_ADD_394_U161, P3_INSTADDRPOINTER_REG_21__SCAN_IN, P3_ADD_394_U42);
  nand ginst20016 (P3_ADD_394_U162, P3_ADD_394_U115, P3_ADD_394_U43);
  nand ginst20017 (P3_ADD_394_U163, P3_INSTADDRPOINTER_REG_20__SCAN_IN, P3_ADD_394_U40);
  nand ginst20018 (P3_ADD_394_U164, P3_ADD_394_U114, P3_ADD_394_U41);
  nand ginst20019 (P3_ADD_394_U165, P3_INSTADDRPOINTER_REG_1__SCAN_IN, P3_ADD_394_U4);
  nand ginst20020 (P3_ADD_394_U166, P3_INSTADDRPOINTER_REG_0__SCAN_IN, P3_ADD_394_U6);
  nand ginst20021 (P3_ADD_394_U167, P3_INSTADDRPOINTER_REG_19__SCAN_IN, P3_ADD_394_U38);
  nand ginst20022 (P3_ADD_394_U168, P3_ADD_394_U113, P3_ADD_394_U39);
  nand ginst20023 (P3_ADD_394_U169, P3_INSTADDRPOINTER_REG_18__SCAN_IN, P3_ADD_394_U36);
  not ginst20024 (P3_ADD_394_U17, P3_INSTADDRPOINTER_REG_8__SCAN_IN);
  nand ginst20025 (P3_ADD_394_U170, P3_ADD_394_U112, P3_ADD_394_U37);
  nand ginst20026 (P3_ADD_394_U171, P3_INSTADDRPOINTER_REG_17__SCAN_IN, P3_ADD_394_U34);
  nand ginst20027 (P3_ADD_394_U172, P3_ADD_394_U111, P3_ADD_394_U35);
  nand ginst20028 (P3_ADD_394_U173, P3_INSTADDRPOINTER_REG_16__SCAN_IN, P3_ADD_394_U32);
  nand ginst20029 (P3_ADD_394_U174, P3_ADD_394_U110, P3_ADD_394_U33);
  nand ginst20030 (P3_ADD_394_U175, P3_INSTADDRPOINTER_REG_15__SCAN_IN, P3_ADD_394_U30);
  nand ginst20031 (P3_ADD_394_U176, P3_ADD_394_U109, P3_ADD_394_U31);
  nand ginst20032 (P3_ADD_394_U177, P3_INSTADDRPOINTER_REG_14__SCAN_IN, P3_ADD_394_U28);
  nand ginst20033 (P3_ADD_394_U178, P3_ADD_394_U108, P3_ADD_394_U29);
  nand ginst20034 (P3_ADD_394_U179, P3_INSTADDRPOINTER_REG_13__SCAN_IN, P3_ADD_394_U26);
  not ginst20035 (P3_ADD_394_U18, P3_INSTADDRPOINTER_REG_9__SCAN_IN);
  nand ginst20036 (P3_ADD_394_U180, P3_ADD_394_U107, P3_ADD_394_U27);
  nand ginst20037 (P3_ADD_394_U181, P3_INSTADDRPOINTER_REG_12__SCAN_IN, P3_ADD_394_U24);
  nand ginst20038 (P3_ADD_394_U182, P3_ADD_394_U106, P3_ADD_394_U25);
  nand ginst20039 (P3_ADD_394_U183, P3_INSTADDRPOINTER_REG_11__SCAN_IN, P3_ADD_394_U22);
  nand ginst20040 (P3_ADD_394_U184, P3_ADD_394_U105, P3_ADD_394_U23);
  nand ginst20041 (P3_ADD_394_U185, P3_INSTADDRPOINTER_REG_10__SCAN_IN, P3_ADD_394_U20);
  nand ginst20042 (P3_ADD_394_U186, P3_ADD_394_U104, P3_ADD_394_U21);
  nand ginst20043 (P3_ADD_394_U19, P3_INSTADDRPOINTER_REG_8__SCAN_IN, P3_ADD_394_U102);
  nand ginst20044 (P3_ADD_394_U20, P3_INSTADDRPOINTER_REG_9__SCAN_IN, P3_ADD_394_U103);
  not ginst20045 (P3_ADD_394_U21, P3_INSTADDRPOINTER_REG_10__SCAN_IN);
  nand ginst20046 (P3_ADD_394_U22, P3_INSTADDRPOINTER_REG_10__SCAN_IN, P3_ADD_394_U104);
  not ginst20047 (P3_ADD_394_U23, P3_INSTADDRPOINTER_REG_11__SCAN_IN);
  nand ginst20048 (P3_ADD_394_U24, P3_INSTADDRPOINTER_REG_11__SCAN_IN, P3_ADD_394_U105);
  not ginst20049 (P3_ADD_394_U25, P3_INSTADDRPOINTER_REG_12__SCAN_IN);
  nand ginst20050 (P3_ADD_394_U26, P3_INSTADDRPOINTER_REG_12__SCAN_IN, P3_ADD_394_U106);
  not ginst20051 (P3_ADD_394_U27, P3_INSTADDRPOINTER_REG_13__SCAN_IN);
  nand ginst20052 (P3_ADD_394_U28, P3_INSTADDRPOINTER_REG_13__SCAN_IN, P3_ADD_394_U107);
  not ginst20053 (P3_ADD_394_U29, P3_INSTADDRPOINTER_REG_14__SCAN_IN);
  nand ginst20054 (P3_ADD_394_U30, P3_INSTADDRPOINTER_REG_14__SCAN_IN, P3_ADD_394_U108);
  not ginst20055 (P3_ADD_394_U31, P3_INSTADDRPOINTER_REG_15__SCAN_IN);
  nand ginst20056 (P3_ADD_394_U32, P3_INSTADDRPOINTER_REG_15__SCAN_IN, P3_ADD_394_U109);
  not ginst20057 (P3_ADD_394_U33, P3_INSTADDRPOINTER_REG_16__SCAN_IN);
  nand ginst20058 (P3_ADD_394_U34, P3_INSTADDRPOINTER_REG_16__SCAN_IN, P3_ADD_394_U110);
  not ginst20059 (P3_ADD_394_U35, P3_INSTADDRPOINTER_REG_17__SCAN_IN);
  nand ginst20060 (P3_ADD_394_U36, P3_INSTADDRPOINTER_REG_17__SCAN_IN, P3_ADD_394_U111);
  not ginst20061 (P3_ADD_394_U37, P3_INSTADDRPOINTER_REG_18__SCAN_IN);
  nand ginst20062 (P3_ADD_394_U38, P3_INSTADDRPOINTER_REG_18__SCAN_IN, P3_ADD_394_U112);
  not ginst20063 (P3_ADD_394_U39, P3_INSTADDRPOINTER_REG_19__SCAN_IN);
  not ginst20064 (P3_ADD_394_U4, P3_INSTADDRPOINTER_REG_0__SCAN_IN);
  nand ginst20065 (P3_ADD_394_U40, P3_INSTADDRPOINTER_REG_19__SCAN_IN, P3_ADD_394_U113);
  not ginst20066 (P3_ADD_394_U41, P3_INSTADDRPOINTER_REG_20__SCAN_IN);
  nand ginst20067 (P3_ADD_394_U42, P3_INSTADDRPOINTER_REG_20__SCAN_IN, P3_ADD_394_U114);
  not ginst20068 (P3_ADD_394_U43, P3_INSTADDRPOINTER_REG_21__SCAN_IN);
  nand ginst20069 (P3_ADD_394_U44, P3_INSTADDRPOINTER_REG_21__SCAN_IN, P3_ADD_394_U115);
  not ginst20070 (P3_ADD_394_U45, P3_INSTADDRPOINTER_REG_22__SCAN_IN);
  nand ginst20071 (P3_ADD_394_U46, P3_INSTADDRPOINTER_REG_22__SCAN_IN, P3_ADD_394_U116);
  not ginst20072 (P3_ADD_394_U47, P3_INSTADDRPOINTER_REG_23__SCAN_IN);
  nand ginst20073 (P3_ADD_394_U48, P3_INSTADDRPOINTER_REG_23__SCAN_IN, P3_ADD_394_U117);
  not ginst20074 (P3_ADD_394_U49, P3_INSTADDRPOINTER_REG_24__SCAN_IN);
  nand ginst20075 (P3_ADD_394_U5, P3_ADD_394_U126, P3_ADD_394_U92);
  nand ginst20076 (P3_ADD_394_U50, P3_INSTADDRPOINTER_REG_24__SCAN_IN, P3_ADD_394_U118);
  not ginst20077 (P3_ADD_394_U51, P3_INSTADDRPOINTER_REG_25__SCAN_IN);
  nand ginst20078 (P3_ADD_394_U52, P3_INSTADDRPOINTER_REG_25__SCAN_IN, P3_ADD_394_U119);
  not ginst20079 (P3_ADD_394_U53, P3_INSTADDRPOINTER_REG_26__SCAN_IN);
  nand ginst20080 (P3_ADD_394_U54, P3_INSTADDRPOINTER_REG_26__SCAN_IN, P3_ADD_394_U120);
  not ginst20081 (P3_ADD_394_U55, P3_INSTADDRPOINTER_REG_27__SCAN_IN);
  nand ginst20082 (P3_ADD_394_U56, P3_INSTADDRPOINTER_REG_27__SCAN_IN, P3_ADD_394_U121);
  not ginst20083 (P3_ADD_394_U57, P3_INSTADDRPOINTER_REG_28__SCAN_IN);
  nand ginst20084 (P3_ADD_394_U58, P3_INSTADDRPOINTER_REG_28__SCAN_IN, P3_ADD_394_U122);
  not ginst20085 (P3_ADD_394_U59, P3_INSTADDRPOINTER_REG_29__SCAN_IN);
  not ginst20086 (P3_ADD_394_U6, P3_INSTADDRPOINTER_REG_1__SCAN_IN);
  nand ginst20087 (P3_ADD_394_U60, P3_INSTADDRPOINTER_REG_29__SCAN_IN, P3_ADD_394_U123);
  not ginst20088 (P3_ADD_394_U61, P3_INSTADDRPOINTER_REG_30__SCAN_IN);
  not ginst20089 (P3_ADD_394_U62, P3_INSTADDRPOINTER_REG_2__SCAN_IN);
  nand ginst20090 (P3_ADD_394_U63, P3_ADD_394_U127, P3_ADD_394_U128);
  nand ginst20091 (P3_ADD_394_U64, P3_ADD_394_U129, P3_ADD_394_U130);
  nand ginst20092 (P3_ADD_394_U65, P3_ADD_394_U131, P3_ADD_394_U132);
  nand ginst20093 (P3_ADD_394_U66, P3_ADD_394_U133, P3_ADD_394_U134);
  nand ginst20094 (P3_ADD_394_U67, P3_ADD_394_U135, P3_ADD_394_U136);
  nand ginst20095 (P3_ADD_394_U68, P3_ADD_394_U137, P3_ADD_394_U138);
  nand ginst20096 (P3_ADD_394_U69, P3_ADD_394_U141, P3_ADD_394_U142);
  not ginst20097 (P3_ADD_394_U7, P3_INSTADDRPOINTER_REG_3__SCAN_IN);
  nand ginst20098 (P3_ADD_394_U70, P3_ADD_394_U143, P3_ADD_394_U144);
  nand ginst20099 (P3_ADD_394_U71, P3_ADD_394_U145, P3_ADD_394_U146);
  nand ginst20100 (P3_ADD_394_U72, P3_ADD_394_U147, P3_ADD_394_U148);
  nand ginst20101 (P3_ADD_394_U73, P3_ADD_394_U149, P3_ADD_394_U150);
  nand ginst20102 (P3_ADD_394_U74, P3_ADD_394_U151, P3_ADD_394_U152);
  nand ginst20103 (P3_ADD_394_U75, P3_ADD_394_U153, P3_ADD_394_U154);
  nand ginst20104 (P3_ADD_394_U76, P3_ADD_394_U155, P3_ADD_394_U156);
  nand ginst20105 (P3_ADD_394_U77, P3_ADD_394_U157, P3_ADD_394_U158);
  nand ginst20106 (P3_ADD_394_U78, P3_ADD_394_U159, P3_ADD_394_U160);
  nand ginst20107 (P3_ADD_394_U79, P3_ADD_394_U161, P3_ADD_394_U162);
  nand ginst20108 (P3_ADD_394_U8, P3_INSTADDRPOINTER_REG_3__SCAN_IN, P3_ADD_394_U92);
  nand ginst20109 (P3_ADD_394_U80, P3_ADD_394_U163, P3_ADD_394_U164);
  nand ginst20110 (P3_ADD_394_U81, P3_ADD_394_U165, P3_ADD_394_U166);
  nand ginst20111 (P3_ADD_394_U82, P3_ADD_394_U167, P3_ADD_394_U168);
  nand ginst20112 (P3_ADD_394_U83, P3_ADD_394_U169, P3_ADD_394_U170);
  nand ginst20113 (P3_ADD_394_U84, P3_ADD_394_U171, P3_ADD_394_U172);
  nand ginst20114 (P3_ADD_394_U85, P3_ADD_394_U173, P3_ADD_394_U174);
  nand ginst20115 (P3_ADD_394_U86, P3_ADD_394_U175, P3_ADD_394_U176);
  nand ginst20116 (P3_ADD_394_U87, P3_ADD_394_U177, P3_ADD_394_U178);
  nand ginst20117 (P3_ADD_394_U88, P3_ADD_394_U179, P3_ADD_394_U180);
  nand ginst20118 (P3_ADD_394_U89, P3_ADD_394_U181, P3_ADD_394_U182);
  not ginst20119 (P3_ADD_394_U9, P3_INSTADDRPOINTER_REG_4__SCAN_IN);
  nand ginst20120 (P3_ADD_394_U90, P3_ADD_394_U183, P3_ADD_394_U184);
  nand ginst20121 (P3_ADD_394_U91, P3_ADD_394_U185, P3_ADD_394_U186);
  nand ginst20122 (P3_ADD_394_U92, P3_ADD_394_U62, P3_ADD_394_U96);
  and ginst20123 (P3_ADD_394_U93, P3_ADD_394_U139, P3_ADD_394_U140);
  not ginst20124 (P3_ADD_394_U94, P3_INSTADDRPOINTER_REG_31__SCAN_IN);
  nand ginst20125 (P3_ADD_394_U95, P3_INSTADDRPOINTER_REG_30__SCAN_IN, P3_ADD_394_U124);
  nand ginst20126 (P3_ADD_394_U96, P3_INSTADDRPOINTER_REG_0__SCAN_IN, P3_INSTADDRPOINTER_REG_1__SCAN_IN);
  not ginst20127 (P3_ADD_394_U97, P3_ADD_394_U92);
  not ginst20128 (P3_ADD_394_U98, P3_ADD_394_U8);
  not ginst20129 (P3_ADD_394_U99, P3_ADD_394_U10);
  nand ginst20130 (P3_ADD_402_1132_U10, P3_ADD_402_1132_U29, P3_U2615);
  not ginst20131 (P3_ADD_402_1132_U11, P3_U2616);
  nand ginst20132 (P3_ADD_402_1132_U12, P3_ADD_402_1132_U30, P3_U2616);
  not ginst20133 (P3_ADD_402_1132_U13, P3_U2617);
  nand ginst20134 (P3_ADD_402_1132_U14, P3_ADD_402_1132_U31, P3_U2617);
  not ginst20135 (P3_ADD_402_1132_U15, P3_U2618);
  nand ginst20136 (P3_ADD_402_1132_U16, P3_ADD_402_1132_U32, P3_U2618);
  not ginst20137 (P3_ADD_402_1132_U17, P3_U2619);
  nand ginst20138 (P3_ADD_402_1132_U18, P3_ADD_402_1132_U35, P3_ADD_402_1132_U36);
  nand ginst20139 (P3_ADD_402_1132_U19, P3_ADD_402_1132_U37, P3_ADD_402_1132_U38);
  nand ginst20140 (P3_ADD_402_1132_U20, P3_ADD_402_1132_U39, P3_ADD_402_1132_U40);
  nand ginst20141 (P3_ADD_402_1132_U21, P3_ADD_402_1132_U41, P3_ADD_402_1132_U42);
  nand ginst20142 (P3_ADD_402_1132_U22, P3_ADD_402_1132_U43, P3_ADD_402_1132_U44);
  nand ginst20143 (P3_ADD_402_1132_U23, P3_ADD_402_1132_U45, P3_ADD_402_1132_U46);
  nand ginst20144 (P3_ADD_402_1132_U24, P3_ADD_402_1132_U47, P3_ADD_402_1132_U48);
  nand ginst20145 (P3_ADD_402_1132_U25, P3_ADD_402_1132_U49, P3_ADD_402_1132_U50);
  not ginst20146 (P3_ADD_402_1132_U26, P3_U2620);
  nand ginst20147 (P3_ADD_402_1132_U27, P3_ADD_402_1132_U33, P3_U2619);
  not ginst20148 (P3_ADD_402_1132_U28, P3_ADD_402_1132_U6);
  not ginst20149 (P3_ADD_402_1132_U29, P3_ADD_402_1132_U8);
  not ginst20150 (P3_ADD_402_1132_U30, P3_ADD_402_1132_U10);
  not ginst20151 (P3_ADD_402_1132_U31, P3_ADD_402_1132_U12);
  not ginst20152 (P3_ADD_402_1132_U32, P3_ADD_402_1132_U14);
  not ginst20153 (P3_ADD_402_1132_U33, P3_ADD_402_1132_U16);
  not ginst20154 (P3_ADD_402_1132_U34, P3_ADD_402_1132_U27);
  nand ginst20155 (P3_ADD_402_1132_U35, P3_ADD_402_1132_U27, P3_U2620);
  nand ginst20156 (P3_ADD_402_1132_U36, P3_ADD_402_1132_U26, P3_ADD_402_1132_U34);
  nand ginst20157 (P3_ADD_402_1132_U37, P3_ADD_402_1132_U16, P3_U2619);
  nand ginst20158 (P3_ADD_402_1132_U38, P3_ADD_402_1132_U17, P3_ADD_402_1132_U33);
  nand ginst20159 (P3_ADD_402_1132_U39, P3_ADD_402_1132_U14, P3_U2618);
  not ginst20160 (P3_ADD_402_1132_U4, P3_U2613);
  nand ginst20161 (P3_ADD_402_1132_U40, P3_ADD_402_1132_U15, P3_ADD_402_1132_U32);
  nand ginst20162 (P3_ADD_402_1132_U41, P3_ADD_402_1132_U12, P3_U2617);
  nand ginst20163 (P3_ADD_402_1132_U42, P3_ADD_402_1132_U13, P3_ADD_402_1132_U31);
  nand ginst20164 (P3_ADD_402_1132_U43, P3_ADD_402_1132_U10, P3_U2616);
  nand ginst20165 (P3_ADD_402_1132_U44, P3_ADD_402_1132_U11, P3_ADD_402_1132_U30);
  nand ginst20166 (P3_ADD_402_1132_U45, P3_ADD_402_1132_U8, P3_U2615);
  nand ginst20167 (P3_ADD_402_1132_U46, P3_ADD_402_1132_U29, P3_ADD_402_1132_U9);
  nand ginst20168 (P3_ADD_402_1132_U47, P3_ADD_402_1132_U6, P3_U2614);
  nand ginst20169 (P3_ADD_402_1132_U48, P3_ADD_402_1132_U28, P3_ADD_402_1132_U7);
  nand ginst20170 (P3_ADD_402_1132_U49, P3_ADD_402_1132_U4, P3_U3069);
  not ginst20171 (P3_ADD_402_1132_U5, P3_U3069);
  nand ginst20172 (P3_ADD_402_1132_U50, P3_ADD_402_1132_U5, P3_U2613);
  nand ginst20173 (P3_ADD_402_1132_U6, P3_U2613, P3_U3069);
  not ginst20174 (P3_ADD_402_1132_U7, P3_U2614);
  nand ginst20175 (P3_ADD_402_1132_U8, P3_ADD_402_1132_U28, P3_U2614);
  not ginst20176 (P3_ADD_402_1132_U9, P3_U2615);
  nand ginst20177 (P3_ADD_405_U10, P3_INSTADDRPOINTER_REG_4__SCAN_IN, P3_ADD_405_U98);
  not ginst20178 (P3_ADD_405_U100, P3_ADD_405_U12);
  not ginst20179 (P3_ADD_405_U101, P3_ADD_405_U14);
  not ginst20180 (P3_ADD_405_U102, P3_ADD_405_U16);
  not ginst20181 (P3_ADD_405_U103, P3_ADD_405_U19);
  not ginst20182 (P3_ADD_405_U104, P3_ADD_405_U20);
  not ginst20183 (P3_ADD_405_U105, P3_ADD_405_U22);
  not ginst20184 (P3_ADD_405_U106, P3_ADD_405_U24);
  not ginst20185 (P3_ADD_405_U107, P3_ADD_405_U26);
  not ginst20186 (P3_ADD_405_U108, P3_ADD_405_U28);
  not ginst20187 (P3_ADD_405_U109, P3_ADD_405_U30);
  not ginst20188 (P3_ADD_405_U11, P3_INSTADDRPOINTER_REG_5__SCAN_IN);
  not ginst20189 (P3_ADD_405_U110, P3_ADD_405_U32);
  not ginst20190 (P3_ADD_405_U111, P3_ADD_405_U34);
  not ginst20191 (P3_ADD_405_U112, P3_ADD_405_U36);
  not ginst20192 (P3_ADD_405_U113, P3_ADD_405_U38);
  not ginst20193 (P3_ADD_405_U114, P3_ADD_405_U40);
  not ginst20194 (P3_ADD_405_U115, P3_ADD_405_U42);
  not ginst20195 (P3_ADD_405_U116, P3_ADD_405_U44);
  not ginst20196 (P3_ADD_405_U117, P3_ADD_405_U46);
  not ginst20197 (P3_ADD_405_U118, P3_ADD_405_U48);
  not ginst20198 (P3_ADD_405_U119, P3_ADD_405_U50);
  nand ginst20199 (P3_ADD_405_U12, P3_INSTADDRPOINTER_REG_5__SCAN_IN, P3_ADD_405_U99);
  not ginst20200 (P3_ADD_405_U120, P3_ADD_405_U52);
  not ginst20201 (P3_ADD_405_U121, P3_ADD_405_U54);
  not ginst20202 (P3_ADD_405_U122, P3_ADD_405_U56);
  not ginst20203 (P3_ADD_405_U123, P3_ADD_405_U58);
  not ginst20204 (P3_ADD_405_U124, P3_ADD_405_U60);
  not ginst20205 (P3_ADD_405_U125, P3_ADD_405_U95);
  nand ginst20206 (P3_ADD_405_U126, P3_INSTADDRPOINTER_REG_0__SCAN_IN, P3_INSTADDRPOINTER_REG_1__SCAN_IN, P3_INSTADDRPOINTER_REG_2__SCAN_IN);
  nand ginst20207 (P3_ADD_405_U127, P3_INSTADDRPOINTER_REG_9__SCAN_IN, P3_ADD_405_U19);
  nand ginst20208 (P3_ADD_405_U128, P3_ADD_405_U103, P3_ADD_405_U18);
  nand ginst20209 (P3_ADD_405_U129, P3_INSTADDRPOINTER_REG_8__SCAN_IN, P3_ADD_405_U16);
  not ginst20210 (P3_ADD_405_U13, P3_INSTADDRPOINTER_REG_6__SCAN_IN);
  nand ginst20211 (P3_ADD_405_U130, P3_ADD_405_U102, P3_ADD_405_U17);
  nand ginst20212 (P3_ADD_405_U131, P3_INSTADDRPOINTER_REG_7__SCAN_IN, P3_ADD_405_U14);
  nand ginst20213 (P3_ADD_405_U132, P3_ADD_405_U101, P3_ADD_405_U15);
  nand ginst20214 (P3_ADD_405_U133, P3_INSTADDRPOINTER_REG_6__SCAN_IN, P3_ADD_405_U12);
  nand ginst20215 (P3_ADD_405_U134, P3_ADD_405_U100, P3_ADD_405_U13);
  nand ginst20216 (P3_ADD_405_U135, P3_INSTADDRPOINTER_REG_5__SCAN_IN, P3_ADD_405_U10);
  nand ginst20217 (P3_ADD_405_U136, P3_ADD_405_U11, P3_ADD_405_U99);
  nand ginst20218 (P3_ADD_405_U137, P3_INSTADDRPOINTER_REG_4__SCAN_IN, P3_ADD_405_U8);
  nand ginst20219 (P3_ADD_405_U138, P3_ADD_405_U9, P3_ADD_405_U98);
  nand ginst20220 (P3_ADD_405_U139, P3_INSTADDRPOINTER_REG_3__SCAN_IN, P3_ADD_405_U92);
  nand ginst20221 (P3_ADD_405_U14, P3_INSTADDRPOINTER_REG_6__SCAN_IN, P3_ADD_405_U100);
  nand ginst20222 (P3_ADD_405_U140, P3_ADD_405_U7, P3_ADD_405_U97);
  nand ginst20223 (P3_ADD_405_U141, P3_INSTADDRPOINTER_REG_31__SCAN_IN, P3_ADD_405_U95);
  nand ginst20224 (P3_ADD_405_U142, P3_ADD_405_U125, P3_ADD_405_U94);
  nand ginst20225 (P3_ADD_405_U143, P3_INSTADDRPOINTER_REG_30__SCAN_IN, P3_ADD_405_U60);
  nand ginst20226 (P3_ADD_405_U144, P3_ADD_405_U124, P3_ADD_405_U61);
  nand ginst20227 (P3_ADD_405_U145, P3_INSTADDRPOINTER_REG_29__SCAN_IN, P3_ADD_405_U58);
  nand ginst20228 (P3_ADD_405_U146, P3_ADD_405_U123, P3_ADD_405_U59);
  nand ginst20229 (P3_ADD_405_U147, P3_INSTADDRPOINTER_REG_28__SCAN_IN, P3_ADD_405_U56);
  nand ginst20230 (P3_ADD_405_U148, P3_ADD_405_U122, P3_ADD_405_U57);
  nand ginst20231 (P3_ADD_405_U149, P3_INSTADDRPOINTER_REG_27__SCAN_IN, P3_ADD_405_U54);
  not ginst20232 (P3_ADD_405_U15, P3_INSTADDRPOINTER_REG_7__SCAN_IN);
  nand ginst20233 (P3_ADD_405_U150, P3_ADD_405_U121, P3_ADD_405_U55);
  nand ginst20234 (P3_ADD_405_U151, P3_INSTADDRPOINTER_REG_26__SCAN_IN, P3_ADD_405_U52);
  nand ginst20235 (P3_ADD_405_U152, P3_ADD_405_U120, P3_ADD_405_U53);
  nand ginst20236 (P3_ADD_405_U153, P3_INSTADDRPOINTER_REG_25__SCAN_IN, P3_ADD_405_U50);
  nand ginst20237 (P3_ADD_405_U154, P3_ADD_405_U119, P3_ADD_405_U51);
  nand ginst20238 (P3_ADD_405_U155, P3_INSTADDRPOINTER_REG_24__SCAN_IN, P3_ADD_405_U48);
  nand ginst20239 (P3_ADD_405_U156, P3_ADD_405_U118, P3_ADD_405_U49);
  nand ginst20240 (P3_ADD_405_U157, P3_INSTADDRPOINTER_REG_23__SCAN_IN, P3_ADD_405_U46);
  nand ginst20241 (P3_ADD_405_U158, P3_ADD_405_U117, P3_ADD_405_U47);
  nand ginst20242 (P3_ADD_405_U159, P3_INSTADDRPOINTER_REG_22__SCAN_IN, P3_ADD_405_U44);
  nand ginst20243 (P3_ADD_405_U16, P3_INSTADDRPOINTER_REG_7__SCAN_IN, P3_ADD_405_U101);
  nand ginst20244 (P3_ADD_405_U160, P3_ADD_405_U116, P3_ADD_405_U45);
  nand ginst20245 (P3_ADD_405_U161, P3_INSTADDRPOINTER_REG_21__SCAN_IN, P3_ADD_405_U42);
  nand ginst20246 (P3_ADD_405_U162, P3_ADD_405_U115, P3_ADD_405_U43);
  nand ginst20247 (P3_ADD_405_U163, P3_INSTADDRPOINTER_REG_20__SCAN_IN, P3_ADD_405_U40);
  nand ginst20248 (P3_ADD_405_U164, P3_ADD_405_U114, P3_ADD_405_U41);
  nand ginst20249 (P3_ADD_405_U165, P3_INSTADDRPOINTER_REG_1__SCAN_IN, P3_ADD_405_U4);
  nand ginst20250 (P3_ADD_405_U166, P3_INSTADDRPOINTER_REG_0__SCAN_IN, P3_ADD_405_U6);
  nand ginst20251 (P3_ADD_405_U167, P3_INSTADDRPOINTER_REG_19__SCAN_IN, P3_ADD_405_U38);
  nand ginst20252 (P3_ADD_405_U168, P3_ADD_405_U113, P3_ADD_405_U39);
  nand ginst20253 (P3_ADD_405_U169, P3_INSTADDRPOINTER_REG_18__SCAN_IN, P3_ADD_405_U36);
  not ginst20254 (P3_ADD_405_U17, P3_INSTADDRPOINTER_REG_8__SCAN_IN);
  nand ginst20255 (P3_ADD_405_U170, P3_ADD_405_U112, P3_ADD_405_U37);
  nand ginst20256 (P3_ADD_405_U171, P3_INSTADDRPOINTER_REG_17__SCAN_IN, P3_ADD_405_U34);
  nand ginst20257 (P3_ADD_405_U172, P3_ADD_405_U111, P3_ADD_405_U35);
  nand ginst20258 (P3_ADD_405_U173, P3_INSTADDRPOINTER_REG_16__SCAN_IN, P3_ADD_405_U32);
  nand ginst20259 (P3_ADD_405_U174, P3_ADD_405_U110, P3_ADD_405_U33);
  nand ginst20260 (P3_ADD_405_U175, P3_INSTADDRPOINTER_REG_15__SCAN_IN, P3_ADD_405_U30);
  nand ginst20261 (P3_ADD_405_U176, P3_ADD_405_U109, P3_ADD_405_U31);
  nand ginst20262 (P3_ADD_405_U177, P3_INSTADDRPOINTER_REG_14__SCAN_IN, P3_ADD_405_U28);
  nand ginst20263 (P3_ADD_405_U178, P3_ADD_405_U108, P3_ADD_405_U29);
  nand ginst20264 (P3_ADD_405_U179, P3_INSTADDRPOINTER_REG_13__SCAN_IN, P3_ADD_405_U26);
  not ginst20265 (P3_ADD_405_U18, P3_INSTADDRPOINTER_REG_9__SCAN_IN);
  nand ginst20266 (P3_ADD_405_U180, P3_ADD_405_U107, P3_ADD_405_U27);
  nand ginst20267 (P3_ADD_405_U181, P3_INSTADDRPOINTER_REG_12__SCAN_IN, P3_ADD_405_U24);
  nand ginst20268 (P3_ADD_405_U182, P3_ADD_405_U106, P3_ADD_405_U25);
  nand ginst20269 (P3_ADD_405_U183, P3_INSTADDRPOINTER_REG_11__SCAN_IN, P3_ADD_405_U22);
  nand ginst20270 (P3_ADD_405_U184, P3_ADD_405_U105, P3_ADD_405_U23);
  nand ginst20271 (P3_ADD_405_U185, P3_INSTADDRPOINTER_REG_10__SCAN_IN, P3_ADD_405_U20);
  nand ginst20272 (P3_ADD_405_U186, P3_ADD_405_U104, P3_ADD_405_U21);
  nand ginst20273 (P3_ADD_405_U19, P3_INSTADDRPOINTER_REG_8__SCAN_IN, P3_ADD_405_U102);
  nand ginst20274 (P3_ADD_405_U20, P3_INSTADDRPOINTER_REG_9__SCAN_IN, P3_ADD_405_U103);
  not ginst20275 (P3_ADD_405_U21, P3_INSTADDRPOINTER_REG_10__SCAN_IN);
  nand ginst20276 (P3_ADD_405_U22, P3_INSTADDRPOINTER_REG_10__SCAN_IN, P3_ADD_405_U104);
  not ginst20277 (P3_ADD_405_U23, P3_INSTADDRPOINTER_REG_11__SCAN_IN);
  nand ginst20278 (P3_ADD_405_U24, P3_INSTADDRPOINTER_REG_11__SCAN_IN, P3_ADD_405_U105);
  not ginst20279 (P3_ADD_405_U25, P3_INSTADDRPOINTER_REG_12__SCAN_IN);
  nand ginst20280 (P3_ADD_405_U26, P3_INSTADDRPOINTER_REG_12__SCAN_IN, P3_ADD_405_U106);
  not ginst20281 (P3_ADD_405_U27, P3_INSTADDRPOINTER_REG_13__SCAN_IN);
  nand ginst20282 (P3_ADD_405_U28, P3_INSTADDRPOINTER_REG_13__SCAN_IN, P3_ADD_405_U107);
  not ginst20283 (P3_ADD_405_U29, P3_INSTADDRPOINTER_REG_14__SCAN_IN);
  nand ginst20284 (P3_ADD_405_U30, P3_INSTADDRPOINTER_REG_14__SCAN_IN, P3_ADD_405_U108);
  not ginst20285 (P3_ADD_405_U31, P3_INSTADDRPOINTER_REG_15__SCAN_IN);
  nand ginst20286 (P3_ADD_405_U32, P3_INSTADDRPOINTER_REG_15__SCAN_IN, P3_ADD_405_U109);
  not ginst20287 (P3_ADD_405_U33, P3_INSTADDRPOINTER_REG_16__SCAN_IN);
  nand ginst20288 (P3_ADD_405_U34, P3_INSTADDRPOINTER_REG_16__SCAN_IN, P3_ADD_405_U110);
  not ginst20289 (P3_ADD_405_U35, P3_INSTADDRPOINTER_REG_17__SCAN_IN);
  nand ginst20290 (P3_ADD_405_U36, P3_INSTADDRPOINTER_REG_17__SCAN_IN, P3_ADD_405_U111);
  not ginst20291 (P3_ADD_405_U37, P3_INSTADDRPOINTER_REG_18__SCAN_IN);
  nand ginst20292 (P3_ADD_405_U38, P3_INSTADDRPOINTER_REG_18__SCAN_IN, P3_ADD_405_U112);
  not ginst20293 (P3_ADD_405_U39, P3_INSTADDRPOINTER_REG_19__SCAN_IN);
  not ginst20294 (P3_ADD_405_U4, P3_INSTADDRPOINTER_REG_0__SCAN_IN);
  nand ginst20295 (P3_ADD_405_U40, P3_INSTADDRPOINTER_REG_19__SCAN_IN, P3_ADD_405_U113);
  not ginst20296 (P3_ADD_405_U41, P3_INSTADDRPOINTER_REG_20__SCAN_IN);
  nand ginst20297 (P3_ADD_405_U42, P3_INSTADDRPOINTER_REG_20__SCAN_IN, P3_ADD_405_U114);
  not ginst20298 (P3_ADD_405_U43, P3_INSTADDRPOINTER_REG_21__SCAN_IN);
  nand ginst20299 (P3_ADD_405_U44, P3_INSTADDRPOINTER_REG_21__SCAN_IN, P3_ADD_405_U115);
  not ginst20300 (P3_ADD_405_U45, P3_INSTADDRPOINTER_REG_22__SCAN_IN);
  nand ginst20301 (P3_ADD_405_U46, P3_INSTADDRPOINTER_REG_22__SCAN_IN, P3_ADD_405_U116);
  not ginst20302 (P3_ADD_405_U47, P3_INSTADDRPOINTER_REG_23__SCAN_IN);
  nand ginst20303 (P3_ADD_405_U48, P3_INSTADDRPOINTER_REG_23__SCAN_IN, P3_ADD_405_U117);
  not ginst20304 (P3_ADD_405_U49, P3_INSTADDRPOINTER_REG_24__SCAN_IN);
  nand ginst20305 (P3_ADD_405_U5, P3_ADD_405_U126, P3_ADD_405_U92);
  nand ginst20306 (P3_ADD_405_U50, P3_INSTADDRPOINTER_REG_24__SCAN_IN, P3_ADD_405_U118);
  not ginst20307 (P3_ADD_405_U51, P3_INSTADDRPOINTER_REG_25__SCAN_IN);
  nand ginst20308 (P3_ADD_405_U52, P3_INSTADDRPOINTER_REG_25__SCAN_IN, P3_ADD_405_U119);
  not ginst20309 (P3_ADD_405_U53, P3_INSTADDRPOINTER_REG_26__SCAN_IN);
  nand ginst20310 (P3_ADD_405_U54, P3_INSTADDRPOINTER_REG_26__SCAN_IN, P3_ADD_405_U120);
  not ginst20311 (P3_ADD_405_U55, P3_INSTADDRPOINTER_REG_27__SCAN_IN);
  nand ginst20312 (P3_ADD_405_U56, P3_INSTADDRPOINTER_REG_27__SCAN_IN, P3_ADD_405_U121);
  not ginst20313 (P3_ADD_405_U57, P3_INSTADDRPOINTER_REG_28__SCAN_IN);
  nand ginst20314 (P3_ADD_405_U58, P3_INSTADDRPOINTER_REG_28__SCAN_IN, P3_ADD_405_U122);
  not ginst20315 (P3_ADD_405_U59, P3_INSTADDRPOINTER_REG_29__SCAN_IN);
  not ginst20316 (P3_ADD_405_U6, P3_INSTADDRPOINTER_REG_1__SCAN_IN);
  nand ginst20317 (P3_ADD_405_U60, P3_INSTADDRPOINTER_REG_29__SCAN_IN, P3_ADD_405_U123);
  not ginst20318 (P3_ADD_405_U61, P3_INSTADDRPOINTER_REG_30__SCAN_IN);
  not ginst20319 (P3_ADD_405_U62, P3_INSTADDRPOINTER_REG_2__SCAN_IN);
  nand ginst20320 (P3_ADD_405_U63, P3_ADD_405_U127, P3_ADD_405_U128);
  nand ginst20321 (P3_ADD_405_U64, P3_ADD_405_U129, P3_ADD_405_U130);
  nand ginst20322 (P3_ADD_405_U65, P3_ADD_405_U131, P3_ADD_405_U132);
  nand ginst20323 (P3_ADD_405_U66, P3_ADD_405_U133, P3_ADD_405_U134);
  nand ginst20324 (P3_ADD_405_U67, P3_ADD_405_U135, P3_ADD_405_U136);
  nand ginst20325 (P3_ADD_405_U68, P3_ADD_405_U137, P3_ADD_405_U138);
  nand ginst20326 (P3_ADD_405_U69, P3_ADD_405_U141, P3_ADD_405_U142);
  not ginst20327 (P3_ADD_405_U7, P3_INSTADDRPOINTER_REG_3__SCAN_IN);
  nand ginst20328 (P3_ADD_405_U70, P3_ADD_405_U143, P3_ADD_405_U144);
  nand ginst20329 (P3_ADD_405_U71, P3_ADD_405_U145, P3_ADD_405_U146);
  nand ginst20330 (P3_ADD_405_U72, P3_ADD_405_U147, P3_ADD_405_U148);
  nand ginst20331 (P3_ADD_405_U73, P3_ADD_405_U149, P3_ADD_405_U150);
  nand ginst20332 (P3_ADD_405_U74, P3_ADD_405_U151, P3_ADD_405_U152);
  nand ginst20333 (P3_ADD_405_U75, P3_ADD_405_U153, P3_ADD_405_U154);
  nand ginst20334 (P3_ADD_405_U76, P3_ADD_405_U155, P3_ADD_405_U156);
  nand ginst20335 (P3_ADD_405_U77, P3_ADD_405_U157, P3_ADD_405_U158);
  nand ginst20336 (P3_ADD_405_U78, P3_ADD_405_U159, P3_ADD_405_U160);
  nand ginst20337 (P3_ADD_405_U79, P3_ADD_405_U161, P3_ADD_405_U162);
  nand ginst20338 (P3_ADD_405_U8, P3_INSTADDRPOINTER_REG_3__SCAN_IN, P3_ADD_405_U92);
  nand ginst20339 (P3_ADD_405_U80, P3_ADD_405_U163, P3_ADD_405_U164);
  nand ginst20340 (P3_ADD_405_U81, P3_ADD_405_U165, P3_ADD_405_U166);
  nand ginst20341 (P3_ADD_405_U82, P3_ADD_405_U167, P3_ADD_405_U168);
  nand ginst20342 (P3_ADD_405_U83, P3_ADD_405_U169, P3_ADD_405_U170);
  nand ginst20343 (P3_ADD_405_U84, P3_ADD_405_U171, P3_ADD_405_U172);
  nand ginst20344 (P3_ADD_405_U85, P3_ADD_405_U173, P3_ADD_405_U174);
  nand ginst20345 (P3_ADD_405_U86, P3_ADD_405_U175, P3_ADD_405_U176);
  nand ginst20346 (P3_ADD_405_U87, P3_ADD_405_U177, P3_ADD_405_U178);
  nand ginst20347 (P3_ADD_405_U88, P3_ADD_405_U179, P3_ADD_405_U180);
  nand ginst20348 (P3_ADD_405_U89, P3_ADD_405_U181, P3_ADD_405_U182);
  not ginst20349 (P3_ADD_405_U9, P3_INSTADDRPOINTER_REG_4__SCAN_IN);
  nand ginst20350 (P3_ADD_405_U90, P3_ADD_405_U183, P3_ADD_405_U184);
  nand ginst20351 (P3_ADD_405_U91, P3_ADD_405_U185, P3_ADD_405_U186);
  nand ginst20352 (P3_ADD_405_U92, P3_ADD_405_U62, P3_ADD_405_U96);
  and ginst20353 (P3_ADD_405_U93, P3_ADD_405_U139, P3_ADD_405_U140);
  not ginst20354 (P3_ADD_405_U94, P3_INSTADDRPOINTER_REG_31__SCAN_IN);
  nand ginst20355 (P3_ADD_405_U95, P3_INSTADDRPOINTER_REG_30__SCAN_IN, P3_ADD_405_U124);
  nand ginst20356 (P3_ADD_405_U96, P3_INSTADDRPOINTER_REG_0__SCAN_IN, P3_INSTADDRPOINTER_REG_1__SCAN_IN);
  not ginst20357 (P3_ADD_405_U97, P3_ADD_405_U92);
  not ginst20358 (P3_ADD_405_U98, P3_ADD_405_U8);
  not ginst20359 (P3_ADD_405_U99, P3_ADD_405_U10);
  nand ginst20360 (P3_ADD_430_U10, P3_REIP_REG_4__SCAN_IN, P3_ADD_430_U95);
  not ginst20361 (P3_ADD_430_U100, P3_ADD_430_U19);
  not ginst20362 (P3_ADD_430_U101, P3_ADD_430_U20);
  not ginst20363 (P3_ADD_430_U102, P3_ADD_430_U22);
  not ginst20364 (P3_ADD_430_U103, P3_ADD_430_U24);
  not ginst20365 (P3_ADD_430_U104, P3_ADD_430_U26);
  not ginst20366 (P3_ADD_430_U105, P3_ADD_430_U28);
  not ginst20367 (P3_ADD_430_U106, P3_ADD_430_U30);
  not ginst20368 (P3_ADD_430_U107, P3_ADD_430_U32);
  not ginst20369 (P3_ADD_430_U108, P3_ADD_430_U34);
  not ginst20370 (P3_ADD_430_U109, P3_ADD_430_U36);
  not ginst20371 (P3_ADD_430_U11, P3_REIP_REG_5__SCAN_IN);
  not ginst20372 (P3_ADD_430_U110, P3_ADD_430_U38);
  not ginst20373 (P3_ADD_430_U111, P3_ADD_430_U40);
  not ginst20374 (P3_ADD_430_U112, P3_ADD_430_U42);
  not ginst20375 (P3_ADD_430_U113, P3_ADD_430_U44);
  not ginst20376 (P3_ADD_430_U114, P3_ADD_430_U46);
  not ginst20377 (P3_ADD_430_U115, P3_ADD_430_U48);
  not ginst20378 (P3_ADD_430_U116, P3_ADD_430_U50);
  not ginst20379 (P3_ADD_430_U117, P3_ADD_430_U52);
  not ginst20380 (P3_ADD_430_U118, P3_ADD_430_U54);
  not ginst20381 (P3_ADD_430_U119, P3_ADD_430_U56);
  nand ginst20382 (P3_ADD_430_U12, P3_REIP_REG_5__SCAN_IN, P3_ADD_430_U96);
  not ginst20383 (P3_ADD_430_U120, P3_ADD_430_U58);
  not ginst20384 (P3_ADD_430_U121, P3_ADD_430_U60);
  not ginst20385 (P3_ADD_430_U122, P3_ADD_430_U93);
  nand ginst20386 (P3_ADD_430_U123, P3_REIP_REG_9__SCAN_IN, P3_ADD_430_U19);
  nand ginst20387 (P3_ADD_430_U124, P3_ADD_430_U100, P3_ADD_430_U18);
  nand ginst20388 (P3_ADD_430_U125, P3_REIP_REG_8__SCAN_IN, P3_ADD_430_U16);
  nand ginst20389 (P3_ADD_430_U126, P3_ADD_430_U17, P3_ADD_430_U99);
  nand ginst20390 (P3_ADD_430_U127, P3_REIP_REG_7__SCAN_IN, P3_ADD_430_U14);
  nand ginst20391 (P3_ADD_430_U128, P3_ADD_430_U15, P3_ADD_430_U98);
  nand ginst20392 (P3_ADD_430_U129, P3_REIP_REG_6__SCAN_IN, P3_ADD_430_U12);
  not ginst20393 (P3_ADD_430_U13, P3_REIP_REG_6__SCAN_IN);
  nand ginst20394 (P3_ADD_430_U130, P3_ADD_430_U13, P3_ADD_430_U97);
  nand ginst20395 (P3_ADD_430_U131, P3_REIP_REG_5__SCAN_IN, P3_ADD_430_U10);
  nand ginst20396 (P3_ADD_430_U132, P3_ADD_430_U11, P3_ADD_430_U96);
  nand ginst20397 (P3_ADD_430_U133, P3_REIP_REG_4__SCAN_IN, P3_ADD_430_U8);
  nand ginst20398 (P3_ADD_430_U134, P3_ADD_430_U9, P3_ADD_430_U95);
  nand ginst20399 (P3_ADD_430_U135, P3_REIP_REG_3__SCAN_IN, P3_ADD_430_U6);
  nand ginst20400 (P3_ADD_430_U136, P3_ADD_430_U7, P3_ADD_430_U94);
  nand ginst20401 (P3_ADD_430_U137, P3_REIP_REG_31__SCAN_IN, P3_ADD_430_U93);
  nand ginst20402 (P3_ADD_430_U138, P3_ADD_430_U122, P3_ADD_430_U92);
  nand ginst20403 (P3_ADD_430_U139, P3_REIP_REG_30__SCAN_IN, P3_ADD_430_U60);
  nand ginst20404 (P3_ADD_430_U14, P3_REIP_REG_6__SCAN_IN, P3_ADD_430_U97);
  nand ginst20405 (P3_ADD_430_U140, P3_ADD_430_U121, P3_ADD_430_U61);
  nand ginst20406 (P3_ADD_430_U141, P3_REIP_REG_2__SCAN_IN, P3_ADD_430_U4);
  nand ginst20407 (P3_ADD_430_U142, P3_REIP_REG_1__SCAN_IN, P3_ADD_430_U5);
  nand ginst20408 (P3_ADD_430_U143, P3_REIP_REG_29__SCAN_IN, P3_ADD_430_U58);
  nand ginst20409 (P3_ADD_430_U144, P3_ADD_430_U120, P3_ADD_430_U59);
  nand ginst20410 (P3_ADD_430_U145, P3_REIP_REG_28__SCAN_IN, P3_ADD_430_U56);
  nand ginst20411 (P3_ADD_430_U146, P3_ADD_430_U119, P3_ADD_430_U57);
  nand ginst20412 (P3_ADD_430_U147, P3_REIP_REG_27__SCAN_IN, P3_ADD_430_U54);
  nand ginst20413 (P3_ADD_430_U148, P3_ADD_430_U118, P3_ADD_430_U55);
  nand ginst20414 (P3_ADD_430_U149, P3_REIP_REG_26__SCAN_IN, P3_ADD_430_U52);
  not ginst20415 (P3_ADD_430_U15, P3_REIP_REG_7__SCAN_IN);
  nand ginst20416 (P3_ADD_430_U150, P3_ADD_430_U117, P3_ADD_430_U53);
  nand ginst20417 (P3_ADD_430_U151, P3_REIP_REG_25__SCAN_IN, P3_ADD_430_U50);
  nand ginst20418 (P3_ADD_430_U152, P3_ADD_430_U116, P3_ADD_430_U51);
  nand ginst20419 (P3_ADD_430_U153, P3_REIP_REG_24__SCAN_IN, P3_ADD_430_U48);
  nand ginst20420 (P3_ADD_430_U154, P3_ADD_430_U115, P3_ADD_430_U49);
  nand ginst20421 (P3_ADD_430_U155, P3_REIP_REG_23__SCAN_IN, P3_ADD_430_U46);
  nand ginst20422 (P3_ADD_430_U156, P3_ADD_430_U114, P3_ADD_430_U47);
  nand ginst20423 (P3_ADD_430_U157, P3_REIP_REG_22__SCAN_IN, P3_ADD_430_U44);
  nand ginst20424 (P3_ADD_430_U158, P3_ADD_430_U113, P3_ADD_430_U45);
  nand ginst20425 (P3_ADD_430_U159, P3_REIP_REG_21__SCAN_IN, P3_ADD_430_U42);
  nand ginst20426 (P3_ADD_430_U16, P3_REIP_REG_7__SCAN_IN, P3_ADD_430_U98);
  nand ginst20427 (P3_ADD_430_U160, P3_ADD_430_U112, P3_ADD_430_U43);
  nand ginst20428 (P3_ADD_430_U161, P3_REIP_REG_20__SCAN_IN, P3_ADD_430_U40);
  nand ginst20429 (P3_ADD_430_U162, P3_ADD_430_U111, P3_ADD_430_U41);
  nand ginst20430 (P3_ADD_430_U163, P3_REIP_REG_19__SCAN_IN, P3_ADD_430_U38);
  nand ginst20431 (P3_ADD_430_U164, P3_ADD_430_U110, P3_ADD_430_U39);
  nand ginst20432 (P3_ADD_430_U165, P3_REIP_REG_18__SCAN_IN, P3_ADD_430_U36);
  nand ginst20433 (P3_ADD_430_U166, P3_ADD_430_U109, P3_ADD_430_U37);
  nand ginst20434 (P3_ADD_430_U167, P3_REIP_REG_17__SCAN_IN, P3_ADD_430_U34);
  nand ginst20435 (P3_ADD_430_U168, P3_ADD_430_U108, P3_ADD_430_U35);
  nand ginst20436 (P3_ADD_430_U169, P3_REIP_REG_16__SCAN_IN, P3_ADD_430_U32);
  not ginst20437 (P3_ADD_430_U17, P3_REIP_REG_8__SCAN_IN);
  nand ginst20438 (P3_ADD_430_U170, P3_ADD_430_U107, P3_ADD_430_U33);
  nand ginst20439 (P3_ADD_430_U171, P3_REIP_REG_15__SCAN_IN, P3_ADD_430_U30);
  nand ginst20440 (P3_ADD_430_U172, P3_ADD_430_U106, P3_ADD_430_U31);
  nand ginst20441 (P3_ADD_430_U173, P3_REIP_REG_14__SCAN_IN, P3_ADD_430_U28);
  nand ginst20442 (P3_ADD_430_U174, P3_ADD_430_U105, P3_ADD_430_U29);
  nand ginst20443 (P3_ADD_430_U175, P3_REIP_REG_13__SCAN_IN, P3_ADD_430_U26);
  nand ginst20444 (P3_ADD_430_U176, P3_ADD_430_U104, P3_ADD_430_U27);
  nand ginst20445 (P3_ADD_430_U177, P3_REIP_REG_12__SCAN_IN, P3_ADD_430_U24);
  nand ginst20446 (P3_ADD_430_U178, P3_ADD_430_U103, P3_ADD_430_U25);
  nand ginst20447 (P3_ADD_430_U179, P3_REIP_REG_11__SCAN_IN, P3_ADD_430_U22);
  not ginst20448 (P3_ADD_430_U18, P3_REIP_REG_9__SCAN_IN);
  nand ginst20449 (P3_ADD_430_U180, P3_ADD_430_U102, P3_ADD_430_U23);
  nand ginst20450 (P3_ADD_430_U181, P3_REIP_REG_10__SCAN_IN, P3_ADD_430_U20);
  nand ginst20451 (P3_ADD_430_U182, P3_ADD_430_U101, P3_ADD_430_U21);
  nand ginst20452 (P3_ADD_430_U19, P3_REIP_REG_8__SCAN_IN, P3_ADD_430_U99);
  nand ginst20453 (P3_ADD_430_U20, P3_REIP_REG_9__SCAN_IN, P3_ADD_430_U100);
  not ginst20454 (P3_ADD_430_U21, P3_REIP_REG_10__SCAN_IN);
  nand ginst20455 (P3_ADD_430_U22, P3_REIP_REG_10__SCAN_IN, P3_ADD_430_U101);
  not ginst20456 (P3_ADD_430_U23, P3_REIP_REG_11__SCAN_IN);
  nand ginst20457 (P3_ADD_430_U24, P3_REIP_REG_11__SCAN_IN, P3_ADD_430_U102);
  not ginst20458 (P3_ADD_430_U25, P3_REIP_REG_12__SCAN_IN);
  nand ginst20459 (P3_ADD_430_U26, P3_REIP_REG_12__SCAN_IN, P3_ADD_430_U103);
  not ginst20460 (P3_ADD_430_U27, P3_REIP_REG_13__SCAN_IN);
  nand ginst20461 (P3_ADD_430_U28, P3_REIP_REG_13__SCAN_IN, P3_ADD_430_U104);
  not ginst20462 (P3_ADD_430_U29, P3_REIP_REG_14__SCAN_IN);
  nand ginst20463 (P3_ADD_430_U30, P3_REIP_REG_14__SCAN_IN, P3_ADD_430_U105);
  not ginst20464 (P3_ADD_430_U31, P3_REIP_REG_15__SCAN_IN);
  nand ginst20465 (P3_ADD_430_U32, P3_REIP_REG_15__SCAN_IN, P3_ADD_430_U106);
  not ginst20466 (P3_ADD_430_U33, P3_REIP_REG_16__SCAN_IN);
  nand ginst20467 (P3_ADD_430_U34, P3_REIP_REG_16__SCAN_IN, P3_ADD_430_U107);
  not ginst20468 (P3_ADD_430_U35, P3_REIP_REG_17__SCAN_IN);
  nand ginst20469 (P3_ADD_430_U36, P3_REIP_REG_17__SCAN_IN, P3_ADD_430_U108);
  not ginst20470 (P3_ADD_430_U37, P3_REIP_REG_18__SCAN_IN);
  nand ginst20471 (P3_ADD_430_U38, P3_REIP_REG_18__SCAN_IN, P3_ADD_430_U109);
  not ginst20472 (P3_ADD_430_U39, P3_REIP_REG_19__SCAN_IN);
  not ginst20473 (P3_ADD_430_U4, P3_REIP_REG_1__SCAN_IN);
  nand ginst20474 (P3_ADD_430_U40, P3_REIP_REG_19__SCAN_IN, P3_ADD_430_U110);
  not ginst20475 (P3_ADD_430_U41, P3_REIP_REG_20__SCAN_IN);
  nand ginst20476 (P3_ADD_430_U42, P3_REIP_REG_20__SCAN_IN, P3_ADD_430_U111);
  not ginst20477 (P3_ADD_430_U43, P3_REIP_REG_21__SCAN_IN);
  nand ginst20478 (P3_ADD_430_U44, P3_REIP_REG_21__SCAN_IN, P3_ADD_430_U112);
  not ginst20479 (P3_ADD_430_U45, P3_REIP_REG_22__SCAN_IN);
  nand ginst20480 (P3_ADD_430_U46, P3_REIP_REG_22__SCAN_IN, P3_ADD_430_U113);
  not ginst20481 (P3_ADD_430_U47, P3_REIP_REG_23__SCAN_IN);
  nand ginst20482 (P3_ADD_430_U48, P3_REIP_REG_23__SCAN_IN, P3_ADD_430_U114);
  not ginst20483 (P3_ADD_430_U49, P3_REIP_REG_24__SCAN_IN);
  not ginst20484 (P3_ADD_430_U5, P3_REIP_REG_2__SCAN_IN);
  nand ginst20485 (P3_ADD_430_U50, P3_REIP_REG_24__SCAN_IN, P3_ADD_430_U115);
  not ginst20486 (P3_ADD_430_U51, P3_REIP_REG_25__SCAN_IN);
  nand ginst20487 (P3_ADD_430_U52, P3_REIP_REG_25__SCAN_IN, P3_ADD_430_U116);
  not ginst20488 (P3_ADD_430_U53, P3_REIP_REG_26__SCAN_IN);
  nand ginst20489 (P3_ADD_430_U54, P3_REIP_REG_26__SCAN_IN, P3_ADD_430_U117);
  not ginst20490 (P3_ADD_430_U55, P3_REIP_REG_27__SCAN_IN);
  nand ginst20491 (P3_ADD_430_U56, P3_REIP_REG_27__SCAN_IN, P3_ADD_430_U118);
  not ginst20492 (P3_ADD_430_U57, P3_REIP_REG_28__SCAN_IN);
  nand ginst20493 (P3_ADD_430_U58, P3_REIP_REG_28__SCAN_IN, P3_ADD_430_U119);
  not ginst20494 (P3_ADD_430_U59, P3_REIP_REG_29__SCAN_IN);
  nand ginst20495 (P3_ADD_430_U6, P3_REIP_REG_1__SCAN_IN, P3_REIP_REG_2__SCAN_IN);
  nand ginst20496 (P3_ADD_430_U60, P3_REIP_REG_29__SCAN_IN, P3_ADD_430_U120);
  not ginst20497 (P3_ADD_430_U61, P3_REIP_REG_30__SCAN_IN);
  nand ginst20498 (P3_ADD_430_U62, P3_ADD_430_U123, P3_ADD_430_U124);
  nand ginst20499 (P3_ADD_430_U63, P3_ADD_430_U125, P3_ADD_430_U126);
  nand ginst20500 (P3_ADD_430_U64, P3_ADD_430_U127, P3_ADD_430_U128);
  nand ginst20501 (P3_ADD_430_U65, P3_ADD_430_U129, P3_ADD_430_U130);
  nand ginst20502 (P3_ADD_430_U66, P3_ADD_430_U131, P3_ADD_430_U132);
  nand ginst20503 (P3_ADD_430_U67, P3_ADD_430_U133, P3_ADD_430_U134);
  nand ginst20504 (P3_ADD_430_U68, P3_ADD_430_U135, P3_ADD_430_U136);
  nand ginst20505 (P3_ADD_430_U69, P3_ADD_430_U137, P3_ADD_430_U138);
  not ginst20506 (P3_ADD_430_U7, P3_REIP_REG_3__SCAN_IN);
  nand ginst20507 (P3_ADD_430_U70, P3_ADD_430_U139, P3_ADD_430_U140);
  nand ginst20508 (P3_ADD_430_U71, P3_ADD_430_U141, P3_ADD_430_U142);
  nand ginst20509 (P3_ADD_430_U72, P3_ADD_430_U143, P3_ADD_430_U144);
  nand ginst20510 (P3_ADD_430_U73, P3_ADD_430_U145, P3_ADD_430_U146);
  nand ginst20511 (P3_ADD_430_U74, P3_ADD_430_U147, P3_ADD_430_U148);
  nand ginst20512 (P3_ADD_430_U75, P3_ADD_430_U149, P3_ADD_430_U150);
  nand ginst20513 (P3_ADD_430_U76, P3_ADD_430_U151, P3_ADD_430_U152);
  nand ginst20514 (P3_ADD_430_U77, P3_ADD_430_U153, P3_ADD_430_U154);
  nand ginst20515 (P3_ADD_430_U78, P3_ADD_430_U155, P3_ADD_430_U156);
  nand ginst20516 (P3_ADD_430_U79, P3_ADD_430_U157, P3_ADD_430_U158);
  nand ginst20517 (P3_ADD_430_U8, P3_REIP_REG_3__SCAN_IN, P3_ADD_430_U94);
  nand ginst20518 (P3_ADD_430_U80, P3_ADD_430_U159, P3_ADD_430_U160);
  nand ginst20519 (P3_ADD_430_U81, P3_ADD_430_U161, P3_ADD_430_U162);
  nand ginst20520 (P3_ADD_430_U82, P3_ADD_430_U163, P3_ADD_430_U164);
  nand ginst20521 (P3_ADD_430_U83, P3_ADD_430_U165, P3_ADD_430_U166);
  nand ginst20522 (P3_ADD_430_U84, P3_ADD_430_U167, P3_ADD_430_U168);
  nand ginst20523 (P3_ADD_430_U85, P3_ADD_430_U169, P3_ADD_430_U170);
  nand ginst20524 (P3_ADD_430_U86, P3_ADD_430_U171, P3_ADD_430_U172);
  nand ginst20525 (P3_ADD_430_U87, P3_ADD_430_U173, P3_ADD_430_U174);
  nand ginst20526 (P3_ADD_430_U88, P3_ADD_430_U175, P3_ADD_430_U176);
  nand ginst20527 (P3_ADD_430_U89, P3_ADD_430_U177, P3_ADD_430_U178);
  not ginst20528 (P3_ADD_430_U9, P3_REIP_REG_4__SCAN_IN);
  nand ginst20529 (P3_ADD_430_U90, P3_ADD_430_U179, P3_ADD_430_U180);
  nand ginst20530 (P3_ADD_430_U91, P3_ADD_430_U181, P3_ADD_430_U182);
  not ginst20531 (P3_ADD_430_U92, P3_REIP_REG_31__SCAN_IN);
  nand ginst20532 (P3_ADD_430_U93, P3_REIP_REG_30__SCAN_IN, P3_ADD_430_U121);
  not ginst20533 (P3_ADD_430_U94, P3_ADD_430_U6);
  not ginst20534 (P3_ADD_430_U95, P3_ADD_430_U8);
  not ginst20535 (P3_ADD_430_U96, P3_ADD_430_U10);
  not ginst20536 (P3_ADD_430_U97, P3_ADD_430_U12);
  not ginst20537 (P3_ADD_430_U98, P3_ADD_430_U14);
  not ginst20538 (P3_ADD_430_U99, P3_ADD_430_U16);
  nand ginst20539 (P3_ADD_441_U10, P3_INSTADDRPOINTER_REG_4__SCAN_IN, P3_ADD_441_U95);
  not ginst20540 (P3_ADD_441_U100, P3_ADD_441_U19);
  not ginst20541 (P3_ADD_441_U101, P3_ADD_441_U20);
  not ginst20542 (P3_ADD_441_U102, P3_ADD_441_U22);
  not ginst20543 (P3_ADD_441_U103, P3_ADD_441_U24);
  not ginst20544 (P3_ADD_441_U104, P3_ADD_441_U26);
  not ginst20545 (P3_ADD_441_U105, P3_ADD_441_U28);
  not ginst20546 (P3_ADD_441_U106, P3_ADD_441_U30);
  not ginst20547 (P3_ADD_441_U107, P3_ADD_441_U32);
  not ginst20548 (P3_ADD_441_U108, P3_ADD_441_U34);
  not ginst20549 (P3_ADD_441_U109, P3_ADD_441_U36);
  not ginst20550 (P3_ADD_441_U11, P3_INSTADDRPOINTER_REG_5__SCAN_IN);
  not ginst20551 (P3_ADD_441_U110, P3_ADD_441_U38);
  not ginst20552 (P3_ADD_441_U111, P3_ADD_441_U40);
  not ginst20553 (P3_ADD_441_U112, P3_ADD_441_U42);
  not ginst20554 (P3_ADD_441_U113, P3_ADD_441_U44);
  not ginst20555 (P3_ADD_441_U114, P3_ADD_441_U46);
  not ginst20556 (P3_ADD_441_U115, P3_ADD_441_U48);
  not ginst20557 (P3_ADD_441_U116, P3_ADD_441_U50);
  not ginst20558 (P3_ADD_441_U117, P3_ADD_441_U52);
  not ginst20559 (P3_ADD_441_U118, P3_ADD_441_U54);
  not ginst20560 (P3_ADD_441_U119, P3_ADD_441_U56);
  nand ginst20561 (P3_ADD_441_U12, P3_INSTADDRPOINTER_REG_5__SCAN_IN, P3_ADD_441_U96);
  not ginst20562 (P3_ADD_441_U120, P3_ADD_441_U58);
  not ginst20563 (P3_ADD_441_U121, P3_ADD_441_U60);
  not ginst20564 (P3_ADD_441_U122, P3_ADD_441_U93);
  nand ginst20565 (P3_ADD_441_U123, P3_INSTADDRPOINTER_REG_9__SCAN_IN, P3_ADD_441_U19);
  nand ginst20566 (P3_ADD_441_U124, P3_ADD_441_U100, P3_ADD_441_U18);
  nand ginst20567 (P3_ADD_441_U125, P3_INSTADDRPOINTER_REG_8__SCAN_IN, P3_ADD_441_U16);
  nand ginst20568 (P3_ADD_441_U126, P3_ADD_441_U17, P3_ADD_441_U99);
  nand ginst20569 (P3_ADD_441_U127, P3_INSTADDRPOINTER_REG_7__SCAN_IN, P3_ADD_441_U14);
  nand ginst20570 (P3_ADD_441_U128, P3_ADD_441_U15, P3_ADD_441_U98);
  nand ginst20571 (P3_ADD_441_U129, P3_INSTADDRPOINTER_REG_6__SCAN_IN, P3_ADD_441_U12);
  not ginst20572 (P3_ADD_441_U13, P3_INSTADDRPOINTER_REG_6__SCAN_IN);
  nand ginst20573 (P3_ADD_441_U130, P3_ADD_441_U13, P3_ADD_441_U97);
  nand ginst20574 (P3_ADD_441_U131, P3_INSTADDRPOINTER_REG_5__SCAN_IN, P3_ADD_441_U10);
  nand ginst20575 (P3_ADD_441_U132, P3_ADD_441_U11, P3_ADD_441_U96);
  nand ginst20576 (P3_ADD_441_U133, P3_INSTADDRPOINTER_REG_4__SCAN_IN, P3_ADD_441_U8);
  nand ginst20577 (P3_ADD_441_U134, P3_ADD_441_U9, P3_ADD_441_U95);
  nand ginst20578 (P3_ADD_441_U135, P3_INSTADDRPOINTER_REG_3__SCAN_IN, P3_ADD_441_U6);
  nand ginst20579 (P3_ADD_441_U136, P3_ADD_441_U7, P3_ADD_441_U94);
  nand ginst20580 (P3_ADD_441_U137, P3_INSTADDRPOINTER_REG_31__SCAN_IN, P3_ADD_441_U93);
  nand ginst20581 (P3_ADD_441_U138, P3_ADD_441_U122, P3_ADD_441_U92);
  nand ginst20582 (P3_ADD_441_U139, P3_INSTADDRPOINTER_REG_30__SCAN_IN, P3_ADD_441_U60);
  nand ginst20583 (P3_ADD_441_U14, P3_INSTADDRPOINTER_REG_6__SCAN_IN, P3_ADD_441_U97);
  nand ginst20584 (P3_ADD_441_U140, P3_ADD_441_U121, P3_ADD_441_U61);
  nand ginst20585 (P3_ADD_441_U141, P3_INSTADDRPOINTER_REG_2__SCAN_IN, P3_ADD_441_U4);
  nand ginst20586 (P3_ADD_441_U142, P3_INSTADDRPOINTER_REG_1__SCAN_IN, P3_ADD_441_U5);
  nand ginst20587 (P3_ADD_441_U143, P3_INSTADDRPOINTER_REG_29__SCAN_IN, P3_ADD_441_U58);
  nand ginst20588 (P3_ADD_441_U144, P3_ADD_441_U120, P3_ADD_441_U59);
  nand ginst20589 (P3_ADD_441_U145, P3_INSTADDRPOINTER_REG_28__SCAN_IN, P3_ADD_441_U56);
  nand ginst20590 (P3_ADD_441_U146, P3_ADD_441_U119, P3_ADD_441_U57);
  nand ginst20591 (P3_ADD_441_U147, P3_INSTADDRPOINTER_REG_27__SCAN_IN, P3_ADD_441_U54);
  nand ginst20592 (P3_ADD_441_U148, P3_ADD_441_U118, P3_ADD_441_U55);
  nand ginst20593 (P3_ADD_441_U149, P3_INSTADDRPOINTER_REG_26__SCAN_IN, P3_ADD_441_U52);
  not ginst20594 (P3_ADD_441_U15, P3_INSTADDRPOINTER_REG_7__SCAN_IN);
  nand ginst20595 (P3_ADD_441_U150, P3_ADD_441_U117, P3_ADD_441_U53);
  nand ginst20596 (P3_ADD_441_U151, P3_INSTADDRPOINTER_REG_25__SCAN_IN, P3_ADD_441_U50);
  nand ginst20597 (P3_ADD_441_U152, P3_ADD_441_U116, P3_ADD_441_U51);
  nand ginst20598 (P3_ADD_441_U153, P3_INSTADDRPOINTER_REG_24__SCAN_IN, P3_ADD_441_U48);
  nand ginst20599 (P3_ADD_441_U154, P3_ADD_441_U115, P3_ADD_441_U49);
  nand ginst20600 (P3_ADD_441_U155, P3_INSTADDRPOINTER_REG_23__SCAN_IN, P3_ADD_441_U46);
  nand ginst20601 (P3_ADD_441_U156, P3_ADD_441_U114, P3_ADD_441_U47);
  nand ginst20602 (P3_ADD_441_U157, P3_INSTADDRPOINTER_REG_22__SCAN_IN, P3_ADD_441_U44);
  nand ginst20603 (P3_ADD_441_U158, P3_ADD_441_U113, P3_ADD_441_U45);
  nand ginst20604 (P3_ADD_441_U159, P3_INSTADDRPOINTER_REG_21__SCAN_IN, P3_ADD_441_U42);
  nand ginst20605 (P3_ADD_441_U16, P3_INSTADDRPOINTER_REG_7__SCAN_IN, P3_ADD_441_U98);
  nand ginst20606 (P3_ADD_441_U160, P3_ADD_441_U112, P3_ADD_441_U43);
  nand ginst20607 (P3_ADD_441_U161, P3_INSTADDRPOINTER_REG_20__SCAN_IN, P3_ADD_441_U40);
  nand ginst20608 (P3_ADD_441_U162, P3_ADD_441_U111, P3_ADD_441_U41);
  nand ginst20609 (P3_ADD_441_U163, P3_INSTADDRPOINTER_REG_19__SCAN_IN, P3_ADD_441_U38);
  nand ginst20610 (P3_ADD_441_U164, P3_ADD_441_U110, P3_ADD_441_U39);
  nand ginst20611 (P3_ADD_441_U165, P3_INSTADDRPOINTER_REG_18__SCAN_IN, P3_ADD_441_U36);
  nand ginst20612 (P3_ADD_441_U166, P3_ADD_441_U109, P3_ADD_441_U37);
  nand ginst20613 (P3_ADD_441_U167, P3_INSTADDRPOINTER_REG_17__SCAN_IN, P3_ADD_441_U34);
  nand ginst20614 (P3_ADD_441_U168, P3_ADD_441_U108, P3_ADD_441_U35);
  nand ginst20615 (P3_ADD_441_U169, P3_INSTADDRPOINTER_REG_16__SCAN_IN, P3_ADD_441_U32);
  not ginst20616 (P3_ADD_441_U17, P3_INSTADDRPOINTER_REG_8__SCAN_IN);
  nand ginst20617 (P3_ADD_441_U170, P3_ADD_441_U107, P3_ADD_441_U33);
  nand ginst20618 (P3_ADD_441_U171, P3_INSTADDRPOINTER_REG_15__SCAN_IN, P3_ADD_441_U30);
  nand ginst20619 (P3_ADD_441_U172, P3_ADD_441_U106, P3_ADD_441_U31);
  nand ginst20620 (P3_ADD_441_U173, P3_INSTADDRPOINTER_REG_14__SCAN_IN, P3_ADD_441_U28);
  nand ginst20621 (P3_ADD_441_U174, P3_ADD_441_U105, P3_ADD_441_U29);
  nand ginst20622 (P3_ADD_441_U175, P3_INSTADDRPOINTER_REG_13__SCAN_IN, P3_ADD_441_U26);
  nand ginst20623 (P3_ADD_441_U176, P3_ADD_441_U104, P3_ADD_441_U27);
  nand ginst20624 (P3_ADD_441_U177, P3_INSTADDRPOINTER_REG_12__SCAN_IN, P3_ADD_441_U24);
  nand ginst20625 (P3_ADD_441_U178, P3_ADD_441_U103, P3_ADD_441_U25);
  nand ginst20626 (P3_ADD_441_U179, P3_INSTADDRPOINTER_REG_11__SCAN_IN, P3_ADD_441_U22);
  not ginst20627 (P3_ADD_441_U18, P3_INSTADDRPOINTER_REG_9__SCAN_IN);
  nand ginst20628 (P3_ADD_441_U180, P3_ADD_441_U102, P3_ADD_441_U23);
  nand ginst20629 (P3_ADD_441_U181, P3_INSTADDRPOINTER_REG_10__SCAN_IN, P3_ADD_441_U20);
  nand ginst20630 (P3_ADD_441_U182, P3_ADD_441_U101, P3_ADD_441_U21);
  nand ginst20631 (P3_ADD_441_U19, P3_INSTADDRPOINTER_REG_8__SCAN_IN, P3_ADD_441_U99);
  nand ginst20632 (P3_ADD_441_U20, P3_INSTADDRPOINTER_REG_9__SCAN_IN, P3_ADD_441_U100);
  not ginst20633 (P3_ADD_441_U21, P3_INSTADDRPOINTER_REG_10__SCAN_IN);
  nand ginst20634 (P3_ADD_441_U22, P3_INSTADDRPOINTER_REG_10__SCAN_IN, P3_ADD_441_U101);
  not ginst20635 (P3_ADD_441_U23, P3_INSTADDRPOINTER_REG_11__SCAN_IN);
  nand ginst20636 (P3_ADD_441_U24, P3_INSTADDRPOINTER_REG_11__SCAN_IN, P3_ADD_441_U102);
  not ginst20637 (P3_ADD_441_U25, P3_INSTADDRPOINTER_REG_12__SCAN_IN);
  nand ginst20638 (P3_ADD_441_U26, P3_INSTADDRPOINTER_REG_12__SCAN_IN, P3_ADD_441_U103);
  not ginst20639 (P3_ADD_441_U27, P3_INSTADDRPOINTER_REG_13__SCAN_IN);
  nand ginst20640 (P3_ADD_441_U28, P3_INSTADDRPOINTER_REG_13__SCAN_IN, P3_ADD_441_U104);
  not ginst20641 (P3_ADD_441_U29, P3_INSTADDRPOINTER_REG_14__SCAN_IN);
  nand ginst20642 (P3_ADD_441_U30, P3_INSTADDRPOINTER_REG_14__SCAN_IN, P3_ADD_441_U105);
  not ginst20643 (P3_ADD_441_U31, P3_INSTADDRPOINTER_REG_15__SCAN_IN);
  nand ginst20644 (P3_ADD_441_U32, P3_INSTADDRPOINTER_REG_15__SCAN_IN, P3_ADD_441_U106);
  not ginst20645 (P3_ADD_441_U33, P3_INSTADDRPOINTER_REG_16__SCAN_IN);
  nand ginst20646 (P3_ADD_441_U34, P3_INSTADDRPOINTER_REG_16__SCAN_IN, P3_ADD_441_U107);
  not ginst20647 (P3_ADD_441_U35, P3_INSTADDRPOINTER_REG_17__SCAN_IN);
  nand ginst20648 (P3_ADD_441_U36, P3_INSTADDRPOINTER_REG_17__SCAN_IN, P3_ADD_441_U108);
  not ginst20649 (P3_ADD_441_U37, P3_INSTADDRPOINTER_REG_18__SCAN_IN);
  nand ginst20650 (P3_ADD_441_U38, P3_INSTADDRPOINTER_REG_18__SCAN_IN, P3_ADD_441_U109);
  not ginst20651 (P3_ADD_441_U39, P3_INSTADDRPOINTER_REG_19__SCAN_IN);
  not ginst20652 (P3_ADD_441_U4, P3_INSTADDRPOINTER_REG_1__SCAN_IN);
  nand ginst20653 (P3_ADD_441_U40, P3_INSTADDRPOINTER_REG_19__SCAN_IN, P3_ADD_441_U110);
  not ginst20654 (P3_ADD_441_U41, P3_INSTADDRPOINTER_REG_20__SCAN_IN);
  nand ginst20655 (P3_ADD_441_U42, P3_INSTADDRPOINTER_REG_20__SCAN_IN, P3_ADD_441_U111);
  not ginst20656 (P3_ADD_441_U43, P3_INSTADDRPOINTER_REG_21__SCAN_IN);
  nand ginst20657 (P3_ADD_441_U44, P3_INSTADDRPOINTER_REG_21__SCAN_IN, P3_ADD_441_U112);
  not ginst20658 (P3_ADD_441_U45, P3_INSTADDRPOINTER_REG_22__SCAN_IN);
  nand ginst20659 (P3_ADD_441_U46, P3_INSTADDRPOINTER_REG_22__SCAN_IN, P3_ADD_441_U113);
  not ginst20660 (P3_ADD_441_U47, P3_INSTADDRPOINTER_REG_23__SCAN_IN);
  nand ginst20661 (P3_ADD_441_U48, P3_INSTADDRPOINTER_REG_23__SCAN_IN, P3_ADD_441_U114);
  not ginst20662 (P3_ADD_441_U49, P3_INSTADDRPOINTER_REG_24__SCAN_IN);
  not ginst20663 (P3_ADD_441_U5, P3_INSTADDRPOINTER_REG_2__SCAN_IN);
  nand ginst20664 (P3_ADD_441_U50, P3_INSTADDRPOINTER_REG_24__SCAN_IN, P3_ADD_441_U115);
  not ginst20665 (P3_ADD_441_U51, P3_INSTADDRPOINTER_REG_25__SCAN_IN);
  nand ginst20666 (P3_ADD_441_U52, P3_INSTADDRPOINTER_REG_25__SCAN_IN, P3_ADD_441_U116);
  not ginst20667 (P3_ADD_441_U53, P3_INSTADDRPOINTER_REG_26__SCAN_IN);
  nand ginst20668 (P3_ADD_441_U54, P3_INSTADDRPOINTER_REG_26__SCAN_IN, P3_ADD_441_U117);
  not ginst20669 (P3_ADD_441_U55, P3_INSTADDRPOINTER_REG_27__SCAN_IN);
  nand ginst20670 (P3_ADD_441_U56, P3_INSTADDRPOINTER_REG_27__SCAN_IN, P3_ADD_441_U118);
  not ginst20671 (P3_ADD_441_U57, P3_INSTADDRPOINTER_REG_28__SCAN_IN);
  nand ginst20672 (P3_ADD_441_U58, P3_INSTADDRPOINTER_REG_28__SCAN_IN, P3_ADD_441_U119);
  not ginst20673 (P3_ADD_441_U59, P3_INSTADDRPOINTER_REG_29__SCAN_IN);
  nand ginst20674 (P3_ADD_441_U6, P3_INSTADDRPOINTER_REG_1__SCAN_IN, P3_INSTADDRPOINTER_REG_2__SCAN_IN);
  nand ginst20675 (P3_ADD_441_U60, P3_INSTADDRPOINTER_REG_29__SCAN_IN, P3_ADD_441_U120);
  not ginst20676 (P3_ADD_441_U61, P3_INSTADDRPOINTER_REG_30__SCAN_IN);
  nand ginst20677 (P3_ADD_441_U62, P3_ADD_441_U123, P3_ADD_441_U124);
  nand ginst20678 (P3_ADD_441_U63, P3_ADD_441_U125, P3_ADD_441_U126);
  nand ginst20679 (P3_ADD_441_U64, P3_ADD_441_U127, P3_ADD_441_U128);
  nand ginst20680 (P3_ADD_441_U65, P3_ADD_441_U129, P3_ADD_441_U130);
  nand ginst20681 (P3_ADD_441_U66, P3_ADD_441_U131, P3_ADD_441_U132);
  nand ginst20682 (P3_ADD_441_U67, P3_ADD_441_U133, P3_ADD_441_U134);
  nand ginst20683 (P3_ADD_441_U68, P3_ADD_441_U135, P3_ADD_441_U136);
  nand ginst20684 (P3_ADD_441_U69, P3_ADD_441_U137, P3_ADD_441_U138);
  not ginst20685 (P3_ADD_441_U7, P3_INSTADDRPOINTER_REG_3__SCAN_IN);
  nand ginst20686 (P3_ADD_441_U70, P3_ADD_441_U139, P3_ADD_441_U140);
  nand ginst20687 (P3_ADD_441_U71, P3_ADD_441_U141, P3_ADD_441_U142);
  nand ginst20688 (P3_ADD_441_U72, P3_ADD_441_U143, P3_ADD_441_U144);
  nand ginst20689 (P3_ADD_441_U73, P3_ADD_441_U145, P3_ADD_441_U146);
  nand ginst20690 (P3_ADD_441_U74, P3_ADD_441_U147, P3_ADD_441_U148);
  nand ginst20691 (P3_ADD_441_U75, P3_ADD_441_U149, P3_ADD_441_U150);
  nand ginst20692 (P3_ADD_441_U76, P3_ADD_441_U151, P3_ADD_441_U152);
  nand ginst20693 (P3_ADD_441_U77, P3_ADD_441_U153, P3_ADD_441_U154);
  nand ginst20694 (P3_ADD_441_U78, P3_ADD_441_U155, P3_ADD_441_U156);
  nand ginst20695 (P3_ADD_441_U79, P3_ADD_441_U157, P3_ADD_441_U158);
  nand ginst20696 (P3_ADD_441_U8, P3_INSTADDRPOINTER_REG_3__SCAN_IN, P3_ADD_441_U94);
  nand ginst20697 (P3_ADD_441_U80, P3_ADD_441_U159, P3_ADD_441_U160);
  nand ginst20698 (P3_ADD_441_U81, P3_ADD_441_U161, P3_ADD_441_U162);
  nand ginst20699 (P3_ADD_441_U82, P3_ADD_441_U163, P3_ADD_441_U164);
  nand ginst20700 (P3_ADD_441_U83, P3_ADD_441_U165, P3_ADD_441_U166);
  nand ginst20701 (P3_ADD_441_U84, P3_ADD_441_U167, P3_ADD_441_U168);
  nand ginst20702 (P3_ADD_441_U85, P3_ADD_441_U169, P3_ADD_441_U170);
  nand ginst20703 (P3_ADD_441_U86, P3_ADD_441_U171, P3_ADD_441_U172);
  nand ginst20704 (P3_ADD_441_U87, P3_ADD_441_U173, P3_ADD_441_U174);
  nand ginst20705 (P3_ADD_441_U88, P3_ADD_441_U175, P3_ADD_441_U176);
  nand ginst20706 (P3_ADD_441_U89, P3_ADD_441_U177, P3_ADD_441_U178);
  not ginst20707 (P3_ADD_441_U9, P3_INSTADDRPOINTER_REG_4__SCAN_IN);
  nand ginst20708 (P3_ADD_441_U90, P3_ADD_441_U179, P3_ADD_441_U180);
  nand ginst20709 (P3_ADD_441_U91, P3_ADD_441_U181, P3_ADD_441_U182);
  not ginst20710 (P3_ADD_441_U92, P3_INSTADDRPOINTER_REG_31__SCAN_IN);
  nand ginst20711 (P3_ADD_441_U93, P3_INSTADDRPOINTER_REG_30__SCAN_IN, P3_ADD_441_U121);
  not ginst20712 (P3_ADD_441_U94, P3_ADD_441_U6);
  not ginst20713 (P3_ADD_441_U95, P3_ADD_441_U8);
  not ginst20714 (P3_ADD_441_U96, P3_ADD_441_U10);
  not ginst20715 (P3_ADD_441_U97, P3_ADD_441_U12);
  not ginst20716 (P3_ADD_441_U98, P3_ADD_441_U14);
  not ginst20717 (P3_ADD_441_U99, P3_ADD_441_U16);
  nand ginst20718 (P3_ADD_467_U10, P3_REIP_REG_4__SCAN_IN, P3_ADD_467_U95);
  not ginst20719 (P3_ADD_467_U100, P3_ADD_467_U19);
  not ginst20720 (P3_ADD_467_U101, P3_ADD_467_U20);
  not ginst20721 (P3_ADD_467_U102, P3_ADD_467_U22);
  not ginst20722 (P3_ADD_467_U103, P3_ADD_467_U24);
  not ginst20723 (P3_ADD_467_U104, P3_ADD_467_U26);
  not ginst20724 (P3_ADD_467_U105, P3_ADD_467_U28);
  not ginst20725 (P3_ADD_467_U106, P3_ADD_467_U30);
  not ginst20726 (P3_ADD_467_U107, P3_ADD_467_U32);
  not ginst20727 (P3_ADD_467_U108, P3_ADD_467_U34);
  not ginst20728 (P3_ADD_467_U109, P3_ADD_467_U36);
  not ginst20729 (P3_ADD_467_U11, P3_REIP_REG_5__SCAN_IN);
  not ginst20730 (P3_ADD_467_U110, P3_ADD_467_U38);
  not ginst20731 (P3_ADD_467_U111, P3_ADD_467_U40);
  not ginst20732 (P3_ADD_467_U112, P3_ADD_467_U42);
  not ginst20733 (P3_ADD_467_U113, P3_ADD_467_U44);
  not ginst20734 (P3_ADD_467_U114, P3_ADD_467_U46);
  not ginst20735 (P3_ADD_467_U115, P3_ADD_467_U48);
  not ginst20736 (P3_ADD_467_U116, P3_ADD_467_U50);
  not ginst20737 (P3_ADD_467_U117, P3_ADD_467_U52);
  not ginst20738 (P3_ADD_467_U118, P3_ADD_467_U54);
  not ginst20739 (P3_ADD_467_U119, P3_ADD_467_U56);
  nand ginst20740 (P3_ADD_467_U12, P3_REIP_REG_5__SCAN_IN, P3_ADD_467_U96);
  not ginst20741 (P3_ADD_467_U120, P3_ADD_467_U58);
  not ginst20742 (P3_ADD_467_U121, P3_ADD_467_U60);
  not ginst20743 (P3_ADD_467_U122, P3_ADD_467_U93);
  nand ginst20744 (P3_ADD_467_U123, P3_REIP_REG_9__SCAN_IN, P3_ADD_467_U19);
  nand ginst20745 (P3_ADD_467_U124, P3_ADD_467_U100, P3_ADD_467_U18);
  nand ginst20746 (P3_ADD_467_U125, P3_REIP_REG_8__SCAN_IN, P3_ADD_467_U16);
  nand ginst20747 (P3_ADD_467_U126, P3_ADD_467_U17, P3_ADD_467_U99);
  nand ginst20748 (P3_ADD_467_U127, P3_REIP_REG_7__SCAN_IN, P3_ADD_467_U14);
  nand ginst20749 (P3_ADD_467_U128, P3_ADD_467_U15, P3_ADD_467_U98);
  nand ginst20750 (P3_ADD_467_U129, P3_REIP_REG_6__SCAN_IN, P3_ADD_467_U12);
  not ginst20751 (P3_ADD_467_U13, P3_REIP_REG_6__SCAN_IN);
  nand ginst20752 (P3_ADD_467_U130, P3_ADD_467_U13, P3_ADD_467_U97);
  nand ginst20753 (P3_ADD_467_U131, P3_REIP_REG_5__SCAN_IN, P3_ADD_467_U10);
  nand ginst20754 (P3_ADD_467_U132, P3_ADD_467_U11, P3_ADD_467_U96);
  nand ginst20755 (P3_ADD_467_U133, P3_REIP_REG_4__SCAN_IN, P3_ADD_467_U8);
  nand ginst20756 (P3_ADD_467_U134, P3_ADD_467_U9, P3_ADD_467_U95);
  nand ginst20757 (P3_ADD_467_U135, P3_REIP_REG_3__SCAN_IN, P3_ADD_467_U6);
  nand ginst20758 (P3_ADD_467_U136, P3_ADD_467_U7, P3_ADD_467_U94);
  nand ginst20759 (P3_ADD_467_U137, P3_REIP_REG_31__SCAN_IN, P3_ADD_467_U93);
  nand ginst20760 (P3_ADD_467_U138, P3_ADD_467_U122, P3_ADD_467_U92);
  nand ginst20761 (P3_ADD_467_U139, P3_REIP_REG_30__SCAN_IN, P3_ADD_467_U60);
  nand ginst20762 (P3_ADD_467_U14, P3_REIP_REG_6__SCAN_IN, P3_ADD_467_U97);
  nand ginst20763 (P3_ADD_467_U140, P3_ADD_467_U121, P3_ADD_467_U61);
  nand ginst20764 (P3_ADD_467_U141, P3_REIP_REG_2__SCAN_IN, P3_ADD_467_U4);
  nand ginst20765 (P3_ADD_467_U142, P3_REIP_REG_1__SCAN_IN, P3_ADD_467_U5);
  nand ginst20766 (P3_ADD_467_U143, P3_REIP_REG_29__SCAN_IN, P3_ADD_467_U58);
  nand ginst20767 (P3_ADD_467_U144, P3_ADD_467_U120, P3_ADD_467_U59);
  nand ginst20768 (P3_ADD_467_U145, P3_REIP_REG_28__SCAN_IN, P3_ADD_467_U56);
  nand ginst20769 (P3_ADD_467_U146, P3_ADD_467_U119, P3_ADD_467_U57);
  nand ginst20770 (P3_ADD_467_U147, P3_REIP_REG_27__SCAN_IN, P3_ADD_467_U54);
  nand ginst20771 (P3_ADD_467_U148, P3_ADD_467_U118, P3_ADD_467_U55);
  nand ginst20772 (P3_ADD_467_U149, P3_REIP_REG_26__SCAN_IN, P3_ADD_467_U52);
  not ginst20773 (P3_ADD_467_U15, P3_REIP_REG_7__SCAN_IN);
  nand ginst20774 (P3_ADD_467_U150, P3_ADD_467_U117, P3_ADD_467_U53);
  nand ginst20775 (P3_ADD_467_U151, P3_REIP_REG_25__SCAN_IN, P3_ADD_467_U50);
  nand ginst20776 (P3_ADD_467_U152, P3_ADD_467_U116, P3_ADD_467_U51);
  nand ginst20777 (P3_ADD_467_U153, P3_REIP_REG_24__SCAN_IN, P3_ADD_467_U48);
  nand ginst20778 (P3_ADD_467_U154, P3_ADD_467_U115, P3_ADD_467_U49);
  nand ginst20779 (P3_ADD_467_U155, P3_REIP_REG_23__SCAN_IN, P3_ADD_467_U46);
  nand ginst20780 (P3_ADD_467_U156, P3_ADD_467_U114, P3_ADD_467_U47);
  nand ginst20781 (P3_ADD_467_U157, P3_REIP_REG_22__SCAN_IN, P3_ADD_467_U44);
  nand ginst20782 (P3_ADD_467_U158, P3_ADD_467_U113, P3_ADD_467_U45);
  nand ginst20783 (P3_ADD_467_U159, P3_REIP_REG_21__SCAN_IN, P3_ADD_467_U42);
  nand ginst20784 (P3_ADD_467_U16, P3_REIP_REG_7__SCAN_IN, P3_ADD_467_U98);
  nand ginst20785 (P3_ADD_467_U160, P3_ADD_467_U112, P3_ADD_467_U43);
  nand ginst20786 (P3_ADD_467_U161, P3_REIP_REG_20__SCAN_IN, P3_ADD_467_U40);
  nand ginst20787 (P3_ADD_467_U162, P3_ADD_467_U111, P3_ADD_467_U41);
  nand ginst20788 (P3_ADD_467_U163, P3_REIP_REG_19__SCAN_IN, P3_ADD_467_U38);
  nand ginst20789 (P3_ADD_467_U164, P3_ADD_467_U110, P3_ADD_467_U39);
  nand ginst20790 (P3_ADD_467_U165, P3_REIP_REG_18__SCAN_IN, P3_ADD_467_U36);
  nand ginst20791 (P3_ADD_467_U166, P3_ADD_467_U109, P3_ADD_467_U37);
  nand ginst20792 (P3_ADD_467_U167, P3_REIP_REG_17__SCAN_IN, P3_ADD_467_U34);
  nand ginst20793 (P3_ADD_467_U168, P3_ADD_467_U108, P3_ADD_467_U35);
  nand ginst20794 (P3_ADD_467_U169, P3_REIP_REG_16__SCAN_IN, P3_ADD_467_U32);
  not ginst20795 (P3_ADD_467_U17, P3_REIP_REG_8__SCAN_IN);
  nand ginst20796 (P3_ADD_467_U170, P3_ADD_467_U107, P3_ADD_467_U33);
  nand ginst20797 (P3_ADD_467_U171, P3_REIP_REG_15__SCAN_IN, P3_ADD_467_U30);
  nand ginst20798 (P3_ADD_467_U172, P3_ADD_467_U106, P3_ADD_467_U31);
  nand ginst20799 (P3_ADD_467_U173, P3_REIP_REG_14__SCAN_IN, P3_ADD_467_U28);
  nand ginst20800 (P3_ADD_467_U174, P3_ADD_467_U105, P3_ADD_467_U29);
  nand ginst20801 (P3_ADD_467_U175, P3_REIP_REG_13__SCAN_IN, P3_ADD_467_U26);
  nand ginst20802 (P3_ADD_467_U176, P3_ADD_467_U104, P3_ADD_467_U27);
  nand ginst20803 (P3_ADD_467_U177, P3_REIP_REG_12__SCAN_IN, P3_ADD_467_U24);
  nand ginst20804 (P3_ADD_467_U178, P3_ADD_467_U103, P3_ADD_467_U25);
  nand ginst20805 (P3_ADD_467_U179, P3_REIP_REG_11__SCAN_IN, P3_ADD_467_U22);
  not ginst20806 (P3_ADD_467_U18, P3_REIP_REG_9__SCAN_IN);
  nand ginst20807 (P3_ADD_467_U180, P3_ADD_467_U102, P3_ADD_467_U23);
  nand ginst20808 (P3_ADD_467_U181, P3_REIP_REG_10__SCAN_IN, P3_ADD_467_U20);
  nand ginst20809 (P3_ADD_467_U182, P3_ADD_467_U101, P3_ADD_467_U21);
  nand ginst20810 (P3_ADD_467_U19, P3_REIP_REG_8__SCAN_IN, P3_ADD_467_U99);
  nand ginst20811 (P3_ADD_467_U20, P3_REIP_REG_9__SCAN_IN, P3_ADD_467_U100);
  not ginst20812 (P3_ADD_467_U21, P3_REIP_REG_10__SCAN_IN);
  nand ginst20813 (P3_ADD_467_U22, P3_REIP_REG_10__SCAN_IN, P3_ADD_467_U101);
  not ginst20814 (P3_ADD_467_U23, P3_REIP_REG_11__SCAN_IN);
  nand ginst20815 (P3_ADD_467_U24, P3_REIP_REG_11__SCAN_IN, P3_ADD_467_U102);
  not ginst20816 (P3_ADD_467_U25, P3_REIP_REG_12__SCAN_IN);
  nand ginst20817 (P3_ADD_467_U26, P3_REIP_REG_12__SCAN_IN, P3_ADD_467_U103);
  not ginst20818 (P3_ADD_467_U27, P3_REIP_REG_13__SCAN_IN);
  nand ginst20819 (P3_ADD_467_U28, P3_REIP_REG_13__SCAN_IN, P3_ADD_467_U104);
  not ginst20820 (P3_ADD_467_U29, P3_REIP_REG_14__SCAN_IN);
  nand ginst20821 (P3_ADD_467_U30, P3_REIP_REG_14__SCAN_IN, P3_ADD_467_U105);
  not ginst20822 (P3_ADD_467_U31, P3_REIP_REG_15__SCAN_IN);
  nand ginst20823 (P3_ADD_467_U32, P3_REIP_REG_15__SCAN_IN, P3_ADD_467_U106);
  not ginst20824 (P3_ADD_467_U33, P3_REIP_REG_16__SCAN_IN);
  nand ginst20825 (P3_ADD_467_U34, P3_REIP_REG_16__SCAN_IN, P3_ADD_467_U107);
  not ginst20826 (P3_ADD_467_U35, P3_REIP_REG_17__SCAN_IN);
  nand ginst20827 (P3_ADD_467_U36, P3_REIP_REG_17__SCAN_IN, P3_ADD_467_U108);
  not ginst20828 (P3_ADD_467_U37, P3_REIP_REG_18__SCAN_IN);
  nand ginst20829 (P3_ADD_467_U38, P3_REIP_REG_18__SCAN_IN, P3_ADD_467_U109);
  not ginst20830 (P3_ADD_467_U39, P3_REIP_REG_19__SCAN_IN);
  not ginst20831 (P3_ADD_467_U4, P3_REIP_REG_1__SCAN_IN);
  nand ginst20832 (P3_ADD_467_U40, P3_REIP_REG_19__SCAN_IN, P3_ADD_467_U110);
  not ginst20833 (P3_ADD_467_U41, P3_REIP_REG_20__SCAN_IN);
  nand ginst20834 (P3_ADD_467_U42, P3_REIP_REG_20__SCAN_IN, P3_ADD_467_U111);
  not ginst20835 (P3_ADD_467_U43, P3_REIP_REG_21__SCAN_IN);
  nand ginst20836 (P3_ADD_467_U44, P3_REIP_REG_21__SCAN_IN, P3_ADD_467_U112);
  not ginst20837 (P3_ADD_467_U45, P3_REIP_REG_22__SCAN_IN);
  nand ginst20838 (P3_ADD_467_U46, P3_REIP_REG_22__SCAN_IN, P3_ADD_467_U113);
  not ginst20839 (P3_ADD_467_U47, P3_REIP_REG_23__SCAN_IN);
  nand ginst20840 (P3_ADD_467_U48, P3_REIP_REG_23__SCAN_IN, P3_ADD_467_U114);
  not ginst20841 (P3_ADD_467_U49, P3_REIP_REG_24__SCAN_IN);
  not ginst20842 (P3_ADD_467_U5, P3_REIP_REG_2__SCAN_IN);
  nand ginst20843 (P3_ADD_467_U50, P3_REIP_REG_24__SCAN_IN, P3_ADD_467_U115);
  not ginst20844 (P3_ADD_467_U51, P3_REIP_REG_25__SCAN_IN);
  nand ginst20845 (P3_ADD_467_U52, P3_REIP_REG_25__SCAN_IN, P3_ADD_467_U116);
  not ginst20846 (P3_ADD_467_U53, P3_REIP_REG_26__SCAN_IN);
  nand ginst20847 (P3_ADD_467_U54, P3_REIP_REG_26__SCAN_IN, P3_ADD_467_U117);
  not ginst20848 (P3_ADD_467_U55, P3_REIP_REG_27__SCAN_IN);
  nand ginst20849 (P3_ADD_467_U56, P3_REIP_REG_27__SCAN_IN, P3_ADD_467_U118);
  not ginst20850 (P3_ADD_467_U57, P3_REIP_REG_28__SCAN_IN);
  nand ginst20851 (P3_ADD_467_U58, P3_REIP_REG_28__SCAN_IN, P3_ADD_467_U119);
  not ginst20852 (P3_ADD_467_U59, P3_REIP_REG_29__SCAN_IN);
  nand ginst20853 (P3_ADD_467_U6, P3_REIP_REG_1__SCAN_IN, P3_REIP_REG_2__SCAN_IN);
  nand ginst20854 (P3_ADD_467_U60, P3_REIP_REG_29__SCAN_IN, P3_ADD_467_U120);
  not ginst20855 (P3_ADD_467_U61, P3_REIP_REG_30__SCAN_IN);
  nand ginst20856 (P3_ADD_467_U62, P3_ADD_467_U123, P3_ADD_467_U124);
  nand ginst20857 (P3_ADD_467_U63, P3_ADD_467_U125, P3_ADD_467_U126);
  nand ginst20858 (P3_ADD_467_U64, P3_ADD_467_U127, P3_ADD_467_U128);
  nand ginst20859 (P3_ADD_467_U65, P3_ADD_467_U129, P3_ADD_467_U130);
  nand ginst20860 (P3_ADD_467_U66, P3_ADD_467_U131, P3_ADD_467_U132);
  nand ginst20861 (P3_ADD_467_U67, P3_ADD_467_U133, P3_ADD_467_U134);
  nand ginst20862 (P3_ADD_467_U68, P3_ADD_467_U135, P3_ADD_467_U136);
  nand ginst20863 (P3_ADD_467_U69, P3_ADD_467_U137, P3_ADD_467_U138);
  not ginst20864 (P3_ADD_467_U7, P3_REIP_REG_3__SCAN_IN);
  nand ginst20865 (P3_ADD_467_U70, P3_ADD_467_U139, P3_ADD_467_U140);
  nand ginst20866 (P3_ADD_467_U71, P3_ADD_467_U141, P3_ADD_467_U142);
  nand ginst20867 (P3_ADD_467_U72, P3_ADD_467_U143, P3_ADD_467_U144);
  nand ginst20868 (P3_ADD_467_U73, P3_ADD_467_U145, P3_ADD_467_U146);
  nand ginst20869 (P3_ADD_467_U74, P3_ADD_467_U147, P3_ADD_467_U148);
  nand ginst20870 (P3_ADD_467_U75, P3_ADD_467_U149, P3_ADD_467_U150);
  nand ginst20871 (P3_ADD_467_U76, P3_ADD_467_U151, P3_ADD_467_U152);
  nand ginst20872 (P3_ADD_467_U77, P3_ADD_467_U153, P3_ADD_467_U154);
  nand ginst20873 (P3_ADD_467_U78, P3_ADD_467_U155, P3_ADD_467_U156);
  nand ginst20874 (P3_ADD_467_U79, P3_ADD_467_U157, P3_ADD_467_U158);
  nand ginst20875 (P3_ADD_467_U8, P3_REIP_REG_3__SCAN_IN, P3_ADD_467_U94);
  nand ginst20876 (P3_ADD_467_U80, P3_ADD_467_U159, P3_ADD_467_U160);
  nand ginst20877 (P3_ADD_467_U81, P3_ADD_467_U161, P3_ADD_467_U162);
  nand ginst20878 (P3_ADD_467_U82, P3_ADD_467_U163, P3_ADD_467_U164);
  nand ginst20879 (P3_ADD_467_U83, P3_ADD_467_U165, P3_ADD_467_U166);
  nand ginst20880 (P3_ADD_467_U84, P3_ADD_467_U167, P3_ADD_467_U168);
  nand ginst20881 (P3_ADD_467_U85, P3_ADD_467_U169, P3_ADD_467_U170);
  nand ginst20882 (P3_ADD_467_U86, P3_ADD_467_U171, P3_ADD_467_U172);
  nand ginst20883 (P3_ADD_467_U87, P3_ADD_467_U173, P3_ADD_467_U174);
  nand ginst20884 (P3_ADD_467_U88, P3_ADD_467_U175, P3_ADD_467_U176);
  nand ginst20885 (P3_ADD_467_U89, P3_ADD_467_U177, P3_ADD_467_U178);
  not ginst20886 (P3_ADD_467_U9, P3_REIP_REG_4__SCAN_IN);
  nand ginst20887 (P3_ADD_467_U90, P3_ADD_467_U179, P3_ADD_467_U180);
  nand ginst20888 (P3_ADD_467_U91, P3_ADD_467_U181, P3_ADD_467_U182);
  not ginst20889 (P3_ADD_467_U92, P3_REIP_REG_31__SCAN_IN);
  nand ginst20890 (P3_ADD_467_U93, P3_REIP_REG_30__SCAN_IN, P3_ADD_467_U121);
  not ginst20891 (P3_ADD_467_U94, P3_ADD_467_U6);
  not ginst20892 (P3_ADD_467_U95, P3_ADD_467_U8);
  not ginst20893 (P3_ADD_467_U96, P3_ADD_467_U10);
  not ginst20894 (P3_ADD_467_U97, P3_ADD_467_U12);
  not ginst20895 (P3_ADD_467_U98, P3_ADD_467_U14);
  not ginst20896 (P3_ADD_467_U99, P3_ADD_467_U16);
  nand ginst20897 (P3_ADD_476_U10, P3_INSTADDRPOINTER_REG_4__SCAN_IN, P3_ADD_476_U95);
  not ginst20898 (P3_ADD_476_U100, P3_ADD_476_U19);
  not ginst20899 (P3_ADD_476_U101, P3_ADD_476_U20);
  not ginst20900 (P3_ADD_476_U102, P3_ADD_476_U22);
  not ginst20901 (P3_ADD_476_U103, P3_ADD_476_U24);
  not ginst20902 (P3_ADD_476_U104, P3_ADD_476_U26);
  not ginst20903 (P3_ADD_476_U105, P3_ADD_476_U28);
  not ginst20904 (P3_ADD_476_U106, P3_ADD_476_U30);
  not ginst20905 (P3_ADD_476_U107, P3_ADD_476_U32);
  not ginst20906 (P3_ADD_476_U108, P3_ADD_476_U34);
  not ginst20907 (P3_ADD_476_U109, P3_ADD_476_U36);
  not ginst20908 (P3_ADD_476_U11, P3_INSTADDRPOINTER_REG_5__SCAN_IN);
  not ginst20909 (P3_ADD_476_U110, P3_ADD_476_U38);
  not ginst20910 (P3_ADD_476_U111, P3_ADD_476_U40);
  not ginst20911 (P3_ADD_476_U112, P3_ADD_476_U42);
  not ginst20912 (P3_ADD_476_U113, P3_ADD_476_U44);
  not ginst20913 (P3_ADD_476_U114, P3_ADD_476_U46);
  not ginst20914 (P3_ADD_476_U115, P3_ADD_476_U48);
  not ginst20915 (P3_ADD_476_U116, P3_ADD_476_U50);
  not ginst20916 (P3_ADD_476_U117, P3_ADD_476_U52);
  not ginst20917 (P3_ADD_476_U118, P3_ADD_476_U54);
  not ginst20918 (P3_ADD_476_U119, P3_ADD_476_U56);
  nand ginst20919 (P3_ADD_476_U12, P3_INSTADDRPOINTER_REG_5__SCAN_IN, P3_ADD_476_U96);
  not ginst20920 (P3_ADD_476_U120, P3_ADD_476_U58);
  not ginst20921 (P3_ADD_476_U121, P3_ADD_476_U60);
  not ginst20922 (P3_ADD_476_U122, P3_ADD_476_U93);
  nand ginst20923 (P3_ADD_476_U123, P3_INSTADDRPOINTER_REG_9__SCAN_IN, P3_ADD_476_U19);
  nand ginst20924 (P3_ADD_476_U124, P3_ADD_476_U100, P3_ADD_476_U18);
  nand ginst20925 (P3_ADD_476_U125, P3_INSTADDRPOINTER_REG_8__SCAN_IN, P3_ADD_476_U16);
  nand ginst20926 (P3_ADD_476_U126, P3_ADD_476_U17, P3_ADD_476_U99);
  nand ginst20927 (P3_ADD_476_U127, P3_INSTADDRPOINTER_REG_7__SCAN_IN, P3_ADD_476_U14);
  nand ginst20928 (P3_ADD_476_U128, P3_ADD_476_U15, P3_ADD_476_U98);
  nand ginst20929 (P3_ADD_476_U129, P3_INSTADDRPOINTER_REG_6__SCAN_IN, P3_ADD_476_U12);
  not ginst20930 (P3_ADD_476_U13, P3_INSTADDRPOINTER_REG_6__SCAN_IN);
  nand ginst20931 (P3_ADD_476_U130, P3_ADD_476_U13, P3_ADD_476_U97);
  nand ginst20932 (P3_ADD_476_U131, P3_INSTADDRPOINTER_REG_5__SCAN_IN, P3_ADD_476_U10);
  nand ginst20933 (P3_ADD_476_U132, P3_ADD_476_U11, P3_ADD_476_U96);
  nand ginst20934 (P3_ADD_476_U133, P3_INSTADDRPOINTER_REG_4__SCAN_IN, P3_ADD_476_U8);
  nand ginst20935 (P3_ADD_476_U134, P3_ADD_476_U9, P3_ADD_476_U95);
  nand ginst20936 (P3_ADD_476_U135, P3_INSTADDRPOINTER_REG_3__SCAN_IN, P3_ADD_476_U6);
  nand ginst20937 (P3_ADD_476_U136, P3_ADD_476_U7, P3_ADD_476_U94);
  nand ginst20938 (P3_ADD_476_U137, P3_INSTADDRPOINTER_REG_31__SCAN_IN, P3_ADD_476_U93);
  nand ginst20939 (P3_ADD_476_U138, P3_ADD_476_U122, P3_ADD_476_U92);
  nand ginst20940 (P3_ADD_476_U139, P3_INSTADDRPOINTER_REG_30__SCAN_IN, P3_ADD_476_U60);
  nand ginst20941 (P3_ADD_476_U14, P3_INSTADDRPOINTER_REG_6__SCAN_IN, P3_ADD_476_U97);
  nand ginst20942 (P3_ADD_476_U140, P3_ADD_476_U121, P3_ADD_476_U61);
  nand ginst20943 (P3_ADD_476_U141, P3_INSTADDRPOINTER_REG_2__SCAN_IN, P3_ADD_476_U4);
  nand ginst20944 (P3_ADD_476_U142, P3_INSTADDRPOINTER_REG_1__SCAN_IN, P3_ADD_476_U5);
  nand ginst20945 (P3_ADD_476_U143, P3_INSTADDRPOINTER_REG_29__SCAN_IN, P3_ADD_476_U58);
  nand ginst20946 (P3_ADD_476_U144, P3_ADD_476_U120, P3_ADD_476_U59);
  nand ginst20947 (P3_ADD_476_U145, P3_INSTADDRPOINTER_REG_28__SCAN_IN, P3_ADD_476_U56);
  nand ginst20948 (P3_ADD_476_U146, P3_ADD_476_U119, P3_ADD_476_U57);
  nand ginst20949 (P3_ADD_476_U147, P3_INSTADDRPOINTER_REG_27__SCAN_IN, P3_ADD_476_U54);
  nand ginst20950 (P3_ADD_476_U148, P3_ADD_476_U118, P3_ADD_476_U55);
  nand ginst20951 (P3_ADD_476_U149, P3_INSTADDRPOINTER_REG_26__SCAN_IN, P3_ADD_476_U52);
  not ginst20952 (P3_ADD_476_U15, P3_INSTADDRPOINTER_REG_7__SCAN_IN);
  nand ginst20953 (P3_ADD_476_U150, P3_ADD_476_U117, P3_ADD_476_U53);
  nand ginst20954 (P3_ADD_476_U151, P3_INSTADDRPOINTER_REG_25__SCAN_IN, P3_ADD_476_U50);
  nand ginst20955 (P3_ADD_476_U152, P3_ADD_476_U116, P3_ADD_476_U51);
  nand ginst20956 (P3_ADD_476_U153, P3_INSTADDRPOINTER_REG_24__SCAN_IN, P3_ADD_476_U48);
  nand ginst20957 (P3_ADD_476_U154, P3_ADD_476_U115, P3_ADD_476_U49);
  nand ginst20958 (P3_ADD_476_U155, P3_INSTADDRPOINTER_REG_23__SCAN_IN, P3_ADD_476_U46);
  nand ginst20959 (P3_ADD_476_U156, P3_ADD_476_U114, P3_ADD_476_U47);
  nand ginst20960 (P3_ADD_476_U157, P3_INSTADDRPOINTER_REG_22__SCAN_IN, P3_ADD_476_U44);
  nand ginst20961 (P3_ADD_476_U158, P3_ADD_476_U113, P3_ADD_476_U45);
  nand ginst20962 (P3_ADD_476_U159, P3_INSTADDRPOINTER_REG_21__SCAN_IN, P3_ADD_476_U42);
  nand ginst20963 (P3_ADD_476_U16, P3_INSTADDRPOINTER_REG_7__SCAN_IN, P3_ADD_476_U98);
  nand ginst20964 (P3_ADD_476_U160, P3_ADD_476_U112, P3_ADD_476_U43);
  nand ginst20965 (P3_ADD_476_U161, P3_INSTADDRPOINTER_REG_20__SCAN_IN, P3_ADD_476_U40);
  nand ginst20966 (P3_ADD_476_U162, P3_ADD_476_U111, P3_ADD_476_U41);
  nand ginst20967 (P3_ADD_476_U163, P3_INSTADDRPOINTER_REG_19__SCAN_IN, P3_ADD_476_U38);
  nand ginst20968 (P3_ADD_476_U164, P3_ADD_476_U110, P3_ADD_476_U39);
  nand ginst20969 (P3_ADD_476_U165, P3_INSTADDRPOINTER_REG_18__SCAN_IN, P3_ADD_476_U36);
  nand ginst20970 (P3_ADD_476_U166, P3_ADD_476_U109, P3_ADD_476_U37);
  nand ginst20971 (P3_ADD_476_U167, P3_INSTADDRPOINTER_REG_17__SCAN_IN, P3_ADD_476_U34);
  nand ginst20972 (P3_ADD_476_U168, P3_ADD_476_U108, P3_ADD_476_U35);
  nand ginst20973 (P3_ADD_476_U169, P3_INSTADDRPOINTER_REG_16__SCAN_IN, P3_ADD_476_U32);
  not ginst20974 (P3_ADD_476_U17, P3_INSTADDRPOINTER_REG_8__SCAN_IN);
  nand ginst20975 (P3_ADD_476_U170, P3_ADD_476_U107, P3_ADD_476_U33);
  nand ginst20976 (P3_ADD_476_U171, P3_INSTADDRPOINTER_REG_15__SCAN_IN, P3_ADD_476_U30);
  nand ginst20977 (P3_ADD_476_U172, P3_ADD_476_U106, P3_ADD_476_U31);
  nand ginst20978 (P3_ADD_476_U173, P3_INSTADDRPOINTER_REG_14__SCAN_IN, P3_ADD_476_U28);
  nand ginst20979 (P3_ADD_476_U174, P3_ADD_476_U105, P3_ADD_476_U29);
  nand ginst20980 (P3_ADD_476_U175, P3_INSTADDRPOINTER_REG_13__SCAN_IN, P3_ADD_476_U26);
  nand ginst20981 (P3_ADD_476_U176, P3_ADD_476_U104, P3_ADD_476_U27);
  nand ginst20982 (P3_ADD_476_U177, P3_INSTADDRPOINTER_REG_12__SCAN_IN, P3_ADD_476_U24);
  nand ginst20983 (P3_ADD_476_U178, P3_ADD_476_U103, P3_ADD_476_U25);
  nand ginst20984 (P3_ADD_476_U179, P3_INSTADDRPOINTER_REG_11__SCAN_IN, P3_ADD_476_U22);
  not ginst20985 (P3_ADD_476_U18, P3_INSTADDRPOINTER_REG_9__SCAN_IN);
  nand ginst20986 (P3_ADD_476_U180, P3_ADD_476_U102, P3_ADD_476_U23);
  nand ginst20987 (P3_ADD_476_U181, P3_INSTADDRPOINTER_REG_10__SCAN_IN, P3_ADD_476_U20);
  nand ginst20988 (P3_ADD_476_U182, P3_ADD_476_U101, P3_ADD_476_U21);
  nand ginst20989 (P3_ADD_476_U19, P3_INSTADDRPOINTER_REG_8__SCAN_IN, P3_ADD_476_U99);
  nand ginst20990 (P3_ADD_476_U20, P3_INSTADDRPOINTER_REG_9__SCAN_IN, P3_ADD_476_U100);
  not ginst20991 (P3_ADD_476_U21, P3_INSTADDRPOINTER_REG_10__SCAN_IN);
  nand ginst20992 (P3_ADD_476_U22, P3_INSTADDRPOINTER_REG_10__SCAN_IN, P3_ADD_476_U101);
  not ginst20993 (P3_ADD_476_U23, P3_INSTADDRPOINTER_REG_11__SCAN_IN);
  nand ginst20994 (P3_ADD_476_U24, P3_INSTADDRPOINTER_REG_11__SCAN_IN, P3_ADD_476_U102);
  not ginst20995 (P3_ADD_476_U25, P3_INSTADDRPOINTER_REG_12__SCAN_IN);
  nand ginst20996 (P3_ADD_476_U26, P3_INSTADDRPOINTER_REG_12__SCAN_IN, P3_ADD_476_U103);
  not ginst20997 (P3_ADD_476_U27, P3_INSTADDRPOINTER_REG_13__SCAN_IN);
  nand ginst20998 (P3_ADD_476_U28, P3_INSTADDRPOINTER_REG_13__SCAN_IN, P3_ADD_476_U104);
  not ginst20999 (P3_ADD_476_U29, P3_INSTADDRPOINTER_REG_14__SCAN_IN);
  nand ginst21000 (P3_ADD_476_U30, P3_INSTADDRPOINTER_REG_14__SCAN_IN, P3_ADD_476_U105);
  not ginst21001 (P3_ADD_476_U31, P3_INSTADDRPOINTER_REG_15__SCAN_IN);
  nand ginst21002 (P3_ADD_476_U32, P3_INSTADDRPOINTER_REG_15__SCAN_IN, P3_ADD_476_U106);
  not ginst21003 (P3_ADD_476_U33, P3_INSTADDRPOINTER_REG_16__SCAN_IN);
  nand ginst21004 (P3_ADD_476_U34, P3_INSTADDRPOINTER_REG_16__SCAN_IN, P3_ADD_476_U107);
  not ginst21005 (P3_ADD_476_U35, P3_INSTADDRPOINTER_REG_17__SCAN_IN);
  nand ginst21006 (P3_ADD_476_U36, P3_INSTADDRPOINTER_REG_17__SCAN_IN, P3_ADD_476_U108);
  not ginst21007 (P3_ADD_476_U37, P3_INSTADDRPOINTER_REG_18__SCAN_IN);
  nand ginst21008 (P3_ADD_476_U38, P3_INSTADDRPOINTER_REG_18__SCAN_IN, P3_ADD_476_U109);
  not ginst21009 (P3_ADD_476_U39, P3_INSTADDRPOINTER_REG_19__SCAN_IN);
  not ginst21010 (P3_ADD_476_U4, P3_INSTADDRPOINTER_REG_1__SCAN_IN);
  nand ginst21011 (P3_ADD_476_U40, P3_INSTADDRPOINTER_REG_19__SCAN_IN, P3_ADD_476_U110);
  not ginst21012 (P3_ADD_476_U41, P3_INSTADDRPOINTER_REG_20__SCAN_IN);
  nand ginst21013 (P3_ADD_476_U42, P3_INSTADDRPOINTER_REG_20__SCAN_IN, P3_ADD_476_U111);
  not ginst21014 (P3_ADD_476_U43, P3_INSTADDRPOINTER_REG_21__SCAN_IN);
  nand ginst21015 (P3_ADD_476_U44, P3_INSTADDRPOINTER_REG_21__SCAN_IN, P3_ADD_476_U112);
  not ginst21016 (P3_ADD_476_U45, P3_INSTADDRPOINTER_REG_22__SCAN_IN);
  nand ginst21017 (P3_ADD_476_U46, P3_INSTADDRPOINTER_REG_22__SCAN_IN, P3_ADD_476_U113);
  not ginst21018 (P3_ADD_476_U47, P3_INSTADDRPOINTER_REG_23__SCAN_IN);
  nand ginst21019 (P3_ADD_476_U48, P3_INSTADDRPOINTER_REG_23__SCAN_IN, P3_ADD_476_U114);
  not ginst21020 (P3_ADD_476_U49, P3_INSTADDRPOINTER_REG_24__SCAN_IN);
  not ginst21021 (P3_ADD_476_U5, P3_INSTADDRPOINTER_REG_2__SCAN_IN);
  nand ginst21022 (P3_ADD_476_U50, P3_INSTADDRPOINTER_REG_24__SCAN_IN, P3_ADD_476_U115);
  not ginst21023 (P3_ADD_476_U51, P3_INSTADDRPOINTER_REG_25__SCAN_IN);
  nand ginst21024 (P3_ADD_476_U52, P3_INSTADDRPOINTER_REG_25__SCAN_IN, P3_ADD_476_U116);
  not ginst21025 (P3_ADD_476_U53, P3_INSTADDRPOINTER_REG_26__SCAN_IN);
  nand ginst21026 (P3_ADD_476_U54, P3_INSTADDRPOINTER_REG_26__SCAN_IN, P3_ADD_476_U117);
  not ginst21027 (P3_ADD_476_U55, P3_INSTADDRPOINTER_REG_27__SCAN_IN);
  nand ginst21028 (P3_ADD_476_U56, P3_INSTADDRPOINTER_REG_27__SCAN_IN, P3_ADD_476_U118);
  not ginst21029 (P3_ADD_476_U57, P3_INSTADDRPOINTER_REG_28__SCAN_IN);
  nand ginst21030 (P3_ADD_476_U58, P3_INSTADDRPOINTER_REG_28__SCAN_IN, P3_ADD_476_U119);
  not ginst21031 (P3_ADD_476_U59, P3_INSTADDRPOINTER_REG_29__SCAN_IN);
  nand ginst21032 (P3_ADD_476_U6, P3_INSTADDRPOINTER_REG_1__SCAN_IN, P3_INSTADDRPOINTER_REG_2__SCAN_IN);
  nand ginst21033 (P3_ADD_476_U60, P3_INSTADDRPOINTER_REG_29__SCAN_IN, P3_ADD_476_U120);
  not ginst21034 (P3_ADD_476_U61, P3_INSTADDRPOINTER_REG_30__SCAN_IN);
  nand ginst21035 (P3_ADD_476_U62, P3_ADD_476_U123, P3_ADD_476_U124);
  nand ginst21036 (P3_ADD_476_U63, P3_ADD_476_U125, P3_ADD_476_U126);
  nand ginst21037 (P3_ADD_476_U64, P3_ADD_476_U127, P3_ADD_476_U128);
  nand ginst21038 (P3_ADD_476_U65, P3_ADD_476_U129, P3_ADD_476_U130);
  nand ginst21039 (P3_ADD_476_U66, P3_ADD_476_U131, P3_ADD_476_U132);
  nand ginst21040 (P3_ADD_476_U67, P3_ADD_476_U133, P3_ADD_476_U134);
  nand ginst21041 (P3_ADD_476_U68, P3_ADD_476_U135, P3_ADD_476_U136);
  nand ginst21042 (P3_ADD_476_U69, P3_ADD_476_U137, P3_ADD_476_U138);
  not ginst21043 (P3_ADD_476_U7, P3_INSTADDRPOINTER_REG_3__SCAN_IN);
  nand ginst21044 (P3_ADD_476_U70, P3_ADD_476_U139, P3_ADD_476_U140);
  nand ginst21045 (P3_ADD_476_U71, P3_ADD_476_U141, P3_ADD_476_U142);
  nand ginst21046 (P3_ADD_476_U72, P3_ADD_476_U143, P3_ADD_476_U144);
  nand ginst21047 (P3_ADD_476_U73, P3_ADD_476_U145, P3_ADD_476_U146);
  nand ginst21048 (P3_ADD_476_U74, P3_ADD_476_U147, P3_ADD_476_U148);
  nand ginst21049 (P3_ADD_476_U75, P3_ADD_476_U149, P3_ADD_476_U150);
  nand ginst21050 (P3_ADD_476_U76, P3_ADD_476_U151, P3_ADD_476_U152);
  nand ginst21051 (P3_ADD_476_U77, P3_ADD_476_U153, P3_ADD_476_U154);
  nand ginst21052 (P3_ADD_476_U78, P3_ADD_476_U155, P3_ADD_476_U156);
  nand ginst21053 (P3_ADD_476_U79, P3_ADD_476_U157, P3_ADD_476_U158);
  nand ginst21054 (P3_ADD_476_U8, P3_INSTADDRPOINTER_REG_3__SCAN_IN, P3_ADD_476_U94);
  nand ginst21055 (P3_ADD_476_U80, P3_ADD_476_U159, P3_ADD_476_U160);
  nand ginst21056 (P3_ADD_476_U81, P3_ADD_476_U161, P3_ADD_476_U162);
  nand ginst21057 (P3_ADD_476_U82, P3_ADD_476_U163, P3_ADD_476_U164);
  nand ginst21058 (P3_ADD_476_U83, P3_ADD_476_U165, P3_ADD_476_U166);
  nand ginst21059 (P3_ADD_476_U84, P3_ADD_476_U167, P3_ADD_476_U168);
  nand ginst21060 (P3_ADD_476_U85, P3_ADD_476_U169, P3_ADD_476_U170);
  nand ginst21061 (P3_ADD_476_U86, P3_ADD_476_U171, P3_ADD_476_U172);
  nand ginst21062 (P3_ADD_476_U87, P3_ADD_476_U173, P3_ADD_476_U174);
  nand ginst21063 (P3_ADD_476_U88, P3_ADD_476_U175, P3_ADD_476_U176);
  nand ginst21064 (P3_ADD_476_U89, P3_ADD_476_U177, P3_ADD_476_U178);
  not ginst21065 (P3_ADD_476_U9, P3_INSTADDRPOINTER_REG_4__SCAN_IN);
  nand ginst21066 (P3_ADD_476_U90, P3_ADD_476_U179, P3_ADD_476_U180);
  nand ginst21067 (P3_ADD_476_U91, P3_ADD_476_U181, P3_ADD_476_U182);
  not ginst21068 (P3_ADD_476_U92, P3_INSTADDRPOINTER_REG_31__SCAN_IN);
  nand ginst21069 (P3_ADD_476_U93, P3_INSTADDRPOINTER_REG_30__SCAN_IN, P3_ADD_476_U121);
  not ginst21070 (P3_ADD_476_U94, P3_ADD_476_U6);
  not ginst21071 (P3_ADD_476_U95, P3_ADD_476_U8);
  not ginst21072 (P3_ADD_476_U96, P3_ADD_476_U10);
  not ginst21073 (P3_ADD_476_U97, P3_ADD_476_U12);
  not ginst21074 (P3_ADD_476_U98, P3_ADD_476_U14);
  not ginst21075 (P3_ADD_476_U99, P3_ADD_476_U16);
  nand ginst21076 (P3_ADD_486_U10, P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN, P3_ADD_486_U18);
  not ginst21077 (P3_ADD_486_U11, P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN);
  nand ginst21078 (P3_ADD_486_U12, P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P3_ADD_486_U19);
  not ginst21079 (P3_ADD_486_U13, P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN);
  nand ginst21080 (P3_ADD_486_U14, P3_ADD_486_U21, P3_ADD_486_U22);
  nand ginst21081 (P3_ADD_486_U15, P3_ADD_486_U23, P3_ADD_486_U24);
  nand ginst21082 (P3_ADD_486_U16, P3_ADD_486_U25, P3_ADD_486_U26);
  nand ginst21083 (P3_ADD_486_U17, P3_ADD_486_U27, P3_ADD_486_U28);
  not ginst21084 (P3_ADD_486_U18, P3_ADD_486_U8);
  not ginst21085 (P3_ADD_486_U19, P3_ADD_486_U10);
  not ginst21086 (P3_ADD_486_U20, P3_ADD_486_U12);
  nand ginst21087 (P3_ADD_486_U21, P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN, P3_ADD_486_U12);
  nand ginst21088 (P3_ADD_486_U22, P3_ADD_486_U13, P3_ADD_486_U20);
  nand ginst21089 (P3_ADD_486_U23, P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P3_ADD_486_U10);
  nand ginst21090 (P3_ADD_486_U24, P3_ADD_486_U11, P3_ADD_486_U19);
  nand ginst21091 (P3_ADD_486_U25, P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN, P3_ADD_486_U8);
  nand ginst21092 (P3_ADD_486_U26, P3_ADD_486_U18, P3_ADD_486_U9);
  nand ginst21093 (P3_ADD_486_U27, P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P3_ADD_486_U5);
  nand ginst21094 (P3_ADD_486_U28, P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN, P3_ADD_486_U7);
  not ginst21095 (P3_ADD_486_U5, P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN);
  and ginst21096 (P3_ADD_486_U6, P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN, P3_ADD_486_U20);
  not ginst21097 (P3_ADD_486_U7, P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN);
  nand ginst21098 (P3_ADD_486_U8, P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN);
  not ginst21099 (P3_ADD_486_U9, P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN);
  nand ginst21100 (P3_ADD_494_U10, P3_INSTADDRPOINTER_REG_4__SCAN_IN, P3_ADD_494_U95);
  not ginst21101 (P3_ADD_494_U100, P3_ADD_494_U19);
  not ginst21102 (P3_ADD_494_U101, P3_ADD_494_U20);
  not ginst21103 (P3_ADD_494_U102, P3_ADD_494_U22);
  not ginst21104 (P3_ADD_494_U103, P3_ADD_494_U24);
  not ginst21105 (P3_ADD_494_U104, P3_ADD_494_U26);
  not ginst21106 (P3_ADD_494_U105, P3_ADD_494_U28);
  not ginst21107 (P3_ADD_494_U106, P3_ADD_494_U30);
  not ginst21108 (P3_ADD_494_U107, P3_ADD_494_U32);
  not ginst21109 (P3_ADD_494_U108, P3_ADD_494_U34);
  not ginst21110 (P3_ADD_494_U109, P3_ADD_494_U36);
  not ginst21111 (P3_ADD_494_U11, P3_INSTADDRPOINTER_REG_5__SCAN_IN);
  not ginst21112 (P3_ADD_494_U110, P3_ADD_494_U38);
  not ginst21113 (P3_ADD_494_U111, P3_ADD_494_U40);
  not ginst21114 (P3_ADD_494_U112, P3_ADD_494_U42);
  not ginst21115 (P3_ADD_494_U113, P3_ADD_494_U44);
  not ginst21116 (P3_ADD_494_U114, P3_ADD_494_U46);
  not ginst21117 (P3_ADD_494_U115, P3_ADD_494_U48);
  not ginst21118 (P3_ADD_494_U116, P3_ADD_494_U50);
  not ginst21119 (P3_ADD_494_U117, P3_ADD_494_U52);
  not ginst21120 (P3_ADD_494_U118, P3_ADD_494_U54);
  not ginst21121 (P3_ADD_494_U119, P3_ADD_494_U56);
  nand ginst21122 (P3_ADD_494_U12, P3_INSTADDRPOINTER_REG_5__SCAN_IN, P3_ADD_494_U96);
  not ginst21123 (P3_ADD_494_U120, P3_ADD_494_U58);
  not ginst21124 (P3_ADD_494_U121, P3_ADD_494_U60);
  not ginst21125 (P3_ADD_494_U122, P3_ADD_494_U93);
  nand ginst21126 (P3_ADD_494_U123, P3_INSTADDRPOINTER_REG_9__SCAN_IN, P3_ADD_494_U19);
  nand ginst21127 (P3_ADD_494_U124, P3_ADD_494_U100, P3_ADD_494_U18);
  nand ginst21128 (P3_ADD_494_U125, P3_INSTADDRPOINTER_REG_8__SCAN_IN, P3_ADD_494_U16);
  nand ginst21129 (P3_ADD_494_U126, P3_ADD_494_U17, P3_ADD_494_U99);
  nand ginst21130 (P3_ADD_494_U127, P3_INSTADDRPOINTER_REG_7__SCAN_IN, P3_ADD_494_U14);
  nand ginst21131 (P3_ADD_494_U128, P3_ADD_494_U15, P3_ADD_494_U98);
  nand ginst21132 (P3_ADD_494_U129, P3_INSTADDRPOINTER_REG_6__SCAN_IN, P3_ADD_494_U12);
  not ginst21133 (P3_ADD_494_U13, P3_INSTADDRPOINTER_REG_6__SCAN_IN);
  nand ginst21134 (P3_ADD_494_U130, P3_ADD_494_U13, P3_ADD_494_U97);
  nand ginst21135 (P3_ADD_494_U131, P3_INSTADDRPOINTER_REG_5__SCAN_IN, P3_ADD_494_U10);
  nand ginst21136 (P3_ADD_494_U132, P3_ADD_494_U11, P3_ADD_494_U96);
  nand ginst21137 (P3_ADD_494_U133, P3_INSTADDRPOINTER_REG_4__SCAN_IN, P3_ADD_494_U8);
  nand ginst21138 (P3_ADD_494_U134, P3_ADD_494_U9, P3_ADD_494_U95);
  nand ginst21139 (P3_ADD_494_U135, P3_INSTADDRPOINTER_REG_3__SCAN_IN, P3_ADD_494_U6);
  nand ginst21140 (P3_ADD_494_U136, P3_ADD_494_U7, P3_ADD_494_U94);
  nand ginst21141 (P3_ADD_494_U137, P3_INSTADDRPOINTER_REG_31__SCAN_IN, P3_ADD_494_U93);
  nand ginst21142 (P3_ADD_494_U138, P3_ADD_494_U122, P3_ADD_494_U92);
  nand ginst21143 (P3_ADD_494_U139, P3_INSTADDRPOINTER_REG_30__SCAN_IN, P3_ADD_494_U60);
  nand ginst21144 (P3_ADD_494_U14, P3_INSTADDRPOINTER_REG_6__SCAN_IN, P3_ADD_494_U97);
  nand ginst21145 (P3_ADD_494_U140, P3_ADD_494_U121, P3_ADD_494_U61);
  nand ginst21146 (P3_ADD_494_U141, P3_INSTADDRPOINTER_REG_2__SCAN_IN, P3_ADD_494_U4);
  nand ginst21147 (P3_ADD_494_U142, P3_INSTADDRPOINTER_REG_1__SCAN_IN, P3_ADD_494_U5);
  nand ginst21148 (P3_ADD_494_U143, P3_INSTADDRPOINTER_REG_29__SCAN_IN, P3_ADD_494_U58);
  nand ginst21149 (P3_ADD_494_U144, P3_ADD_494_U120, P3_ADD_494_U59);
  nand ginst21150 (P3_ADD_494_U145, P3_INSTADDRPOINTER_REG_28__SCAN_IN, P3_ADD_494_U56);
  nand ginst21151 (P3_ADD_494_U146, P3_ADD_494_U119, P3_ADD_494_U57);
  nand ginst21152 (P3_ADD_494_U147, P3_INSTADDRPOINTER_REG_27__SCAN_IN, P3_ADD_494_U54);
  nand ginst21153 (P3_ADD_494_U148, P3_ADD_494_U118, P3_ADD_494_U55);
  nand ginst21154 (P3_ADD_494_U149, P3_INSTADDRPOINTER_REG_26__SCAN_IN, P3_ADD_494_U52);
  not ginst21155 (P3_ADD_494_U15, P3_INSTADDRPOINTER_REG_7__SCAN_IN);
  nand ginst21156 (P3_ADD_494_U150, P3_ADD_494_U117, P3_ADD_494_U53);
  nand ginst21157 (P3_ADD_494_U151, P3_INSTADDRPOINTER_REG_25__SCAN_IN, P3_ADD_494_U50);
  nand ginst21158 (P3_ADD_494_U152, P3_ADD_494_U116, P3_ADD_494_U51);
  nand ginst21159 (P3_ADD_494_U153, P3_INSTADDRPOINTER_REG_24__SCAN_IN, P3_ADD_494_U48);
  nand ginst21160 (P3_ADD_494_U154, P3_ADD_494_U115, P3_ADD_494_U49);
  nand ginst21161 (P3_ADD_494_U155, P3_INSTADDRPOINTER_REG_23__SCAN_IN, P3_ADD_494_U46);
  nand ginst21162 (P3_ADD_494_U156, P3_ADD_494_U114, P3_ADD_494_U47);
  nand ginst21163 (P3_ADD_494_U157, P3_INSTADDRPOINTER_REG_22__SCAN_IN, P3_ADD_494_U44);
  nand ginst21164 (P3_ADD_494_U158, P3_ADD_494_U113, P3_ADD_494_U45);
  nand ginst21165 (P3_ADD_494_U159, P3_INSTADDRPOINTER_REG_21__SCAN_IN, P3_ADD_494_U42);
  nand ginst21166 (P3_ADD_494_U16, P3_INSTADDRPOINTER_REG_7__SCAN_IN, P3_ADD_494_U98);
  nand ginst21167 (P3_ADD_494_U160, P3_ADD_494_U112, P3_ADD_494_U43);
  nand ginst21168 (P3_ADD_494_U161, P3_INSTADDRPOINTER_REG_20__SCAN_IN, P3_ADD_494_U40);
  nand ginst21169 (P3_ADD_494_U162, P3_ADD_494_U111, P3_ADD_494_U41);
  nand ginst21170 (P3_ADD_494_U163, P3_INSTADDRPOINTER_REG_19__SCAN_IN, P3_ADD_494_U38);
  nand ginst21171 (P3_ADD_494_U164, P3_ADD_494_U110, P3_ADD_494_U39);
  nand ginst21172 (P3_ADD_494_U165, P3_INSTADDRPOINTER_REG_18__SCAN_IN, P3_ADD_494_U36);
  nand ginst21173 (P3_ADD_494_U166, P3_ADD_494_U109, P3_ADD_494_U37);
  nand ginst21174 (P3_ADD_494_U167, P3_INSTADDRPOINTER_REG_17__SCAN_IN, P3_ADD_494_U34);
  nand ginst21175 (P3_ADD_494_U168, P3_ADD_494_U108, P3_ADD_494_U35);
  nand ginst21176 (P3_ADD_494_U169, P3_INSTADDRPOINTER_REG_16__SCAN_IN, P3_ADD_494_U32);
  not ginst21177 (P3_ADD_494_U17, P3_INSTADDRPOINTER_REG_8__SCAN_IN);
  nand ginst21178 (P3_ADD_494_U170, P3_ADD_494_U107, P3_ADD_494_U33);
  nand ginst21179 (P3_ADD_494_U171, P3_INSTADDRPOINTER_REG_15__SCAN_IN, P3_ADD_494_U30);
  nand ginst21180 (P3_ADD_494_U172, P3_ADD_494_U106, P3_ADD_494_U31);
  nand ginst21181 (P3_ADD_494_U173, P3_INSTADDRPOINTER_REG_14__SCAN_IN, P3_ADD_494_U28);
  nand ginst21182 (P3_ADD_494_U174, P3_ADD_494_U105, P3_ADD_494_U29);
  nand ginst21183 (P3_ADD_494_U175, P3_INSTADDRPOINTER_REG_13__SCAN_IN, P3_ADD_494_U26);
  nand ginst21184 (P3_ADD_494_U176, P3_ADD_494_U104, P3_ADD_494_U27);
  nand ginst21185 (P3_ADD_494_U177, P3_INSTADDRPOINTER_REG_12__SCAN_IN, P3_ADD_494_U24);
  nand ginst21186 (P3_ADD_494_U178, P3_ADD_494_U103, P3_ADD_494_U25);
  nand ginst21187 (P3_ADD_494_U179, P3_INSTADDRPOINTER_REG_11__SCAN_IN, P3_ADD_494_U22);
  not ginst21188 (P3_ADD_494_U18, P3_INSTADDRPOINTER_REG_9__SCAN_IN);
  nand ginst21189 (P3_ADD_494_U180, P3_ADD_494_U102, P3_ADD_494_U23);
  nand ginst21190 (P3_ADD_494_U181, P3_INSTADDRPOINTER_REG_10__SCAN_IN, P3_ADD_494_U20);
  nand ginst21191 (P3_ADD_494_U182, P3_ADD_494_U101, P3_ADD_494_U21);
  nand ginst21192 (P3_ADD_494_U19, P3_INSTADDRPOINTER_REG_8__SCAN_IN, P3_ADD_494_U99);
  nand ginst21193 (P3_ADD_494_U20, P3_INSTADDRPOINTER_REG_9__SCAN_IN, P3_ADD_494_U100);
  not ginst21194 (P3_ADD_494_U21, P3_INSTADDRPOINTER_REG_10__SCAN_IN);
  nand ginst21195 (P3_ADD_494_U22, P3_INSTADDRPOINTER_REG_10__SCAN_IN, P3_ADD_494_U101);
  not ginst21196 (P3_ADD_494_U23, P3_INSTADDRPOINTER_REG_11__SCAN_IN);
  nand ginst21197 (P3_ADD_494_U24, P3_INSTADDRPOINTER_REG_11__SCAN_IN, P3_ADD_494_U102);
  not ginst21198 (P3_ADD_494_U25, P3_INSTADDRPOINTER_REG_12__SCAN_IN);
  nand ginst21199 (P3_ADD_494_U26, P3_INSTADDRPOINTER_REG_12__SCAN_IN, P3_ADD_494_U103);
  not ginst21200 (P3_ADD_494_U27, P3_INSTADDRPOINTER_REG_13__SCAN_IN);
  nand ginst21201 (P3_ADD_494_U28, P3_INSTADDRPOINTER_REG_13__SCAN_IN, P3_ADD_494_U104);
  not ginst21202 (P3_ADD_494_U29, P3_INSTADDRPOINTER_REG_14__SCAN_IN);
  nand ginst21203 (P3_ADD_494_U30, P3_INSTADDRPOINTER_REG_14__SCAN_IN, P3_ADD_494_U105);
  not ginst21204 (P3_ADD_494_U31, P3_INSTADDRPOINTER_REG_15__SCAN_IN);
  nand ginst21205 (P3_ADD_494_U32, P3_INSTADDRPOINTER_REG_15__SCAN_IN, P3_ADD_494_U106);
  not ginst21206 (P3_ADD_494_U33, P3_INSTADDRPOINTER_REG_16__SCAN_IN);
  nand ginst21207 (P3_ADD_494_U34, P3_INSTADDRPOINTER_REG_16__SCAN_IN, P3_ADD_494_U107);
  not ginst21208 (P3_ADD_494_U35, P3_INSTADDRPOINTER_REG_17__SCAN_IN);
  nand ginst21209 (P3_ADD_494_U36, P3_INSTADDRPOINTER_REG_17__SCAN_IN, P3_ADD_494_U108);
  not ginst21210 (P3_ADD_494_U37, P3_INSTADDRPOINTER_REG_18__SCAN_IN);
  nand ginst21211 (P3_ADD_494_U38, P3_INSTADDRPOINTER_REG_18__SCAN_IN, P3_ADD_494_U109);
  not ginst21212 (P3_ADD_494_U39, P3_INSTADDRPOINTER_REG_19__SCAN_IN);
  not ginst21213 (P3_ADD_494_U4, P3_INSTADDRPOINTER_REG_1__SCAN_IN);
  nand ginst21214 (P3_ADD_494_U40, P3_INSTADDRPOINTER_REG_19__SCAN_IN, P3_ADD_494_U110);
  not ginst21215 (P3_ADD_494_U41, P3_INSTADDRPOINTER_REG_20__SCAN_IN);
  nand ginst21216 (P3_ADD_494_U42, P3_INSTADDRPOINTER_REG_20__SCAN_IN, P3_ADD_494_U111);
  not ginst21217 (P3_ADD_494_U43, P3_INSTADDRPOINTER_REG_21__SCAN_IN);
  nand ginst21218 (P3_ADD_494_U44, P3_INSTADDRPOINTER_REG_21__SCAN_IN, P3_ADD_494_U112);
  not ginst21219 (P3_ADD_494_U45, P3_INSTADDRPOINTER_REG_22__SCAN_IN);
  nand ginst21220 (P3_ADD_494_U46, P3_INSTADDRPOINTER_REG_22__SCAN_IN, P3_ADD_494_U113);
  not ginst21221 (P3_ADD_494_U47, P3_INSTADDRPOINTER_REG_23__SCAN_IN);
  nand ginst21222 (P3_ADD_494_U48, P3_INSTADDRPOINTER_REG_23__SCAN_IN, P3_ADD_494_U114);
  not ginst21223 (P3_ADD_494_U49, P3_INSTADDRPOINTER_REG_24__SCAN_IN);
  not ginst21224 (P3_ADD_494_U5, P3_INSTADDRPOINTER_REG_2__SCAN_IN);
  nand ginst21225 (P3_ADD_494_U50, P3_INSTADDRPOINTER_REG_24__SCAN_IN, P3_ADD_494_U115);
  not ginst21226 (P3_ADD_494_U51, P3_INSTADDRPOINTER_REG_25__SCAN_IN);
  nand ginst21227 (P3_ADD_494_U52, P3_INSTADDRPOINTER_REG_25__SCAN_IN, P3_ADD_494_U116);
  not ginst21228 (P3_ADD_494_U53, P3_INSTADDRPOINTER_REG_26__SCAN_IN);
  nand ginst21229 (P3_ADD_494_U54, P3_INSTADDRPOINTER_REG_26__SCAN_IN, P3_ADD_494_U117);
  not ginst21230 (P3_ADD_494_U55, P3_INSTADDRPOINTER_REG_27__SCAN_IN);
  nand ginst21231 (P3_ADD_494_U56, P3_INSTADDRPOINTER_REG_27__SCAN_IN, P3_ADD_494_U118);
  not ginst21232 (P3_ADD_494_U57, P3_INSTADDRPOINTER_REG_28__SCAN_IN);
  nand ginst21233 (P3_ADD_494_U58, P3_INSTADDRPOINTER_REG_28__SCAN_IN, P3_ADD_494_U119);
  not ginst21234 (P3_ADD_494_U59, P3_INSTADDRPOINTER_REG_29__SCAN_IN);
  nand ginst21235 (P3_ADD_494_U6, P3_INSTADDRPOINTER_REG_1__SCAN_IN, P3_INSTADDRPOINTER_REG_2__SCAN_IN);
  nand ginst21236 (P3_ADD_494_U60, P3_INSTADDRPOINTER_REG_29__SCAN_IN, P3_ADD_494_U120);
  not ginst21237 (P3_ADD_494_U61, P3_INSTADDRPOINTER_REG_30__SCAN_IN);
  nand ginst21238 (P3_ADD_494_U62, P3_ADD_494_U123, P3_ADD_494_U124);
  nand ginst21239 (P3_ADD_494_U63, P3_ADD_494_U125, P3_ADD_494_U126);
  nand ginst21240 (P3_ADD_494_U64, P3_ADD_494_U127, P3_ADD_494_U128);
  nand ginst21241 (P3_ADD_494_U65, P3_ADD_494_U129, P3_ADD_494_U130);
  nand ginst21242 (P3_ADD_494_U66, P3_ADD_494_U131, P3_ADD_494_U132);
  nand ginst21243 (P3_ADD_494_U67, P3_ADD_494_U133, P3_ADD_494_U134);
  nand ginst21244 (P3_ADD_494_U68, P3_ADD_494_U135, P3_ADD_494_U136);
  nand ginst21245 (P3_ADD_494_U69, P3_ADD_494_U137, P3_ADD_494_U138);
  not ginst21246 (P3_ADD_494_U7, P3_INSTADDRPOINTER_REG_3__SCAN_IN);
  nand ginst21247 (P3_ADD_494_U70, P3_ADD_494_U139, P3_ADD_494_U140);
  nand ginst21248 (P3_ADD_494_U71, P3_ADD_494_U141, P3_ADD_494_U142);
  nand ginst21249 (P3_ADD_494_U72, P3_ADD_494_U143, P3_ADD_494_U144);
  nand ginst21250 (P3_ADD_494_U73, P3_ADD_494_U145, P3_ADD_494_U146);
  nand ginst21251 (P3_ADD_494_U74, P3_ADD_494_U147, P3_ADD_494_U148);
  nand ginst21252 (P3_ADD_494_U75, P3_ADD_494_U149, P3_ADD_494_U150);
  nand ginst21253 (P3_ADD_494_U76, P3_ADD_494_U151, P3_ADD_494_U152);
  nand ginst21254 (P3_ADD_494_U77, P3_ADD_494_U153, P3_ADD_494_U154);
  nand ginst21255 (P3_ADD_494_U78, P3_ADD_494_U155, P3_ADD_494_U156);
  nand ginst21256 (P3_ADD_494_U79, P3_ADD_494_U157, P3_ADD_494_U158);
  nand ginst21257 (P3_ADD_494_U8, P3_INSTADDRPOINTER_REG_3__SCAN_IN, P3_ADD_494_U94);
  nand ginst21258 (P3_ADD_494_U80, P3_ADD_494_U159, P3_ADD_494_U160);
  nand ginst21259 (P3_ADD_494_U81, P3_ADD_494_U161, P3_ADD_494_U162);
  nand ginst21260 (P3_ADD_494_U82, P3_ADD_494_U163, P3_ADD_494_U164);
  nand ginst21261 (P3_ADD_494_U83, P3_ADD_494_U165, P3_ADD_494_U166);
  nand ginst21262 (P3_ADD_494_U84, P3_ADD_494_U167, P3_ADD_494_U168);
  nand ginst21263 (P3_ADD_494_U85, P3_ADD_494_U169, P3_ADD_494_U170);
  nand ginst21264 (P3_ADD_494_U86, P3_ADD_494_U171, P3_ADD_494_U172);
  nand ginst21265 (P3_ADD_494_U87, P3_ADD_494_U173, P3_ADD_494_U174);
  nand ginst21266 (P3_ADD_494_U88, P3_ADD_494_U175, P3_ADD_494_U176);
  nand ginst21267 (P3_ADD_494_U89, P3_ADD_494_U177, P3_ADD_494_U178);
  not ginst21268 (P3_ADD_494_U9, P3_INSTADDRPOINTER_REG_4__SCAN_IN);
  nand ginst21269 (P3_ADD_494_U90, P3_ADD_494_U179, P3_ADD_494_U180);
  nand ginst21270 (P3_ADD_494_U91, P3_ADD_494_U181, P3_ADD_494_U182);
  not ginst21271 (P3_ADD_494_U92, P3_INSTADDRPOINTER_REG_31__SCAN_IN);
  nand ginst21272 (P3_ADD_494_U93, P3_INSTADDRPOINTER_REG_30__SCAN_IN, P3_ADD_494_U121);
  not ginst21273 (P3_ADD_494_U94, P3_ADD_494_U6);
  not ginst21274 (P3_ADD_494_U95, P3_ADD_494_U8);
  not ginst21275 (P3_ADD_494_U96, P3_ADD_494_U10);
  not ginst21276 (P3_ADD_494_U97, P3_ADD_494_U12);
  not ginst21277 (P3_ADD_494_U98, P3_ADD_494_U14);
  not ginst21278 (P3_ADD_494_U99, P3_ADD_494_U16);
  nand ginst21279 (P3_ADD_495_U10, P3_ADD_495_U19, P3_ADD_495_U20);
  not ginst21280 (P3_ADD_495_U11, P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN);
  nand ginst21281 (P3_ADD_495_U12, P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P3_ADD_495_U13);
  not ginst21282 (P3_ADD_495_U13, P3_ADD_495_U6);
  not ginst21283 (P3_ADD_495_U14, P3_ADD_495_U12);
  nand ginst21284 (P3_ADD_495_U15, P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN, P3_ADD_495_U12);
  nand ginst21285 (P3_ADD_495_U16, P3_ADD_495_U11, P3_ADD_495_U14);
  nand ginst21286 (P3_ADD_495_U17, P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P3_ADD_495_U6);
  nand ginst21287 (P3_ADD_495_U18, P3_ADD_495_U13, P3_ADD_495_U7);
  nand ginst21288 (P3_ADD_495_U19, P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN, P3_ADD_495_U4);
  nand ginst21289 (P3_ADD_495_U20, P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P3_ADD_495_U5);
  not ginst21290 (P3_ADD_495_U4, P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN);
  not ginst21291 (P3_ADD_495_U5, P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN);
  nand ginst21292 (P3_ADD_495_U6, P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN, P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN);
  not ginst21293 (P3_ADD_495_U7, P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN);
  nand ginst21294 (P3_ADD_495_U8, P3_ADD_495_U15, P3_ADD_495_U16);
  nand ginst21295 (P3_ADD_495_U9, P3_ADD_495_U17, P3_ADD_495_U18);
  nand ginst21296 (P3_ADD_505_U10, P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN, P3_ADD_505_U18);
  not ginst21297 (P3_ADD_505_U11, P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN);
  nand ginst21298 (P3_ADD_505_U12, P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P3_ADD_505_U19);
  not ginst21299 (P3_ADD_505_U13, P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN);
  nand ginst21300 (P3_ADD_505_U14, P3_ADD_505_U21, P3_ADD_505_U22);
  nand ginst21301 (P3_ADD_505_U15, P3_ADD_505_U23, P3_ADD_505_U24);
  nand ginst21302 (P3_ADD_505_U16, P3_ADD_505_U25, P3_ADD_505_U26);
  nand ginst21303 (P3_ADD_505_U17, P3_ADD_505_U27, P3_ADD_505_U28);
  not ginst21304 (P3_ADD_505_U18, P3_ADD_505_U8);
  not ginst21305 (P3_ADD_505_U19, P3_ADD_505_U10);
  not ginst21306 (P3_ADD_505_U20, P3_ADD_505_U12);
  nand ginst21307 (P3_ADD_505_U21, P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN, P3_ADD_505_U12);
  nand ginst21308 (P3_ADD_505_U22, P3_ADD_505_U13, P3_ADD_505_U20);
  nand ginst21309 (P3_ADD_505_U23, P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P3_ADD_505_U10);
  nand ginst21310 (P3_ADD_505_U24, P3_ADD_505_U11, P3_ADD_505_U19);
  nand ginst21311 (P3_ADD_505_U25, P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN, P3_ADD_505_U8);
  nand ginst21312 (P3_ADD_505_U26, P3_ADD_505_U18, P3_ADD_505_U9);
  nand ginst21313 (P3_ADD_505_U27, P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P3_ADD_505_U5);
  nand ginst21314 (P3_ADD_505_U28, P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN, P3_ADD_505_U7);
  not ginst21315 (P3_ADD_505_U5, P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN);
  and ginst21316 (P3_ADD_505_U6, P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN, P3_ADD_505_U20);
  not ginst21317 (P3_ADD_505_U7, P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN);
  nand ginst21318 (P3_ADD_505_U8, P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN);
  not ginst21319 (P3_ADD_505_U9, P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN);
  nand ginst21320 (P3_ADD_515_U10, P3_INSTADDRPOINTER_REG_4__SCAN_IN, P3_ADD_515_U95);
  not ginst21321 (P3_ADD_515_U100, P3_ADD_515_U19);
  not ginst21322 (P3_ADD_515_U101, P3_ADD_515_U20);
  not ginst21323 (P3_ADD_515_U102, P3_ADD_515_U22);
  not ginst21324 (P3_ADD_515_U103, P3_ADD_515_U24);
  not ginst21325 (P3_ADD_515_U104, P3_ADD_515_U26);
  not ginst21326 (P3_ADD_515_U105, P3_ADD_515_U28);
  not ginst21327 (P3_ADD_515_U106, P3_ADD_515_U30);
  not ginst21328 (P3_ADD_515_U107, P3_ADD_515_U32);
  not ginst21329 (P3_ADD_515_U108, P3_ADD_515_U34);
  not ginst21330 (P3_ADD_515_U109, P3_ADD_515_U36);
  not ginst21331 (P3_ADD_515_U11, P3_INSTADDRPOINTER_REG_5__SCAN_IN);
  not ginst21332 (P3_ADD_515_U110, P3_ADD_515_U38);
  not ginst21333 (P3_ADD_515_U111, P3_ADD_515_U40);
  not ginst21334 (P3_ADD_515_U112, P3_ADD_515_U42);
  not ginst21335 (P3_ADD_515_U113, P3_ADD_515_U44);
  not ginst21336 (P3_ADD_515_U114, P3_ADD_515_U46);
  not ginst21337 (P3_ADD_515_U115, P3_ADD_515_U48);
  not ginst21338 (P3_ADD_515_U116, P3_ADD_515_U50);
  not ginst21339 (P3_ADD_515_U117, P3_ADD_515_U52);
  not ginst21340 (P3_ADD_515_U118, P3_ADD_515_U54);
  not ginst21341 (P3_ADD_515_U119, P3_ADD_515_U56);
  nand ginst21342 (P3_ADD_515_U12, P3_INSTADDRPOINTER_REG_5__SCAN_IN, P3_ADD_515_U96);
  not ginst21343 (P3_ADD_515_U120, P3_ADD_515_U58);
  not ginst21344 (P3_ADD_515_U121, P3_ADD_515_U60);
  not ginst21345 (P3_ADD_515_U122, P3_ADD_515_U93);
  nand ginst21346 (P3_ADD_515_U123, P3_INSTADDRPOINTER_REG_9__SCAN_IN, P3_ADD_515_U19);
  nand ginst21347 (P3_ADD_515_U124, P3_ADD_515_U100, P3_ADD_515_U18);
  nand ginst21348 (P3_ADD_515_U125, P3_INSTADDRPOINTER_REG_8__SCAN_IN, P3_ADD_515_U16);
  nand ginst21349 (P3_ADD_515_U126, P3_ADD_515_U17, P3_ADD_515_U99);
  nand ginst21350 (P3_ADD_515_U127, P3_INSTADDRPOINTER_REG_7__SCAN_IN, P3_ADD_515_U14);
  nand ginst21351 (P3_ADD_515_U128, P3_ADD_515_U15, P3_ADD_515_U98);
  nand ginst21352 (P3_ADD_515_U129, P3_INSTADDRPOINTER_REG_6__SCAN_IN, P3_ADD_515_U12);
  not ginst21353 (P3_ADD_515_U13, P3_INSTADDRPOINTER_REG_6__SCAN_IN);
  nand ginst21354 (P3_ADD_515_U130, P3_ADD_515_U13, P3_ADD_515_U97);
  nand ginst21355 (P3_ADD_515_U131, P3_INSTADDRPOINTER_REG_5__SCAN_IN, P3_ADD_515_U10);
  nand ginst21356 (P3_ADD_515_U132, P3_ADD_515_U11, P3_ADD_515_U96);
  nand ginst21357 (P3_ADD_515_U133, P3_INSTADDRPOINTER_REG_4__SCAN_IN, P3_ADD_515_U8);
  nand ginst21358 (P3_ADD_515_U134, P3_ADD_515_U9, P3_ADD_515_U95);
  nand ginst21359 (P3_ADD_515_U135, P3_INSTADDRPOINTER_REG_3__SCAN_IN, P3_ADD_515_U6);
  nand ginst21360 (P3_ADD_515_U136, P3_ADD_515_U7, P3_ADD_515_U94);
  nand ginst21361 (P3_ADD_515_U137, P3_INSTADDRPOINTER_REG_31__SCAN_IN, P3_ADD_515_U93);
  nand ginst21362 (P3_ADD_515_U138, P3_ADD_515_U122, P3_ADD_515_U92);
  nand ginst21363 (P3_ADD_515_U139, P3_INSTADDRPOINTER_REG_30__SCAN_IN, P3_ADD_515_U60);
  nand ginst21364 (P3_ADD_515_U14, P3_INSTADDRPOINTER_REG_6__SCAN_IN, P3_ADD_515_U97);
  nand ginst21365 (P3_ADD_515_U140, P3_ADD_515_U121, P3_ADD_515_U61);
  nand ginst21366 (P3_ADD_515_U141, P3_INSTADDRPOINTER_REG_2__SCAN_IN, P3_ADD_515_U4);
  nand ginst21367 (P3_ADD_515_U142, P3_INSTADDRPOINTER_REG_1__SCAN_IN, P3_ADD_515_U5);
  nand ginst21368 (P3_ADD_515_U143, P3_INSTADDRPOINTER_REG_29__SCAN_IN, P3_ADD_515_U58);
  nand ginst21369 (P3_ADD_515_U144, P3_ADD_515_U120, P3_ADD_515_U59);
  nand ginst21370 (P3_ADD_515_U145, P3_INSTADDRPOINTER_REG_28__SCAN_IN, P3_ADD_515_U56);
  nand ginst21371 (P3_ADD_515_U146, P3_ADD_515_U119, P3_ADD_515_U57);
  nand ginst21372 (P3_ADD_515_U147, P3_INSTADDRPOINTER_REG_27__SCAN_IN, P3_ADD_515_U54);
  nand ginst21373 (P3_ADD_515_U148, P3_ADD_515_U118, P3_ADD_515_U55);
  nand ginst21374 (P3_ADD_515_U149, P3_INSTADDRPOINTER_REG_26__SCAN_IN, P3_ADD_515_U52);
  not ginst21375 (P3_ADD_515_U15, P3_INSTADDRPOINTER_REG_7__SCAN_IN);
  nand ginst21376 (P3_ADD_515_U150, P3_ADD_515_U117, P3_ADD_515_U53);
  nand ginst21377 (P3_ADD_515_U151, P3_INSTADDRPOINTER_REG_25__SCAN_IN, P3_ADD_515_U50);
  nand ginst21378 (P3_ADD_515_U152, P3_ADD_515_U116, P3_ADD_515_U51);
  nand ginst21379 (P3_ADD_515_U153, P3_INSTADDRPOINTER_REG_24__SCAN_IN, P3_ADD_515_U48);
  nand ginst21380 (P3_ADD_515_U154, P3_ADD_515_U115, P3_ADD_515_U49);
  nand ginst21381 (P3_ADD_515_U155, P3_INSTADDRPOINTER_REG_23__SCAN_IN, P3_ADD_515_U46);
  nand ginst21382 (P3_ADD_515_U156, P3_ADD_515_U114, P3_ADD_515_U47);
  nand ginst21383 (P3_ADD_515_U157, P3_INSTADDRPOINTER_REG_22__SCAN_IN, P3_ADD_515_U44);
  nand ginst21384 (P3_ADD_515_U158, P3_ADD_515_U113, P3_ADD_515_U45);
  nand ginst21385 (P3_ADD_515_U159, P3_INSTADDRPOINTER_REG_21__SCAN_IN, P3_ADD_515_U42);
  nand ginst21386 (P3_ADD_515_U16, P3_INSTADDRPOINTER_REG_7__SCAN_IN, P3_ADD_515_U98);
  nand ginst21387 (P3_ADD_515_U160, P3_ADD_515_U112, P3_ADD_515_U43);
  nand ginst21388 (P3_ADD_515_U161, P3_INSTADDRPOINTER_REG_20__SCAN_IN, P3_ADD_515_U40);
  nand ginst21389 (P3_ADD_515_U162, P3_ADD_515_U111, P3_ADD_515_U41);
  nand ginst21390 (P3_ADD_515_U163, P3_INSTADDRPOINTER_REG_19__SCAN_IN, P3_ADD_515_U38);
  nand ginst21391 (P3_ADD_515_U164, P3_ADD_515_U110, P3_ADD_515_U39);
  nand ginst21392 (P3_ADD_515_U165, P3_INSTADDRPOINTER_REG_18__SCAN_IN, P3_ADD_515_U36);
  nand ginst21393 (P3_ADD_515_U166, P3_ADD_515_U109, P3_ADD_515_U37);
  nand ginst21394 (P3_ADD_515_U167, P3_INSTADDRPOINTER_REG_17__SCAN_IN, P3_ADD_515_U34);
  nand ginst21395 (P3_ADD_515_U168, P3_ADD_515_U108, P3_ADD_515_U35);
  nand ginst21396 (P3_ADD_515_U169, P3_INSTADDRPOINTER_REG_16__SCAN_IN, P3_ADD_515_U32);
  not ginst21397 (P3_ADD_515_U17, P3_INSTADDRPOINTER_REG_8__SCAN_IN);
  nand ginst21398 (P3_ADD_515_U170, P3_ADD_515_U107, P3_ADD_515_U33);
  nand ginst21399 (P3_ADD_515_U171, P3_INSTADDRPOINTER_REG_15__SCAN_IN, P3_ADD_515_U30);
  nand ginst21400 (P3_ADD_515_U172, P3_ADD_515_U106, P3_ADD_515_U31);
  nand ginst21401 (P3_ADD_515_U173, P3_INSTADDRPOINTER_REG_14__SCAN_IN, P3_ADD_515_U28);
  nand ginst21402 (P3_ADD_515_U174, P3_ADD_515_U105, P3_ADD_515_U29);
  nand ginst21403 (P3_ADD_515_U175, P3_INSTADDRPOINTER_REG_13__SCAN_IN, P3_ADD_515_U26);
  nand ginst21404 (P3_ADD_515_U176, P3_ADD_515_U104, P3_ADD_515_U27);
  nand ginst21405 (P3_ADD_515_U177, P3_INSTADDRPOINTER_REG_12__SCAN_IN, P3_ADD_515_U24);
  nand ginst21406 (P3_ADD_515_U178, P3_ADD_515_U103, P3_ADD_515_U25);
  nand ginst21407 (P3_ADD_515_U179, P3_INSTADDRPOINTER_REG_11__SCAN_IN, P3_ADD_515_U22);
  not ginst21408 (P3_ADD_515_U18, P3_INSTADDRPOINTER_REG_9__SCAN_IN);
  nand ginst21409 (P3_ADD_515_U180, P3_ADD_515_U102, P3_ADD_515_U23);
  nand ginst21410 (P3_ADD_515_U181, P3_INSTADDRPOINTER_REG_10__SCAN_IN, P3_ADD_515_U20);
  nand ginst21411 (P3_ADD_515_U182, P3_ADD_515_U101, P3_ADD_515_U21);
  nand ginst21412 (P3_ADD_515_U19, P3_INSTADDRPOINTER_REG_8__SCAN_IN, P3_ADD_515_U99);
  nand ginst21413 (P3_ADD_515_U20, P3_INSTADDRPOINTER_REG_9__SCAN_IN, P3_ADD_515_U100);
  not ginst21414 (P3_ADD_515_U21, P3_INSTADDRPOINTER_REG_10__SCAN_IN);
  nand ginst21415 (P3_ADD_515_U22, P3_INSTADDRPOINTER_REG_10__SCAN_IN, P3_ADD_515_U101);
  not ginst21416 (P3_ADD_515_U23, P3_INSTADDRPOINTER_REG_11__SCAN_IN);
  nand ginst21417 (P3_ADD_515_U24, P3_INSTADDRPOINTER_REG_11__SCAN_IN, P3_ADD_515_U102);
  not ginst21418 (P3_ADD_515_U25, P3_INSTADDRPOINTER_REG_12__SCAN_IN);
  nand ginst21419 (P3_ADD_515_U26, P3_INSTADDRPOINTER_REG_12__SCAN_IN, P3_ADD_515_U103);
  not ginst21420 (P3_ADD_515_U27, P3_INSTADDRPOINTER_REG_13__SCAN_IN);
  nand ginst21421 (P3_ADD_515_U28, P3_INSTADDRPOINTER_REG_13__SCAN_IN, P3_ADD_515_U104);
  not ginst21422 (P3_ADD_515_U29, P3_INSTADDRPOINTER_REG_14__SCAN_IN);
  nand ginst21423 (P3_ADD_515_U30, P3_INSTADDRPOINTER_REG_14__SCAN_IN, P3_ADD_515_U105);
  not ginst21424 (P3_ADD_515_U31, P3_INSTADDRPOINTER_REG_15__SCAN_IN);
  nand ginst21425 (P3_ADD_515_U32, P3_INSTADDRPOINTER_REG_15__SCAN_IN, P3_ADD_515_U106);
  not ginst21426 (P3_ADD_515_U33, P3_INSTADDRPOINTER_REG_16__SCAN_IN);
  nand ginst21427 (P3_ADD_515_U34, P3_INSTADDRPOINTER_REG_16__SCAN_IN, P3_ADD_515_U107);
  not ginst21428 (P3_ADD_515_U35, P3_INSTADDRPOINTER_REG_17__SCAN_IN);
  nand ginst21429 (P3_ADD_515_U36, P3_INSTADDRPOINTER_REG_17__SCAN_IN, P3_ADD_515_U108);
  not ginst21430 (P3_ADD_515_U37, P3_INSTADDRPOINTER_REG_18__SCAN_IN);
  nand ginst21431 (P3_ADD_515_U38, P3_INSTADDRPOINTER_REG_18__SCAN_IN, P3_ADD_515_U109);
  not ginst21432 (P3_ADD_515_U39, P3_INSTADDRPOINTER_REG_19__SCAN_IN);
  not ginst21433 (P3_ADD_515_U4, P3_INSTADDRPOINTER_REG_1__SCAN_IN);
  nand ginst21434 (P3_ADD_515_U40, P3_INSTADDRPOINTER_REG_19__SCAN_IN, P3_ADD_515_U110);
  not ginst21435 (P3_ADD_515_U41, P3_INSTADDRPOINTER_REG_20__SCAN_IN);
  nand ginst21436 (P3_ADD_515_U42, P3_INSTADDRPOINTER_REG_20__SCAN_IN, P3_ADD_515_U111);
  not ginst21437 (P3_ADD_515_U43, P3_INSTADDRPOINTER_REG_21__SCAN_IN);
  nand ginst21438 (P3_ADD_515_U44, P3_INSTADDRPOINTER_REG_21__SCAN_IN, P3_ADD_515_U112);
  not ginst21439 (P3_ADD_515_U45, P3_INSTADDRPOINTER_REG_22__SCAN_IN);
  nand ginst21440 (P3_ADD_515_U46, P3_INSTADDRPOINTER_REG_22__SCAN_IN, P3_ADD_515_U113);
  not ginst21441 (P3_ADD_515_U47, P3_INSTADDRPOINTER_REG_23__SCAN_IN);
  nand ginst21442 (P3_ADD_515_U48, P3_INSTADDRPOINTER_REG_23__SCAN_IN, P3_ADD_515_U114);
  not ginst21443 (P3_ADD_515_U49, P3_INSTADDRPOINTER_REG_24__SCAN_IN);
  not ginst21444 (P3_ADD_515_U5, P3_INSTADDRPOINTER_REG_2__SCAN_IN);
  nand ginst21445 (P3_ADD_515_U50, P3_INSTADDRPOINTER_REG_24__SCAN_IN, P3_ADD_515_U115);
  not ginst21446 (P3_ADD_515_U51, P3_INSTADDRPOINTER_REG_25__SCAN_IN);
  nand ginst21447 (P3_ADD_515_U52, P3_INSTADDRPOINTER_REG_25__SCAN_IN, P3_ADD_515_U116);
  not ginst21448 (P3_ADD_515_U53, P3_INSTADDRPOINTER_REG_26__SCAN_IN);
  nand ginst21449 (P3_ADD_515_U54, P3_INSTADDRPOINTER_REG_26__SCAN_IN, P3_ADD_515_U117);
  not ginst21450 (P3_ADD_515_U55, P3_INSTADDRPOINTER_REG_27__SCAN_IN);
  nand ginst21451 (P3_ADD_515_U56, P3_INSTADDRPOINTER_REG_27__SCAN_IN, P3_ADD_515_U118);
  not ginst21452 (P3_ADD_515_U57, P3_INSTADDRPOINTER_REG_28__SCAN_IN);
  nand ginst21453 (P3_ADD_515_U58, P3_INSTADDRPOINTER_REG_28__SCAN_IN, P3_ADD_515_U119);
  not ginst21454 (P3_ADD_515_U59, P3_INSTADDRPOINTER_REG_29__SCAN_IN);
  nand ginst21455 (P3_ADD_515_U6, P3_INSTADDRPOINTER_REG_1__SCAN_IN, P3_INSTADDRPOINTER_REG_2__SCAN_IN);
  nand ginst21456 (P3_ADD_515_U60, P3_INSTADDRPOINTER_REG_29__SCAN_IN, P3_ADD_515_U120);
  not ginst21457 (P3_ADD_515_U61, P3_INSTADDRPOINTER_REG_30__SCAN_IN);
  nand ginst21458 (P3_ADD_515_U62, P3_ADD_515_U123, P3_ADD_515_U124);
  nand ginst21459 (P3_ADD_515_U63, P3_ADD_515_U125, P3_ADD_515_U126);
  nand ginst21460 (P3_ADD_515_U64, P3_ADD_515_U127, P3_ADD_515_U128);
  nand ginst21461 (P3_ADD_515_U65, P3_ADD_515_U129, P3_ADD_515_U130);
  nand ginst21462 (P3_ADD_515_U66, P3_ADD_515_U131, P3_ADD_515_U132);
  nand ginst21463 (P3_ADD_515_U67, P3_ADD_515_U133, P3_ADD_515_U134);
  nand ginst21464 (P3_ADD_515_U68, P3_ADD_515_U135, P3_ADD_515_U136);
  nand ginst21465 (P3_ADD_515_U69, P3_ADD_515_U137, P3_ADD_515_U138);
  not ginst21466 (P3_ADD_515_U7, P3_INSTADDRPOINTER_REG_3__SCAN_IN);
  nand ginst21467 (P3_ADD_515_U70, P3_ADD_515_U139, P3_ADD_515_U140);
  nand ginst21468 (P3_ADD_515_U71, P3_ADD_515_U141, P3_ADD_515_U142);
  nand ginst21469 (P3_ADD_515_U72, P3_ADD_515_U143, P3_ADD_515_U144);
  nand ginst21470 (P3_ADD_515_U73, P3_ADD_515_U145, P3_ADD_515_U146);
  nand ginst21471 (P3_ADD_515_U74, P3_ADD_515_U147, P3_ADD_515_U148);
  nand ginst21472 (P3_ADD_515_U75, P3_ADD_515_U149, P3_ADD_515_U150);
  nand ginst21473 (P3_ADD_515_U76, P3_ADD_515_U151, P3_ADD_515_U152);
  nand ginst21474 (P3_ADD_515_U77, P3_ADD_515_U153, P3_ADD_515_U154);
  nand ginst21475 (P3_ADD_515_U78, P3_ADD_515_U155, P3_ADD_515_U156);
  nand ginst21476 (P3_ADD_515_U79, P3_ADD_515_U157, P3_ADD_515_U158);
  nand ginst21477 (P3_ADD_515_U8, P3_INSTADDRPOINTER_REG_3__SCAN_IN, P3_ADD_515_U94);
  nand ginst21478 (P3_ADD_515_U80, P3_ADD_515_U159, P3_ADD_515_U160);
  nand ginst21479 (P3_ADD_515_U81, P3_ADD_515_U161, P3_ADD_515_U162);
  nand ginst21480 (P3_ADD_515_U82, P3_ADD_515_U163, P3_ADD_515_U164);
  nand ginst21481 (P3_ADD_515_U83, P3_ADD_515_U165, P3_ADD_515_U166);
  nand ginst21482 (P3_ADD_515_U84, P3_ADD_515_U167, P3_ADD_515_U168);
  nand ginst21483 (P3_ADD_515_U85, P3_ADD_515_U169, P3_ADD_515_U170);
  nand ginst21484 (P3_ADD_515_U86, P3_ADD_515_U171, P3_ADD_515_U172);
  nand ginst21485 (P3_ADD_515_U87, P3_ADD_515_U173, P3_ADD_515_U174);
  nand ginst21486 (P3_ADD_515_U88, P3_ADD_515_U175, P3_ADD_515_U176);
  nand ginst21487 (P3_ADD_515_U89, P3_ADD_515_U177, P3_ADD_515_U178);
  not ginst21488 (P3_ADD_515_U9, P3_INSTADDRPOINTER_REG_4__SCAN_IN);
  nand ginst21489 (P3_ADD_515_U90, P3_ADD_515_U179, P3_ADD_515_U180);
  nand ginst21490 (P3_ADD_515_U91, P3_ADD_515_U181, P3_ADD_515_U182);
  not ginst21491 (P3_ADD_515_U92, P3_INSTADDRPOINTER_REG_31__SCAN_IN);
  nand ginst21492 (P3_ADD_515_U93, P3_INSTADDRPOINTER_REG_30__SCAN_IN, P3_ADD_515_U121);
  not ginst21493 (P3_ADD_515_U94, P3_ADD_515_U6);
  not ginst21494 (P3_ADD_515_U95, P3_ADD_515_U8);
  not ginst21495 (P3_ADD_515_U96, P3_ADD_515_U10);
  not ginst21496 (P3_ADD_515_U97, P3_ADD_515_U12);
  not ginst21497 (P3_ADD_515_U98, P3_ADD_515_U14);
  not ginst21498 (P3_ADD_515_U99, P3_ADD_515_U16);
  nand ginst21499 (P3_ADD_526_U10, P3_INSTADDRPOINTER_REG_0__SCAN_IN, P3_INSTADDRPOINTER_REG_1__SCAN_IN, P3_INSTADDRPOINTER_REG_2__SCAN_IN);
  nand ginst21500 (P3_ADD_526_U100, P3_INSTADDRPOINTER_REG_0__SCAN_IN, P3_INSTADDRPOINTER_REG_1__SCAN_IN);
  nand ginst21501 (P3_ADD_526_U101, P3_INSTADDRPOINTER_REG_27__SCAN_IN, P3_ADD_526_U122);
  nand ginst21502 (P3_ADD_526_U102, P3_INSTADDRPOINTER_REG_25__SCAN_IN, P3_ADD_526_U116);
  nand ginst21503 (P3_ADD_526_U103, P3_INSTADDRPOINTER_REG_23__SCAN_IN, P3_ADD_526_U115);
  nand ginst21504 (P3_ADD_526_U104, P3_INSTADDRPOINTER_REG_21__SCAN_IN, P3_ADD_526_U121);
  nand ginst21505 (P3_ADD_526_U105, P3_INSTADDRPOINTER_REG_19__SCAN_IN, P3_ADD_526_U114);
  nand ginst21506 (P3_ADD_526_U106, P3_INSTADDRPOINTER_REG_17__SCAN_IN, P3_ADD_526_U117);
  nand ginst21507 (P3_ADD_526_U107, P3_INSTADDRPOINTER_REG_15__SCAN_IN, P3_ADD_526_U124);
  nand ginst21508 (P3_ADD_526_U108, P3_INSTADDRPOINTER_REG_13__SCAN_IN, P3_ADD_526_U119);
  nand ginst21509 (P3_ADD_526_U109, P3_INSTADDRPOINTER_REG_11__SCAN_IN, P3_ADD_526_U113);
  not ginst21510 (P3_ADD_526_U11, P3_INSTADDRPOINTER_REG_6__SCAN_IN);
  nand ginst21511 (P3_ADD_526_U110, P3_INSTADDRPOINTER_REG_9__SCAN_IN, P3_ADD_526_U120);
  not ginst21512 (P3_ADD_526_U111, P3_ADD_526_U10);
  not ginst21513 (P3_ADD_526_U112, P3_ADD_526_U13);
  not ginst21514 (P3_ADD_526_U113, P3_ADD_526_U22);
  not ginst21515 (P3_ADD_526_U114, P3_ADD_526_U34);
  not ginst21516 (P3_ADD_526_U115, P3_ADD_526_U40);
  not ginst21517 (P3_ADD_526_U116, P3_ADD_526_U43);
  not ginst21518 (P3_ADD_526_U117, P3_ADD_526_U31);
  not ginst21519 (P3_ADD_526_U118, P3_ADD_526_U16);
  not ginst21520 (P3_ADD_526_U119, P3_ADD_526_U25);
  not ginst21521 (P3_ADD_526_U12, P3_INSTADDRPOINTER_REG_5__SCAN_IN);
  not ginst21522 (P3_ADD_526_U120, P3_ADD_526_U17);
  not ginst21523 (P3_ADD_526_U121, P3_ADD_526_U36);
  not ginst21524 (P3_ADD_526_U122, P3_ADD_526_U46);
  not ginst21525 (P3_ADD_526_U123, P3_ADD_526_U48);
  not ginst21526 (P3_ADD_526_U124, P3_ADD_526_U27);
  not ginst21527 (P3_ADD_526_U125, P3_ADD_526_U95);
  not ginst21528 (P3_ADD_526_U126, P3_ADD_526_U96);
  not ginst21529 (P3_ADD_526_U127, P3_ADD_526_U97);
  not ginst21530 (P3_ADD_526_U128, P3_ADD_526_U49);
  not ginst21531 (P3_ADD_526_U129, P3_ADD_526_U99);
  nand ginst21532 (P3_ADD_526_U13, P3_ADD_526_U111, P3_ADD_526_U82);
  not ginst21533 (P3_ADD_526_U130, P3_ADD_526_U100);
  not ginst21534 (P3_ADD_526_U131, P3_ADD_526_U101);
  not ginst21535 (P3_ADD_526_U132, P3_ADD_526_U102);
  not ginst21536 (P3_ADD_526_U133, P3_ADD_526_U103);
  not ginst21537 (P3_ADD_526_U134, P3_ADD_526_U104);
  not ginst21538 (P3_ADD_526_U135, P3_ADD_526_U105);
  not ginst21539 (P3_ADD_526_U136, P3_ADD_526_U106);
  not ginst21540 (P3_ADD_526_U137, P3_ADD_526_U107);
  not ginst21541 (P3_ADD_526_U138, P3_ADD_526_U108);
  not ginst21542 (P3_ADD_526_U139, P3_ADD_526_U109);
  not ginst21543 (P3_ADD_526_U14, P3_INSTADDRPOINTER_REG_8__SCAN_IN);
  not ginst21544 (P3_ADD_526_U140, P3_ADD_526_U110);
  nand ginst21545 (P3_ADD_526_U141, P3_ADD_526_U120, P3_ADD_526_U18);
  nand ginst21546 (P3_ADD_526_U142, P3_INSTADDRPOINTER_REG_9__SCAN_IN, P3_ADD_526_U17);
  nand ginst21547 (P3_ADD_526_U143, P3_INSTADDRPOINTER_REG_8__SCAN_IN, P3_ADD_526_U95);
  nand ginst21548 (P3_ADD_526_U144, P3_ADD_526_U125, P3_ADD_526_U14);
  nand ginst21549 (P3_ADD_526_U145, P3_ADD_526_U118, P3_ADD_526_U15);
  nand ginst21550 (P3_ADD_526_U146, P3_INSTADDRPOINTER_REG_7__SCAN_IN, P3_ADD_526_U16);
  nand ginst21551 (P3_ADD_526_U147, P3_INSTADDRPOINTER_REG_6__SCAN_IN, P3_ADD_526_U96);
  nand ginst21552 (P3_ADD_526_U148, P3_ADD_526_U11, P3_ADD_526_U126);
  nand ginst21553 (P3_ADD_526_U149, P3_ADD_526_U112, P3_ADD_526_U12);
  not ginst21554 (P3_ADD_526_U15, P3_INSTADDRPOINTER_REG_7__SCAN_IN);
  nand ginst21555 (P3_ADD_526_U150, P3_INSTADDRPOINTER_REG_5__SCAN_IN, P3_ADD_526_U13);
  nand ginst21556 (P3_ADD_526_U151, P3_INSTADDRPOINTER_REG_4__SCAN_IN, P3_ADD_526_U97);
  nand ginst21557 (P3_ADD_526_U152, P3_ADD_526_U127, P3_ADD_526_U8);
  nand ginst21558 (P3_ADD_526_U153, P3_ADD_526_U111, P3_ADD_526_U9);
  nand ginst21559 (P3_ADD_526_U154, P3_INSTADDRPOINTER_REG_3__SCAN_IN, P3_ADD_526_U10);
  nand ginst21560 (P3_ADD_526_U155, P3_INSTADDRPOINTER_REG_31__SCAN_IN, P3_ADD_526_U99);
  nand ginst21561 (P3_ADD_526_U156, P3_ADD_526_U129, P3_ADD_526_U98);
  nand ginst21562 (P3_ADD_526_U157, P3_INSTADDRPOINTER_REG_30__SCAN_IN, P3_ADD_526_U49);
  nand ginst21563 (P3_ADD_526_U158, P3_ADD_526_U128, P3_ADD_526_U50);
  nand ginst21564 (P3_ADD_526_U159, P3_INSTADDRPOINTER_REG_2__SCAN_IN, P3_ADD_526_U100);
  nand ginst21565 (P3_ADD_526_U16, P3_ADD_526_U112, P3_ADD_526_U83);
  nand ginst21566 (P3_ADD_526_U160, P3_ADD_526_U130, P3_ADD_526_U6);
  nand ginst21567 (P3_ADD_526_U161, P3_ADD_526_U123, P3_ADD_526_U47);
  nand ginst21568 (P3_ADD_526_U162, P3_INSTADDRPOINTER_REG_29__SCAN_IN, P3_ADD_526_U48);
  nand ginst21569 (P3_ADD_526_U163, P3_INSTADDRPOINTER_REG_28__SCAN_IN, P3_ADD_526_U101);
  nand ginst21570 (P3_ADD_526_U164, P3_ADD_526_U131, P3_ADD_526_U45);
  nand ginst21571 (P3_ADD_526_U165, P3_ADD_526_U122, P3_ADD_526_U44);
  nand ginst21572 (P3_ADD_526_U166, P3_INSTADDRPOINTER_REG_27__SCAN_IN, P3_ADD_526_U46);
  nand ginst21573 (P3_ADD_526_U167, P3_INSTADDRPOINTER_REG_26__SCAN_IN, P3_ADD_526_U102);
  nand ginst21574 (P3_ADD_526_U168, P3_ADD_526_U132, P3_ADD_526_U41);
  nand ginst21575 (P3_ADD_526_U169, P3_ADD_526_U116, P3_ADD_526_U42);
  nand ginst21576 (P3_ADD_526_U17, P3_ADD_526_U118, P3_ADD_526_U84);
  nand ginst21577 (P3_ADD_526_U170, P3_INSTADDRPOINTER_REG_25__SCAN_IN, P3_ADD_526_U43);
  nand ginst21578 (P3_ADD_526_U171, P3_INSTADDRPOINTER_REG_24__SCAN_IN, P3_ADD_526_U103);
  nand ginst21579 (P3_ADD_526_U172, P3_ADD_526_U133, P3_ADD_526_U38);
  nand ginst21580 (P3_ADD_526_U173, P3_ADD_526_U115, P3_ADD_526_U39);
  nand ginst21581 (P3_ADD_526_U174, P3_INSTADDRPOINTER_REG_23__SCAN_IN, P3_ADD_526_U40);
  nand ginst21582 (P3_ADD_526_U175, P3_INSTADDRPOINTER_REG_22__SCAN_IN, P3_ADD_526_U104);
  nand ginst21583 (P3_ADD_526_U176, P3_ADD_526_U134, P3_ADD_526_U37);
  nand ginst21584 (P3_ADD_526_U177, P3_ADD_526_U121, P3_ADD_526_U35);
  nand ginst21585 (P3_ADD_526_U178, P3_INSTADDRPOINTER_REG_21__SCAN_IN, P3_ADD_526_U36);
  nand ginst21586 (P3_ADD_526_U179, P3_INSTADDRPOINTER_REG_20__SCAN_IN, P3_ADD_526_U105);
  not ginst21587 (P3_ADD_526_U18, P3_INSTADDRPOINTER_REG_9__SCAN_IN);
  nand ginst21588 (P3_ADD_526_U180, P3_ADD_526_U135, P3_ADD_526_U32);
  nand ginst21589 (P3_ADD_526_U181, P3_INSTADDRPOINTER_REG_0__SCAN_IN, P3_ADD_526_U7);
  nand ginst21590 (P3_ADD_526_U182, P3_INSTADDRPOINTER_REG_1__SCAN_IN, P3_ADD_526_U5);
  nand ginst21591 (P3_ADD_526_U183, P3_ADD_526_U114, P3_ADD_526_U33);
  nand ginst21592 (P3_ADD_526_U184, P3_INSTADDRPOINTER_REG_19__SCAN_IN, P3_ADD_526_U34);
  nand ginst21593 (P3_ADD_526_U185, P3_INSTADDRPOINTER_REG_18__SCAN_IN, P3_ADD_526_U106);
  nand ginst21594 (P3_ADD_526_U186, P3_ADD_526_U136, P3_ADD_526_U29);
  nand ginst21595 (P3_ADD_526_U187, P3_ADD_526_U117, P3_ADD_526_U30);
  nand ginst21596 (P3_ADD_526_U188, P3_INSTADDRPOINTER_REG_17__SCAN_IN, P3_ADD_526_U31);
  nand ginst21597 (P3_ADD_526_U189, P3_INSTADDRPOINTER_REG_16__SCAN_IN, P3_ADD_526_U107);
  not ginst21598 (P3_ADD_526_U19, P3_INSTADDRPOINTER_REG_10__SCAN_IN);
  nand ginst21599 (P3_ADD_526_U190, P3_ADD_526_U137, P3_ADD_526_U28);
  nand ginst21600 (P3_ADD_526_U191, P3_ADD_526_U124, P3_ADD_526_U26);
  nand ginst21601 (P3_ADD_526_U192, P3_INSTADDRPOINTER_REG_15__SCAN_IN, P3_ADD_526_U27);
  nand ginst21602 (P3_ADD_526_U193, P3_INSTADDRPOINTER_REG_14__SCAN_IN, P3_ADD_526_U108);
  nand ginst21603 (P3_ADD_526_U194, P3_ADD_526_U138, P3_ADD_526_U23);
  nand ginst21604 (P3_ADD_526_U195, P3_ADD_526_U119, P3_ADD_526_U24);
  nand ginst21605 (P3_ADD_526_U196, P3_INSTADDRPOINTER_REG_13__SCAN_IN, P3_ADD_526_U25);
  nand ginst21606 (P3_ADD_526_U197, P3_INSTADDRPOINTER_REG_12__SCAN_IN, P3_ADD_526_U109);
  nand ginst21607 (P3_ADD_526_U198, P3_ADD_526_U139, P3_ADD_526_U20);
  nand ginst21608 (P3_ADD_526_U199, P3_ADD_526_U113, P3_ADD_526_U21);
  not ginst21609 (P3_ADD_526_U20, P3_INSTADDRPOINTER_REG_12__SCAN_IN);
  nand ginst21610 (P3_ADD_526_U200, P3_INSTADDRPOINTER_REG_11__SCAN_IN, P3_ADD_526_U22);
  nand ginst21611 (P3_ADD_526_U201, P3_INSTADDRPOINTER_REG_10__SCAN_IN, P3_ADD_526_U110);
  nand ginst21612 (P3_ADD_526_U202, P3_ADD_526_U140, P3_ADD_526_U19);
  not ginst21613 (P3_ADD_526_U21, P3_INSTADDRPOINTER_REG_11__SCAN_IN);
  nand ginst21614 (P3_ADD_526_U22, P3_ADD_526_U120, P3_ADD_526_U85);
  not ginst21615 (P3_ADD_526_U23, P3_INSTADDRPOINTER_REG_14__SCAN_IN);
  not ginst21616 (P3_ADD_526_U24, P3_INSTADDRPOINTER_REG_13__SCAN_IN);
  nand ginst21617 (P3_ADD_526_U25, P3_ADD_526_U113, P3_ADD_526_U86);
  not ginst21618 (P3_ADD_526_U26, P3_INSTADDRPOINTER_REG_15__SCAN_IN);
  nand ginst21619 (P3_ADD_526_U27, P3_ADD_526_U119, P3_ADD_526_U87);
  not ginst21620 (P3_ADD_526_U28, P3_INSTADDRPOINTER_REG_16__SCAN_IN);
  not ginst21621 (P3_ADD_526_U29, P3_INSTADDRPOINTER_REG_18__SCAN_IN);
  not ginst21622 (P3_ADD_526_U30, P3_INSTADDRPOINTER_REG_17__SCAN_IN);
  nand ginst21623 (P3_ADD_526_U31, P3_ADD_526_U124, P3_ADD_526_U88);
  not ginst21624 (P3_ADD_526_U32, P3_INSTADDRPOINTER_REG_20__SCAN_IN);
  not ginst21625 (P3_ADD_526_U33, P3_INSTADDRPOINTER_REG_19__SCAN_IN);
  nand ginst21626 (P3_ADD_526_U34, P3_ADD_526_U117, P3_ADD_526_U89);
  not ginst21627 (P3_ADD_526_U35, P3_INSTADDRPOINTER_REG_21__SCAN_IN);
  nand ginst21628 (P3_ADD_526_U36, P3_ADD_526_U114, P3_ADD_526_U90);
  not ginst21629 (P3_ADD_526_U37, P3_INSTADDRPOINTER_REG_22__SCAN_IN);
  not ginst21630 (P3_ADD_526_U38, P3_INSTADDRPOINTER_REG_24__SCAN_IN);
  not ginst21631 (P3_ADD_526_U39, P3_INSTADDRPOINTER_REG_23__SCAN_IN);
  nand ginst21632 (P3_ADD_526_U40, P3_ADD_526_U121, P3_ADD_526_U91);
  not ginst21633 (P3_ADD_526_U41, P3_INSTADDRPOINTER_REG_26__SCAN_IN);
  not ginst21634 (P3_ADD_526_U42, P3_INSTADDRPOINTER_REG_25__SCAN_IN);
  nand ginst21635 (P3_ADD_526_U43, P3_ADD_526_U115, P3_ADD_526_U92);
  not ginst21636 (P3_ADD_526_U44, P3_INSTADDRPOINTER_REG_27__SCAN_IN);
  not ginst21637 (P3_ADD_526_U45, P3_INSTADDRPOINTER_REG_28__SCAN_IN);
  nand ginst21638 (P3_ADD_526_U46, P3_ADD_526_U116, P3_ADD_526_U93);
  not ginst21639 (P3_ADD_526_U47, P3_INSTADDRPOINTER_REG_29__SCAN_IN);
  nand ginst21640 (P3_ADD_526_U48, P3_ADD_526_U122, P3_ADD_526_U94);
  nand ginst21641 (P3_ADD_526_U49, P3_INSTADDRPOINTER_REG_29__SCAN_IN, P3_ADD_526_U123);
  not ginst21642 (P3_ADD_526_U5, P3_INSTADDRPOINTER_REG_0__SCAN_IN);
  not ginst21643 (P3_ADD_526_U50, P3_INSTADDRPOINTER_REG_30__SCAN_IN);
  nand ginst21644 (P3_ADD_526_U51, P3_ADD_526_U141, P3_ADD_526_U142);
  nand ginst21645 (P3_ADD_526_U52, P3_ADD_526_U143, P3_ADD_526_U144);
  nand ginst21646 (P3_ADD_526_U53, P3_ADD_526_U145, P3_ADD_526_U146);
  nand ginst21647 (P3_ADD_526_U54, P3_ADD_526_U147, P3_ADD_526_U148);
  nand ginst21648 (P3_ADD_526_U55, P3_ADD_526_U149, P3_ADD_526_U150);
  nand ginst21649 (P3_ADD_526_U56, P3_ADD_526_U151, P3_ADD_526_U152);
  nand ginst21650 (P3_ADD_526_U57, P3_ADD_526_U153, P3_ADD_526_U154);
  nand ginst21651 (P3_ADD_526_U58, P3_ADD_526_U155, P3_ADD_526_U156);
  nand ginst21652 (P3_ADD_526_U59, P3_ADD_526_U157, P3_ADD_526_U158);
  not ginst21653 (P3_ADD_526_U6, P3_INSTADDRPOINTER_REG_2__SCAN_IN);
  nand ginst21654 (P3_ADD_526_U60, P3_ADD_526_U159, P3_ADD_526_U160);
  nand ginst21655 (P3_ADD_526_U61, P3_ADD_526_U161, P3_ADD_526_U162);
  nand ginst21656 (P3_ADD_526_U62, P3_ADD_526_U163, P3_ADD_526_U164);
  nand ginst21657 (P3_ADD_526_U63, P3_ADD_526_U165, P3_ADD_526_U166);
  nand ginst21658 (P3_ADD_526_U64, P3_ADD_526_U167, P3_ADD_526_U168);
  nand ginst21659 (P3_ADD_526_U65, P3_ADD_526_U169, P3_ADD_526_U170);
  nand ginst21660 (P3_ADD_526_U66, P3_ADD_526_U171, P3_ADD_526_U172);
  nand ginst21661 (P3_ADD_526_U67, P3_ADD_526_U173, P3_ADD_526_U174);
  nand ginst21662 (P3_ADD_526_U68, P3_ADD_526_U175, P3_ADD_526_U176);
  nand ginst21663 (P3_ADD_526_U69, P3_ADD_526_U177, P3_ADD_526_U178);
  not ginst21664 (P3_ADD_526_U7, P3_INSTADDRPOINTER_REG_1__SCAN_IN);
  nand ginst21665 (P3_ADD_526_U70, P3_ADD_526_U179, P3_ADD_526_U180);
  nand ginst21666 (P3_ADD_526_U71, P3_ADD_526_U181, P3_ADD_526_U182);
  nand ginst21667 (P3_ADD_526_U72, P3_ADD_526_U183, P3_ADD_526_U184);
  nand ginst21668 (P3_ADD_526_U73, P3_ADD_526_U185, P3_ADD_526_U186);
  nand ginst21669 (P3_ADD_526_U74, P3_ADD_526_U187, P3_ADD_526_U188);
  nand ginst21670 (P3_ADD_526_U75, P3_ADD_526_U189, P3_ADD_526_U190);
  nand ginst21671 (P3_ADD_526_U76, P3_ADD_526_U191, P3_ADD_526_U192);
  nand ginst21672 (P3_ADD_526_U77, P3_ADD_526_U193, P3_ADD_526_U194);
  nand ginst21673 (P3_ADD_526_U78, P3_ADD_526_U195, P3_ADD_526_U196);
  nand ginst21674 (P3_ADD_526_U79, P3_ADD_526_U197, P3_ADD_526_U198);
  not ginst21675 (P3_ADD_526_U8, P3_INSTADDRPOINTER_REG_4__SCAN_IN);
  nand ginst21676 (P3_ADD_526_U80, P3_ADD_526_U199, P3_ADD_526_U200);
  nand ginst21677 (P3_ADD_526_U81, P3_ADD_526_U201, P3_ADD_526_U202);
  and ginst21678 (P3_ADD_526_U82, P3_INSTADDRPOINTER_REG_3__SCAN_IN, P3_INSTADDRPOINTER_REG_4__SCAN_IN);
  and ginst21679 (P3_ADD_526_U83, P3_INSTADDRPOINTER_REG_5__SCAN_IN, P3_INSTADDRPOINTER_REG_6__SCAN_IN);
  and ginst21680 (P3_ADD_526_U84, P3_INSTADDRPOINTER_REG_7__SCAN_IN, P3_INSTADDRPOINTER_REG_8__SCAN_IN);
  and ginst21681 (P3_ADD_526_U85, P3_INSTADDRPOINTER_REG_9__SCAN_IN, P3_INSTADDRPOINTER_REG_10__SCAN_IN);
  and ginst21682 (P3_ADD_526_U86, P3_INSTADDRPOINTER_REG_11__SCAN_IN, P3_INSTADDRPOINTER_REG_12__SCAN_IN);
  and ginst21683 (P3_ADD_526_U87, P3_INSTADDRPOINTER_REG_13__SCAN_IN, P3_INSTADDRPOINTER_REG_14__SCAN_IN);
  and ginst21684 (P3_ADD_526_U88, P3_INSTADDRPOINTER_REG_15__SCAN_IN, P3_INSTADDRPOINTER_REG_16__SCAN_IN);
  and ginst21685 (P3_ADD_526_U89, P3_INSTADDRPOINTER_REG_17__SCAN_IN, P3_INSTADDRPOINTER_REG_18__SCAN_IN);
  not ginst21686 (P3_ADD_526_U9, P3_INSTADDRPOINTER_REG_3__SCAN_IN);
  and ginst21687 (P3_ADD_526_U90, P3_INSTADDRPOINTER_REG_19__SCAN_IN, P3_INSTADDRPOINTER_REG_20__SCAN_IN);
  and ginst21688 (P3_ADD_526_U91, P3_INSTADDRPOINTER_REG_21__SCAN_IN, P3_INSTADDRPOINTER_REG_22__SCAN_IN);
  and ginst21689 (P3_ADD_526_U92, P3_INSTADDRPOINTER_REG_23__SCAN_IN, P3_INSTADDRPOINTER_REG_24__SCAN_IN);
  and ginst21690 (P3_ADD_526_U93, P3_INSTADDRPOINTER_REG_25__SCAN_IN, P3_INSTADDRPOINTER_REG_26__SCAN_IN);
  and ginst21691 (P3_ADD_526_U94, P3_INSTADDRPOINTER_REG_27__SCAN_IN, P3_INSTADDRPOINTER_REG_28__SCAN_IN);
  nand ginst21692 (P3_ADD_526_U95, P3_INSTADDRPOINTER_REG_7__SCAN_IN, P3_ADD_526_U118);
  nand ginst21693 (P3_ADD_526_U96, P3_INSTADDRPOINTER_REG_5__SCAN_IN, P3_ADD_526_U112);
  nand ginst21694 (P3_ADD_526_U97, P3_INSTADDRPOINTER_REG_3__SCAN_IN, P3_ADD_526_U111);
  not ginst21695 (P3_ADD_526_U98, P3_INSTADDRPOINTER_REG_31__SCAN_IN);
  nand ginst21696 (P3_ADD_526_U99, P3_INSTADDRPOINTER_REG_30__SCAN_IN, P3_ADD_526_U128);
  not ginst21697 (P3_ADD_531_U10, P3_INSTADDRPOINTER_REG_3__SCAN_IN);
  not ginst21698 (P3_ADD_531_U100, P3_ADD_531_U11);
  not ginst21699 (P3_ADD_531_U101, P3_ADD_531_U13);
  not ginst21700 (P3_ADD_531_U102, P3_ADD_531_U15);
  not ginst21701 (P3_ADD_531_U103, P3_ADD_531_U17);
  not ginst21702 (P3_ADD_531_U104, P3_ADD_531_U19);
  not ginst21703 (P3_ADD_531_U105, P3_ADD_531_U22);
  not ginst21704 (P3_ADD_531_U106, P3_ADD_531_U23);
  not ginst21705 (P3_ADD_531_U107, P3_ADD_531_U25);
  not ginst21706 (P3_ADD_531_U108, P3_ADD_531_U27);
  not ginst21707 (P3_ADD_531_U109, P3_ADD_531_U29);
  nand ginst21708 (P3_ADD_531_U11, P3_INSTADDRPOINTER_REG_3__SCAN_IN, P3_ADD_531_U99);
  not ginst21709 (P3_ADD_531_U110, P3_ADD_531_U31);
  not ginst21710 (P3_ADD_531_U111, P3_ADD_531_U33);
  not ginst21711 (P3_ADD_531_U112, P3_ADD_531_U35);
  not ginst21712 (P3_ADD_531_U113, P3_ADD_531_U37);
  not ginst21713 (P3_ADD_531_U114, P3_ADD_531_U39);
  not ginst21714 (P3_ADD_531_U115, P3_ADD_531_U41);
  not ginst21715 (P3_ADD_531_U116, P3_ADD_531_U43);
  not ginst21716 (P3_ADD_531_U117, P3_ADD_531_U45);
  not ginst21717 (P3_ADD_531_U118, P3_ADD_531_U47);
  not ginst21718 (P3_ADD_531_U119, P3_ADD_531_U49);
  not ginst21719 (P3_ADD_531_U12, P3_INSTADDRPOINTER_REG_4__SCAN_IN);
  not ginst21720 (P3_ADD_531_U120, P3_ADD_531_U51);
  not ginst21721 (P3_ADD_531_U121, P3_ADD_531_U53);
  not ginst21722 (P3_ADD_531_U122, P3_ADD_531_U55);
  not ginst21723 (P3_ADD_531_U123, P3_ADD_531_U57);
  not ginst21724 (P3_ADD_531_U124, P3_ADD_531_U59);
  not ginst21725 (P3_ADD_531_U125, P3_ADD_531_U61);
  not ginst21726 (P3_ADD_531_U126, P3_ADD_531_U63);
  not ginst21727 (P3_ADD_531_U127, P3_ADD_531_U97);
  nand ginst21728 (P3_ADD_531_U128, P3_INSTADDRPOINTER_REG_9__SCAN_IN, P3_ADD_531_U22);
  nand ginst21729 (P3_ADD_531_U129, P3_ADD_531_U105, P3_ADD_531_U21);
  nand ginst21730 (P3_ADD_531_U13, P3_INSTADDRPOINTER_REG_4__SCAN_IN, P3_ADD_531_U100);
  nand ginst21731 (P3_ADD_531_U130, P3_INSTADDRPOINTER_REG_8__SCAN_IN, P3_ADD_531_U19);
  nand ginst21732 (P3_ADD_531_U131, P3_ADD_531_U104, P3_ADD_531_U20);
  nand ginst21733 (P3_ADD_531_U132, P3_INSTADDRPOINTER_REG_7__SCAN_IN, P3_ADD_531_U17);
  nand ginst21734 (P3_ADD_531_U133, P3_ADD_531_U103, P3_ADD_531_U18);
  nand ginst21735 (P3_ADD_531_U134, P3_INSTADDRPOINTER_REG_6__SCAN_IN, P3_ADD_531_U15);
  nand ginst21736 (P3_ADD_531_U135, P3_ADD_531_U102, P3_ADD_531_U16);
  nand ginst21737 (P3_ADD_531_U136, P3_INSTADDRPOINTER_REG_5__SCAN_IN, P3_ADD_531_U13);
  nand ginst21738 (P3_ADD_531_U137, P3_ADD_531_U101, P3_ADD_531_U14);
  nand ginst21739 (P3_ADD_531_U138, P3_INSTADDRPOINTER_REG_4__SCAN_IN, P3_ADD_531_U11);
  nand ginst21740 (P3_ADD_531_U139, P3_ADD_531_U100, P3_ADD_531_U12);
  not ginst21741 (P3_ADD_531_U14, P3_INSTADDRPOINTER_REG_5__SCAN_IN);
  nand ginst21742 (P3_ADD_531_U140, P3_INSTADDRPOINTER_REG_3__SCAN_IN, P3_ADD_531_U9);
  nand ginst21743 (P3_ADD_531_U141, P3_ADD_531_U10, P3_ADD_531_U99);
  nand ginst21744 (P3_ADD_531_U142, P3_INSTADDRPOINTER_REG_31__SCAN_IN, P3_ADD_531_U97);
  nand ginst21745 (P3_ADD_531_U143, P3_ADD_531_U127, P3_ADD_531_U96);
  nand ginst21746 (P3_ADD_531_U144, P3_INSTADDRPOINTER_REG_30__SCAN_IN, P3_ADD_531_U63);
  nand ginst21747 (P3_ADD_531_U145, P3_ADD_531_U126, P3_ADD_531_U64);
  nand ginst21748 (P3_ADD_531_U146, P3_INSTADDRPOINTER_REG_2__SCAN_IN, P3_ADD_531_U7);
  nand ginst21749 (P3_ADD_531_U147, P3_ADD_531_U8, P3_ADD_531_U98);
  nand ginst21750 (P3_ADD_531_U148, P3_INSTADDRPOINTER_REG_29__SCAN_IN, P3_ADD_531_U61);
  nand ginst21751 (P3_ADD_531_U149, P3_ADD_531_U125, P3_ADD_531_U62);
  nand ginst21752 (P3_ADD_531_U15, P3_INSTADDRPOINTER_REG_5__SCAN_IN, P3_ADD_531_U101);
  nand ginst21753 (P3_ADD_531_U150, P3_INSTADDRPOINTER_REG_28__SCAN_IN, P3_ADD_531_U59);
  nand ginst21754 (P3_ADD_531_U151, P3_ADD_531_U124, P3_ADD_531_U60);
  nand ginst21755 (P3_ADD_531_U152, P3_INSTADDRPOINTER_REG_27__SCAN_IN, P3_ADD_531_U57);
  nand ginst21756 (P3_ADD_531_U153, P3_ADD_531_U123, P3_ADD_531_U58);
  nand ginst21757 (P3_ADD_531_U154, P3_INSTADDRPOINTER_REG_26__SCAN_IN, P3_ADD_531_U55);
  nand ginst21758 (P3_ADD_531_U155, P3_ADD_531_U122, P3_ADD_531_U56);
  nand ginst21759 (P3_ADD_531_U156, P3_INSTADDRPOINTER_REG_25__SCAN_IN, P3_ADD_531_U53);
  nand ginst21760 (P3_ADD_531_U157, P3_ADD_531_U121, P3_ADD_531_U54);
  nand ginst21761 (P3_ADD_531_U158, P3_INSTADDRPOINTER_REG_24__SCAN_IN, P3_ADD_531_U51);
  nand ginst21762 (P3_ADD_531_U159, P3_ADD_531_U120, P3_ADD_531_U52);
  not ginst21763 (P3_ADD_531_U16, P3_INSTADDRPOINTER_REG_6__SCAN_IN);
  nand ginst21764 (P3_ADD_531_U160, P3_INSTADDRPOINTER_REG_23__SCAN_IN, P3_ADD_531_U49);
  nand ginst21765 (P3_ADD_531_U161, P3_ADD_531_U119, P3_ADD_531_U50);
  nand ginst21766 (P3_ADD_531_U162, P3_INSTADDRPOINTER_REG_22__SCAN_IN, P3_ADD_531_U47);
  nand ginst21767 (P3_ADD_531_U163, P3_ADD_531_U118, P3_ADD_531_U48);
  nand ginst21768 (P3_ADD_531_U164, P3_INSTADDRPOINTER_REG_21__SCAN_IN, P3_ADD_531_U45);
  nand ginst21769 (P3_ADD_531_U165, P3_ADD_531_U117, P3_ADD_531_U46);
  nand ginst21770 (P3_ADD_531_U166, P3_INSTADDRPOINTER_REG_20__SCAN_IN, P3_ADD_531_U43);
  nand ginst21771 (P3_ADD_531_U167, P3_ADD_531_U116, P3_ADD_531_U44);
  nand ginst21772 (P3_ADD_531_U168, P3_INSTADDRPOINTER_REG_1__SCAN_IN, P3_ADD_531_U5);
  nand ginst21773 (P3_ADD_531_U169, P3_INSTADDRPOINTER_REG_0__SCAN_IN, P3_ADD_531_U6);
  nand ginst21774 (P3_ADD_531_U17, P3_INSTADDRPOINTER_REG_6__SCAN_IN, P3_ADD_531_U102);
  nand ginst21775 (P3_ADD_531_U170, P3_INSTADDRPOINTER_REG_19__SCAN_IN, P3_ADD_531_U41);
  nand ginst21776 (P3_ADD_531_U171, P3_ADD_531_U115, P3_ADD_531_U42);
  nand ginst21777 (P3_ADD_531_U172, P3_INSTADDRPOINTER_REG_18__SCAN_IN, P3_ADD_531_U39);
  nand ginst21778 (P3_ADD_531_U173, P3_ADD_531_U114, P3_ADD_531_U40);
  nand ginst21779 (P3_ADD_531_U174, P3_INSTADDRPOINTER_REG_17__SCAN_IN, P3_ADD_531_U37);
  nand ginst21780 (P3_ADD_531_U175, P3_ADD_531_U113, P3_ADD_531_U38);
  nand ginst21781 (P3_ADD_531_U176, P3_INSTADDRPOINTER_REG_16__SCAN_IN, P3_ADD_531_U35);
  nand ginst21782 (P3_ADD_531_U177, P3_ADD_531_U112, P3_ADD_531_U36);
  nand ginst21783 (P3_ADD_531_U178, P3_INSTADDRPOINTER_REG_15__SCAN_IN, P3_ADD_531_U33);
  nand ginst21784 (P3_ADD_531_U179, P3_ADD_531_U111, P3_ADD_531_U34);
  not ginst21785 (P3_ADD_531_U18, P3_INSTADDRPOINTER_REG_7__SCAN_IN);
  nand ginst21786 (P3_ADD_531_U180, P3_INSTADDRPOINTER_REG_14__SCAN_IN, P3_ADD_531_U31);
  nand ginst21787 (P3_ADD_531_U181, P3_ADD_531_U110, P3_ADD_531_U32);
  nand ginst21788 (P3_ADD_531_U182, P3_INSTADDRPOINTER_REG_13__SCAN_IN, P3_ADD_531_U29);
  nand ginst21789 (P3_ADD_531_U183, P3_ADD_531_U109, P3_ADD_531_U30);
  nand ginst21790 (P3_ADD_531_U184, P3_INSTADDRPOINTER_REG_12__SCAN_IN, P3_ADD_531_U27);
  nand ginst21791 (P3_ADD_531_U185, P3_ADD_531_U108, P3_ADD_531_U28);
  nand ginst21792 (P3_ADD_531_U186, P3_INSTADDRPOINTER_REG_11__SCAN_IN, P3_ADD_531_U25);
  nand ginst21793 (P3_ADD_531_U187, P3_ADD_531_U107, P3_ADD_531_U26);
  nand ginst21794 (P3_ADD_531_U188, P3_INSTADDRPOINTER_REG_10__SCAN_IN, P3_ADD_531_U23);
  nand ginst21795 (P3_ADD_531_U189, P3_ADD_531_U106, P3_ADD_531_U24);
  nand ginst21796 (P3_ADD_531_U19, P3_INSTADDRPOINTER_REG_7__SCAN_IN, P3_ADD_531_U103);
  not ginst21797 (P3_ADD_531_U20, P3_INSTADDRPOINTER_REG_8__SCAN_IN);
  not ginst21798 (P3_ADD_531_U21, P3_INSTADDRPOINTER_REG_9__SCAN_IN);
  nand ginst21799 (P3_ADD_531_U22, P3_INSTADDRPOINTER_REG_8__SCAN_IN, P3_ADD_531_U104);
  nand ginst21800 (P3_ADD_531_U23, P3_INSTADDRPOINTER_REG_9__SCAN_IN, P3_ADD_531_U105);
  not ginst21801 (P3_ADD_531_U24, P3_INSTADDRPOINTER_REG_10__SCAN_IN);
  nand ginst21802 (P3_ADD_531_U25, P3_INSTADDRPOINTER_REG_10__SCAN_IN, P3_ADD_531_U106);
  not ginst21803 (P3_ADD_531_U26, P3_INSTADDRPOINTER_REG_11__SCAN_IN);
  nand ginst21804 (P3_ADD_531_U27, P3_INSTADDRPOINTER_REG_11__SCAN_IN, P3_ADD_531_U107);
  not ginst21805 (P3_ADD_531_U28, P3_INSTADDRPOINTER_REG_12__SCAN_IN);
  nand ginst21806 (P3_ADD_531_U29, P3_INSTADDRPOINTER_REG_12__SCAN_IN, P3_ADD_531_U108);
  not ginst21807 (P3_ADD_531_U30, P3_INSTADDRPOINTER_REG_13__SCAN_IN);
  nand ginst21808 (P3_ADD_531_U31, P3_INSTADDRPOINTER_REG_13__SCAN_IN, P3_ADD_531_U109);
  not ginst21809 (P3_ADD_531_U32, P3_INSTADDRPOINTER_REG_14__SCAN_IN);
  nand ginst21810 (P3_ADD_531_U33, P3_INSTADDRPOINTER_REG_14__SCAN_IN, P3_ADD_531_U110);
  not ginst21811 (P3_ADD_531_U34, P3_INSTADDRPOINTER_REG_15__SCAN_IN);
  nand ginst21812 (P3_ADD_531_U35, P3_INSTADDRPOINTER_REG_15__SCAN_IN, P3_ADD_531_U111);
  not ginst21813 (P3_ADD_531_U36, P3_INSTADDRPOINTER_REG_16__SCAN_IN);
  nand ginst21814 (P3_ADD_531_U37, P3_INSTADDRPOINTER_REG_16__SCAN_IN, P3_ADD_531_U112);
  not ginst21815 (P3_ADD_531_U38, P3_INSTADDRPOINTER_REG_17__SCAN_IN);
  nand ginst21816 (P3_ADD_531_U39, P3_INSTADDRPOINTER_REG_17__SCAN_IN, P3_ADD_531_U113);
  not ginst21817 (P3_ADD_531_U40, P3_INSTADDRPOINTER_REG_18__SCAN_IN);
  nand ginst21818 (P3_ADD_531_U41, P3_INSTADDRPOINTER_REG_18__SCAN_IN, P3_ADD_531_U114);
  not ginst21819 (P3_ADD_531_U42, P3_INSTADDRPOINTER_REG_19__SCAN_IN);
  nand ginst21820 (P3_ADD_531_U43, P3_INSTADDRPOINTER_REG_19__SCAN_IN, P3_ADD_531_U115);
  not ginst21821 (P3_ADD_531_U44, P3_INSTADDRPOINTER_REG_20__SCAN_IN);
  nand ginst21822 (P3_ADD_531_U45, P3_INSTADDRPOINTER_REG_20__SCAN_IN, P3_ADD_531_U116);
  not ginst21823 (P3_ADD_531_U46, P3_INSTADDRPOINTER_REG_21__SCAN_IN);
  nand ginst21824 (P3_ADD_531_U47, P3_INSTADDRPOINTER_REG_21__SCAN_IN, P3_ADD_531_U117);
  not ginst21825 (P3_ADD_531_U48, P3_INSTADDRPOINTER_REG_22__SCAN_IN);
  nand ginst21826 (P3_ADD_531_U49, P3_INSTADDRPOINTER_REG_22__SCAN_IN, P3_ADD_531_U118);
  not ginst21827 (P3_ADD_531_U5, P3_INSTADDRPOINTER_REG_0__SCAN_IN);
  not ginst21828 (P3_ADD_531_U50, P3_INSTADDRPOINTER_REG_23__SCAN_IN);
  nand ginst21829 (P3_ADD_531_U51, P3_INSTADDRPOINTER_REG_23__SCAN_IN, P3_ADD_531_U119);
  not ginst21830 (P3_ADD_531_U52, P3_INSTADDRPOINTER_REG_24__SCAN_IN);
  nand ginst21831 (P3_ADD_531_U53, P3_INSTADDRPOINTER_REG_24__SCAN_IN, P3_ADD_531_U120);
  not ginst21832 (P3_ADD_531_U54, P3_INSTADDRPOINTER_REG_25__SCAN_IN);
  nand ginst21833 (P3_ADD_531_U55, P3_INSTADDRPOINTER_REG_25__SCAN_IN, P3_ADD_531_U121);
  not ginst21834 (P3_ADD_531_U56, P3_INSTADDRPOINTER_REG_26__SCAN_IN);
  nand ginst21835 (P3_ADD_531_U57, P3_INSTADDRPOINTER_REG_26__SCAN_IN, P3_ADD_531_U122);
  not ginst21836 (P3_ADD_531_U58, P3_INSTADDRPOINTER_REG_27__SCAN_IN);
  nand ginst21837 (P3_ADD_531_U59, P3_INSTADDRPOINTER_REG_27__SCAN_IN, P3_ADD_531_U123);
  not ginst21838 (P3_ADD_531_U6, P3_INSTADDRPOINTER_REG_1__SCAN_IN);
  not ginst21839 (P3_ADD_531_U60, P3_INSTADDRPOINTER_REG_28__SCAN_IN);
  nand ginst21840 (P3_ADD_531_U61, P3_INSTADDRPOINTER_REG_28__SCAN_IN, P3_ADD_531_U124);
  not ginst21841 (P3_ADD_531_U62, P3_INSTADDRPOINTER_REG_29__SCAN_IN);
  nand ginst21842 (P3_ADD_531_U63, P3_INSTADDRPOINTER_REG_29__SCAN_IN, P3_ADD_531_U125);
  not ginst21843 (P3_ADD_531_U64, P3_INSTADDRPOINTER_REG_30__SCAN_IN);
  nand ginst21844 (P3_ADD_531_U65, P3_ADD_531_U128, P3_ADD_531_U129);
  nand ginst21845 (P3_ADD_531_U66, P3_ADD_531_U130, P3_ADD_531_U131);
  nand ginst21846 (P3_ADD_531_U67, P3_ADD_531_U132, P3_ADD_531_U133);
  nand ginst21847 (P3_ADD_531_U68, P3_ADD_531_U134, P3_ADD_531_U135);
  nand ginst21848 (P3_ADD_531_U69, P3_ADD_531_U136, P3_ADD_531_U137);
  nand ginst21849 (P3_ADD_531_U7, P3_INSTADDRPOINTER_REG_0__SCAN_IN, P3_INSTADDRPOINTER_REG_1__SCAN_IN);
  nand ginst21850 (P3_ADD_531_U70, P3_ADD_531_U138, P3_ADD_531_U139);
  nand ginst21851 (P3_ADD_531_U71, P3_ADD_531_U140, P3_ADD_531_U141);
  nand ginst21852 (P3_ADD_531_U72, P3_ADD_531_U142, P3_ADD_531_U143);
  nand ginst21853 (P3_ADD_531_U73, P3_ADD_531_U144, P3_ADD_531_U145);
  nand ginst21854 (P3_ADD_531_U74, P3_ADD_531_U146, P3_ADD_531_U147);
  nand ginst21855 (P3_ADD_531_U75, P3_ADD_531_U148, P3_ADD_531_U149);
  nand ginst21856 (P3_ADD_531_U76, P3_ADD_531_U150, P3_ADD_531_U151);
  nand ginst21857 (P3_ADD_531_U77, P3_ADD_531_U152, P3_ADD_531_U153);
  nand ginst21858 (P3_ADD_531_U78, P3_ADD_531_U154, P3_ADD_531_U155);
  nand ginst21859 (P3_ADD_531_U79, P3_ADD_531_U156, P3_ADD_531_U157);
  not ginst21860 (P3_ADD_531_U8, P3_INSTADDRPOINTER_REG_2__SCAN_IN);
  nand ginst21861 (P3_ADD_531_U80, P3_ADD_531_U158, P3_ADD_531_U159);
  nand ginst21862 (P3_ADD_531_U81, P3_ADD_531_U160, P3_ADD_531_U161);
  nand ginst21863 (P3_ADD_531_U82, P3_ADD_531_U162, P3_ADD_531_U163);
  nand ginst21864 (P3_ADD_531_U83, P3_ADD_531_U164, P3_ADD_531_U165);
  nand ginst21865 (P3_ADD_531_U84, P3_ADD_531_U166, P3_ADD_531_U167);
  nand ginst21866 (P3_ADD_531_U85, P3_ADD_531_U168, P3_ADD_531_U169);
  nand ginst21867 (P3_ADD_531_U86, P3_ADD_531_U170, P3_ADD_531_U171);
  nand ginst21868 (P3_ADD_531_U87, P3_ADD_531_U172, P3_ADD_531_U173);
  nand ginst21869 (P3_ADD_531_U88, P3_ADD_531_U174, P3_ADD_531_U175);
  nand ginst21870 (P3_ADD_531_U89, P3_ADD_531_U176, P3_ADD_531_U177);
  nand ginst21871 (P3_ADD_531_U9, P3_INSTADDRPOINTER_REG_2__SCAN_IN, P3_ADD_531_U98);
  nand ginst21872 (P3_ADD_531_U90, P3_ADD_531_U178, P3_ADD_531_U179);
  nand ginst21873 (P3_ADD_531_U91, P3_ADD_531_U180, P3_ADD_531_U181);
  nand ginst21874 (P3_ADD_531_U92, P3_ADD_531_U182, P3_ADD_531_U183);
  nand ginst21875 (P3_ADD_531_U93, P3_ADD_531_U184, P3_ADD_531_U185);
  nand ginst21876 (P3_ADD_531_U94, P3_ADD_531_U186, P3_ADD_531_U187);
  nand ginst21877 (P3_ADD_531_U95, P3_ADD_531_U188, P3_ADD_531_U189);
  not ginst21878 (P3_ADD_531_U96, P3_INSTADDRPOINTER_REG_31__SCAN_IN);
  nand ginst21879 (P3_ADD_531_U97, P3_INSTADDRPOINTER_REG_30__SCAN_IN, P3_ADD_531_U126);
  not ginst21880 (P3_ADD_531_U98, P3_ADD_531_U7);
  not ginst21881 (P3_ADD_531_U99, P3_ADD_531_U9);
  nand ginst21882 (P3_ADD_536_U10, P3_INSTADDRPOINTER_REG_4__SCAN_IN, P3_ADD_536_U95);
  not ginst21883 (P3_ADD_536_U100, P3_ADD_536_U19);
  not ginst21884 (P3_ADD_536_U101, P3_ADD_536_U20);
  not ginst21885 (P3_ADD_536_U102, P3_ADD_536_U22);
  not ginst21886 (P3_ADD_536_U103, P3_ADD_536_U24);
  not ginst21887 (P3_ADD_536_U104, P3_ADD_536_U26);
  not ginst21888 (P3_ADD_536_U105, P3_ADD_536_U28);
  not ginst21889 (P3_ADD_536_U106, P3_ADD_536_U30);
  not ginst21890 (P3_ADD_536_U107, P3_ADD_536_U32);
  not ginst21891 (P3_ADD_536_U108, P3_ADD_536_U34);
  not ginst21892 (P3_ADD_536_U109, P3_ADD_536_U36);
  not ginst21893 (P3_ADD_536_U11, P3_INSTADDRPOINTER_REG_5__SCAN_IN);
  not ginst21894 (P3_ADD_536_U110, P3_ADD_536_U38);
  not ginst21895 (P3_ADD_536_U111, P3_ADD_536_U40);
  not ginst21896 (P3_ADD_536_U112, P3_ADD_536_U42);
  not ginst21897 (P3_ADD_536_U113, P3_ADD_536_U44);
  not ginst21898 (P3_ADD_536_U114, P3_ADD_536_U46);
  not ginst21899 (P3_ADD_536_U115, P3_ADD_536_U48);
  not ginst21900 (P3_ADD_536_U116, P3_ADD_536_U50);
  not ginst21901 (P3_ADD_536_U117, P3_ADD_536_U52);
  not ginst21902 (P3_ADD_536_U118, P3_ADD_536_U54);
  not ginst21903 (P3_ADD_536_U119, P3_ADD_536_U56);
  nand ginst21904 (P3_ADD_536_U12, P3_INSTADDRPOINTER_REG_5__SCAN_IN, P3_ADD_536_U96);
  not ginst21905 (P3_ADD_536_U120, P3_ADD_536_U58);
  not ginst21906 (P3_ADD_536_U121, P3_ADD_536_U60);
  not ginst21907 (P3_ADD_536_U122, P3_ADD_536_U93);
  nand ginst21908 (P3_ADD_536_U123, P3_INSTADDRPOINTER_REG_9__SCAN_IN, P3_ADD_536_U19);
  nand ginst21909 (P3_ADD_536_U124, P3_ADD_536_U100, P3_ADD_536_U18);
  nand ginst21910 (P3_ADD_536_U125, P3_INSTADDRPOINTER_REG_8__SCAN_IN, P3_ADD_536_U16);
  nand ginst21911 (P3_ADD_536_U126, P3_ADD_536_U17, P3_ADD_536_U99);
  nand ginst21912 (P3_ADD_536_U127, P3_INSTADDRPOINTER_REG_7__SCAN_IN, P3_ADD_536_U14);
  nand ginst21913 (P3_ADD_536_U128, P3_ADD_536_U15, P3_ADD_536_U98);
  nand ginst21914 (P3_ADD_536_U129, P3_INSTADDRPOINTER_REG_6__SCAN_IN, P3_ADD_536_U12);
  not ginst21915 (P3_ADD_536_U13, P3_INSTADDRPOINTER_REG_6__SCAN_IN);
  nand ginst21916 (P3_ADD_536_U130, P3_ADD_536_U13, P3_ADD_536_U97);
  nand ginst21917 (P3_ADD_536_U131, P3_INSTADDRPOINTER_REG_5__SCAN_IN, P3_ADD_536_U10);
  nand ginst21918 (P3_ADD_536_U132, P3_ADD_536_U11, P3_ADD_536_U96);
  nand ginst21919 (P3_ADD_536_U133, P3_INSTADDRPOINTER_REG_4__SCAN_IN, P3_ADD_536_U8);
  nand ginst21920 (P3_ADD_536_U134, P3_ADD_536_U9, P3_ADD_536_U95);
  nand ginst21921 (P3_ADD_536_U135, P3_INSTADDRPOINTER_REG_3__SCAN_IN, P3_ADD_536_U6);
  nand ginst21922 (P3_ADD_536_U136, P3_ADD_536_U7, P3_ADD_536_U94);
  nand ginst21923 (P3_ADD_536_U137, P3_INSTADDRPOINTER_REG_31__SCAN_IN, P3_ADD_536_U93);
  nand ginst21924 (P3_ADD_536_U138, P3_ADD_536_U122, P3_ADD_536_U92);
  nand ginst21925 (P3_ADD_536_U139, P3_INSTADDRPOINTER_REG_30__SCAN_IN, P3_ADD_536_U60);
  nand ginst21926 (P3_ADD_536_U14, P3_INSTADDRPOINTER_REG_6__SCAN_IN, P3_ADD_536_U97);
  nand ginst21927 (P3_ADD_536_U140, P3_ADD_536_U121, P3_ADD_536_U61);
  nand ginst21928 (P3_ADD_536_U141, P3_INSTADDRPOINTER_REG_2__SCAN_IN, P3_ADD_536_U4);
  nand ginst21929 (P3_ADD_536_U142, P3_INSTADDRPOINTER_REG_1__SCAN_IN, P3_ADD_536_U5);
  nand ginst21930 (P3_ADD_536_U143, P3_INSTADDRPOINTER_REG_29__SCAN_IN, P3_ADD_536_U58);
  nand ginst21931 (P3_ADD_536_U144, P3_ADD_536_U120, P3_ADD_536_U59);
  nand ginst21932 (P3_ADD_536_U145, P3_INSTADDRPOINTER_REG_28__SCAN_IN, P3_ADD_536_U56);
  nand ginst21933 (P3_ADD_536_U146, P3_ADD_536_U119, P3_ADD_536_U57);
  nand ginst21934 (P3_ADD_536_U147, P3_INSTADDRPOINTER_REG_27__SCAN_IN, P3_ADD_536_U54);
  nand ginst21935 (P3_ADD_536_U148, P3_ADD_536_U118, P3_ADD_536_U55);
  nand ginst21936 (P3_ADD_536_U149, P3_INSTADDRPOINTER_REG_26__SCAN_IN, P3_ADD_536_U52);
  not ginst21937 (P3_ADD_536_U15, P3_INSTADDRPOINTER_REG_7__SCAN_IN);
  nand ginst21938 (P3_ADD_536_U150, P3_ADD_536_U117, P3_ADD_536_U53);
  nand ginst21939 (P3_ADD_536_U151, P3_INSTADDRPOINTER_REG_25__SCAN_IN, P3_ADD_536_U50);
  nand ginst21940 (P3_ADD_536_U152, P3_ADD_536_U116, P3_ADD_536_U51);
  nand ginst21941 (P3_ADD_536_U153, P3_INSTADDRPOINTER_REG_24__SCAN_IN, P3_ADD_536_U48);
  nand ginst21942 (P3_ADD_536_U154, P3_ADD_536_U115, P3_ADD_536_U49);
  nand ginst21943 (P3_ADD_536_U155, P3_INSTADDRPOINTER_REG_23__SCAN_IN, P3_ADD_536_U46);
  nand ginst21944 (P3_ADD_536_U156, P3_ADD_536_U114, P3_ADD_536_U47);
  nand ginst21945 (P3_ADD_536_U157, P3_INSTADDRPOINTER_REG_22__SCAN_IN, P3_ADD_536_U44);
  nand ginst21946 (P3_ADD_536_U158, P3_ADD_536_U113, P3_ADD_536_U45);
  nand ginst21947 (P3_ADD_536_U159, P3_INSTADDRPOINTER_REG_21__SCAN_IN, P3_ADD_536_U42);
  nand ginst21948 (P3_ADD_536_U16, P3_INSTADDRPOINTER_REG_7__SCAN_IN, P3_ADD_536_U98);
  nand ginst21949 (P3_ADD_536_U160, P3_ADD_536_U112, P3_ADD_536_U43);
  nand ginst21950 (P3_ADD_536_U161, P3_INSTADDRPOINTER_REG_20__SCAN_IN, P3_ADD_536_U40);
  nand ginst21951 (P3_ADD_536_U162, P3_ADD_536_U111, P3_ADD_536_U41);
  nand ginst21952 (P3_ADD_536_U163, P3_INSTADDRPOINTER_REG_19__SCAN_IN, P3_ADD_536_U38);
  nand ginst21953 (P3_ADD_536_U164, P3_ADD_536_U110, P3_ADD_536_U39);
  nand ginst21954 (P3_ADD_536_U165, P3_INSTADDRPOINTER_REG_18__SCAN_IN, P3_ADD_536_U36);
  nand ginst21955 (P3_ADD_536_U166, P3_ADD_536_U109, P3_ADD_536_U37);
  nand ginst21956 (P3_ADD_536_U167, P3_INSTADDRPOINTER_REG_17__SCAN_IN, P3_ADD_536_U34);
  nand ginst21957 (P3_ADD_536_U168, P3_ADD_536_U108, P3_ADD_536_U35);
  nand ginst21958 (P3_ADD_536_U169, P3_INSTADDRPOINTER_REG_16__SCAN_IN, P3_ADD_536_U32);
  not ginst21959 (P3_ADD_536_U17, P3_INSTADDRPOINTER_REG_8__SCAN_IN);
  nand ginst21960 (P3_ADD_536_U170, P3_ADD_536_U107, P3_ADD_536_U33);
  nand ginst21961 (P3_ADD_536_U171, P3_INSTADDRPOINTER_REG_15__SCAN_IN, P3_ADD_536_U30);
  nand ginst21962 (P3_ADD_536_U172, P3_ADD_536_U106, P3_ADD_536_U31);
  nand ginst21963 (P3_ADD_536_U173, P3_INSTADDRPOINTER_REG_14__SCAN_IN, P3_ADD_536_U28);
  nand ginst21964 (P3_ADD_536_U174, P3_ADD_536_U105, P3_ADD_536_U29);
  nand ginst21965 (P3_ADD_536_U175, P3_INSTADDRPOINTER_REG_13__SCAN_IN, P3_ADD_536_U26);
  nand ginst21966 (P3_ADD_536_U176, P3_ADD_536_U104, P3_ADD_536_U27);
  nand ginst21967 (P3_ADD_536_U177, P3_INSTADDRPOINTER_REG_12__SCAN_IN, P3_ADD_536_U24);
  nand ginst21968 (P3_ADD_536_U178, P3_ADD_536_U103, P3_ADD_536_U25);
  nand ginst21969 (P3_ADD_536_U179, P3_INSTADDRPOINTER_REG_11__SCAN_IN, P3_ADD_536_U22);
  not ginst21970 (P3_ADD_536_U18, P3_INSTADDRPOINTER_REG_9__SCAN_IN);
  nand ginst21971 (P3_ADD_536_U180, P3_ADD_536_U102, P3_ADD_536_U23);
  nand ginst21972 (P3_ADD_536_U181, P3_INSTADDRPOINTER_REG_10__SCAN_IN, P3_ADD_536_U20);
  nand ginst21973 (P3_ADD_536_U182, P3_ADD_536_U101, P3_ADD_536_U21);
  nand ginst21974 (P3_ADD_536_U19, P3_INSTADDRPOINTER_REG_8__SCAN_IN, P3_ADD_536_U99);
  nand ginst21975 (P3_ADD_536_U20, P3_INSTADDRPOINTER_REG_9__SCAN_IN, P3_ADD_536_U100);
  not ginst21976 (P3_ADD_536_U21, P3_INSTADDRPOINTER_REG_10__SCAN_IN);
  nand ginst21977 (P3_ADD_536_U22, P3_INSTADDRPOINTER_REG_10__SCAN_IN, P3_ADD_536_U101);
  not ginst21978 (P3_ADD_536_U23, P3_INSTADDRPOINTER_REG_11__SCAN_IN);
  nand ginst21979 (P3_ADD_536_U24, P3_INSTADDRPOINTER_REG_11__SCAN_IN, P3_ADD_536_U102);
  not ginst21980 (P3_ADD_536_U25, P3_INSTADDRPOINTER_REG_12__SCAN_IN);
  nand ginst21981 (P3_ADD_536_U26, P3_INSTADDRPOINTER_REG_12__SCAN_IN, P3_ADD_536_U103);
  not ginst21982 (P3_ADD_536_U27, P3_INSTADDRPOINTER_REG_13__SCAN_IN);
  nand ginst21983 (P3_ADD_536_U28, P3_INSTADDRPOINTER_REG_13__SCAN_IN, P3_ADD_536_U104);
  not ginst21984 (P3_ADD_536_U29, P3_INSTADDRPOINTER_REG_14__SCAN_IN);
  nand ginst21985 (P3_ADD_536_U30, P3_INSTADDRPOINTER_REG_14__SCAN_IN, P3_ADD_536_U105);
  not ginst21986 (P3_ADD_536_U31, P3_INSTADDRPOINTER_REG_15__SCAN_IN);
  nand ginst21987 (P3_ADD_536_U32, P3_INSTADDRPOINTER_REG_15__SCAN_IN, P3_ADD_536_U106);
  not ginst21988 (P3_ADD_536_U33, P3_INSTADDRPOINTER_REG_16__SCAN_IN);
  nand ginst21989 (P3_ADD_536_U34, P3_INSTADDRPOINTER_REG_16__SCAN_IN, P3_ADD_536_U107);
  not ginst21990 (P3_ADD_536_U35, P3_INSTADDRPOINTER_REG_17__SCAN_IN);
  nand ginst21991 (P3_ADD_536_U36, P3_INSTADDRPOINTER_REG_17__SCAN_IN, P3_ADD_536_U108);
  not ginst21992 (P3_ADD_536_U37, P3_INSTADDRPOINTER_REG_18__SCAN_IN);
  nand ginst21993 (P3_ADD_536_U38, P3_INSTADDRPOINTER_REG_18__SCAN_IN, P3_ADD_536_U109);
  not ginst21994 (P3_ADD_536_U39, P3_INSTADDRPOINTER_REG_19__SCAN_IN);
  not ginst21995 (P3_ADD_536_U4, P3_INSTADDRPOINTER_REG_1__SCAN_IN);
  nand ginst21996 (P3_ADD_536_U40, P3_INSTADDRPOINTER_REG_19__SCAN_IN, P3_ADD_536_U110);
  not ginst21997 (P3_ADD_536_U41, P3_INSTADDRPOINTER_REG_20__SCAN_IN);
  nand ginst21998 (P3_ADD_536_U42, P3_INSTADDRPOINTER_REG_20__SCAN_IN, P3_ADD_536_U111);
  not ginst21999 (P3_ADD_536_U43, P3_INSTADDRPOINTER_REG_21__SCAN_IN);
  nand ginst22000 (P3_ADD_536_U44, P3_INSTADDRPOINTER_REG_21__SCAN_IN, P3_ADD_536_U112);
  not ginst22001 (P3_ADD_536_U45, P3_INSTADDRPOINTER_REG_22__SCAN_IN);
  nand ginst22002 (P3_ADD_536_U46, P3_INSTADDRPOINTER_REG_22__SCAN_IN, P3_ADD_536_U113);
  not ginst22003 (P3_ADD_536_U47, P3_INSTADDRPOINTER_REG_23__SCAN_IN);
  nand ginst22004 (P3_ADD_536_U48, P3_INSTADDRPOINTER_REG_23__SCAN_IN, P3_ADD_536_U114);
  not ginst22005 (P3_ADD_536_U49, P3_INSTADDRPOINTER_REG_24__SCAN_IN);
  not ginst22006 (P3_ADD_536_U5, P3_INSTADDRPOINTER_REG_2__SCAN_IN);
  nand ginst22007 (P3_ADD_536_U50, P3_INSTADDRPOINTER_REG_24__SCAN_IN, P3_ADD_536_U115);
  not ginst22008 (P3_ADD_536_U51, P3_INSTADDRPOINTER_REG_25__SCAN_IN);
  nand ginst22009 (P3_ADD_536_U52, P3_INSTADDRPOINTER_REG_25__SCAN_IN, P3_ADD_536_U116);
  not ginst22010 (P3_ADD_536_U53, P3_INSTADDRPOINTER_REG_26__SCAN_IN);
  nand ginst22011 (P3_ADD_536_U54, P3_INSTADDRPOINTER_REG_26__SCAN_IN, P3_ADD_536_U117);
  not ginst22012 (P3_ADD_536_U55, P3_INSTADDRPOINTER_REG_27__SCAN_IN);
  nand ginst22013 (P3_ADD_536_U56, P3_INSTADDRPOINTER_REG_27__SCAN_IN, P3_ADD_536_U118);
  not ginst22014 (P3_ADD_536_U57, P3_INSTADDRPOINTER_REG_28__SCAN_IN);
  nand ginst22015 (P3_ADD_536_U58, P3_INSTADDRPOINTER_REG_28__SCAN_IN, P3_ADD_536_U119);
  not ginst22016 (P3_ADD_536_U59, P3_INSTADDRPOINTER_REG_29__SCAN_IN);
  nand ginst22017 (P3_ADD_536_U6, P3_INSTADDRPOINTER_REG_1__SCAN_IN, P3_INSTADDRPOINTER_REG_2__SCAN_IN);
  nand ginst22018 (P3_ADD_536_U60, P3_INSTADDRPOINTER_REG_29__SCAN_IN, P3_ADD_536_U120);
  not ginst22019 (P3_ADD_536_U61, P3_INSTADDRPOINTER_REG_30__SCAN_IN);
  nand ginst22020 (P3_ADD_536_U62, P3_ADD_536_U123, P3_ADD_536_U124);
  nand ginst22021 (P3_ADD_536_U63, P3_ADD_536_U125, P3_ADD_536_U126);
  nand ginst22022 (P3_ADD_536_U64, P3_ADD_536_U127, P3_ADD_536_U128);
  nand ginst22023 (P3_ADD_536_U65, P3_ADD_536_U129, P3_ADD_536_U130);
  nand ginst22024 (P3_ADD_536_U66, P3_ADD_536_U131, P3_ADD_536_U132);
  nand ginst22025 (P3_ADD_536_U67, P3_ADD_536_U133, P3_ADD_536_U134);
  nand ginst22026 (P3_ADD_536_U68, P3_ADD_536_U135, P3_ADD_536_U136);
  nand ginst22027 (P3_ADD_536_U69, P3_ADD_536_U137, P3_ADD_536_U138);
  not ginst22028 (P3_ADD_536_U7, P3_INSTADDRPOINTER_REG_3__SCAN_IN);
  nand ginst22029 (P3_ADD_536_U70, P3_ADD_536_U139, P3_ADD_536_U140);
  nand ginst22030 (P3_ADD_536_U71, P3_ADD_536_U141, P3_ADD_536_U142);
  nand ginst22031 (P3_ADD_536_U72, P3_ADD_536_U143, P3_ADD_536_U144);
  nand ginst22032 (P3_ADD_536_U73, P3_ADD_536_U145, P3_ADD_536_U146);
  nand ginst22033 (P3_ADD_536_U74, P3_ADD_536_U147, P3_ADD_536_U148);
  nand ginst22034 (P3_ADD_536_U75, P3_ADD_536_U149, P3_ADD_536_U150);
  nand ginst22035 (P3_ADD_536_U76, P3_ADD_536_U151, P3_ADD_536_U152);
  nand ginst22036 (P3_ADD_536_U77, P3_ADD_536_U153, P3_ADD_536_U154);
  nand ginst22037 (P3_ADD_536_U78, P3_ADD_536_U155, P3_ADD_536_U156);
  nand ginst22038 (P3_ADD_536_U79, P3_ADD_536_U157, P3_ADD_536_U158);
  nand ginst22039 (P3_ADD_536_U8, P3_INSTADDRPOINTER_REG_3__SCAN_IN, P3_ADD_536_U94);
  nand ginst22040 (P3_ADD_536_U80, P3_ADD_536_U159, P3_ADD_536_U160);
  nand ginst22041 (P3_ADD_536_U81, P3_ADD_536_U161, P3_ADD_536_U162);
  nand ginst22042 (P3_ADD_536_U82, P3_ADD_536_U163, P3_ADD_536_U164);
  nand ginst22043 (P3_ADD_536_U83, P3_ADD_536_U165, P3_ADD_536_U166);
  nand ginst22044 (P3_ADD_536_U84, P3_ADD_536_U167, P3_ADD_536_U168);
  nand ginst22045 (P3_ADD_536_U85, P3_ADD_536_U169, P3_ADD_536_U170);
  nand ginst22046 (P3_ADD_536_U86, P3_ADD_536_U171, P3_ADD_536_U172);
  nand ginst22047 (P3_ADD_536_U87, P3_ADD_536_U173, P3_ADD_536_U174);
  nand ginst22048 (P3_ADD_536_U88, P3_ADD_536_U175, P3_ADD_536_U176);
  nand ginst22049 (P3_ADD_536_U89, P3_ADD_536_U177, P3_ADD_536_U178);
  not ginst22050 (P3_ADD_536_U9, P3_INSTADDRPOINTER_REG_4__SCAN_IN);
  nand ginst22051 (P3_ADD_536_U90, P3_ADD_536_U179, P3_ADD_536_U180);
  nand ginst22052 (P3_ADD_536_U91, P3_ADD_536_U181, P3_ADD_536_U182);
  not ginst22053 (P3_ADD_536_U92, P3_INSTADDRPOINTER_REG_31__SCAN_IN);
  nand ginst22054 (P3_ADD_536_U93, P3_INSTADDRPOINTER_REG_30__SCAN_IN, P3_ADD_536_U121);
  not ginst22055 (P3_ADD_536_U94, P3_ADD_536_U6);
  not ginst22056 (P3_ADD_536_U95, P3_ADD_536_U8);
  not ginst22057 (P3_ADD_536_U96, P3_ADD_536_U10);
  not ginst22058 (P3_ADD_536_U97, P3_ADD_536_U12);
  not ginst22059 (P3_ADD_536_U98, P3_ADD_536_U14);
  not ginst22060 (P3_ADD_536_U99, P3_ADD_536_U16);
  nand ginst22061 (P3_ADD_541_U10, P3_INSTADDRPOINTER_REG_4__SCAN_IN, P3_ADD_541_U95);
  not ginst22062 (P3_ADD_541_U100, P3_ADD_541_U19);
  not ginst22063 (P3_ADD_541_U101, P3_ADD_541_U20);
  not ginst22064 (P3_ADD_541_U102, P3_ADD_541_U22);
  not ginst22065 (P3_ADD_541_U103, P3_ADD_541_U24);
  not ginst22066 (P3_ADD_541_U104, P3_ADD_541_U26);
  not ginst22067 (P3_ADD_541_U105, P3_ADD_541_U28);
  not ginst22068 (P3_ADD_541_U106, P3_ADD_541_U30);
  not ginst22069 (P3_ADD_541_U107, P3_ADD_541_U32);
  not ginst22070 (P3_ADD_541_U108, P3_ADD_541_U34);
  not ginst22071 (P3_ADD_541_U109, P3_ADD_541_U36);
  not ginst22072 (P3_ADD_541_U11, P3_INSTADDRPOINTER_REG_5__SCAN_IN);
  not ginst22073 (P3_ADD_541_U110, P3_ADD_541_U38);
  not ginst22074 (P3_ADD_541_U111, P3_ADD_541_U40);
  not ginst22075 (P3_ADD_541_U112, P3_ADD_541_U42);
  not ginst22076 (P3_ADD_541_U113, P3_ADD_541_U44);
  not ginst22077 (P3_ADD_541_U114, P3_ADD_541_U46);
  not ginst22078 (P3_ADD_541_U115, P3_ADD_541_U48);
  not ginst22079 (P3_ADD_541_U116, P3_ADD_541_U50);
  not ginst22080 (P3_ADD_541_U117, P3_ADD_541_U52);
  not ginst22081 (P3_ADD_541_U118, P3_ADD_541_U54);
  not ginst22082 (P3_ADD_541_U119, P3_ADD_541_U56);
  nand ginst22083 (P3_ADD_541_U12, P3_INSTADDRPOINTER_REG_5__SCAN_IN, P3_ADD_541_U96);
  not ginst22084 (P3_ADD_541_U120, P3_ADD_541_U58);
  not ginst22085 (P3_ADD_541_U121, P3_ADD_541_U60);
  not ginst22086 (P3_ADD_541_U122, P3_ADD_541_U93);
  nand ginst22087 (P3_ADD_541_U123, P3_INSTADDRPOINTER_REG_9__SCAN_IN, P3_ADD_541_U19);
  nand ginst22088 (P3_ADD_541_U124, P3_ADD_541_U100, P3_ADD_541_U18);
  nand ginst22089 (P3_ADD_541_U125, P3_INSTADDRPOINTER_REG_8__SCAN_IN, P3_ADD_541_U16);
  nand ginst22090 (P3_ADD_541_U126, P3_ADD_541_U17, P3_ADD_541_U99);
  nand ginst22091 (P3_ADD_541_U127, P3_INSTADDRPOINTER_REG_7__SCAN_IN, P3_ADD_541_U14);
  nand ginst22092 (P3_ADD_541_U128, P3_ADD_541_U15, P3_ADD_541_U98);
  nand ginst22093 (P3_ADD_541_U129, P3_INSTADDRPOINTER_REG_6__SCAN_IN, P3_ADD_541_U12);
  not ginst22094 (P3_ADD_541_U13, P3_INSTADDRPOINTER_REG_6__SCAN_IN);
  nand ginst22095 (P3_ADD_541_U130, P3_ADD_541_U13, P3_ADD_541_U97);
  nand ginst22096 (P3_ADD_541_U131, P3_INSTADDRPOINTER_REG_5__SCAN_IN, P3_ADD_541_U10);
  nand ginst22097 (P3_ADD_541_U132, P3_ADD_541_U11, P3_ADD_541_U96);
  nand ginst22098 (P3_ADD_541_U133, P3_INSTADDRPOINTER_REG_4__SCAN_IN, P3_ADD_541_U8);
  nand ginst22099 (P3_ADD_541_U134, P3_ADD_541_U9, P3_ADD_541_U95);
  nand ginst22100 (P3_ADD_541_U135, P3_INSTADDRPOINTER_REG_3__SCAN_IN, P3_ADD_541_U6);
  nand ginst22101 (P3_ADD_541_U136, P3_ADD_541_U7, P3_ADD_541_U94);
  nand ginst22102 (P3_ADD_541_U137, P3_INSTADDRPOINTER_REG_31__SCAN_IN, P3_ADD_541_U93);
  nand ginst22103 (P3_ADD_541_U138, P3_ADD_541_U122, P3_ADD_541_U92);
  nand ginst22104 (P3_ADD_541_U139, P3_INSTADDRPOINTER_REG_30__SCAN_IN, P3_ADD_541_U60);
  nand ginst22105 (P3_ADD_541_U14, P3_INSTADDRPOINTER_REG_6__SCAN_IN, P3_ADD_541_U97);
  nand ginst22106 (P3_ADD_541_U140, P3_ADD_541_U121, P3_ADD_541_U61);
  nand ginst22107 (P3_ADD_541_U141, P3_INSTADDRPOINTER_REG_2__SCAN_IN, P3_ADD_541_U4);
  nand ginst22108 (P3_ADD_541_U142, P3_INSTADDRPOINTER_REG_1__SCAN_IN, P3_ADD_541_U5);
  nand ginst22109 (P3_ADD_541_U143, P3_INSTADDRPOINTER_REG_29__SCAN_IN, P3_ADD_541_U58);
  nand ginst22110 (P3_ADD_541_U144, P3_ADD_541_U120, P3_ADD_541_U59);
  nand ginst22111 (P3_ADD_541_U145, P3_INSTADDRPOINTER_REG_28__SCAN_IN, P3_ADD_541_U56);
  nand ginst22112 (P3_ADD_541_U146, P3_ADD_541_U119, P3_ADD_541_U57);
  nand ginst22113 (P3_ADD_541_U147, P3_INSTADDRPOINTER_REG_27__SCAN_IN, P3_ADD_541_U54);
  nand ginst22114 (P3_ADD_541_U148, P3_ADD_541_U118, P3_ADD_541_U55);
  nand ginst22115 (P3_ADD_541_U149, P3_INSTADDRPOINTER_REG_26__SCAN_IN, P3_ADD_541_U52);
  not ginst22116 (P3_ADD_541_U15, P3_INSTADDRPOINTER_REG_7__SCAN_IN);
  nand ginst22117 (P3_ADD_541_U150, P3_ADD_541_U117, P3_ADD_541_U53);
  nand ginst22118 (P3_ADD_541_U151, P3_INSTADDRPOINTER_REG_25__SCAN_IN, P3_ADD_541_U50);
  nand ginst22119 (P3_ADD_541_U152, P3_ADD_541_U116, P3_ADD_541_U51);
  nand ginst22120 (P3_ADD_541_U153, P3_INSTADDRPOINTER_REG_24__SCAN_IN, P3_ADD_541_U48);
  nand ginst22121 (P3_ADD_541_U154, P3_ADD_541_U115, P3_ADD_541_U49);
  nand ginst22122 (P3_ADD_541_U155, P3_INSTADDRPOINTER_REG_23__SCAN_IN, P3_ADD_541_U46);
  nand ginst22123 (P3_ADD_541_U156, P3_ADD_541_U114, P3_ADD_541_U47);
  nand ginst22124 (P3_ADD_541_U157, P3_INSTADDRPOINTER_REG_22__SCAN_IN, P3_ADD_541_U44);
  nand ginst22125 (P3_ADD_541_U158, P3_ADD_541_U113, P3_ADD_541_U45);
  nand ginst22126 (P3_ADD_541_U159, P3_INSTADDRPOINTER_REG_21__SCAN_IN, P3_ADD_541_U42);
  nand ginst22127 (P3_ADD_541_U16, P3_INSTADDRPOINTER_REG_7__SCAN_IN, P3_ADD_541_U98);
  nand ginst22128 (P3_ADD_541_U160, P3_ADD_541_U112, P3_ADD_541_U43);
  nand ginst22129 (P3_ADD_541_U161, P3_INSTADDRPOINTER_REG_20__SCAN_IN, P3_ADD_541_U40);
  nand ginst22130 (P3_ADD_541_U162, P3_ADD_541_U111, P3_ADD_541_U41);
  nand ginst22131 (P3_ADD_541_U163, P3_INSTADDRPOINTER_REG_19__SCAN_IN, P3_ADD_541_U38);
  nand ginst22132 (P3_ADD_541_U164, P3_ADD_541_U110, P3_ADD_541_U39);
  nand ginst22133 (P3_ADD_541_U165, P3_INSTADDRPOINTER_REG_18__SCAN_IN, P3_ADD_541_U36);
  nand ginst22134 (P3_ADD_541_U166, P3_ADD_541_U109, P3_ADD_541_U37);
  nand ginst22135 (P3_ADD_541_U167, P3_INSTADDRPOINTER_REG_17__SCAN_IN, P3_ADD_541_U34);
  nand ginst22136 (P3_ADD_541_U168, P3_ADD_541_U108, P3_ADD_541_U35);
  nand ginst22137 (P3_ADD_541_U169, P3_INSTADDRPOINTER_REG_16__SCAN_IN, P3_ADD_541_U32);
  not ginst22138 (P3_ADD_541_U17, P3_INSTADDRPOINTER_REG_8__SCAN_IN);
  nand ginst22139 (P3_ADD_541_U170, P3_ADD_541_U107, P3_ADD_541_U33);
  nand ginst22140 (P3_ADD_541_U171, P3_INSTADDRPOINTER_REG_15__SCAN_IN, P3_ADD_541_U30);
  nand ginst22141 (P3_ADD_541_U172, P3_ADD_541_U106, P3_ADD_541_U31);
  nand ginst22142 (P3_ADD_541_U173, P3_INSTADDRPOINTER_REG_14__SCAN_IN, P3_ADD_541_U28);
  nand ginst22143 (P3_ADD_541_U174, P3_ADD_541_U105, P3_ADD_541_U29);
  nand ginst22144 (P3_ADD_541_U175, P3_INSTADDRPOINTER_REG_13__SCAN_IN, P3_ADD_541_U26);
  nand ginst22145 (P3_ADD_541_U176, P3_ADD_541_U104, P3_ADD_541_U27);
  nand ginst22146 (P3_ADD_541_U177, P3_INSTADDRPOINTER_REG_12__SCAN_IN, P3_ADD_541_U24);
  nand ginst22147 (P3_ADD_541_U178, P3_ADD_541_U103, P3_ADD_541_U25);
  nand ginst22148 (P3_ADD_541_U179, P3_INSTADDRPOINTER_REG_11__SCAN_IN, P3_ADD_541_U22);
  not ginst22149 (P3_ADD_541_U18, P3_INSTADDRPOINTER_REG_9__SCAN_IN);
  nand ginst22150 (P3_ADD_541_U180, P3_ADD_541_U102, P3_ADD_541_U23);
  nand ginst22151 (P3_ADD_541_U181, P3_INSTADDRPOINTER_REG_10__SCAN_IN, P3_ADD_541_U20);
  nand ginst22152 (P3_ADD_541_U182, P3_ADD_541_U101, P3_ADD_541_U21);
  nand ginst22153 (P3_ADD_541_U19, P3_INSTADDRPOINTER_REG_8__SCAN_IN, P3_ADD_541_U99);
  nand ginst22154 (P3_ADD_541_U20, P3_INSTADDRPOINTER_REG_9__SCAN_IN, P3_ADD_541_U100);
  not ginst22155 (P3_ADD_541_U21, P3_INSTADDRPOINTER_REG_10__SCAN_IN);
  nand ginst22156 (P3_ADD_541_U22, P3_INSTADDRPOINTER_REG_10__SCAN_IN, P3_ADD_541_U101);
  not ginst22157 (P3_ADD_541_U23, P3_INSTADDRPOINTER_REG_11__SCAN_IN);
  nand ginst22158 (P3_ADD_541_U24, P3_INSTADDRPOINTER_REG_11__SCAN_IN, P3_ADD_541_U102);
  not ginst22159 (P3_ADD_541_U25, P3_INSTADDRPOINTER_REG_12__SCAN_IN);
  nand ginst22160 (P3_ADD_541_U26, P3_INSTADDRPOINTER_REG_12__SCAN_IN, P3_ADD_541_U103);
  not ginst22161 (P3_ADD_541_U27, P3_INSTADDRPOINTER_REG_13__SCAN_IN);
  nand ginst22162 (P3_ADD_541_U28, P3_INSTADDRPOINTER_REG_13__SCAN_IN, P3_ADD_541_U104);
  not ginst22163 (P3_ADD_541_U29, P3_INSTADDRPOINTER_REG_14__SCAN_IN);
  nand ginst22164 (P3_ADD_541_U30, P3_INSTADDRPOINTER_REG_14__SCAN_IN, P3_ADD_541_U105);
  not ginst22165 (P3_ADD_541_U31, P3_INSTADDRPOINTER_REG_15__SCAN_IN);
  nand ginst22166 (P3_ADD_541_U32, P3_INSTADDRPOINTER_REG_15__SCAN_IN, P3_ADD_541_U106);
  not ginst22167 (P3_ADD_541_U33, P3_INSTADDRPOINTER_REG_16__SCAN_IN);
  nand ginst22168 (P3_ADD_541_U34, P3_INSTADDRPOINTER_REG_16__SCAN_IN, P3_ADD_541_U107);
  not ginst22169 (P3_ADD_541_U35, P3_INSTADDRPOINTER_REG_17__SCAN_IN);
  nand ginst22170 (P3_ADD_541_U36, P3_INSTADDRPOINTER_REG_17__SCAN_IN, P3_ADD_541_U108);
  not ginst22171 (P3_ADD_541_U37, P3_INSTADDRPOINTER_REG_18__SCAN_IN);
  nand ginst22172 (P3_ADD_541_U38, P3_INSTADDRPOINTER_REG_18__SCAN_IN, P3_ADD_541_U109);
  not ginst22173 (P3_ADD_541_U39, P3_INSTADDRPOINTER_REG_19__SCAN_IN);
  not ginst22174 (P3_ADD_541_U4, P3_INSTADDRPOINTER_REG_1__SCAN_IN);
  nand ginst22175 (P3_ADD_541_U40, P3_INSTADDRPOINTER_REG_19__SCAN_IN, P3_ADD_541_U110);
  not ginst22176 (P3_ADD_541_U41, P3_INSTADDRPOINTER_REG_20__SCAN_IN);
  nand ginst22177 (P3_ADD_541_U42, P3_INSTADDRPOINTER_REG_20__SCAN_IN, P3_ADD_541_U111);
  not ginst22178 (P3_ADD_541_U43, P3_INSTADDRPOINTER_REG_21__SCAN_IN);
  nand ginst22179 (P3_ADD_541_U44, P3_INSTADDRPOINTER_REG_21__SCAN_IN, P3_ADD_541_U112);
  not ginst22180 (P3_ADD_541_U45, P3_INSTADDRPOINTER_REG_22__SCAN_IN);
  nand ginst22181 (P3_ADD_541_U46, P3_INSTADDRPOINTER_REG_22__SCAN_IN, P3_ADD_541_U113);
  not ginst22182 (P3_ADD_541_U47, P3_INSTADDRPOINTER_REG_23__SCAN_IN);
  nand ginst22183 (P3_ADD_541_U48, P3_INSTADDRPOINTER_REG_23__SCAN_IN, P3_ADD_541_U114);
  not ginst22184 (P3_ADD_541_U49, P3_INSTADDRPOINTER_REG_24__SCAN_IN);
  not ginst22185 (P3_ADD_541_U5, P3_INSTADDRPOINTER_REG_2__SCAN_IN);
  nand ginst22186 (P3_ADD_541_U50, P3_INSTADDRPOINTER_REG_24__SCAN_IN, P3_ADD_541_U115);
  not ginst22187 (P3_ADD_541_U51, P3_INSTADDRPOINTER_REG_25__SCAN_IN);
  nand ginst22188 (P3_ADD_541_U52, P3_INSTADDRPOINTER_REG_25__SCAN_IN, P3_ADD_541_U116);
  not ginst22189 (P3_ADD_541_U53, P3_INSTADDRPOINTER_REG_26__SCAN_IN);
  nand ginst22190 (P3_ADD_541_U54, P3_INSTADDRPOINTER_REG_26__SCAN_IN, P3_ADD_541_U117);
  not ginst22191 (P3_ADD_541_U55, P3_INSTADDRPOINTER_REG_27__SCAN_IN);
  nand ginst22192 (P3_ADD_541_U56, P3_INSTADDRPOINTER_REG_27__SCAN_IN, P3_ADD_541_U118);
  not ginst22193 (P3_ADD_541_U57, P3_INSTADDRPOINTER_REG_28__SCAN_IN);
  nand ginst22194 (P3_ADD_541_U58, P3_INSTADDRPOINTER_REG_28__SCAN_IN, P3_ADD_541_U119);
  not ginst22195 (P3_ADD_541_U59, P3_INSTADDRPOINTER_REG_29__SCAN_IN);
  nand ginst22196 (P3_ADD_541_U6, P3_INSTADDRPOINTER_REG_1__SCAN_IN, P3_INSTADDRPOINTER_REG_2__SCAN_IN);
  nand ginst22197 (P3_ADD_541_U60, P3_INSTADDRPOINTER_REG_29__SCAN_IN, P3_ADD_541_U120);
  not ginst22198 (P3_ADD_541_U61, P3_INSTADDRPOINTER_REG_30__SCAN_IN);
  nand ginst22199 (P3_ADD_541_U62, P3_ADD_541_U123, P3_ADD_541_U124);
  nand ginst22200 (P3_ADD_541_U63, P3_ADD_541_U125, P3_ADD_541_U126);
  nand ginst22201 (P3_ADD_541_U64, P3_ADD_541_U127, P3_ADD_541_U128);
  nand ginst22202 (P3_ADD_541_U65, P3_ADD_541_U129, P3_ADD_541_U130);
  nand ginst22203 (P3_ADD_541_U66, P3_ADD_541_U131, P3_ADD_541_U132);
  nand ginst22204 (P3_ADD_541_U67, P3_ADD_541_U133, P3_ADD_541_U134);
  nand ginst22205 (P3_ADD_541_U68, P3_ADD_541_U135, P3_ADD_541_U136);
  nand ginst22206 (P3_ADD_541_U69, P3_ADD_541_U137, P3_ADD_541_U138);
  not ginst22207 (P3_ADD_541_U7, P3_INSTADDRPOINTER_REG_3__SCAN_IN);
  nand ginst22208 (P3_ADD_541_U70, P3_ADD_541_U139, P3_ADD_541_U140);
  nand ginst22209 (P3_ADD_541_U71, P3_ADD_541_U141, P3_ADD_541_U142);
  nand ginst22210 (P3_ADD_541_U72, P3_ADD_541_U143, P3_ADD_541_U144);
  nand ginst22211 (P3_ADD_541_U73, P3_ADD_541_U145, P3_ADD_541_U146);
  nand ginst22212 (P3_ADD_541_U74, P3_ADD_541_U147, P3_ADD_541_U148);
  nand ginst22213 (P3_ADD_541_U75, P3_ADD_541_U149, P3_ADD_541_U150);
  nand ginst22214 (P3_ADD_541_U76, P3_ADD_541_U151, P3_ADD_541_U152);
  nand ginst22215 (P3_ADD_541_U77, P3_ADD_541_U153, P3_ADD_541_U154);
  nand ginst22216 (P3_ADD_541_U78, P3_ADD_541_U155, P3_ADD_541_U156);
  nand ginst22217 (P3_ADD_541_U79, P3_ADD_541_U157, P3_ADD_541_U158);
  nand ginst22218 (P3_ADD_541_U8, P3_INSTADDRPOINTER_REG_3__SCAN_IN, P3_ADD_541_U94);
  nand ginst22219 (P3_ADD_541_U80, P3_ADD_541_U159, P3_ADD_541_U160);
  nand ginst22220 (P3_ADD_541_U81, P3_ADD_541_U161, P3_ADD_541_U162);
  nand ginst22221 (P3_ADD_541_U82, P3_ADD_541_U163, P3_ADD_541_U164);
  nand ginst22222 (P3_ADD_541_U83, P3_ADD_541_U165, P3_ADD_541_U166);
  nand ginst22223 (P3_ADD_541_U84, P3_ADD_541_U167, P3_ADD_541_U168);
  nand ginst22224 (P3_ADD_541_U85, P3_ADD_541_U169, P3_ADD_541_U170);
  nand ginst22225 (P3_ADD_541_U86, P3_ADD_541_U171, P3_ADD_541_U172);
  nand ginst22226 (P3_ADD_541_U87, P3_ADD_541_U173, P3_ADD_541_U174);
  nand ginst22227 (P3_ADD_541_U88, P3_ADD_541_U175, P3_ADD_541_U176);
  nand ginst22228 (P3_ADD_541_U89, P3_ADD_541_U177, P3_ADD_541_U178);
  not ginst22229 (P3_ADD_541_U9, P3_INSTADDRPOINTER_REG_4__SCAN_IN);
  nand ginst22230 (P3_ADD_541_U90, P3_ADD_541_U179, P3_ADD_541_U180);
  nand ginst22231 (P3_ADD_541_U91, P3_ADD_541_U181, P3_ADD_541_U182);
  not ginst22232 (P3_ADD_541_U92, P3_INSTADDRPOINTER_REG_31__SCAN_IN);
  nand ginst22233 (P3_ADD_541_U93, P3_INSTADDRPOINTER_REG_30__SCAN_IN, P3_ADD_541_U121);
  not ginst22234 (P3_ADD_541_U94, P3_ADD_541_U6);
  not ginst22235 (P3_ADD_541_U95, P3_ADD_541_U8);
  not ginst22236 (P3_ADD_541_U96, P3_ADD_541_U10);
  not ginst22237 (P3_ADD_541_U97, P3_ADD_541_U12);
  not ginst22238 (P3_ADD_541_U98, P3_ADD_541_U14);
  not ginst22239 (P3_ADD_541_U99, P3_ADD_541_U16);
  nand ginst22240 (P3_ADD_546_U10, P3_EAX_REG_0__SCAN_IN, P3_EAX_REG_1__SCAN_IN, P3_EAX_REG_2__SCAN_IN);
  nand ginst22241 (P3_ADD_546_U100, P3_EAX_REG_0__SCAN_IN, P3_EAX_REG_1__SCAN_IN);
  nand ginst22242 (P3_ADD_546_U101, P3_EAX_REG_27__SCAN_IN, P3_ADD_546_U122);
  nand ginst22243 (P3_ADD_546_U102, P3_EAX_REG_25__SCAN_IN, P3_ADD_546_U116);
  nand ginst22244 (P3_ADD_546_U103, P3_EAX_REG_23__SCAN_IN, P3_ADD_546_U115);
  nand ginst22245 (P3_ADD_546_U104, P3_EAX_REG_21__SCAN_IN, P3_ADD_546_U121);
  nand ginst22246 (P3_ADD_546_U105, P3_EAX_REG_19__SCAN_IN, P3_ADD_546_U114);
  nand ginst22247 (P3_ADD_546_U106, P3_EAX_REG_17__SCAN_IN, P3_ADD_546_U117);
  nand ginst22248 (P3_ADD_546_U107, P3_EAX_REG_15__SCAN_IN, P3_ADD_546_U124);
  nand ginst22249 (P3_ADD_546_U108, P3_EAX_REG_13__SCAN_IN, P3_ADD_546_U119);
  nand ginst22250 (P3_ADD_546_U109, P3_EAX_REG_11__SCAN_IN, P3_ADD_546_U113);
  not ginst22251 (P3_ADD_546_U11, P3_EAX_REG_6__SCAN_IN);
  nand ginst22252 (P3_ADD_546_U110, P3_EAX_REG_9__SCAN_IN, P3_ADD_546_U120);
  not ginst22253 (P3_ADD_546_U111, P3_ADD_546_U10);
  not ginst22254 (P3_ADD_546_U112, P3_ADD_546_U13);
  not ginst22255 (P3_ADD_546_U113, P3_ADD_546_U22);
  not ginst22256 (P3_ADD_546_U114, P3_ADD_546_U34);
  not ginst22257 (P3_ADD_546_U115, P3_ADD_546_U40);
  not ginst22258 (P3_ADD_546_U116, P3_ADD_546_U43);
  not ginst22259 (P3_ADD_546_U117, P3_ADD_546_U31);
  not ginst22260 (P3_ADD_546_U118, P3_ADD_546_U16);
  not ginst22261 (P3_ADD_546_U119, P3_ADD_546_U25);
  not ginst22262 (P3_ADD_546_U12, P3_EAX_REG_5__SCAN_IN);
  not ginst22263 (P3_ADD_546_U120, P3_ADD_546_U17);
  not ginst22264 (P3_ADD_546_U121, P3_ADD_546_U36);
  not ginst22265 (P3_ADD_546_U122, P3_ADD_546_U46);
  not ginst22266 (P3_ADD_546_U123, P3_ADD_546_U48);
  not ginst22267 (P3_ADD_546_U124, P3_ADD_546_U27);
  not ginst22268 (P3_ADD_546_U125, P3_ADD_546_U95);
  not ginst22269 (P3_ADD_546_U126, P3_ADD_546_U96);
  not ginst22270 (P3_ADD_546_U127, P3_ADD_546_U97);
  not ginst22271 (P3_ADD_546_U128, P3_ADD_546_U49);
  not ginst22272 (P3_ADD_546_U129, P3_ADD_546_U99);
  nand ginst22273 (P3_ADD_546_U13, P3_ADD_546_U111, P3_ADD_546_U82);
  not ginst22274 (P3_ADD_546_U130, P3_ADD_546_U100);
  not ginst22275 (P3_ADD_546_U131, P3_ADD_546_U101);
  not ginst22276 (P3_ADD_546_U132, P3_ADD_546_U102);
  not ginst22277 (P3_ADD_546_U133, P3_ADD_546_U103);
  not ginst22278 (P3_ADD_546_U134, P3_ADD_546_U104);
  not ginst22279 (P3_ADD_546_U135, P3_ADD_546_U105);
  not ginst22280 (P3_ADD_546_U136, P3_ADD_546_U106);
  not ginst22281 (P3_ADD_546_U137, P3_ADD_546_U107);
  not ginst22282 (P3_ADD_546_U138, P3_ADD_546_U108);
  not ginst22283 (P3_ADD_546_U139, P3_ADD_546_U109);
  not ginst22284 (P3_ADD_546_U14, P3_EAX_REG_8__SCAN_IN);
  not ginst22285 (P3_ADD_546_U140, P3_ADD_546_U110);
  nand ginst22286 (P3_ADD_546_U141, P3_ADD_546_U120, P3_ADD_546_U18);
  nand ginst22287 (P3_ADD_546_U142, P3_EAX_REG_9__SCAN_IN, P3_ADD_546_U17);
  nand ginst22288 (P3_ADD_546_U143, P3_EAX_REG_8__SCAN_IN, P3_ADD_546_U95);
  nand ginst22289 (P3_ADD_546_U144, P3_ADD_546_U125, P3_ADD_546_U14);
  nand ginst22290 (P3_ADD_546_U145, P3_ADD_546_U118, P3_ADD_546_U15);
  nand ginst22291 (P3_ADD_546_U146, P3_EAX_REG_7__SCAN_IN, P3_ADD_546_U16);
  nand ginst22292 (P3_ADD_546_U147, P3_EAX_REG_6__SCAN_IN, P3_ADD_546_U96);
  nand ginst22293 (P3_ADD_546_U148, P3_ADD_546_U11, P3_ADD_546_U126);
  nand ginst22294 (P3_ADD_546_U149, P3_ADD_546_U112, P3_ADD_546_U12);
  not ginst22295 (P3_ADD_546_U15, P3_EAX_REG_7__SCAN_IN);
  nand ginst22296 (P3_ADD_546_U150, P3_EAX_REG_5__SCAN_IN, P3_ADD_546_U13);
  nand ginst22297 (P3_ADD_546_U151, P3_EAX_REG_4__SCAN_IN, P3_ADD_546_U97);
  nand ginst22298 (P3_ADD_546_U152, P3_ADD_546_U127, P3_ADD_546_U8);
  nand ginst22299 (P3_ADD_546_U153, P3_ADD_546_U111, P3_ADD_546_U9);
  nand ginst22300 (P3_ADD_546_U154, P3_EAX_REG_3__SCAN_IN, P3_ADD_546_U10);
  nand ginst22301 (P3_ADD_546_U155, P3_EAX_REG_31__SCAN_IN, P3_ADD_546_U99);
  nand ginst22302 (P3_ADD_546_U156, P3_ADD_546_U129, P3_ADD_546_U98);
  nand ginst22303 (P3_ADD_546_U157, P3_EAX_REG_30__SCAN_IN, P3_ADD_546_U49);
  nand ginst22304 (P3_ADD_546_U158, P3_ADD_546_U128, P3_ADD_546_U50);
  nand ginst22305 (P3_ADD_546_U159, P3_EAX_REG_2__SCAN_IN, P3_ADD_546_U100);
  nand ginst22306 (P3_ADD_546_U16, P3_ADD_546_U112, P3_ADD_546_U83);
  nand ginst22307 (P3_ADD_546_U160, P3_ADD_546_U130, P3_ADD_546_U6);
  nand ginst22308 (P3_ADD_546_U161, P3_ADD_546_U123, P3_ADD_546_U47);
  nand ginst22309 (P3_ADD_546_U162, P3_EAX_REG_29__SCAN_IN, P3_ADD_546_U48);
  nand ginst22310 (P3_ADD_546_U163, P3_EAX_REG_28__SCAN_IN, P3_ADD_546_U101);
  nand ginst22311 (P3_ADD_546_U164, P3_ADD_546_U131, P3_ADD_546_U45);
  nand ginst22312 (P3_ADD_546_U165, P3_ADD_546_U122, P3_ADD_546_U44);
  nand ginst22313 (P3_ADD_546_U166, P3_EAX_REG_27__SCAN_IN, P3_ADD_546_U46);
  nand ginst22314 (P3_ADD_546_U167, P3_EAX_REG_26__SCAN_IN, P3_ADD_546_U102);
  nand ginst22315 (P3_ADD_546_U168, P3_ADD_546_U132, P3_ADD_546_U41);
  nand ginst22316 (P3_ADD_546_U169, P3_ADD_546_U116, P3_ADD_546_U42);
  nand ginst22317 (P3_ADD_546_U17, P3_ADD_546_U118, P3_ADD_546_U84);
  nand ginst22318 (P3_ADD_546_U170, P3_EAX_REG_25__SCAN_IN, P3_ADD_546_U43);
  nand ginst22319 (P3_ADD_546_U171, P3_EAX_REG_24__SCAN_IN, P3_ADD_546_U103);
  nand ginst22320 (P3_ADD_546_U172, P3_ADD_546_U133, P3_ADD_546_U38);
  nand ginst22321 (P3_ADD_546_U173, P3_ADD_546_U115, P3_ADD_546_U39);
  nand ginst22322 (P3_ADD_546_U174, P3_EAX_REG_23__SCAN_IN, P3_ADD_546_U40);
  nand ginst22323 (P3_ADD_546_U175, P3_EAX_REG_22__SCAN_IN, P3_ADD_546_U104);
  nand ginst22324 (P3_ADD_546_U176, P3_ADD_546_U134, P3_ADD_546_U37);
  nand ginst22325 (P3_ADD_546_U177, P3_ADD_546_U121, P3_ADD_546_U35);
  nand ginst22326 (P3_ADD_546_U178, P3_EAX_REG_21__SCAN_IN, P3_ADD_546_U36);
  nand ginst22327 (P3_ADD_546_U179, P3_EAX_REG_20__SCAN_IN, P3_ADD_546_U105);
  not ginst22328 (P3_ADD_546_U18, P3_EAX_REG_9__SCAN_IN);
  nand ginst22329 (P3_ADD_546_U180, P3_ADD_546_U135, P3_ADD_546_U32);
  nand ginst22330 (P3_ADD_546_U181, P3_EAX_REG_0__SCAN_IN, P3_ADD_546_U7);
  nand ginst22331 (P3_ADD_546_U182, P3_EAX_REG_1__SCAN_IN, P3_ADD_546_U5);
  nand ginst22332 (P3_ADD_546_U183, P3_ADD_546_U114, P3_ADD_546_U33);
  nand ginst22333 (P3_ADD_546_U184, P3_EAX_REG_19__SCAN_IN, P3_ADD_546_U34);
  nand ginst22334 (P3_ADD_546_U185, P3_EAX_REG_18__SCAN_IN, P3_ADD_546_U106);
  nand ginst22335 (P3_ADD_546_U186, P3_ADD_546_U136, P3_ADD_546_U29);
  nand ginst22336 (P3_ADD_546_U187, P3_ADD_546_U117, P3_ADD_546_U30);
  nand ginst22337 (P3_ADD_546_U188, P3_EAX_REG_17__SCAN_IN, P3_ADD_546_U31);
  nand ginst22338 (P3_ADD_546_U189, P3_EAX_REG_16__SCAN_IN, P3_ADD_546_U107);
  not ginst22339 (P3_ADD_546_U19, P3_EAX_REG_10__SCAN_IN);
  nand ginst22340 (P3_ADD_546_U190, P3_ADD_546_U137, P3_ADD_546_U28);
  nand ginst22341 (P3_ADD_546_U191, P3_ADD_546_U124, P3_ADD_546_U26);
  nand ginst22342 (P3_ADD_546_U192, P3_EAX_REG_15__SCAN_IN, P3_ADD_546_U27);
  nand ginst22343 (P3_ADD_546_U193, P3_EAX_REG_14__SCAN_IN, P3_ADD_546_U108);
  nand ginst22344 (P3_ADD_546_U194, P3_ADD_546_U138, P3_ADD_546_U23);
  nand ginst22345 (P3_ADD_546_U195, P3_ADD_546_U119, P3_ADD_546_U24);
  nand ginst22346 (P3_ADD_546_U196, P3_EAX_REG_13__SCAN_IN, P3_ADD_546_U25);
  nand ginst22347 (P3_ADD_546_U197, P3_EAX_REG_12__SCAN_IN, P3_ADD_546_U109);
  nand ginst22348 (P3_ADD_546_U198, P3_ADD_546_U139, P3_ADD_546_U20);
  nand ginst22349 (P3_ADD_546_U199, P3_ADD_546_U113, P3_ADD_546_U21);
  not ginst22350 (P3_ADD_546_U20, P3_EAX_REG_12__SCAN_IN);
  nand ginst22351 (P3_ADD_546_U200, P3_EAX_REG_11__SCAN_IN, P3_ADD_546_U22);
  nand ginst22352 (P3_ADD_546_U201, P3_EAX_REG_10__SCAN_IN, P3_ADD_546_U110);
  nand ginst22353 (P3_ADD_546_U202, P3_ADD_546_U140, P3_ADD_546_U19);
  not ginst22354 (P3_ADD_546_U21, P3_EAX_REG_11__SCAN_IN);
  nand ginst22355 (P3_ADD_546_U22, P3_ADD_546_U120, P3_ADD_546_U85);
  not ginst22356 (P3_ADD_546_U23, P3_EAX_REG_14__SCAN_IN);
  not ginst22357 (P3_ADD_546_U24, P3_EAX_REG_13__SCAN_IN);
  nand ginst22358 (P3_ADD_546_U25, P3_ADD_546_U113, P3_ADD_546_U86);
  not ginst22359 (P3_ADD_546_U26, P3_EAX_REG_15__SCAN_IN);
  nand ginst22360 (P3_ADD_546_U27, P3_ADD_546_U119, P3_ADD_546_U87);
  not ginst22361 (P3_ADD_546_U28, P3_EAX_REG_16__SCAN_IN);
  not ginst22362 (P3_ADD_546_U29, P3_EAX_REG_18__SCAN_IN);
  not ginst22363 (P3_ADD_546_U30, P3_EAX_REG_17__SCAN_IN);
  nand ginst22364 (P3_ADD_546_U31, P3_ADD_546_U124, P3_ADD_546_U88);
  not ginst22365 (P3_ADD_546_U32, P3_EAX_REG_20__SCAN_IN);
  not ginst22366 (P3_ADD_546_U33, P3_EAX_REG_19__SCAN_IN);
  nand ginst22367 (P3_ADD_546_U34, P3_ADD_546_U117, P3_ADD_546_U89);
  not ginst22368 (P3_ADD_546_U35, P3_EAX_REG_21__SCAN_IN);
  nand ginst22369 (P3_ADD_546_U36, P3_ADD_546_U114, P3_ADD_546_U90);
  not ginst22370 (P3_ADD_546_U37, P3_EAX_REG_22__SCAN_IN);
  not ginst22371 (P3_ADD_546_U38, P3_EAX_REG_24__SCAN_IN);
  not ginst22372 (P3_ADD_546_U39, P3_EAX_REG_23__SCAN_IN);
  nand ginst22373 (P3_ADD_546_U40, P3_ADD_546_U121, P3_ADD_546_U91);
  not ginst22374 (P3_ADD_546_U41, P3_EAX_REG_26__SCAN_IN);
  not ginst22375 (P3_ADD_546_U42, P3_EAX_REG_25__SCAN_IN);
  nand ginst22376 (P3_ADD_546_U43, P3_ADD_546_U115, P3_ADD_546_U92);
  not ginst22377 (P3_ADD_546_U44, P3_EAX_REG_27__SCAN_IN);
  not ginst22378 (P3_ADD_546_U45, P3_EAX_REG_28__SCAN_IN);
  nand ginst22379 (P3_ADD_546_U46, P3_ADD_546_U116, P3_ADD_546_U93);
  not ginst22380 (P3_ADD_546_U47, P3_EAX_REG_29__SCAN_IN);
  nand ginst22381 (P3_ADD_546_U48, P3_ADD_546_U122, P3_ADD_546_U94);
  nand ginst22382 (P3_ADD_546_U49, P3_EAX_REG_29__SCAN_IN, P3_ADD_546_U123);
  not ginst22383 (P3_ADD_546_U5, P3_EAX_REG_0__SCAN_IN);
  not ginst22384 (P3_ADD_546_U50, P3_EAX_REG_30__SCAN_IN);
  nand ginst22385 (P3_ADD_546_U51, P3_ADD_546_U141, P3_ADD_546_U142);
  nand ginst22386 (P3_ADD_546_U52, P3_ADD_546_U143, P3_ADD_546_U144);
  nand ginst22387 (P3_ADD_546_U53, P3_ADD_546_U145, P3_ADD_546_U146);
  nand ginst22388 (P3_ADD_546_U54, P3_ADD_546_U147, P3_ADD_546_U148);
  nand ginst22389 (P3_ADD_546_U55, P3_ADD_546_U149, P3_ADD_546_U150);
  nand ginst22390 (P3_ADD_546_U56, P3_ADD_546_U151, P3_ADD_546_U152);
  nand ginst22391 (P3_ADD_546_U57, P3_ADD_546_U153, P3_ADD_546_U154);
  nand ginst22392 (P3_ADD_546_U58, P3_ADD_546_U155, P3_ADD_546_U156);
  nand ginst22393 (P3_ADD_546_U59, P3_ADD_546_U157, P3_ADD_546_U158);
  not ginst22394 (P3_ADD_546_U6, P3_EAX_REG_2__SCAN_IN);
  nand ginst22395 (P3_ADD_546_U60, P3_ADD_546_U159, P3_ADD_546_U160);
  nand ginst22396 (P3_ADD_546_U61, P3_ADD_546_U161, P3_ADD_546_U162);
  nand ginst22397 (P3_ADD_546_U62, P3_ADD_546_U163, P3_ADD_546_U164);
  nand ginst22398 (P3_ADD_546_U63, P3_ADD_546_U165, P3_ADD_546_U166);
  nand ginst22399 (P3_ADD_546_U64, P3_ADD_546_U167, P3_ADD_546_U168);
  nand ginst22400 (P3_ADD_546_U65, P3_ADD_546_U169, P3_ADD_546_U170);
  nand ginst22401 (P3_ADD_546_U66, P3_ADD_546_U171, P3_ADD_546_U172);
  nand ginst22402 (P3_ADD_546_U67, P3_ADD_546_U173, P3_ADD_546_U174);
  nand ginst22403 (P3_ADD_546_U68, P3_ADD_546_U175, P3_ADD_546_U176);
  nand ginst22404 (P3_ADD_546_U69, P3_ADD_546_U177, P3_ADD_546_U178);
  not ginst22405 (P3_ADD_546_U7, P3_EAX_REG_1__SCAN_IN);
  nand ginst22406 (P3_ADD_546_U70, P3_ADD_546_U179, P3_ADD_546_U180);
  nand ginst22407 (P3_ADD_546_U71, P3_ADD_546_U181, P3_ADD_546_U182);
  nand ginst22408 (P3_ADD_546_U72, P3_ADD_546_U183, P3_ADD_546_U184);
  nand ginst22409 (P3_ADD_546_U73, P3_ADD_546_U185, P3_ADD_546_U186);
  nand ginst22410 (P3_ADD_546_U74, P3_ADD_546_U187, P3_ADD_546_U188);
  nand ginst22411 (P3_ADD_546_U75, P3_ADD_546_U189, P3_ADD_546_U190);
  nand ginst22412 (P3_ADD_546_U76, P3_ADD_546_U191, P3_ADD_546_U192);
  nand ginst22413 (P3_ADD_546_U77, P3_ADD_546_U193, P3_ADD_546_U194);
  nand ginst22414 (P3_ADD_546_U78, P3_ADD_546_U195, P3_ADD_546_U196);
  nand ginst22415 (P3_ADD_546_U79, P3_ADD_546_U197, P3_ADD_546_U198);
  not ginst22416 (P3_ADD_546_U8, P3_EAX_REG_4__SCAN_IN);
  nand ginst22417 (P3_ADD_546_U80, P3_ADD_546_U199, P3_ADD_546_U200);
  nand ginst22418 (P3_ADD_546_U81, P3_ADD_546_U201, P3_ADD_546_U202);
  and ginst22419 (P3_ADD_546_U82, P3_EAX_REG_3__SCAN_IN, P3_EAX_REG_4__SCAN_IN);
  and ginst22420 (P3_ADD_546_U83, P3_EAX_REG_5__SCAN_IN, P3_EAX_REG_6__SCAN_IN);
  and ginst22421 (P3_ADD_546_U84, P3_EAX_REG_7__SCAN_IN, P3_EAX_REG_8__SCAN_IN);
  and ginst22422 (P3_ADD_546_U85, P3_EAX_REG_9__SCAN_IN, P3_EAX_REG_10__SCAN_IN);
  and ginst22423 (P3_ADD_546_U86, P3_EAX_REG_11__SCAN_IN, P3_EAX_REG_12__SCAN_IN);
  and ginst22424 (P3_ADD_546_U87, P3_EAX_REG_13__SCAN_IN, P3_EAX_REG_14__SCAN_IN);
  and ginst22425 (P3_ADD_546_U88, P3_EAX_REG_15__SCAN_IN, P3_EAX_REG_16__SCAN_IN);
  and ginst22426 (P3_ADD_546_U89, P3_EAX_REG_17__SCAN_IN, P3_EAX_REG_18__SCAN_IN);
  not ginst22427 (P3_ADD_546_U9, P3_EAX_REG_3__SCAN_IN);
  and ginst22428 (P3_ADD_546_U90, P3_EAX_REG_19__SCAN_IN, P3_EAX_REG_20__SCAN_IN);
  and ginst22429 (P3_ADD_546_U91, P3_EAX_REG_21__SCAN_IN, P3_EAX_REG_22__SCAN_IN);
  and ginst22430 (P3_ADD_546_U92, P3_EAX_REG_23__SCAN_IN, P3_EAX_REG_24__SCAN_IN);
  and ginst22431 (P3_ADD_546_U93, P3_EAX_REG_25__SCAN_IN, P3_EAX_REG_26__SCAN_IN);
  and ginst22432 (P3_ADD_546_U94, P3_EAX_REG_27__SCAN_IN, P3_EAX_REG_28__SCAN_IN);
  nand ginst22433 (P3_ADD_546_U95, P3_EAX_REG_7__SCAN_IN, P3_ADD_546_U118);
  nand ginst22434 (P3_ADD_546_U96, P3_EAX_REG_5__SCAN_IN, P3_ADD_546_U112);
  nand ginst22435 (P3_ADD_546_U97, P3_EAX_REG_3__SCAN_IN, P3_ADD_546_U111);
  not ginst22436 (P3_ADD_546_U98, P3_EAX_REG_31__SCAN_IN);
  nand ginst22437 (P3_ADD_546_U99, P3_EAX_REG_30__SCAN_IN, P3_ADD_546_U128);
  not ginst22438 (P3_ADD_547_U10, P3_INSTADDRPOINTER_REG_3__SCAN_IN);
  not ginst22439 (P3_ADD_547_U100, P3_ADD_547_U11);
  not ginst22440 (P3_ADD_547_U101, P3_ADD_547_U13);
  not ginst22441 (P3_ADD_547_U102, P3_ADD_547_U15);
  not ginst22442 (P3_ADD_547_U103, P3_ADD_547_U17);
  not ginst22443 (P3_ADD_547_U104, P3_ADD_547_U19);
  not ginst22444 (P3_ADD_547_U105, P3_ADD_547_U22);
  not ginst22445 (P3_ADD_547_U106, P3_ADD_547_U23);
  not ginst22446 (P3_ADD_547_U107, P3_ADD_547_U25);
  not ginst22447 (P3_ADD_547_U108, P3_ADD_547_U27);
  not ginst22448 (P3_ADD_547_U109, P3_ADD_547_U29);
  nand ginst22449 (P3_ADD_547_U11, P3_INSTADDRPOINTER_REG_3__SCAN_IN, P3_ADD_547_U99);
  not ginst22450 (P3_ADD_547_U110, P3_ADD_547_U31);
  not ginst22451 (P3_ADD_547_U111, P3_ADD_547_U33);
  not ginst22452 (P3_ADD_547_U112, P3_ADD_547_U35);
  not ginst22453 (P3_ADD_547_U113, P3_ADD_547_U37);
  not ginst22454 (P3_ADD_547_U114, P3_ADD_547_U39);
  not ginst22455 (P3_ADD_547_U115, P3_ADD_547_U41);
  not ginst22456 (P3_ADD_547_U116, P3_ADD_547_U43);
  not ginst22457 (P3_ADD_547_U117, P3_ADD_547_U45);
  not ginst22458 (P3_ADD_547_U118, P3_ADD_547_U47);
  not ginst22459 (P3_ADD_547_U119, P3_ADD_547_U49);
  not ginst22460 (P3_ADD_547_U12, P3_INSTADDRPOINTER_REG_4__SCAN_IN);
  not ginst22461 (P3_ADD_547_U120, P3_ADD_547_U51);
  not ginst22462 (P3_ADD_547_U121, P3_ADD_547_U53);
  not ginst22463 (P3_ADD_547_U122, P3_ADD_547_U55);
  not ginst22464 (P3_ADD_547_U123, P3_ADD_547_U57);
  not ginst22465 (P3_ADD_547_U124, P3_ADD_547_U59);
  not ginst22466 (P3_ADD_547_U125, P3_ADD_547_U61);
  not ginst22467 (P3_ADD_547_U126, P3_ADD_547_U63);
  not ginst22468 (P3_ADD_547_U127, P3_ADD_547_U97);
  nand ginst22469 (P3_ADD_547_U128, P3_INSTADDRPOINTER_REG_9__SCAN_IN, P3_ADD_547_U22);
  nand ginst22470 (P3_ADD_547_U129, P3_ADD_547_U105, P3_ADD_547_U21);
  nand ginst22471 (P3_ADD_547_U13, P3_INSTADDRPOINTER_REG_4__SCAN_IN, P3_ADD_547_U100);
  nand ginst22472 (P3_ADD_547_U130, P3_INSTADDRPOINTER_REG_8__SCAN_IN, P3_ADD_547_U19);
  nand ginst22473 (P3_ADD_547_U131, P3_ADD_547_U104, P3_ADD_547_U20);
  nand ginst22474 (P3_ADD_547_U132, P3_INSTADDRPOINTER_REG_7__SCAN_IN, P3_ADD_547_U17);
  nand ginst22475 (P3_ADD_547_U133, P3_ADD_547_U103, P3_ADD_547_U18);
  nand ginst22476 (P3_ADD_547_U134, P3_INSTADDRPOINTER_REG_6__SCAN_IN, P3_ADD_547_U15);
  nand ginst22477 (P3_ADD_547_U135, P3_ADD_547_U102, P3_ADD_547_U16);
  nand ginst22478 (P3_ADD_547_U136, P3_INSTADDRPOINTER_REG_5__SCAN_IN, P3_ADD_547_U13);
  nand ginst22479 (P3_ADD_547_U137, P3_ADD_547_U101, P3_ADD_547_U14);
  nand ginst22480 (P3_ADD_547_U138, P3_INSTADDRPOINTER_REG_4__SCAN_IN, P3_ADD_547_U11);
  nand ginst22481 (P3_ADD_547_U139, P3_ADD_547_U100, P3_ADD_547_U12);
  not ginst22482 (P3_ADD_547_U14, P3_INSTADDRPOINTER_REG_5__SCAN_IN);
  nand ginst22483 (P3_ADD_547_U140, P3_INSTADDRPOINTER_REG_3__SCAN_IN, P3_ADD_547_U9);
  nand ginst22484 (P3_ADD_547_U141, P3_ADD_547_U10, P3_ADD_547_U99);
  nand ginst22485 (P3_ADD_547_U142, P3_INSTADDRPOINTER_REG_31__SCAN_IN, P3_ADD_547_U97);
  nand ginst22486 (P3_ADD_547_U143, P3_ADD_547_U127, P3_ADD_547_U96);
  nand ginst22487 (P3_ADD_547_U144, P3_INSTADDRPOINTER_REG_30__SCAN_IN, P3_ADD_547_U63);
  nand ginst22488 (P3_ADD_547_U145, P3_ADD_547_U126, P3_ADD_547_U64);
  nand ginst22489 (P3_ADD_547_U146, P3_INSTADDRPOINTER_REG_2__SCAN_IN, P3_ADD_547_U7);
  nand ginst22490 (P3_ADD_547_U147, P3_ADD_547_U8, P3_ADD_547_U98);
  nand ginst22491 (P3_ADD_547_U148, P3_INSTADDRPOINTER_REG_29__SCAN_IN, P3_ADD_547_U61);
  nand ginst22492 (P3_ADD_547_U149, P3_ADD_547_U125, P3_ADD_547_U62);
  nand ginst22493 (P3_ADD_547_U15, P3_INSTADDRPOINTER_REG_5__SCAN_IN, P3_ADD_547_U101);
  nand ginst22494 (P3_ADD_547_U150, P3_INSTADDRPOINTER_REG_28__SCAN_IN, P3_ADD_547_U59);
  nand ginst22495 (P3_ADD_547_U151, P3_ADD_547_U124, P3_ADD_547_U60);
  nand ginst22496 (P3_ADD_547_U152, P3_INSTADDRPOINTER_REG_27__SCAN_IN, P3_ADD_547_U57);
  nand ginst22497 (P3_ADD_547_U153, P3_ADD_547_U123, P3_ADD_547_U58);
  nand ginst22498 (P3_ADD_547_U154, P3_INSTADDRPOINTER_REG_26__SCAN_IN, P3_ADD_547_U55);
  nand ginst22499 (P3_ADD_547_U155, P3_ADD_547_U122, P3_ADD_547_U56);
  nand ginst22500 (P3_ADD_547_U156, P3_INSTADDRPOINTER_REG_25__SCAN_IN, P3_ADD_547_U53);
  nand ginst22501 (P3_ADD_547_U157, P3_ADD_547_U121, P3_ADD_547_U54);
  nand ginst22502 (P3_ADD_547_U158, P3_INSTADDRPOINTER_REG_24__SCAN_IN, P3_ADD_547_U51);
  nand ginst22503 (P3_ADD_547_U159, P3_ADD_547_U120, P3_ADD_547_U52);
  not ginst22504 (P3_ADD_547_U16, P3_INSTADDRPOINTER_REG_6__SCAN_IN);
  nand ginst22505 (P3_ADD_547_U160, P3_INSTADDRPOINTER_REG_23__SCAN_IN, P3_ADD_547_U49);
  nand ginst22506 (P3_ADD_547_U161, P3_ADD_547_U119, P3_ADD_547_U50);
  nand ginst22507 (P3_ADD_547_U162, P3_INSTADDRPOINTER_REG_22__SCAN_IN, P3_ADD_547_U47);
  nand ginst22508 (P3_ADD_547_U163, P3_ADD_547_U118, P3_ADD_547_U48);
  nand ginst22509 (P3_ADD_547_U164, P3_INSTADDRPOINTER_REG_21__SCAN_IN, P3_ADD_547_U45);
  nand ginst22510 (P3_ADD_547_U165, P3_ADD_547_U117, P3_ADD_547_U46);
  nand ginst22511 (P3_ADD_547_U166, P3_INSTADDRPOINTER_REG_20__SCAN_IN, P3_ADD_547_U43);
  nand ginst22512 (P3_ADD_547_U167, P3_ADD_547_U116, P3_ADD_547_U44);
  nand ginst22513 (P3_ADD_547_U168, P3_INSTADDRPOINTER_REG_1__SCAN_IN, P3_ADD_547_U5);
  nand ginst22514 (P3_ADD_547_U169, P3_INSTADDRPOINTER_REG_0__SCAN_IN, P3_ADD_547_U6);
  nand ginst22515 (P3_ADD_547_U17, P3_INSTADDRPOINTER_REG_6__SCAN_IN, P3_ADD_547_U102);
  nand ginst22516 (P3_ADD_547_U170, P3_INSTADDRPOINTER_REG_19__SCAN_IN, P3_ADD_547_U41);
  nand ginst22517 (P3_ADD_547_U171, P3_ADD_547_U115, P3_ADD_547_U42);
  nand ginst22518 (P3_ADD_547_U172, P3_INSTADDRPOINTER_REG_18__SCAN_IN, P3_ADD_547_U39);
  nand ginst22519 (P3_ADD_547_U173, P3_ADD_547_U114, P3_ADD_547_U40);
  nand ginst22520 (P3_ADD_547_U174, P3_INSTADDRPOINTER_REG_17__SCAN_IN, P3_ADD_547_U37);
  nand ginst22521 (P3_ADD_547_U175, P3_ADD_547_U113, P3_ADD_547_U38);
  nand ginst22522 (P3_ADD_547_U176, P3_INSTADDRPOINTER_REG_16__SCAN_IN, P3_ADD_547_U35);
  nand ginst22523 (P3_ADD_547_U177, P3_ADD_547_U112, P3_ADD_547_U36);
  nand ginst22524 (P3_ADD_547_U178, P3_INSTADDRPOINTER_REG_15__SCAN_IN, P3_ADD_547_U33);
  nand ginst22525 (P3_ADD_547_U179, P3_ADD_547_U111, P3_ADD_547_U34);
  not ginst22526 (P3_ADD_547_U18, P3_INSTADDRPOINTER_REG_7__SCAN_IN);
  nand ginst22527 (P3_ADD_547_U180, P3_INSTADDRPOINTER_REG_14__SCAN_IN, P3_ADD_547_U31);
  nand ginst22528 (P3_ADD_547_U181, P3_ADD_547_U110, P3_ADD_547_U32);
  nand ginst22529 (P3_ADD_547_U182, P3_INSTADDRPOINTER_REG_13__SCAN_IN, P3_ADD_547_U29);
  nand ginst22530 (P3_ADD_547_U183, P3_ADD_547_U109, P3_ADD_547_U30);
  nand ginst22531 (P3_ADD_547_U184, P3_INSTADDRPOINTER_REG_12__SCAN_IN, P3_ADD_547_U27);
  nand ginst22532 (P3_ADD_547_U185, P3_ADD_547_U108, P3_ADD_547_U28);
  nand ginst22533 (P3_ADD_547_U186, P3_INSTADDRPOINTER_REG_11__SCAN_IN, P3_ADD_547_U25);
  nand ginst22534 (P3_ADD_547_U187, P3_ADD_547_U107, P3_ADD_547_U26);
  nand ginst22535 (P3_ADD_547_U188, P3_INSTADDRPOINTER_REG_10__SCAN_IN, P3_ADD_547_U23);
  nand ginst22536 (P3_ADD_547_U189, P3_ADD_547_U106, P3_ADD_547_U24);
  nand ginst22537 (P3_ADD_547_U19, P3_INSTADDRPOINTER_REG_7__SCAN_IN, P3_ADD_547_U103);
  not ginst22538 (P3_ADD_547_U20, P3_INSTADDRPOINTER_REG_8__SCAN_IN);
  not ginst22539 (P3_ADD_547_U21, P3_INSTADDRPOINTER_REG_9__SCAN_IN);
  nand ginst22540 (P3_ADD_547_U22, P3_INSTADDRPOINTER_REG_8__SCAN_IN, P3_ADD_547_U104);
  nand ginst22541 (P3_ADD_547_U23, P3_INSTADDRPOINTER_REG_9__SCAN_IN, P3_ADD_547_U105);
  not ginst22542 (P3_ADD_547_U24, P3_INSTADDRPOINTER_REG_10__SCAN_IN);
  nand ginst22543 (P3_ADD_547_U25, P3_INSTADDRPOINTER_REG_10__SCAN_IN, P3_ADD_547_U106);
  not ginst22544 (P3_ADD_547_U26, P3_INSTADDRPOINTER_REG_11__SCAN_IN);
  nand ginst22545 (P3_ADD_547_U27, P3_INSTADDRPOINTER_REG_11__SCAN_IN, P3_ADD_547_U107);
  not ginst22546 (P3_ADD_547_U28, P3_INSTADDRPOINTER_REG_12__SCAN_IN);
  nand ginst22547 (P3_ADD_547_U29, P3_INSTADDRPOINTER_REG_12__SCAN_IN, P3_ADD_547_U108);
  not ginst22548 (P3_ADD_547_U30, P3_INSTADDRPOINTER_REG_13__SCAN_IN);
  nand ginst22549 (P3_ADD_547_U31, P3_INSTADDRPOINTER_REG_13__SCAN_IN, P3_ADD_547_U109);
  not ginst22550 (P3_ADD_547_U32, P3_INSTADDRPOINTER_REG_14__SCAN_IN);
  nand ginst22551 (P3_ADD_547_U33, P3_INSTADDRPOINTER_REG_14__SCAN_IN, P3_ADD_547_U110);
  not ginst22552 (P3_ADD_547_U34, P3_INSTADDRPOINTER_REG_15__SCAN_IN);
  nand ginst22553 (P3_ADD_547_U35, P3_INSTADDRPOINTER_REG_15__SCAN_IN, P3_ADD_547_U111);
  not ginst22554 (P3_ADD_547_U36, P3_INSTADDRPOINTER_REG_16__SCAN_IN);
  nand ginst22555 (P3_ADD_547_U37, P3_INSTADDRPOINTER_REG_16__SCAN_IN, P3_ADD_547_U112);
  not ginst22556 (P3_ADD_547_U38, P3_INSTADDRPOINTER_REG_17__SCAN_IN);
  nand ginst22557 (P3_ADD_547_U39, P3_INSTADDRPOINTER_REG_17__SCAN_IN, P3_ADD_547_U113);
  not ginst22558 (P3_ADD_547_U40, P3_INSTADDRPOINTER_REG_18__SCAN_IN);
  nand ginst22559 (P3_ADD_547_U41, P3_INSTADDRPOINTER_REG_18__SCAN_IN, P3_ADD_547_U114);
  not ginst22560 (P3_ADD_547_U42, P3_INSTADDRPOINTER_REG_19__SCAN_IN);
  nand ginst22561 (P3_ADD_547_U43, P3_INSTADDRPOINTER_REG_19__SCAN_IN, P3_ADD_547_U115);
  not ginst22562 (P3_ADD_547_U44, P3_INSTADDRPOINTER_REG_20__SCAN_IN);
  nand ginst22563 (P3_ADD_547_U45, P3_INSTADDRPOINTER_REG_20__SCAN_IN, P3_ADD_547_U116);
  not ginst22564 (P3_ADD_547_U46, P3_INSTADDRPOINTER_REG_21__SCAN_IN);
  nand ginst22565 (P3_ADD_547_U47, P3_INSTADDRPOINTER_REG_21__SCAN_IN, P3_ADD_547_U117);
  not ginst22566 (P3_ADD_547_U48, P3_INSTADDRPOINTER_REG_22__SCAN_IN);
  nand ginst22567 (P3_ADD_547_U49, P3_INSTADDRPOINTER_REG_22__SCAN_IN, P3_ADD_547_U118);
  not ginst22568 (P3_ADD_547_U5, P3_INSTADDRPOINTER_REG_0__SCAN_IN);
  not ginst22569 (P3_ADD_547_U50, P3_INSTADDRPOINTER_REG_23__SCAN_IN);
  nand ginst22570 (P3_ADD_547_U51, P3_INSTADDRPOINTER_REG_23__SCAN_IN, P3_ADD_547_U119);
  not ginst22571 (P3_ADD_547_U52, P3_INSTADDRPOINTER_REG_24__SCAN_IN);
  nand ginst22572 (P3_ADD_547_U53, P3_INSTADDRPOINTER_REG_24__SCAN_IN, P3_ADD_547_U120);
  not ginst22573 (P3_ADD_547_U54, P3_INSTADDRPOINTER_REG_25__SCAN_IN);
  nand ginst22574 (P3_ADD_547_U55, P3_INSTADDRPOINTER_REG_25__SCAN_IN, P3_ADD_547_U121);
  not ginst22575 (P3_ADD_547_U56, P3_INSTADDRPOINTER_REG_26__SCAN_IN);
  nand ginst22576 (P3_ADD_547_U57, P3_INSTADDRPOINTER_REG_26__SCAN_IN, P3_ADD_547_U122);
  not ginst22577 (P3_ADD_547_U58, P3_INSTADDRPOINTER_REG_27__SCAN_IN);
  nand ginst22578 (P3_ADD_547_U59, P3_INSTADDRPOINTER_REG_27__SCAN_IN, P3_ADD_547_U123);
  not ginst22579 (P3_ADD_547_U6, P3_INSTADDRPOINTER_REG_1__SCAN_IN);
  not ginst22580 (P3_ADD_547_U60, P3_INSTADDRPOINTER_REG_28__SCAN_IN);
  nand ginst22581 (P3_ADD_547_U61, P3_INSTADDRPOINTER_REG_28__SCAN_IN, P3_ADD_547_U124);
  not ginst22582 (P3_ADD_547_U62, P3_INSTADDRPOINTER_REG_29__SCAN_IN);
  nand ginst22583 (P3_ADD_547_U63, P3_INSTADDRPOINTER_REG_29__SCAN_IN, P3_ADD_547_U125);
  not ginst22584 (P3_ADD_547_U64, P3_INSTADDRPOINTER_REG_30__SCAN_IN);
  nand ginst22585 (P3_ADD_547_U65, P3_ADD_547_U128, P3_ADD_547_U129);
  nand ginst22586 (P3_ADD_547_U66, P3_ADD_547_U130, P3_ADD_547_U131);
  nand ginst22587 (P3_ADD_547_U67, P3_ADD_547_U132, P3_ADD_547_U133);
  nand ginst22588 (P3_ADD_547_U68, P3_ADD_547_U134, P3_ADD_547_U135);
  nand ginst22589 (P3_ADD_547_U69, P3_ADD_547_U136, P3_ADD_547_U137);
  nand ginst22590 (P3_ADD_547_U7, P3_INSTADDRPOINTER_REG_0__SCAN_IN, P3_INSTADDRPOINTER_REG_1__SCAN_IN);
  nand ginst22591 (P3_ADD_547_U70, P3_ADD_547_U138, P3_ADD_547_U139);
  nand ginst22592 (P3_ADD_547_U71, P3_ADD_547_U140, P3_ADD_547_U141);
  nand ginst22593 (P3_ADD_547_U72, P3_ADD_547_U142, P3_ADD_547_U143);
  nand ginst22594 (P3_ADD_547_U73, P3_ADD_547_U144, P3_ADD_547_U145);
  nand ginst22595 (P3_ADD_547_U74, P3_ADD_547_U146, P3_ADD_547_U147);
  nand ginst22596 (P3_ADD_547_U75, P3_ADD_547_U148, P3_ADD_547_U149);
  nand ginst22597 (P3_ADD_547_U76, P3_ADD_547_U150, P3_ADD_547_U151);
  nand ginst22598 (P3_ADD_547_U77, P3_ADD_547_U152, P3_ADD_547_U153);
  nand ginst22599 (P3_ADD_547_U78, P3_ADD_547_U154, P3_ADD_547_U155);
  nand ginst22600 (P3_ADD_547_U79, P3_ADD_547_U156, P3_ADD_547_U157);
  not ginst22601 (P3_ADD_547_U8, P3_INSTADDRPOINTER_REG_2__SCAN_IN);
  nand ginst22602 (P3_ADD_547_U80, P3_ADD_547_U158, P3_ADD_547_U159);
  nand ginst22603 (P3_ADD_547_U81, P3_ADD_547_U160, P3_ADD_547_U161);
  nand ginst22604 (P3_ADD_547_U82, P3_ADD_547_U162, P3_ADD_547_U163);
  nand ginst22605 (P3_ADD_547_U83, P3_ADD_547_U164, P3_ADD_547_U165);
  nand ginst22606 (P3_ADD_547_U84, P3_ADD_547_U166, P3_ADD_547_U167);
  nand ginst22607 (P3_ADD_547_U85, P3_ADD_547_U168, P3_ADD_547_U169);
  nand ginst22608 (P3_ADD_547_U86, P3_ADD_547_U170, P3_ADD_547_U171);
  nand ginst22609 (P3_ADD_547_U87, P3_ADD_547_U172, P3_ADD_547_U173);
  nand ginst22610 (P3_ADD_547_U88, P3_ADD_547_U174, P3_ADD_547_U175);
  nand ginst22611 (P3_ADD_547_U89, P3_ADD_547_U176, P3_ADD_547_U177);
  nand ginst22612 (P3_ADD_547_U9, P3_INSTADDRPOINTER_REG_2__SCAN_IN, P3_ADD_547_U98);
  nand ginst22613 (P3_ADD_547_U90, P3_ADD_547_U178, P3_ADD_547_U179);
  nand ginst22614 (P3_ADD_547_U91, P3_ADD_547_U180, P3_ADD_547_U181);
  nand ginst22615 (P3_ADD_547_U92, P3_ADD_547_U182, P3_ADD_547_U183);
  nand ginst22616 (P3_ADD_547_U93, P3_ADD_547_U184, P3_ADD_547_U185);
  nand ginst22617 (P3_ADD_547_U94, P3_ADD_547_U186, P3_ADD_547_U187);
  nand ginst22618 (P3_ADD_547_U95, P3_ADD_547_U188, P3_ADD_547_U189);
  not ginst22619 (P3_ADD_547_U96, P3_INSTADDRPOINTER_REG_31__SCAN_IN);
  nand ginst22620 (P3_ADD_547_U97, P3_INSTADDRPOINTER_REG_30__SCAN_IN, P3_ADD_547_U126);
  not ginst22621 (P3_ADD_547_U98, P3_ADD_547_U7);
  not ginst22622 (P3_ADD_547_U99, P3_ADD_547_U9);
  nand ginst22623 (P3_ADD_552_U10, P3_EBX_REG_0__SCAN_IN, P3_EBX_REG_1__SCAN_IN, P3_EBX_REG_2__SCAN_IN);
  nand ginst22624 (P3_ADD_552_U100, P3_EBX_REG_0__SCAN_IN, P3_EBX_REG_1__SCAN_IN);
  nand ginst22625 (P3_ADD_552_U101, P3_EBX_REG_27__SCAN_IN, P3_ADD_552_U122);
  nand ginst22626 (P3_ADD_552_U102, P3_EBX_REG_25__SCAN_IN, P3_ADD_552_U116);
  nand ginst22627 (P3_ADD_552_U103, P3_EBX_REG_23__SCAN_IN, P3_ADD_552_U115);
  nand ginst22628 (P3_ADD_552_U104, P3_EBX_REG_21__SCAN_IN, P3_ADD_552_U121);
  nand ginst22629 (P3_ADD_552_U105, P3_EBX_REG_19__SCAN_IN, P3_ADD_552_U114);
  nand ginst22630 (P3_ADD_552_U106, P3_EBX_REG_17__SCAN_IN, P3_ADD_552_U117);
  nand ginst22631 (P3_ADD_552_U107, P3_EBX_REG_15__SCAN_IN, P3_ADD_552_U124);
  nand ginst22632 (P3_ADD_552_U108, P3_EBX_REG_13__SCAN_IN, P3_ADD_552_U119);
  nand ginst22633 (P3_ADD_552_U109, P3_EBX_REG_11__SCAN_IN, P3_ADD_552_U113);
  not ginst22634 (P3_ADD_552_U11, P3_EBX_REG_6__SCAN_IN);
  nand ginst22635 (P3_ADD_552_U110, P3_EBX_REG_9__SCAN_IN, P3_ADD_552_U120);
  not ginst22636 (P3_ADD_552_U111, P3_ADD_552_U10);
  not ginst22637 (P3_ADD_552_U112, P3_ADD_552_U13);
  not ginst22638 (P3_ADD_552_U113, P3_ADD_552_U22);
  not ginst22639 (P3_ADD_552_U114, P3_ADD_552_U34);
  not ginst22640 (P3_ADD_552_U115, P3_ADD_552_U40);
  not ginst22641 (P3_ADD_552_U116, P3_ADD_552_U43);
  not ginst22642 (P3_ADD_552_U117, P3_ADD_552_U31);
  not ginst22643 (P3_ADD_552_U118, P3_ADD_552_U16);
  not ginst22644 (P3_ADD_552_U119, P3_ADD_552_U25);
  not ginst22645 (P3_ADD_552_U12, P3_EBX_REG_5__SCAN_IN);
  not ginst22646 (P3_ADD_552_U120, P3_ADD_552_U17);
  not ginst22647 (P3_ADD_552_U121, P3_ADD_552_U36);
  not ginst22648 (P3_ADD_552_U122, P3_ADD_552_U46);
  not ginst22649 (P3_ADD_552_U123, P3_ADD_552_U48);
  not ginst22650 (P3_ADD_552_U124, P3_ADD_552_U27);
  not ginst22651 (P3_ADD_552_U125, P3_ADD_552_U95);
  not ginst22652 (P3_ADD_552_U126, P3_ADD_552_U96);
  not ginst22653 (P3_ADD_552_U127, P3_ADD_552_U97);
  not ginst22654 (P3_ADD_552_U128, P3_ADD_552_U49);
  not ginst22655 (P3_ADD_552_U129, P3_ADD_552_U99);
  nand ginst22656 (P3_ADD_552_U13, P3_ADD_552_U111, P3_ADD_552_U82);
  not ginst22657 (P3_ADD_552_U130, P3_ADD_552_U100);
  not ginst22658 (P3_ADD_552_U131, P3_ADD_552_U101);
  not ginst22659 (P3_ADD_552_U132, P3_ADD_552_U102);
  not ginst22660 (P3_ADD_552_U133, P3_ADD_552_U103);
  not ginst22661 (P3_ADD_552_U134, P3_ADD_552_U104);
  not ginst22662 (P3_ADD_552_U135, P3_ADD_552_U105);
  not ginst22663 (P3_ADD_552_U136, P3_ADD_552_U106);
  not ginst22664 (P3_ADD_552_U137, P3_ADD_552_U107);
  not ginst22665 (P3_ADD_552_U138, P3_ADD_552_U108);
  not ginst22666 (P3_ADD_552_U139, P3_ADD_552_U109);
  not ginst22667 (P3_ADD_552_U14, P3_EBX_REG_8__SCAN_IN);
  not ginst22668 (P3_ADD_552_U140, P3_ADD_552_U110);
  nand ginst22669 (P3_ADD_552_U141, P3_ADD_552_U120, P3_ADD_552_U18);
  nand ginst22670 (P3_ADD_552_U142, P3_EBX_REG_9__SCAN_IN, P3_ADD_552_U17);
  nand ginst22671 (P3_ADD_552_U143, P3_EBX_REG_8__SCAN_IN, P3_ADD_552_U95);
  nand ginst22672 (P3_ADD_552_U144, P3_ADD_552_U125, P3_ADD_552_U14);
  nand ginst22673 (P3_ADD_552_U145, P3_ADD_552_U118, P3_ADD_552_U15);
  nand ginst22674 (P3_ADD_552_U146, P3_EBX_REG_7__SCAN_IN, P3_ADD_552_U16);
  nand ginst22675 (P3_ADD_552_U147, P3_EBX_REG_6__SCAN_IN, P3_ADD_552_U96);
  nand ginst22676 (P3_ADD_552_U148, P3_ADD_552_U11, P3_ADD_552_U126);
  nand ginst22677 (P3_ADD_552_U149, P3_ADD_552_U112, P3_ADD_552_U12);
  not ginst22678 (P3_ADD_552_U15, P3_EBX_REG_7__SCAN_IN);
  nand ginst22679 (P3_ADD_552_U150, P3_EBX_REG_5__SCAN_IN, P3_ADD_552_U13);
  nand ginst22680 (P3_ADD_552_U151, P3_EBX_REG_4__SCAN_IN, P3_ADD_552_U97);
  nand ginst22681 (P3_ADD_552_U152, P3_ADD_552_U127, P3_ADD_552_U8);
  nand ginst22682 (P3_ADD_552_U153, P3_ADD_552_U111, P3_ADD_552_U9);
  nand ginst22683 (P3_ADD_552_U154, P3_EBX_REG_3__SCAN_IN, P3_ADD_552_U10);
  nand ginst22684 (P3_ADD_552_U155, P3_EBX_REG_31__SCAN_IN, P3_ADD_552_U99);
  nand ginst22685 (P3_ADD_552_U156, P3_ADD_552_U129, P3_ADD_552_U98);
  nand ginst22686 (P3_ADD_552_U157, P3_EBX_REG_30__SCAN_IN, P3_ADD_552_U49);
  nand ginst22687 (P3_ADD_552_U158, P3_ADD_552_U128, P3_ADD_552_U50);
  nand ginst22688 (P3_ADD_552_U159, P3_EBX_REG_2__SCAN_IN, P3_ADD_552_U100);
  nand ginst22689 (P3_ADD_552_U16, P3_ADD_552_U112, P3_ADD_552_U83);
  nand ginst22690 (P3_ADD_552_U160, P3_ADD_552_U130, P3_ADD_552_U6);
  nand ginst22691 (P3_ADD_552_U161, P3_ADD_552_U123, P3_ADD_552_U47);
  nand ginst22692 (P3_ADD_552_U162, P3_EBX_REG_29__SCAN_IN, P3_ADD_552_U48);
  nand ginst22693 (P3_ADD_552_U163, P3_EBX_REG_28__SCAN_IN, P3_ADD_552_U101);
  nand ginst22694 (P3_ADD_552_U164, P3_ADD_552_U131, P3_ADD_552_U45);
  nand ginst22695 (P3_ADD_552_U165, P3_ADD_552_U122, P3_ADD_552_U44);
  nand ginst22696 (P3_ADD_552_U166, P3_EBX_REG_27__SCAN_IN, P3_ADD_552_U46);
  nand ginst22697 (P3_ADD_552_U167, P3_EBX_REG_26__SCAN_IN, P3_ADD_552_U102);
  nand ginst22698 (P3_ADD_552_U168, P3_ADD_552_U132, P3_ADD_552_U41);
  nand ginst22699 (P3_ADD_552_U169, P3_ADD_552_U116, P3_ADD_552_U42);
  nand ginst22700 (P3_ADD_552_U17, P3_ADD_552_U118, P3_ADD_552_U84);
  nand ginst22701 (P3_ADD_552_U170, P3_EBX_REG_25__SCAN_IN, P3_ADD_552_U43);
  nand ginst22702 (P3_ADD_552_U171, P3_EBX_REG_24__SCAN_IN, P3_ADD_552_U103);
  nand ginst22703 (P3_ADD_552_U172, P3_ADD_552_U133, P3_ADD_552_U38);
  nand ginst22704 (P3_ADD_552_U173, P3_ADD_552_U115, P3_ADD_552_U39);
  nand ginst22705 (P3_ADD_552_U174, P3_EBX_REG_23__SCAN_IN, P3_ADD_552_U40);
  nand ginst22706 (P3_ADD_552_U175, P3_EBX_REG_22__SCAN_IN, P3_ADD_552_U104);
  nand ginst22707 (P3_ADD_552_U176, P3_ADD_552_U134, P3_ADD_552_U37);
  nand ginst22708 (P3_ADD_552_U177, P3_ADD_552_U121, P3_ADD_552_U35);
  nand ginst22709 (P3_ADD_552_U178, P3_EBX_REG_21__SCAN_IN, P3_ADD_552_U36);
  nand ginst22710 (P3_ADD_552_U179, P3_EBX_REG_20__SCAN_IN, P3_ADD_552_U105);
  not ginst22711 (P3_ADD_552_U18, P3_EBX_REG_9__SCAN_IN);
  nand ginst22712 (P3_ADD_552_U180, P3_ADD_552_U135, P3_ADD_552_U32);
  nand ginst22713 (P3_ADD_552_U181, P3_EBX_REG_0__SCAN_IN, P3_ADD_552_U7);
  nand ginst22714 (P3_ADD_552_U182, P3_EBX_REG_1__SCAN_IN, P3_ADD_552_U5);
  nand ginst22715 (P3_ADD_552_U183, P3_ADD_552_U114, P3_ADD_552_U33);
  nand ginst22716 (P3_ADD_552_U184, P3_EBX_REG_19__SCAN_IN, P3_ADD_552_U34);
  nand ginst22717 (P3_ADD_552_U185, P3_EBX_REG_18__SCAN_IN, P3_ADD_552_U106);
  nand ginst22718 (P3_ADD_552_U186, P3_ADD_552_U136, P3_ADD_552_U29);
  nand ginst22719 (P3_ADD_552_U187, P3_ADD_552_U117, P3_ADD_552_U30);
  nand ginst22720 (P3_ADD_552_U188, P3_EBX_REG_17__SCAN_IN, P3_ADD_552_U31);
  nand ginst22721 (P3_ADD_552_U189, P3_EBX_REG_16__SCAN_IN, P3_ADD_552_U107);
  not ginst22722 (P3_ADD_552_U19, P3_EBX_REG_10__SCAN_IN);
  nand ginst22723 (P3_ADD_552_U190, P3_ADD_552_U137, P3_ADD_552_U28);
  nand ginst22724 (P3_ADD_552_U191, P3_ADD_552_U124, P3_ADD_552_U26);
  nand ginst22725 (P3_ADD_552_U192, P3_EBX_REG_15__SCAN_IN, P3_ADD_552_U27);
  nand ginst22726 (P3_ADD_552_U193, P3_EBX_REG_14__SCAN_IN, P3_ADD_552_U108);
  nand ginst22727 (P3_ADD_552_U194, P3_ADD_552_U138, P3_ADD_552_U23);
  nand ginst22728 (P3_ADD_552_U195, P3_ADD_552_U119, P3_ADD_552_U24);
  nand ginst22729 (P3_ADD_552_U196, P3_EBX_REG_13__SCAN_IN, P3_ADD_552_U25);
  nand ginst22730 (P3_ADD_552_U197, P3_EBX_REG_12__SCAN_IN, P3_ADD_552_U109);
  nand ginst22731 (P3_ADD_552_U198, P3_ADD_552_U139, P3_ADD_552_U20);
  nand ginst22732 (P3_ADD_552_U199, P3_ADD_552_U113, P3_ADD_552_U21);
  not ginst22733 (P3_ADD_552_U20, P3_EBX_REG_12__SCAN_IN);
  nand ginst22734 (P3_ADD_552_U200, P3_EBX_REG_11__SCAN_IN, P3_ADD_552_U22);
  nand ginst22735 (P3_ADD_552_U201, P3_EBX_REG_10__SCAN_IN, P3_ADD_552_U110);
  nand ginst22736 (P3_ADD_552_U202, P3_ADD_552_U140, P3_ADD_552_U19);
  not ginst22737 (P3_ADD_552_U21, P3_EBX_REG_11__SCAN_IN);
  nand ginst22738 (P3_ADD_552_U22, P3_ADD_552_U120, P3_ADD_552_U85);
  not ginst22739 (P3_ADD_552_U23, P3_EBX_REG_14__SCAN_IN);
  not ginst22740 (P3_ADD_552_U24, P3_EBX_REG_13__SCAN_IN);
  nand ginst22741 (P3_ADD_552_U25, P3_ADD_552_U113, P3_ADD_552_U86);
  not ginst22742 (P3_ADD_552_U26, P3_EBX_REG_15__SCAN_IN);
  nand ginst22743 (P3_ADD_552_U27, P3_ADD_552_U119, P3_ADD_552_U87);
  not ginst22744 (P3_ADD_552_U28, P3_EBX_REG_16__SCAN_IN);
  not ginst22745 (P3_ADD_552_U29, P3_EBX_REG_18__SCAN_IN);
  not ginst22746 (P3_ADD_552_U30, P3_EBX_REG_17__SCAN_IN);
  nand ginst22747 (P3_ADD_552_U31, P3_ADD_552_U124, P3_ADD_552_U88);
  not ginst22748 (P3_ADD_552_U32, P3_EBX_REG_20__SCAN_IN);
  not ginst22749 (P3_ADD_552_U33, P3_EBX_REG_19__SCAN_IN);
  nand ginst22750 (P3_ADD_552_U34, P3_ADD_552_U117, P3_ADD_552_U89);
  not ginst22751 (P3_ADD_552_U35, P3_EBX_REG_21__SCAN_IN);
  nand ginst22752 (P3_ADD_552_U36, P3_ADD_552_U114, P3_ADD_552_U90);
  not ginst22753 (P3_ADD_552_U37, P3_EBX_REG_22__SCAN_IN);
  not ginst22754 (P3_ADD_552_U38, P3_EBX_REG_24__SCAN_IN);
  not ginst22755 (P3_ADD_552_U39, P3_EBX_REG_23__SCAN_IN);
  nand ginst22756 (P3_ADD_552_U40, P3_ADD_552_U121, P3_ADD_552_U91);
  not ginst22757 (P3_ADD_552_U41, P3_EBX_REG_26__SCAN_IN);
  not ginst22758 (P3_ADD_552_U42, P3_EBX_REG_25__SCAN_IN);
  nand ginst22759 (P3_ADD_552_U43, P3_ADD_552_U115, P3_ADD_552_U92);
  not ginst22760 (P3_ADD_552_U44, P3_EBX_REG_27__SCAN_IN);
  not ginst22761 (P3_ADD_552_U45, P3_EBX_REG_28__SCAN_IN);
  nand ginst22762 (P3_ADD_552_U46, P3_ADD_552_U116, P3_ADD_552_U93);
  not ginst22763 (P3_ADD_552_U47, P3_EBX_REG_29__SCAN_IN);
  nand ginst22764 (P3_ADD_552_U48, P3_ADD_552_U122, P3_ADD_552_U94);
  nand ginst22765 (P3_ADD_552_U49, P3_EBX_REG_29__SCAN_IN, P3_ADD_552_U123);
  not ginst22766 (P3_ADD_552_U5, P3_EBX_REG_0__SCAN_IN);
  not ginst22767 (P3_ADD_552_U50, P3_EBX_REG_30__SCAN_IN);
  nand ginst22768 (P3_ADD_552_U51, P3_ADD_552_U141, P3_ADD_552_U142);
  nand ginst22769 (P3_ADD_552_U52, P3_ADD_552_U143, P3_ADD_552_U144);
  nand ginst22770 (P3_ADD_552_U53, P3_ADD_552_U145, P3_ADD_552_U146);
  nand ginst22771 (P3_ADD_552_U54, P3_ADD_552_U147, P3_ADD_552_U148);
  nand ginst22772 (P3_ADD_552_U55, P3_ADD_552_U149, P3_ADD_552_U150);
  nand ginst22773 (P3_ADD_552_U56, P3_ADD_552_U151, P3_ADD_552_U152);
  nand ginst22774 (P3_ADD_552_U57, P3_ADD_552_U153, P3_ADD_552_U154);
  nand ginst22775 (P3_ADD_552_U58, P3_ADD_552_U155, P3_ADD_552_U156);
  nand ginst22776 (P3_ADD_552_U59, P3_ADD_552_U157, P3_ADD_552_U158);
  not ginst22777 (P3_ADD_552_U6, P3_EBX_REG_2__SCAN_IN);
  nand ginst22778 (P3_ADD_552_U60, P3_ADD_552_U159, P3_ADD_552_U160);
  nand ginst22779 (P3_ADD_552_U61, P3_ADD_552_U161, P3_ADD_552_U162);
  nand ginst22780 (P3_ADD_552_U62, P3_ADD_552_U163, P3_ADD_552_U164);
  nand ginst22781 (P3_ADD_552_U63, P3_ADD_552_U165, P3_ADD_552_U166);
  nand ginst22782 (P3_ADD_552_U64, P3_ADD_552_U167, P3_ADD_552_U168);
  nand ginst22783 (P3_ADD_552_U65, P3_ADD_552_U169, P3_ADD_552_U170);
  nand ginst22784 (P3_ADD_552_U66, P3_ADD_552_U171, P3_ADD_552_U172);
  nand ginst22785 (P3_ADD_552_U67, P3_ADD_552_U173, P3_ADD_552_U174);
  nand ginst22786 (P3_ADD_552_U68, P3_ADD_552_U175, P3_ADD_552_U176);
  nand ginst22787 (P3_ADD_552_U69, P3_ADD_552_U177, P3_ADD_552_U178);
  not ginst22788 (P3_ADD_552_U7, P3_EBX_REG_1__SCAN_IN);
  nand ginst22789 (P3_ADD_552_U70, P3_ADD_552_U179, P3_ADD_552_U180);
  nand ginst22790 (P3_ADD_552_U71, P3_ADD_552_U181, P3_ADD_552_U182);
  nand ginst22791 (P3_ADD_552_U72, P3_ADD_552_U183, P3_ADD_552_U184);
  nand ginst22792 (P3_ADD_552_U73, P3_ADD_552_U185, P3_ADD_552_U186);
  nand ginst22793 (P3_ADD_552_U74, P3_ADD_552_U187, P3_ADD_552_U188);
  nand ginst22794 (P3_ADD_552_U75, P3_ADD_552_U189, P3_ADD_552_U190);
  nand ginst22795 (P3_ADD_552_U76, P3_ADD_552_U191, P3_ADD_552_U192);
  nand ginst22796 (P3_ADD_552_U77, P3_ADD_552_U193, P3_ADD_552_U194);
  nand ginst22797 (P3_ADD_552_U78, P3_ADD_552_U195, P3_ADD_552_U196);
  nand ginst22798 (P3_ADD_552_U79, P3_ADD_552_U197, P3_ADD_552_U198);
  not ginst22799 (P3_ADD_552_U8, P3_EBX_REG_4__SCAN_IN);
  nand ginst22800 (P3_ADD_552_U80, P3_ADD_552_U199, P3_ADD_552_U200);
  nand ginst22801 (P3_ADD_552_U81, P3_ADD_552_U201, P3_ADD_552_U202);
  and ginst22802 (P3_ADD_552_U82, P3_EBX_REG_3__SCAN_IN, P3_EBX_REG_4__SCAN_IN);
  and ginst22803 (P3_ADD_552_U83, P3_EBX_REG_5__SCAN_IN, P3_EBX_REG_6__SCAN_IN);
  and ginst22804 (P3_ADD_552_U84, P3_EBX_REG_7__SCAN_IN, P3_EBX_REG_8__SCAN_IN);
  and ginst22805 (P3_ADD_552_U85, P3_EBX_REG_9__SCAN_IN, P3_EBX_REG_10__SCAN_IN);
  and ginst22806 (P3_ADD_552_U86, P3_EBX_REG_11__SCAN_IN, P3_EBX_REG_12__SCAN_IN);
  and ginst22807 (P3_ADD_552_U87, P3_EBX_REG_13__SCAN_IN, P3_EBX_REG_14__SCAN_IN);
  and ginst22808 (P3_ADD_552_U88, P3_EBX_REG_15__SCAN_IN, P3_EBX_REG_16__SCAN_IN);
  and ginst22809 (P3_ADD_552_U89, P3_EBX_REG_17__SCAN_IN, P3_EBX_REG_18__SCAN_IN);
  not ginst22810 (P3_ADD_552_U9, P3_EBX_REG_3__SCAN_IN);
  and ginst22811 (P3_ADD_552_U90, P3_EBX_REG_19__SCAN_IN, P3_EBX_REG_20__SCAN_IN);
  and ginst22812 (P3_ADD_552_U91, P3_EBX_REG_21__SCAN_IN, P3_EBX_REG_22__SCAN_IN);
  and ginst22813 (P3_ADD_552_U92, P3_EBX_REG_23__SCAN_IN, P3_EBX_REG_24__SCAN_IN);
  and ginst22814 (P3_ADD_552_U93, P3_EBX_REG_25__SCAN_IN, P3_EBX_REG_26__SCAN_IN);
  and ginst22815 (P3_ADD_552_U94, P3_EBX_REG_27__SCAN_IN, P3_EBX_REG_28__SCAN_IN);
  nand ginst22816 (P3_ADD_552_U95, P3_EBX_REG_7__SCAN_IN, P3_ADD_552_U118);
  nand ginst22817 (P3_ADD_552_U96, P3_EBX_REG_5__SCAN_IN, P3_ADD_552_U112);
  nand ginst22818 (P3_ADD_552_U97, P3_EBX_REG_3__SCAN_IN, P3_ADD_552_U111);
  not ginst22819 (P3_ADD_552_U98, P3_EBX_REG_31__SCAN_IN);
  nand ginst22820 (P3_ADD_552_U99, P3_EBX_REG_30__SCAN_IN, P3_ADD_552_U128);
  not ginst22821 (P3_ADD_553_U10, P3_INSTADDRPOINTER_REG_3__SCAN_IN);
  not ginst22822 (P3_ADD_553_U100, P3_ADD_553_U11);
  not ginst22823 (P3_ADD_553_U101, P3_ADD_553_U13);
  not ginst22824 (P3_ADD_553_U102, P3_ADD_553_U15);
  not ginst22825 (P3_ADD_553_U103, P3_ADD_553_U17);
  not ginst22826 (P3_ADD_553_U104, P3_ADD_553_U19);
  not ginst22827 (P3_ADD_553_U105, P3_ADD_553_U22);
  not ginst22828 (P3_ADD_553_U106, P3_ADD_553_U23);
  not ginst22829 (P3_ADD_553_U107, P3_ADD_553_U25);
  not ginst22830 (P3_ADD_553_U108, P3_ADD_553_U27);
  not ginst22831 (P3_ADD_553_U109, P3_ADD_553_U29);
  nand ginst22832 (P3_ADD_553_U11, P3_INSTADDRPOINTER_REG_3__SCAN_IN, P3_ADD_553_U99);
  not ginst22833 (P3_ADD_553_U110, P3_ADD_553_U31);
  not ginst22834 (P3_ADD_553_U111, P3_ADD_553_U33);
  not ginst22835 (P3_ADD_553_U112, P3_ADD_553_U35);
  not ginst22836 (P3_ADD_553_U113, P3_ADD_553_U37);
  not ginst22837 (P3_ADD_553_U114, P3_ADD_553_U39);
  not ginst22838 (P3_ADD_553_U115, P3_ADD_553_U41);
  not ginst22839 (P3_ADD_553_U116, P3_ADD_553_U43);
  not ginst22840 (P3_ADD_553_U117, P3_ADD_553_U45);
  not ginst22841 (P3_ADD_553_U118, P3_ADD_553_U47);
  not ginst22842 (P3_ADD_553_U119, P3_ADD_553_U49);
  not ginst22843 (P3_ADD_553_U12, P3_INSTADDRPOINTER_REG_4__SCAN_IN);
  not ginst22844 (P3_ADD_553_U120, P3_ADD_553_U51);
  not ginst22845 (P3_ADD_553_U121, P3_ADD_553_U53);
  not ginst22846 (P3_ADD_553_U122, P3_ADD_553_U55);
  not ginst22847 (P3_ADD_553_U123, P3_ADD_553_U57);
  not ginst22848 (P3_ADD_553_U124, P3_ADD_553_U59);
  not ginst22849 (P3_ADD_553_U125, P3_ADD_553_U61);
  not ginst22850 (P3_ADD_553_U126, P3_ADD_553_U63);
  not ginst22851 (P3_ADD_553_U127, P3_ADD_553_U97);
  nand ginst22852 (P3_ADD_553_U128, P3_INSTADDRPOINTER_REG_9__SCAN_IN, P3_ADD_553_U22);
  nand ginst22853 (P3_ADD_553_U129, P3_ADD_553_U105, P3_ADD_553_U21);
  nand ginst22854 (P3_ADD_553_U13, P3_INSTADDRPOINTER_REG_4__SCAN_IN, P3_ADD_553_U100);
  nand ginst22855 (P3_ADD_553_U130, P3_INSTADDRPOINTER_REG_8__SCAN_IN, P3_ADD_553_U19);
  nand ginst22856 (P3_ADD_553_U131, P3_ADD_553_U104, P3_ADD_553_U20);
  nand ginst22857 (P3_ADD_553_U132, P3_INSTADDRPOINTER_REG_7__SCAN_IN, P3_ADD_553_U17);
  nand ginst22858 (P3_ADD_553_U133, P3_ADD_553_U103, P3_ADD_553_U18);
  nand ginst22859 (P3_ADD_553_U134, P3_INSTADDRPOINTER_REG_6__SCAN_IN, P3_ADD_553_U15);
  nand ginst22860 (P3_ADD_553_U135, P3_ADD_553_U102, P3_ADD_553_U16);
  nand ginst22861 (P3_ADD_553_U136, P3_INSTADDRPOINTER_REG_5__SCAN_IN, P3_ADD_553_U13);
  nand ginst22862 (P3_ADD_553_U137, P3_ADD_553_U101, P3_ADD_553_U14);
  nand ginst22863 (P3_ADD_553_U138, P3_INSTADDRPOINTER_REG_4__SCAN_IN, P3_ADD_553_U11);
  nand ginst22864 (P3_ADD_553_U139, P3_ADD_553_U100, P3_ADD_553_U12);
  not ginst22865 (P3_ADD_553_U14, P3_INSTADDRPOINTER_REG_5__SCAN_IN);
  nand ginst22866 (P3_ADD_553_U140, P3_INSTADDRPOINTER_REG_3__SCAN_IN, P3_ADD_553_U9);
  nand ginst22867 (P3_ADD_553_U141, P3_ADD_553_U10, P3_ADD_553_U99);
  nand ginst22868 (P3_ADD_553_U142, P3_INSTADDRPOINTER_REG_31__SCAN_IN, P3_ADD_553_U97);
  nand ginst22869 (P3_ADD_553_U143, P3_ADD_553_U127, P3_ADD_553_U96);
  nand ginst22870 (P3_ADD_553_U144, P3_INSTADDRPOINTER_REG_30__SCAN_IN, P3_ADD_553_U63);
  nand ginst22871 (P3_ADD_553_U145, P3_ADD_553_U126, P3_ADD_553_U64);
  nand ginst22872 (P3_ADD_553_U146, P3_INSTADDRPOINTER_REG_2__SCAN_IN, P3_ADD_553_U7);
  nand ginst22873 (P3_ADD_553_U147, P3_ADD_553_U8, P3_ADD_553_U98);
  nand ginst22874 (P3_ADD_553_U148, P3_INSTADDRPOINTER_REG_29__SCAN_IN, P3_ADD_553_U61);
  nand ginst22875 (P3_ADD_553_U149, P3_ADD_553_U125, P3_ADD_553_U62);
  nand ginst22876 (P3_ADD_553_U15, P3_INSTADDRPOINTER_REG_5__SCAN_IN, P3_ADD_553_U101);
  nand ginst22877 (P3_ADD_553_U150, P3_INSTADDRPOINTER_REG_28__SCAN_IN, P3_ADD_553_U59);
  nand ginst22878 (P3_ADD_553_U151, P3_ADD_553_U124, P3_ADD_553_U60);
  nand ginst22879 (P3_ADD_553_U152, P3_INSTADDRPOINTER_REG_27__SCAN_IN, P3_ADD_553_U57);
  nand ginst22880 (P3_ADD_553_U153, P3_ADD_553_U123, P3_ADD_553_U58);
  nand ginst22881 (P3_ADD_553_U154, P3_INSTADDRPOINTER_REG_26__SCAN_IN, P3_ADD_553_U55);
  nand ginst22882 (P3_ADD_553_U155, P3_ADD_553_U122, P3_ADD_553_U56);
  nand ginst22883 (P3_ADD_553_U156, P3_INSTADDRPOINTER_REG_25__SCAN_IN, P3_ADD_553_U53);
  nand ginst22884 (P3_ADD_553_U157, P3_ADD_553_U121, P3_ADD_553_U54);
  nand ginst22885 (P3_ADD_553_U158, P3_INSTADDRPOINTER_REG_24__SCAN_IN, P3_ADD_553_U51);
  nand ginst22886 (P3_ADD_553_U159, P3_ADD_553_U120, P3_ADD_553_U52);
  not ginst22887 (P3_ADD_553_U16, P3_INSTADDRPOINTER_REG_6__SCAN_IN);
  nand ginst22888 (P3_ADD_553_U160, P3_INSTADDRPOINTER_REG_23__SCAN_IN, P3_ADD_553_U49);
  nand ginst22889 (P3_ADD_553_U161, P3_ADD_553_U119, P3_ADD_553_U50);
  nand ginst22890 (P3_ADD_553_U162, P3_INSTADDRPOINTER_REG_22__SCAN_IN, P3_ADD_553_U47);
  nand ginst22891 (P3_ADD_553_U163, P3_ADD_553_U118, P3_ADD_553_U48);
  nand ginst22892 (P3_ADD_553_U164, P3_INSTADDRPOINTER_REG_21__SCAN_IN, P3_ADD_553_U45);
  nand ginst22893 (P3_ADD_553_U165, P3_ADD_553_U117, P3_ADD_553_U46);
  nand ginst22894 (P3_ADD_553_U166, P3_INSTADDRPOINTER_REG_20__SCAN_IN, P3_ADD_553_U43);
  nand ginst22895 (P3_ADD_553_U167, P3_ADD_553_U116, P3_ADD_553_U44);
  nand ginst22896 (P3_ADD_553_U168, P3_INSTADDRPOINTER_REG_1__SCAN_IN, P3_ADD_553_U5);
  nand ginst22897 (P3_ADD_553_U169, P3_INSTADDRPOINTER_REG_0__SCAN_IN, P3_ADD_553_U6);
  nand ginst22898 (P3_ADD_553_U17, P3_INSTADDRPOINTER_REG_6__SCAN_IN, P3_ADD_553_U102);
  nand ginst22899 (P3_ADD_553_U170, P3_INSTADDRPOINTER_REG_19__SCAN_IN, P3_ADD_553_U41);
  nand ginst22900 (P3_ADD_553_U171, P3_ADD_553_U115, P3_ADD_553_U42);
  nand ginst22901 (P3_ADD_553_U172, P3_INSTADDRPOINTER_REG_18__SCAN_IN, P3_ADD_553_U39);
  nand ginst22902 (P3_ADD_553_U173, P3_ADD_553_U114, P3_ADD_553_U40);
  nand ginst22903 (P3_ADD_553_U174, P3_INSTADDRPOINTER_REG_17__SCAN_IN, P3_ADD_553_U37);
  nand ginst22904 (P3_ADD_553_U175, P3_ADD_553_U113, P3_ADD_553_U38);
  nand ginst22905 (P3_ADD_553_U176, P3_INSTADDRPOINTER_REG_16__SCAN_IN, P3_ADD_553_U35);
  nand ginst22906 (P3_ADD_553_U177, P3_ADD_553_U112, P3_ADD_553_U36);
  nand ginst22907 (P3_ADD_553_U178, P3_INSTADDRPOINTER_REG_15__SCAN_IN, P3_ADD_553_U33);
  nand ginst22908 (P3_ADD_553_U179, P3_ADD_553_U111, P3_ADD_553_U34);
  not ginst22909 (P3_ADD_553_U18, P3_INSTADDRPOINTER_REG_7__SCAN_IN);
  nand ginst22910 (P3_ADD_553_U180, P3_INSTADDRPOINTER_REG_14__SCAN_IN, P3_ADD_553_U31);
  nand ginst22911 (P3_ADD_553_U181, P3_ADD_553_U110, P3_ADD_553_U32);
  nand ginst22912 (P3_ADD_553_U182, P3_INSTADDRPOINTER_REG_13__SCAN_IN, P3_ADD_553_U29);
  nand ginst22913 (P3_ADD_553_U183, P3_ADD_553_U109, P3_ADD_553_U30);
  nand ginst22914 (P3_ADD_553_U184, P3_INSTADDRPOINTER_REG_12__SCAN_IN, P3_ADD_553_U27);
  nand ginst22915 (P3_ADD_553_U185, P3_ADD_553_U108, P3_ADD_553_U28);
  nand ginst22916 (P3_ADD_553_U186, P3_INSTADDRPOINTER_REG_11__SCAN_IN, P3_ADD_553_U25);
  nand ginst22917 (P3_ADD_553_U187, P3_ADD_553_U107, P3_ADD_553_U26);
  nand ginst22918 (P3_ADD_553_U188, P3_INSTADDRPOINTER_REG_10__SCAN_IN, P3_ADD_553_U23);
  nand ginst22919 (P3_ADD_553_U189, P3_ADD_553_U106, P3_ADD_553_U24);
  nand ginst22920 (P3_ADD_553_U19, P3_INSTADDRPOINTER_REG_7__SCAN_IN, P3_ADD_553_U103);
  not ginst22921 (P3_ADD_553_U20, P3_INSTADDRPOINTER_REG_8__SCAN_IN);
  not ginst22922 (P3_ADD_553_U21, P3_INSTADDRPOINTER_REG_9__SCAN_IN);
  nand ginst22923 (P3_ADD_553_U22, P3_INSTADDRPOINTER_REG_8__SCAN_IN, P3_ADD_553_U104);
  nand ginst22924 (P3_ADD_553_U23, P3_INSTADDRPOINTER_REG_9__SCAN_IN, P3_ADD_553_U105);
  not ginst22925 (P3_ADD_553_U24, P3_INSTADDRPOINTER_REG_10__SCAN_IN);
  nand ginst22926 (P3_ADD_553_U25, P3_INSTADDRPOINTER_REG_10__SCAN_IN, P3_ADD_553_U106);
  not ginst22927 (P3_ADD_553_U26, P3_INSTADDRPOINTER_REG_11__SCAN_IN);
  nand ginst22928 (P3_ADD_553_U27, P3_INSTADDRPOINTER_REG_11__SCAN_IN, P3_ADD_553_U107);
  not ginst22929 (P3_ADD_553_U28, P3_INSTADDRPOINTER_REG_12__SCAN_IN);
  nand ginst22930 (P3_ADD_553_U29, P3_INSTADDRPOINTER_REG_12__SCAN_IN, P3_ADD_553_U108);
  not ginst22931 (P3_ADD_553_U30, P3_INSTADDRPOINTER_REG_13__SCAN_IN);
  nand ginst22932 (P3_ADD_553_U31, P3_INSTADDRPOINTER_REG_13__SCAN_IN, P3_ADD_553_U109);
  not ginst22933 (P3_ADD_553_U32, P3_INSTADDRPOINTER_REG_14__SCAN_IN);
  nand ginst22934 (P3_ADD_553_U33, P3_INSTADDRPOINTER_REG_14__SCAN_IN, P3_ADD_553_U110);
  not ginst22935 (P3_ADD_553_U34, P3_INSTADDRPOINTER_REG_15__SCAN_IN);
  nand ginst22936 (P3_ADD_553_U35, P3_INSTADDRPOINTER_REG_15__SCAN_IN, P3_ADD_553_U111);
  not ginst22937 (P3_ADD_553_U36, P3_INSTADDRPOINTER_REG_16__SCAN_IN);
  nand ginst22938 (P3_ADD_553_U37, P3_INSTADDRPOINTER_REG_16__SCAN_IN, P3_ADD_553_U112);
  not ginst22939 (P3_ADD_553_U38, P3_INSTADDRPOINTER_REG_17__SCAN_IN);
  nand ginst22940 (P3_ADD_553_U39, P3_INSTADDRPOINTER_REG_17__SCAN_IN, P3_ADD_553_U113);
  not ginst22941 (P3_ADD_553_U40, P3_INSTADDRPOINTER_REG_18__SCAN_IN);
  nand ginst22942 (P3_ADD_553_U41, P3_INSTADDRPOINTER_REG_18__SCAN_IN, P3_ADD_553_U114);
  not ginst22943 (P3_ADD_553_U42, P3_INSTADDRPOINTER_REG_19__SCAN_IN);
  nand ginst22944 (P3_ADD_553_U43, P3_INSTADDRPOINTER_REG_19__SCAN_IN, P3_ADD_553_U115);
  not ginst22945 (P3_ADD_553_U44, P3_INSTADDRPOINTER_REG_20__SCAN_IN);
  nand ginst22946 (P3_ADD_553_U45, P3_INSTADDRPOINTER_REG_20__SCAN_IN, P3_ADD_553_U116);
  not ginst22947 (P3_ADD_553_U46, P3_INSTADDRPOINTER_REG_21__SCAN_IN);
  nand ginst22948 (P3_ADD_553_U47, P3_INSTADDRPOINTER_REG_21__SCAN_IN, P3_ADD_553_U117);
  not ginst22949 (P3_ADD_553_U48, P3_INSTADDRPOINTER_REG_22__SCAN_IN);
  nand ginst22950 (P3_ADD_553_U49, P3_INSTADDRPOINTER_REG_22__SCAN_IN, P3_ADD_553_U118);
  not ginst22951 (P3_ADD_553_U5, P3_INSTADDRPOINTER_REG_0__SCAN_IN);
  not ginst22952 (P3_ADD_553_U50, P3_INSTADDRPOINTER_REG_23__SCAN_IN);
  nand ginst22953 (P3_ADD_553_U51, P3_INSTADDRPOINTER_REG_23__SCAN_IN, P3_ADD_553_U119);
  not ginst22954 (P3_ADD_553_U52, P3_INSTADDRPOINTER_REG_24__SCAN_IN);
  nand ginst22955 (P3_ADD_553_U53, P3_INSTADDRPOINTER_REG_24__SCAN_IN, P3_ADD_553_U120);
  not ginst22956 (P3_ADD_553_U54, P3_INSTADDRPOINTER_REG_25__SCAN_IN);
  nand ginst22957 (P3_ADD_553_U55, P3_INSTADDRPOINTER_REG_25__SCAN_IN, P3_ADD_553_U121);
  not ginst22958 (P3_ADD_553_U56, P3_INSTADDRPOINTER_REG_26__SCAN_IN);
  nand ginst22959 (P3_ADD_553_U57, P3_INSTADDRPOINTER_REG_26__SCAN_IN, P3_ADD_553_U122);
  not ginst22960 (P3_ADD_553_U58, P3_INSTADDRPOINTER_REG_27__SCAN_IN);
  nand ginst22961 (P3_ADD_553_U59, P3_INSTADDRPOINTER_REG_27__SCAN_IN, P3_ADD_553_U123);
  not ginst22962 (P3_ADD_553_U6, P3_INSTADDRPOINTER_REG_1__SCAN_IN);
  not ginst22963 (P3_ADD_553_U60, P3_INSTADDRPOINTER_REG_28__SCAN_IN);
  nand ginst22964 (P3_ADD_553_U61, P3_INSTADDRPOINTER_REG_28__SCAN_IN, P3_ADD_553_U124);
  not ginst22965 (P3_ADD_553_U62, P3_INSTADDRPOINTER_REG_29__SCAN_IN);
  nand ginst22966 (P3_ADD_553_U63, P3_INSTADDRPOINTER_REG_29__SCAN_IN, P3_ADD_553_U125);
  not ginst22967 (P3_ADD_553_U64, P3_INSTADDRPOINTER_REG_30__SCAN_IN);
  nand ginst22968 (P3_ADD_553_U65, P3_ADD_553_U128, P3_ADD_553_U129);
  nand ginst22969 (P3_ADD_553_U66, P3_ADD_553_U130, P3_ADD_553_U131);
  nand ginst22970 (P3_ADD_553_U67, P3_ADD_553_U132, P3_ADD_553_U133);
  nand ginst22971 (P3_ADD_553_U68, P3_ADD_553_U134, P3_ADD_553_U135);
  nand ginst22972 (P3_ADD_553_U69, P3_ADD_553_U136, P3_ADD_553_U137);
  nand ginst22973 (P3_ADD_553_U7, P3_INSTADDRPOINTER_REG_0__SCAN_IN, P3_INSTADDRPOINTER_REG_1__SCAN_IN);
  nand ginst22974 (P3_ADD_553_U70, P3_ADD_553_U138, P3_ADD_553_U139);
  nand ginst22975 (P3_ADD_553_U71, P3_ADD_553_U140, P3_ADD_553_U141);
  nand ginst22976 (P3_ADD_553_U72, P3_ADD_553_U142, P3_ADD_553_U143);
  nand ginst22977 (P3_ADD_553_U73, P3_ADD_553_U144, P3_ADD_553_U145);
  nand ginst22978 (P3_ADD_553_U74, P3_ADD_553_U146, P3_ADD_553_U147);
  nand ginst22979 (P3_ADD_553_U75, P3_ADD_553_U148, P3_ADD_553_U149);
  nand ginst22980 (P3_ADD_553_U76, P3_ADD_553_U150, P3_ADD_553_U151);
  nand ginst22981 (P3_ADD_553_U77, P3_ADD_553_U152, P3_ADD_553_U153);
  nand ginst22982 (P3_ADD_553_U78, P3_ADD_553_U154, P3_ADD_553_U155);
  nand ginst22983 (P3_ADD_553_U79, P3_ADD_553_U156, P3_ADD_553_U157);
  not ginst22984 (P3_ADD_553_U8, P3_INSTADDRPOINTER_REG_2__SCAN_IN);
  nand ginst22985 (P3_ADD_553_U80, P3_ADD_553_U158, P3_ADD_553_U159);
  nand ginst22986 (P3_ADD_553_U81, P3_ADD_553_U160, P3_ADD_553_U161);
  nand ginst22987 (P3_ADD_553_U82, P3_ADD_553_U162, P3_ADD_553_U163);
  nand ginst22988 (P3_ADD_553_U83, P3_ADD_553_U164, P3_ADD_553_U165);
  nand ginst22989 (P3_ADD_553_U84, P3_ADD_553_U166, P3_ADD_553_U167);
  nand ginst22990 (P3_ADD_553_U85, P3_ADD_553_U168, P3_ADD_553_U169);
  nand ginst22991 (P3_ADD_553_U86, P3_ADD_553_U170, P3_ADD_553_U171);
  nand ginst22992 (P3_ADD_553_U87, P3_ADD_553_U172, P3_ADD_553_U173);
  nand ginst22993 (P3_ADD_553_U88, P3_ADD_553_U174, P3_ADD_553_U175);
  nand ginst22994 (P3_ADD_553_U89, P3_ADD_553_U176, P3_ADD_553_U177);
  nand ginst22995 (P3_ADD_553_U9, P3_INSTADDRPOINTER_REG_2__SCAN_IN, P3_ADD_553_U98);
  nand ginst22996 (P3_ADD_553_U90, P3_ADD_553_U178, P3_ADD_553_U179);
  nand ginst22997 (P3_ADD_553_U91, P3_ADD_553_U180, P3_ADD_553_U181);
  nand ginst22998 (P3_ADD_553_U92, P3_ADD_553_U182, P3_ADD_553_U183);
  nand ginst22999 (P3_ADD_553_U93, P3_ADD_553_U184, P3_ADD_553_U185);
  nand ginst23000 (P3_ADD_553_U94, P3_ADD_553_U186, P3_ADD_553_U187);
  nand ginst23001 (P3_ADD_553_U95, P3_ADD_553_U188, P3_ADD_553_U189);
  not ginst23002 (P3_ADD_553_U96, P3_INSTADDRPOINTER_REG_31__SCAN_IN);
  nand ginst23003 (P3_ADD_553_U97, P3_INSTADDRPOINTER_REG_30__SCAN_IN, P3_ADD_553_U126);
  not ginst23004 (P3_ADD_553_U98, P3_ADD_553_U7);
  not ginst23005 (P3_ADD_553_U99, P3_ADD_553_U9);
  not ginst23006 (P3_ADD_558_U10, P3_INSTADDRPOINTER_REG_3__SCAN_IN);
  not ginst23007 (P3_ADD_558_U100, P3_ADD_558_U11);
  not ginst23008 (P3_ADD_558_U101, P3_ADD_558_U13);
  not ginst23009 (P3_ADD_558_U102, P3_ADD_558_U15);
  not ginst23010 (P3_ADD_558_U103, P3_ADD_558_U17);
  not ginst23011 (P3_ADD_558_U104, P3_ADD_558_U19);
  not ginst23012 (P3_ADD_558_U105, P3_ADD_558_U22);
  not ginst23013 (P3_ADD_558_U106, P3_ADD_558_U23);
  not ginst23014 (P3_ADD_558_U107, P3_ADD_558_U25);
  not ginst23015 (P3_ADD_558_U108, P3_ADD_558_U27);
  not ginst23016 (P3_ADD_558_U109, P3_ADD_558_U29);
  nand ginst23017 (P3_ADD_558_U11, P3_INSTADDRPOINTER_REG_3__SCAN_IN, P3_ADD_558_U99);
  not ginst23018 (P3_ADD_558_U110, P3_ADD_558_U31);
  not ginst23019 (P3_ADD_558_U111, P3_ADD_558_U33);
  not ginst23020 (P3_ADD_558_U112, P3_ADD_558_U35);
  not ginst23021 (P3_ADD_558_U113, P3_ADD_558_U37);
  not ginst23022 (P3_ADD_558_U114, P3_ADD_558_U39);
  not ginst23023 (P3_ADD_558_U115, P3_ADD_558_U41);
  not ginst23024 (P3_ADD_558_U116, P3_ADD_558_U43);
  not ginst23025 (P3_ADD_558_U117, P3_ADD_558_U45);
  not ginst23026 (P3_ADD_558_U118, P3_ADD_558_U47);
  not ginst23027 (P3_ADD_558_U119, P3_ADD_558_U49);
  not ginst23028 (P3_ADD_558_U12, P3_INSTADDRPOINTER_REG_4__SCAN_IN);
  not ginst23029 (P3_ADD_558_U120, P3_ADD_558_U51);
  not ginst23030 (P3_ADD_558_U121, P3_ADD_558_U53);
  not ginst23031 (P3_ADD_558_U122, P3_ADD_558_U55);
  not ginst23032 (P3_ADD_558_U123, P3_ADD_558_U57);
  not ginst23033 (P3_ADD_558_U124, P3_ADD_558_U59);
  not ginst23034 (P3_ADD_558_U125, P3_ADD_558_U61);
  not ginst23035 (P3_ADD_558_U126, P3_ADD_558_U63);
  not ginst23036 (P3_ADD_558_U127, P3_ADD_558_U97);
  nand ginst23037 (P3_ADD_558_U128, P3_INSTADDRPOINTER_REG_9__SCAN_IN, P3_ADD_558_U22);
  nand ginst23038 (P3_ADD_558_U129, P3_ADD_558_U105, P3_ADD_558_U21);
  nand ginst23039 (P3_ADD_558_U13, P3_INSTADDRPOINTER_REG_4__SCAN_IN, P3_ADD_558_U100);
  nand ginst23040 (P3_ADD_558_U130, P3_INSTADDRPOINTER_REG_8__SCAN_IN, P3_ADD_558_U19);
  nand ginst23041 (P3_ADD_558_U131, P3_ADD_558_U104, P3_ADD_558_U20);
  nand ginst23042 (P3_ADD_558_U132, P3_INSTADDRPOINTER_REG_7__SCAN_IN, P3_ADD_558_U17);
  nand ginst23043 (P3_ADD_558_U133, P3_ADD_558_U103, P3_ADD_558_U18);
  nand ginst23044 (P3_ADD_558_U134, P3_INSTADDRPOINTER_REG_6__SCAN_IN, P3_ADD_558_U15);
  nand ginst23045 (P3_ADD_558_U135, P3_ADD_558_U102, P3_ADD_558_U16);
  nand ginst23046 (P3_ADD_558_U136, P3_INSTADDRPOINTER_REG_5__SCAN_IN, P3_ADD_558_U13);
  nand ginst23047 (P3_ADD_558_U137, P3_ADD_558_U101, P3_ADD_558_U14);
  nand ginst23048 (P3_ADD_558_U138, P3_INSTADDRPOINTER_REG_4__SCAN_IN, P3_ADD_558_U11);
  nand ginst23049 (P3_ADD_558_U139, P3_ADD_558_U100, P3_ADD_558_U12);
  not ginst23050 (P3_ADD_558_U14, P3_INSTADDRPOINTER_REG_5__SCAN_IN);
  nand ginst23051 (P3_ADD_558_U140, P3_INSTADDRPOINTER_REG_3__SCAN_IN, P3_ADD_558_U9);
  nand ginst23052 (P3_ADD_558_U141, P3_ADD_558_U10, P3_ADD_558_U99);
  nand ginst23053 (P3_ADD_558_U142, P3_INSTADDRPOINTER_REG_31__SCAN_IN, P3_ADD_558_U97);
  nand ginst23054 (P3_ADD_558_U143, P3_ADD_558_U127, P3_ADD_558_U96);
  nand ginst23055 (P3_ADD_558_U144, P3_INSTADDRPOINTER_REG_30__SCAN_IN, P3_ADD_558_U63);
  nand ginst23056 (P3_ADD_558_U145, P3_ADD_558_U126, P3_ADD_558_U64);
  nand ginst23057 (P3_ADD_558_U146, P3_INSTADDRPOINTER_REG_2__SCAN_IN, P3_ADD_558_U7);
  nand ginst23058 (P3_ADD_558_U147, P3_ADD_558_U8, P3_ADD_558_U98);
  nand ginst23059 (P3_ADD_558_U148, P3_INSTADDRPOINTER_REG_29__SCAN_IN, P3_ADD_558_U61);
  nand ginst23060 (P3_ADD_558_U149, P3_ADD_558_U125, P3_ADD_558_U62);
  nand ginst23061 (P3_ADD_558_U15, P3_INSTADDRPOINTER_REG_5__SCAN_IN, P3_ADD_558_U101);
  nand ginst23062 (P3_ADD_558_U150, P3_INSTADDRPOINTER_REG_28__SCAN_IN, P3_ADD_558_U59);
  nand ginst23063 (P3_ADD_558_U151, P3_ADD_558_U124, P3_ADD_558_U60);
  nand ginst23064 (P3_ADD_558_U152, P3_INSTADDRPOINTER_REG_27__SCAN_IN, P3_ADD_558_U57);
  nand ginst23065 (P3_ADD_558_U153, P3_ADD_558_U123, P3_ADD_558_U58);
  nand ginst23066 (P3_ADD_558_U154, P3_INSTADDRPOINTER_REG_26__SCAN_IN, P3_ADD_558_U55);
  nand ginst23067 (P3_ADD_558_U155, P3_ADD_558_U122, P3_ADD_558_U56);
  nand ginst23068 (P3_ADD_558_U156, P3_INSTADDRPOINTER_REG_25__SCAN_IN, P3_ADD_558_U53);
  nand ginst23069 (P3_ADD_558_U157, P3_ADD_558_U121, P3_ADD_558_U54);
  nand ginst23070 (P3_ADD_558_U158, P3_INSTADDRPOINTER_REG_24__SCAN_IN, P3_ADD_558_U51);
  nand ginst23071 (P3_ADD_558_U159, P3_ADD_558_U120, P3_ADD_558_U52);
  not ginst23072 (P3_ADD_558_U16, P3_INSTADDRPOINTER_REG_6__SCAN_IN);
  nand ginst23073 (P3_ADD_558_U160, P3_INSTADDRPOINTER_REG_23__SCAN_IN, P3_ADD_558_U49);
  nand ginst23074 (P3_ADD_558_U161, P3_ADD_558_U119, P3_ADD_558_U50);
  nand ginst23075 (P3_ADD_558_U162, P3_INSTADDRPOINTER_REG_22__SCAN_IN, P3_ADD_558_U47);
  nand ginst23076 (P3_ADD_558_U163, P3_ADD_558_U118, P3_ADD_558_U48);
  nand ginst23077 (P3_ADD_558_U164, P3_INSTADDRPOINTER_REG_21__SCAN_IN, P3_ADD_558_U45);
  nand ginst23078 (P3_ADD_558_U165, P3_ADD_558_U117, P3_ADD_558_U46);
  nand ginst23079 (P3_ADD_558_U166, P3_INSTADDRPOINTER_REG_20__SCAN_IN, P3_ADD_558_U43);
  nand ginst23080 (P3_ADD_558_U167, P3_ADD_558_U116, P3_ADD_558_U44);
  nand ginst23081 (P3_ADD_558_U168, P3_INSTADDRPOINTER_REG_1__SCAN_IN, P3_ADD_558_U5);
  nand ginst23082 (P3_ADD_558_U169, P3_INSTADDRPOINTER_REG_0__SCAN_IN, P3_ADD_558_U6);
  nand ginst23083 (P3_ADD_558_U17, P3_INSTADDRPOINTER_REG_6__SCAN_IN, P3_ADD_558_U102);
  nand ginst23084 (P3_ADD_558_U170, P3_INSTADDRPOINTER_REG_19__SCAN_IN, P3_ADD_558_U41);
  nand ginst23085 (P3_ADD_558_U171, P3_ADD_558_U115, P3_ADD_558_U42);
  nand ginst23086 (P3_ADD_558_U172, P3_INSTADDRPOINTER_REG_18__SCAN_IN, P3_ADD_558_U39);
  nand ginst23087 (P3_ADD_558_U173, P3_ADD_558_U114, P3_ADD_558_U40);
  nand ginst23088 (P3_ADD_558_U174, P3_INSTADDRPOINTER_REG_17__SCAN_IN, P3_ADD_558_U37);
  nand ginst23089 (P3_ADD_558_U175, P3_ADD_558_U113, P3_ADD_558_U38);
  nand ginst23090 (P3_ADD_558_U176, P3_INSTADDRPOINTER_REG_16__SCAN_IN, P3_ADD_558_U35);
  nand ginst23091 (P3_ADD_558_U177, P3_ADD_558_U112, P3_ADD_558_U36);
  nand ginst23092 (P3_ADD_558_U178, P3_INSTADDRPOINTER_REG_15__SCAN_IN, P3_ADD_558_U33);
  nand ginst23093 (P3_ADD_558_U179, P3_ADD_558_U111, P3_ADD_558_U34);
  not ginst23094 (P3_ADD_558_U18, P3_INSTADDRPOINTER_REG_7__SCAN_IN);
  nand ginst23095 (P3_ADD_558_U180, P3_INSTADDRPOINTER_REG_14__SCAN_IN, P3_ADD_558_U31);
  nand ginst23096 (P3_ADD_558_U181, P3_ADD_558_U110, P3_ADD_558_U32);
  nand ginst23097 (P3_ADD_558_U182, P3_INSTADDRPOINTER_REG_13__SCAN_IN, P3_ADD_558_U29);
  nand ginst23098 (P3_ADD_558_U183, P3_ADD_558_U109, P3_ADD_558_U30);
  nand ginst23099 (P3_ADD_558_U184, P3_INSTADDRPOINTER_REG_12__SCAN_IN, P3_ADD_558_U27);
  nand ginst23100 (P3_ADD_558_U185, P3_ADD_558_U108, P3_ADD_558_U28);
  nand ginst23101 (P3_ADD_558_U186, P3_INSTADDRPOINTER_REG_11__SCAN_IN, P3_ADD_558_U25);
  nand ginst23102 (P3_ADD_558_U187, P3_ADD_558_U107, P3_ADD_558_U26);
  nand ginst23103 (P3_ADD_558_U188, P3_INSTADDRPOINTER_REG_10__SCAN_IN, P3_ADD_558_U23);
  nand ginst23104 (P3_ADD_558_U189, P3_ADD_558_U106, P3_ADD_558_U24);
  nand ginst23105 (P3_ADD_558_U19, P3_INSTADDRPOINTER_REG_7__SCAN_IN, P3_ADD_558_U103);
  not ginst23106 (P3_ADD_558_U20, P3_INSTADDRPOINTER_REG_8__SCAN_IN);
  not ginst23107 (P3_ADD_558_U21, P3_INSTADDRPOINTER_REG_9__SCAN_IN);
  nand ginst23108 (P3_ADD_558_U22, P3_INSTADDRPOINTER_REG_8__SCAN_IN, P3_ADD_558_U104);
  nand ginst23109 (P3_ADD_558_U23, P3_INSTADDRPOINTER_REG_9__SCAN_IN, P3_ADD_558_U105);
  not ginst23110 (P3_ADD_558_U24, P3_INSTADDRPOINTER_REG_10__SCAN_IN);
  nand ginst23111 (P3_ADD_558_U25, P3_INSTADDRPOINTER_REG_10__SCAN_IN, P3_ADD_558_U106);
  not ginst23112 (P3_ADD_558_U26, P3_INSTADDRPOINTER_REG_11__SCAN_IN);
  nand ginst23113 (P3_ADD_558_U27, P3_INSTADDRPOINTER_REG_11__SCAN_IN, P3_ADD_558_U107);
  not ginst23114 (P3_ADD_558_U28, P3_INSTADDRPOINTER_REG_12__SCAN_IN);
  nand ginst23115 (P3_ADD_558_U29, P3_INSTADDRPOINTER_REG_12__SCAN_IN, P3_ADD_558_U108);
  not ginst23116 (P3_ADD_558_U30, P3_INSTADDRPOINTER_REG_13__SCAN_IN);
  nand ginst23117 (P3_ADD_558_U31, P3_INSTADDRPOINTER_REG_13__SCAN_IN, P3_ADD_558_U109);
  not ginst23118 (P3_ADD_558_U32, P3_INSTADDRPOINTER_REG_14__SCAN_IN);
  nand ginst23119 (P3_ADD_558_U33, P3_INSTADDRPOINTER_REG_14__SCAN_IN, P3_ADD_558_U110);
  not ginst23120 (P3_ADD_558_U34, P3_INSTADDRPOINTER_REG_15__SCAN_IN);
  nand ginst23121 (P3_ADD_558_U35, P3_INSTADDRPOINTER_REG_15__SCAN_IN, P3_ADD_558_U111);
  not ginst23122 (P3_ADD_558_U36, P3_INSTADDRPOINTER_REG_16__SCAN_IN);
  nand ginst23123 (P3_ADD_558_U37, P3_INSTADDRPOINTER_REG_16__SCAN_IN, P3_ADD_558_U112);
  not ginst23124 (P3_ADD_558_U38, P3_INSTADDRPOINTER_REG_17__SCAN_IN);
  nand ginst23125 (P3_ADD_558_U39, P3_INSTADDRPOINTER_REG_17__SCAN_IN, P3_ADD_558_U113);
  not ginst23126 (P3_ADD_558_U40, P3_INSTADDRPOINTER_REG_18__SCAN_IN);
  nand ginst23127 (P3_ADD_558_U41, P3_INSTADDRPOINTER_REG_18__SCAN_IN, P3_ADD_558_U114);
  not ginst23128 (P3_ADD_558_U42, P3_INSTADDRPOINTER_REG_19__SCAN_IN);
  nand ginst23129 (P3_ADD_558_U43, P3_INSTADDRPOINTER_REG_19__SCAN_IN, P3_ADD_558_U115);
  not ginst23130 (P3_ADD_558_U44, P3_INSTADDRPOINTER_REG_20__SCAN_IN);
  nand ginst23131 (P3_ADD_558_U45, P3_INSTADDRPOINTER_REG_20__SCAN_IN, P3_ADD_558_U116);
  not ginst23132 (P3_ADD_558_U46, P3_INSTADDRPOINTER_REG_21__SCAN_IN);
  nand ginst23133 (P3_ADD_558_U47, P3_INSTADDRPOINTER_REG_21__SCAN_IN, P3_ADD_558_U117);
  not ginst23134 (P3_ADD_558_U48, P3_INSTADDRPOINTER_REG_22__SCAN_IN);
  nand ginst23135 (P3_ADD_558_U49, P3_INSTADDRPOINTER_REG_22__SCAN_IN, P3_ADD_558_U118);
  not ginst23136 (P3_ADD_558_U5, P3_INSTADDRPOINTER_REG_0__SCAN_IN);
  not ginst23137 (P3_ADD_558_U50, P3_INSTADDRPOINTER_REG_23__SCAN_IN);
  nand ginst23138 (P3_ADD_558_U51, P3_INSTADDRPOINTER_REG_23__SCAN_IN, P3_ADD_558_U119);
  not ginst23139 (P3_ADD_558_U52, P3_INSTADDRPOINTER_REG_24__SCAN_IN);
  nand ginst23140 (P3_ADD_558_U53, P3_INSTADDRPOINTER_REG_24__SCAN_IN, P3_ADD_558_U120);
  not ginst23141 (P3_ADD_558_U54, P3_INSTADDRPOINTER_REG_25__SCAN_IN);
  nand ginst23142 (P3_ADD_558_U55, P3_INSTADDRPOINTER_REG_25__SCAN_IN, P3_ADD_558_U121);
  not ginst23143 (P3_ADD_558_U56, P3_INSTADDRPOINTER_REG_26__SCAN_IN);
  nand ginst23144 (P3_ADD_558_U57, P3_INSTADDRPOINTER_REG_26__SCAN_IN, P3_ADD_558_U122);
  not ginst23145 (P3_ADD_558_U58, P3_INSTADDRPOINTER_REG_27__SCAN_IN);
  nand ginst23146 (P3_ADD_558_U59, P3_INSTADDRPOINTER_REG_27__SCAN_IN, P3_ADD_558_U123);
  not ginst23147 (P3_ADD_558_U6, P3_INSTADDRPOINTER_REG_1__SCAN_IN);
  not ginst23148 (P3_ADD_558_U60, P3_INSTADDRPOINTER_REG_28__SCAN_IN);
  nand ginst23149 (P3_ADD_558_U61, P3_INSTADDRPOINTER_REG_28__SCAN_IN, P3_ADD_558_U124);
  not ginst23150 (P3_ADD_558_U62, P3_INSTADDRPOINTER_REG_29__SCAN_IN);
  nand ginst23151 (P3_ADD_558_U63, P3_INSTADDRPOINTER_REG_29__SCAN_IN, P3_ADD_558_U125);
  not ginst23152 (P3_ADD_558_U64, P3_INSTADDRPOINTER_REG_30__SCAN_IN);
  nand ginst23153 (P3_ADD_558_U65, P3_ADD_558_U128, P3_ADD_558_U129);
  nand ginst23154 (P3_ADD_558_U66, P3_ADD_558_U130, P3_ADD_558_U131);
  nand ginst23155 (P3_ADD_558_U67, P3_ADD_558_U132, P3_ADD_558_U133);
  nand ginst23156 (P3_ADD_558_U68, P3_ADD_558_U134, P3_ADD_558_U135);
  nand ginst23157 (P3_ADD_558_U69, P3_ADD_558_U136, P3_ADD_558_U137);
  nand ginst23158 (P3_ADD_558_U7, P3_INSTADDRPOINTER_REG_0__SCAN_IN, P3_INSTADDRPOINTER_REG_1__SCAN_IN);
  nand ginst23159 (P3_ADD_558_U70, P3_ADD_558_U138, P3_ADD_558_U139);
  nand ginst23160 (P3_ADD_558_U71, P3_ADD_558_U140, P3_ADD_558_U141);
  nand ginst23161 (P3_ADD_558_U72, P3_ADD_558_U142, P3_ADD_558_U143);
  nand ginst23162 (P3_ADD_558_U73, P3_ADD_558_U144, P3_ADD_558_U145);
  nand ginst23163 (P3_ADD_558_U74, P3_ADD_558_U146, P3_ADD_558_U147);
  nand ginst23164 (P3_ADD_558_U75, P3_ADD_558_U148, P3_ADD_558_U149);
  nand ginst23165 (P3_ADD_558_U76, P3_ADD_558_U150, P3_ADD_558_U151);
  nand ginst23166 (P3_ADD_558_U77, P3_ADD_558_U152, P3_ADD_558_U153);
  nand ginst23167 (P3_ADD_558_U78, P3_ADD_558_U154, P3_ADD_558_U155);
  nand ginst23168 (P3_ADD_558_U79, P3_ADD_558_U156, P3_ADD_558_U157);
  not ginst23169 (P3_ADD_558_U8, P3_INSTADDRPOINTER_REG_2__SCAN_IN);
  nand ginst23170 (P3_ADD_558_U80, P3_ADD_558_U158, P3_ADD_558_U159);
  nand ginst23171 (P3_ADD_558_U81, P3_ADD_558_U160, P3_ADD_558_U161);
  nand ginst23172 (P3_ADD_558_U82, P3_ADD_558_U162, P3_ADD_558_U163);
  nand ginst23173 (P3_ADD_558_U83, P3_ADD_558_U164, P3_ADD_558_U165);
  nand ginst23174 (P3_ADD_558_U84, P3_ADD_558_U166, P3_ADD_558_U167);
  nand ginst23175 (P3_ADD_558_U85, P3_ADD_558_U168, P3_ADD_558_U169);
  nand ginst23176 (P3_ADD_558_U86, P3_ADD_558_U170, P3_ADD_558_U171);
  nand ginst23177 (P3_ADD_558_U87, P3_ADD_558_U172, P3_ADD_558_U173);
  nand ginst23178 (P3_ADD_558_U88, P3_ADD_558_U174, P3_ADD_558_U175);
  nand ginst23179 (P3_ADD_558_U89, P3_ADD_558_U176, P3_ADD_558_U177);
  nand ginst23180 (P3_ADD_558_U9, P3_INSTADDRPOINTER_REG_2__SCAN_IN, P3_ADD_558_U98);
  nand ginst23181 (P3_ADD_558_U90, P3_ADD_558_U178, P3_ADD_558_U179);
  nand ginst23182 (P3_ADD_558_U91, P3_ADD_558_U180, P3_ADD_558_U181);
  nand ginst23183 (P3_ADD_558_U92, P3_ADD_558_U182, P3_ADD_558_U183);
  nand ginst23184 (P3_ADD_558_U93, P3_ADD_558_U184, P3_ADD_558_U185);
  nand ginst23185 (P3_ADD_558_U94, P3_ADD_558_U186, P3_ADD_558_U187);
  nand ginst23186 (P3_ADD_558_U95, P3_ADD_558_U188, P3_ADD_558_U189);
  not ginst23187 (P3_ADD_558_U96, P3_INSTADDRPOINTER_REG_31__SCAN_IN);
  nand ginst23188 (P3_ADD_558_U97, P3_INSTADDRPOINTER_REG_30__SCAN_IN, P3_ADD_558_U126);
  not ginst23189 (P3_ADD_558_U98, P3_ADD_558_U7);
  not ginst23190 (P3_ADD_558_U99, P3_ADD_558_U9);
  nor ginst23191 (P3_GTE_355_U6, P3_GTE_355_U8, P3_SUB_355_U6);
  and ginst23192 (P3_GTE_355_U7, P3_SUB_355_U22, P3_SUB_355_U7);
  nor ginst23193 (P3_GTE_355_U8, P3_GTE_355_U7, P3_SUB_355_U19, P3_SUB_355_U20, P3_SUB_355_U21);
  nor ginst23194 (P3_GTE_370_U6, P3_GTE_370_U8, P3_SUB_370_U6);
  and ginst23195 (P3_GTE_370_U7, P3_GTE_370_U9, P3_SUB_370_U21);
  nor ginst23196 (P3_GTE_370_U8, P3_GTE_370_U7, P3_SUB_370_U19, P3_SUB_370_U20);
  or ginst23197 (P3_GTE_370_U9, P3_SUB_370_U22, P3_SUB_370_U7);
  nor ginst23198 (P3_GTE_390_U6, P3_GTE_390_U8, P3_SUB_390_U6);
  and ginst23199 (P3_GTE_390_U7, P3_GTE_390_U9, P3_SUB_390_U21);
  nor ginst23200 (P3_GTE_390_U8, P3_GTE_390_U7, P3_SUB_390_U19, P3_SUB_390_U20);
  or ginst23201 (P3_GTE_390_U9, P3_SUB_390_U22, P3_SUB_390_U7);
  nor ginst23202 (P3_GTE_401_U6, P3_GTE_401_U8, P3_SUB_401_U6);
  and ginst23203 (P3_GTE_401_U7, P3_GTE_401_U9, P3_SUB_401_U21);
  nor ginst23204 (P3_GTE_401_U8, P3_GTE_401_U7, P3_SUB_401_U19, P3_SUB_401_U20);
  or ginst23205 (P3_GTE_401_U9, P3_SUB_401_U22, P3_SUB_401_U7);
  nor ginst23206 (P3_GTE_412_U6, P3_GTE_412_U7, P3_SUB_412_U6);
  nor ginst23207 (P3_GTE_412_U7, P3_SUB_412_U16, P3_SUB_412_U17, P3_SUB_412_U18, P3_SUB_412_U19);
  nor ginst23208 (P3_GTE_450_U6, P3_GTE_450_U7, P3_SUB_450_U6);
  nor ginst23209 (P3_GTE_450_U7, P3_SUB_450_U16, P3_SUB_450_U17, P3_SUB_450_U18, P3_SUB_450_U19);
  nor ginst23210 (P3_GTE_485_U6, P3_GTE_485_U7, P3_SUB_485_U6);
  nor ginst23211 (P3_GTE_485_U7, P3_SUB_485_U16, P3_SUB_485_U17, P3_SUB_485_U18, P3_SUB_485_U19);
  nor ginst23212 (P3_GTE_504_U6, P3_GTE_504_U7, P3_SUB_504_U6);
  nor ginst23213 (P3_GTE_504_U7, P3_SUB_504_U16, P3_SUB_504_U17, P3_SUB_504_U18, P3_SUB_504_U19);
  not ginst23214 (P3_LTE_597_U6, P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN);
  or ginst23215 (P3_LT_563_1260_U6, P3_LT_563_1260_U7, P3_U3304);
  nor ginst23216 (P3_LT_563_1260_U7, P3_SUB_563_U6, P3_SUB_563_U7);
  not ginst23217 (P3_LT_563_U10, P3_U3306);
  not ginst23218 (P3_LT_563_U11, P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN);
  not ginst23219 (P3_LT_563_U12, P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN);
  not ginst23220 (P3_LT_563_U13, P3_U3305);
  not ginst23221 (P3_LT_563_U14, P3_U3304);
  not ginst23222 (P3_LT_563_U15, P3_U3308);
  not ginst23223 (P3_LT_563_U16, P3_LT_563_U8);
  nand ginst23224 (P3_LT_563_U17, P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN, P3_LT_563_U16);
  nand ginst23225 (P3_LT_563_U18, P3_LT_563_U17, P3_U3307);
  nand ginst23226 (P3_LT_563_U19, P3_LT_563_U8, P3_LT_563_U9);
  nand ginst23227 (P3_LT_563_U20, P3_LT_563_U11, P3_U3306);
  nand ginst23228 (P3_LT_563_U21, P3_LT_563_U18, P3_LT_563_U19, P3_LT_563_U20);
  nand ginst23229 (P3_LT_563_U22, P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN, P3_LT_563_U10);
  nand ginst23230 (P3_LT_563_U23, P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN, P3_LT_563_U13);
  nand ginst23231 (P3_LT_563_U24, P3_LT_563_U21, P3_LT_563_U22, P3_LT_563_U23);
  nand ginst23232 (P3_LT_563_U25, P3_LT_563_U12, P3_U3305);
  nand ginst23233 (P3_LT_563_U26, P3_LT_563_U7, P3_U3304);
  nand ginst23234 (P3_LT_563_U27, P3_LT_563_U24, P3_LT_563_U25, P3_LT_563_U26);
  nand ginst23235 (P3_LT_563_U28, P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN, P3_LT_563_U14);
  nand ginst23236 (P3_LT_563_U6, P3_LT_563_U27, P3_LT_563_U28);
  not ginst23237 (P3_LT_563_U7, P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN);
  nand ginst23238 (P3_LT_563_U8, P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P3_LT_563_U15);
  not ginst23239 (P3_LT_563_U9, P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN);
  or ginst23240 (P3_LT_589_U6, P3_LT_589_U8, P3_U2629);
  and ginst23241 (P3_LT_589_U7, P3_SUB_589_U6, P3_SUB_589_U7);
  nor ginst23242 (P3_LT_589_U8, P3_LT_589_U7, P3_SUB_589_U8, P3_SUB_589_U9);
  and ginst23243 (P3_SUB_320_U10, P3_SUB_320_U118, P3_SUB_320_U32);
  not ginst23244 (P3_SUB_320_U100, P3_SUB_320_U35);
  not ginst23245 (P3_SUB_320_U101, P3_SUB_320_U36);
  not ginst23246 (P3_SUB_320_U102, P3_SUB_320_U37);
  not ginst23247 (P3_SUB_320_U103, P3_SUB_320_U38);
  or ginst23248 (P3_SUB_320_U104, P3_PHYADDRPOINTER_REG_0__SCAN_IN, P3_ADD_318_U4);
  nand ginst23249 (P3_SUB_320_U105, P3_ADD_318_U71, P3_SUB_320_U104);
  nand ginst23250 (P3_SUB_320_U106, P3_ADD_318_U72, P3_SUB_320_U37);
  nand ginst23251 (P3_SUB_320_U107, P3_SUB_320_U101, P3_SUB_320_U63);
  nand ginst23252 (P3_SUB_320_U108, P3_ADD_318_U73, P3_SUB_320_U107);
  nand ginst23253 (P3_SUB_320_U109, P3_SUB_320_U100, P3_SUB_320_U65);
  and ginst23254 (P3_SUB_320_U11, P3_SUB_320_U116, P3_SUB_320_U33);
  nand ginst23255 (P3_SUB_320_U110, P3_ADD_318_U75, P3_SUB_320_U109);
  nand ginst23256 (P3_SUB_320_U111, P3_SUB_320_U67, P3_SUB_320_U99);
  nand ginst23257 (P3_SUB_320_U112, P3_ADD_318_U77, P3_SUB_320_U111);
  nand ginst23258 (P3_SUB_320_U113, P3_SUB_320_U69, P3_SUB_320_U98);
  nand ginst23259 (P3_SUB_320_U114, P3_ADD_318_U79, P3_SUB_320_U113);
  nand ginst23260 (P3_SUB_320_U115, P3_SUB_320_U73, P3_SUB_320_U97);
  nand ginst23261 (P3_SUB_320_U116, P3_ADD_318_U81, P3_SUB_320_U115);
  nand ginst23262 (P3_SUB_320_U117, P3_SUB_320_U75, P3_SUB_320_U96);
  nand ginst23263 (P3_SUB_320_U118, P3_ADD_318_U83, P3_SUB_320_U117);
  nand ginst23264 (P3_SUB_320_U119, P3_SUB_320_U77, P3_SUB_320_U95);
  and ginst23265 (P3_SUB_320_U12, P3_SUB_320_U114, P3_SUB_320_U34);
  nand ginst23266 (P3_SUB_320_U120, P3_ADD_318_U85, P3_SUB_320_U119);
  nand ginst23267 (P3_SUB_320_U121, P3_SUB_320_U79, P3_SUB_320_U94);
  nand ginst23268 (P3_SUB_320_U122, P3_ADD_318_U87, P3_SUB_320_U121);
  nand ginst23269 (P3_SUB_320_U123, P3_SUB_320_U81, P3_SUB_320_U93);
  nand ginst23270 (P3_SUB_320_U124, P3_ADD_318_U89, P3_SUB_320_U123);
  nand ginst23271 (P3_SUB_320_U125, P3_SUB_320_U52, P3_SUB_320_U86);
  nand ginst23272 (P3_SUB_320_U126, P3_ADD_318_U91, P3_SUB_320_U125);
  nand ginst23273 (P3_SUB_320_U127, P3_SUB_320_U103, P3_SUB_320_U61);
  nand ginst23274 (P3_SUB_320_U128, P3_ADD_318_U62, P3_SUB_320_U24);
  nand ginst23275 (P3_SUB_320_U129, P3_SUB_320_U52, P3_SUB_320_U86);
  and ginst23276 (P3_SUB_320_U13, P3_SUB_320_U112, P3_SUB_320_U35);
  nand ginst23277 (P3_SUB_320_U130, P3_ADD_318_U64, P3_SUB_320_U23);
  nand ginst23278 (P3_SUB_320_U131, P3_SUB_320_U54, P3_SUB_320_U85);
  nand ginst23279 (P3_SUB_320_U132, P3_ADD_318_U66, P3_SUB_320_U22);
  nand ginst23280 (P3_SUB_320_U133, P3_SUB_320_U56, P3_SUB_320_U84);
  nand ginst23281 (P3_SUB_320_U134, P3_ADD_318_U68, P3_SUB_320_U21);
  nand ginst23282 (P3_SUB_320_U135, P3_SUB_320_U58, P3_SUB_320_U83);
  nand ginst23283 (P3_SUB_320_U136, P3_SUB_320_U127, P3_SUB_320_U60);
  nand ginst23284 (P3_SUB_320_U137, P3_ADD_318_U69, P3_SUB_320_U103, P3_SUB_320_U61);
  nand ginst23285 (P3_SUB_320_U138, P3_ADD_318_U70, P3_SUB_320_U38);
  nand ginst23286 (P3_SUB_320_U139, P3_SUB_320_U103, P3_SUB_320_U61);
  and ginst23287 (P3_SUB_320_U14, P3_SUB_320_U110, P3_SUB_320_U36);
  nand ginst23288 (P3_SUB_320_U140, P3_ADD_318_U74, P3_SUB_320_U36);
  nand ginst23289 (P3_SUB_320_U141, P3_SUB_320_U101, P3_SUB_320_U63);
  nand ginst23290 (P3_SUB_320_U142, P3_ADD_318_U76, P3_SUB_320_U35);
  nand ginst23291 (P3_SUB_320_U143, P3_SUB_320_U100, P3_SUB_320_U65);
  nand ginst23292 (P3_SUB_320_U144, P3_ADD_318_U78, P3_SUB_320_U34);
  nand ginst23293 (P3_SUB_320_U145, P3_SUB_320_U67, P3_SUB_320_U99);
  nand ginst23294 (P3_SUB_320_U146, P3_ADD_318_U80, P3_SUB_320_U33);
  nand ginst23295 (P3_SUB_320_U147, P3_SUB_320_U69, P3_SUB_320_U98);
  nand ginst23296 (P3_SUB_320_U148, P3_ADD_318_U4, P3_SUB_320_U72);
  nand ginst23297 (P3_SUB_320_U149, P3_PHYADDRPOINTER_REG_0__SCAN_IN, P3_SUB_320_U71);
  and ginst23298 (P3_SUB_320_U15, P3_SUB_320_U108, P3_SUB_320_U37);
  nand ginst23299 (P3_SUB_320_U150, P3_ADD_318_U82, P3_SUB_320_U32);
  nand ginst23300 (P3_SUB_320_U151, P3_SUB_320_U73, P3_SUB_320_U97);
  nand ginst23301 (P3_SUB_320_U152, P3_ADD_318_U84, P3_SUB_320_U31);
  nand ginst23302 (P3_SUB_320_U153, P3_SUB_320_U75, P3_SUB_320_U96);
  nand ginst23303 (P3_SUB_320_U154, P3_ADD_318_U86, P3_SUB_320_U30);
  nand ginst23304 (P3_SUB_320_U155, P3_SUB_320_U77, P3_SUB_320_U95);
  nand ginst23305 (P3_SUB_320_U156, P3_ADD_318_U88, P3_SUB_320_U29);
  nand ginst23306 (P3_SUB_320_U157, P3_SUB_320_U79, P3_SUB_320_U94);
  nand ginst23307 (P3_SUB_320_U158, P3_ADD_318_U90, P3_SUB_320_U28);
  nand ginst23308 (P3_SUB_320_U159, P3_SUB_320_U81, P3_SUB_320_U93);
  and ginst23309 (P3_SUB_320_U16, P3_SUB_320_U106, P3_SUB_320_U38);
  and ginst23310 (P3_SUB_320_U17, P3_SUB_320_U105, P3_SUB_320_U21);
  and ginst23311 (P3_SUB_320_U18, P3_SUB_320_U22, P3_SUB_320_U92);
  and ginst23312 (P3_SUB_320_U19, P3_SUB_320_U23, P3_SUB_320_U90);
  and ginst23313 (P3_SUB_320_U20, P3_SUB_320_U24, P3_SUB_320_U88);
  or ginst23314 (P3_SUB_320_U21, P3_PHYADDRPOINTER_REG_0__SCAN_IN, P3_ADD_318_U4, P3_ADD_318_U71);
  nand ginst23315 (P3_SUB_320_U22, P3_SUB_320_U27, P3_SUB_320_U58, P3_SUB_320_U83);
  nand ginst23316 (P3_SUB_320_U23, P3_SUB_320_U26, P3_SUB_320_U56, P3_SUB_320_U84);
  nand ginst23317 (P3_SUB_320_U24, P3_SUB_320_U25, P3_SUB_320_U54, P3_SUB_320_U85);
  not ginst23318 (P3_SUB_320_U25, P3_ADD_318_U63);
  not ginst23319 (P3_SUB_320_U26, P3_ADD_318_U65);
  not ginst23320 (P3_SUB_320_U27, P3_ADD_318_U67);
  nand ginst23321 (P3_SUB_320_U28, P3_SUB_320_U49, P3_SUB_320_U52, P3_SUB_320_U86);
  nand ginst23322 (P3_SUB_320_U29, P3_SUB_320_U48, P3_SUB_320_U81, P3_SUB_320_U93);
  nand ginst23323 (P3_SUB_320_U30, P3_SUB_320_U47, P3_SUB_320_U79, P3_SUB_320_U94);
  nand ginst23324 (P3_SUB_320_U31, P3_SUB_320_U46, P3_SUB_320_U77, P3_SUB_320_U95);
  nand ginst23325 (P3_SUB_320_U32, P3_SUB_320_U45, P3_SUB_320_U75, P3_SUB_320_U96);
  nand ginst23326 (P3_SUB_320_U33, P3_SUB_320_U44, P3_SUB_320_U73, P3_SUB_320_U97);
  nand ginst23327 (P3_SUB_320_U34, P3_SUB_320_U43, P3_SUB_320_U69, P3_SUB_320_U98);
  nand ginst23328 (P3_SUB_320_U35, P3_SUB_320_U42, P3_SUB_320_U67, P3_SUB_320_U99);
  nand ginst23329 (P3_SUB_320_U36, P3_SUB_320_U100, P3_SUB_320_U41, P3_SUB_320_U65);
  nand ginst23330 (P3_SUB_320_U37, P3_SUB_320_U101, P3_SUB_320_U40, P3_SUB_320_U63);
  nand ginst23331 (P3_SUB_320_U38, P3_SUB_320_U102, P3_SUB_320_U39);
  not ginst23332 (P3_SUB_320_U39, P3_ADD_318_U72);
  not ginst23333 (P3_SUB_320_U40, P3_ADD_318_U73);
  not ginst23334 (P3_SUB_320_U41, P3_ADD_318_U75);
  not ginst23335 (P3_SUB_320_U42, P3_ADD_318_U77);
  not ginst23336 (P3_SUB_320_U43, P3_ADD_318_U79);
  not ginst23337 (P3_SUB_320_U44, P3_ADD_318_U81);
  not ginst23338 (P3_SUB_320_U45, P3_ADD_318_U83);
  not ginst23339 (P3_SUB_320_U46, P3_ADD_318_U85);
  not ginst23340 (P3_SUB_320_U47, P3_ADD_318_U87);
  not ginst23341 (P3_SUB_320_U48, P3_ADD_318_U89);
  not ginst23342 (P3_SUB_320_U49, P3_ADD_318_U91);
  nand ginst23343 (P3_SUB_320_U50, P3_SUB_320_U148, P3_SUB_320_U149);
  nand ginst23344 (P3_SUB_320_U51, P3_SUB_320_U136, P3_SUB_320_U137);
  not ginst23345 (P3_SUB_320_U52, P3_ADD_318_U62);
  and ginst23346 (P3_SUB_320_U53, P3_SUB_320_U128, P3_SUB_320_U129);
  not ginst23347 (P3_SUB_320_U54, P3_ADD_318_U64);
  and ginst23348 (P3_SUB_320_U55, P3_SUB_320_U130, P3_SUB_320_U131);
  not ginst23349 (P3_SUB_320_U56, P3_ADD_318_U66);
  and ginst23350 (P3_SUB_320_U57, P3_SUB_320_U132, P3_SUB_320_U133);
  not ginst23351 (P3_SUB_320_U58, P3_ADD_318_U68);
  and ginst23352 (P3_SUB_320_U59, P3_SUB_320_U134, P3_SUB_320_U135);
  and ginst23353 (P3_SUB_320_U6, P3_SUB_320_U126, P3_SUB_320_U28);
  not ginst23354 (P3_SUB_320_U60, P3_ADD_318_U69);
  not ginst23355 (P3_SUB_320_U61, P3_ADD_318_U70);
  and ginst23356 (P3_SUB_320_U62, P3_SUB_320_U138, P3_SUB_320_U139);
  not ginst23357 (P3_SUB_320_U63, P3_ADD_318_U74);
  and ginst23358 (P3_SUB_320_U64, P3_SUB_320_U140, P3_SUB_320_U141);
  not ginst23359 (P3_SUB_320_U65, P3_ADD_318_U76);
  and ginst23360 (P3_SUB_320_U66, P3_SUB_320_U142, P3_SUB_320_U143);
  not ginst23361 (P3_SUB_320_U67, P3_ADD_318_U78);
  and ginst23362 (P3_SUB_320_U68, P3_SUB_320_U144, P3_SUB_320_U145);
  not ginst23363 (P3_SUB_320_U69, P3_ADD_318_U80);
  and ginst23364 (P3_SUB_320_U7, P3_SUB_320_U124, P3_SUB_320_U29);
  and ginst23365 (P3_SUB_320_U70, P3_SUB_320_U146, P3_SUB_320_U147);
  not ginst23366 (P3_SUB_320_U71, P3_ADD_318_U4);
  not ginst23367 (P3_SUB_320_U72, P3_PHYADDRPOINTER_REG_0__SCAN_IN);
  not ginst23368 (P3_SUB_320_U73, P3_ADD_318_U82);
  and ginst23369 (P3_SUB_320_U74, P3_SUB_320_U150, P3_SUB_320_U151);
  not ginst23370 (P3_SUB_320_U75, P3_ADD_318_U84);
  and ginst23371 (P3_SUB_320_U76, P3_SUB_320_U152, P3_SUB_320_U153);
  not ginst23372 (P3_SUB_320_U77, P3_ADD_318_U86);
  and ginst23373 (P3_SUB_320_U78, P3_SUB_320_U154, P3_SUB_320_U155);
  not ginst23374 (P3_SUB_320_U79, P3_ADD_318_U88);
  and ginst23375 (P3_SUB_320_U8, P3_SUB_320_U122, P3_SUB_320_U30);
  and ginst23376 (P3_SUB_320_U80, P3_SUB_320_U156, P3_SUB_320_U157);
  not ginst23377 (P3_SUB_320_U81, P3_ADD_318_U90);
  and ginst23378 (P3_SUB_320_U82, P3_SUB_320_U158, P3_SUB_320_U159);
  not ginst23379 (P3_SUB_320_U83, P3_SUB_320_U21);
  not ginst23380 (P3_SUB_320_U84, P3_SUB_320_U22);
  not ginst23381 (P3_SUB_320_U85, P3_SUB_320_U23);
  not ginst23382 (P3_SUB_320_U86, P3_SUB_320_U24);
  nand ginst23383 (P3_SUB_320_U87, P3_SUB_320_U54, P3_SUB_320_U85);
  nand ginst23384 (P3_SUB_320_U88, P3_ADD_318_U63, P3_SUB_320_U87);
  nand ginst23385 (P3_SUB_320_U89, P3_SUB_320_U56, P3_SUB_320_U84);
  and ginst23386 (P3_SUB_320_U9, P3_SUB_320_U120, P3_SUB_320_U31);
  nand ginst23387 (P3_SUB_320_U90, P3_ADD_318_U65, P3_SUB_320_U89);
  nand ginst23388 (P3_SUB_320_U91, P3_SUB_320_U58, P3_SUB_320_U83);
  nand ginst23389 (P3_SUB_320_U92, P3_ADD_318_U67, P3_SUB_320_U91);
  not ginst23390 (P3_SUB_320_U93, P3_SUB_320_U28);
  not ginst23391 (P3_SUB_320_U94, P3_SUB_320_U29);
  not ginst23392 (P3_SUB_320_U95, P3_SUB_320_U30);
  not ginst23393 (P3_SUB_320_U96, P3_SUB_320_U31);
  not ginst23394 (P3_SUB_320_U97, P3_SUB_320_U32);
  not ginst23395 (P3_SUB_320_U98, P3_SUB_320_U33);
  not ginst23396 (P3_SUB_320_U99, P3_SUB_320_U34);
  not ginst23397 (P3_SUB_355_U10, P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN);
  not ginst23398 (P3_SUB_355_U11, P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN);
  not ginst23399 (P3_SUB_355_U12, P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN);
  not ginst23400 (P3_SUB_355_U13, P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN);
  not ginst23401 (P3_SUB_355_U14, P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN);
  not ginst23402 (P3_SUB_355_U15, P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN);
  nand ginst23403 (P3_SUB_355_U16, P3_SUB_355_U40, P3_SUB_355_U41);
  not ginst23404 (P3_SUB_355_U17, P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN);
  not ginst23405 (P3_SUB_355_U18, P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN);
  nand ginst23406 (P3_SUB_355_U19, P3_SUB_355_U50, P3_SUB_355_U51);
  nand ginst23407 (P3_SUB_355_U20, P3_SUB_355_U55, P3_SUB_355_U56);
  nand ginst23408 (P3_SUB_355_U21, P3_SUB_355_U60, P3_SUB_355_U61);
  nand ginst23409 (P3_SUB_355_U22, P3_SUB_355_U65, P3_SUB_355_U66);
  nand ginst23410 (P3_SUB_355_U23, P3_SUB_355_U47, P3_SUB_355_U48);
  nand ginst23411 (P3_SUB_355_U24, P3_SUB_355_U52, P3_SUB_355_U53);
  nand ginst23412 (P3_SUB_355_U25, P3_SUB_355_U57, P3_SUB_355_U58);
  nand ginst23413 (P3_SUB_355_U26, P3_SUB_355_U62, P3_SUB_355_U63);
  nand ginst23414 (P3_SUB_355_U27, P3_SUB_355_U36, P3_SUB_355_U37);
  nand ginst23415 (P3_SUB_355_U28, P3_SUB_355_U32, P3_SUB_355_U33);
  not ginst23416 (P3_SUB_355_U29, P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN);
  not ginst23417 (P3_SUB_355_U30, P3_SUB_355_U9);
  nand ginst23418 (P3_SUB_355_U31, P3_SUB_355_U10, P3_SUB_355_U30);
  nand ginst23419 (P3_SUB_355_U32, P3_SUB_355_U29, P3_SUB_355_U31);
  nand ginst23420 (P3_SUB_355_U33, P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN, P3_SUB_355_U9);
  not ginst23421 (P3_SUB_355_U34, P3_SUB_355_U28);
  nand ginst23422 (P3_SUB_355_U35, P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN, P3_SUB_355_U12);
  nand ginst23423 (P3_SUB_355_U36, P3_SUB_355_U28, P3_SUB_355_U35);
  nand ginst23424 (P3_SUB_355_U37, P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN, P3_SUB_355_U11);
  not ginst23425 (P3_SUB_355_U38, P3_SUB_355_U27);
  nand ginst23426 (P3_SUB_355_U39, P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P3_SUB_355_U14);
  nand ginst23427 (P3_SUB_355_U40, P3_SUB_355_U27, P3_SUB_355_U39);
  nand ginst23428 (P3_SUB_355_U41, P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN, P3_SUB_355_U13);
  not ginst23429 (P3_SUB_355_U42, P3_SUB_355_U16);
  nand ginst23430 (P3_SUB_355_U43, P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN, P3_SUB_355_U17);
  nand ginst23431 (P3_SUB_355_U44, P3_SUB_355_U42, P3_SUB_355_U43);
  nand ginst23432 (P3_SUB_355_U45, P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN, P3_SUB_355_U15);
  nand ginst23433 (P3_SUB_355_U46, P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P3_SUB_355_U8);
  nand ginst23434 (P3_SUB_355_U47, P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN, P3_SUB_355_U15);
  nand ginst23435 (P3_SUB_355_U48, P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN, P3_SUB_355_U17);
  not ginst23436 (P3_SUB_355_U49, P3_SUB_355_U23);
  nand ginst23437 (P3_SUB_355_U50, P3_SUB_355_U42, P3_SUB_355_U49);
  nand ginst23438 (P3_SUB_355_U51, P3_SUB_355_U16, P3_SUB_355_U23);
  nand ginst23439 (P3_SUB_355_U52, P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P3_SUB_355_U14);
  nand ginst23440 (P3_SUB_355_U53, P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN, P3_SUB_355_U13);
  not ginst23441 (P3_SUB_355_U54, P3_SUB_355_U24);
  nand ginst23442 (P3_SUB_355_U55, P3_SUB_355_U38, P3_SUB_355_U54);
  nand ginst23443 (P3_SUB_355_U56, P3_SUB_355_U24, P3_SUB_355_U27);
  nand ginst23444 (P3_SUB_355_U57, P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN, P3_SUB_355_U12);
  nand ginst23445 (P3_SUB_355_U58, P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN, P3_SUB_355_U11);
  not ginst23446 (P3_SUB_355_U59, P3_SUB_355_U25);
  nand ginst23447 (P3_SUB_355_U6, P3_SUB_355_U44, P3_SUB_355_U45);
  nand ginst23448 (P3_SUB_355_U60, P3_SUB_355_U34, P3_SUB_355_U59);
  nand ginst23449 (P3_SUB_355_U61, P3_SUB_355_U25, P3_SUB_355_U28);
  nand ginst23450 (P3_SUB_355_U62, P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P3_SUB_355_U10);
  nand ginst23451 (P3_SUB_355_U63, P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN, P3_SUB_355_U29);
  not ginst23452 (P3_SUB_355_U64, P3_SUB_355_U26);
  nand ginst23453 (P3_SUB_355_U65, P3_SUB_355_U30, P3_SUB_355_U64);
  nand ginst23454 (P3_SUB_355_U66, P3_SUB_355_U26, P3_SUB_355_U9);
  nand ginst23455 (P3_SUB_355_U7, P3_SUB_355_U46, P3_SUB_355_U9);
  not ginst23456 (P3_SUB_355_U8, P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN);
  nand ginst23457 (P3_SUB_355_U9, P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN, P3_SUB_355_U18);
  and ginst23458 (P3_SUB_357_1258_U10, P3_SUB_357_1258_U156, P3_SUB_357_1258_U205, P3_SUB_357_1258_U206, P3_SUB_357_1258_U210);
  and ginst23459 (P3_SUB_357_1258_U100, P3_SUB_357_1258_U8, P3_SUB_357_1258_U99);
  and ginst23460 (P3_SUB_357_1258_U101, P3_INSTADDRPOINTER_REG_16__SCAN_IN, P3_INSTADDRPOINTER_REG_17__SCAN_IN);
  and ginst23461 (P3_SUB_357_1258_U102, P3_SUB_357_1258_U199, P3_SUB_357_1258_U56);
  and ginst23462 (P3_SUB_357_1258_U103, P3_SUB_357_1258_U13, P3_SUB_357_1258_U215);
  and ginst23463 (P3_SUB_357_1258_U104, P3_SUB_357_1258_U14, P3_SUB_357_1258_U216);
  and ginst23464 (P3_SUB_357_1258_U105, P3_SUB_357_1258_U157, P3_SUB_357_1258_U219, P3_SUB_357_1258_U58);
  and ginst23465 (P3_SUB_357_1258_U106, P3_SUB_357_1258_U157, P3_SUB_357_1258_U219);
  and ginst23466 (P3_SUB_357_1258_U107, P3_INSTADDRPOINTER_REG_31__SCAN_IN, P3_SUB_357_1258_U269, P3_SUB_357_1258_U60);
  and ginst23467 (P3_SUB_357_1258_U108, P3_INSTADDRPOINTER_REG_30__SCAN_IN, P3_INSTADDRPOINTER_REG_31__SCAN_IN);
  and ginst23468 (P3_SUB_357_1258_U109, P3_SUB_357_1258_U157, P3_SUB_357_1258_U385, P3_SUB_357_1258_U386);
  and ginst23469 (P3_SUB_357_1258_U11, P3_SUB_357_1258_U211, P3_SUB_357_1258_U9);
  and ginst23470 (P3_SUB_357_1258_U110, P3_SUB_357_1258_U153, P3_SUB_357_1258_U232);
  and ginst23471 (P3_SUB_357_1258_U111, P3_SUB_357_1258_U156, P3_SUB_357_1258_U237);
  and ginst23472 (P3_SUB_357_1258_U112, P3_SUB_357_1258_U156, P3_SUB_357_1258_U243);
  and ginst23473 (P3_SUB_357_1258_U113, P3_SUB_357_1258_U155, P3_SUB_357_1258_U464, P3_SUB_357_1258_U465);
  and ginst23474 (P3_SUB_357_1258_U114, P3_SUB_357_1258_U154, P3_SUB_357_1258_U254);
  nand ginst23475 (P3_SUB_357_1258_U115, P3_SUB_357_1258_U152, P3_SUB_357_1258_U176, P3_SUB_357_1258_U268);
  and ginst23476 (P3_SUB_357_1258_U116, P3_SUB_357_1258_U313, P3_SUB_357_1258_U314);
  nand ginst23477 (P3_SUB_357_1258_U117, P3_SUB_357_1258_U267, P3_SUB_357_1258_U300);
  and ginst23478 (P3_SUB_357_1258_U118, P3_SUB_357_1258_U320, P3_SUB_357_1258_U321);
  nand ginst23479 (P3_SUB_357_1258_U119, P3_SUB_357_1258_U172, P3_SUB_357_1258_U173);
  and ginst23480 (P3_SUB_357_1258_U12, P3_SUB_357_1258_U10, P3_SUB_357_1258_U212);
  and ginst23481 (P3_SUB_357_1258_U120, P3_SUB_357_1258_U327, P3_SUB_357_1258_U328);
  nand ginst23482 (P3_SUB_357_1258_U121, P3_SUB_357_1258_U266, P3_SUB_357_1258_U298);
  and ginst23483 (P3_SUB_357_1258_U122, P3_SUB_357_1258_U334, P3_SUB_357_1258_U335);
  nand ginst23484 (P3_SUB_357_1258_U123, P3_SUB_357_1258_U167, P3_SUB_357_1258_U96);
  nand ginst23485 (P3_SUB_357_1258_U124, P3_SUB_357_1258_U180, P3_SUB_357_1258_U181);
  nand ginst23486 (P3_SUB_357_1258_U125, P3_SUB_357_1258_U159, P3_SUB_357_1258_U183);
  and ginst23487 (P3_SUB_357_1258_U126, P3_SUB_357_1258_U355, P3_SUB_357_1258_U356);
  nand ginst23488 (P3_SUB_357_1258_U127, P3_SUB_357_1258_U270, P3_SUB_357_1258_U271, P3_SUB_357_1258_U66);
  and ginst23489 (P3_SUB_357_1258_U128, P3_SUB_357_1258_U367, P3_SUB_357_1258_U368);
  nand ginst23490 (P3_SUB_357_1258_U129, P3_SUB_357_1258_U274, P3_SUB_357_1258_U275, P3_SUB_357_1258_U304);
  and ginst23491 (P3_SUB_357_1258_U13, P3_SUB_357_1258_U11, P3_SUB_357_1258_U213);
  and ginst23492 (P3_SUB_357_1258_U130, P3_SUB_357_1258_U378, P3_SUB_357_1258_U379);
  nand ginst23493 (P3_SUB_357_1258_U131, P3_SUB_357_1258_U106, P3_SUB_357_1258_U218);
  and ginst23494 (P3_SUB_357_1258_U132, P3_SUB_357_1258_U392, P3_SUB_357_1258_U393);
  nand ginst23495 (P3_SUB_357_1258_U133, P3_SUB_357_1258_U14, P3_SUB_357_1258_U282);
  and ginst23496 (P3_SUB_357_1258_U134, P3_SUB_357_1258_U399, P3_SUB_357_1258_U400);
  nand ginst23497 (P3_SUB_357_1258_U135, P3_SUB_357_1258_U12, P3_SUB_357_1258_U280);
  and ginst23498 (P3_SUB_357_1258_U136, P3_SUB_357_1258_U406, P3_SUB_357_1258_U407);
  nand ginst23499 (P3_SUB_357_1258_U137, P3_SUB_357_1258_U10, P3_SUB_357_1258_U278);
  and ginst23500 (P3_SUB_357_1258_U138, P3_SUB_357_1258_U413, P3_SUB_357_1258_U414);
  nand ginst23501 (P3_SUB_357_1258_U139, P3_SUB_357_1258_U111, P3_SUB_357_1258_U236);
  and ginst23502 (P3_SUB_357_1258_U14, P3_SUB_357_1258_U12, P3_SUB_357_1258_U214);
  and ginst23503 (P3_SUB_357_1258_U140, P3_SUB_357_1258_U432, P3_SUB_357_1258_U433);
  nand ginst23504 (P3_SUB_357_1258_U141, P3_SUB_357_1258_U201, P3_SUB_357_1258_U272, P3_SUB_357_1258_U273);
  and ginst23505 (P3_SUB_357_1258_U142, P3_SUB_357_1258_U443, P3_SUB_357_1258_U444);
  nand ginst23506 (P3_SUB_357_1258_U143, P3_SUB_357_1258_U198, P3_SUB_357_1258_U199);
  and ginst23507 (P3_SUB_357_1258_U144, P3_SUB_357_1258_U450, P3_SUB_357_1258_U451);
  nand ginst23508 (P3_SUB_357_1258_U145, P3_SUB_357_1258_U194, P3_SUB_357_1258_U195);
  and ginst23509 (P3_SUB_357_1258_U146, P3_SUB_357_1258_U457, P3_SUB_357_1258_U458);
  nand ginst23510 (P3_SUB_357_1258_U147, P3_SUB_357_1258_U100, P3_SUB_357_1258_U292);
  and ginst23511 (P3_SUB_357_1258_U148, P3_SUB_357_1258_U471, P3_SUB_357_1258_U472);
  nand ginst23512 (P3_SUB_357_1258_U149, P3_SUB_357_1258_U288, P3_SUB_357_1258_U5);
  and ginst23513 (P3_SUB_357_1258_U15, P3_SUB_357_1258_U252, P3_SUB_357_1258_U255);
  nand ginst23514 (P3_SUB_357_1258_U150, P3_SUB_357_1258_U186, P3_SUB_357_1258_U286);
  nand ginst23515 (P3_SUB_357_1258_U151, P3_ADD_357_U6, P3_SUB_357_1258_U129);
  nand ginst23516 (P3_SUB_357_1258_U152, P3_ADD_357_U6, P3_SUB_357_1258_U117);
  nand ginst23517 (P3_SUB_357_1258_U153, P3_SUB_357_1258_U217, P3_SUB_357_1258_U39);
  nand ginst23518 (P3_SUB_357_1258_U154, P3_SUB_357_1258_U191, P3_SUB_357_1258_U39);
  nand ginst23519 (P3_SUB_357_1258_U155, P3_INSTADDRPOINTER_REG_12__SCAN_IN, P3_ADD_357_U6);
  nand ginst23520 (P3_SUB_357_1258_U156, P3_INSTADDRPOINTER_REG_20__SCAN_IN, P3_ADD_357_U6);
  nand ginst23521 (P3_SUB_357_1258_U157, P3_INSTADDRPOINTER_REG_25__SCAN_IN, P3_ADD_357_U6);
  not ginst23522 (P3_SUB_357_1258_U158, P3_SUB_357_1258_U66);
  nand ginst23523 (P3_SUB_357_1258_U159, P3_INSTADDRPOINTER_REG_2__SCAN_IN, P3_ADD_357_U13);
  and ginst23524 (P3_SUB_357_1258_U16, P3_SUB_357_1258_U248, P3_SUB_357_1258_U249);
  or ginst23525 (P3_SUB_357_1258_U160, P3_INSTADDRPOINTER_REG_4__SCAN_IN, P3_ADD_357_U19);
  not ginst23526 (P3_SUB_357_1258_U161, P3_SUB_357_1258_U30);
  nand ginst23527 (P3_SUB_357_1258_U162, P3_INSTADDRPOINTER_REG_4__SCAN_IN, P3_ADD_357_U19);
  or ginst23528 (P3_SUB_357_1258_U163, P3_INSTADDRPOINTER_REG_3__SCAN_IN, P3_ADD_357_U7);
  or ginst23529 (P3_SUB_357_1258_U164, P3_INSTADDRPOINTER_REG_2__SCAN_IN, P3_ADD_357_U13);
  not ginst23530 (P3_SUB_357_1258_U165, P3_SUB_357_1258_U127);
  nand ginst23531 (P3_SUB_357_1258_U166, P3_SUB_357_1258_U159, P3_SUB_357_1258_U270, P3_SUB_357_1258_U271, P3_SUB_357_1258_U66);
  nand ginst23532 (P3_SUB_357_1258_U167, P3_SUB_357_1258_U166, P3_SUB_357_1258_U94);
  nand ginst23533 (P3_SUB_357_1258_U168, P3_SUB_357_1258_U160, P3_SUB_357_1258_U95);
  not ginst23534 (P3_SUB_357_1258_U169, P3_SUB_357_1258_U123);
  and ginst23535 (P3_SUB_357_1258_U17, P3_SUB_357_1258_U241, P3_SUB_357_1258_U244);
  or ginst23536 (P3_SUB_357_1258_U170, P3_INSTADDRPOINTER_REG_5__SCAN_IN, P3_ADD_357_U8);
  or ginst23537 (P3_SUB_357_1258_U171, P3_INSTADDRPOINTER_REG_6__SCAN_IN, P3_ADD_357_U17);
  nand ginst23538 (P3_SUB_357_1258_U172, P3_SUB_357_1258_U121, P3_SUB_357_1258_U171);
  nand ginst23539 (P3_SUB_357_1258_U173, P3_INSTADDRPOINTER_REG_6__SCAN_IN, P3_ADD_357_U17);
  not ginst23540 (P3_SUB_357_1258_U174, P3_SUB_357_1258_U119);
  or ginst23541 (P3_SUB_357_1258_U175, P3_INSTADDRPOINTER_REG_7__SCAN_IN, P3_ADD_357_U9);
  nand ginst23542 (P3_SUB_357_1258_U176, P3_INSTADDRPOINTER_REG_8__SCAN_IN, P3_SUB_357_1258_U117);
  not ginst23543 (P3_SUB_357_1258_U177, P3_SUB_357_1258_U115);
  or ginst23544 (P3_SUB_357_1258_U178, P3_INSTADDRPOINTER_REG_9__SCAN_IN, P3_ADD_357_U6);
  nand ginst23545 (P3_SUB_357_1258_U179, P3_INSTADDRPOINTER_REG_9__SCAN_IN, P3_ADD_357_U6);
  and ginst23546 (P3_SUB_357_1258_U18, P3_SUB_357_1258_U230, P3_SUB_357_1258_U233);
  nand ginst23547 (P3_SUB_357_1258_U180, P3_SUB_357_1258_U166, P3_SUB_357_1258_U97);
  nand ginst23548 (P3_SUB_357_1258_U181, P3_INSTADDRPOINTER_REG_3__SCAN_IN, P3_ADD_357_U7);
  not ginst23549 (P3_SUB_357_1258_U182, P3_SUB_357_1258_U124);
  nand ginst23550 (P3_SUB_357_1258_U183, P3_SUB_357_1258_U127, P3_SUB_357_1258_U164);
  not ginst23551 (P3_SUB_357_1258_U184, P3_SUB_357_1258_U125);
  nand ginst23552 (P3_SUB_357_1258_U185, P3_INSTADDRPOINTER_REG_3__SCAN_IN, P3_ADD_357_U7);
  nand ginst23553 (P3_SUB_357_1258_U186, P3_INSTADDRPOINTER_REG_9__SCAN_IN, P3_ADD_357_U6);
  or ginst23554 (P3_SUB_357_1258_U187, P3_INSTADDRPOINTER_REG_10__SCAN_IN, P3_ADD_357_U6);
  nand ginst23555 (P3_SUB_357_1258_U188, P3_INSTADDRPOINTER_REG_10__SCAN_IN, P3_ADD_357_U6);
  or ginst23556 (P3_SUB_357_1258_U189, P3_INSTADDRPOINTER_REG_11__SCAN_IN, P3_ADD_357_U6);
  and ginst23557 (P3_SUB_357_1258_U19, P3_SUB_357_1258_U227, P3_SUB_357_1258_U303);
  nand ginst23558 (P3_SUB_357_1258_U190, P3_INSTADDRPOINTER_REG_11__SCAN_IN, P3_ADD_357_U6);
  nand ginst23559 (P3_SUB_357_1258_U191, P3_INSTADDRPOINTER_REG_12__SCAN_IN, P3_INSTADDRPOINTER_REG_13__SCAN_IN);
  nand ginst23560 (P3_SUB_357_1258_U192, P3_INSTADDRPOINTER_REG_13__SCAN_IN, P3_ADD_357_U6);
  or ginst23561 (P3_SUB_357_1258_U193, P3_INSTADDRPOINTER_REG_14__SCAN_IN, P3_ADD_357_U6);
  nand ginst23562 (P3_SUB_357_1258_U194, P3_SUB_357_1258_U147, P3_SUB_357_1258_U193);
  nand ginst23563 (P3_SUB_357_1258_U195, P3_INSTADDRPOINTER_REG_14__SCAN_IN, P3_ADD_357_U6);
  not ginst23564 (P3_SUB_357_1258_U196, P3_SUB_357_1258_U145);
  or ginst23565 (P3_SUB_357_1258_U197, P3_INSTADDRPOINTER_REG_15__SCAN_IN, P3_ADD_357_U6);
  nand ginst23566 (P3_SUB_357_1258_U198, P3_SUB_357_1258_U145, P3_SUB_357_1258_U197);
  nand ginst23567 (P3_SUB_357_1258_U199, P3_INSTADDRPOINTER_REG_15__SCAN_IN, P3_ADD_357_U6);
  and ginst23568 (P3_SUB_357_1258_U20, P3_SUB_357_1258_U225, P3_SUB_357_1258_U296);
  not ginst23569 (P3_SUB_357_1258_U200, P3_SUB_357_1258_U143);
  nand ginst23570 (P3_SUB_357_1258_U201, P3_SUB_357_1258_U101, P3_SUB_357_1258_U143);
  not ginst23571 (P3_SUB_357_1258_U202, P3_SUB_357_1258_U67);
  not ginst23572 (P3_SUB_357_1258_U203, P3_SUB_357_1258_U141);
  or ginst23573 (P3_SUB_357_1258_U204, P3_INSTADDRPOINTER_REG_18__SCAN_IN, P3_ADD_357_U6);
  nand ginst23574 (P3_SUB_357_1258_U205, P3_INSTADDRPOINTER_REG_18__SCAN_IN, P3_ADD_357_U6);
  nand ginst23575 (P3_SUB_357_1258_U206, P3_INSTADDRPOINTER_REG_19__SCAN_IN, P3_ADD_357_U6);
  not ginst23576 (P3_SUB_357_1258_U207, P3_SUB_357_1258_U57);
  nand ginst23577 (P3_SUB_357_1258_U208, P3_INSTADDRPOINTER_REG_21__SCAN_IN, P3_SUB_357_1258_U207);
  nand ginst23578 (P3_SUB_357_1258_U209, P3_SUB_357_1258_U208, P3_SUB_357_1258_U39);
  nand ginst23579 (P3_SUB_357_1258_U21, P3_SUB_357_1258_U307, P3_SUB_357_1258_U425, P3_SUB_357_1258_U426);
  nand ginst23580 (P3_SUB_357_1258_U210, P3_INSTADDRPOINTER_REG_21__SCAN_IN, P3_ADD_357_U6);
  or ginst23581 (P3_SUB_357_1258_U211, P3_INSTADDRPOINTER_REG_22__SCAN_IN, P3_ADD_357_U6);
  nand ginst23582 (P3_SUB_357_1258_U212, P3_INSTADDRPOINTER_REG_22__SCAN_IN, P3_ADD_357_U6);
  or ginst23583 (P3_SUB_357_1258_U213, P3_INSTADDRPOINTER_REG_23__SCAN_IN, P3_ADD_357_U6);
  nand ginst23584 (P3_SUB_357_1258_U214, P3_INSTADDRPOINTER_REG_23__SCAN_IN, P3_ADD_357_U6);
  or ginst23585 (P3_SUB_357_1258_U215, P3_INSTADDRPOINTER_REG_24__SCAN_IN, P3_ADD_357_U6);
  nand ginst23586 (P3_SUB_357_1258_U216, P3_INSTADDRPOINTER_REG_24__SCAN_IN, P3_ADD_357_U6);
  nand ginst23587 (P3_SUB_357_1258_U217, P3_INSTADDRPOINTER_REG_25__SCAN_IN, P3_INSTADDRPOINTER_REG_26__SCAN_IN);
  nand ginst23588 (P3_SUB_357_1258_U218, P3_SUB_357_1258_U153, P3_SUB_357_1258_U63);
  nand ginst23589 (P3_SUB_357_1258_U219, P3_INSTADDRPOINTER_REG_26__SCAN_IN, P3_ADD_357_U6);
  not ginst23590 (P3_SUB_357_1258_U22, P3_ADD_357_U9);
  not ginst23591 (P3_SUB_357_1258_U220, P3_SUB_357_1258_U131);
  not ginst23592 (P3_SUB_357_1258_U221, P3_SUB_357_1258_U62);
  nand ginst23593 (P3_SUB_357_1258_U222, P3_INSTADDRPOINTER_REG_29__SCAN_IN, P3_SUB_357_1258_U129);
  not ginst23594 (P3_SUB_357_1258_U223, P3_SUB_357_1258_U61);
  nand ginst23595 (P3_SUB_357_1258_U224, P3_SUB_357_1258_U107, P3_SUB_357_1258_U151);
  nand ginst23596 (P3_SUB_357_1258_U225, P3_SUB_357_1258_U294, P3_SUB_357_1258_U353, P3_SUB_357_1258_U354);
  nand ginst23597 (P3_SUB_357_1258_U226, P3_INSTADDRPOINTER_REG_28__SCAN_IN, P3_SUB_357_1258_U221);
  nand ginst23598 (P3_SUB_357_1258_U227, P3_SUB_357_1258_U376, P3_SUB_357_1258_U377, P3_SUB_357_1258_U62);
  or ginst23599 (P3_SUB_357_1258_U228, P3_INSTADDRPOINTER_REG_25__SCAN_IN, P3_ADD_357_U6);
  nand ginst23600 (P3_SUB_357_1258_U229, P3_SUB_357_1258_U228, P3_SUB_357_1258_U63);
  not ginst23601 (P3_SUB_357_1258_U23, P3_INSTADDRPOINTER_REG_7__SCAN_IN);
  nand ginst23602 (P3_SUB_357_1258_U230, P3_SUB_357_1258_U109, P3_SUB_357_1258_U229);
  nand ginst23603 (P3_SUB_357_1258_U231, P3_SUB_357_1258_U157, P3_SUB_357_1258_U285);
  nand ginst23604 (P3_SUB_357_1258_U232, P3_INSTADDRPOINTER_REG_26__SCAN_IN, P3_ADD_357_U6);
  nand ginst23605 (P3_SUB_357_1258_U233, P3_SUB_357_1258_U110, P3_SUB_357_1258_U231);
  or ginst23606 (P3_SUB_357_1258_U234, P3_INSTADDRPOINTER_REG_25__SCAN_IN, P3_ADD_357_U6);
  not ginst23607 (P3_SUB_357_1258_U235, P3_SUB_357_1258_U65);
  nand ginst23608 (P3_SUB_357_1258_U236, P3_ADD_357_U6, P3_SUB_357_1258_U65);
  nand ginst23609 (P3_SUB_357_1258_U237, P3_SUB_357_1258_U207, P3_SUB_357_1258_U64);
  not ginst23610 (P3_SUB_357_1258_U238, P3_SUB_357_1258_U139);
  nand ginst23611 (P3_SUB_357_1258_U239, P3_INSTADDRPOINTER_REG_20__SCAN_IN, P3_SUB_357_1258_U235);
  not ginst23612 (P3_SUB_357_1258_U24, P3_ADD_357_U8);
  nand ginst23613 (P3_SUB_357_1258_U240, P3_INSTADDRPOINTER_REG_19__SCAN_IN, P3_SUB_357_1258_U64);
  nand ginst23614 (P3_SUB_357_1258_U241, P3_SUB_357_1258_U240, P3_SUB_357_1258_U420, P3_SUB_357_1258_U421);
  nand ginst23615 (P3_SUB_357_1258_U242, P3_SUB_357_1258_U206, P3_SUB_357_1258_U277);
  nand ginst23616 (P3_SUB_357_1258_U243, P3_SUB_357_1258_U39, P3_SUB_357_1258_U57);
  nand ginst23617 (P3_SUB_357_1258_U244, P3_SUB_357_1258_U112, P3_SUB_357_1258_U242);
  or ginst23618 (P3_SUB_357_1258_U245, P3_INSTADDRPOINTER_REG_19__SCAN_IN, P3_ADD_357_U6);
  nand ginst23619 (P3_SUB_357_1258_U246, P3_INSTADDRPOINTER_REG_17__SCAN_IN, P3_SUB_357_1258_U202);
  nand ginst23620 (P3_SUB_357_1258_U247, P3_INSTADDRPOINTER_REG_16__SCAN_IN, P3_SUB_357_1258_U143);
  nand ginst23621 (P3_SUB_357_1258_U248, P3_SUB_357_1258_U247, P3_SUB_357_1258_U439, P3_SUB_357_1258_U440);
  nand ginst23622 (P3_SUB_357_1258_U249, P3_SUB_357_1258_U441, P3_SUB_357_1258_U442, P3_SUB_357_1258_U67);
  not ginst23623 (P3_SUB_357_1258_U25, P3_INSTADDRPOINTER_REG_5__SCAN_IN);
  or ginst23624 (P3_SUB_357_1258_U250, P3_INSTADDRPOINTER_REG_12__SCAN_IN, P3_ADD_357_U6);
  nand ginst23625 (P3_SUB_357_1258_U251, P3_SUB_357_1258_U250, P3_SUB_357_1258_U68);
  nand ginst23626 (P3_SUB_357_1258_U252, P3_SUB_357_1258_U113, P3_SUB_357_1258_U251);
  nand ginst23627 (P3_SUB_357_1258_U253, P3_SUB_357_1258_U155, P3_SUB_357_1258_U291);
  nand ginst23628 (P3_SUB_357_1258_U254, P3_INSTADDRPOINTER_REG_13__SCAN_IN, P3_ADD_357_U6);
  nand ginst23629 (P3_SUB_357_1258_U255, P3_SUB_357_1258_U114, P3_SUB_357_1258_U253);
  or ginst23630 (P3_SUB_357_1258_U256, P3_INSTADDRPOINTER_REG_12__SCAN_IN, P3_ADD_357_U6);
  nand ginst23631 (P3_SUB_357_1258_U257, P3_INSTADDRPOINTER_REG_10__SCAN_IN, P3_ADD_357_U6);
  nand ginst23632 (P3_SUB_357_1258_U258, P3_SUB_357_1258_U178, P3_SUB_357_1258_U179);
  nand ginst23633 (P3_SUB_357_1258_U259, P3_SUB_357_1258_U160, P3_SUB_357_1258_U162);
  not ginst23634 (P3_SUB_357_1258_U26, P3_ADD_357_U19);
  nand ginst23635 (P3_SUB_357_1258_U260, P3_SUB_357_1258_U163, P3_SUB_357_1258_U185);
  nand ginst23636 (P3_SUB_357_1258_U261, P3_SUB_357_1258_U159, P3_SUB_357_1258_U164);
  nand ginst23637 (P3_SUB_357_1258_U262, P3_SUB_357_1258_U157, P3_SUB_357_1258_U234);
  nand ginst23638 (P3_SUB_357_1258_U263, P3_SUB_357_1258_U206, P3_SUB_357_1258_U245);
  nand ginst23639 (P3_SUB_357_1258_U264, P3_SUB_357_1258_U155, P3_SUB_357_1258_U256);
  nand ginst23640 (P3_SUB_357_1258_U265, P3_SUB_357_1258_U187, P3_SUB_357_1258_U257);
  nand ginst23641 (P3_SUB_357_1258_U266, P3_INSTADDRPOINTER_REG_5__SCAN_IN, P3_ADD_357_U8);
  nand ginst23642 (P3_SUB_357_1258_U267, P3_INSTADDRPOINTER_REG_7__SCAN_IN, P3_ADD_357_U9);
  nand ginst23643 (P3_SUB_357_1258_U268, P3_INSTADDRPOINTER_REG_8__SCAN_IN, P3_ADD_357_U6);
  nand ginst23644 (P3_SUB_357_1258_U269, P3_INSTADDRPOINTER_REG_29__SCAN_IN, P3_ADD_357_U6);
  not ginst23645 (P3_SUB_357_1258_U27, P3_INSTADDRPOINTER_REG_4__SCAN_IN);
  nand ginst23646 (P3_SUB_357_1258_U270, P3_INSTADDRPOINTER_REG_1__SCAN_IN, P3_SUB_357_1258_U161);
  nand ginst23647 (P3_SUB_357_1258_U271, P3_INSTADDRPOINTER_REG_1__SCAN_IN, P3_SUB_357_U7);
  nand ginst23648 (P3_SUB_357_1258_U272, P3_ADD_357_U6, P3_SUB_357_1258_U67);
  nand ginst23649 (P3_SUB_357_1258_U273, P3_INSTADDRPOINTER_REG_17__SCAN_IN, P3_ADD_357_U6);
  nand ginst23650 (P3_SUB_357_1258_U274, P3_ADD_357_U6, P3_SUB_357_1258_U62);
  nand ginst23651 (P3_SUB_357_1258_U275, P3_INSTADDRPOINTER_REG_28__SCAN_IN, P3_ADD_357_U6);
  nand ginst23652 (P3_SUB_357_1258_U276, P3_SUB_357_1258_U141, P3_SUB_357_1258_U204);
  not ginst23653 (P3_SUB_357_1258_U277, P3_SUB_357_1258_U64);
  nand ginst23654 (P3_SUB_357_1258_U278, P3_SUB_357_1258_U141, P3_SUB_357_1258_U9);
  not ginst23655 (P3_SUB_357_1258_U279, P3_SUB_357_1258_U137);
  not ginst23656 (P3_SUB_357_1258_U28, P3_ADD_357_U10);
  nand ginst23657 (P3_SUB_357_1258_U280, P3_SUB_357_1258_U11, P3_SUB_357_1258_U141);
  not ginst23658 (P3_SUB_357_1258_U281, P3_SUB_357_1258_U135);
  nand ginst23659 (P3_SUB_357_1258_U282, P3_SUB_357_1258_U13, P3_SUB_357_1258_U141);
  not ginst23660 (P3_SUB_357_1258_U283, P3_SUB_357_1258_U133);
  nand ginst23661 (P3_SUB_357_1258_U284, P3_SUB_357_1258_U103, P3_SUB_357_1258_U141);
  not ginst23662 (P3_SUB_357_1258_U285, P3_SUB_357_1258_U63);
  nand ginst23663 (P3_SUB_357_1258_U286, P3_SUB_357_1258_U115, P3_SUB_357_1258_U178);
  not ginst23664 (P3_SUB_357_1258_U287, P3_SUB_357_1258_U150);
  nand ginst23665 (P3_SUB_357_1258_U288, P3_SUB_357_1258_U115, P3_SUB_357_1258_U6);
  not ginst23666 (P3_SUB_357_1258_U289, P3_SUB_357_1258_U149);
  not ginst23667 (P3_SUB_357_1258_U29, P3_INSTADDRPOINTER_REG_0__SCAN_IN);
  nand ginst23668 (P3_SUB_357_1258_U290, P3_SUB_357_1258_U115, P3_SUB_357_1258_U7);
  not ginst23669 (P3_SUB_357_1258_U291, P3_SUB_357_1258_U68);
  nand ginst23670 (P3_SUB_357_1258_U292, P3_SUB_357_1258_U115, P3_SUB_357_1258_U98);
  not ginst23671 (P3_SUB_357_1258_U293, P3_SUB_357_1258_U147);
  nand ginst23672 (P3_SUB_357_1258_U294, P3_SUB_357_1258_U223, P3_SUB_357_1258_U60);
  nand ginst23673 (P3_SUB_357_1258_U295, P3_INSTADDRPOINTER_REG_30__SCAN_IN, P3_SUB_357_1258_U61);
  nand ginst23674 (P3_SUB_357_1258_U296, P3_SUB_357_1258_U295, P3_SUB_357_1258_U351, P3_SUB_357_1258_U352);
  nand ginst23675 (P3_SUB_357_1258_U297, P3_SUB_357_1258_U108, P3_SUB_357_1258_U61);
  nand ginst23676 (P3_SUB_357_1258_U298, P3_SUB_357_1258_U123, P3_SUB_357_1258_U170);
  not ginst23677 (P3_SUB_357_1258_U299, P3_SUB_357_1258_U121);
  nand ginst23678 (P3_SUB_357_1258_U30, P3_INSTADDRPOINTER_REG_0__SCAN_IN, P3_ADD_357_U10);
  nand ginst23679 (P3_SUB_357_1258_U300, P3_SUB_357_1258_U119, P3_SUB_357_1258_U175);
  not ginst23680 (P3_SUB_357_1258_U301, P3_SUB_357_1258_U117);
  nand ginst23681 (P3_SUB_357_1258_U302, P3_INSTADDRPOINTER_REG_27__SCAN_IN, P3_SUB_357_1258_U131);
  nand ginst23682 (P3_SUB_357_1258_U303, P3_SUB_357_1258_U302, P3_SUB_357_1258_U374, P3_SUB_357_1258_U375);
  nand ginst23683 (P3_SUB_357_1258_U304, P3_SUB_357_1258_U131, P3_SUB_357_1258_U4);
  not ginst23684 (P3_SUB_357_1258_U305, P3_SUB_357_1258_U129);
  nand ginst23685 (P3_SUB_357_1258_U306, P3_SUB_357_1258_U131, P3_SUB_357_1258_U4);
  nand ginst23686 (P3_SUB_357_1258_U307, P3_INSTADDRPOINTER_REG_1__SCAN_IN, P3_SUB_357_1258_U158);
  nand ginst23687 (P3_SUB_357_1258_U308, P3_ADD_357_U6, P3_SUB_357_1258_U41);
  nand ginst23688 (P3_SUB_357_1258_U309, P3_INSTADDRPOINTER_REG_9__SCAN_IN, P3_SUB_357_1258_U39);
  not ginst23689 (P3_SUB_357_1258_U31, P3_SUB_357_U7);
  nand ginst23690 (P3_SUB_357_1258_U310, P3_SUB_357_1258_U308, P3_SUB_357_1258_U309);
  nand ginst23691 (P3_SUB_357_1258_U311, P3_SUB_357_1258_U115, P3_SUB_357_1258_U258);
  nand ginst23692 (P3_SUB_357_1258_U312, P3_SUB_357_1258_U177, P3_SUB_357_1258_U310);
  nand ginst23693 (P3_SUB_357_1258_U313, P3_ADD_357_U6, P3_SUB_357_1258_U40);
  nand ginst23694 (P3_SUB_357_1258_U314, P3_INSTADDRPOINTER_REG_8__SCAN_IN, P3_SUB_357_1258_U39);
  nand ginst23695 (P3_SUB_357_1258_U315, P3_ADD_357_U6, P3_SUB_357_1258_U40);
  nand ginst23696 (P3_SUB_357_1258_U316, P3_INSTADDRPOINTER_REG_8__SCAN_IN, P3_SUB_357_1258_U39);
  nand ginst23697 (P3_SUB_357_1258_U317, P3_SUB_357_1258_U315, P3_SUB_357_1258_U316);
  nand ginst23698 (P3_SUB_357_1258_U318, P3_SUB_357_1258_U116, P3_SUB_357_1258_U117);
  nand ginst23699 (P3_SUB_357_1258_U319, P3_SUB_357_1258_U301, P3_SUB_357_1258_U317);
  not ginst23700 (P3_SUB_357_1258_U32, P3_ADD_357_U13);
  nand ginst23701 (P3_SUB_357_1258_U320, P3_INSTADDRPOINTER_REG_7__SCAN_IN, P3_SUB_357_1258_U22);
  nand ginst23702 (P3_SUB_357_1258_U321, P3_ADD_357_U9, P3_SUB_357_1258_U23);
  nand ginst23703 (P3_SUB_357_1258_U322, P3_INSTADDRPOINTER_REG_7__SCAN_IN, P3_SUB_357_1258_U22);
  nand ginst23704 (P3_SUB_357_1258_U323, P3_ADD_357_U9, P3_SUB_357_1258_U23);
  nand ginst23705 (P3_SUB_357_1258_U324, P3_SUB_357_1258_U322, P3_SUB_357_1258_U323);
  nand ginst23706 (P3_SUB_357_1258_U325, P3_SUB_357_1258_U118, P3_SUB_357_1258_U119);
  nand ginst23707 (P3_SUB_357_1258_U326, P3_SUB_357_1258_U174, P3_SUB_357_1258_U324);
  nand ginst23708 (P3_SUB_357_1258_U327, P3_INSTADDRPOINTER_REG_6__SCAN_IN, P3_SUB_357_1258_U37);
  nand ginst23709 (P3_SUB_357_1258_U328, P3_ADD_357_U17, P3_SUB_357_1258_U38);
  nand ginst23710 (P3_SUB_357_1258_U329, P3_INSTADDRPOINTER_REG_6__SCAN_IN, P3_SUB_357_1258_U37);
  not ginst23711 (P3_SUB_357_1258_U33, P3_INSTADDRPOINTER_REG_2__SCAN_IN);
  nand ginst23712 (P3_SUB_357_1258_U330, P3_ADD_357_U17, P3_SUB_357_1258_U38);
  nand ginst23713 (P3_SUB_357_1258_U331, P3_SUB_357_1258_U329, P3_SUB_357_1258_U330);
  nand ginst23714 (P3_SUB_357_1258_U332, P3_SUB_357_1258_U120, P3_SUB_357_1258_U121);
  nand ginst23715 (P3_SUB_357_1258_U333, P3_SUB_357_1258_U299, P3_SUB_357_1258_U331);
  nand ginst23716 (P3_SUB_357_1258_U334, P3_INSTADDRPOINTER_REG_5__SCAN_IN, P3_SUB_357_1258_U24);
  nand ginst23717 (P3_SUB_357_1258_U335, P3_ADD_357_U8, P3_SUB_357_1258_U25);
  nand ginst23718 (P3_SUB_357_1258_U336, P3_INSTADDRPOINTER_REG_5__SCAN_IN, P3_SUB_357_1258_U24);
  nand ginst23719 (P3_SUB_357_1258_U337, P3_ADD_357_U8, P3_SUB_357_1258_U25);
  nand ginst23720 (P3_SUB_357_1258_U338, P3_SUB_357_1258_U336, P3_SUB_357_1258_U337);
  nand ginst23721 (P3_SUB_357_1258_U339, P3_SUB_357_1258_U122, P3_SUB_357_1258_U123);
  not ginst23722 (P3_SUB_357_1258_U34, P3_INSTADDRPOINTER_REG_1__SCAN_IN);
  nand ginst23723 (P3_SUB_357_1258_U340, P3_SUB_357_1258_U169, P3_SUB_357_1258_U338);
  nand ginst23724 (P3_SUB_357_1258_U341, P3_INSTADDRPOINTER_REG_4__SCAN_IN, P3_SUB_357_1258_U26);
  nand ginst23725 (P3_SUB_357_1258_U342, P3_ADD_357_U19, P3_SUB_357_1258_U27);
  nand ginst23726 (P3_SUB_357_1258_U343, P3_SUB_357_1258_U341, P3_SUB_357_1258_U342);
  nand ginst23727 (P3_SUB_357_1258_U344, P3_SUB_357_1258_U124, P3_SUB_357_1258_U259);
  nand ginst23728 (P3_SUB_357_1258_U345, P3_SUB_357_1258_U182, P3_SUB_357_1258_U343);
  nand ginst23729 (P3_SUB_357_1258_U346, P3_INSTADDRPOINTER_REG_3__SCAN_IN, P3_SUB_357_1258_U35);
  nand ginst23730 (P3_SUB_357_1258_U347, P3_ADD_357_U7, P3_SUB_357_1258_U36);
  nand ginst23731 (P3_SUB_357_1258_U348, P3_SUB_357_1258_U346, P3_SUB_357_1258_U347);
  nand ginst23732 (P3_SUB_357_1258_U349, P3_SUB_357_1258_U125, P3_SUB_357_1258_U260);
  not ginst23733 (P3_SUB_357_1258_U35, P3_ADD_357_U7);
  nand ginst23734 (P3_SUB_357_1258_U350, P3_SUB_357_1258_U184, P3_SUB_357_1258_U348);
  nand ginst23735 (P3_SUB_357_1258_U351, P3_INSTADDRPOINTER_REG_31__SCAN_IN, P3_SUB_357_1258_U39);
  nand ginst23736 (P3_SUB_357_1258_U352, P3_ADD_357_U6, P3_SUB_357_1258_U224);
  nand ginst23737 (P3_SUB_357_1258_U353, P3_INSTADDRPOINTER_REG_31__SCAN_IN, P3_ADD_357_U6);
  nand ginst23738 (P3_SUB_357_1258_U354, P3_SUB_357_1258_U297, P3_SUB_357_1258_U39);
  nand ginst23739 (P3_SUB_357_1258_U355, P3_ADD_357_U6, P3_SUB_357_1258_U60);
  nand ginst23740 (P3_SUB_357_1258_U356, P3_INSTADDRPOINTER_REG_30__SCAN_IN, P3_SUB_357_1258_U39);
  nand ginst23741 (P3_SUB_357_1258_U357, P3_ADD_357_U6, P3_SUB_357_1258_U60);
  nand ginst23742 (P3_SUB_357_1258_U358, P3_INSTADDRPOINTER_REG_30__SCAN_IN, P3_SUB_357_1258_U39);
  nand ginst23743 (P3_SUB_357_1258_U359, P3_SUB_357_1258_U357, P3_SUB_357_1258_U358);
  not ginst23744 (P3_SUB_357_1258_U36, P3_INSTADDRPOINTER_REG_3__SCAN_IN);
  nand ginst23745 (P3_SUB_357_1258_U360, P3_SUB_357_1258_U126, P3_SUB_357_1258_U61);
  nand ginst23746 (P3_SUB_357_1258_U361, P3_SUB_357_1258_U223, P3_SUB_357_1258_U359);
  nand ginst23747 (P3_SUB_357_1258_U362, P3_INSTADDRPOINTER_REG_2__SCAN_IN, P3_SUB_357_1258_U32);
  nand ginst23748 (P3_SUB_357_1258_U363, P3_ADD_357_U13, P3_SUB_357_1258_U33);
  nand ginst23749 (P3_SUB_357_1258_U364, P3_SUB_357_1258_U362, P3_SUB_357_1258_U363);
  nand ginst23750 (P3_SUB_357_1258_U365, P3_SUB_357_1258_U127, P3_SUB_357_1258_U261);
  nand ginst23751 (P3_SUB_357_1258_U366, P3_SUB_357_1258_U165, P3_SUB_357_1258_U364);
  nand ginst23752 (P3_SUB_357_1258_U367, P3_ADD_357_U6, P3_SUB_357_1258_U59);
  nand ginst23753 (P3_SUB_357_1258_U368, P3_INSTADDRPOINTER_REG_29__SCAN_IN, P3_SUB_357_1258_U39);
  nand ginst23754 (P3_SUB_357_1258_U369, P3_ADD_357_U6, P3_SUB_357_1258_U59);
  not ginst23755 (P3_SUB_357_1258_U37, P3_ADD_357_U17);
  nand ginst23756 (P3_SUB_357_1258_U370, P3_INSTADDRPOINTER_REG_29__SCAN_IN, P3_SUB_357_1258_U39);
  nand ginst23757 (P3_SUB_357_1258_U371, P3_SUB_357_1258_U369, P3_SUB_357_1258_U370);
  nand ginst23758 (P3_SUB_357_1258_U372, P3_SUB_357_1258_U128, P3_SUB_357_1258_U129);
  nand ginst23759 (P3_SUB_357_1258_U373, P3_SUB_357_1258_U305, P3_SUB_357_1258_U371);
  nand ginst23760 (P3_SUB_357_1258_U374, P3_INSTADDRPOINTER_REG_28__SCAN_IN, P3_SUB_357_1258_U39);
  nand ginst23761 (P3_SUB_357_1258_U375, P3_ADD_357_U6, P3_SUB_357_1258_U226);
  nand ginst23762 (P3_SUB_357_1258_U376, P3_INSTADDRPOINTER_REG_28__SCAN_IN, P3_ADD_357_U6);
  nand ginst23763 (P3_SUB_357_1258_U377, P3_SUB_357_1258_U306, P3_SUB_357_1258_U39);
  nand ginst23764 (P3_SUB_357_1258_U378, P3_INSTADDRPOINTER_REG_27__SCAN_IN, P3_SUB_357_1258_U39);
  nand ginst23765 (P3_SUB_357_1258_U379, P3_ADD_357_U6, P3_SUB_357_1258_U58);
  not ginst23766 (P3_SUB_357_1258_U38, P3_INSTADDRPOINTER_REG_6__SCAN_IN);
  nand ginst23767 (P3_SUB_357_1258_U380, P3_INSTADDRPOINTER_REG_27__SCAN_IN, P3_SUB_357_1258_U39);
  nand ginst23768 (P3_SUB_357_1258_U381, P3_ADD_357_U6, P3_SUB_357_1258_U58);
  nand ginst23769 (P3_SUB_357_1258_U382, P3_SUB_357_1258_U380, P3_SUB_357_1258_U381);
  nand ginst23770 (P3_SUB_357_1258_U383, P3_SUB_357_1258_U130, P3_SUB_357_1258_U131);
  nand ginst23771 (P3_SUB_357_1258_U384, P3_SUB_357_1258_U220, P3_SUB_357_1258_U382);
  nand ginst23772 (P3_SUB_357_1258_U385, P3_INSTADDRPOINTER_REG_26__SCAN_IN, P3_SUB_357_1258_U39);
  nand ginst23773 (P3_SUB_357_1258_U386, P3_ADD_357_U6, P3_SUB_357_1258_U43);
  nand ginst23774 (P3_SUB_357_1258_U387, P3_INSTADDRPOINTER_REG_25__SCAN_IN, P3_SUB_357_1258_U39);
  nand ginst23775 (P3_SUB_357_1258_U388, P3_ADD_357_U6, P3_SUB_357_1258_U42);
  nand ginst23776 (P3_SUB_357_1258_U389, P3_SUB_357_1258_U387, P3_SUB_357_1258_U388);
  not ginst23777 (P3_SUB_357_1258_U39, P3_ADD_357_U6);
  nand ginst23778 (P3_SUB_357_1258_U390, P3_SUB_357_1258_U262, P3_SUB_357_1258_U63);
  nand ginst23779 (P3_SUB_357_1258_U391, P3_SUB_357_1258_U285, P3_SUB_357_1258_U389);
  nand ginst23780 (P3_SUB_357_1258_U392, P3_INSTADDRPOINTER_REG_24__SCAN_IN, P3_SUB_357_1258_U39);
  nand ginst23781 (P3_SUB_357_1258_U393, P3_ADD_357_U6, P3_SUB_357_1258_U44);
  nand ginst23782 (P3_SUB_357_1258_U394, P3_INSTADDRPOINTER_REG_24__SCAN_IN, P3_SUB_357_1258_U39);
  nand ginst23783 (P3_SUB_357_1258_U395, P3_ADD_357_U6, P3_SUB_357_1258_U44);
  nand ginst23784 (P3_SUB_357_1258_U396, P3_SUB_357_1258_U394, P3_SUB_357_1258_U395);
  nand ginst23785 (P3_SUB_357_1258_U397, P3_SUB_357_1258_U132, P3_SUB_357_1258_U133);
  nand ginst23786 (P3_SUB_357_1258_U398, P3_SUB_357_1258_U283, P3_SUB_357_1258_U396);
  nand ginst23787 (P3_SUB_357_1258_U399, P3_INSTADDRPOINTER_REG_23__SCAN_IN, P3_SUB_357_1258_U39);
  and ginst23788 (P3_SUB_357_1258_U4, P3_INSTADDRPOINTER_REG_27__SCAN_IN, P3_INSTADDRPOINTER_REG_28__SCAN_IN);
  not ginst23789 (P3_SUB_357_1258_U40, P3_INSTADDRPOINTER_REG_8__SCAN_IN);
  nand ginst23790 (P3_SUB_357_1258_U400, P3_ADD_357_U6, P3_SUB_357_1258_U45);
  nand ginst23791 (P3_SUB_357_1258_U401, P3_INSTADDRPOINTER_REG_23__SCAN_IN, P3_SUB_357_1258_U39);
  nand ginst23792 (P3_SUB_357_1258_U402, P3_ADD_357_U6, P3_SUB_357_1258_U45);
  nand ginst23793 (P3_SUB_357_1258_U403, P3_SUB_357_1258_U401, P3_SUB_357_1258_U402);
  nand ginst23794 (P3_SUB_357_1258_U404, P3_SUB_357_1258_U134, P3_SUB_357_1258_U135);
  nand ginst23795 (P3_SUB_357_1258_U405, P3_SUB_357_1258_U281, P3_SUB_357_1258_U403);
  nand ginst23796 (P3_SUB_357_1258_U406, P3_INSTADDRPOINTER_REG_22__SCAN_IN, P3_SUB_357_1258_U39);
  nand ginst23797 (P3_SUB_357_1258_U407, P3_ADD_357_U6, P3_SUB_357_1258_U46);
  nand ginst23798 (P3_SUB_357_1258_U408, P3_INSTADDRPOINTER_REG_22__SCAN_IN, P3_SUB_357_1258_U39);
  nand ginst23799 (P3_SUB_357_1258_U409, P3_ADD_357_U6, P3_SUB_357_1258_U46);
  not ginst23800 (P3_SUB_357_1258_U41, P3_INSTADDRPOINTER_REG_9__SCAN_IN);
  nand ginst23801 (P3_SUB_357_1258_U410, P3_SUB_357_1258_U408, P3_SUB_357_1258_U409);
  nand ginst23802 (P3_SUB_357_1258_U411, P3_SUB_357_1258_U136, P3_SUB_357_1258_U137);
  nand ginst23803 (P3_SUB_357_1258_U412, P3_SUB_357_1258_U279, P3_SUB_357_1258_U410);
  nand ginst23804 (P3_SUB_357_1258_U413, P3_INSTADDRPOINTER_REG_21__SCAN_IN, P3_SUB_357_1258_U39);
  nand ginst23805 (P3_SUB_357_1258_U414, P3_ADD_357_U6, P3_SUB_357_1258_U48);
  nand ginst23806 (P3_SUB_357_1258_U415, P3_INSTADDRPOINTER_REG_21__SCAN_IN, P3_SUB_357_1258_U39);
  nand ginst23807 (P3_SUB_357_1258_U416, P3_ADD_357_U6, P3_SUB_357_1258_U48);
  nand ginst23808 (P3_SUB_357_1258_U417, P3_SUB_357_1258_U415, P3_SUB_357_1258_U416);
  nand ginst23809 (P3_SUB_357_1258_U418, P3_SUB_357_1258_U138, P3_SUB_357_1258_U139);
  nand ginst23810 (P3_SUB_357_1258_U419, P3_SUB_357_1258_U238, P3_SUB_357_1258_U417);
  not ginst23811 (P3_SUB_357_1258_U42, P3_INSTADDRPOINTER_REG_25__SCAN_IN);
  nand ginst23812 (P3_SUB_357_1258_U420, P3_INSTADDRPOINTER_REG_20__SCAN_IN, P3_SUB_357_1258_U39);
  nand ginst23813 (P3_SUB_357_1258_U421, P3_ADD_357_U6, P3_SUB_357_1258_U239);
  nand ginst23814 (P3_SUB_357_1258_U422, P3_INSTADDRPOINTER_REG_1__SCAN_IN, P3_SUB_357_1258_U30);
  nand ginst23815 (P3_SUB_357_1258_U423, P3_SUB_357_1258_U161, P3_SUB_357_1258_U34);
  nand ginst23816 (P3_SUB_357_1258_U424, P3_SUB_357_1258_U422, P3_SUB_357_1258_U423);
  nand ginst23817 (P3_SUB_357_1258_U425, P3_SUB_357_1258_U30, P3_SUB_357_1258_U34, P3_SUB_357_U7);
  nand ginst23818 (P3_SUB_357_1258_U426, P3_SUB_357_1258_U31, P3_SUB_357_1258_U424);
  nand ginst23819 (P3_SUB_357_1258_U427, P3_INSTADDRPOINTER_REG_19__SCAN_IN, P3_SUB_357_1258_U39);
  nand ginst23820 (P3_SUB_357_1258_U428, P3_ADD_357_U6, P3_SUB_357_1258_U47);
  nand ginst23821 (P3_SUB_357_1258_U429, P3_SUB_357_1258_U427, P3_SUB_357_1258_U428);
  not ginst23822 (P3_SUB_357_1258_U43, P3_INSTADDRPOINTER_REG_26__SCAN_IN);
  nand ginst23823 (P3_SUB_357_1258_U430, P3_SUB_357_1258_U263, P3_SUB_357_1258_U64);
  nand ginst23824 (P3_SUB_357_1258_U431, P3_SUB_357_1258_U277, P3_SUB_357_1258_U429);
  nand ginst23825 (P3_SUB_357_1258_U432, P3_INSTADDRPOINTER_REG_18__SCAN_IN, P3_SUB_357_1258_U39);
  nand ginst23826 (P3_SUB_357_1258_U433, P3_ADD_357_U6, P3_SUB_357_1258_U49);
  nand ginst23827 (P3_SUB_357_1258_U434, P3_INSTADDRPOINTER_REG_18__SCAN_IN, P3_SUB_357_1258_U39);
  nand ginst23828 (P3_SUB_357_1258_U435, P3_ADD_357_U6, P3_SUB_357_1258_U49);
  nand ginst23829 (P3_SUB_357_1258_U436, P3_SUB_357_1258_U434, P3_SUB_357_1258_U435);
  nand ginst23830 (P3_SUB_357_1258_U437, P3_SUB_357_1258_U140, P3_SUB_357_1258_U141);
  nand ginst23831 (P3_SUB_357_1258_U438, P3_SUB_357_1258_U203, P3_SUB_357_1258_U436);
  nand ginst23832 (P3_SUB_357_1258_U439, P3_INSTADDRPOINTER_REG_17__SCAN_IN, P3_SUB_357_1258_U39);
  not ginst23833 (P3_SUB_357_1258_U44, P3_INSTADDRPOINTER_REG_24__SCAN_IN);
  nand ginst23834 (P3_SUB_357_1258_U440, P3_ADD_357_U6, P3_SUB_357_1258_U246);
  nand ginst23835 (P3_SUB_357_1258_U441, P3_INSTADDRPOINTER_REG_17__SCAN_IN, P3_ADD_357_U6);
  nand ginst23836 (P3_SUB_357_1258_U442, P3_SUB_357_1258_U201, P3_SUB_357_1258_U39);
  nand ginst23837 (P3_SUB_357_1258_U443, P3_INSTADDRPOINTER_REG_16__SCAN_IN, P3_SUB_357_1258_U39);
  nand ginst23838 (P3_SUB_357_1258_U444, P3_ADD_357_U6, P3_SUB_357_1258_U56);
  nand ginst23839 (P3_SUB_357_1258_U445, P3_INSTADDRPOINTER_REG_16__SCAN_IN, P3_SUB_357_1258_U39);
  nand ginst23840 (P3_SUB_357_1258_U446, P3_ADD_357_U6, P3_SUB_357_1258_U56);
  nand ginst23841 (P3_SUB_357_1258_U447, P3_SUB_357_1258_U445, P3_SUB_357_1258_U446);
  nand ginst23842 (P3_SUB_357_1258_U448, P3_SUB_357_1258_U142, P3_SUB_357_1258_U143);
  nand ginst23843 (P3_SUB_357_1258_U449, P3_SUB_357_1258_U200, P3_SUB_357_1258_U447);
  not ginst23844 (P3_SUB_357_1258_U45, P3_INSTADDRPOINTER_REG_23__SCAN_IN);
  nand ginst23845 (P3_SUB_357_1258_U450, P3_INSTADDRPOINTER_REG_15__SCAN_IN, P3_SUB_357_1258_U39);
  nand ginst23846 (P3_SUB_357_1258_U451, P3_ADD_357_U6, P3_SUB_357_1258_U55);
  nand ginst23847 (P3_SUB_357_1258_U452, P3_INSTADDRPOINTER_REG_15__SCAN_IN, P3_SUB_357_1258_U39);
  nand ginst23848 (P3_SUB_357_1258_U453, P3_ADD_357_U6, P3_SUB_357_1258_U55);
  nand ginst23849 (P3_SUB_357_1258_U454, P3_SUB_357_1258_U452, P3_SUB_357_1258_U453);
  nand ginst23850 (P3_SUB_357_1258_U455, P3_SUB_357_1258_U144, P3_SUB_357_1258_U145);
  nand ginst23851 (P3_SUB_357_1258_U456, P3_SUB_357_1258_U196, P3_SUB_357_1258_U454);
  nand ginst23852 (P3_SUB_357_1258_U457, P3_INSTADDRPOINTER_REG_14__SCAN_IN, P3_SUB_357_1258_U39);
  nand ginst23853 (P3_SUB_357_1258_U458, P3_ADD_357_U6, P3_SUB_357_1258_U54);
  nand ginst23854 (P3_SUB_357_1258_U459, P3_INSTADDRPOINTER_REG_14__SCAN_IN, P3_SUB_357_1258_U39);
  not ginst23855 (P3_SUB_357_1258_U46, P3_INSTADDRPOINTER_REG_22__SCAN_IN);
  nand ginst23856 (P3_SUB_357_1258_U460, P3_ADD_357_U6, P3_SUB_357_1258_U54);
  nand ginst23857 (P3_SUB_357_1258_U461, P3_SUB_357_1258_U459, P3_SUB_357_1258_U460);
  nand ginst23858 (P3_SUB_357_1258_U462, P3_SUB_357_1258_U146, P3_SUB_357_1258_U147);
  nand ginst23859 (P3_SUB_357_1258_U463, P3_SUB_357_1258_U293, P3_SUB_357_1258_U461);
  nand ginst23860 (P3_SUB_357_1258_U464, P3_INSTADDRPOINTER_REG_13__SCAN_IN, P3_SUB_357_1258_U39);
  nand ginst23861 (P3_SUB_357_1258_U465, P3_ADD_357_U6, P3_SUB_357_1258_U51);
  nand ginst23862 (P3_SUB_357_1258_U466, P3_INSTADDRPOINTER_REG_12__SCAN_IN, P3_SUB_357_1258_U39);
  nand ginst23863 (P3_SUB_357_1258_U467, P3_ADD_357_U6, P3_SUB_357_1258_U50);
  nand ginst23864 (P3_SUB_357_1258_U468, P3_SUB_357_1258_U466, P3_SUB_357_1258_U467);
  nand ginst23865 (P3_SUB_357_1258_U469, P3_SUB_357_1258_U264, P3_SUB_357_1258_U68);
  not ginst23866 (P3_SUB_357_1258_U47, P3_INSTADDRPOINTER_REG_19__SCAN_IN);
  nand ginst23867 (P3_SUB_357_1258_U470, P3_SUB_357_1258_U291, P3_SUB_357_1258_U468);
  nand ginst23868 (P3_SUB_357_1258_U471, P3_INSTADDRPOINTER_REG_11__SCAN_IN, P3_SUB_357_1258_U39);
  nand ginst23869 (P3_SUB_357_1258_U472, P3_ADD_357_U6, P3_SUB_357_1258_U52);
  nand ginst23870 (P3_SUB_357_1258_U473, P3_INSTADDRPOINTER_REG_11__SCAN_IN, P3_SUB_357_1258_U39);
  nand ginst23871 (P3_SUB_357_1258_U474, P3_ADD_357_U6, P3_SUB_357_1258_U52);
  nand ginst23872 (P3_SUB_357_1258_U475, P3_SUB_357_1258_U473, P3_SUB_357_1258_U474);
  nand ginst23873 (P3_SUB_357_1258_U476, P3_SUB_357_1258_U148, P3_SUB_357_1258_U149);
  nand ginst23874 (P3_SUB_357_1258_U477, P3_SUB_357_1258_U289, P3_SUB_357_1258_U475);
  nand ginst23875 (P3_SUB_357_1258_U478, P3_INSTADDRPOINTER_REG_10__SCAN_IN, P3_SUB_357_1258_U39);
  nand ginst23876 (P3_SUB_357_1258_U479, P3_ADD_357_U6, P3_SUB_357_1258_U53);
  not ginst23877 (P3_SUB_357_1258_U48, P3_INSTADDRPOINTER_REG_21__SCAN_IN);
  nand ginst23878 (P3_SUB_357_1258_U480, P3_SUB_357_1258_U478, P3_SUB_357_1258_U479);
  nand ginst23879 (P3_SUB_357_1258_U481, P3_SUB_357_1258_U150, P3_SUB_357_1258_U265);
  nand ginst23880 (P3_SUB_357_1258_U482, P3_SUB_357_1258_U287, P3_SUB_357_1258_U480);
  nand ginst23881 (P3_SUB_357_1258_U483, P3_INSTADDRPOINTER_REG_0__SCAN_IN, P3_SUB_357_1258_U28);
  nand ginst23882 (P3_SUB_357_1258_U484, P3_ADD_357_U10, P3_SUB_357_1258_U29);
  not ginst23883 (P3_SUB_357_1258_U49, P3_INSTADDRPOINTER_REG_18__SCAN_IN);
  and ginst23884 (P3_SUB_357_1258_U5, P3_SUB_357_1258_U186, P3_SUB_357_1258_U188);
  not ginst23885 (P3_SUB_357_1258_U50, P3_INSTADDRPOINTER_REG_12__SCAN_IN);
  not ginst23886 (P3_SUB_357_1258_U51, P3_INSTADDRPOINTER_REG_13__SCAN_IN);
  not ginst23887 (P3_SUB_357_1258_U52, P3_INSTADDRPOINTER_REG_11__SCAN_IN);
  not ginst23888 (P3_SUB_357_1258_U53, P3_INSTADDRPOINTER_REG_10__SCAN_IN);
  not ginst23889 (P3_SUB_357_1258_U54, P3_INSTADDRPOINTER_REG_14__SCAN_IN);
  not ginst23890 (P3_SUB_357_1258_U55, P3_INSTADDRPOINTER_REG_15__SCAN_IN);
  not ginst23891 (P3_SUB_357_1258_U56, P3_INSTADDRPOINTER_REG_16__SCAN_IN);
  nand ginst23892 (P3_SUB_357_1258_U57, P3_INSTADDRPOINTER_REG_19__SCAN_IN, P3_INSTADDRPOINTER_REG_20__SCAN_IN);
  not ginst23893 (P3_SUB_357_1258_U58, P3_INSTADDRPOINTER_REG_27__SCAN_IN);
  not ginst23894 (P3_SUB_357_1258_U59, P3_INSTADDRPOINTER_REG_29__SCAN_IN);
  and ginst23895 (P3_SUB_357_1258_U6, P3_SUB_357_1258_U178, P3_SUB_357_1258_U187);
  not ginst23896 (P3_SUB_357_1258_U60, P3_INSTADDRPOINTER_REG_30__SCAN_IN);
  nand ginst23897 (P3_SUB_357_1258_U61, P3_SUB_357_1258_U151, P3_SUB_357_1258_U222, P3_SUB_357_1258_U269);
  nand ginst23898 (P3_SUB_357_1258_U62, P3_SUB_357_1258_U105, P3_SUB_357_1258_U218);
  nand ginst23899 (P3_SUB_357_1258_U63, P3_SUB_357_1258_U104, P3_SUB_357_1258_U284);
  nand ginst23900 (P3_SUB_357_1258_U64, P3_SUB_357_1258_U205, P3_SUB_357_1258_U276);
  nand ginst23901 (P3_SUB_357_1258_U65, P3_SUB_357_1258_U277, P3_SUB_357_1258_U47);
  nand ginst23902 (P3_SUB_357_1258_U66, P3_SUB_357_1258_U161, P3_SUB_357_U7);
  nand ginst23903 (P3_SUB_357_1258_U67, P3_SUB_357_1258_U102, P3_SUB_357_1258_U198);
  nand ginst23904 (P3_SUB_357_1258_U68, P3_SUB_357_1258_U290, P3_SUB_357_1258_U8);
  nand ginst23905 (P3_SUB_357_1258_U69, P3_SUB_357_1258_U483, P3_SUB_357_1258_U484);
  and ginst23906 (P3_SUB_357_1258_U7, P3_SUB_357_1258_U189, P3_SUB_357_1258_U6);
  nand ginst23907 (P3_SUB_357_1258_U70, P3_SUB_357_1258_U311, P3_SUB_357_1258_U312);
  nand ginst23908 (P3_SUB_357_1258_U71, P3_SUB_357_1258_U318, P3_SUB_357_1258_U319);
  nand ginst23909 (P3_SUB_357_1258_U72, P3_SUB_357_1258_U325, P3_SUB_357_1258_U326);
  nand ginst23910 (P3_SUB_357_1258_U73, P3_SUB_357_1258_U332, P3_SUB_357_1258_U333);
  nand ginst23911 (P3_SUB_357_1258_U74, P3_SUB_357_1258_U339, P3_SUB_357_1258_U340);
  nand ginst23912 (P3_SUB_357_1258_U75, P3_SUB_357_1258_U344, P3_SUB_357_1258_U345);
  nand ginst23913 (P3_SUB_357_1258_U76, P3_SUB_357_1258_U349, P3_SUB_357_1258_U350);
  nand ginst23914 (P3_SUB_357_1258_U77, P3_SUB_357_1258_U360, P3_SUB_357_1258_U361);
  nand ginst23915 (P3_SUB_357_1258_U78, P3_SUB_357_1258_U365, P3_SUB_357_1258_U366);
  nand ginst23916 (P3_SUB_357_1258_U79, P3_SUB_357_1258_U372, P3_SUB_357_1258_U373);
  and ginst23917 (P3_SUB_357_1258_U8, P3_SUB_357_1258_U190, P3_SUB_357_1258_U5);
  nand ginst23918 (P3_SUB_357_1258_U80, P3_SUB_357_1258_U383, P3_SUB_357_1258_U384);
  nand ginst23919 (P3_SUB_357_1258_U81, P3_SUB_357_1258_U390, P3_SUB_357_1258_U391);
  nand ginst23920 (P3_SUB_357_1258_U82, P3_SUB_357_1258_U397, P3_SUB_357_1258_U398);
  nand ginst23921 (P3_SUB_357_1258_U83, P3_SUB_357_1258_U404, P3_SUB_357_1258_U405);
  nand ginst23922 (P3_SUB_357_1258_U84, P3_SUB_357_1258_U411, P3_SUB_357_1258_U412);
  nand ginst23923 (P3_SUB_357_1258_U85, P3_SUB_357_1258_U418, P3_SUB_357_1258_U419);
  nand ginst23924 (P3_SUB_357_1258_U86, P3_SUB_357_1258_U430, P3_SUB_357_1258_U431);
  nand ginst23925 (P3_SUB_357_1258_U87, P3_SUB_357_1258_U437, P3_SUB_357_1258_U438);
  nand ginst23926 (P3_SUB_357_1258_U88, P3_SUB_357_1258_U448, P3_SUB_357_1258_U449);
  nand ginst23927 (P3_SUB_357_1258_U89, P3_SUB_357_1258_U455, P3_SUB_357_1258_U456);
  and ginst23928 (P3_SUB_357_1258_U9, P3_SUB_357_1258_U204, P3_SUB_357_1258_U209);
  nand ginst23929 (P3_SUB_357_1258_U90, P3_SUB_357_1258_U462, P3_SUB_357_1258_U463);
  nand ginst23930 (P3_SUB_357_1258_U91, P3_SUB_357_1258_U469, P3_SUB_357_1258_U470);
  nand ginst23931 (P3_SUB_357_1258_U92, P3_SUB_357_1258_U476, P3_SUB_357_1258_U477);
  nand ginst23932 (P3_SUB_357_1258_U93, P3_SUB_357_1258_U481, P3_SUB_357_1258_U482);
  and ginst23933 (P3_SUB_357_1258_U94, P3_SUB_357_1258_U160, P3_SUB_357_1258_U163, P3_SUB_357_1258_U164);
  and ginst23934 (P3_SUB_357_1258_U95, P3_INSTADDRPOINTER_REG_3__SCAN_IN, P3_ADD_357_U7);
  and ginst23935 (P3_SUB_357_1258_U96, P3_SUB_357_1258_U162, P3_SUB_357_1258_U168);
  and ginst23936 (P3_SUB_357_1258_U97, P3_SUB_357_1258_U163, P3_SUB_357_1258_U164);
  and ginst23937 (P3_SUB_357_1258_U98, P3_SUB_357_1258_U154, P3_SUB_357_1258_U7);
  and ginst23938 (P3_SUB_357_1258_U99, P3_SUB_357_1258_U155, P3_SUB_357_1258_U192);
  not ginst23939 (P3_SUB_357_U10, P3_U2621);
  not ginst23940 (P3_SUB_357_U11, P3_U2624);
  not ginst23941 (P3_SUB_357_U12, P3_U2623);
  not ginst23942 (P3_SUB_357_U13, P3_U2625);
  not ginst23943 (P3_SUB_357_U6, P3_U2627);
  not ginst23944 (P3_SUB_357_U7, P3_U2622);
  not ginst23945 (P3_SUB_357_U8, P3_U2628);
  not ginst23946 (P3_SUB_357_U9, P3_U2626);
  not ginst23947 (P3_SUB_370_U10, P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN);
  not ginst23948 (P3_SUB_370_U11, P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN);
  not ginst23949 (P3_SUB_370_U12, P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN);
  not ginst23950 (P3_SUB_370_U13, P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN);
  not ginst23951 (P3_SUB_370_U14, P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN);
  not ginst23952 (P3_SUB_370_U15, P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN);
  nand ginst23953 (P3_SUB_370_U16, P3_SUB_370_U40, P3_SUB_370_U41);
  not ginst23954 (P3_SUB_370_U17, P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN);
  not ginst23955 (P3_SUB_370_U18, P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN);
  nand ginst23956 (P3_SUB_370_U19, P3_SUB_370_U50, P3_SUB_370_U51);
  nand ginst23957 (P3_SUB_370_U20, P3_SUB_370_U55, P3_SUB_370_U56);
  nand ginst23958 (P3_SUB_370_U21, P3_SUB_370_U60, P3_SUB_370_U61);
  nand ginst23959 (P3_SUB_370_U22, P3_SUB_370_U65, P3_SUB_370_U66);
  nand ginst23960 (P3_SUB_370_U23, P3_SUB_370_U47, P3_SUB_370_U48);
  nand ginst23961 (P3_SUB_370_U24, P3_SUB_370_U52, P3_SUB_370_U53);
  nand ginst23962 (P3_SUB_370_U25, P3_SUB_370_U57, P3_SUB_370_U58);
  nand ginst23963 (P3_SUB_370_U26, P3_SUB_370_U62, P3_SUB_370_U63);
  nand ginst23964 (P3_SUB_370_U27, P3_SUB_370_U36, P3_SUB_370_U37);
  nand ginst23965 (P3_SUB_370_U28, P3_SUB_370_U32, P3_SUB_370_U33);
  not ginst23966 (P3_SUB_370_U29, P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN);
  not ginst23967 (P3_SUB_370_U30, P3_SUB_370_U9);
  nand ginst23968 (P3_SUB_370_U31, P3_SUB_370_U10, P3_SUB_370_U30);
  nand ginst23969 (P3_SUB_370_U32, P3_SUB_370_U29, P3_SUB_370_U31);
  nand ginst23970 (P3_SUB_370_U33, P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN, P3_SUB_370_U9);
  not ginst23971 (P3_SUB_370_U34, P3_SUB_370_U28);
  nand ginst23972 (P3_SUB_370_U35, P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN, P3_SUB_370_U12);
  nand ginst23973 (P3_SUB_370_U36, P3_SUB_370_U28, P3_SUB_370_U35);
  nand ginst23974 (P3_SUB_370_U37, P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN, P3_SUB_370_U11);
  not ginst23975 (P3_SUB_370_U38, P3_SUB_370_U27);
  nand ginst23976 (P3_SUB_370_U39, P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P3_SUB_370_U14);
  nand ginst23977 (P3_SUB_370_U40, P3_SUB_370_U27, P3_SUB_370_U39);
  nand ginst23978 (P3_SUB_370_U41, P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN, P3_SUB_370_U13);
  not ginst23979 (P3_SUB_370_U42, P3_SUB_370_U16);
  nand ginst23980 (P3_SUB_370_U43, P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN, P3_SUB_370_U17);
  nand ginst23981 (P3_SUB_370_U44, P3_SUB_370_U42, P3_SUB_370_U43);
  nand ginst23982 (P3_SUB_370_U45, P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN, P3_SUB_370_U15);
  nand ginst23983 (P3_SUB_370_U46, P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P3_SUB_370_U8);
  nand ginst23984 (P3_SUB_370_U47, P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN, P3_SUB_370_U15);
  nand ginst23985 (P3_SUB_370_U48, P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN, P3_SUB_370_U17);
  not ginst23986 (P3_SUB_370_U49, P3_SUB_370_U23);
  nand ginst23987 (P3_SUB_370_U50, P3_SUB_370_U42, P3_SUB_370_U49);
  nand ginst23988 (P3_SUB_370_U51, P3_SUB_370_U16, P3_SUB_370_U23);
  nand ginst23989 (P3_SUB_370_U52, P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P3_SUB_370_U14);
  nand ginst23990 (P3_SUB_370_U53, P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN, P3_SUB_370_U13);
  not ginst23991 (P3_SUB_370_U54, P3_SUB_370_U24);
  nand ginst23992 (P3_SUB_370_U55, P3_SUB_370_U38, P3_SUB_370_U54);
  nand ginst23993 (P3_SUB_370_U56, P3_SUB_370_U24, P3_SUB_370_U27);
  nand ginst23994 (P3_SUB_370_U57, P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN, P3_SUB_370_U12);
  nand ginst23995 (P3_SUB_370_U58, P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN, P3_SUB_370_U11);
  not ginst23996 (P3_SUB_370_U59, P3_SUB_370_U25);
  nand ginst23997 (P3_SUB_370_U6, P3_SUB_370_U44, P3_SUB_370_U45);
  nand ginst23998 (P3_SUB_370_U60, P3_SUB_370_U34, P3_SUB_370_U59);
  nand ginst23999 (P3_SUB_370_U61, P3_SUB_370_U25, P3_SUB_370_U28);
  nand ginst24000 (P3_SUB_370_U62, P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P3_SUB_370_U10);
  nand ginst24001 (P3_SUB_370_U63, P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN, P3_SUB_370_U29);
  not ginst24002 (P3_SUB_370_U64, P3_SUB_370_U26);
  nand ginst24003 (P3_SUB_370_U65, P3_SUB_370_U30, P3_SUB_370_U64);
  nand ginst24004 (P3_SUB_370_U66, P3_SUB_370_U26, P3_SUB_370_U9);
  nand ginst24005 (P3_SUB_370_U7, P3_SUB_370_U46, P3_SUB_370_U9);
  not ginst24006 (P3_SUB_370_U8, P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN);
  nand ginst24007 (P3_SUB_370_U9, P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN, P3_SUB_370_U18);
  not ginst24008 (P3_SUB_390_U10, P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN);
  not ginst24009 (P3_SUB_390_U11, P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN);
  not ginst24010 (P3_SUB_390_U12, P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN);
  not ginst24011 (P3_SUB_390_U13, P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN);
  not ginst24012 (P3_SUB_390_U14, P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN);
  not ginst24013 (P3_SUB_390_U15, P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN);
  nand ginst24014 (P3_SUB_390_U16, P3_SUB_390_U40, P3_SUB_390_U41);
  not ginst24015 (P3_SUB_390_U17, P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN);
  not ginst24016 (P3_SUB_390_U18, P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN);
  nand ginst24017 (P3_SUB_390_U19, P3_SUB_390_U50, P3_SUB_390_U51);
  nand ginst24018 (P3_SUB_390_U20, P3_SUB_390_U55, P3_SUB_390_U56);
  nand ginst24019 (P3_SUB_390_U21, P3_SUB_390_U60, P3_SUB_390_U61);
  nand ginst24020 (P3_SUB_390_U22, P3_SUB_390_U65, P3_SUB_390_U66);
  nand ginst24021 (P3_SUB_390_U23, P3_SUB_390_U47, P3_SUB_390_U48);
  nand ginst24022 (P3_SUB_390_U24, P3_SUB_390_U52, P3_SUB_390_U53);
  nand ginst24023 (P3_SUB_390_U25, P3_SUB_390_U57, P3_SUB_390_U58);
  nand ginst24024 (P3_SUB_390_U26, P3_SUB_390_U62, P3_SUB_390_U63);
  nand ginst24025 (P3_SUB_390_U27, P3_SUB_390_U36, P3_SUB_390_U37);
  nand ginst24026 (P3_SUB_390_U28, P3_SUB_390_U32, P3_SUB_390_U33);
  not ginst24027 (P3_SUB_390_U29, P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN);
  not ginst24028 (P3_SUB_390_U30, P3_SUB_390_U9);
  nand ginst24029 (P3_SUB_390_U31, P3_SUB_390_U10, P3_SUB_390_U30);
  nand ginst24030 (P3_SUB_390_U32, P3_SUB_390_U29, P3_SUB_390_U31);
  nand ginst24031 (P3_SUB_390_U33, P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN, P3_SUB_390_U9);
  not ginst24032 (P3_SUB_390_U34, P3_SUB_390_U28);
  nand ginst24033 (P3_SUB_390_U35, P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN, P3_SUB_390_U12);
  nand ginst24034 (P3_SUB_390_U36, P3_SUB_390_U28, P3_SUB_390_U35);
  nand ginst24035 (P3_SUB_390_U37, P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN, P3_SUB_390_U11);
  not ginst24036 (P3_SUB_390_U38, P3_SUB_390_U27);
  nand ginst24037 (P3_SUB_390_U39, P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P3_SUB_390_U14);
  nand ginst24038 (P3_SUB_390_U40, P3_SUB_390_U27, P3_SUB_390_U39);
  nand ginst24039 (P3_SUB_390_U41, P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN, P3_SUB_390_U13);
  not ginst24040 (P3_SUB_390_U42, P3_SUB_390_U16);
  nand ginst24041 (P3_SUB_390_U43, P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN, P3_SUB_390_U17);
  nand ginst24042 (P3_SUB_390_U44, P3_SUB_390_U42, P3_SUB_390_U43);
  nand ginst24043 (P3_SUB_390_U45, P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN, P3_SUB_390_U15);
  nand ginst24044 (P3_SUB_390_U46, P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P3_SUB_390_U8);
  nand ginst24045 (P3_SUB_390_U47, P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN, P3_SUB_390_U15);
  nand ginst24046 (P3_SUB_390_U48, P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN, P3_SUB_390_U17);
  not ginst24047 (P3_SUB_390_U49, P3_SUB_390_U23);
  nand ginst24048 (P3_SUB_390_U50, P3_SUB_390_U42, P3_SUB_390_U49);
  nand ginst24049 (P3_SUB_390_U51, P3_SUB_390_U16, P3_SUB_390_U23);
  nand ginst24050 (P3_SUB_390_U52, P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P3_SUB_390_U14);
  nand ginst24051 (P3_SUB_390_U53, P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN, P3_SUB_390_U13);
  not ginst24052 (P3_SUB_390_U54, P3_SUB_390_U24);
  nand ginst24053 (P3_SUB_390_U55, P3_SUB_390_U38, P3_SUB_390_U54);
  nand ginst24054 (P3_SUB_390_U56, P3_SUB_390_U24, P3_SUB_390_U27);
  nand ginst24055 (P3_SUB_390_U57, P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN, P3_SUB_390_U12);
  nand ginst24056 (P3_SUB_390_U58, P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN, P3_SUB_390_U11);
  not ginst24057 (P3_SUB_390_U59, P3_SUB_390_U25);
  nand ginst24058 (P3_SUB_390_U6, P3_SUB_390_U44, P3_SUB_390_U45);
  nand ginst24059 (P3_SUB_390_U60, P3_SUB_390_U34, P3_SUB_390_U59);
  nand ginst24060 (P3_SUB_390_U61, P3_SUB_390_U25, P3_SUB_390_U28);
  nand ginst24061 (P3_SUB_390_U62, P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P3_SUB_390_U10);
  nand ginst24062 (P3_SUB_390_U63, P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN, P3_SUB_390_U29);
  not ginst24063 (P3_SUB_390_U64, P3_SUB_390_U26);
  nand ginst24064 (P3_SUB_390_U65, P3_SUB_390_U30, P3_SUB_390_U64);
  nand ginst24065 (P3_SUB_390_U66, P3_SUB_390_U26, P3_SUB_390_U9);
  nand ginst24066 (P3_SUB_390_U7, P3_SUB_390_U46, P3_SUB_390_U9);
  not ginst24067 (P3_SUB_390_U8, P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN);
  nand ginst24068 (P3_SUB_390_U9, P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN, P3_SUB_390_U18);
  not ginst24069 (P3_SUB_401_U10, P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN);
  not ginst24070 (P3_SUB_401_U11, P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN);
  not ginst24071 (P3_SUB_401_U12, P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN);
  not ginst24072 (P3_SUB_401_U13, P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN);
  not ginst24073 (P3_SUB_401_U14, P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN);
  not ginst24074 (P3_SUB_401_U15, P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN);
  nand ginst24075 (P3_SUB_401_U16, P3_SUB_401_U40, P3_SUB_401_U41);
  not ginst24076 (P3_SUB_401_U17, P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN);
  not ginst24077 (P3_SUB_401_U18, P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN);
  nand ginst24078 (P3_SUB_401_U19, P3_SUB_401_U50, P3_SUB_401_U51);
  nand ginst24079 (P3_SUB_401_U20, P3_SUB_401_U55, P3_SUB_401_U56);
  nand ginst24080 (P3_SUB_401_U21, P3_SUB_401_U60, P3_SUB_401_U61);
  nand ginst24081 (P3_SUB_401_U22, P3_SUB_401_U65, P3_SUB_401_U66);
  nand ginst24082 (P3_SUB_401_U23, P3_SUB_401_U47, P3_SUB_401_U48);
  nand ginst24083 (P3_SUB_401_U24, P3_SUB_401_U52, P3_SUB_401_U53);
  nand ginst24084 (P3_SUB_401_U25, P3_SUB_401_U57, P3_SUB_401_U58);
  nand ginst24085 (P3_SUB_401_U26, P3_SUB_401_U62, P3_SUB_401_U63);
  nand ginst24086 (P3_SUB_401_U27, P3_SUB_401_U36, P3_SUB_401_U37);
  nand ginst24087 (P3_SUB_401_U28, P3_SUB_401_U32, P3_SUB_401_U33);
  not ginst24088 (P3_SUB_401_U29, P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN);
  not ginst24089 (P3_SUB_401_U30, P3_SUB_401_U9);
  nand ginst24090 (P3_SUB_401_U31, P3_SUB_401_U10, P3_SUB_401_U30);
  nand ginst24091 (P3_SUB_401_U32, P3_SUB_401_U29, P3_SUB_401_U31);
  nand ginst24092 (P3_SUB_401_U33, P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN, P3_SUB_401_U9);
  not ginst24093 (P3_SUB_401_U34, P3_SUB_401_U28);
  nand ginst24094 (P3_SUB_401_U35, P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN, P3_SUB_401_U12);
  nand ginst24095 (P3_SUB_401_U36, P3_SUB_401_U28, P3_SUB_401_U35);
  nand ginst24096 (P3_SUB_401_U37, P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN, P3_SUB_401_U11);
  not ginst24097 (P3_SUB_401_U38, P3_SUB_401_U27);
  nand ginst24098 (P3_SUB_401_U39, P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P3_SUB_401_U14);
  nand ginst24099 (P3_SUB_401_U40, P3_SUB_401_U27, P3_SUB_401_U39);
  nand ginst24100 (P3_SUB_401_U41, P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN, P3_SUB_401_U13);
  not ginst24101 (P3_SUB_401_U42, P3_SUB_401_U16);
  nand ginst24102 (P3_SUB_401_U43, P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN, P3_SUB_401_U17);
  nand ginst24103 (P3_SUB_401_U44, P3_SUB_401_U42, P3_SUB_401_U43);
  nand ginst24104 (P3_SUB_401_U45, P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN, P3_SUB_401_U15);
  nand ginst24105 (P3_SUB_401_U46, P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P3_SUB_401_U8);
  nand ginst24106 (P3_SUB_401_U47, P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN, P3_SUB_401_U15);
  nand ginst24107 (P3_SUB_401_U48, P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN, P3_SUB_401_U17);
  not ginst24108 (P3_SUB_401_U49, P3_SUB_401_U23);
  nand ginst24109 (P3_SUB_401_U50, P3_SUB_401_U42, P3_SUB_401_U49);
  nand ginst24110 (P3_SUB_401_U51, P3_SUB_401_U16, P3_SUB_401_U23);
  nand ginst24111 (P3_SUB_401_U52, P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P3_SUB_401_U14);
  nand ginst24112 (P3_SUB_401_U53, P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN, P3_SUB_401_U13);
  not ginst24113 (P3_SUB_401_U54, P3_SUB_401_U24);
  nand ginst24114 (P3_SUB_401_U55, P3_SUB_401_U38, P3_SUB_401_U54);
  nand ginst24115 (P3_SUB_401_U56, P3_SUB_401_U24, P3_SUB_401_U27);
  nand ginst24116 (P3_SUB_401_U57, P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN, P3_SUB_401_U12);
  nand ginst24117 (P3_SUB_401_U58, P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN, P3_SUB_401_U11);
  not ginst24118 (P3_SUB_401_U59, P3_SUB_401_U25);
  nand ginst24119 (P3_SUB_401_U6, P3_SUB_401_U44, P3_SUB_401_U45);
  nand ginst24120 (P3_SUB_401_U60, P3_SUB_401_U34, P3_SUB_401_U59);
  nand ginst24121 (P3_SUB_401_U61, P3_SUB_401_U25, P3_SUB_401_U28);
  nand ginst24122 (P3_SUB_401_U62, P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P3_SUB_401_U10);
  nand ginst24123 (P3_SUB_401_U63, P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN, P3_SUB_401_U29);
  not ginst24124 (P3_SUB_401_U64, P3_SUB_401_U26);
  nand ginst24125 (P3_SUB_401_U65, P3_SUB_401_U30, P3_SUB_401_U64);
  nand ginst24126 (P3_SUB_401_U66, P3_SUB_401_U26, P3_SUB_401_U9);
  nand ginst24127 (P3_SUB_401_U7, P3_SUB_401_U46, P3_SUB_401_U9);
  not ginst24128 (P3_SUB_401_U8, P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN);
  nand ginst24129 (P3_SUB_401_U9, P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN, P3_SUB_401_U18);
  not ginst24130 (P3_SUB_412_U10, P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN);
  not ginst24131 (P3_SUB_412_U11, P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN);
  not ginst24132 (P3_SUB_412_U12, P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN);
  not ginst24133 (P3_SUB_412_U13, P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN);
  nand ginst24134 (P3_SUB_412_U14, P3_SUB_412_U38, P3_SUB_412_U39);
  not ginst24135 (P3_SUB_412_U15, P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN);
  nand ginst24136 (P3_SUB_412_U16, P3_SUB_412_U47, P3_SUB_412_U48);
  nand ginst24137 (P3_SUB_412_U17, P3_SUB_412_U52, P3_SUB_412_U53);
  nand ginst24138 (P3_SUB_412_U18, P3_SUB_412_U57, P3_SUB_412_U58);
  nand ginst24139 (P3_SUB_412_U19, P3_SUB_412_U62, P3_SUB_412_U63);
  nand ginst24140 (P3_SUB_412_U20, P3_SUB_412_U44, P3_SUB_412_U45);
  nand ginst24141 (P3_SUB_412_U21, P3_SUB_412_U49, P3_SUB_412_U50);
  nand ginst24142 (P3_SUB_412_U22, P3_SUB_412_U54, P3_SUB_412_U55);
  nand ginst24143 (P3_SUB_412_U23, P3_SUB_412_U59, P3_SUB_412_U60);
  nand ginst24144 (P3_SUB_412_U24, P3_SUB_412_U34, P3_SUB_412_U35);
  nand ginst24145 (P3_SUB_412_U25, P3_SUB_412_U30, P3_SUB_412_U31);
  not ginst24146 (P3_SUB_412_U26, P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN);
  not ginst24147 (P3_SUB_412_U27, P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN);
  not ginst24148 (P3_SUB_412_U28, P3_SUB_412_U7);
  nand ginst24149 (P3_SUB_412_U29, P3_SUB_412_U28, P3_SUB_412_U8);
  nand ginst24150 (P3_SUB_412_U30, P3_SUB_412_U26, P3_SUB_412_U29);
  nand ginst24151 (P3_SUB_412_U31, P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN, P3_SUB_412_U7);
  not ginst24152 (P3_SUB_412_U32, P3_SUB_412_U25);
  nand ginst24153 (P3_SUB_412_U33, P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN, P3_SUB_412_U10);
  nand ginst24154 (P3_SUB_412_U34, P3_SUB_412_U25, P3_SUB_412_U33);
  nand ginst24155 (P3_SUB_412_U35, P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN, P3_SUB_412_U9);
  not ginst24156 (P3_SUB_412_U36, P3_SUB_412_U24);
  nand ginst24157 (P3_SUB_412_U37, P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P3_SUB_412_U12);
  nand ginst24158 (P3_SUB_412_U38, P3_SUB_412_U24, P3_SUB_412_U37);
  nand ginst24159 (P3_SUB_412_U39, P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN, P3_SUB_412_U11);
  not ginst24160 (P3_SUB_412_U40, P3_SUB_412_U14);
  nand ginst24161 (P3_SUB_412_U41, P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN, P3_SUB_412_U15);
  nand ginst24162 (P3_SUB_412_U42, P3_SUB_412_U40, P3_SUB_412_U41);
  nand ginst24163 (P3_SUB_412_U43, P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN, P3_SUB_412_U13);
  nand ginst24164 (P3_SUB_412_U44, P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN, P3_SUB_412_U13);
  nand ginst24165 (P3_SUB_412_U45, P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN, P3_SUB_412_U15);
  not ginst24166 (P3_SUB_412_U46, P3_SUB_412_U20);
  nand ginst24167 (P3_SUB_412_U47, P3_SUB_412_U40, P3_SUB_412_U46);
  nand ginst24168 (P3_SUB_412_U48, P3_SUB_412_U14, P3_SUB_412_U20);
  nand ginst24169 (P3_SUB_412_U49, P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P3_SUB_412_U12);
  nand ginst24170 (P3_SUB_412_U50, P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN, P3_SUB_412_U11);
  not ginst24171 (P3_SUB_412_U51, P3_SUB_412_U21);
  nand ginst24172 (P3_SUB_412_U52, P3_SUB_412_U36, P3_SUB_412_U51);
  nand ginst24173 (P3_SUB_412_U53, P3_SUB_412_U21, P3_SUB_412_U24);
  nand ginst24174 (P3_SUB_412_U54, P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN, P3_SUB_412_U10);
  nand ginst24175 (P3_SUB_412_U55, P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN, P3_SUB_412_U9);
  not ginst24176 (P3_SUB_412_U56, P3_SUB_412_U22);
  nand ginst24177 (P3_SUB_412_U57, P3_SUB_412_U32, P3_SUB_412_U56);
  nand ginst24178 (P3_SUB_412_U58, P3_SUB_412_U22, P3_SUB_412_U25);
  nand ginst24179 (P3_SUB_412_U59, P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P3_SUB_412_U8);
  nand ginst24180 (P3_SUB_412_U6, P3_SUB_412_U42, P3_SUB_412_U43);
  nand ginst24181 (P3_SUB_412_U60, P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN, P3_SUB_412_U26);
  not ginst24182 (P3_SUB_412_U61, P3_SUB_412_U23);
  nand ginst24183 (P3_SUB_412_U62, P3_SUB_412_U28, P3_SUB_412_U61);
  nand ginst24184 (P3_SUB_412_U63, P3_SUB_412_U23, P3_SUB_412_U7);
  nand ginst24185 (P3_SUB_412_U7, P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN, P3_SUB_412_U27);
  not ginst24186 (P3_SUB_412_U8, P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN);
  not ginst24187 (P3_SUB_412_U9, P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN);
  and ginst24188 (P3_SUB_414_U10, P3_SUB_414_U118, P3_SUB_414_U32);
  not ginst24189 (P3_SUB_414_U100, P3_SUB_414_U35);
  not ginst24190 (P3_SUB_414_U101, P3_SUB_414_U36);
  not ginst24191 (P3_SUB_414_U102, P3_SUB_414_U37);
  not ginst24192 (P3_SUB_414_U103, P3_SUB_414_U38);
  or ginst24193 (P3_SUB_414_U104, P3_EBX_REG_0__SCAN_IN, P3_EBX_REG_1__SCAN_IN);
  nand ginst24194 (P3_SUB_414_U105, P3_EBX_REG_2__SCAN_IN, P3_SUB_414_U104);
  nand ginst24195 (P3_SUB_414_U106, P3_EBX_REG_29__SCAN_IN, P3_SUB_414_U37);
  nand ginst24196 (P3_SUB_414_U107, P3_SUB_414_U101, P3_SUB_414_U63);
  nand ginst24197 (P3_SUB_414_U108, P3_EBX_REG_28__SCAN_IN, P3_SUB_414_U107);
  nand ginst24198 (P3_SUB_414_U109, P3_SUB_414_U100, P3_SUB_414_U65);
  and ginst24199 (P3_SUB_414_U11, P3_SUB_414_U116, P3_SUB_414_U33);
  nand ginst24200 (P3_SUB_414_U110, P3_EBX_REG_26__SCAN_IN, P3_SUB_414_U109);
  nand ginst24201 (P3_SUB_414_U111, P3_SUB_414_U67, P3_SUB_414_U99);
  nand ginst24202 (P3_SUB_414_U112, P3_EBX_REG_24__SCAN_IN, P3_SUB_414_U111);
  nand ginst24203 (P3_SUB_414_U113, P3_SUB_414_U69, P3_SUB_414_U98);
  nand ginst24204 (P3_SUB_414_U114, P3_EBX_REG_22__SCAN_IN, P3_SUB_414_U113);
  nand ginst24205 (P3_SUB_414_U115, P3_SUB_414_U73, P3_SUB_414_U97);
  nand ginst24206 (P3_SUB_414_U116, P3_EBX_REG_20__SCAN_IN, P3_SUB_414_U115);
  nand ginst24207 (P3_SUB_414_U117, P3_SUB_414_U75, P3_SUB_414_U96);
  nand ginst24208 (P3_SUB_414_U118, P3_EBX_REG_18__SCAN_IN, P3_SUB_414_U117);
  nand ginst24209 (P3_SUB_414_U119, P3_SUB_414_U77, P3_SUB_414_U95);
  and ginst24210 (P3_SUB_414_U12, P3_SUB_414_U114, P3_SUB_414_U34);
  nand ginst24211 (P3_SUB_414_U120, P3_EBX_REG_16__SCAN_IN, P3_SUB_414_U119);
  nand ginst24212 (P3_SUB_414_U121, P3_SUB_414_U79, P3_SUB_414_U94);
  nand ginst24213 (P3_SUB_414_U122, P3_EBX_REG_14__SCAN_IN, P3_SUB_414_U121);
  nand ginst24214 (P3_SUB_414_U123, P3_SUB_414_U81, P3_SUB_414_U93);
  nand ginst24215 (P3_SUB_414_U124, P3_EBX_REG_12__SCAN_IN, P3_SUB_414_U123);
  nand ginst24216 (P3_SUB_414_U125, P3_SUB_414_U52, P3_SUB_414_U86);
  nand ginst24217 (P3_SUB_414_U126, P3_EBX_REG_10__SCAN_IN, P3_SUB_414_U125);
  nand ginst24218 (P3_SUB_414_U127, P3_SUB_414_U103, P3_SUB_414_U61);
  nand ginst24219 (P3_SUB_414_U128, P3_EBX_REG_9__SCAN_IN, P3_SUB_414_U24);
  nand ginst24220 (P3_SUB_414_U129, P3_SUB_414_U52, P3_SUB_414_U86);
  and ginst24221 (P3_SUB_414_U13, P3_SUB_414_U112, P3_SUB_414_U35);
  nand ginst24222 (P3_SUB_414_U130, P3_EBX_REG_7__SCAN_IN, P3_SUB_414_U23);
  nand ginst24223 (P3_SUB_414_U131, P3_SUB_414_U54, P3_SUB_414_U85);
  nand ginst24224 (P3_SUB_414_U132, P3_EBX_REG_5__SCAN_IN, P3_SUB_414_U22);
  nand ginst24225 (P3_SUB_414_U133, P3_SUB_414_U56, P3_SUB_414_U84);
  nand ginst24226 (P3_SUB_414_U134, P3_EBX_REG_3__SCAN_IN, P3_SUB_414_U21);
  nand ginst24227 (P3_SUB_414_U135, P3_SUB_414_U58, P3_SUB_414_U83);
  nand ginst24228 (P3_SUB_414_U136, P3_SUB_414_U127, P3_SUB_414_U60);
  nand ginst24229 (P3_SUB_414_U137, P3_EBX_REG_31__SCAN_IN, P3_SUB_414_U103, P3_SUB_414_U61);
  nand ginst24230 (P3_SUB_414_U138, P3_EBX_REG_30__SCAN_IN, P3_SUB_414_U38);
  nand ginst24231 (P3_SUB_414_U139, P3_SUB_414_U103, P3_SUB_414_U61);
  and ginst24232 (P3_SUB_414_U14, P3_SUB_414_U110, P3_SUB_414_U36);
  nand ginst24233 (P3_SUB_414_U140, P3_EBX_REG_27__SCAN_IN, P3_SUB_414_U36);
  nand ginst24234 (P3_SUB_414_U141, P3_SUB_414_U101, P3_SUB_414_U63);
  nand ginst24235 (P3_SUB_414_U142, P3_EBX_REG_25__SCAN_IN, P3_SUB_414_U35);
  nand ginst24236 (P3_SUB_414_U143, P3_SUB_414_U100, P3_SUB_414_U65);
  nand ginst24237 (P3_SUB_414_U144, P3_EBX_REG_23__SCAN_IN, P3_SUB_414_U34);
  nand ginst24238 (P3_SUB_414_U145, P3_SUB_414_U67, P3_SUB_414_U99);
  nand ginst24239 (P3_SUB_414_U146, P3_EBX_REG_21__SCAN_IN, P3_SUB_414_U33);
  nand ginst24240 (P3_SUB_414_U147, P3_SUB_414_U69, P3_SUB_414_U98);
  nand ginst24241 (P3_SUB_414_U148, P3_EBX_REG_1__SCAN_IN, P3_SUB_414_U72);
  nand ginst24242 (P3_SUB_414_U149, P3_EBX_REG_0__SCAN_IN, P3_SUB_414_U71);
  and ginst24243 (P3_SUB_414_U15, P3_SUB_414_U108, P3_SUB_414_U37);
  nand ginst24244 (P3_SUB_414_U150, P3_EBX_REG_19__SCAN_IN, P3_SUB_414_U32);
  nand ginst24245 (P3_SUB_414_U151, P3_SUB_414_U73, P3_SUB_414_U97);
  nand ginst24246 (P3_SUB_414_U152, P3_EBX_REG_17__SCAN_IN, P3_SUB_414_U31);
  nand ginst24247 (P3_SUB_414_U153, P3_SUB_414_U75, P3_SUB_414_U96);
  nand ginst24248 (P3_SUB_414_U154, P3_EBX_REG_15__SCAN_IN, P3_SUB_414_U30);
  nand ginst24249 (P3_SUB_414_U155, P3_SUB_414_U77, P3_SUB_414_U95);
  nand ginst24250 (P3_SUB_414_U156, P3_EBX_REG_13__SCAN_IN, P3_SUB_414_U29);
  nand ginst24251 (P3_SUB_414_U157, P3_SUB_414_U79, P3_SUB_414_U94);
  nand ginst24252 (P3_SUB_414_U158, P3_EBX_REG_11__SCAN_IN, P3_SUB_414_U28);
  nand ginst24253 (P3_SUB_414_U159, P3_SUB_414_U81, P3_SUB_414_U93);
  and ginst24254 (P3_SUB_414_U16, P3_SUB_414_U106, P3_SUB_414_U38);
  and ginst24255 (P3_SUB_414_U17, P3_SUB_414_U105, P3_SUB_414_U21);
  and ginst24256 (P3_SUB_414_U18, P3_SUB_414_U22, P3_SUB_414_U92);
  and ginst24257 (P3_SUB_414_U19, P3_SUB_414_U23, P3_SUB_414_U90);
  and ginst24258 (P3_SUB_414_U20, P3_SUB_414_U24, P3_SUB_414_U88);
  or ginst24259 (P3_SUB_414_U21, P3_EBX_REG_0__SCAN_IN, P3_EBX_REG_1__SCAN_IN, P3_EBX_REG_2__SCAN_IN);
  nand ginst24260 (P3_SUB_414_U22, P3_SUB_414_U27, P3_SUB_414_U58, P3_SUB_414_U83);
  nand ginst24261 (P3_SUB_414_U23, P3_SUB_414_U26, P3_SUB_414_U56, P3_SUB_414_U84);
  nand ginst24262 (P3_SUB_414_U24, P3_SUB_414_U25, P3_SUB_414_U54, P3_SUB_414_U85);
  not ginst24263 (P3_SUB_414_U25, P3_EBX_REG_8__SCAN_IN);
  not ginst24264 (P3_SUB_414_U26, P3_EBX_REG_6__SCAN_IN);
  not ginst24265 (P3_SUB_414_U27, P3_EBX_REG_4__SCAN_IN);
  nand ginst24266 (P3_SUB_414_U28, P3_SUB_414_U49, P3_SUB_414_U52, P3_SUB_414_U86);
  nand ginst24267 (P3_SUB_414_U29, P3_SUB_414_U48, P3_SUB_414_U81, P3_SUB_414_U93);
  nand ginst24268 (P3_SUB_414_U30, P3_SUB_414_U47, P3_SUB_414_U79, P3_SUB_414_U94);
  nand ginst24269 (P3_SUB_414_U31, P3_SUB_414_U46, P3_SUB_414_U77, P3_SUB_414_U95);
  nand ginst24270 (P3_SUB_414_U32, P3_SUB_414_U45, P3_SUB_414_U75, P3_SUB_414_U96);
  nand ginst24271 (P3_SUB_414_U33, P3_SUB_414_U44, P3_SUB_414_U73, P3_SUB_414_U97);
  nand ginst24272 (P3_SUB_414_U34, P3_SUB_414_U43, P3_SUB_414_U69, P3_SUB_414_U98);
  nand ginst24273 (P3_SUB_414_U35, P3_SUB_414_U42, P3_SUB_414_U67, P3_SUB_414_U99);
  nand ginst24274 (P3_SUB_414_U36, P3_SUB_414_U100, P3_SUB_414_U41, P3_SUB_414_U65);
  nand ginst24275 (P3_SUB_414_U37, P3_SUB_414_U101, P3_SUB_414_U40, P3_SUB_414_U63);
  nand ginst24276 (P3_SUB_414_U38, P3_SUB_414_U102, P3_SUB_414_U39);
  not ginst24277 (P3_SUB_414_U39, P3_EBX_REG_29__SCAN_IN);
  not ginst24278 (P3_SUB_414_U40, P3_EBX_REG_28__SCAN_IN);
  not ginst24279 (P3_SUB_414_U41, P3_EBX_REG_26__SCAN_IN);
  not ginst24280 (P3_SUB_414_U42, P3_EBX_REG_24__SCAN_IN);
  not ginst24281 (P3_SUB_414_U43, P3_EBX_REG_22__SCAN_IN);
  not ginst24282 (P3_SUB_414_U44, P3_EBX_REG_20__SCAN_IN);
  not ginst24283 (P3_SUB_414_U45, P3_EBX_REG_18__SCAN_IN);
  not ginst24284 (P3_SUB_414_U46, P3_EBX_REG_16__SCAN_IN);
  not ginst24285 (P3_SUB_414_U47, P3_EBX_REG_14__SCAN_IN);
  not ginst24286 (P3_SUB_414_U48, P3_EBX_REG_12__SCAN_IN);
  not ginst24287 (P3_SUB_414_U49, P3_EBX_REG_10__SCAN_IN);
  nand ginst24288 (P3_SUB_414_U50, P3_SUB_414_U148, P3_SUB_414_U149);
  nand ginst24289 (P3_SUB_414_U51, P3_SUB_414_U136, P3_SUB_414_U137);
  not ginst24290 (P3_SUB_414_U52, P3_EBX_REG_9__SCAN_IN);
  and ginst24291 (P3_SUB_414_U53, P3_SUB_414_U128, P3_SUB_414_U129);
  not ginst24292 (P3_SUB_414_U54, P3_EBX_REG_7__SCAN_IN);
  and ginst24293 (P3_SUB_414_U55, P3_SUB_414_U130, P3_SUB_414_U131);
  not ginst24294 (P3_SUB_414_U56, P3_EBX_REG_5__SCAN_IN);
  and ginst24295 (P3_SUB_414_U57, P3_SUB_414_U132, P3_SUB_414_U133);
  not ginst24296 (P3_SUB_414_U58, P3_EBX_REG_3__SCAN_IN);
  and ginst24297 (P3_SUB_414_U59, P3_SUB_414_U134, P3_SUB_414_U135);
  and ginst24298 (P3_SUB_414_U6, P3_SUB_414_U126, P3_SUB_414_U28);
  not ginst24299 (P3_SUB_414_U60, P3_EBX_REG_31__SCAN_IN);
  not ginst24300 (P3_SUB_414_U61, P3_EBX_REG_30__SCAN_IN);
  and ginst24301 (P3_SUB_414_U62, P3_SUB_414_U138, P3_SUB_414_U139);
  not ginst24302 (P3_SUB_414_U63, P3_EBX_REG_27__SCAN_IN);
  and ginst24303 (P3_SUB_414_U64, P3_SUB_414_U140, P3_SUB_414_U141);
  not ginst24304 (P3_SUB_414_U65, P3_EBX_REG_25__SCAN_IN);
  and ginst24305 (P3_SUB_414_U66, P3_SUB_414_U142, P3_SUB_414_U143);
  not ginst24306 (P3_SUB_414_U67, P3_EBX_REG_23__SCAN_IN);
  and ginst24307 (P3_SUB_414_U68, P3_SUB_414_U144, P3_SUB_414_U145);
  not ginst24308 (P3_SUB_414_U69, P3_EBX_REG_21__SCAN_IN);
  and ginst24309 (P3_SUB_414_U7, P3_SUB_414_U124, P3_SUB_414_U29);
  and ginst24310 (P3_SUB_414_U70, P3_SUB_414_U146, P3_SUB_414_U147);
  not ginst24311 (P3_SUB_414_U71, P3_EBX_REG_1__SCAN_IN);
  not ginst24312 (P3_SUB_414_U72, P3_EBX_REG_0__SCAN_IN);
  not ginst24313 (P3_SUB_414_U73, P3_EBX_REG_19__SCAN_IN);
  and ginst24314 (P3_SUB_414_U74, P3_SUB_414_U150, P3_SUB_414_U151);
  not ginst24315 (P3_SUB_414_U75, P3_EBX_REG_17__SCAN_IN);
  and ginst24316 (P3_SUB_414_U76, P3_SUB_414_U152, P3_SUB_414_U153);
  not ginst24317 (P3_SUB_414_U77, P3_EBX_REG_15__SCAN_IN);
  and ginst24318 (P3_SUB_414_U78, P3_SUB_414_U154, P3_SUB_414_U155);
  not ginst24319 (P3_SUB_414_U79, P3_EBX_REG_13__SCAN_IN);
  and ginst24320 (P3_SUB_414_U8, P3_SUB_414_U122, P3_SUB_414_U30);
  and ginst24321 (P3_SUB_414_U80, P3_SUB_414_U156, P3_SUB_414_U157);
  not ginst24322 (P3_SUB_414_U81, P3_EBX_REG_11__SCAN_IN);
  and ginst24323 (P3_SUB_414_U82, P3_SUB_414_U158, P3_SUB_414_U159);
  not ginst24324 (P3_SUB_414_U83, P3_SUB_414_U21);
  not ginst24325 (P3_SUB_414_U84, P3_SUB_414_U22);
  not ginst24326 (P3_SUB_414_U85, P3_SUB_414_U23);
  not ginst24327 (P3_SUB_414_U86, P3_SUB_414_U24);
  nand ginst24328 (P3_SUB_414_U87, P3_SUB_414_U54, P3_SUB_414_U85);
  nand ginst24329 (P3_SUB_414_U88, P3_EBX_REG_8__SCAN_IN, P3_SUB_414_U87);
  nand ginst24330 (P3_SUB_414_U89, P3_SUB_414_U56, P3_SUB_414_U84);
  and ginst24331 (P3_SUB_414_U9, P3_SUB_414_U120, P3_SUB_414_U31);
  nand ginst24332 (P3_SUB_414_U90, P3_EBX_REG_6__SCAN_IN, P3_SUB_414_U89);
  nand ginst24333 (P3_SUB_414_U91, P3_SUB_414_U58, P3_SUB_414_U83);
  nand ginst24334 (P3_SUB_414_U92, P3_EBX_REG_4__SCAN_IN, P3_SUB_414_U91);
  not ginst24335 (P3_SUB_414_U93, P3_SUB_414_U28);
  not ginst24336 (P3_SUB_414_U94, P3_SUB_414_U29);
  not ginst24337 (P3_SUB_414_U95, P3_SUB_414_U30);
  not ginst24338 (P3_SUB_414_U96, P3_SUB_414_U31);
  not ginst24339 (P3_SUB_414_U97, P3_SUB_414_U32);
  not ginst24340 (P3_SUB_414_U98, P3_SUB_414_U33);
  not ginst24341 (P3_SUB_414_U99, P3_SUB_414_U34);
  not ginst24342 (P3_SUB_450_U10, P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN);
  not ginst24343 (P3_SUB_450_U11, P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN);
  not ginst24344 (P3_SUB_450_U12, P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN);
  not ginst24345 (P3_SUB_450_U13, P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN);
  nand ginst24346 (P3_SUB_450_U14, P3_SUB_450_U38, P3_SUB_450_U39);
  not ginst24347 (P3_SUB_450_U15, P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN);
  nand ginst24348 (P3_SUB_450_U16, P3_SUB_450_U47, P3_SUB_450_U48);
  nand ginst24349 (P3_SUB_450_U17, P3_SUB_450_U52, P3_SUB_450_U53);
  nand ginst24350 (P3_SUB_450_U18, P3_SUB_450_U57, P3_SUB_450_U58);
  nand ginst24351 (P3_SUB_450_U19, P3_SUB_450_U62, P3_SUB_450_U63);
  nand ginst24352 (P3_SUB_450_U20, P3_SUB_450_U44, P3_SUB_450_U45);
  nand ginst24353 (P3_SUB_450_U21, P3_SUB_450_U49, P3_SUB_450_U50);
  nand ginst24354 (P3_SUB_450_U22, P3_SUB_450_U54, P3_SUB_450_U55);
  nand ginst24355 (P3_SUB_450_U23, P3_SUB_450_U59, P3_SUB_450_U60);
  nand ginst24356 (P3_SUB_450_U24, P3_SUB_450_U34, P3_SUB_450_U35);
  nand ginst24357 (P3_SUB_450_U25, P3_SUB_450_U30, P3_SUB_450_U31);
  not ginst24358 (P3_SUB_450_U26, P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN);
  not ginst24359 (P3_SUB_450_U27, P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN);
  not ginst24360 (P3_SUB_450_U28, P3_SUB_450_U7);
  nand ginst24361 (P3_SUB_450_U29, P3_SUB_450_U28, P3_SUB_450_U8);
  nand ginst24362 (P3_SUB_450_U30, P3_SUB_450_U26, P3_SUB_450_U29);
  nand ginst24363 (P3_SUB_450_U31, P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN, P3_SUB_450_U7);
  not ginst24364 (P3_SUB_450_U32, P3_SUB_450_U25);
  nand ginst24365 (P3_SUB_450_U33, P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN, P3_SUB_450_U10);
  nand ginst24366 (P3_SUB_450_U34, P3_SUB_450_U25, P3_SUB_450_U33);
  nand ginst24367 (P3_SUB_450_U35, P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN, P3_SUB_450_U9);
  not ginst24368 (P3_SUB_450_U36, P3_SUB_450_U24);
  nand ginst24369 (P3_SUB_450_U37, P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P3_SUB_450_U12);
  nand ginst24370 (P3_SUB_450_U38, P3_SUB_450_U24, P3_SUB_450_U37);
  nand ginst24371 (P3_SUB_450_U39, P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN, P3_SUB_450_U11);
  not ginst24372 (P3_SUB_450_U40, P3_SUB_450_U14);
  nand ginst24373 (P3_SUB_450_U41, P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN, P3_SUB_450_U15);
  nand ginst24374 (P3_SUB_450_U42, P3_SUB_450_U40, P3_SUB_450_U41);
  nand ginst24375 (P3_SUB_450_U43, P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN, P3_SUB_450_U13);
  nand ginst24376 (P3_SUB_450_U44, P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN, P3_SUB_450_U13);
  nand ginst24377 (P3_SUB_450_U45, P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN, P3_SUB_450_U15);
  not ginst24378 (P3_SUB_450_U46, P3_SUB_450_U20);
  nand ginst24379 (P3_SUB_450_U47, P3_SUB_450_U40, P3_SUB_450_U46);
  nand ginst24380 (P3_SUB_450_U48, P3_SUB_450_U14, P3_SUB_450_U20);
  nand ginst24381 (P3_SUB_450_U49, P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P3_SUB_450_U12);
  nand ginst24382 (P3_SUB_450_U50, P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN, P3_SUB_450_U11);
  not ginst24383 (P3_SUB_450_U51, P3_SUB_450_U21);
  nand ginst24384 (P3_SUB_450_U52, P3_SUB_450_U36, P3_SUB_450_U51);
  nand ginst24385 (P3_SUB_450_U53, P3_SUB_450_U21, P3_SUB_450_U24);
  nand ginst24386 (P3_SUB_450_U54, P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN, P3_SUB_450_U10);
  nand ginst24387 (P3_SUB_450_U55, P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN, P3_SUB_450_U9);
  not ginst24388 (P3_SUB_450_U56, P3_SUB_450_U22);
  nand ginst24389 (P3_SUB_450_U57, P3_SUB_450_U32, P3_SUB_450_U56);
  nand ginst24390 (P3_SUB_450_U58, P3_SUB_450_U22, P3_SUB_450_U25);
  nand ginst24391 (P3_SUB_450_U59, P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P3_SUB_450_U8);
  nand ginst24392 (P3_SUB_450_U6, P3_SUB_450_U42, P3_SUB_450_U43);
  nand ginst24393 (P3_SUB_450_U60, P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN, P3_SUB_450_U26);
  not ginst24394 (P3_SUB_450_U61, P3_SUB_450_U23);
  nand ginst24395 (P3_SUB_450_U62, P3_SUB_450_U28, P3_SUB_450_U61);
  nand ginst24396 (P3_SUB_450_U63, P3_SUB_450_U23, P3_SUB_450_U7);
  nand ginst24397 (P3_SUB_450_U7, P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN, P3_SUB_450_U27);
  not ginst24398 (P3_SUB_450_U8, P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN);
  not ginst24399 (P3_SUB_450_U9, P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN);
  not ginst24400 (P3_SUB_485_U10, P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN);
  not ginst24401 (P3_SUB_485_U11, P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN);
  not ginst24402 (P3_SUB_485_U12, P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN);
  not ginst24403 (P3_SUB_485_U13, P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN);
  nand ginst24404 (P3_SUB_485_U14, P3_SUB_485_U38, P3_SUB_485_U39);
  not ginst24405 (P3_SUB_485_U15, P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN);
  nand ginst24406 (P3_SUB_485_U16, P3_SUB_485_U47, P3_SUB_485_U48);
  nand ginst24407 (P3_SUB_485_U17, P3_SUB_485_U52, P3_SUB_485_U53);
  nand ginst24408 (P3_SUB_485_U18, P3_SUB_485_U57, P3_SUB_485_U58);
  nand ginst24409 (P3_SUB_485_U19, P3_SUB_485_U62, P3_SUB_485_U63);
  nand ginst24410 (P3_SUB_485_U20, P3_SUB_485_U44, P3_SUB_485_U45);
  nand ginst24411 (P3_SUB_485_U21, P3_SUB_485_U49, P3_SUB_485_U50);
  nand ginst24412 (P3_SUB_485_U22, P3_SUB_485_U54, P3_SUB_485_U55);
  nand ginst24413 (P3_SUB_485_U23, P3_SUB_485_U59, P3_SUB_485_U60);
  nand ginst24414 (P3_SUB_485_U24, P3_SUB_485_U34, P3_SUB_485_U35);
  nand ginst24415 (P3_SUB_485_U25, P3_SUB_485_U30, P3_SUB_485_U31);
  not ginst24416 (P3_SUB_485_U26, P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN);
  not ginst24417 (P3_SUB_485_U27, P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN);
  not ginst24418 (P3_SUB_485_U28, P3_SUB_485_U7);
  nand ginst24419 (P3_SUB_485_U29, P3_SUB_485_U28, P3_SUB_485_U8);
  nand ginst24420 (P3_SUB_485_U30, P3_SUB_485_U26, P3_SUB_485_U29);
  nand ginst24421 (P3_SUB_485_U31, P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN, P3_SUB_485_U7);
  not ginst24422 (P3_SUB_485_U32, P3_SUB_485_U25);
  nand ginst24423 (P3_SUB_485_U33, P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN, P3_SUB_485_U10);
  nand ginst24424 (P3_SUB_485_U34, P3_SUB_485_U25, P3_SUB_485_U33);
  nand ginst24425 (P3_SUB_485_U35, P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN, P3_SUB_485_U9);
  not ginst24426 (P3_SUB_485_U36, P3_SUB_485_U24);
  nand ginst24427 (P3_SUB_485_U37, P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P3_SUB_485_U12);
  nand ginst24428 (P3_SUB_485_U38, P3_SUB_485_U24, P3_SUB_485_U37);
  nand ginst24429 (P3_SUB_485_U39, P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN, P3_SUB_485_U11);
  not ginst24430 (P3_SUB_485_U40, P3_SUB_485_U14);
  nand ginst24431 (P3_SUB_485_U41, P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN, P3_SUB_485_U15);
  nand ginst24432 (P3_SUB_485_U42, P3_SUB_485_U40, P3_SUB_485_U41);
  nand ginst24433 (P3_SUB_485_U43, P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN, P3_SUB_485_U13);
  nand ginst24434 (P3_SUB_485_U44, P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN, P3_SUB_485_U13);
  nand ginst24435 (P3_SUB_485_U45, P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN, P3_SUB_485_U15);
  not ginst24436 (P3_SUB_485_U46, P3_SUB_485_U20);
  nand ginst24437 (P3_SUB_485_U47, P3_SUB_485_U40, P3_SUB_485_U46);
  nand ginst24438 (P3_SUB_485_U48, P3_SUB_485_U14, P3_SUB_485_U20);
  nand ginst24439 (P3_SUB_485_U49, P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P3_SUB_485_U12);
  nand ginst24440 (P3_SUB_485_U50, P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN, P3_SUB_485_U11);
  not ginst24441 (P3_SUB_485_U51, P3_SUB_485_U21);
  nand ginst24442 (P3_SUB_485_U52, P3_SUB_485_U36, P3_SUB_485_U51);
  nand ginst24443 (P3_SUB_485_U53, P3_SUB_485_U21, P3_SUB_485_U24);
  nand ginst24444 (P3_SUB_485_U54, P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN, P3_SUB_485_U10);
  nand ginst24445 (P3_SUB_485_U55, P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN, P3_SUB_485_U9);
  not ginst24446 (P3_SUB_485_U56, P3_SUB_485_U22);
  nand ginst24447 (P3_SUB_485_U57, P3_SUB_485_U32, P3_SUB_485_U56);
  nand ginst24448 (P3_SUB_485_U58, P3_SUB_485_U22, P3_SUB_485_U25);
  nand ginst24449 (P3_SUB_485_U59, P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P3_SUB_485_U8);
  nand ginst24450 (P3_SUB_485_U6, P3_SUB_485_U42, P3_SUB_485_U43);
  nand ginst24451 (P3_SUB_485_U60, P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN, P3_SUB_485_U26);
  not ginst24452 (P3_SUB_485_U61, P3_SUB_485_U23);
  nand ginst24453 (P3_SUB_485_U62, P3_SUB_485_U28, P3_SUB_485_U61);
  nand ginst24454 (P3_SUB_485_U63, P3_SUB_485_U23, P3_SUB_485_U7);
  nand ginst24455 (P3_SUB_485_U7, P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN, P3_SUB_485_U27);
  not ginst24456 (P3_SUB_485_U8, P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN);
  not ginst24457 (P3_SUB_485_U9, P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN);
  not ginst24458 (P3_SUB_504_U10, P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN);
  not ginst24459 (P3_SUB_504_U11, P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN);
  not ginst24460 (P3_SUB_504_U12, P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN);
  not ginst24461 (P3_SUB_504_U13, P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN);
  nand ginst24462 (P3_SUB_504_U14, P3_SUB_504_U38, P3_SUB_504_U39);
  not ginst24463 (P3_SUB_504_U15, P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN);
  nand ginst24464 (P3_SUB_504_U16, P3_SUB_504_U47, P3_SUB_504_U48);
  nand ginst24465 (P3_SUB_504_U17, P3_SUB_504_U52, P3_SUB_504_U53);
  nand ginst24466 (P3_SUB_504_U18, P3_SUB_504_U57, P3_SUB_504_U58);
  nand ginst24467 (P3_SUB_504_U19, P3_SUB_504_U62, P3_SUB_504_U63);
  nand ginst24468 (P3_SUB_504_U20, P3_SUB_504_U44, P3_SUB_504_U45);
  nand ginst24469 (P3_SUB_504_U21, P3_SUB_504_U49, P3_SUB_504_U50);
  nand ginst24470 (P3_SUB_504_U22, P3_SUB_504_U54, P3_SUB_504_U55);
  nand ginst24471 (P3_SUB_504_U23, P3_SUB_504_U59, P3_SUB_504_U60);
  nand ginst24472 (P3_SUB_504_U24, P3_SUB_504_U34, P3_SUB_504_U35);
  nand ginst24473 (P3_SUB_504_U25, P3_SUB_504_U30, P3_SUB_504_U31);
  not ginst24474 (P3_SUB_504_U26, P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN);
  not ginst24475 (P3_SUB_504_U27, P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN);
  not ginst24476 (P3_SUB_504_U28, P3_SUB_504_U7);
  nand ginst24477 (P3_SUB_504_U29, P3_SUB_504_U28, P3_SUB_504_U8);
  nand ginst24478 (P3_SUB_504_U30, P3_SUB_504_U26, P3_SUB_504_U29);
  nand ginst24479 (P3_SUB_504_U31, P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN, P3_SUB_504_U7);
  not ginst24480 (P3_SUB_504_U32, P3_SUB_504_U25);
  nand ginst24481 (P3_SUB_504_U33, P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN, P3_SUB_504_U10);
  nand ginst24482 (P3_SUB_504_U34, P3_SUB_504_U25, P3_SUB_504_U33);
  nand ginst24483 (P3_SUB_504_U35, P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN, P3_SUB_504_U9);
  not ginst24484 (P3_SUB_504_U36, P3_SUB_504_U24);
  nand ginst24485 (P3_SUB_504_U37, P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P3_SUB_504_U12);
  nand ginst24486 (P3_SUB_504_U38, P3_SUB_504_U24, P3_SUB_504_U37);
  nand ginst24487 (P3_SUB_504_U39, P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN, P3_SUB_504_U11);
  not ginst24488 (P3_SUB_504_U40, P3_SUB_504_U14);
  nand ginst24489 (P3_SUB_504_U41, P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN, P3_SUB_504_U15);
  nand ginst24490 (P3_SUB_504_U42, P3_SUB_504_U40, P3_SUB_504_U41);
  nand ginst24491 (P3_SUB_504_U43, P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN, P3_SUB_504_U13);
  nand ginst24492 (P3_SUB_504_U44, P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN, P3_SUB_504_U13);
  nand ginst24493 (P3_SUB_504_U45, P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN, P3_SUB_504_U15);
  not ginst24494 (P3_SUB_504_U46, P3_SUB_504_U20);
  nand ginst24495 (P3_SUB_504_U47, P3_SUB_504_U40, P3_SUB_504_U46);
  nand ginst24496 (P3_SUB_504_U48, P3_SUB_504_U14, P3_SUB_504_U20);
  nand ginst24497 (P3_SUB_504_U49, P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P3_SUB_504_U12);
  nand ginst24498 (P3_SUB_504_U50, P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN, P3_SUB_504_U11);
  not ginst24499 (P3_SUB_504_U51, P3_SUB_504_U21);
  nand ginst24500 (P3_SUB_504_U52, P3_SUB_504_U36, P3_SUB_504_U51);
  nand ginst24501 (P3_SUB_504_U53, P3_SUB_504_U21, P3_SUB_504_U24);
  nand ginst24502 (P3_SUB_504_U54, P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN, P3_SUB_504_U10);
  nand ginst24503 (P3_SUB_504_U55, P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN, P3_SUB_504_U9);
  not ginst24504 (P3_SUB_504_U56, P3_SUB_504_U22);
  nand ginst24505 (P3_SUB_504_U57, P3_SUB_504_U32, P3_SUB_504_U56);
  nand ginst24506 (P3_SUB_504_U58, P3_SUB_504_U22, P3_SUB_504_U25);
  nand ginst24507 (P3_SUB_504_U59, P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P3_SUB_504_U8);
  nand ginst24508 (P3_SUB_504_U6, P3_SUB_504_U42, P3_SUB_504_U43);
  nand ginst24509 (P3_SUB_504_U60, P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN, P3_SUB_504_U26);
  not ginst24510 (P3_SUB_504_U61, P3_SUB_504_U23);
  nand ginst24511 (P3_SUB_504_U62, P3_SUB_504_U28, P3_SUB_504_U61);
  nand ginst24512 (P3_SUB_504_U63, P3_SUB_504_U23, P3_SUB_504_U7);
  nand ginst24513 (P3_SUB_504_U7, P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN, P3_SUB_504_U27);
  not ginst24514 (P3_SUB_504_U8, P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN);
  not ginst24515 (P3_SUB_504_U9, P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN);
  not ginst24516 (P3_SUB_563_U6, P3_U3305);
  not ginst24517 (P3_SUB_563_U7, P3_U3306);
  nand ginst24518 (P3_SUB_580_U10, P3_INSTADDRPOINTER_REG_0__SCAN_IN, P3_SUB_580_U7);
  nand ginst24519 (P3_SUB_580_U6, P3_SUB_580_U10, P3_SUB_580_U9);
  not ginst24520 (P3_SUB_580_U7, P3_INSTADDRPOINTER_REG_1__SCAN_IN);
  not ginst24521 (P3_SUB_580_U8, P3_INSTADDRPOINTER_REG_0__SCAN_IN);
  nand ginst24522 (P3_SUB_580_U9, P3_INSTADDRPOINTER_REG_1__SCAN_IN, P3_SUB_580_U8);
  not ginst24523 (P3_SUB_589_U6, P3_U3301);
  not ginst24524 (P3_SUB_589_U7, P3_U3302);
  not ginst24525 (P3_SUB_589_U8, P3_U2632);
  not ginst24526 (P3_SUB_589_U9, P3_U3300);
  nor ginst24527 (P3_U2352, P3_STATEBS16_REG_SCAN_IN, U209);
  and ginst24528 (P3_U2353, P3_U2449, P3_U3354);
  and ginst24529 (P3_U2354, P3_U3688, P3_U4325);
  and ginst24530 (P3_U2355, P3_U3689, P3_U4325);
  and ginst24531 (P3_U2356, P3_U2353, P3_U3355);
  and ginst24532 (P3_U2357, P3_U2451, P3_U4323);
  and ginst24533 (P3_U2358, P3_U3690, P3_U4341);
  and ginst24534 (P3_U2359, P3_U2462, P3_U4324);
  and ginst24535 (P3_U2360, P3_U2462, P3_U4296);
  and ginst24536 (P3_U2361, P3_U2462, P3_U4297);
  and ginst24537 (P3_U2362, P3_U3691, P3_U4341);
  and ginst24538 (P3_U2363, P3_U5435, P3_U5442);
  and ginst24539 (P3_U2364, P3_U3204, P3_U5392);
  and ginst24540 (P3_U2365, P3_U3201, P3_U5341);
  and ginst24541 (P3_U2366, P3_U3198, P3_U5290);
  and ginst24542 (P3_U2367, P3_U5232, P3_U5239);
  and ginst24543 (P3_U2368, P3_U3193, P3_U5189);
  and ginst24544 (P3_U2369, P3_U3189, P3_U5137);
  and ginst24545 (P3_U2370, P3_U3185, P3_U5085);
  and ginst24546 (P3_U2371, P3_U5028, P3_U5036);
  and ginst24547 (P3_U2372, P3_U3176, P3_U4985);
  and ginst24548 (P3_U2373, P3_U3172, P3_U4933);
  and ginst24549 (P3_U2374, P3_U3168, P3_U4881);
  and ginst24550 (P3_U2375, P3_U4821, P3_U4829);
  and ginst24551 (P3_U2376, P3_U3160, P3_U4778);
  and ginst24552 (P3_U2377, P3_U3152, P3_U4726);
  and ginst24553 (P3_U2378, P3_U3146, P3_U4674);
  and ginst24554 (P3_U2379, P3_U4312, P3_U4322);
  and ginst24555 (P3_U2380, P3_STATE2_REG_2__SCAN_IN, P3_U3260);
  and ginst24556 (P3_U2381, P3_STATE2_REG_3__SCAN_IN, P3_U4312);
  and ginst24557 (P3_U2382, P3_U3249, P3_U3951);
  and ginst24558 (P3_U2383, P3_U2380, P3_U4296);
  and ginst24559 (P3_U2384, P3_U2380, P3_U4297);
  and ginst24560 (P3_U2385, P3_STATE2_REG_1__SCAN_IN, P3_U3260);
  and ginst24561 (P3_U2386, P3_STATE2_REG_1__SCAN_IN, P3_U3249);
  and ginst24562 (P3_U2387, P3_U3249, P3_U3953);
  and ginst24563 (P3_U2388, P3_U3249, P3_U3952);
  and ginst24564 (P3_U2389, P3_U3249, P3_U4354);
  and ginst24565 (P3_U2390, P3_STATE2_REG_0__SCAN_IN, P3_U4353);
  and ginst24566 (P3_U2391, P3_U3218, P3_U4310);
  and ginst24567 (P3_U2392, P3_U2383, P3_U4293);
  and ginst24568 (P3_U2393, P3_U2361, P3_U2628);
  and ginst24569 (P3_U2394, P3_U2382, P3_U2628);
  and ginst24570 (P3_U2395, P3_U2361, P3_U3241);
  and ginst24571 (P3_U2396, P3_U2382, P3_U3241);
  and ginst24572 (P3_U2397, P3_STATEBS16_REG_SCAN_IN, P3_U2386);
  and ginst24573 (P3_U2398, P3_U2386, P3_U2631);
  and ginst24574 (P3_U2399, P3_U4309, P3_U4573);
  and ginst24575 (P3_U2400, P3_U4310, P3_U4573);
  and ginst24576 (P3_U2401, P3_STATE2_REG_3__SCAN_IN, P3_U3260);
  and ginst24577 (P3_U2402, P3_U3090, P3_U3248);
  and ginst24578 (P3_U2403, P3_U2385, P3_U3258);
  and ginst24579 (P3_U2404, P3_U2384, P3_U3257);
  and ginst24580 (P3_U2405, P3_U2384, P3_U7095);
  and ginst24581 (P3_U2406, P3_U3104, P3_U4311);
  and ginst24582 (P3_U2407, P3_U4311, P3_U4505);
  and ginst24583 (P3_U2408, P3_U3218, P3_U4309);
  and ginst24584 (P3_U2409, P3_STATE2_REG_0__SCAN_IN, P3_U3251);
  and ginst24585 (P3_U2410, P3_U3121, P3_U3251);
  and ginst24586 (P3_U2411, P3_U4310, P3_U4608);
  and ginst24587 (P3_U2412, P3_U3107, P3_U3218, P3_U4539);
  and ginst24588 (P3_U2413, BUF2_REG_0__SCAN_IN, P3_U4312);
  and ginst24589 (P3_U2414, BUF2_REG_1__SCAN_IN, P3_U4312);
  and ginst24590 (P3_U2415, BUF2_REG_2__SCAN_IN, P3_U4312);
  and ginst24591 (P3_U2416, BUF2_REG_3__SCAN_IN, P3_U4312);
  and ginst24592 (P3_U2417, BUF2_REG_4__SCAN_IN, P3_U4312);
  and ginst24593 (P3_U2418, BUF2_REG_5__SCAN_IN, P3_U4312);
  and ginst24594 (P3_U2419, BUF2_REG_6__SCAN_IN, P3_U4312);
  and ginst24595 (P3_U2420, BUF2_REG_7__SCAN_IN, P3_U4312);
  and ginst24596 (P3_U2421, BUF2_REG_24__SCAN_IN, P3_U2379);
  and ginst24597 (P3_U2422, BUF2_REG_16__SCAN_IN, P3_U2379);
  and ginst24598 (P3_U2423, BUF2_REG_25__SCAN_IN, P3_U2379);
  and ginst24599 (P3_U2424, BUF2_REG_17__SCAN_IN, P3_U2379);
  and ginst24600 (P3_U2425, BUF2_REG_26__SCAN_IN, P3_U2379);
  and ginst24601 (P3_U2426, BUF2_REG_18__SCAN_IN, P3_U2379);
  and ginst24602 (P3_U2427, BUF2_REG_27__SCAN_IN, P3_U2379);
  and ginst24603 (P3_U2428, BUF2_REG_19__SCAN_IN, P3_U2379);
  and ginst24604 (P3_U2429, BUF2_REG_28__SCAN_IN, P3_U2379);
  and ginst24605 (P3_U2430, BUF2_REG_20__SCAN_IN, P3_U2379);
  and ginst24606 (P3_U2431, BUF2_REG_29__SCAN_IN, P3_U2379);
  and ginst24607 (P3_U2432, BUF2_REG_21__SCAN_IN, P3_U2379);
  and ginst24608 (P3_U2433, BUF2_REG_30__SCAN_IN, P3_U2379);
  and ginst24609 (P3_U2434, BUF2_REG_22__SCAN_IN, P3_U2379);
  and ginst24610 (P3_U2435, BUF2_REG_31__SCAN_IN, P3_U2379);
  and ginst24611 (P3_U2436, BUF2_REG_23__SCAN_IN, P3_U2379);
  and ginst24612 (P3_U2437, P3_U2381, P3_U3108);
  and ginst24613 (P3_U2438, P3_U2381, P3_U3104);
  and ginst24614 (P3_U2439, P3_U2381, P3_U3101);
  and ginst24615 (P3_U2440, P3_U2381, P3_U3107);
  and ginst24616 (P3_U2441, P3_U2381, P3_U3102);
  and ginst24617 (P3_U2442, P3_U2381, P3_U3110);
  and ginst24618 (P3_U2443, P3_U2381, P3_U3074);
  and ginst24619 (P3_U2444, P3_U2391, P3_U3074);
  and ginst24620 (P3_U2445, P3_U2381, P3_U3218);
  and ginst24621 (P3_U2446, P3_U2391, P3_U3113);
  and ginst24622 (P3_U2447, P3_U2409, P3_U3108);
  and ginst24623 (P3_U2448, P3_U2391, P3_U4590);
  and ginst24624 (P3_U2449, P3_U4344, P3_U4522);
  and ginst24625 (P3_U2450, P3_U3660, P3_U4351);
  and ginst24626 (P3_U2451, P3_U2412, P3_U3102, P3_U4608);
  and ginst24627 (P3_U2452, P3_U2412, P3_U2463, P3_U4522);
  and ginst24628 (P3_U2453, P3_STATE2_REG_2__SCAN_IN, P3_STATE2_REG_1__SCAN_IN);
  and ginst24629 (P3_U2454, P3_U2380, P3_U4323);
  and ginst24630 (P3_U2455, P3_U2380, P3_U4324);
  and ginst24631 (P3_U2456, P3_U4556, P3_U4607);
  and ginst24632 (P3_U2457, P3_U3139, P3_U3269);
  and ginst24633 (P3_U2458, P3_U3269, P3_U4652);
  and ginst24634 (P3_U2459, P3_U3139, P3_U7962);
  and ginst24635 (P3_U2460, P3_U4652, P3_U7962);
  and ginst24636 (P3_U2461, P3_U4522, P3_U4573);
  and ginst24637 (P3_U2462, P3_U2412, P3_U2449);
  and ginst24638 (P3_U2463, P3_U4590, P3_U4607);
  and ginst24639 (P3_U2464, P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN);
  and ginst24640 (P3_U2465, P3_U2464, P3_U4332);
  and ginst24641 (P3_U2466, P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P3_U3093);
  and ginst24642 (P3_U2467, P3_U2464, P3_U2466);
  and ginst24643 (P3_U2468, P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN, P3_U3094);
  and ginst24644 (P3_U2469, P3_U2464, P3_U2468);
  and ginst24645 (P3_U2470, P3_U2464, P3_U4467);
  and ginst24646 (P3_U2471, P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P3_U4468);
  and ginst24647 (P3_U2472, P3_U2466, P3_U3097);
  and ginst24648 (P3_U2473, P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P3_U2472);
  and ginst24649 (P3_U2474, P3_U2468, P3_U3097);
  and ginst24650 (P3_U2475, P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P3_U2474);
  and ginst24651 (P3_U2476, P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P3_U4469);
  and ginst24652 (P3_U2477, P3_U2466, P3_U4470);
  and ginst24653 (P3_U2478, P3_U2468, P3_U4470);
  and ginst24654 (P3_U2479, P3_U4467, P3_U4470);
  and ginst24655 (P3_U2480, P3_U3100, P3_U4468);
  nor ginst24656 (P3_U2481, P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN);
  and ginst24657 (P3_U2482, P3_U2466, P3_U2481);
  and ginst24658 (P3_U2483, P3_U2468, P3_U2481);
  and ginst24659 (P3_U2484, P3_U3100, P3_U4469);
  and ginst24660 (P3_U2485, P3_U3270, P3_U4656);
  and ginst24661 (P3_U2486, P3_U3182, P3_U3271);
  and ginst24662 (P3_U2487, P3_U3142, P3_U3270);
  and ginst24663 (P3_U2488, P3_U2487, P3_U4657);
  and ginst24664 (P3_U2489, P3_U3090, P3_U4315);
  and ginst24665 (P3_U2490, P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P3_U3156);
  and ginst24666 (P3_U2491, P3_U2487, P3_U4644);
  and ginst24667 (P3_U2492, P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN, P3_U3128);
  and ginst24668 (P3_U2493, P3_U3128, P3_U4646);
  and ginst24669 (P3_U2494, P3_U2487, P3_U4645);
  and ginst24670 (P3_U2495, P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P3_U4646);
  and ginst24671 (P3_U2496, P3_U3128, P3_U4643);
  and ginst24672 (P3_U2497, P3_U2487, P3_U2496);
  and ginst24673 (P3_U2498, P3_U3182, P3_U7968);
  and ginst24674 (P3_U2499, P3_U4657, P3_U4658);
  and ginst24675 (P3_U2500, P3_U4644, P3_U4658);
  nor ginst24676 (P3_U2501, P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN, P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN);
  and ginst24677 (P3_U2502, P3_U4645, P3_U4658);
  and ginst24678 (P3_U2503, P3_U2496, P3_U4658);
  and ginst24679 (P3_U2504, P3_U3271, P3_U4660);
  and ginst24680 (P3_U2505, P3_U2485, P3_U4644);
  and ginst24681 (P3_U2506, P3_U2485, P3_U4645);
  and ginst24682 (P3_U2507, P3_U2485, P3_U2496);
  and ginst24683 (P3_U2508, P3_U4660, P3_U7968);
  and ginst24684 (P3_U2509, P3_U4656, P3_U7965);
  and ginst24685 (P3_U2510, P3_U2509, P3_U4657);
  and ginst24686 (P3_U2511, P3_U2509, P3_U4644);
  and ginst24687 (P3_U2512, P3_U2509, P3_U4645);
  and ginst24688 (P3_U2513, P3_U2496, P3_U2509);
  and ginst24689 (P3_U2514, P3_U3216, P3_U3218);
  and ginst24690 (P3_U2515, P3_U5485, P3_U7969, P3_U7970);
  and ginst24691 (P3_U2516, P3_U5492, P3_U5493);
  and ginst24692 (P3_U2517, P3_U3246, P3_U5526);
  and ginst24693 (P3_U2518, P3_U3668, P3_U5522);
  and ginst24694 (P3_U2519, P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN, P3_U3228);
  and ginst24695 (P3_U2520, P3_U5543, P3_U5548);
  and ginst24696 (P3_U2521, P3_U2519, P3_U2520);
  and ginst24697 (P3_U2522, P3_U3093, P3_U3228);
  and ginst24698 (P3_U2523, P3_U2520, P3_U2522);
  and ginst24699 (P3_U2524, P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN, P3_U5558);
  and ginst24700 (P3_U2525, P3_U2520, P3_U2524);
  and ginst24701 (P3_U2526, P3_U3093, P3_U5558);
  and ginst24702 (P3_U2527, P3_U2520, P3_U2526);
  and ginst24703 (P3_U2528, P3_U3225, P3_U5543);
  and ginst24704 (P3_U2529, P3_U2519, P3_U2528);
  and ginst24705 (P3_U2530, P3_U2522, P3_U2528);
  and ginst24706 (P3_U2531, P3_U2524, P3_U2528);
  and ginst24707 (P3_U2532, P3_U2526, P3_U2528);
  and ginst24708 (P3_U2533, P3_U3265, P3_U5548);
  and ginst24709 (P3_U2534, P3_U2519, P3_U2533);
  and ginst24710 (P3_U2535, P3_U2522, P3_U2533);
  and ginst24711 (P3_U2536, P3_U2524, P3_U2533);
  and ginst24712 (P3_U2537, P3_U2526, P3_U2533);
  and ginst24713 (P3_U2538, P3_U3225, P3_U3265);
  and ginst24714 (P3_U2539, P3_U2519, P3_U2538);
  and ginst24715 (P3_U2540, P3_U2522, P3_U2538);
  and ginst24716 (P3_U2541, P3_U2524, P3_U2538);
  and ginst24717 (P3_U2542, P3_U2526, P3_U2538);
  and ginst24718 (P3_U2543, P3_U3266, P3_U3272);
  and ginst24719 (P3_U2544, P3_U2468, P3_U2543);
  and ginst24720 (P3_U2545, P3_U2543, P3_U4467);
  and ginst24721 (P3_U2546, P3_U2543, P3_U4332);
  and ginst24722 (P3_U2547, P3_U2466, P3_U2543);
  and ginst24723 (P3_U2548, P3_U3266, P3_U8034);
  and ginst24724 (P3_U2549, P3_U2468, P3_U2548);
  and ginst24725 (P3_U2550, P3_U2548, P3_U4467);
  and ginst24726 (P3_U2551, P3_U2548, P3_U4332);
  and ginst24727 (P3_U2552, P3_U2466, P3_U2548);
  and ginst24728 (P3_U2553, P3_U3272, P3_U7516);
  and ginst24729 (P3_U2554, P3_U2468, P3_U2553);
  and ginst24730 (P3_U2555, P3_U2553, P3_U4467);
  and ginst24731 (P3_U2556, P3_U2553, P3_U4332);
  and ginst24732 (P3_U2557, P3_U2466, P3_U2553);
  and ginst24733 (P3_U2558, P3_U7516, P3_U8034);
  and ginst24734 (P3_U2559, P3_U2468, P3_U2558);
  and ginst24735 (P3_U2560, P3_U2558, P3_U4467);
  and ginst24736 (P3_U2561, P3_U2558, P3_U4332);
  and ginst24737 (P3_U2562, P3_U2466, P3_U2558);
  and ginst24738 (P3_U2563, P3_U4291, P3_U8037);
  and ginst24739 (P3_U2564, P3_U2522, P3_U2563);
  and ginst24740 (P3_U2565, P3_U2519, P3_U2563);
  and ginst24741 (P3_U2566, P3_U2526, P3_U2563);
  and ginst24742 (P3_U2567, P3_U2524, P3_U2563);
  and ginst24743 (P3_U2568, P3_U3267, P3_U8037);
  and ginst24744 (P3_U2569, P3_U2522, P3_U2568);
  and ginst24745 (P3_U2570, P3_U2519, P3_U2568);
  and ginst24746 (P3_U2571, P3_U2526, P3_U2568);
  and ginst24747 (P3_U2572, P3_U2524, P3_U2568);
  and ginst24748 (P3_U2573, P3_U3273, P3_U4291);
  and ginst24749 (P3_U2574, P3_U2522, P3_U2573);
  and ginst24750 (P3_U2575, P3_U2519, P3_U2573);
  and ginst24751 (P3_U2576, P3_U2526, P3_U2573);
  and ginst24752 (P3_U2577, P3_U2524, P3_U2573);
  and ginst24753 (P3_U2578, P3_U3267, P3_U3273);
  and ginst24754 (P3_U2579, P3_U2522, P3_U2578);
  and ginst24755 (P3_U2580, P3_U2519, P3_U2578);
  and ginst24756 (P3_U2581, P3_U2526, P3_U2578);
  and ginst24757 (P3_U2582, P3_U2524, P3_U2578);
  and ginst24758 (P3_U2583, P3_U4468, P3_U7775);
  and ginst24759 (P3_U2584, P3_U2472, P3_U7775);
  and ginst24760 (P3_U2585, P3_U2474, P3_U7775);
  and ginst24761 (P3_U2586, P3_U4469, P3_U7775);
  and ginst24762 (P3_U2587, P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN, P3_U7775);
  and ginst24763 (P3_U2588, P3_U2587, P3_U4332);
  and ginst24764 (P3_U2589, P3_U2466, P3_U2587);
  and ginst24765 (P3_U2590, P3_U2468, P3_U2587);
  and ginst24766 (P3_U2591, P3_U2587, P3_U4467);
  and ginst24767 (P3_U2592, P3_U3268, P3_U4468);
  and ginst24768 (P3_U2593, P3_U2472, P3_U3268);
  and ginst24769 (P3_U2594, P3_U2474, P3_U3268);
  and ginst24770 (P3_U2595, P3_U3268, P3_U4469);
  and ginst24771 (P3_U2596, P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN, P3_U3268);
  and ginst24772 (P3_U2597, P3_U2596, P3_U4332);
  and ginst24773 (P3_U2598, P3_U2466, P3_U2596);
  and ginst24774 (P3_U2599, P3_U2468, P3_U2596);
  and ginst24775 (P3_U2600, P3_U2596, P3_U4467);
  and ginst24776 (P3_U2601, P3_U2352, P3_U2392);
  and ginst24777 (P3_U2602, P3_EBX_REG_31__SCAN_IN, P3_U2404);
  and ginst24778 (P3_U2603, P3_U4133, P3_U7358, P3_U7359, P3_U7360);
  and ginst24779 (P3_U2604, P3_U7946, P3_U7947);
  nand ginst24780 (P3_U2605, P3_U4212, P3_U4213, P3_U4214, P3_U4215);
  nand ginst24781 (P3_U2606, P3_U4208, P3_U4209, P3_U4210, P3_U4211);
  nand ginst24782 (P3_U2607, P3_U4204, P3_U4205, P3_U4206, P3_U4207);
  nand ginst24783 (P3_U2608, P3_U4200, P3_U4201, P3_U4202, P3_U4203);
  nand ginst24784 (P3_U2609, P3_U4196, P3_U4197, P3_U4198, P3_U4199);
  nand ginst24785 (P3_U2610, P3_U4192, P3_U4193, P3_U4194, P3_U4195);
  nand ginst24786 (P3_U2611, P3_U4188, P3_U4189, P3_U4190, P3_U4191);
  nand ginst24787 (P3_U2612, P3_U4184, P3_U4185, P3_U4186, P3_U4187);
  nand ginst24788 (P3_U2613, P3_U4276, P3_U4277, P3_U4278, P3_U4279);
  nand ginst24789 (P3_U2614, P3_U4272, P3_U4273, P3_U4274, P3_U4275);
  nand ginst24790 (P3_U2615, P3_U4268, P3_U4269, P3_U4270, P3_U4271);
  nand ginst24791 (P3_U2616, P3_U4264, P3_U4265, P3_U4266, P3_U4267);
  nand ginst24792 (P3_U2617, P3_U4260, P3_U4261, P3_U4262, P3_U4263);
  nand ginst24793 (P3_U2618, P3_U4256, P3_U4257, P3_U4258, P3_U4259);
  nand ginst24794 (P3_U2619, P3_U4252, P3_U4253, P3_U4254, P3_U4255);
  nand ginst24795 (P3_U2620, P3_U4248, P3_U4249, P3_U4250, P3_U4251);
  nand ginst24796 (P3_U2621, P3_U4180, P3_U4181, P3_U4182, P3_U4183);
  nand ginst24797 (P3_U2622, P3_U4176, P3_U4177, P3_U4178, P3_U4179);
  nand ginst24798 (P3_U2623, P3_U4172, P3_U4173, P3_U4174, P3_U4175);
  nand ginst24799 (P3_U2624, P3_U4168, P3_U4169, P3_U4170, P3_U4171);
  nand ginst24800 (P3_U2625, P3_U4164, P3_U4165, P3_U4166, P3_U4167);
  nand ginst24801 (P3_U2626, P3_U4160, P3_U4161, P3_U4162, P3_U4163);
  nand ginst24802 (P3_U2627, P3_U4156, P3_U4157, P3_U4158, P3_U4159);
  nand ginst24803 (P3_U2628, P3_U4152, P3_U4153, P3_U4154, P3_U4155);
  and ginst24804 (P3_U2629, P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN, P3_U3207);
  not ginst24805 (P3_U2630, U209);
  not ginst24806 (P3_U2631, P3_STATEBS16_REG_SCAN_IN);
  and ginst24807 (P3_U2632, P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P3_U3207);
  nand ginst24808 (P3_U2633, P3_U7383, P3_U7937);
  nand ginst24809 (P3_U2634, P3_U7381, P3_U7382);
  nand ginst24810 (P3_U2635, P3_U4335, P3_U8024, P3_U8025);
  nand ginst24811 (P3_U2636, P3_U4335, P3_U8020, P3_U8021);
  nand ginst24812 (P3_U2637, P3_U7369, P3_U7370);
  nand ginst24813 (P3_U2638, P3_U4327, P3_U8012, P3_U8013);
  nand ginst24814 (P3_U2639, P3_U4327, P3_U8002, P3_U8003);
  and ginst24815 (P3_U2640, P3_U7357, P3_U7907);
  nand ginst24816 (P3_U2641, P3_U4129, P3_U4130, P3_U7351, P3_U7352, P3_U7354);
  nand ginst24817 (P3_U2642, P3_U4126, P3_U4127, P3_U7343, P3_U7344, P3_U7346);
  nand ginst24818 (P3_U2643, P3_U4123, P3_U4124, P3_U7335, P3_U7336, P3_U7338);
  nand ginst24819 (P3_U2644, P3_U4120, P3_U4121, P3_U7327, P3_U7328, P3_U7330);
  nand ginst24820 (P3_U2645, P3_U4117, P3_U4118, P3_U7319, P3_U7320, P3_U7322);
  nand ginst24821 (P3_U2646, P3_U4114, P3_U4115, P3_U7311, P3_U7312, P3_U7314);
  nand ginst24822 (P3_U2647, P3_U4111, P3_U4112, P3_U7303, P3_U7304, P3_U7306);
  nand ginst24823 (P3_U2648, P3_U4108, P3_U4109, P3_U7295, P3_U7296, P3_U7298);
  nand ginst24824 (P3_U2649, P3_U4105, P3_U4106, P3_U7287, P3_U7288, P3_U7290);
  nand ginst24825 (P3_U2650, P3_U4102, P3_U4103, P3_U7279, P3_U7280, P3_U7282);
  nand ginst24826 (P3_U2651, P3_U4099, P3_U4100, P3_U7271, P3_U7272, P3_U7274);
  nand ginst24827 (P3_U2652, P3_U4096, P3_U4097, P3_U7263, P3_U7264, P3_U7266);
  nand ginst24828 (P3_U2653, P3_U4093, P3_U4094, P3_U7255, P3_U7256, P3_U7258);
  nand ginst24829 (P3_U2654, P3_U4090, P3_U4091, P3_U7247, P3_U7248, P3_U7250);
  nand ginst24830 (P3_U2655, P3_U4087, P3_U4088, P3_U7239, P3_U7240, P3_U7242);
  nand ginst24831 (P3_U2656, P3_U4084, P3_U4085, P3_U7231, P3_U7232, P3_U7234);
  nand ginst24832 (P3_U2657, P3_U4081, P3_U4082, P3_U7223, P3_U7224, P3_U7226);
  nand ginst24833 (P3_U2658, P3_U4078, P3_U4079, P3_U7215, P3_U7216, P3_U7218);
  nand ginst24834 (P3_U2659, P3_U4075, P3_U4076, P3_U7207, P3_U7208, P3_U7210);
  nand ginst24835 (P3_U2660, P3_U4072, P3_U4073, P3_U7199, P3_U7200, P3_U7202);
  nand ginst24836 (P3_U2661, P3_U4069, P3_U4070, P3_U7191, P3_U7192, P3_U7194);
  nand ginst24837 (P3_U2662, P3_U4066, P3_U4067, P3_U7183, P3_U7184, P3_U7186);
  nand ginst24838 (P3_U2663, P3_U4063, P3_U4064, P3_U7175, P3_U7176, P3_U7178);
  nand ginst24839 (P3_U2664, P3_U4060, P3_U4061, P3_U7167, P3_U7168, P3_U7170);
  nand ginst24840 (P3_U2665, P3_U4057, P3_U4058, P3_U7159, P3_U7160, P3_U7162);
  nand ginst24841 (P3_U2666, P3_U4054, P3_U4056);
  nand ginst24842 (P3_U2667, P3_U4049, P3_U4051);
  nand ginst24843 (P3_U2668, P3_U4043, P3_U4045, P3_U7129, P3_U7132, P3_U7133);
  nand ginst24844 (P3_U2669, P3_U4039, P3_U4041, P3_U7119, P3_U7122, P3_U7123);
  nand ginst24845 (P3_U2670, P3_U4035, P3_U4037, P3_U7109, P3_U7112, P3_U7113);
  nand ginst24846 (P3_U2671, P3_U4031, P3_U4033, P3_U7099, P3_U7102, P3_U7103);
  nand ginst24847 (P3_U2672, P3_U7091, P3_U7092);
  nand ginst24848 (P3_U2673, P3_U7088, P3_U7089, P3_U7090);
  nand ginst24849 (P3_U2674, P3_U7085, P3_U7086, P3_U7087);
  nand ginst24850 (P3_U2675, P3_U7082, P3_U7083, P3_U7084);
  nand ginst24851 (P3_U2676, P3_U7079, P3_U7080, P3_U7081);
  nand ginst24852 (P3_U2677, P3_U7076, P3_U7077, P3_U7078);
  nand ginst24853 (P3_U2678, P3_U7073, P3_U7074, P3_U7075);
  nand ginst24854 (P3_U2679, P3_U7070, P3_U7071, P3_U7072);
  nand ginst24855 (P3_U2680, P3_U7067, P3_U7068, P3_U7069);
  nand ginst24856 (P3_U2681, P3_U7064, P3_U7065, P3_U7066);
  nand ginst24857 (P3_U2682, P3_U7061, P3_U7062, P3_U7063);
  nand ginst24858 (P3_U2683, P3_U7058, P3_U7059, P3_U7060);
  nand ginst24859 (P3_U2684, P3_U7055, P3_U7056, P3_U7057);
  nand ginst24860 (P3_U2685, P3_U7052, P3_U7053, P3_U7054);
  nand ginst24861 (P3_U2686, P3_U7049, P3_U7050, P3_U7051);
  nand ginst24862 (P3_U2687, P3_U7046, P3_U7047, P3_U7048);
  nand ginst24863 (P3_U2688, P3_U7043, P3_U7044, P3_U7045);
  nand ginst24864 (P3_U2689, P3_U7040, P3_U7041, P3_U7042);
  nand ginst24865 (P3_U2690, P3_U7037, P3_U7038, P3_U7039);
  nand ginst24866 (P3_U2691, P3_U7034, P3_U7035, P3_U7036);
  nand ginst24867 (P3_U2692, P3_U7031, P3_U7032, P3_U7033);
  nand ginst24868 (P3_U2693, P3_U7028, P3_U7029, P3_U7030);
  nand ginst24869 (P3_U2694, P3_U7025, P3_U7026, P3_U7027);
  nand ginst24870 (P3_U2695, P3_U7022, P3_U7023, P3_U7024);
  nand ginst24871 (P3_U2696, P3_U7019, P3_U7020, P3_U7021);
  nand ginst24872 (P3_U2697, P3_U7016, P3_U7017, P3_U7018);
  nand ginst24873 (P3_U2698, P3_U7013, P3_U7014, P3_U7015);
  nand ginst24874 (P3_U2699, P3_U7010, P3_U7011, P3_U7012);
  nand ginst24875 (P3_U2700, P3_U7007, P3_U7008, P3_U7009);
  nand ginst24876 (P3_U2701, P3_U7004, P3_U7005, P3_U7006);
  nand ginst24877 (P3_U2702, P3_U7001, P3_U7002, P3_U7003);
  nand ginst24878 (P3_U2703, P3_U6998, P3_U6999, P3_U7000);
  nand ginst24879 (P3_U2704, P3_U6993, P3_U6994, P3_U6995);
  nand ginst24880 (P3_U2705, P3_U6988, P3_U6989, P3_U6990, P3_U6991, P3_U6992);
  nand ginst24881 (P3_U2706, P3_U6983, P3_U6984, P3_U6985, P3_U6986, P3_U6987);
  nand ginst24882 (P3_U2707, P3_U6978, P3_U6979, P3_U6980, P3_U6981, P3_U6982);
  nand ginst24883 (P3_U2708, P3_U4029, P3_U6973, P3_U6974, P3_U6976);
  nand ginst24884 (P3_U2709, P3_U4028, P3_U6968, P3_U6969, P3_U6971);
  nand ginst24885 (P3_U2710, P3_U4027, P3_U6963, P3_U6964, P3_U6966);
  nand ginst24886 (P3_U2711, P3_U4026, P3_U6958, P3_U6959, P3_U6961);
  nand ginst24887 (P3_U2712, P3_U4025, P3_U6953, P3_U6954, P3_U6956);
  nand ginst24888 (P3_U2713, P3_U4024, P3_U6948, P3_U6949, P3_U6951);
  nand ginst24889 (P3_U2714, P3_U4023, P3_U6943, P3_U6944, P3_U6946);
  nand ginst24890 (P3_U2715, P3_U4022, P3_U6938, P3_U6939, P3_U6941);
  nand ginst24891 (P3_U2716, P3_U4021, P3_U6933, P3_U6934, P3_U6936);
  nand ginst24892 (P3_U2717, P3_U4020, P3_U6928, P3_U6929, P3_U6931);
  nand ginst24893 (P3_U2718, P3_U4019, P3_U6923, P3_U6924, P3_U6926);
  nand ginst24894 (P3_U2719, P3_U4018, P3_U6918, P3_U6919, P3_U6921);
  nand ginst24895 (P3_U2720, P3_U4017, P3_U6914, P3_U6916);
  nand ginst24896 (P3_U2721, P3_U4016, P3_U6910, P3_U6912);
  nand ginst24897 (P3_U2722, P3_U4015, P3_U6906, P3_U6908);
  nand ginst24898 (P3_U2723, P3_U4014, P3_U6902, P3_U6903);
  nand ginst24899 (P3_U2724, P3_U4013, P3_U6898, P3_U6899);
  nand ginst24900 (P3_U2725, P3_U4012, P3_U6894, P3_U6895);
  nand ginst24901 (P3_U2726, P3_U4011, P3_U6890, P3_U6891);
  nand ginst24902 (P3_U2727, P3_U4010, P3_U6886, P3_U6887);
  nand ginst24903 (P3_U2728, P3_U4009, P3_U6882, P3_U6883);
  nand ginst24904 (P3_U2729, P3_U4008, P3_U6878, P3_U6879);
  nand ginst24905 (P3_U2730, P3_U4007, P3_U6874, P3_U6875);
  nand ginst24906 (P3_U2731, P3_U4006, P3_U6870, P3_U6871);
  nand ginst24907 (P3_U2732, P3_U4005, P3_U6866, P3_U6867);
  nand ginst24908 (P3_U2733, P3_U4004, P3_U6862, P3_U6863);
  nand ginst24909 (P3_U2734, P3_U4003, P3_U6858, P3_U6859);
  nand ginst24910 (P3_U2735, P3_U4002, P3_U6854, P3_U6855);
  and ginst24911 (P3_U2736, P3_DATAO_REG_31__SCAN_IN, P3_U6759);
  nand ginst24912 (P3_U2737, P3_U4001, P3_U6850);
  nand ginst24913 (P3_U2738, P3_U4000, P3_U6847);
  nand ginst24914 (P3_U2739, P3_U3999, P3_U6844);
  nand ginst24915 (P3_U2740, P3_U3998, P3_U6841);
  nand ginst24916 (P3_U2741, P3_U3997, P3_U6838);
  nand ginst24917 (P3_U2742, P3_U3996, P3_U6835);
  nand ginst24918 (P3_U2743, P3_U3995, P3_U6832);
  nand ginst24919 (P3_U2744, P3_U3994, P3_U6829);
  nand ginst24920 (P3_U2745, P3_U3993, P3_U6826);
  nand ginst24921 (P3_U2746, P3_U3992, P3_U6823);
  nand ginst24922 (P3_U2747, P3_U3991, P3_U6820);
  nand ginst24923 (P3_U2748, P3_U3990, P3_U6817);
  nand ginst24924 (P3_U2749, P3_U3989, P3_U6814);
  nand ginst24925 (P3_U2750, P3_U3988, P3_U6811);
  nand ginst24926 (P3_U2751, P3_U3987, P3_U6808);
  nand ginst24927 (P3_U2752, P3_U6805, P3_U6806, P3_U6807);
  nand ginst24928 (P3_U2753, P3_U6802, P3_U6803, P3_U6804);
  nand ginst24929 (P3_U2754, P3_U6799, P3_U6800, P3_U6801);
  nand ginst24930 (P3_U2755, P3_U6796, P3_U6797, P3_U6798);
  nand ginst24931 (P3_U2756, P3_U6793, P3_U6794, P3_U6795);
  nand ginst24932 (P3_U2757, P3_U6790, P3_U6791, P3_U6792);
  nand ginst24933 (P3_U2758, P3_U6787, P3_U6788, P3_U6789);
  nand ginst24934 (P3_U2759, P3_U6784, P3_U6785, P3_U6786);
  nand ginst24935 (P3_U2760, P3_U6781, P3_U6782, P3_U6783);
  nand ginst24936 (P3_U2761, P3_U6778, P3_U6779, P3_U6780);
  nand ginst24937 (P3_U2762, P3_U6775, P3_U6776, P3_U6777);
  nand ginst24938 (P3_U2763, P3_U6772, P3_U6773, P3_U6774);
  nand ginst24939 (P3_U2764, P3_U6769, P3_U6770, P3_U6771);
  nand ginst24940 (P3_U2765, P3_U6766, P3_U6767, P3_U6768);
  nand ginst24941 (P3_U2766, P3_U6763, P3_U6764, P3_U6765);
  nand ginst24942 (P3_U2767, P3_U6760, P3_U6761, P3_U6762);
  nand ginst24943 (P3_U2768, P3_U6754, P3_U6755, P3_U6756);
  nand ginst24944 (P3_U2769, P3_U6751, P3_U6752, P3_U6753);
  nand ginst24945 (P3_U2770, P3_U6748, P3_U6749, P3_U6750);
  nand ginst24946 (P3_U2771, P3_U6745, P3_U6746, P3_U6747);
  nand ginst24947 (P3_U2772, P3_U6742, P3_U6743, P3_U6744);
  nand ginst24948 (P3_U2773, P3_U6739, P3_U6740, P3_U6741);
  nand ginst24949 (P3_U2774, P3_U6736, P3_U6737, P3_U6738);
  nand ginst24950 (P3_U2775, P3_U6733, P3_U6734, P3_U6735);
  nand ginst24951 (P3_U2776, P3_U6730, P3_U6731, P3_U6732);
  nand ginst24952 (P3_U2777, P3_U6727, P3_U6728, P3_U6729);
  nand ginst24953 (P3_U2778, P3_U6724, P3_U6725, P3_U6726);
  nand ginst24954 (P3_U2779, P3_U6721, P3_U6722, P3_U6723);
  nand ginst24955 (P3_U2780, P3_U6718, P3_U6719, P3_U6720);
  nand ginst24956 (P3_U2781, P3_U6715, P3_U6716, P3_U6717);
  nand ginst24957 (P3_U2782, P3_U6712, P3_U6713, P3_U6714);
  nand ginst24958 (P3_U2783, P3_U6709, P3_U6710, P3_U6711);
  nand ginst24959 (P3_U2784, P3_U6706, P3_U6707, P3_U6708);
  nand ginst24960 (P3_U2785, P3_U6703, P3_U6704, P3_U6705);
  nand ginst24961 (P3_U2786, P3_U6700, P3_U6701, P3_U6702);
  nand ginst24962 (P3_U2787, P3_U6697, P3_U6698, P3_U6699);
  nand ginst24963 (P3_U2788, P3_U6694, P3_U6695, P3_U6696);
  nand ginst24964 (P3_U2789, P3_U6691, P3_U6692, P3_U6693);
  nand ginst24965 (P3_U2790, P3_U6688, P3_U6689, P3_U6690);
  nand ginst24966 (P3_U2791, P3_U6685, P3_U6686, P3_U6687);
  nand ginst24967 (P3_U2792, P3_U6682, P3_U6683, P3_U6684);
  nand ginst24968 (P3_U2793, P3_U6679, P3_U6680, P3_U6681);
  nand ginst24969 (P3_U2794, P3_U6676, P3_U6677, P3_U6678);
  nand ginst24970 (P3_U2795, P3_U6673, P3_U6674, P3_U6675);
  nand ginst24971 (P3_U2796, P3_U6670, P3_U6671, P3_U6672);
  nand ginst24972 (P3_U2797, P3_U6667, P3_U6668, P3_U6669);
  nand ginst24973 (P3_U2798, P3_U6664, P3_U6665, P3_U6666);
  nand ginst24974 (P3_U2799, P3_U3985, P3_U6653, P3_U6654, P3_U6655, P3_U6656);
  nand ginst24975 (P3_U2800, P3_U3984, P3_U6645, P3_U6646, P3_U6647, P3_U6648);
  nand ginst24976 (P3_U2801, P3_U3983, P3_U6637, P3_U6638, P3_U6639, P3_U6640);
  nand ginst24977 (P3_U2802, P3_U3982, P3_U6629, P3_U6630, P3_U6631, P3_U6632);
  nand ginst24978 (P3_U2803, P3_U3981, P3_U6621, P3_U6622, P3_U6623, P3_U6624);
  nand ginst24979 (P3_U2804, P3_U3980, P3_U6613, P3_U6614, P3_U6615, P3_U6616);
  nand ginst24980 (P3_U2805, P3_U3979, P3_U6605, P3_U6606, P3_U6607, P3_U6608);
  nand ginst24981 (P3_U2806, P3_U3978, P3_U6597, P3_U6598, P3_U6599, P3_U6600);
  nand ginst24982 (P3_U2807, P3_U3977, P3_U6589, P3_U6590, P3_U6591, P3_U6592);
  nand ginst24983 (P3_U2808, P3_U3976, P3_U6581, P3_U6582, P3_U6583, P3_U6584);
  nand ginst24984 (P3_U2809, P3_U3975, P3_U6573, P3_U6574, P3_U6575, P3_U6576);
  nand ginst24985 (P3_U2810, P3_U3974, P3_U6565, P3_U6566, P3_U6567, P3_U6568);
  nand ginst24986 (P3_U2811, P3_U3973, P3_U6557, P3_U6558, P3_U6559, P3_U6560);
  nand ginst24987 (P3_U2812, P3_U3972, P3_U6549, P3_U6550, P3_U6551, P3_U6552);
  nand ginst24988 (P3_U2813, P3_U3971, P3_U6541, P3_U6542, P3_U6543, P3_U6544);
  nand ginst24989 (P3_U2814, P3_U3970, P3_U6533, P3_U6534, P3_U6535, P3_U6536);
  nand ginst24990 (P3_U2815, P3_U3969, P3_U6525, P3_U6526, P3_U6527, P3_U6528);
  nand ginst24991 (P3_U2816, P3_U3968, P3_U6517, P3_U6518, P3_U6519, P3_U6520);
  nand ginst24992 (P3_U2817, P3_U3967, P3_U6509, P3_U6510, P3_U6511, P3_U6512);
  nand ginst24993 (P3_U2818, P3_U3966, P3_U6501, P3_U6502, P3_U6503, P3_U6504);
  nand ginst24994 (P3_U2819, P3_U3965, P3_U6493, P3_U6494, P3_U6495, P3_U6496);
  nand ginst24995 (P3_U2820, P3_U3964, P3_U6485, P3_U6486, P3_U6487, P3_U6488);
  nand ginst24996 (P3_U2821, P3_U3963, P3_U6477, P3_U6478, P3_U6479, P3_U6480);
  nand ginst24997 (P3_U2822, P3_U3962, P3_U6469, P3_U6470, P3_U6471, P3_U6472);
  nand ginst24998 (P3_U2823, P3_U3961, P3_U6461, P3_U6462, P3_U6463, P3_U6464);
  nand ginst24999 (P3_U2824, P3_U3960, P3_U6453, P3_U6454, P3_U6455, P3_U6456);
  nand ginst25000 (P3_U2825, P3_U3959, P3_U6445, P3_U6446, P3_U6447, P3_U6448);
  nand ginst25001 (P3_U2826, P3_U3958, P3_U6437, P3_U6438, P3_U6439, P3_U6440);
  nand ginst25002 (P3_U2827, P3_U3957, P3_U6429, P3_U6430, P3_U6431, P3_U6432);
  nand ginst25003 (P3_U2828, P3_U3956, P3_U6421, P3_U6422, P3_U6423, P3_U6424);
  nand ginst25004 (P3_U2829, P3_U3955, P3_U6413, P3_U6414, P3_U6415, P3_U6416);
  nand ginst25005 (P3_U2830, P3_U3954, P3_U6405, P3_U6406, P3_U6407, P3_U6408);
  and ginst25006 (P3_U2831, P3_U6396, P3_U7906);
  nand ginst25007 (P3_U2832, P3_U6373, P3_U6374, P3_U6375);
  nand ginst25008 (P3_U2833, P3_U6349, P3_U6350, P3_U6351);
  nand ginst25009 (P3_U2834, P3_U6325, P3_U6326, P3_U6327);
  nand ginst25010 (P3_U2835, P3_U6301, P3_U6302, P3_U6303);
  nand ginst25011 (P3_U2836, P3_U6277, P3_U6278, P3_U6279);
  nand ginst25012 (P3_U2837, P3_U3893, P3_U6254);
  nand ginst25013 (P3_U2838, P3_U3883, P3_U6230);
  nand ginst25014 (P3_U2839, P3_U3873, P3_U6206);
  nand ginst25015 (P3_U2840, P3_U3863, P3_U6182);
  nand ginst25016 (P3_U2841, P3_U3853, P3_U6158);
  nand ginst25017 (P3_U2842, P3_U3845, P3_U6134);
  nand ginst25018 (P3_U2843, P3_U6109, P3_U6110, P3_U6111);
  nand ginst25019 (P3_U2844, P3_U6085, P3_U6086, P3_U6087);
  nand ginst25020 (P3_U2845, P3_U6061, P3_U6062, P3_U6063);
  nand ginst25021 (P3_U2846, P3_U6037, P3_U6038, P3_U6039);
  nand ginst25022 (P3_U2847, P3_U3811, P3_U6014);
  nand ginst25023 (P3_U2848, P3_U3803, P3_U5990);
  nand ginst25024 (P3_U2849, P3_U5965, P3_U5966, P3_U5967);
  nand ginst25025 (P3_U2850, P3_U5941, P3_U5942, P3_U5943);
  nand ginst25026 (P3_U2851, P3_U5917, P3_U5918, P3_U5919);
  nand ginst25027 (P3_U2852, P3_U5893, P3_U5894, P3_U5895);
  nand ginst25028 (P3_U2853, P3_U5869, P3_U5870, P3_U5871);
  nand ginst25029 (P3_U2854, P3_U5845, P3_U5846, P3_U5847);
  nand ginst25030 (P3_U2855, P3_U5821, P3_U5822, P3_U5823);
  nand ginst25031 (P3_U2856, P3_U5797, P3_U5798, P3_U5799);
  nand ginst25032 (P3_U2857, P3_U5773, P3_U5774, P3_U5775);
  nand ginst25033 (P3_U2858, P3_U5749, P3_U5750, P3_U5751);
  nand ginst25034 (P3_U2859, P3_U5725, P3_U5726, P3_U5727);
  nand ginst25035 (P3_U2860, P3_U5701, P3_U5702, P3_U5703);
  nand ginst25036 (P3_U2861, P3_U5677, P3_U5678, P3_U5679);
  nand ginst25037 (P3_U2862, P3_U5653, P3_U5654, P3_U5655);
  nand ginst25038 (P3_U2863, P3_U5615, P3_U5616);
  nand ginst25039 (P3_U2864, P3_U5609, P3_U5610);
  nand ginst25040 (P3_U2865, P3_U5598, P3_U5599);
  nand ginst25041 (P3_U2866, P3_U5590, P3_U5591);
  and ginst25042 (P3_U2867, P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN, P3_U5579);
  nand ginst25043 (P3_U2868, P3_U3651, P3_U5482);
  nand ginst25044 (P3_U2869, P3_U3649, P3_U5477);
  nand ginst25045 (P3_U2870, P3_U3647, P3_U5472);
  nand ginst25046 (P3_U2871, P3_U3645, P3_U5467);
  nand ginst25047 (P3_U2872, P3_U3643, P3_U5462);
  nand ginst25048 (P3_U2873, P3_U3641, P3_U5457);
  nand ginst25049 (P3_U2874, P3_U3639, P3_U5452);
  nand ginst25050 (P3_U2875, P3_U3637, P3_U5447);
  nand ginst25051 (P3_U2876, P3_U3633, P3_U5432);
  nand ginst25052 (P3_U2877, P3_U3631, P3_U5427);
  nand ginst25053 (P3_U2878, P3_U3629, P3_U5422);
  nand ginst25054 (P3_U2879, P3_U3627, P3_U5417);
  nand ginst25055 (P3_U2880, P3_U3625, P3_U5412);
  nand ginst25056 (P3_U2881, P3_U3623, P3_U5407);
  nand ginst25057 (P3_U2882, P3_U3621, P3_U5402);
  nand ginst25058 (P3_U2883, P3_U3619, P3_U5397);
  nand ginst25059 (P3_U2884, P3_U3615, P3_U5381);
  nand ginst25060 (P3_U2885, P3_U3613, P3_U5376);
  nand ginst25061 (P3_U2886, P3_U3611, P3_U5371);
  nand ginst25062 (P3_U2887, P3_U3609, P3_U5366);
  nand ginst25063 (P3_U2888, P3_U3607, P3_U5361);
  nand ginst25064 (P3_U2889, P3_U3605, P3_U5356);
  nand ginst25065 (P3_U2890, P3_U3603, P3_U5351);
  nand ginst25066 (P3_U2891, P3_U3601, P3_U5346);
  nand ginst25067 (P3_U2892, P3_U3598, P3_U5330);
  nand ginst25068 (P3_U2893, P3_U3596, P3_U5325);
  nand ginst25069 (P3_U2894, P3_U3594, P3_U5320);
  nand ginst25070 (P3_U2895, P3_U3592, P3_U5315);
  nand ginst25071 (P3_U2896, P3_U3590, P3_U5310);
  nand ginst25072 (P3_U2897, P3_U3588, P3_U5305);
  nand ginst25073 (P3_U2898, P3_U3586, P3_U5300);
  nand ginst25074 (P3_U2899, P3_U3584, P3_U5295);
  nand ginst25075 (P3_U2900, P3_U3580, P3_U5279);
  nand ginst25076 (P3_U2901, P3_U3578, P3_U5274);
  nand ginst25077 (P3_U2902, P3_U3576, P3_U5269);
  nand ginst25078 (P3_U2903, P3_U3574, P3_U5264);
  nand ginst25079 (P3_U2904, P3_U3572, P3_U5259);
  nand ginst25080 (P3_U2905, P3_U3570, P3_U5254);
  nand ginst25081 (P3_U2906, P3_U3568, P3_U5249);
  nand ginst25082 (P3_U2907, P3_U3566, P3_U5244);
  nand ginst25083 (P3_U2908, P3_U3562, P3_U5228, P3_U5229);
  nand ginst25084 (P3_U2909, P3_U3560, P3_U5223, P3_U5224);
  nand ginst25085 (P3_U2910, P3_U3558, P3_U5218, P3_U5219);
  nand ginst25086 (P3_U2911, P3_U3556, P3_U5213, P3_U5214);
  nand ginst25087 (P3_U2912, P3_U3554, P3_U5208, P3_U5209);
  nand ginst25088 (P3_U2913, P3_U3552, P3_U5203, P3_U5204);
  nand ginst25089 (P3_U2914, P3_U3550, P3_U5198, P3_U5199);
  nand ginst25090 (P3_U2915, P3_U3548, P3_U5193, P3_U5194);
  nand ginst25091 (P3_U2916, P3_U3544, P3_U5176, P3_U5177);
  nand ginst25092 (P3_U2917, P3_U3542, P3_U5171, P3_U5172);
  nand ginst25093 (P3_U2918, P3_U3540, P3_U5166, P3_U5167);
  nand ginst25094 (P3_U2919, P3_U3538, P3_U5161, P3_U5162);
  nand ginst25095 (P3_U2920, P3_U3536, P3_U5156, P3_U5157);
  nand ginst25096 (P3_U2921, P3_U3534, P3_U5151, P3_U5152);
  nand ginst25097 (P3_U2922, P3_U3532, P3_U5146, P3_U5147);
  nand ginst25098 (P3_U2923, P3_U3530, P3_U5141, P3_U5142);
  nand ginst25099 (P3_U2924, P3_U3526, P3_U5124, P3_U5125);
  nand ginst25100 (P3_U2925, P3_U3524, P3_U5119, P3_U5120);
  nand ginst25101 (P3_U2926, P3_U3522, P3_U5114, P3_U5115);
  nand ginst25102 (P3_U2927, P3_U3520, P3_U5109, P3_U5110);
  nand ginst25103 (P3_U2928, P3_U3518, P3_U5104, P3_U5105);
  nand ginst25104 (P3_U2929, P3_U3516, P3_U5099, P3_U5100);
  nand ginst25105 (P3_U2930, P3_U3514, P3_U5094, P3_U5095);
  nand ginst25106 (P3_U2931, P3_U3512, P3_U5089, P3_U5090);
  nand ginst25107 (P3_U2932, P3_U3509, P3_U5075, P3_U5076);
  nand ginst25108 (P3_U2933, P3_U3507, P3_U5070, P3_U5071);
  nand ginst25109 (P3_U2934, P3_U3505, P3_U5065, P3_U5066);
  nand ginst25110 (P3_U2935, P3_U3503, P3_U5060, P3_U5061);
  nand ginst25111 (P3_U2936, P3_U3501, P3_U5055, P3_U5056);
  nand ginst25112 (P3_U2937, P3_U3499, P3_U5050, P3_U5051);
  nand ginst25113 (P3_U2938, P3_U3497, P3_U5045, P3_U5046);
  nand ginst25114 (P3_U2939, P3_U3495, P3_U5040, P3_U5041);
  nand ginst25115 (P3_U2940, P3_U3492, P3_U5024, P3_U5025);
  nand ginst25116 (P3_U2941, P3_U3490, P3_U5019, P3_U5020);
  nand ginst25117 (P3_U2942, P3_U3488, P3_U5014, P3_U5015);
  nand ginst25118 (P3_U2943, P3_U3486, P3_U5009, P3_U5010);
  nand ginst25119 (P3_U2944, P3_U3484, P3_U5004, P3_U5005);
  nand ginst25120 (P3_U2945, P3_U3482, P3_U4999, P3_U5000);
  nand ginst25121 (P3_U2946, P3_U3480, P3_U4994, P3_U4995);
  nand ginst25122 (P3_U2947, P3_U3478, P3_U4989, P3_U4990);
  nand ginst25123 (P3_U2948, P3_U3474, P3_U4972, P3_U4973);
  nand ginst25124 (P3_U2949, P3_U3472, P3_U4967, P3_U4968);
  nand ginst25125 (P3_U2950, P3_U3470, P3_U4962, P3_U4963);
  nand ginst25126 (P3_U2951, P3_U3468, P3_U4957, P3_U4958);
  nand ginst25127 (P3_U2952, P3_U3466, P3_U4952, P3_U4953);
  nand ginst25128 (P3_U2953, P3_U3464, P3_U4947, P3_U4948);
  nand ginst25129 (P3_U2954, P3_U3462, P3_U4942, P3_U4943);
  nand ginst25130 (P3_U2955, P3_U3460, P3_U4937, P3_U4938);
  nand ginst25131 (P3_U2956, P3_U3456, P3_U4920, P3_U4921);
  nand ginst25132 (P3_U2957, P3_U3454, P3_U4915, P3_U4916);
  nand ginst25133 (P3_U2958, P3_U3452, P3_U4910, P3_U4911);
  nand ginst25134 (P3_U2959, P3_U3450, P3_U4905, P3_U4906);
  nand ginst25135 (P3_U2960, P3_U3448, P3_U4900, P3_U4901);
  nand ginst25136 (P3_U2961, P3_U3446, P3_U4895, P3_U4896);
  nand ginst25137 (P3_U2962, P3_U3444, P3_U4890, P3_U4891);
  nand ginst25138 (P3_U2963, P3_U3442, P3_U4885, P3_U4886);
  nand ginst25139 (P3_U2964, P3_U3439, P3_U4868, P3_U4869);
  nand ginst25140 (P3_U2965, P3_U3437, P3_U4863, P3_U4864);
  nand ginst25141 (P3_U2966, P3_U3435, P3_U4858, P3_U4859);
  nand ginst25142 (P3_U2967, P3_U3433, P3_U4853, P3_U4854);
  nand ginst25143 (P3_U2968, P3_U3431, P3_U4848, P3_U4849);
  nand ginst25144 (P3_U2969, P3_U3429, P3_U4843, P3_U4844);
  nand ginst25145 (P3_U2970, P3_U3427, P3_U4838, P3_U4839);
  nand ginst25146 (P3_U2971, P3_U3425, P3_U4833, P3_U4834);
  nand ginst25147 (P3_U2972, P3_U3421, P3_U4817, P3_U4818);
  nand ginst25148 (P3_U2973, P3_U3419, P3_U4812, P3_U4813);
  nand ginst25149 (P3_U2974, P3_U3417, P3_U4807, P3_U4808);
  nand ginst25150 (P3_U2975, P3_U3415, P3_U4802, P3_U4803);
  nand ginst25151 (P3_U2976, P3_U3413, P3_U4797, P3_U4798);
  nand ginst25152 (P3_U2977, P3_U3411, P3_U4792, P3_U4793);
  nand ginst25153 (P3_U2978, P3_U3409, P3_U4787, P3_U4788);
  nand ginst25154 (P3_U2979, P3_U3407, P3_U4782, P3_U4783);
  nand ginst25155 (P3_U2980, P3_U3403, P3_U4765, P3_U4766);
  nand ginst25156 (P3_U2981, P3_U3401, P3_U4760, P3_U4761);
  nand ginst25157 (P3_U2982, P3_U3399, P3_U4755, P3_U4756);
  nand ginst25158 (P3_U2983, P3_U3397, P3_U4750, P3_U4751);
  nand ginst25159 (P3_U2984, P3_U3395, P3_U4745, P3_U4746);
  nand ginst25160 (P3_U2985, P3_U3393, P3_U4740, P3_U4741);
  nand ginst25161 (P3_U2986, P3_U3391, P3_U4735, P3_U4736);
  nand ginst25162 (P3_U2987, P3_U3389, P3_U4730, P3_U4731);
  nand ginst25163 (P3_U2988, P3_U3385, P3_U4713, P3_U4714);
  nand ginst25164 (P3_U2989, P3_U3383, P3_U4708, P3_U4709);
  nand ginst25165 (P3_U2990, P3_U3381, P3_U4703, P3_U4704);
  nand ginst25166 (P3_U2991, P3_U3379, P3_U4698, P3_U4699);
  nand ginst25167 (P3_U2992, P3_U3377, P3_U4693, P3_U4694);
  nand ginst25168 (P3_U2993, P3_U3375, P3_U4688, P3_U4689);
  nand ginst25169 (P3_U2994, P3_U3373, P3_U4683, P3_U4684);
  nand ginst25170 (P3_U2995, P3_U3371, P3_U4678, P3_U4679);
  nand ginst25171 (P3_U2996, P3_U3367, P3_U7958, P3_U7959);
  nand ginst25172 (P3_U2997, P3_U4329, P3_U4634, P3_U4635, P3_U4636);
  nand ginst25173 (P3_U2998, P3_U3363, P3_U4632);
  and ginst25174 (P3_U2999, P3_DATAWIDTH_REG_31__SCAN_IN, P3_U7937);
  and ginst25175 (P3_U3000, P3_DATAWIDTH_REG_30__SCAN_IN, P3_U7937);
  and ginst25176 (P3_U3001, P3_DATAWIDTH_REG_29__SCAN_IN, P3_U7937);
  and ginst25177 (P3_U3002, P3_DATAWIDTH_REG_28__SCAN_IN, P3_U7937);
  and ginst25178 (P3_U3003, P3_DATAWIDTH_REG_27__SCAN_IN, P3_U7937);
  and ginst25179 (P3_U3004, P3_DATAWIDTH_REG_26__SCAN_IN, P3_U7937);
  and ginst25180 (P3_U3005, P3_DATAWIDTH_REG_25__SCAN_IN, P3_U7937);
  and ginst25181 (P3_U3006, P3_DATAWIDTH_REG_24__SCAN_IN, P3_U7937);
  and ginst25182 (P3_U3007, P3_DATAWIDTH_REG_23__SCAN_IN, P3_U7937);
  and ginst25183 (P3_U3008, P3_DATAWIDTH_REG_22__SCAN_IN, P3_U7937);
  and ginst25184 (P3_U3009, P3_DATAWIDTH_REG_21__SCAN_IN, P3_U7937);
  and ginst25185 (P3_U3010, P3_DATAWIDTH_REG_20__SCAN_IN, P3_U7937);
  and ginst25186 (P3_U3011, P3_DATAWIDTH_REG_19__SCAN_IN, P3_U7937);
  and ginst25187 (P3_U3012, P3_DATAWIDTH_REG_18__SCAN_IN, P3_U7937);
  and ginst25188 (P3_U3013, P3_DATAWIDTH_REG_17__SCAN_IN, P3_U7937);
  and ginst25189 (P3_U3014, P3_DATAWIDTH_REG_16__SCAN_IN, P3_U7937);
  and ginst25190 (P3_U3015, P3_DATAWIDTH_REG_15__SCAN_IN, P3_U7937);
  and ginst25191 (P3_U3016, P3_DATAWIDTH_REG_14__SCAN_IN, P3_U7937);
  and ginst25192 (P3_U3017, P3_DATAWIDTH_REG_13__SCAN_IN, P3_U7937);
  and ginst25193 (P3_U3018, P3_DATAWIDTH_REG_12__SCAN_IN, P3_U7937);
  and ginst25194 (P3_U3019, P3_DATAWIDTH_REG_11__SCAN_IN, P3_U7937);
  and ginst25195 (P3_U3020, P3_DATAWIDTH_REG_10__SCAN_IN, P3_U7937);
  and ginst25196 (P3_U3021, P3_DATAWIDTH_REG_9__SCAN_IN, P3_U7937);
  and ginst25197 (P3_U3022, P3_DATAWIDTH_REG_8__SCAN_IN, P3_U7937);
  and ginst25198 (P3_U3023, P3_DATAWIDTH_REG_7__SCAN_IN, P3_U7937);
  and ginst25199 (P3_U3024, P3_DATAWIDTH_REG_6__SCAN_IN, P3_U7937);
  and ginst25200 (P3_U3025, P3_DATAWIDTH_REG_5__SCAN_IN, P3_U7937);
  and ginst25201 (P3_U3026, P3_DATAWIDTH_REG_4__SCAN_IN, P3_U7937);
  and ginst25202 (P3_U3027, P3_DATAWIDTH_REG_3__SCAN_IN, P3_U7937);
  and ginst25203 (P3_U3028, P3_DATAWIDTH_REG_2__SCAN_IN, P3_U7937);
  nand ginst25204 (P3_U3029, P3_U4463, P3_U7933, P3_U7934);
  nand ginst25205 (P3_U3030, P3_U3311, P3_U7931, P3_U7932);
  nand ginst25206 (P3_U3031, P3_U3310, P3_U4457);
  nand ginst25207 (P3_U3032, P3_U4442, P3_U4443, P3_U4444);
  nand ginst25208 (P3_U3033, P3_U4439, P3_U4440, P3_U4441);
  nand ginst25209 (P3_U3034, P3_U4436, P3_U4437, P3_U4438);
  nand ginst25210 (P3_U3035, P3_U4433, P3_U4434, P3_U4435);
  nand ginst25211 (P3_U3036, P3_U4430, P3_U4431, P3_U4432);
  nand ginst25212 (P3_U3037, P3_U4427, P3_U4428, P3_U4429);
  nand ginst25213 (P3_U3038, P3_U4424, P3_U4425, P3_U4426);
  nand ginst25214 (P3_U3039, P3_U4421, P3_U4422, P3_U4423);
  nand ginst25215 (P3_U3040, P3_U4418, P3_U4419, P3_U4420);
  nand ginst25216 (P3_U3041, P3_U4415, P3_U4416, P3_U4417);
  nand ginst25217 (P3_U3042, P3_U4412, P3_U4413, P3_U4414);
  nand ginst25218 (P3_U3043, P3_U4409, P3_U4410, P3_U4411);
  nand ginst25219 (P3_U3044, P3_U4406, P3_U4407, P3_U4408);
  nand ginst25220 (P3_U3045, P3_U4403, P3_U4404, P3_U4405);
  nand ginst25221 (P3_U3046, P3_U4400, P3_U4401, P3_U4402);
  nand ginst25222 (P3_U3047, P3_U4397, P3_U4398, P3_U4399);
  nand ginst25223 (P3_U3048, P3_U4394, P3_U4395, P3_U4396);
  nand ginst25224 (P3_U3049, P3_U4391, P3_U4392, P3_U4393);
  nand ginst25225 (P3_U3050, P3_U4388, P3_U4389, P3_U4390);
  nand ginst25226 (P3_U3051, P3_U4385, P3_U4386, P3_U4387);
  nand ginst25227 (P3_U3052, P3_U4382, P3_U4383, P3_U4384);
  nand ginst25228 (P3_U3053, P3_U4379, P3_U4380, P3_U4381);
  nand ginst25229 (P3_U3054, P3_U4376, P3_U4377, P3_U4378);
  nand ginst25230 (P3_U3055, P3_U4373, P3_U4374, P3_U4375);
  nand ginst25231 (P3_U3056, P3_U4370, P3_U4371, P3_U4372);
  nand ginst25232 (P3_U3057, P3_U4367, P3_U4368, P3_U4369);
  nand ginst25233 (P3_U3058, P3_U4364, P3_U4365, P3_U4366);
  nand ginst25234 (P3_U3059, P3_U4361, P3_U4362, P3_U4363);
  nand ginst25235 (P3_U3060, P3_U4358, P3_U4359, P3_U4360);
  nand ginst25236 (P3_U3061, P3_U4355, P3_U4356, P3_U4357);
  nand ginst25237 (P3_U3062, P3_U4244, P3_U4245, P3_U4246, P3_U4247);
  nand ginst25238 (P3_U3063, P3_U4240, P3_U4241, P3_U4242, P3_U4243);
  nand ginst25239 (P3_U3064, P3_U4236, P3_U4237, P3_U4238, P3_U4239);
  nand ginst25240 (P3_U3065, P3_U4232, P3_U4233, P3_U4234, P3_U4235);
  nand ginst25241 (P3_U3066, P3_U4228, P3_U4229, P3_U4230, P3_U4231);
  nand ginst25242 (P3_U3067, P3_U4224, P3_U4225, P3_U4226, P3_U4227);
  nand ginst25243 (P3_U3068, P3_U4220, P3_U4221, P3_U4222, P3_U4223);
  nand ginst25244 (P3_U3069, P3_U4216, P3_U4217, P3_U4218, P3_U4219);
  nand ginst25245 (P3_U3070, P3_U2457, P3_U4642);
  nand ginst25246 (P3_U3071, P3_U2459, P3_U4642);
  nand ginst25247 (P3_U3072, P3_U2458, P3_U4642);
  nand ginst25248 (P3_U3073, P3_U2460, P3_U4642);
  nand ginst25249 (P3_U3074, P3_U3343, P3_U3344, P3_U3345, P3_U3346, P3_U3347);
  not ginst25250 (P3_U3075, P3_REQUESTPENDING_REG_SCAN_IN);
  not ginst25251 (P3_U3076, P3_STATE_REG_1__SCAN_IN);
  nand ginst25252 (P3_U3077, P3_STATE_REG_1__SCAN_IN, P3_U3085);
  nand ginst25253 (P3_U3078, P3_U3079, P3_U4308);
  not ginst25254 (P3_U3079, P3_STATE_REG_2__SCAN_IN);
  nand ginst25255 (P3_U3080, P3_STATE_REG_2__SCAN_IN, P3_U4308);
  not ginst25256 (P3_U3081, P3_REIP_REG_1__SCAN_IN);
  nand ginst25257 (P3_U3082, P3_STATE_REG_1__SCAN_IN, P3_U3079);
  or ginst25258 (P3_U3083, P3_STATE_REG_2__SCAN_IN, P3_STATE_REG_1__SCAN_IN);
  not ginst25259 (P3_U3084, HOLD);
  not ginst25260 (P3_U3085, P3_STATE_REG_0__SCAN_IN);
  nand ginst25261 (P3_U3086, P3_STATE_REG_0__SCAN_IN, P3_U3087);
  nand ginst25262 (P3_U3087, P3_REQUESTPENDING_REG_SCAN_IN, P3_U3084);
  or ginst25263 (P3_U3088, HOLD, P3_REQUESTPENDING_REG_SCAN_IN);
  not ginst25264 (P3_U3089, P3_STATE2_REG_1__SCAN_IN);
  not ginst25265 (P3_U3090, P3_STATE2_REG_2__SCAN_IN);
  or ginst25266 (P3_U3091, P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN);
  nand ginst25267 (P3_U3092, P3_U3097, P3_U4467);
  not ginst25268 (P3_U3093, P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN);
  not ginst25269 (P3_U3094, P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN);
  nand ginst25270 (P3_U3095, P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN);
  nand ginst25271 (P3_U3096, P3_U3097, P3_U4332);
  not ginst25272 (P3_U3097, P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN);
  nand ginst25273 (P3_U3098, P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN, P3_U3100);
  nand ginst25274 (P3_U3099, P3_U4332, P3_U4470);
  not ginst25275 (P3_U3100, P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN);
  nand ginst25276 (P3_U3101, P3_U3338, P3_U3339, P3_U3340, P3_U3341, P3_U3342);
  nand ginst25277 (P3_U3102, P3_U3323, P3_U3324, P3_U3325, P3_U3326, P3_U3327);
  nand ginst25278 (P3_U3103, P3_U3074, P3_U3110);
  nand ginst25279 (P3_U3104, P3_U3318, P3_U3319, P3_U3320, P3_U3321, P3_U3322);
  nand ginst25280 (P3_U3105, P3_U3085, P3_U4466);
  nand ginst25281 (P3_U3106, P3_U2630, P3_U4293);
  nand ginst25282 (P3_U3107, P3_U3328, P3_U3329, P3_U3330, P3_U3331, P3_U3332);
  nand ginst25283 (P3_U3108, P3_U3313, P3_U3314, P3_U3315, P3_U3316, P3_U3317);
  nand ginst25284 (P3_U3109, P3_U2353, P3_U4488);
  nand ginst25285 (P3_U3110, P3_U3348, P3_U3349, P3_U3350, P3_U3351, P3_U3352);
  nand ginst25286 (P3_U3111, P3_U3104, P3_U3108);
  nand ginst25287 (P3_U3112, P3_U3108, P3_U4505);
  nand ginst25288 (P3_U3113, P3_U3110, P3_U4607);
  nand ginst25289 (P3_U3114, P3_U4488, P3_U4505);
  nand ginst25290 (P3_U3115, P3_U2451, P3_U4297);
  nand ginst25291 (P3_U3116, P3_U2452, P3_U4297);
  nand ginst25292 (P3_U3117, P3_U2452, P3_U4296);
  nand ginst25293 (P3_U3118, P3_U3104, P3_U4488);
  nand ginst25294 (P3_U3119, P3_U2353, P3_U3356);
  nand ginst25295 (P3_U3120, P3_LT_563_U6, P3_U3262, P3_U4313, P3_U7948, P3_U7949);
  not ginst25296 (P3_U3121, P3_STATE2_REG_0__SCAN_IN);
  nand ginst25297 (P3_U3122, P3_STATE2_REG_0__SCAN_IN, P3_U4629);
  or ginst25298 (P3_U3123, P3_STATE2_REG_3__SCAN_IN, P3_STATE2_REG_1__SCAN_IN);
  nand ginst25299 (P3_U3124, P3_STATE2_REG_2__SCAN_IN, P3_U3089);
  or ginst25300 (P3_U3125, P3_STATE2_REG_2__SCAN_IN, P3_STATE2_REG_1__SCAN_IN);
  nand ginst25301 (P3_U3126, P3_STATE2_REG_3__SCAN_IN, P3_LTE_597_U6);
  nand ginst25302 (P3_U3127, P3_U3121, P3_U4666);
  not ginst25303 (P3_U3128, P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN);
  not ginst25304 (P3_U3129, P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN);
  nand ginst25305 (P3_U3130, P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN, P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN);
  not ginst25306 (P3_U3131, P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN);
  nand ginst25307 (P3_U3132, P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN, P3_U4648);
  not ginst25308 (P3_U3133, P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN);
  nand ginst25309 (P3_U3134, P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN, P3_U4649);
  or ginst25310 (P3_U3135, P3_STATE2_REG_3__SCAN_IN, P3_STATE2_REG_2__SCAN_IN);
  nand ginst25311 (P3_U3136, P3_STATEBS16_REG_SCAN_IN, P3_U4295);
  nand ginst25312 (P3_U3137, P3_U3153, P3_U4641);
  nand ginst25313 (P3_U3138, P3_U3128, P3_U3137);
  nand ginst25314 (P3_U3139, P3_U3180, P3_U4651);
  nand ginst25315 (P3_U3140, P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P3_U3141);
  nand ginst25316 (P3_U3141, P3_U3150, P3_U3158);
  nand ginst25317 (P3_U3142, P3_U4331, P3_U4655);
  nand ginst25318 (P3_U3143, P3_U3128, P3_U3156);
  nand ginst25319 (P3_U3144, P3_U2486, P3_U4647);
  nand ginst25320 (P3_U3145, P3_U3144, P3_U4667);
  nand ginst25321 (P3_U3146, P3_U3134, P3_U4663);
  nand ginst25322 (P3_U3147, P3_U2492, P3_U3386);
  nand ginst25323 (P3_U3148, P3_U3128, P3_U3141);
  nand ginst25324 (P3_U3149, P3_U2486, P3_U2490);
  nand ginst25325 (P3_U3150, P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P3_U3137);
  nand ginst25326 (P3_U3151, P3_U3149, P3_U4719);
  nand ginst25327 (P3_U3152, P3_U3147, P3_U4717);
  nand ginst25328 (P3_U3153, P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P3_U3129);
  nand ginst25329 (P3_U3154, P3_U3404, P3_U4640);
  nand ginst25330 (P3_U3155, P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P3_U4643);
  nand ginst25331 (P3_U3156, P3_U3148, P3_U3155);
  nand ginst25332 (P3_U3157, P3_U2486, P3_U2493);
  nand ginst25333 (P3_U3158, P3_U3128, P3_U4642);
  nand ginst25334 (P3_U3159, P3_U3157, P3_U4771);
  nand ginst25335 (P3_U3160, P3_U3154, P3_U4769);
  nand ginst25336 (P3_U3161, P3_U2492, P3_U3422);
  nand ginst25337 (P3_U3162, P3_U2486, P3_U2495);
  nand ginst25338 (P3_U3163, P3_U3162, P3_U4822);
  nand ginst25339 (P3_U3164, P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN, P3_U3131, P3_U4648);
  nand ginst25340 (P3_U3165, P3_U3142, P3_U7965);
  nand ginst25341 (P3_U3166, P3_U2498, P3_U4647);
  nand ginst25342 (P3_U3167, P3_U3166, P3_U4874);
  nand ginst25343 (P3_U3168, P3_U3164, P3_U4872);
  nand ginst25344 (P3_U3169, P3_U2501, P3_U3457);
  nand ginst25345 (P3_U3170, P3_U2490, P3_U2498);
  nand ginst25346 (P3_U3171, P3_U3170, P3_U4926);
  nand ginst25347 (P3_U3172, P3_U3169, P3_U4924);
  nand ginst25348 (P3_U3173, P3_U3475, P3_U4640);
  nand ginst25349 (P3_U3174, P3_U2493, P3_U2498);
  nand ginst25350 (P3_U3175, P3_U3174, P3_U4978);
  nand ginst25351 (P3_U3176, P3_U3173, P3_U4976);
  nand ginst25352 (P3_U3177, P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN, P3_U2501, P3_U3129);
  nand ginst25353 (P3_U3178, P3_U2495, P3_U2498);
  nand ginst25354 (P3_U3179, P3_U3178, P3_U5029);
  nand ginst25355 (P3_U3180, P3_U3133, P3_U4649);
  nand ginst25356 (P3_U3181, P3_U2485, P3_U4657);
  nand ginst25357 (P3_U3182, P3_U3181, P3_U3368);
  nand ginst25358 (P3_U3183, P3_U2504, P3_U4647);
  nand ginst25359 (P3_U3184, P3_U3181, P3_U3183);
  nand ginst25360 (P3_U3185, P3_U3180, P3_U4331);
  nand ginst25361 (P3_U3186, P3_U2492, P3_U3527);
  nand ginst25362 (P3_U3187, P3_U2490, P3_U2504);
  nand ginst25363 (P3_U3188, P3_U3187, P3_U5130);
  nand ginst25364 (P3_U3189, P3_U3186, P3_U5128);
  nand ginst25365 (P3_U3190, P3_U3545, P3_U4640);
  nand ginst25366 (P3_U3191, P3_U2493, P3_U2504);
  nand ginst25367 (P3_U3192, P3_U3191, P3_U5182);
  nand ginst25368 (P3_U3193, P3_U3190, P3_U5180);
  nand ginst25369 (P3_U3194, P3_U2492, P3_U3563);
  nand ginst25370 (P3_U3195, P3_U2495, P3_U2504);
  nand ginst25371 (P3_U3196, P3_U3581, P3_U4648);
  nand ginst25372 (P3_U3197, P3_U2508, P3_U4647);
  nand ginst25373 (P3_U3198, P3_U3196, P3_U5282);
  nand ginst25374 (P3_U3199, P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN, P3_U2501, P3_U3133);
  nand ginst25375 (P3_U3200, P3_U2490, P3_U2508);
  nand ginst25376 (P3_U3201, P3_U3199, P3_U5333);
  nand ginst25377 (P3_U3202, P3_U3616, P3_U4640);
  nand ginst25378 (P3_U3203, P3_U2493, P3_U2508);
  nand ginst25379 (P3_U3204, P3_U3202, P3_U5384);
  nand ginst25380 (P3_U3205, P3_U2501, P3_U3634);
  nand ginst25381 (P3_U3206, P3_U2495, P3_U2508);
  not ginst25382 (P3_U3207, P3_FLUSH_REG_SCAN_IN);
  nand ginst25383 (P3_U3208, P3_U3102, P3_U4539);
  nand ginst25384 (P3_U3209, P3_U2514, P3_U3113);
  not ginst25385 (P3_U3210, P3_GTE_412_U6);
  not ginst25386 (P3_U3211, P3_GTE_485_U6);
  not ginst25387 (P3_U3212, P3_GTE_390_U6);
  not ginst25388 (P3_U3213, P3_GTE_450_U6);
  not ginst25389 (P3_U3214, P3_GTE_504_U6);
  not ginst25390 (P3_U3215, P3_GTE_401_U6);
  nand ginst25391 (P3_U3216, P3_U3074, P3_U4590);
  nand ginst25392 (P3_U3217, P3_U2450, P3_U4323);
  nand ginst25393 (P3_U3218, P3_U3333, P3_U3334, P3_U3335, P3_U3336, P3_U3337);
  nand ginst25394 (P3_U3219, P3_U2461, P3_U3662);
  nand ginst25395 (P3_U3220, P3_U3667, P3_U7975, P3_U7976);
  nand ginst25396 (P3_U3221, P3_U3119, P3_U3222, P3_U5524);
  nand ginst25397 (P3_U3222, P3_U3218, P3_U4314);
  nand ginst25398 (P3_U3223, P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P3_U5503);
  nand ginst25399 (P3_U3224, P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P3_U5505);
  nand ginst25400 (P3_U3225, P3_U3096, P3_U3227);
  nand ginst25401 (P3_U3226, P3_U2517, P3_U3674);
  nand ginst25402 (P3_U3227, P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN, P3_U3095);
  nand ginst25403 (P3_U3228, P3_U3091, P3_U3095);
  nand ginst25404 (P3_U3229, P3_U3218, P3_U4323, P3_U4350);
  nand ginst25405 (P3_U3230, P3_U2518, P3_U3243);
  nand ginst25406 (P3_U3231, P3_U3115, P3_U5559);
  not ginst25407 (P3_U3232, P3_LT_589_U6);
  nand ginst25408 (P3_U3233, P3_U3127, P3_U4330, P3_U5578);
  nand ginst25409 (P3_U3234, P3_U3123, P3_U3135);
  nand ginst25410 (P3_U3235, P3_U3101, P3_U3104, P3_U4294);
  nand ginst25411 (P3_U3236, P3_U2630, P3_U3101, P3_U4505);
  not ginst25412 (P3_U3237, P3_GTE_370_U6);
  not ginst25413 (P3_U3238, P3_GTE_355_U6);
  nand ginst25414 (P3_U3239, P3_U3089, P3_U4295);
  not ginst25415 (P3_U3240, P3_REIP_REG_0__SCAN_IN);
  not ginst25416 (P3_U3241, P3_U2628);
  nand ginst25417 (P3_U3242, P3_U2450, P3_U3661);
  nand ginst25418 (P3_U3243, P3_U2461, P3_U4314);
  nand ginst25419 (P3_U3244, P3_U4352, P3_U4522);
  nand ginst25420 (P3_U3245, P3_U3102, P3_U4352);
  nand ginst25421 (P3_U3246, P3_U2449, P3_U3663, P3_U3664);
  nand ginst25422 (P3_U3247, P3_STATE2_REG_2__SCAN_IN, P3_U3248);
  nand ginst25423 (P3_U3248, P3_U4336, P3_U5630);
  nand ginst25424 (P3_U3249, P3_U6402, P3_U6403);
  nand ginst25425 (P3_U3250, P3_U2390, P3_U6663);
  nand ginst25426 (P3_U3251, P3_U6757, P3_U6758);
  nand ginst25427 (P3_U3252, P3_U2390, P3_U6853);
  nand ginst25428 (P3_U3253, P3_U2390, P3_U6997);
  nand ginst25429 (P3_U3254, P3_U5489, P3_U5490);
  nand ginst25430 (P3_U3255, P3_U5486, P3_U5487);
  not ginst25431 (P3_U3256, P3_EBX_REG_31__SCAN_IN);
  or ginst25432 (P3_U3257, P3_STATEBS16_REG_SCAN_IN, U209);
  not ginst25433 (P3_U3258, P3_ADD_318_U69);
  nand ginst25434 (P3_U3259, P3_ADD_318_U69, P3_U2385);
  nand ginst25435 (P3_U3260, P3_U4030, P3_U4334);
  nand ginst25436 (P3_U3261, P3_U4138, P3_U4141, P3_U4144, P3_U4148);
  nand ginst25437 (P3_U3262, P3_U2462, P3_U3108, P3_U4282);
  not ginst25438 (P3_U3263, P3_CODEFETCH_REG_SCAN_IN);
  not ginst25439 (P3_U3264, P3_READREQUEST_REG_SCAN_IN);
  nand ginst25440 (P3_U3265, P3_U3099, P3_U3224);
  nand ginst25441 (P3_U3266, P3_U3223, P3_U7515);
  nand ginst25442 (P3_U3267, P3_U3092, P3_U4289);
  nand ginst25443 (P3_U3268, P3_U3098, P3_U7774);
  nand ginst25444 (P3_U3269, P3_U7960, P3_U7961);
  nand ginst25445 (P3_U3270, P3_U7963, P3_U7964);
  nand ginst25446 (P3_U3271, P3_U7966, P3_U7967);
  nand ginst25447 (P3_U3272, P3_U8032, P3_U8033);
  nand ginst25448 (P3_U3273, P3_U8035, P3_U8036);
  nand ginst25449 (P3_U3274, P3_U7920, P3_U7921);
  nand ginst25450 (P3_U3275, P3_U7922, P3_U7923);
  nand ginst25451 (P3_U3276, P3_U7924, P3_U7925);
  nand ginst25452 (P3_U3277, P3_U7926, P3_U7927);
  nand ginst25453 (P3_U3278, P3_U7935, P3_U7936);
  and ginst25454 (P3_U3279, P3_U3083, P3_U4286);
  nand ginst25455 (P3_U3280, P3_U7938, P3_U7939);
  nand ginst25456 (P3_U3281, P3_U7940, P3_U7941);
  nand ginst25457 (P3_U3282, P3_U7954, P3_U7955);
  and ginst25458 (P3_U3283, P3_U2356, P3_U3652);
  nand ginst25459 (P3_U3284, P3_U7971, P3_U7972);
  nand ginst25460 (P3_U3285, P3_U7979, P3_U7980);
  nand ginst25461 (P3_U3286, P3_U7986, P3_U7987);
  nand ginst25462 (P3_U3287, P3_U7983, P3_U7984);
  nand ginst25463 (P3_U3288, P3_U7989, P3_U7990);
  nand ginst25464 (P3_U3289, P3_U7991, P3_U7992);
  nand ginst25465 (P3_U3290, P3_U7995, P3_U7996);
  nor ginst25466 (P3_U3291, P3_DATAWIDTH_REG_1__SCAN_IN, P3_REIP_REG_1__SCAN_IN);
  nand ginst25467 (P3_U3292, P3_U8010, P3_U8011);
  nand ginst25468 (P3_U3293, P3_U8014, P3_U8015);
  nand ginst25469 (P3_U3294, P3_U8016, P3_U8017);
  nand ginst25470 (P3_U3295, P3_U8018, P3_U8019);
  nand ginst25471 (P3_U3296, P3_U8022, P3_U8023);
  nand ginst25472 (P3_U3297, P3_U8026, P3_U8027);
  nand ginst25473 (P3_U3298, P3_U8028, P3_U8029);
  nand ginst25474 (P3_U3299, P3_U8030, P3_U8031);
  nand ginst25475 (P3_U3300, P3_U8038, P3_U8039);
  nand ginst25476 (P3_U3301, P3_U8040, P3_U8041);
  nand ginst25477 (P3_U3302, P3_U8042, P3_U8043);
  and ginst25478 (P3_U3303, P3_ADD_495_U8, P3_U2356);
  nand ginst25479 (P3_U3304, P3_U8044, P3_U8045);
  nand ginst25480 (P3_U3305, P3_U8046, P3_U8047);
  nand ginst25481 (P3_U3306, P3_U8048, P3_U8049);
  nand ginst25482 (P3_U3307, P3_U8050, P3_U8051);
  nand ginst25483 (P3_U3308, P3_U8052, P3_U8053);
  and ginst25484 (P3_U3309, P3_STATE_REG_0__SCAN_IN, P3_U4447);
  and ginst25485 (P3_U3310, P3_U3080, P3_U4456);
  and ginst25486 (P3_U3311, P3_U3078, P3_U4458);
  and ginst25487 (P3_U3312, P3_STATE_REG_0__SCAN_IN, P3_REQUESTPENDING_REG_SCAN_IN);
  and ginst25488 (P3_U3313, P3_U4472, P3_U4473, P3_U4474, P3_U4475);
  and ginst25489 (P3_U3314, P3_U4476, P3_U4477, P3_U4478, P3_U4479);
  and ginst25490 (P3_U3315, P3_U4480, P3_U4481);
  and ginst25491 (P3_U3316, P3_U4482, P3_U4483);
  and ginst25492 (P3_U3317, P3_U4484, P3_U4485, P3_U4486, P3_U4487);
  and ginst25493 (P3_U3318, P3_U4489, P3_U4490, P3_U4491, P3_U4492);
  and ginst25494 (P3_U3319, P3_U4493, P3_U4494, P3_U4495, P3_U4496);
  and ginst25495 (P3_U3320, P3_U4497, P3_U4498);
  and ginst25496 (P3_U3321, P3_U4499, P3_U4500);
  and ginst25497 (P3_U3322, P3_U4501, P3_U4502, P3_U4503, P3_U4504);
  and ginst25498 (P3_U3323, P3_U4506, P3_U4507, P3_U4508, P3_U4509);
  and ginst25499 (P3_U3324, P3_U4510, P3_U4511, P3_U4512, P3_U4513);
  and ginst25500 (P3_U3325, P3_U4514, P3_U4515);
  and ginst25501 (P3_U3326, P3_U4516, P3_U4517);
  and ginst25502 (P3_U3327, P3_U4518, P3_U4519, P3_U4520, P3_U4521);
  and ginst25503 (P3_U3328, P3_U4540, P3_U4541, P3_U4542, P3_U4543);
  and ginst25504 (P3_U3329, P3_U4544, P3_U4545, P3_U4546, P3_U4547);
  and ginst25505 (P3_U3330, P3_U4548, P3_U4549);
  and ginst25506 (P3_U3331, P3_U4550, P3_U4551);
  and ginst25507 (P3_U3332, P3_U4552, P3_U4553, P3_U4554, P3_U4555);
  and ginst25508 (P3_U3333, P3_U4557, P3_U4558, P3_U4559, P3_U4560);
  and ginst25509 (P3_U3334, P3_U4561, P3_U4562, P3_U4563, P3_U4564);
  and ginst25510 (P3_U3335, P3_U4565, P3_U4566);
  and ginst25511 (P3_U3336, P3_U4567, P3_U4568);
  and ginst25512 (P3_U3337, P3_U4569, P3_U4570, P3_U4571, P3_U4572);
  and ginst25513 (P3_U3338, P3_U4523, P3_U4524, P3_U4525, P3_U4526);
  and ginst25514 (P3_U3339, P3_U4527, P3_U4528, P3_U4529, P3_U4530);
  and ginst25515 (P3_U3340, P3_U4531, P3_U4532);
  and ginst25516 (P3_U3341, P3_U4533, P3_U4534);
  and ginst25517 (P3_U3342, P3_U4535, P3_U4536, P3_U4537, P3_U4538);
  and ginst25518 (P3_U3343, P3_U4591, P3_U4592, P3_U4593, P3_U4594);
  and ginst25519 (P3_U3344, P3_U4595, P3_U4596, P3_U4597, P3_U4598);
  and ginst25520 (P3_U3345, P3_U4599, P3_U4600);
  and ginst25521 (P3_U3346, P3_U4601, P3_U4602);
  and ginst25522 (P3_U3347, P3_U4603, P3_U4604, P3_U4605, P3_U4606);
  and ginst25523 (P3_U3348, P3_U4574, P3_U4575, P3_U4576, P3_U4577);
  and ginst25524 (P3_U3349, P3_U4578, P3_U4579, P3_U4580, P3_U4581);
  and ginst25525 (P3_U3350, P3_U4582, P3_U4583);
  and ginst25526 (P3_U3351, P3_U4584, P3_U4585);
  and ginst25527 (P3_U3352, P3_U4586, P3_U4587, P3_U4588, P3_U4589);
  and ginst25528 (P3_U3353, P3_U2352, P3_U4293);
  and ginst25529 (P3_U3354, P3_U3218, P3_U4556);
  and ginst25530 (P3_U3355, P3_U3101, P3_U4323);
  and ginst25531 (P3_U3356, P3_U3101, P3_U4324);
  and ginst25532 (P3_U3357, P3_U4609, P3_U4610, P3_U4611, P3_U4612);
  and ginst25533 (P3_U3358, P3_U4613, P3_U4614, P3_U4615, P3_U4616);
  and ginst25534 (P3_U3359, P3_U2630, P3_U4539);
  and ginst25535 (P3_U3360, P3_U3107, P3_U3108, P3_U3218);
  and ginst25536 (P3_U3361, P3_U3235, P3_U3236, P3_U4621);
  and ginst25537 (P3_U3362, P3_U3089, P3_U4626);
  and ginst25538 (P3_U3363, P3_U3124, P3_U4631);
  and ginst25539 (P3_U3364, P3_U2630, P3_U4340);
  and ginst25540 (P3_U3365, P3_STATE2_REG_3__SCAN_IN, P3_STATE2_REG_0__SCAN_IN);
  and ginst25541 (P3_U3366, P3_U4328, P3_U4338);
  and ginst25542 (P3_U3367, P3_U3366, P3_U4639);
  and ginst25543 (P3_U3368, P3_U3165, P3_U4659);
  and ginst25544 (P3_U3369, P3_U4312, P3_U4671);
  and ginst25545 (P3_U3370, P3_U4675, P3_U4676);
  and ginst25546 (P3_U3371, P3_U3370, P3_U4677);
  and ginst25547 (P3_U3372, P3_U4680, P3_U4681);
  and ginst25548 (P3_U3373, P3_U3372, P3_U4682);
  and ginst25549 (P3_U3374, P3_U4685, P3_U4686);
  and ginst25550 (P3_U3375, P3_U3374, P3_U4687);
  and ginst25551 (P3_U3376, P3_U4690, P3_U4691);
  and ginst25552 (P3_U3377, P3_U3376, P3_U4692);
  and ginst25553 (P3_U3378, P3_U4695, P3_U4696);
  and ginst25554 (P3_U3379, P3_U3378, P3_U4697);
  and ginst25555 (P3_U3380, P3_U4700, P3_U4701);
  and ginst25556 (P3_U3381, P3_U3380, P3_U4702);
  and ginst25557 (P3_U3382, P3_U4705, P3_U4706);
  and ginst25558 (P3_U3383, P3_U3382, P3_U4707);
  and ginst25559 (P3_U3384, P3_U4710, P3_U4711);
  and ginst25560 (P3_U3385, P3_U3384, P3_U4712);
  and ginst25561 (P3_U3386, P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN, P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN);
  and ginst25562 (P3_U3387, P3_U4312, P3_U4723);
  and ginst25563 (P3_U3388, P3_U4727, P3_U4728);
  and ginst25564 (P3_U3389, P3_U3388, P3_U4729);
  and ginst25565 (P3_U3390, P3_U4732, P3_U4733);
  and ginst25566 (P3_U3391, P3_U3390, P3_U4734);
  and ginst25567 (P3_U3392, P3_U4737, P3_U4738);
  and ginst25568 (P3_U3393, P3_U3392, P3_U4739);
  and ginst25569 (P3_U3394, P3_U4742, P3_U4743);
  and ginst25570 (P3_U3395, P3_U3394, P3_U4744);
  and ginst25571 (P3_U3396, P3_U4747, P3_U4748);
  and ginst25572 (P3_U3397, P3_U3396, P3_U4749);
  and ginst25573 (P3_U3398, P3_U4752, P3_U4753);
  and ginst25574 (P3_U3399, P3_U3398, P3_U4754);
  and ginst25575 (P3_U3400, P3_U4757, P3_U4758);
  and ginst25576 (P3_U3401, P3_U3400, P3_U4759);
  and ginst25577 (P3_U3402, P3_U4762, P3_U4763);
  and ginst25578 (P3_U3403, P3_U3402, P3_U4764);
  and ginst25579 (P3_U3404, P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN, P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN);
  and ginst25580 (P3_U3405, P3_U4312, P3_U4775);
  and ginst25581 (P3_U3406, P3_U4779, P3_U4780);
  and ginst25582 (P3_U3407, P3_U3406, P3_U4781);
  and ginst25583 (P3_U3408, P3_U4784, P3_U4785);
  and ginst25584 (P3_U3409, P3_U3408, P3_U4786);
  and ginst25585 (P3_U3410, P3_U4789, P3_U4790);
  and ginst25586 (P3_U3411, P3_U3410, P3_U4791);
  and ginst25587 (P3_U3412, P3_U4794, P3_U4795);
  and ginst25588 (P3_U3413, P3_U3412, P3_U4796);
  and ginst25589 (P3_U3414, P3_U4799, P3_U4800);
  and ginst25590 (P3_U3415, P3_U3414, P3_U4801);
  and ginst25591 (P3_U3416, P3_U4804, P3_U4805);
  and ginst25592 (P3_U3417, P3_U3416, P3_U4806);
  and ginst25593 (P3_U3418, P3_U4809, P3_U4810);
  and ginst25594 (P3_U3419, P3_U3418, P3_U4811);
  and ginst25595 (P3_U3420, P3_U4814, P3_U4815);
  and ginst25596 (P3_U3421, P3_U3420, P3_U4816);
  and ginst25597 (P3_U3422, P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN, P3_U3129);
  and ginst25598 (P3_U3423, P3_U4312, P3_U4826);
  and ginst25599 (P3_U3424, P3_U4830, P3_U4831);
  and ginst25600 (P3_U3425, P3_U3424, P3_U4832);
  and ginst25601 (P3_U3426, P3_U4835, P3_U4836);
  and ginst25602 (P3_U3427, P3_U3426, P3_U4837);
  and ginst25603 (P3_U3428, P3_U4840, P3_U4841);
  and ginst25604 (P3_U3429, P3_U3428, P3_U4842);
  and ginst25605 (P3_U3430, P3_U4845, P3_U4846);
  and ginst25606 (P3_U3431, P3_U3430, P3_U4847);
  and ginst25607 (P3_U3432, P3_U4850, P3_U4851);
  and ginst25608 (P3_U3433, P3_U3432, P3_U4852);
  and ginst25609 (P3_U3434, P3_U4855, P3_U4856);
  and ginst25610 (P3_U3435, P3_U3434, P3_U4857);
  and ginst25611 (P3_U3436, P3_U4860, P3_U4861);
  and ginst25612 (P3_U3437, P3_U3436, P3_U4862);
  and ginst25613 (P3_U3438, P3_U4865, P3_U4866);
  and ginst25614 (P3_U3439, P3_U3438, P3_U4867);
  and ginst25615 (P3_U3440, P3_U4312, P3_U4878);
  and ginst25616 (P3_U3441, P3_U4882, P3_U4883);
  and ginst25617 (P3_U3442, P3_U3441, P3_U4884);
  and ginst25618 (P3_U3443, P3_U4887, P3_U4888);
  and ginst25619 (P3_U3444, P3_U3443, P3_U4889);
  and ginst25620 (P3_U3445, P3_U4892, P3_U4893);
  and ginst25621 (P3_U3446, P3_U3445, P3_U4894);
  and ginst25622 (P3_U3447, P3_U4897, P3_U4898);
  and ginst25623 (P3_U3448, P3_U3447, P3_U4899);
  and ginst25624 (P3_U3449, P3_U4902, P3_U4903);
  and ginst25625 (P3_U3450, P3_U3449, P3_U4904);
  and ginst25626 (P3_U3451, P3_U4907, P3_U4908);
  and ginst25627 (P3_U3452, P3_U3451, P3_U4909);
  and ginst25628 (P3_U3453, P3_U4912, P3_U4913);
  and ginst25629 (P3_U3454, P3_U3453, P3_U4914);
  and ginst25630 (P3_U3455, P3_U4917, P3_U4918);
  and ginst25631 (P3_U3456, P3_U3455, P3_U4919);
  and ginst25632 (P3_U3457, P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN, P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN);
  and ginst25633 (P3_U3458, P3_U4312, P3_U4930);
  and ginst25634 (P3_U3459, P3_U4934, P3_U4935);
  and ginst25635 (P3_U3460, P3_U3459, P3_U4936);
  and ginst25636 (P3_U3461, P3_U4939, P3_U4940);
  and ginst25637 (P3_U3462, P3_U3461, P3_U4941);
  and ginst25638 (P3_U3463, P3_U4944, P3_U4945);
  and ginst25639 (P3_U3464, P3_U3463, P3_U4946);
  and ginst25640 (P3_U3465, P3_U4949, P3_U4950);
  and ginst25641 (P3_U3466, P3_U3465, P3_U4951);
  and ginst25642 (P3_U3467, P3_U4954, P3_U4955);
  and ginst25643 (P3_U3468, P3_U3467, P3_U4956);
  and ginst25644 (P3_U3469, P3_U4959, P3_U4960);
  and ginst25645 (P3_U3470, P3_U3469, P3_U4961);
  and ginst25646 (P3_U3471, P3_U4964, P3_U4965);
  and ginst25647 (P3_U3472, P3_U3471, P3_U4966);
  and ginst25648 (P3_U3473, P3_U4969, P3_U4970);
  and ginst25649 (P3_U3474, P3_U3473, P3_U4971);
  and ginst25650 (P3_U3475, P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN, P3_U3131);
  and ginst25651 (P3_U3476, P3_U4312, P3_U4982);
  and ginst25652 (P3_U3477, P3_U4986, P3_U4987);
  and ginst25653 (P3_U3478, P3_U3477, P3_U4988);
  and ginst25654 (P3_U3479, P3_U4991, P3_U4992);
  and ginst25655 (P3_U3480, P3_U3479, P3_U4993);
  and ginst25656 (P3_U3481, P3_U4996, P3_U4997);
  and ginst25657 (P3_U3482, P3_U3481, P3_U4998);
  and ginst25658 (P3_U3483, P3_U5001, P3_U5002);
  and ginst25659 (P3_U3484, P3_U3483, P3_U5003);
  and ginst25660 (P3_U3485, P3_U5006, P3_U5007);
  and ginst25661 (P3_U3486, P3_U3485, P3_U5008);
  and ginst25662 (P3_U3487, P3_U5011, P3_U5012);
  and ginst25663 (P3_U3488, P3_U3487, P3_U5013);
  and ginst25664 (P3_U3489, P3_U5016, P3_U5017);
  and ginst25665 (P3_U3490, P3_U3489, P3_U5018);
  and ginst25666 (P3_U3491, P3_U5021, P3_U5022);
  and ginst25667 (P3_U3492, P3_U3491, P3_U5023);
  and ginst25668 (P3_U3493, P3_U4312, P3_U5033);
  and ginst25669 (P3_U3494, P3_U5037, P3_U5038);
  and ginst25670 (P3_U3495, P3_U3494, P3_U5039);
  and ginst25671 (P3_U3496, P3_U5042, P3_U5043);
  and ginst25672 (P3_U3497, P3_U3496, P3_U5044);
  and ginst25673 (P3_U3498, P3_U5047, P3_U5048);
  and ginst25674 (P3_U3499, P3_U3498, P3_U5049);
  and ginst25675 (P3_U3500, P3_U5052, P3_U5053);
  and ginst25676 (P3_U3501, P3_U3500, P3_U5054);
  and ginst25677 (P3_U3502, P3_U5057, P3_U5058);
  and ginst25678 (P3_U3503, P3_U3502, P3_U5059);
  and ginst25679 (P3_U3504, P3_U5062, P3_U5063);
  and ginst25680 (P3_U3505, P3_U3504, P3_U5064);
  and ginst25681 (P3_U3506, P3_U5067, P3_U5068);
  and ginst25682 (P3_U3507, P3_U3506, P3_U5069);
  and ginst25683 (P3_U3508, P3_U5072, P3_U5073);
  and ginst25684 (P3_U3509, P3_U3508, P3_U5074);
  and ginst25685 (P3_U3510, P3_U4312, P3_U5082);
  and ginst25686 (P3_U3511, P3_U5086, P3_U5087);
  and ginst25687 (P3_U3512, P3_U3511, P3_U5088);
  and ginst25688 (P3_U3513, P3_U5091, P3_U5092);
  and ginst25689 (P3_U3514, P3_U3513, P3_U5093);
  and ginst25690 (P3_U3515, P3_U5096, P3_U5097);
  and ginst25691 (P3_U3516, P3_U3515, P3_U5098);
  and ginst25692 (P3_U3517, P3_U5101, P3_U5102);
  and ginst25693 (P3_U3518, P3_U3517, P3_U5103);
  and ginst25694 (P3_U3519, P3_U5106, P3_U5107);
  and ginst25695 (P3_U3520, P3_U3519, P3_U5108);
  and ginst25696 (P3_U3521, P3_U5111, P3_U5112);
  and ginst25697 (P3_U3522, P3_U3521, P3_U5113);
  and ginst25698 (P3_U3523, P3_U5116, P3_U5117);
  and ginst25699 (P3_U3524, P3_U3523, P3_U5118);
  and ginst25700 (P3_U3525, P3_U5121, P3_U5122);
  and ginst25701 (P3_U3526, P3_U3525, P3_U5123);
  and ginst25702 (P3_U3527, P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN, P3_U3133);
  and ginst25703 (P3_U3528, P3_U4312, P3_U5134);
  and ginst25704 (P3_U3529, P3_U5138, P3_U5139);
  and ginst25705 (P3_U3530, P3_U3529, P3_U5140);
  and ginst25706 (P3_U3531, P3_U5143, P3_U5144);
  and ginst25707 (P3_U3532, P3_U3531, P3_U5145);
  and ginst25708 (P3_U3533, P3_U5148, P3_U5149);
  and ginst25709 (P3_U3534, P3_U3533, P3_U5150);
  and ginst25710 (P3_U3535, P3_U5153, P3_U5154);
  and ginst25711 (P3_U3536, P3_U3535, P3_U5155);
  and ginst25712 (P3_U3537, P3_U5158, P3_U5159);
  and ginst25713 (P3_U3538, P3_U3537, P3_U5160);
  and ginst25714 (P3_U3539, P3_U5163, P3_U5164);
  and ginst25715 (P3_U3540, P3_U3539, P3_U5165);
  and ginst25716 (P3_U3541, P3_U5168, P3_U5169);
  and ginst25717 (P3_U3542, P3_U3541, P3_U5170);
  and ginst25718 (P3_U3543, P3_U5173, P3_U5174);
  and ginst25719 (P3_U3544, P3_U3543, P3_U5175);
  and ginst25720 (P3_U3545, P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN, P3_U3133);
  and ginst25721 (P3_U3546, P3_U4312, P3_U5186);
  and ginst25722 (P3_U3547, P3_U5190, P3_U5191);
  and ginst25723 (P3_U3548, P3_U3547, P3_U5192);
  and ginst25724 (P3_U3549, P3_U5195, P3_U5196);
  and ginst25725 (P3_U3550, P3_U3549, P3_U5197);
  and ginst25726 (P3_U3551, P3_U5200, P3_U5201);
  and ginst25727 (P3_U3552, P3_U3551, P3_U5202);
  and ginst25728 (P3_U3553, P3_U5205, P3_U5206);
  and ginst25729 (P3_U3554, P3_U3553, P3_U5207);
  and ginst25730 (P3_U3555, P3_U5210, P3_U5211);
  and ginst25731 (P3_U3556, P3_U3555, P3_U5212);
  and ginst25732 (P3_U3557, P3_U5215, P3_U5216);
  and ginst25733 (P3_U3558, P3_U3557, P3_U5217);
  and ginst25734 (P3_U3559, P3_U5220, P3_U5221);
  and ginst25735 (P3_U3560, P3_U3559, P3_U5222);
  and ginst25736 (P3_U3561, P3_U5225, P3_U5226);
  and ginst25737 (P3_U3562, P3_U3561, P3_U5227);
  nor ginst25738 (P3_U3563, P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN, P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN);
  and ginst25739 (P3_U3564, P3_U4312, P3_U5237);
  and ginst25740 (P3_U3565, P3_U5240, P3_U5241, P3_U5243);
  and ginst25741 (P3_U3566, P3_U3565, P3_U5242);
  and ginst25742 (P3_U3567, P3_U5245, P3_U5246, P3_U5248);
  and ginst25743 (P3_U3568, P3_U3567, P3_U5247);
  and ginst25744 (P3_U3569, P3_U5250, P3_U5251, P3_U5253);
  and ginst25745 (P3_U3570, P3_U3569, P3_U5252);
  and ginst25746 (P3_U3571, P3_U5255, P3_U5256, P3_U5258);
  and ginst25747 (P3_U3572, P3_U3571, P3_U5257);
  and ginst25748 (P3_U3573, P3_U5260, P3_U5261, P3_U5263);
  and ginst25749 (P3_U3574, P3_U3573, P3_U5262);
  and ginst25750 (P3_U3575, P3_U5265, P3_U5266, P3_U5268);
  and ginst25751 (P3_U3576, P3_U3575, P3_U5267);
  and ginst25752 (P3_U3577, P3_U5270, P3_U5271, P3_U5273);
  and ginst25753 (P3_U3578, P3_U3577, P3_U5272);
  and ginst25754 (P3_U3579, P3_U5275, P3_U5276, P3_U5278);
  and ginst25755 (P3_U3580, P3_U3579, P3_U5277);
  nor ginst25756 (P3_U3581, P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN, P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN);
  and ginst25757 (P3_U3582, P3_U4312, P3_U5288);
  and ginst25758 (P3_U3583, P3_U5291, P3_U5292, P3_U5294);
  and ginst25759 (P3_U3584, P3_U3583, P3_U5293);
  and ginst25760 (P3_U3585, P3_U5296, P3_U5297, P3_U5299);
  and ginst25761 (P3_U3586, P3_U3585, P3_U5298);
  and ginst25762 (P3_U3587, P3_U5301, P3_U5302, P3_U5304);
  and ginst25763 (P3_U3588, P3_U3587, P3_U5303);
  and ginst25764 (P3_U3589, P3_U5306, P3_U5307, P3_U5309);
  and ginst25765 (P3_U3590, P3_U3589, P3_U5308);
  and ginst25766 (P3_U3591, P3_U5311, P3_U5312, P3_U5314);
  and ginst25767 (P3_U3592, P3_U3591, P3_U5313);
  and ginst25768 (P3_U3593, P3_U5316, P3_U5317, P3_U5319);
  and ginst25769 (P3_U3594, P3_U3593, P3_U5318);
  and ginst25770 (P3_U3595, P3_U5321, P3_U5322, P3_U5324);
  and ginst25771 (P3_U3596, P3_U3595, P3_U5323);
  and ginst25772 (P3_U3597, P3_U5326, P3_U5327, P3_U5329);
  and ginst25773 (P3_U3598, P3_U3597, P3_U5328);
  and ginst25774 (P3_U3599, P3_U4312, P3_U5339);
  and ginst25775 (P3_U3600, P3_U5342, P3_U5343, P3_U5345);
  and ginst25776 (P3_U3601, P3_U3600, P3_U5344);
  and ginst25777 (P3_U3602, P3_U5347, P3_U5348, P3_U5350);
  and ginst25778 (P3_U3603, P3_U3602, P3_U5349);
  and ginst25779 (P3_U3604, P3_U5352, P3_U5353, P3_U5355);
  and ginst25780 (P3_U3605, P3_U3604, P3_U5354);
  and ginst25781 (P3_U3606, P3_U5357, P3_U5358, P3_U5360);
  and ginst25782 (P3_U3607, P3_U3606, P3_U5359);
  and ginst25783 (P3_U3608, P3_U5362, P3_U5363, P3_U5365);
  and ginst25784 (P3_U3609, P3_U3608, P3_U5364);
  and ginst25785 (P3_U3610, P3_U5367, P3_U5368, P3_U5370);
  and ginst25786 (P3_U3611, P3_U3610, P3_U5369);
  and ginst25787 (P3_U3612, P3_U5372, P3_U5373, P3_U5375);
  and ginst25788 (P3_U3613, P3_U3612, P3_U5374);
  and ginst25789 (P3_U3614, P3_U5377, P3_U5378, P3_U5380);
  and ginst25790 (P3_U3615, P3_U3614, P3_U5379);
  nor ginst25791 (P3_U3616, P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN, P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN);
  and ginst25792 (P3_U3617, P3_U4312, P3_U5390);
  and ginst25793 (P3_U3618, P3_U5393, P3_U5394, P3_U5396);
  and ginst25794 (P3_U3619, P3_U3618, P3_U5395);
  and ginst25795 (P3_U3620, P3_U5398, P3_U5399, P3_U5401);
  and ginst25796 (P3_U3621, P3_U3620, P3_U5400);
  and ginst25797 (P3_U3622, P3_U5403, P3_U5404, P3_U5406);
  and ginst25798 (P3_U3623, P3_U3622, P3_U5405);
  and ginst25799 (P3_U3624, P3_U5408, P3_U5409, P3_U5411);
  and ginst25800 (P3_U3625, P3_U3624, P3_U5410);
  and ginst25801 (P3_U3626, P3_U5413, P3_U5414, P3_U5416);
  and ginst25802 (P3_U3627, P3_U3626, P3_U5415);
  and ginst25803 (P3_U3628, P3_U5418, P3_U5419, P3_U5421);
  and ginst25804 (P3_U3629, P3_U3628, P3_U5420);
  and ginst25805 (P3_U3630, P3_U5423, P3_U5424, P3_U5426);
  and ginst25806 (P3_U3631, P3_U3630, P3_U5425);
  and ginst25807 (P3_U3632, P3_U5428, P3_U5429, P3_U5431);
  and ginst25808 (P3_U3633, P3_U3632, P3_U5430);
  nor ginst25809 (P3_U3634, P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN, P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN);
  and ginst25810 (P3_U3635, P3_U4312, P3_U5440);
  and ginst25811 (P3_U3636, P3_U5443, P3_U5444, P3_U5446);
  and ginst25812 (P3_U3637, P3_U3636, P3_U5445);
  and ginst25813 (P3_U3638, P3_U5448, P3_U5449, P3_U5451);
  and ginst25814 (P3_U3639, P3_U3638, P3_U5450);
  and ginst25815 (P3_U3640, P3_U5453, P3_U5454, P3_U5456);
  and ginst25816 (P3_U3641, P3_U3640, P3_U5455);
  and ginst25817 (P3_U3642, P3_U5458, P3_U5459, P3_U5461);
  and ginst25818 (P3_U3643, P3_U3642, P3_U5460);
  and ginst25819 (P3_U3644, P3_U5463, P3_U5464, P3_U5466);
  and ginst25820 (P3_U3645, P3_U3644, P3_U5465);
  and ginst25821 (P3_U3646, P3_U5468, P3_U5469, P3_U5471);
  and ginst25822 (P3_U3647, P3_U3646, P3_U5470);
  and ginst25823 (P3_U3648, P3_U5473, P3_U5474, P3_U5476);
  and ginst25824 (P3_U3649, P3_U3648, P3_U5475);
  and ginst25825 (P3_U3650, P3_U5478, P3_U5479, P3_U5481);
  and ginst25826 (P3_U3651, P3_U3650, P3_U5480);
  and ginst25827 (P3_U3652, P3_ADD_495_U8, P3_U4340);
  and ginst25828 (P3_U3653, P3_STATE2_REG_0__SCAN_IN, P3_FLUSH_REG_SCAN_IN);
  and ginst25829 (P3_U3654, P3_U3104, P3_U4522);
  and ginst25830 (P3_U3655, P3_U3107, P3_U3118);
  and ginst25831 (P3_U3656, P3_U4333, P3_U5495);
  and ginst25832 (P3_U3657, P3_U3656, P3_U5494);
  and ginst25833 (P3_U3658, P3_U4330, P3_U5498);
  and ginst25834 (P3_U3659, P3_U5501, P3_U5502);
  and ginst25835 (P3_U3660, P3_U4539, P3_U4556);
  and ginst25836 (P3_U3661, P3_U2461, P3_U4297);
  and ginst25837 (P3_U3662, P3_U3101, P3_U4590);
  and ginst25838 (P3_U3663, P3_U3101, P3_U4556);
  and ginst25839 (P3_U3664, P3_U4324, P3_U4573);
  and ginst25840 (P3_U3665, P3_U5508, P3_U5510, P3_U5511);
  and ginst25841 (P3_U3666, P3_U4339, P3_U5519, P3_U5520);
  and ginst25842 (P3_U3667, P3_U3666, P3_U5521, P3_U7977, P3_U7978);
  and ginst25843 (P3_U3668, P3_U2517, P3_U3242, P3_U5528);
  and ginst25844 (P3_U3669, P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P3_U4470);
  and ginst25845 (P3_U3670, P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P3_U3093);
  and ginst25846 (P3_U3671, P3_U3116, P3_U3117, P3_U3119);
  and ginst25847 (P3_U3672, P3_U3244, P3_U3245, P3_U3671);
  and ginst25848 (P3_U3673, P3_U2456, P3_U4505);
  and ginst25849 (P3_U3674, P3_U5532, P3_U5533);
  and ginst25850 (P3_U3675, P3_U5536, P3_U5538);
  and ginst25851 (P3_U3676, P3_U3675, P3_U3677, P3_U5539);
  and ginst25852 (P3_U3677, P3_U5540, P3_U5541);
  and ginst25853 (P3_U3678, P3_U5550, P3_U5552);
  and ginst25854 (P3_U3679, P3_U3678, P3_U5551);
  and ginst25855 (P3_U3680, P3_U5554, P3_U5555);
  and ginst25856 (P3_U3681, P3_U3682, P3_U5562);
  and ginst25857 (P3_U3682, P3_U5564, P3_U5565);
  and ginst25858 (P3_U3683, P3_U5567, P3_U5568);
  and ginst25859 (P3_U3684, P3_U5574, P3_U5576);
  and ginst25860 (P3_U3685, P3_U5587, P3_U5588);
  and ginst25861 (P3_U3686, P3_U5592, P3_U5594);
  and ginst25862 (P3_U3687, P3_U4333, P3_U5625, P3_U5626);
  and ginst25863 (P3_U3688, P3_U2456, P3_U4296);
  and ginst25864 (P3_U3689, P3_U2456, P3_U4323);
  and ginst25865 (P3_U3690, P3_U4556, P3_U4608);
  and ginst25866 (P3_U3691, P3_U2456, P3_U4590);
  and ginst25867 (P3_U3692, P3_U5635, P3_U5636);
  and ginst25868 (P3_U3693, P3_U3694, P3_U5632, P3_U5633, P3_U5637, P3_U5638);
  and ginst25869 (P3_U3694, P3_U3695, P3_U5641);
  and ginst25870 (P3_U3695, P3_U5639, P3_U5640);
  and ginst25871 (P3_U3696, P3_U5642, P3_U5643, P3_U5644, P3_U5645, P3_U5646);
  and ginst25872 (P3_U3697, P3_U5647, P3_U5648, P3_U5649, P3_U5650, P3_U5651);
  and ginst25873 (P3_U3698, P3_U3696, P3_U3697);
  and ginst25874 (P3_U3699, P3_U5659, P3_U5660);
  and ginst25875 (P3_U3700, P3_U3701, P3_U5657, P3_U5661, P3_U5662);
  and ginst25876 (P3_U3701, P3_U3702, P3_U5665);
  and ginst25877 (P3_U3702, P3_U5663, P3_U5664);
  and ginst25878 (P3_U3703, P3_U5666, P3_U5667, P3_U5668, P3_U5669, P3_U5670);
  and ginst25879 (P3_U3704, P3_U5671, P3_U5672, P3_U5673, P3_U5674);
  and ginst25880 (P3_U3705, P3_U3703, P3_U3704, P3_U5675);
  and ginst25881 (P3_U3706, P3_U3707, P3_U5681);
  and ginst25882 (P3_U3707, P3_U5683, P3_U5684);
  and ginst25883 (P3_U3708, P3_U3709, P3_U5689);
  and ginst25884 (P3_U3709, P3_U5687, P3_U5688);
  and ginst25885 (P3_U3710, P3_U3708, P3_U5685, P3_U5686);
  and ginst25886 (P3_U3711, P3_U5690, P3_U5691, P3_U5692, P3_U5693, P3_U5694);
  and ginst25887 (P3_U3712, P3_U5695, P3_U5696, P3_U5697, P3_U5698);
  and ginst25888 (P3_U3713, P3_U3711, P3_U3712, P3_U5699);
  and ginst25889 (P3_U3714, P3_U5704, P3_U5705);
  and ginst25890 (P3_U3715, P3_U5707, P3_U5708);
  and ginst25891 (P3_U3716, P3_U3717, P3_U5713);
  and ginst25892 (P3_U3717, P3_U5711, P3_U5712);
  and ginst25893 (P3_U3718, P3_U3716, P3_U5709, P3_U5710);
  and ginst25894 (P3_U3719, P3_U5714, P3_U5715, P3_U5716, P3_U5717, P3_U5718);
  and ginst25895 (P3_U3720, P3_U5719, P3_U5720, P3_U5721, P3_U5722);
  and ginst25896 (P3_U3721, P3_U3719, P3_U3720, P3_U5723);
  and ginst25897 (P3_U3722, P3_U3723, P3_U5729);
  and ginst25898 (P3_U3723, P3_U5731, P3_U5732);
  and ginst25899 (P3_U3724, P3_U3725, P3_U5737);
  and ginst25900 (P3_U3725, P3_U5735, P3_U5736);
  and ginst25901 (P3_U3726, P3_U3724, P3_U5733, P3_U5734);
  and ginst25902 (P3_U3727, P3_U5738, P3_U5739, P3_U5740, P3_U5741, P3_U5742);
  and ginst25903 (P3_U3728, P3_U5743, P3_U5744, P3_U5745, P3_U5746);
  and ginst25904 (P3_U3729, P3_U3727, P3_U3728, P3_U5747);
  and ginst25905 (P3_U3730, P3_U3731, P3_U5752);
  and ginst25906 (P3_U3731, P3_U5755, P3_U5756);
  and ginst25907 (P3_U3732, P3_U3733, P3_U5761);
  and ginst25908 (P3_U3733, P3_U5759, P3_U5760);
  and ginst25909 (P3_U3734, P3_U3732, P3_U5757, P3_U5758);
  and ginst25910 (P3_U3735, P3_U5762, P3_U5763, P3_U5764, P3_U5765, P3_U5766);
  and ginst25911 (P3_U3736, P3_U5767, P3_U5768, P3_U5769, P3_U5770);
  and ginst25912 (P3_U3737, P3_U3735, P3_U3736, P3_U5771);
  and ginst25913 (P3_U3738, P3_U3739, P3_U5776);
  and ginst25914 (P3_U3739, P3_U5779, P3_U5780);
  and ginst25915 (P3_U3740, P3_U3741, P3_U5785);
  and ginst25916 (P3_U3741, P3_U5783, P3_U5784);
  and ginst25917 (P3_U3742, P3_U3740, P3_U5781, P3_U5782);
  and ginst25918 (P3_U3743, P3_U5786, P3_U5787, P3_U5788, P3_U5789, P3_U5790);
  and ginst25919 (P3_U3744, P3_U5791, P3_U5792, P3_U5793, P3_U5794);
  and ginst25920 (P3_U3745, P3_U3743, P3_U3744, P3_U5795);
  and ginst25921 (P3_U3746, P3_U3747, P3_U5800);
  and ginst25922 (P3_U3747, P3_U5803, P3_U5804);
  and ginst25923 (P3_U3748, P3_U3749, P3_U5809);
  and ginst25924 (P3_U3749, P3_U5807, P3_U5808);
  and ginst25925 (P3_U3750, P3_U3748, P3_U5805, P3_U5806);
  and ginst25926 (P3_U3751, P3_U5810, P3_U5811, P3_U5812, P3_U5813, P3_U5814);
  and ginst25927 (P3_U3752, P3_U5815, P3_U5816, P3_U5817, P3_U5818);
  and ginst25928 (P3_U3753, P3_U3751, P3_U3752, P3_U5819);
  and ginst25929 (P3_U3754, P3_U3755, P3_U5824);
  and ginst25930 (P3_U3755, P3_U5827, P3_U5828);
  and ginst25931 (P3_U3756, P3_U5831, P3_U5832, P3_U5833);
  and ginst25932 (P3_U3757, P3_U3756, P3_U5829, P3_U5830);
  and ginst25933 (P3_U3758, P3_U5834, P3_U5835, P3_U5836, P3_U5837, P3_U5838);
  and ginst25934 (P3_U3759, P3_U5839, P3_U5840, P3_U5841, P3_U5842);
  and ginst25935 (P3_U3760, P3_U3758, P3_U3759, P3_U5843);
  and ginst25936 (P3_U3761, P3_U3762, P3_U5848);
  and ginst25937 (P3_U3762, P3_U5851, P3_U5852);
  and ginst25938 (P3_U3763, P3_U5856, P3_U5857);
  and ginst25939 (P3_U3764, P3_U3763, P3_U5853, P3_U5854, P3_U5855);
  and ginst25940 (P3_U3765, P3_U5858, P3_U5859, P3_U5860, P3_U5861, P3_U5862);
  and ginst25941 (P3_U3766, P3_U5863, P3_U5864, P3_U5865, P3_U5866);
  and ginst25942 (P3_U3767, P3_U3765, P3_U3766, P3_U5867);
  and ginst25943 (P3_U3768, P3_U3769, P3_U5873);
  and ginst25944 (P3_U3769, P3_U5875, P3_U5876);
  and ginst25945 (P3_U3770, P3_U5880, P3_U5881);
  and ginst25946 (P3_U3771, P3_U3770, P3_U5877, P3_U5878, P3_U5879);
  and ginst25947 (P3_U3772, P3_U5882, P3_U5883, P3_U5884, P3_U5885, P3_U5886);
  and ginst25948 (P3_U3773, P3_U5887, P3_U5888, P3_U5889, P3_U5890);
  and ginst25949 (P3_U3774, P3_U3772, P3_U3773, P3_U5891);
  and ginst25950 (P3_U3775, P3_U3776, P3_U5897);
  and ginst25951 (P3_U3776, P3_U5899, P3_U5900);
  and ginst25952 (P3_U3777, P3_U5904, P3_U5905);
  and ginst25953 (P3_U3778, P3_U3777, P3_U5901, P3_U5902, P3_U5903);
  and ginst25954 (P3_U3779, P3_U5906, P3_U5907, P3_U5908, P3_U5909, P3_U5910);
  and ginst25955 (P3_U3780, P3_U5911, P3_U5912, P3_U5913, P3_U5914);
  and ginst25956 (P3_U3781, P3_U3779, P3_U3780, P3_U5915);
  and ginst25957 (P3_U3782, P3_U3783, P3_U5920);
  and ginst25958 (P3_U3783, P3_U5923, P3_U5924);
  and ginst25959 (P3_U3784, P3_U5928, P3_U5929);
  and ginst25960 (P3_U3785, P3_U3784, P3_U5925, P3_U5926, P3_U5927);
  and ginst25961 (P3_U3786, P3_U5930, P3_U5931, P3_U5932, P3_U5933, P3_U5934);
  and ginst25962 (P3_U3787, P3_U5935, P3_U5936, P3_U5937, P3_U5938);
  and ginst25963 (P3_U3788, P3_U3786, P3_U3787, P3_U5939);
  and ginst25964 (P3_U3789, P3_U3790, P3_U5944);
  and ginst25965 (P3_U3790, P3_U5947, P3_U5948);
  and ginst25966 (P3_U3791, P3_U5952, P3_U5953);
  and ginst25967 (P3_U3792, P3_U3791, P3_U5949, P3_U5950, P3_U5951);
  and ginst25968 (P3_U3793, P3_U5954, P3_U5955, P3_U5956, P3_U5957, P3_U5958);
  and ginst25969 (P3_U3794, P3_U5959, P3_U5960, P3_U5961, P3_U5962);
  and ginst25970 (P3_U3795, P3_U3793, P3_U3794, P3_U5963);
  and ginst25971 (P3_U3796, P3_U5971, P3_U5972);
  and ginst25972 (P3_U3797, P3_U5976, P3_U5977);
  and ginst25973 (P3_U3798, P3_U3797, P3_U5973, P3_U5974, P3_U5975);
  and ginst25974 (P3_U3799, P3_U3796, P3_U3798, P3_U5968, P3_U5969, P3_U5970);
  and ginst25975 (P3_U3800, P3_U5978, P3_U5979, P3_U5980, P3_U5981, P3_U5982);
  and ginst25976 (P3_U3801, P3_U5983, P3_U5984, P3_U5985, P3_U5986);
  and ginst25977 (P3_U3802, P3_U3800, P3_U3801, P3_U5987);
  and ginst25978 (P3_U3803, P3_U5989, P3_U5991);
  and ginst25979 (P3_U3804, P3_U5995, P3_U5996);
  and ginst25980 (P3_U3805, P3_U6000, P3_U6001);
  and ginst25981 (P3_U3806, P3_U3805, P3_U5997, P3_U5998, P3_U5999);
  and ginst25982 (P3_U3807, P3_U3804, P3_U3806, P3_U5992, P3_U5993, P3_U5994);
  and ginst25983 (P3_U3808, P3_U6002, P3_U6003, P3_U6004, P3_U6005, P3_U6006);
  and ginst25984 (P3_U3809, P3_U6007, P3_U6008, P3_U6009, P3_U6010);
  and ginst25985 (P3_U3810, P3_U3808, P3_U3809, P3_U6011);
  and ginst25986 (P3_U3811, P3_U6013, P3_U6015);
  and ginst25987 (P3_U3812, P3_U3813, P3_U6017);
  and ginst25988 (P3_U3813, P3_U6019, P3_U6020);
  and ginst25989 (P3_U3814, P3_U6024, P3_U6025);
  and ginst25990 (P3_U3815, P3_U3814, P3_U6021, P3_U6022, P3_U6023);
  and ginst25991 (P3_U3816, P3_U6026, P3_U6027, P3_U6028, P3_U6029, P3_U6030);
  and ginst25992 (P3_U3817, P3_U6031, P3_U6032, P3_U6033, P3_U6034);
  and ginst25993 (P3_U3818, P3_U3816, P3_U3817, P3_U6035);
  and ginst25994 (P3_U3819, P3_U6043, P3_U6044);
  and ginst25995 (P3_U3820, P3_U3821, P3_U6041, P3_U6045, P3_U6046, P3_U6047);
  and ginst25996 (P3_U3821, P3_U6048, P3_U6049);
  and ginst25997 (P3_U3822, P3_U6050, P3_U6051, P3_U6052, P3_U6053, P3_U6054);
  and ginst25998 (P3_U3823, P3_U6055, P3_U6056, P3_U6057, P3_U6058);
  and ginst25999 (P3_U3824, P3_U3822, P3_U3823, P3_U6059);
  and ginst26000 (P3_U3825, P3_U3826, P3_U6065);
  and ginst26001 (P3_U3826, P3_U6067, P3_U6068);
  and ginst26002 (P3_U3827, P3_U6072, P3_U6073);
  and ginst26003 (P3_U3828, P3_U3827, P3_U6069, P3_U6070, P3_U6071);
  and ginst26004 (P3_U3829, P3_U6074, P3_U6075, P3_U6076, P3_U6077, P3_U6078);
  and ginst26005 (P3_U3830, P3_U6079, P3_U6080, P3_U6081, P3_U6082);
  and ginst26006 (P3_U3831, P3_U3829, P3_U3830, P3_U6083);
  and ginst26007 (P3_U3832, P3_U6091, P3_U6092);
  and ginst26008 (P3_U3833, P3_U3834, P3_U6089, P3_U6093, P3_U6094, P3_U6095);
  and ginst26009 (P3_U3834, P3_U6096, P3_U6097);
  and ginst26010 (P3_U3835, P3_U6098, P3_U6099, P3_U6100, P3_U6101, P3_U6102);
  and ginst26011 (P3_U3836, P3_U6103, P3_U6104, P3_U6105, P3_U6106);
  and ginst26012 (P3_U3837, P3_U3835, P3_U3836, P3_U6107);
  and ginst26013 (P3_U3838, P3_U6115, P3_U6116);
  and ginst26014 (P3_U3839, P3_U6120, P3_U6121);
  and ginst26015 (P3_U3840, P3_U3839, P3_U6117, P3_U6118, P3_U6119);
  and ginst26016 (P3_U3841, P3_U3838, P3_U3840, P3_U3844, P3_U6112, P3_U6114);
  and ginst26017 (P3_U3842, P3_U6122, P3_U6123, P3_U6124, P3_U6125, P3_U6126);
  and ginst26018 (P3_U3843, P3_U6127, P3_U6128, P3_U6129, P3_U6130);
  and ginst26019 (P3_U3844, P3_U3842, P3_U3843, P3_U6131);
  and ginst26020 (P3_U3845, P3_U6133, P3_U6135);
  and ginst26021 (P3_U3846, P3_U6139, P3_U6140);
  and ginst26022 (P3_U3847, P3_U6144, P3_U6145);
  and ginst26023 (P3_U3848, P3_U3847, P3_U6141, P3_U6142, P3_U6143);
  and ginst26024 (P3_U3849, P3_U3846, P3_U3848, P3_U3852, P3_U6136, P3_U6138);
  and ginst26025 (P3_U3850, P3_U6146, P3_U6147, P3_U6148, P3_U6149, P3_U6150);
  and ginst26026 (P3_U3851, P3_U6151, P3_U6152, P3_U6153, P3_U6154);
  and ginst26027 (P3_U3852, P3_U3850, P3_U3851, P3_U6155);
  and ginst26028 (P3_U3853, P3_U6157, P3_U6159);
  and ginst26029 (P3_U3854, P3_U6163, P3_U6164);
  and ginst26030 (P3_U3855, P3_U6168, P3_U6169);
  and ginst26031 (P3_U3856, P3_U3855, P3_U6165, P3_U6166, P3_U6167);
  and ginst26032 (P3_U3857, P3_U3854, P3_U3856, P3_U6160, P3_U6161, P3_U6162);
  and ginst26033 (P3_U3858, P3_U6170, P3_U6171, P3_U6172);
  and ginst26034 (P3_U3859, P3_U6173, P3_U6174);
  and ginst26035 (P3_U3860, P3_U6175, P3_U6176, P3_U6177);
  and ginst26036 (P3_U3861, P3_U6178, P3_U6179);
  and ginst26037 (P3_U3862, P3_U3858, P3_U3859, P3_U3860, P3_U3861);
  and ginst26038 (P3_U3863, P3_U6181, P3_U6183);
  and ginst26039 (P3_U3864, P3_U6187, P3_U6188);
  and ginst26040 (P3_U3865, P3_U6192, P3_U6193);
  and ginst26041 (P3_U3866, P3_U3865, P3_U6189, P3_U6190, P3_U6191);
  and ginst26042 (P3_U3867, P3_U3864, P3_U3866, P3_U6184, P3_U6185, P3_U6186);
  and ginst26043 (P3_U3868, P3_U6194, P3_U6195, P3_U6196);
  and ginst26044 (P3_U3869, P3_U6197, P3_U6198);
  and ginst26045 (P3_U3870, P3_U6199, P3_U6200, P3_U6201);
  and ginst26046 (P3_U3871, P3_U6202, P3_U6203);
  and ginst26047 (P3_U3872, P3_U3868, P3_U3869, P3_U3870, P3_U3871);
  and ginst26048 (P3_U3873, P3_U6205, P3_U6207);
  and ginst26049 (P3_U3874, P3_U6211, P3_U6212);
  and ginst26050 (P3_U3875, P3_U6216, P3_U6217);
  and ginst26051 (P3_U3876, P3_U3875, P3_U6213, P3_U6214, P3_U6215);
  and ginst26052 (P3_U3877, P3_U3874, P3_U3876, P3_U6208, P3_U6209, P3_U6210);
  and ginst26053 (P3_U3878, P3_U6218, P3_U6219, P3_U6220);
  and ginst26054 (P3_U3879, P3_U6221, P3_U6222);
  and ginst26055 (P3_U3880, P3_U6223, P3_U6224, P3_U6225);
  and ginst26056 (P3_U3881, P3_U6226, P3_U6227);
  and ginst26057 (P3_U3882, P3_U3878, P3_U3879, P3_U3880, P3_U3881);
  and ginst26058 (P3_U3883, P3_U6229, P3_U6231);
  and ginst26059 (P3_U3884, P3_U6235, P3_U6236);
  and ginst26060 (P3_U3885, P3_U6240, P3_U6241);
  and ginst26061 (P3_U3886, P3_U3885, P3_U6237, P3_U6238, P3_U6239);
  and ginst26062 (P3_U3887, P3_U3884, P3_U3886, P3_U6232, P3_U6233, P3_U6234);
  and ginst26063 (P3_U3888, P3_U6242, P3_U6243, P3_U6244);
  and ginst26064 (P3_U3889, P3_U6245, P3_U6246);
  and ginst26065 (P3_U3890, P3_U6247, P3_U6248, P3_U6249);
  and ginst26066 (P3_U3891, P3_U6250, P3_U6251);
  and ginst26067 (P3_U3892, P3_U3888, P3_U3889, P3_U3890, P3_U3891);
  and ginst26068 (P3_U3893, P3_U6253, P3_U6255);
  and ginst26069 (P3_U3894, P3_U6256, P3_U6257);
  and ginst26070 (P3_U3895, P3_U6259, P3_U6260);
  and ginst26071 (P3_U3896, P3_U6264, P3_U6265);
  and ginst26072 (P3_U3897, P3_U3896, P3_U6261, P3_U6262, P3_U6263);
  and ginst26073 (P3_U3898, P3_U6266, P3_U6267, P3_U6268);
  and ginst26074 (P3_U3899, P3_U6269, P3_U6270);
  and ginst26075 (P3_U3900, P3_U6271, P3_U6272, P3_U6273);
  and ginst26076 (P3_U3901, P3_U6274, P3_U6275);
  and ginst26077 (P3_U3902, P3_U3898, P3_U3899, P3_U3900, P3_U3901);
  and ginst26078 (P3_U3903, P3_U6280, P3_U6281);
  and ginst26079 (P3_U3904, P3_U6283, P3_U6284);
  and ginst26080 (P3_U3905, P3_U6288, P3_U6289);
  and ginst26081 (P3_U3906, P3_U3905, P3_U6285, P3_U6286, P3_U6287);
  and ginst26082 (P3_U3907, P3_U6290, P3_U6291, P3_U6292);
  and ginst26083 (P3_U3908, P3_U6293, P3_U6294);
  and ginst26084 (P3_U3909, P3_U6295, P3_U6296, P3_U6297);
  and ginst26085 (P3_U3910, P3_U6298, P3_U6299);
  and ginst26086 (P3_U3911, P3_U3907, P3_U3908, P3_U3909, P3_U3910);
  and ginst26087 (P3_U3912, P3_U6304, P3_U6305);
  and ginst26088 (P3_U3913, P3_U6307, P3_U6308);
  and ginst26089 (P3_U3914, P3_U6312, P3_U6313);
  and ginst26090 (P3_U3915, P3_U3914, P3_U6309, P3_U6310, P3_U6311);
  and ginst26091 (P3_U3916, P3_U6314, P3_U6315, P3_U6316);
  and ginst26092 (P3_U3917, P3_U6317, P3_U6318);
  and ginst26093 (P3_U3918, P3_U6319, P3_U6320, P3_U6321);
  and ginst26094 (P3_U3919, P3_U6322, P3_U6323);
  and ginst26095 (P3_U3920, P3_U3916, P3_U3917, P3_U3918, P3_U3919);
  and ginst26096 (P3_U3921, P3_U6328, P3_U6329);
  and ginst26097 (P3_U3922, P3_U6331, P3_U6332);
  and ginst26098 (P3_U3923, P3_U6336, P3_U6337);
  and ginst26099 (P3_U3924, P3_U3923, P3_U6333, P3_U6334, P3_U6335);
  and ginst26100 (P3_U3925, P3_U6338, P3_U6339, P3_U6340);
  and ginst26101 (P3_U3926, P3_U6341, P3_U6342);
  and ginst26102 (P3_U3927, P3_U6343, P3_U6344, P3_U6345);
  and ginst26103 (P3_U3928, P3_U6346, P3_U6347);
  and ginst26104 (P3_U3929, P3_U3925, P3_U3926, P3_U3927, P3_U3928);
  and ginst26105 (P3_U3930, P3_U6352, P3_U6353);
  and ginst26106 (P3_U3931, P3_U6355, P3_U6356);
  and ginst26107 (P3_U3932, P3_U6360, P3_U6361);
  and ginst26108 (P3_U3933, P3_U3932, P3_U6357, P3_U6358, P3_U6359);
  and ginst26109 (P3_U3934, P3_U6362, P3_U6363, P3_U6364);
  and ginst26110 (P3_U3935, P3_U6365, P3_U6366);
  and ginst26111 (P3_U3936, P3_U6367, P3_U6368, P3_U6369);
  and ginst26112 (P3_U3937, P3_U6370, P3_U6371);
  and ginst26113 (P3_U3938, P3_U3934, P3_U3935, P3_U3936, P3_U3937);
  and ginst26114 (P3_U3939, P3_U3247, P3_U6398);
  and ginst26115 (P3_U3940, P3_U6376, P3_U6377);
  and ginst26116 (P3_U3941, P3_U6379, P3_U6380);
  and ginst26117 (P3_U3942, P3_U3941, P3_U6381);
  and ginst26118 (P3_U3943, P3_U6384, P3_U6385, P3_U6386);
  and ginst26119 (P3_U3944, P3_U3943, P3_U6382, P3_U6383);
  and ginst26120 (P3_U3945, P3_U3940, P3_U3942, P3_U3944, P3_U6378);
  and ginst26121 (P3_U3946, P3_U6387, P3_U6388, P3_U6389);
  and ginst26122 (P3_U3947, P3_U6390, P3_U6391);
  and ginst26123 (P3_U3948, P3_U3946, P3_U3947, P3_U6392);
  and ginst26124 (P3_U3949, P3_U6393, P3_U6394);
  and ginst26125 (P3_U3950, P3_U3948, P3_U3949, P3_U6395, P3_U6397, P3_U6398);
  and ginst26126 (P3_U3951, P3_STATE2_REG_0__SCAN_IN, P3_U3104);
  and ginst26127 (P3_U3952, P3_STATE2_REG_2__SCAN_IN, P3_U3121);
  and ginst26128 (P3_U3953, P3_STATE2_REG_0__SCAN_IN, P3_U4505);
  and ginst26129 (P3_U3954, P3_U6409, P3_U6410, P3_U6411, P3_U6412);
  and ginst26130 (P3_U3955, P3_U6417, P3_U6418, P3_U6419, P3_U6420);
  and ginst26131 (P3_U3956, P3_U6425, P3_U6426, P3_U6427, P3_U6428);
  and ginst26132 (P3_U3957, P3_U6433, P3_U6434, P3_U6435, P3_U6436);
  and ginst26133 (P3_U3958, P3_U6441, P3_U6442, P3_U6443, P3_U6444);
  and ginst26134 (P3_U3959, P3_U6449, P3_U6450, P3_U6451, P3_U6452);
  and ginst26135 (P3_U3960, P3_U6457, P3_U6458, P3_U6459, P3_U6460);
  and ginst26136 (P3_U3961, P3_U6465, P3_U6466, P3_U6467, P3_U6468);
  and ginst26137 (P3_U3962, P3_U6473, P3_U6474, P3_U6475, P3_U6476);
  and ginst26138 (P3_U3963, P3_U6481, P3_U6482, P3_U6483, P3_U6484);
  and ginst26139 (P3_U3964, P3_U6489, P3_U6490, P3_U6491, P3_U6492);
  and ginst26140 (P3_U3965, P3_U6497, P3_U6498, P3_U6499, P3_U6500);
  and ginst26141 (P3_U3966, P3_U6505, P3_U6506, P3_U6507, P3_U6508);
  and ginst26142 (P3_U3967, P3_U6513, P3_U6514, P3_U6515, P3_U6516);
  and ginst26143 (P3_U3968, P3_U6521, P3_U6522, P3_U6523, P3_U6524);
  and ginst26144 (P3_U3969, P3_U6529, P3_U6530, P3_U6531, P3_U6532);
  and ginst26145 (P3_U3970, P3_U6537, P3_U6538, P3_U6539, P3_U6540);
  and ginst26146 (P3_U3971, P3_U6545, P3_U6546, P3_U6547, P3_U6548);
  and ginst26147 (P3_U3972, P3_U6553, P3_U6554, P3_U6555, P3_U6556);
  and ginst26148 (P3_U3973, P3_U6561, P3_U6562, P3_U6563, P3_U6564);
  and ginst26149 (P3_U3974, P3_U6569, P3_U6570, P3_U6571, P3_U6572);
  and ginst26150 (P3_U3975, P3_U6577, P3_U6578, P3_U6579, P3_U6580);
  and ginst26151 (P3_U3976, P3_U6585, P3_U6586, P3_U6587, P3_U6588);
  and ginst26152 (P3_U3977, P3_U6593, P3_U6594, P3_U6595, P3_U6596);
  and ginst26153 (P3_U3978, P3_U6601, P3_U6602, P3_U6603, P3_U6604);
  and ginst26154 (P3_U3979, P3_U6609, P3_U6610, P3_U6611, P3_U6612);
  and ginst26155 (P3_U3980, P3_U6617, P3_U6618, P3_U6619, P3_U6620);
  and ginst26156 (P3_U3981, P3_U6625, P3_U6626, P3_U6627, P3_U6628);
  and ginst26157 (P3_U3982, P3_U6633, P3_U6634, P3_U6635, P3_U6636);
  and ginst26158 (P3_U3983, P3_U6641, P3_U6642, P3_U6643, P3_U6644);
  and ginst26159 (P3_U3984, P3_U6649, P3_U6650, P3_U6651, P3_U6652);
  and ginst26160 (P3_U3985, P3_U6657, P3_U6658, P3_U6659, P3_U6660);
  and ginst26161 (P3_U3986, P3_U2390, P3_U4293);
  and ginst26162 (P3_U3987, P3_U6809, P3_U6810);
  and ginst26163 (P3_U3988, P3_U6812, P3_U6813);
  and ginst26164 (P3_U3989, P3_U6815, P3_U6816);
  and ginst26165 (P3_U3990, P3_U6818, P3_U6819);
  and ginst26166 (P3_U3991, P3_U6821, P3_U6822);
  and ginst26167 (P3_U3992, P3_U6824, P3_U6825);
  and ginst26168 (P3_U3993, P3_U6827, P3_U6828);
  and ginst26169 (P3_U3994, P3_U6830, P3_U6831);
  and ginst26170 (P3_U3995, P3_U6833, P3_U6834);
  and ginst26171 (P3_U3996, P3_U6836, P3_U6837);
  and ginst26172 (P3_U3997, P3_U6839, P3_U6840);
  and ginst26173 (P3_U3998, P3_U6842, P3_U6843);
  and ginst26174 (P3_U3999, P3_U6845, P3_U6846);
  and ginst26175 (P3_U4000, P3_U6848, P3_U6849);
  and ginst26176 (P3_U4001, P3_U6851, P3_U6852);
  and ginst26177 (P3_U4002, P3_U6856, P3_U6857);
  and ginst26178 (P3_U4003, P3_U6860, P3_U6861);
  and ginst26179 (P3_U4004, P3_U6864, P3_U6865);
  and ginst26180 (P3_U4005, P3_U6868, P3_U6869);
  and ginst26181 (P3_U4006, P3_U6872, P3_U6873);
  and ginst26182 (P3_U4007, P3_U6876, P3_U6877);
  and ginst26183 (P3_U4008, P3_U6880, P3_U6881);
  and ginst26184 (P3_U4009, P3_U6884, P3_U6885);
  and ginst26185 (P3_U4010, P3_U6888, P3_U6889);
  and ginst26186 (P3_U4011, P3_U6892, P3_U6893);
  and ginst26187 (P3_U4012, P3_U6896, P3_U6897);
  and ginst26188 (P3_U4013, P3_U6900, P3_U6901);
  and ginst26189 (P3_U4014, P3_U6904, P3_U6905);
  and ginst26190 (P3_U4015, P3_U6907, P3_U6909);
  and ginst26191 (P3_U4016, P3_U6911, P3_U6913);
  and ginst26192 (P3_U4017, P3_U6915, P3_U6917);
  and ginst26193 (P3_U4018, P3_U6920, P3_U6922);
  and ginst26194 (P3_U4019, P3_U6925, P3_U6927);
  and ginst26195 (P3_U4020, P3_U6930, P3_U6932);
  and ginst26196 (P3_U4021, P3_U6935, P3_U6937);
  and ginst26197 (P3_U4022, P3_U6940, P3_U6942);
  and ginst26198 (P3_U4023, P3_U6945, P3_U6947);
  and ginst26199 (P3_U4024, P3_U6950, P3_U6952);
  and ginst26200 (P3_U4025, P3_U6955, P3_U6957);
  and ginst26201 (P3_U4026, P3_U6960, P3_U6962);
  and ginst26202 (P3_U4027, P3_U6965, P3_U6967);
  and ginst26203 (P3_U4028, P3_U6970, P3_U6972);
  and ginst26204 (P3_U4029, P3_U6975, P3_U6977);
  and ginst26205 (P3_U4030, P3_U4328, P3_U4329, P3_U4336);
  and ginst26206 (P3_U4031, P3_U4032, P3_U7097, P3_U7098);
  and ginst26207 (P3_U4032, P3_U7100, P3_U7101);
  and ginst26208 (P3_U4033, P3_U4034, P3_U7104);
  and ginst26209 (P3_U4034, P3_U7105, P3_U7106);
  and ginst26210 (P3_U4035, P3_U4036, P3_U7107, P3_U7108);
  and ginst26211 (P3_U4036, P3_U7110, P3_U7111);
  and ginst26212 (P3_U4037, P3_U4038, P3_U7114);
  and ginst26213 (P3_U4038, P3_U7115, P3_U7116);
  and ginst26214 (P3_U4039, P3_U4040, P3_U7117, P3_U7118);
  and ginst26215 (P3_U4040, P3_U7120, P3_U7121);
  and ginst26216 (P3_U4041, P3_U4042, P3_U7124);
  and ginst26217 (P3_U4042, P3_U7125, P3_U7126);
  and ginst26218 (P3_U4043, P3_U4044, P3_U7127, P3_U7128);
  and ginst26219 (P3_U4044, P3_U7130, P3_U7131);
  and ginst26220 (P3_U4045, P3_U4046, P3_U7134);
  and ginst26221 (P3_U4046, P3_U7135, P3_U7136);
  and ginst26222 (P3_U4047, P3_U4316, P3_U7137, P3_U7138);
  and ginst26223 (P3_U4048, P3_U7140, P3_U7141);
  and ginst26224 (P3_U4049, P3_U4050, P3_U7144);
  and ginst26225 (P3_U4050, P3_U7145, P3_U7146);
  and ginst26226 (P3_U4051, P3_U4047, P3_U4048, P3_U7139, P3_U7142, P3_U7143);
  and ginst26227 (P3_U4052, P3_U4316, P3_U7147, P3_U7148);
  and ginst26228 (P3_U4053, P3_U7150, P3_U7151);
  and ginst26229 (P3_U4054, P3_U4055, P3_U7154);
  and ginst26230 (P3_U4055, P3_U7155, P3_U7156);
  and ginst26231 (P3_U4056, P3_U4052, P3_U4053, P3_U7149, P3_U7152, P3_U7153);
  and ginst26232 (P3_U4057, P3_U4316, P3_U7157, P3_U7158);
  and ginst26233 (P3_U4058, P3_U4059, P3_U7161);
  and ginst26234 (P3_U4059, P3_U7163, P3_U7164);
  and ginst26235 (P3_U4060, P3_U4316, P3_U7165, P3_U7166);
  and ginst26236 (P3_U4061, P3_U4062, P3_U7169);
  and ginst26237 (P3_U4062, P3_U7171, P3_U7172);
  and ginst26238 (P3_U4063, P3_U4316, P3_U7173, P3_U7174);
  and ginst26239 (P3_U4064, P3_U4065, P3_U7177);
  and ginst26240 (P3_U4065, P3_U7179, P3_U7180);
  and ginst26241 (P3_U4066, P3_U4316, P3_U7181, P3_U7182);
  and ginst26242 (P3_U4067, P3_U4068, P3_U7185);
  and ginst26243 (P3_U4068, P3_U7187, P3_U7188);
  and ginst26244 (P3_U4069, P3_U4316, P3_U7189, P3_U7190);
  and ginst26245 (P3_U4070, P3_U4071, P3_U7193);
  and ginst26246 (P3_U4071, P3_U7195, P3_U7196);
  and ginst26247 (P3_U4072, P3_U4316, P3_U7197, P3_U7198);
  and ginst26248 (P3_U4073, P3_U4074, P3_U7201);
  and ginst26249 (P3_U4074, P3_U7203, P3_U7204);
  and ginst26250 (P3_U4075, P3_U4316, P3_U7205, P3_U7206);
  and ginst26251 (P3_U4076, P3_U4077, P3_U7209);
  and ginst26252 (P3_U4077, P3_U7211, P3_U7212);
  and ginst26253 (P3_U4078, P3_U4316, P3_U7213, P3_U7214);
  and ginst26254 (P3_U4079, P3_U4080, P3_U7217);
  and ginst26255 (P3_U4080, P3_U7219, P3_U7220);
  and ginst26256 (P3_U4081, P3_U4316, P3_U7221, P3_U7222);
  and ginst26257 (P3_U4082, P3_U4083, P3_U7225);
  and ginst26258 (P3_U4083, P3_U7227, P3_U7228);
  and ginst26259 (P3_U4084, P3_U4316, P3_U7229, P3_U7230);
  and ginst26260 (P3_U4085, P3_U4086, P3_U7233);
  and ginst26261 (P3_U4086, P3_U7235, P3_U7236);
  and ginst26262 (P3_U4087, P3_U4316, P3_U7237, P3_U7238);
  and ginst26263 (P3_U4088, P3_U4089, P3_U7241);
  and ginst26264 (P3_U4089, P3_U7243, P3_U7244);
  and ginst26265 (P3_U4090, P3_U4316, P3_U7245, P3_U7246);
  and ginst26266 (P3_U4091, P3_U4092, P3_U7249);
  and ginst26267 (P3_U4092, P3_U7251, P3_U7252);
  and ginst26268 (P3_U4093, P3_U4316, P3_U7253, P3_U7254);
  and ginst26269 (P3_U4094, P3_U4095, P3_U7257);
  and ginst26270 (P3_U4095, P3_U7259, P3_U7260);
  and ginst26271 (P3_U4096, P3_U4316, P3_U7261, P3_U7262);
  and ginst26272 (P3_U4097, P3_U4098, P3_U7265);
  and ginst26273 (P3_U4098, P3_U7267, P3_U7268);
  and ginst26274 (P3_U4099, P3_U7269, P3_U7270);
  and ginst26275 (P3_U4100, P3_U4101, P3_U7273);
  and ginst26276 (P3_U4101, P3_U7275, P3_U7276);
  and ginst26277 (P3_U4102, P3_U7277, P3_U7278);
  and ginst26278 (P3_U4103, P3_U4104, P3_U7281);
  and ginst26279 (P3_U4104, P3_U7283, P3_U7284);
  and ginst26280 (P3_U4105, P3_U7285, P3_U7286);
  and ginst26281 (P3_U4106, P3_U4107, P3_U7289);
  and ginst26282 (P3_U4107, P3_U7291, P3_U7292);
  and ginst26283 (P3_U4108, P3_U7293, P3_U7294);
  and ginst26284 (P3_U4109, P3_U4110, P3_U7297);
  and ginst26285 (P3_U4110, P3_U7299, P3_U7300);
  and ginst26286 (P3_U4111, P3_U7301, P3_U7302);
  and ginst26287 (P3_U4112, P3_U4113, P3_U7305);
  and ginst26288 (P3_U4113, P3_U7307, P3_U7308);
  and ginst26289 (P3_U4114, P3_U7309, P3_U7310);
  and ginst26290 (P3_U4115, P3_U4116, P3_U7313);
  and ginst26291 (P3_U4116, P3_U7315, P3_U7316);
  and ginst26292 (P3_U4117, P3_U7317, P3_U7318);
  and ginst26293 (P3_U4118, P3_U4119, P3_U7321);
  and ginst26294 (P3_U4119, P3_U7323, P3_U7324);
  and ginst26295 (P3_U4120, P3_U7325, P3_U7326);
  and ginst26296 (P3_U4121, P3_U4122, P3_U7329);
  and ginst26297 (P3_U4122, P3_U7331, P3_U7332);
  and ginst26298 (P3_U4123, P3_U7333, P3_U7334);
  and ginst26299 (P3_U4124, P3_U4125, P3_U7337);
  and ginst26300 (P3_U4125, P3_U7339, P3_U7340);
  and ginst26301 (P3_U4126, P3_U7341, P3_U7342);
  and ginst26302 (P3_U4127, P3_U4128, P3_U7345);
  and ginst26303 (P3_U4128, P3_U7347, P3_U7348);
  and ginst26304 (P3_U4129, P3_U7349, P3_U7350);
  and ginst26305 (P3_U4130, P3_U4131, P3_U7353);
  and ginst26306 (P3_U4131, P3_U7355, P3_U7356);
  and ginst26307 (P3_U4132, P3_U7364, P3_U7365);
  and ginst26308 (P3_U4133, P3_U4132, P3_U7361);
  and ginst26309 (P3_U4134, P3_U3259, P3_U7362);
  nor ginst26310 (P3_U4135, P3_SUB_320_U51, P3_U7363);
  nor ginst26311 (P3_U4136, P3_DATAWIDTH_REG_2__SCAN_IN, P3_DATAWIDTH_REG_3__SCAN_IN, P3_DATAWIDTH_REG_4__SCAN_IN, P3_DATAWIDTH_REG_5__SCAN_IN);
  nor ginst26312 (P3_U4137, P3_DATAWIDTH_REG_6__SCAN_IN, P3_DATAWIDTH_REG_7__SCAN_IN, P3_DATAWIDTH_REG_8__SCAN_IN, P3_DATAWIDTH_REG_9__SCAN_IN);
  and ginst26313 (P3_U4138, P3_U4136, P3_U4137);
  nor ginst26314 (P3_U4139, P3_DATAWIDTH_REG_10__SCAN_IN, P3_DATAWIDTH_REG_11__SCAN_IN, P3_DATAWIDTH_REG_12__SCAN_IN, P3_DATAWIDTH_REG_13__SCAN_IN);
  nor ginst26315 (P3_U4140, P3_DATAWIDTH_REG_14__SCAN_IN, P3_DATAWIDTH_REG_15__SCAN_IN, P3_DATAWIDTH_REG_16__SCAN_IN, P3_DATAWIDTH_REG_17__SCAN_IN);
  and ginst26316 (P3_U4141, P3_U4139, P3_U4140);
  nor ginst26317 (P3_U4142, P3_DATAWIDTH_REG_18__SCAN_IN, P3_DATAWIDTH_REG_19__SCAN_IN, P3_DATAWIDTH_REG_20__SCAN_IN, P3_DATAWIDTH_REG_21__SCAN_IN);
  nor ginst26318 (P3_U4143, P3_DATAWIDTH_REG_22__SCAN_IN, P3_DATAWIDTH_REG_23__SCAN_IN, P3_DATAWIDTH_REG_24__SCAN_IN, P3_DATAWIDTH_REG_25__SCAN_IN);
  and ginst26319 (P3_U4144, P3_U4142, P3_U4143);
  nor ginst26320 (P3_U4145, P3_DATAWIDTH_REG_26__SCAN_IN, P3_DATAWIDTH_REG_27__SCAN_IN);
  nor ginst26321 (P3_U4146, P3_DATAWIDTH_REG_28__SCAN_IN, P3_DATAWIDTH_REG_29__SCAN_IN);
  nor ginst26322 (P3_U4147, P3_DATAWIDTH_REG_30__SCAN_IN, P3_DATAWIDTH_REG_31__SCAN_IN);
  and ginst26323 (P3_U4148, P3_U4145, P3_U4146, P3_U4147, P3_U7366);
  nor ginst26324 (P3_U4149, P3_DATAWIDTH_REG_0__SCAN_IN, P3_DATAWIDTH_REG_1__SCAN_IN, P3_REIP_REG_0__SCAN_IN);
  and ginst26325 (P3_U4150, P3_U2630, P3_U7375);
  and ginst26326 (P3_U4151, P3_U3135, P3_U7373);
  and ginst26327 (P3_U4152, P3_U7387, P3_U7388, P3_U7389, P3_U7390);
  and ginst26328 (P3_U4153, P3_U7391, P3_U7392, P3_U7393, P3_U7394);
  and ginst26329 (P3_U4154, P3_U7395, P3_U7396, P3_U7397, P3_U7398);
  and ginst26330 (P3_U4155, P3_U7399, P3_U7400, P3_U7401, P3_U7402);
  and ginst26331 (P3_U4156, P3_U7403, P3_U7404, P3_U7405, P3_U7406);
  and ginst26332 (P3_U4157, P3_U7407, P3_U7408, P3_U7409, P3_U7410);
  and ginst26333 (P3_U4158, P3_U7411, P3_U7412, P3_U7413, P3_U7414);
  and ginst26334 (P3_U4159, P3_U7415, P3_U7416, P3_U7417, P3_U7418);
  and ginst26335 (P3_U4160, P3_U7419, P3_U7420, P3_U7421, P3_U7422);
  and ginst26336 (P3_U4161, P3_U7423, P3_U7424, P3_U7425, P3_U7426);
  and ginst26337 (P3_U4162, P3_U7427, P3_U7428, P3_U7429, P3_U7430);
  and ginst26338 (P3_U4163, P3_U7431, P3_U7432, P3_U7433, P3_U7434);
  and ginst26339 (P3_U4164, P3_U7435, P3_U7436, P3_U7437, P3_U7438);
  and ginst26340 (P3_U4165, P3_U7439, P3_U7440, P3_U7441, P3_U7442);
  and ginst26341 (P3_U4166, P3_U7443, P3_U7444, P3_U7445, P3_U7446);
  and ginst26342 (P3_U4167, P3_U7447, P3_U7448, P3_U7449, P3_U7450);
  and ginst26343 (P3_U4168, P3_U7451, P3_U7452, P3_U7453, P3_U7454);
  and ginst26344 (P3_U4169, P3_U7455, P3_U7456, P3_U7457, P3_U7458);
  and ginst26345 (P3_U4170, P3_U7459, P3_U7460, P3_U7461, P3_U7462);
  and ginst26346 (P3_U4171, P3_U7463, P3_U7464, P3_U7465, P3_U7466);
  and ginst26347 (P3_U4172, P3_U7467, P3_U7468, P3_U7469, P3_U7470);
  and ginst26348 (P3_U4173, P3_U7471, P3_U7472, P3_U7473, P3_U7474);
  and ginst26349 (P3_U4174, P3_U7475, P3_U7476, P3_U7477, P3_U7478);
  and ginst26350 (P3_U4175, P3_U7479, P3_U7480, P3_U7481, P3_U7482);
  and ginst26351 (P3_U4176, P3_U7483, P3_U7484, P3_U7485, P3_U7486);
  and ginst26352 (P3_U4177, P3_U7487, P3_U7488, P3_U7489, P3_U7490);
  and ginst26353 (P3_U4178, P3_U7491, P3_U7492, P3_U7493, P3_U7494);
  and ginst26354 (P3_U4179, P3_U7495, P3_U7496, P3_U7497, P3_U7498);
  and ginst26355 (P3_U4180, P3_U7499, P3_U7500, P3_U7501, P3_U7502);
  and ginst26356 (P3_U4181, P3_U7503, P3_U7504, P3_U7505, P3_U7506);
  and ginst26357 (P3_U4182, P3_U7507, P3_U7508, P3_U7509, P3_U7510);
  and ginst26358 (P3_U4183, P3_U7511, P3_U7512, P3_U7513, P3_U7514);
  and ginst26359 (P3_U4184, P3_U7517, P3_U7518, P3_U7519, P3_U7520);
  and ginst26360 (P3_U4185, P3_U7521, P3_U7522, P3_U7523, P3_U7524);
  and ginst26361 (P3_U4186, P3_U7525, P3_U7526, P3_U7527, P3_U7528);
  and ginst26362 (P3_U4187, P3_U7529, P3_U7530, P3_U7531, P3_U7532);
  and ginst26363 (P3_U4188, P3_U7533, P3_U7534, P3_U7535, P3_U7536);
  and ginst26364 (P3_U4189, P3_U7537, P3_U7538, P3_U7539, P3_U7540);
  and ginst26365 (P3_U4190, P3_U7541, P3_U7542, P3_U7543, P3_U7544);
  and ginst26366 (P3_U4191, P3_U7545, P3_U7546, P3_U7547, P3_U7548);
  and ginst26367 (P3_U4192, P3_U7549, P3_U7550, P3_U7551, P3_U7552);
  and ginst26368 (P3_U4193, P3_U7553, P3_U7554, P3_U7555, P3_U7556);
  and ginst26369 (P3_U4194, P3_U7557, P3_U7558, P3_U7559, P3_U7560);
  and ginst26370 (P3_U4195, P3_U7561, P3_U7562, P3_U7563, P3_U7564);
  and ginst26371 (P3_U4196, P3_U7565, P3_U7566, P3_U7567, P3_U7568);
  and ginst26372 (P3_U4197, P3_U7569, P3_U7570, P3_U7571, P3_U7572);
  and ginst26373 (P3_U4198, P3_U7573, P3_U7574, P3_U7575, P3_U7576);
  and ginst26374 (P3_U4199, P3_U7577, P3_U7578, P3_U7579, P3_U7580);
  and ginst26375 (P3_U4200, P3_U7581, P3_U7582, P3_U7583, P3_U7584);
  and ginst26376 (P3_U4201, P3_U7585, P3_U7586, P3_U7587, P3_U7588);
  and ginst26377 (P3_U4202, P3_U7589, P3_U7590, P3_U7591, P3_U7592);
  and ginst26378 (P3_U4203, P3_U7593, P3_U7594, P3_U7595, P3_U7596);
  and ginst26379 (P3_U4204, P3_U7597, P3_U7598, P3_U7599, P3_U7600);
  and ginst26380 (P3_U4205, P3_U7601, P3_U7602, P3_U7603, P3_U7604);
  and ginst26381 (P3_U4206, P3_U7605, P3_U7606, P3_U7607, P3_U7608);
  and ginst26382 (P3_U4207, P3_U7609, P3_U7610, P3_U7611, P3_U7612);
  and ginst26383 (P3_U4208, P3_U7613, P3_U7614, P3_U7615, P3_U7616);
  and ginst26384 (P3_U4209, P3_U7617, P3_U7618, P3_U7619, P3_U7620);
  and ginst26385 (P3_U4210, P3_U7621, P3_U7622, P3_U7623, P3_U7624);
  and ginst26386 (P3_U4211, P3_U7625, P3_U7626, P3_U7627, P3_U7628);
  and ginst26387 (P3_U4212, P3_U7629, P3_U7630, P3_U7631, P3_U7632);
  and ginst26388 (P3_U4213, P3_U7633, P3_U7634, P3_U7635, P3_U7636);
  and ginst26389 (P3_U4214, P3_U7637, P3_U7638, P3_U7639, P3_U7640);
  and ginst26390 (P3_U4215, P3_U7641, P3_U7642, P3_U7643, P3_U7644);
  and ginst26391 (P3_U4216, P3_U7646, P3_U7647, P3_U7648, P3_U7649);
  and ginst26392 (P3_U4217, P3_U7650, P3_U7651, P3_U7652, P3_U7653);
  and ginst26393 (P3_U4218, P3_U7654, P3_U7655, P3_U7656, P3_U7657);
  and ginst26394 (P3_U4219, P3_U7658, P3_U7659, P3_U7660, P3_U7661);
  and ginst26395 (P3_U4220, P3_U7662, P3_U7663, P3_U7664, P3_U7665);
  and ginst26396 (P3_U4221, P3_U7666, P3_U7667, P3_U7668, P3_U7669);
  and ginst26397 (P3_U4222, P3_U7670, P3_U7671, P3_U7672, P3_U7673);
  and ginst26398 (P3_U4223, P3_U7674, P3_U7675, P3_U7676, P3_U7677);
  and ginst26399 (P3_U4224, P3_U7678, P3_U7679, P3_U7680, P3_U7681);
  and ginst26400 (P3_U4225, P3_U7682, P3_U7683, P3_U7684, P3_U7685);
  and ginst26401 (P3_U4226, P3_U7686, P3_U7687, P3_U7688, P3_U7689);
  and ginst26402 (P3_U4227, P3_U7690, P3_U7691, P3_U7692, P3_U7693);
  and ginst26403 (P3_U4228, P3_U7694, P3_U7695, P3_U7696, P3_U7697);
  and ginst26404 (P3_U4229, P3_U7698, P3_U7699, P3_U7700, P3_U7701);
  and ginst26405 (P3_U4230, P3_U7702, P3_U7703, P3_U7704, P3_U7705);
  and ginst26406 (P3_U4231, P3_U7706, P3_U7707, P3_U7708, P3_U7709);
  and ginst26407 (P3_U4232, P3_U7710, P3_U7711, P3_U7712, P3_U7713);
  and ginst26408 (P3_U4233, P3_U7714, P3_U7715, P3_U7716, P3_U7717);
  and ginst26409 (P3_U4234, P3_U7718, P3_U7719, P3_U7720, P3_U7721);
  and ginst26410 (P3_U4235, P3_U7722, P3_U7723, P3_U7724, P3_U7725);
  and ginst26411 (P3_U4236, P3_U7726, P3_U7727, P3_U7728, P3_U7729);
  and ginst26412 (P3_U4237, P3_U7730, P3_U7731, P3_U7732, P3_U7733);
  and ginst26413 (P3_U4238, P3_U7734, P3_U7735, P3_U7736, P3_U7737);
  and ginst26414 (P3_U4239, P3_U7738, P3_U7739, P3_U7740, P3_U7741);
  and ginst26415 (P3_U4240, P3_U7742, P3_U7743, P3_U7744, P3_U7745);
  and ginst26416 (P3_U4241, P3_U7746, P3_U7747, P3_U7748, P3_U7749);
  and ginst26417 (P3_U4242, P3_U7750, P3_U7751, P3_U7752, P3_U7753);
  and ginst26418 (P3_U4243, P3_U7754, P3_U7755, P3_U7756, P3_U7757);
  and ginst26419 (P3_U4244, P3_U7758, P3_U7759, P3_U7760, P3_U7761);
  and ginst26420 (P3_U4245, P3_U7762, P3_U7763, P3_U7764, P3_U7765);
  and ginst26421 (P3_U4246, P3_U7766, P3_U7767, P3_U7768, P3_U7769);
  and ginst26422 (P3_U4247, P3_U7770, P3_U7771, P3_U7772, P3_U7773);
  and ginst26423 (P3_U4248, P3_U7776, P3_U7777, P3_U7778, P3_U7779);
  and ginst26424 (P3_U4249, P3_U7780, P3_U7781, P3_U7782, P3_U7783);
  and ginst26425 (P3_U4250, P3_U7784, P3_U7785, P3_U7786, P3_U7787);
  and ginst26426 (P3_U4251, P3_U7788, P3_U7789, P3_U7790, P3_U7791);
  and ginst26427 (P3_U4252, P3_U7792, P3_U7793, P3_U7794, P3_U7795);
  and ginst26428 (P3_U4253, P3_U7796, P3_U7797, P3_U7798, P3_U7799);
  and ginst26429 (P3_U4254, P3_U7800, P3_U7801, P3_U7802, P3_U7803);
  and ginst26430 (P3_U4255, P3_U7804, P3_U7805, P3_U7806, P3_U7807);
  and ginst26431 (P3_U4256, P3_U7808, P3_U7809, P3_U7810, P3_U7811);
  and ginst26432 (P3_U4257, P3_U7812, P3_U7813, P3_U7814, P3_U7815);
  and ginst26433 (P3_U4258, P3_U7816, P3_U7817, P3_U7818, P3_U7819);
  and ginst26434 (P3_U4259, P3_U7820, P3_U7821, P3_U7822, P3_U7823);
  and ginst26435 (P3_U4260, P3_U7824, P3_U7825, P3_U7826, P3_U7827);
  and ginst26436 (P3_U4261, P3_U7828, P3_U7829, P3_U7830, P3_U7831);
  and ginst26437 (P3_U4262, P3_U7832, P3_U7833, P3_U7834, P3_U7835);
  and ginst26438 (P3_U4263, P3_U7836, P3_U7837, P3_U7838, P3_U7839);
  and ginst26439 (P3_U4264, P3_U7840, P3_U7841, P3_U7842, P3_U7843);
  and ginst26440 (P3_U4265, P3_U7844, P3_U7845, P3_U7846, P3_U7847);
  and ginst26441 (P3_U4266, P3_U7848, P3_U7849, P3_U7850, P3_U7851);
  and ginst26442 (P3_U4267, P3_U7852, P3_U7853, P3_U7854, P3_U7855);
  and ginst26443 (P3_U4268, P3_U7856, P3_U7857, P3_U7858, P3_U7859);
  and ginst26444 (P3_U4269, P3_U7860, P3_U7861, P3_U7862, P3_U7863);
  and ginst26445 (P3_U4270, P3_U7864, P3_U7865, P3_U7866, P3_U7867);
  and ginst26446 (P3_U4271, P3_U7868, P3_U7869, P3_U7870, P3_U7871);
  and ginst26447 (P3_U4272, P3_U7872, P3_U7873, P3_U7874, P3_U7875);
  and ginst26448 (P3_U4273, P3_U7876, P3_U7877, P3_U7878, P3_U7879);
  and ginst26449 (P3_U4274, P3_U7880, P3_U7881, P3_U7882, P3_U7883);
  and ginst26450 (P3_U4275, P3_U7884, P3_U7885, P3_U7886, P3_U7887);
  and ginst26451 (P3_U4276, P3_U7888, P3_U7889, P3_U7890, P3_U7891);
  and ginst26452 (P3_U4277, P3_U7892, P3_U7893, P3_U7894, P3_U7895);
  and ginst26453 (P3_U4278, P3_U7896, P3_U7897, P3_U7898, P3_U7899);
  and ginst26454 (P3_U4279, P3_U7900, P3_U7901, P3_U7902, P3_U7903);
  and ginst26455 (P3_U4280, P3_U7942, P3_U7943);
  nand ginst26456 (P3_U4281, P3_U2604, P3_U3361);
  and ginst26457 (P3_U4282, P3_U7950, P3_U7951);
  nand ginst26458 (P3_U4283, P3_U3658, P3_U5497);
  not ginst26459 (P3_U4284, P3_INSTADDRPOINTER_REG_31__SCAN_IN);
  nand ginst26460 (P3_U4285, P3_U2390, P3_U4281);
  not ginst26461 (P3_U4286, BS16);
  nand ginst26462 (P3_U4287, P3_U4151, P3_U4334);
  nand ginst26463 (P3_U4288, P3_U3239, P3_U4334);
  nand ginst26464 (P3_U4289, P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN, P3_U3091);
  nand ginst26465 (P3_U4290, P3_U2515, P3_U2516, P3_U3657);
  not ginst26466 (P3_U4291, P3_U3267);
  nand ginst26467 (P3_U4292, HOLD, P3_U2630);
  not ginst26468 (P3_U4293, P3_U3105);
  not ginst26469 (P3_U4294, P3_U3106);
  not ginst26470 (P3_U4295, P3_U3135);
  not ginst26471 (P3_U4296, P3_U3112);
  not ginst26472 (P3_U4297, P3_U3111);
  not ginst26473 (P3_U4298, P3_U3242);
  not ginst26474 (P3_U4299, P3_U3243);
  not ginst26475 (P3_U4300, P3_U3244);
  not ginst26476 (P3_U4301, P3_U3245);
  not ginst26477 (P3_U4302, P3_U3119);
  not ginst26478 (P3_U4303, P3_U3117);
  not ginst26479 (P3_U4304, P3_U3116);
  not ginst26480 (P3_U4305, P3_U3115);
  not ginst26481 (P3_U4306, P3_U3246);
  not ginst26482 (P3_U4307, P3_U3261);
  not ginst26483 (P3_U4308, P3_U3077);
  not ginst26484 (P3_U4309, P3_U3253);
  not ginst26485 (P3_U4310, P3_U3252);
  not ginst26486 (P3_U4311, P3_U3250);
  not ginst26487 (P3_U4312, P3_U3127);
  not ginst26488 (P3_U4313, P3_LT_563_1260_U6);
  not ginst26489 (P3_U4314, P3_U3217);
  nand ginst26490 (P3_U4315, P3_U2631, P3_U4295);
  nand ginst26491 (P3_U4316, P3_U3260, P3_U4347);
  nand ginst26492 (P3_U4317, P3_U2383, P3_U3105);
  not ginst26493 (P3_U4318, P3_U3247);
  not ginst26494 (P3_U4319, P3_U3259);
  not ginst26495 (P3_U4320, P3_U3080);
  not ginst26496 (P3_U4321, P3_U3078);
  not ginst26497 (P3_U4322, P3_U3136);
  not ginst26498 (P3_U4323, P3_U3114);
  not ginst26499 (P3_U4324, P3_U3118);
  not ginst26500 (P3_U4325, P3_U3219);
  not ginst26501 (P3_U4326, P3_U3181);
  nand ginst26502 (P3_U4327, P3_U4149, P3_U4307);
  nand ginst26503 (P3_U4328, P3_U3365, P3_U4354);
  nand ginst26504 (P3_U4329, P3_STATE2_REG_1__SCAN_IN, P3_U2631, P3_U3090, P3_U3121);
  nand ginst26505 (P3_U4330, P3_U2453, P3_U3653);
  nand ginst26506 (P3_U4331, P3_U2458, P3_U4653);
  not ginst26507 (P3_U4332, P3_U3095);
  nand ginst26508 (P3_U4333, P3_U3113, P3_U4350);
  nand ginst26509 (P3_U4334, P3_U2390, P3_U7093);
  nand ginst26510 (P3_U4335, P3_U3085, P3_U4452);
  nand ginst26511 (P3_U4336, P3_U3121, P3_U4347);
  nand ginst26512 (P3_U4337, P3_U2453, P3_U3232);
  nand ginst26513 (P3_U4338, P3_STATE2_REG_0__SCAN_IN, P3_U3090, U209);
  nand ginst26514 (P3_U4339, P3_U3654, P3_U4608);
  not ginst26515 (P3_U4340, P3_U3123);
  not ginst26516 (P3_U4341, P3_U3229);
  not ginst26517 (P3_U4342, P3_U3150);
  not ginst26518 (P3_U4343, P3_U3158);
  not ginst26519 (P3_U4344, P3_U3103);
  not ginst26520 (P3_U4345, P3_U3126);
  not ginst26521 (P3_U4346, P3_U3082);
  not ginst26522 (P3_U4347, P3_U3239);
  not ginst26523 (P3_U4348, P3_U3236);
  not ginst26524 (P3_U4349, P3_U3235);
  not ginst26525 (P3_U4350, P3_U3208);
  not ginst26526 (P3_U4351, P3_U3216);
  not ginst26527 (P3_U4352, P3_U3222);
  not ginst26528 (P3_U4353, P3_U3124);
  not ginst26529 (P3_U4354, P3_U3125);
  nand ginst26530 (P3_U4355, P3_REIP_REG_31__SCAN_IN, P3_U4321);
  nand ginst26531 (P3_U4356, P3_REIP_REG_30__SCAN_IN, P3_U4320);
  nand ginst26532 (P3_U4357, P3_ADDRESS_REG_29__SCAN_IN, P3_U3077);
  nand ginst26533 (P3_U4358, P3_REIP_REG_30__SCAN_IN, P3_U4321);
  nand ginst26534 (P3_U4359, P3_REIP_REG_29__SCAN_IN, P3_U4320);
  nand ginst26535 (P3_U4360, P3_ADDRESS_REG_28__SCAN_IN, P3_U3077);
  nand ginst26536 (P3_U4361, P3_REIP_REG_29__SCAN_IN, P3_U4321);
  nand ginst26537 (P3_U4362, P3_REIP_REG_28__SCAN_IN, P3_U4320);
  nand ginst26538 (P3_U4363, P3_ADDRESS_REG_27__SCAN_IN, P3_U3077);
  nand ginst26539 (P3_U4364, P3_REIP_REG_28__SCAN_IN, P3_U4321);
  nand ginst26540 (P3_U4365, P3_REIP_REG_27__SCAN_IN, P3_U4320);
  nand ginst26541 (P3_U4366, P3_ADDRESS_REG_26__SCAN_IN, P3_U3077);
  nand ginst26542 (P3_U4367, P3_REIP_REG_27__SCAN_IN, P3_U4321);
  nand ginst26543 (P3_U4368, P3_REIP_REG_26__SCAN_IN, P3_U4320);
  nand ginst26544 (P3_U4369, P3_ADDRESS_REG_25__SCAN_IN, P3_U3077);
  nand ginst26545 (P3_U4370, P3_REIP_REG_26__SCAN_IN, P3_U4321);
  nand ginst26546 (P3_U4371, P3_REIP_REG_25__SCAN_IN, P3_U4320);
  nand ginst26547 (P3_U4372, P3_ADDRESS_REG_24__SCAN_IN, P3_U3077);
  nand ginst26548 (P3_U4373, P3_REIP_REG_25__SCAN_IN, P3_U4321);
  nand ginst26549 (P3_U4374, P3_REIP_REG_24__SCAN_IN, P3_U4320);
  nand ginst26550 (P3_U4375, P3_ADDRESS_REG_23__SCAN_IN, P3_U3077);
  nand ginst26551 (P3_U4376, P3_REIP_REG_24__SCAN_IN, P3_U4321);
  nand ginst26552 (P3_U4377, P3_REIP_REG_23__SCAN_IN, P3_U4320);
  nand ginst26553 (P3_U4378, P3_ADDRESS_REG_22__SCAN_IN, P3_U3077);
  nand ginst26554 (P3_U4379, P3_REIP_REG_23__SCAN_IN, P3_U4321);
  nand ginst26555 (P3_U4380, P3_REIP_REG_22__SCAN_IN, P3_U4320);
  nand ginst26556 (P3_U4381, P3_ADDRESS_REG_21__SCAN_IN, P3_U3077);
  nand ginst26557 (P3_U4382, P3_REIP_REG_22__SCAN_IN, P3_U4321);
  nand ginst26558 (P3_U4383, P3_REIP_REG_21__SCAN_IN, P3_U4320);
  nand ginst26559 (P3_U4384, P3_ADDRESS_REG_20__SCAN_IN, P3_U3077);
  nand ginst26560 (P3_U4385, P3_REIP_REG_21__SCAN_IN, P3_U4321);
  nand ginst26561 (P3_U4386, P3_REIP_REG_20__SCAN_IN, P3_U4320);
  nand ginst26562 (P3_U4387, P3_ADDRESS_REG_19__SCAN_IN, P3_U3077);
  nand ginst26563 (P3_U4388, P3_REIP_REG_20__SCAN_IN, P3_U4321);
  nand ginst26564 (P3_U4389, P3_REIP_REG_19__SCAN_IN, P3_U4320);
  nand ginst26565 (P3_U4390, P3_ADDRESS_REG_18__SCAN_IN, P3_U3077);
  nand ginst26566 (P3_U4391, P3_REIP_REG_19__SCAN_IN, P3_U4321);
  nand ginst26567 (P3_U4392, P3_REIP_REG_18__SCAN_IN, P3_U4320);
  nand ginst26568 (P3_U4393, P3_ADDRESS_REG_17__SCAN_IN, P3_U3077);
  nand ginst26569 (P3_U4394, P3_REIP_REG_18__SCAN_IN, P3_U4321);
  nand ginst26570 (P3_U4395, P3_REIP_REG_17__SCAN_IN, P3_U4320);
  nand ginst26571 (P3_U4396, P3_ADDRESS_REG_16__SCAN_IN, P3_U3077);
  nand ginst26572 (P3_U4397, P3_REIP_REG_17__SCAN_IN, P3_U4321);
  nand ginst26573 (P3_U4398, P3_REIP_REG_16__SCAN_IN, P3_U4320);
  nand ginst26574 (P3_U4399, P3_ADDRESS_REG_15__SCAN_IN, P3_U3077);
  nand ginst26575 (P3_U4400, P3_REIP_REG_16__SCAN_IN, P3_U4321);
  nand ginst26576 (P3_U4401, P3_REIP_REG_15__SCAN_IN, P3_U4320);
  nand ginst26577 (P3_U4402, P3_ADDRESS_REG_14__SCAN_IN, P3_U3077);
  nand ginst26578 (P3_U4403, P3_REIP_REG_15__SCAN_IN, P3_U4321);
  nand ginst26579 (P3_U4404, P3_REIP_REG_14__SCAN_IN, P3_U4320);
  nand ginst26580 (P3_U4405, P3_ADDRESS_REG_13__SCAN_IN, P3_U3077);
  nand ginst26581 (P3_U4406, P3_REIP_REG_14__SCAN_IN, P3_U4321);
  nand ginst26582 (P3_U4407, P3_REIP_REG_13__SCAN_IN, P3_U4320);
  nand ginst26583 (P3_U4408, P3_ADDRESS_REG_12__SCAN_IN, P3_U3077);
  nand ginst26584 (P3_U4409, P3_REIP_REG_13__SCAN_IN, P3_U4321);
  nand ginst26585 (P3_U4410, P3_REIP_REG_12__SCAN_IN, P3_U4320);
  nand ginst26586 (P3_U4411, P3_ADDRESS_REG_11__SCAN_IN, P3_U3077);
  nand ginst26587 (P3_U4412, P3_REIP_REG_12__SCAN_IN, P3_U4321);
  nand ginst26588 (P3_U4413, P3_REIP_REG_11__SCAN_IN, P3_U4320);
  nand ginst26589 (P3_U4414, P3_ADDRESS_REG_10__SCAN_IN, P3_U3077);
  nand ginst26590 (P3_U4415, P3_REIP_REG_11__SCAN_IN, P3_U4321);
  nand ginst26591 (P3_U4416, P3_REIP_REG_10__SCAN_IN, P3_U4320);
  nand ginst26592 (P3_U4417, P3_ADDRESS_REG_9__SCAN_IN, P3_U3077);
  nand ginst26593 (P3_U4418, P3_REIP_REG_10__SCAN_IN, P3_U4321);
  nand ginst26594 (P3_U4419, P3_REIP_REG_9__SCAN_IN, P3_U4320);
  nand ginst26595 (P3_U4420, P3_ADDRESS_REG_8__SCAN_IN, P3_U3077);
  nand ginst26596 (P3_U4421, P3_REIP_REG_9__SCAN_IN, P3_U4321);
  nand ginst26597 (P3_U4422, P3_REIP_REG_8__SCAN_IN, P3_U4320);
  nand ginst26598 (P3_U4423, P3_ADDRESS_REG_7__SCAN_IN, P3_U3077);
  nand ginst26599 (P3_U4424, P3_REIP_REG_8__SCAN_IN, P3_U4321);
  nand ginst26600 (P3_U4425, P3_REIP_REG_7__SCAN_IN, P3_U4320);
  nand ginst26601 (P3_U4426, P3_ADDRESS_REG_6__SCAN_IN, P3_U3077);
  nand ginst26602 (P3_U4427, P3_REIP_REG_7__SCAN_IN, P3_U4321);
  nand ginst26603 (P3_U4428, P3_REIP_REG_6__SCAN_IN, P3_U4320);
  nand ginst26604 (P3_U4429, P3_ADDRESS_REG_5__SCAN_IN, P3_U3077);
  nand ginst26605 (P3_U4430, P3_REIP_REG_6__SCAN_IN, P3_U4321);
  nand ginst26606 (P3_U4431, P3_REIP_REG_5__SCAN_IN, P3_U4320);
  nand ginst26607 (P3_U4432, P3_ADDRESS_REG_4__SCAN_IN, P3_U3077);
  nand ginst26608 (P3_U4433, P3_REIP_REG_5__SCAN_IN, P3_U4321);
  nand ginst26609 (P3_U4434, P3_REIP_REG_4__SCAN_IN, P3_U4320);
  nand ginst26610 (P3_U4435, P3_ADDRESS_REG_3__SCAN_IN, P3_U3077);
  nand ginst26611 (P3_U4436, P3_REIP_REG_4__SCAN_IN, P3_U4321);
  nand ginst26612 (P3_U4437, P3_REIP_REG_3__SCAN_IN, P3_U4320);
  nand ginst26613 (P3_U4438, P3_ADDRESS_REG_2__SCAN_IN, P3_U3077);
  nand ginst26614 (P3_U4439, P3_REIP_REG_3__SCAN_IN, P3_U4321);
  nand ginst26615 (P3_U4440, P3_REIP_REG_2__SCAN_IN, P3_U4320);
  nand ginst26616 (P3_U4441, P3_ADDRESS_REG_1__SCAN_IN, P3_U3077);
  nand ginst26617 (P3_U4442, P3_REIP_REG_2__SCAN_IN, P3_U4321);
  nand ginst26618 (P3_U4443, P3_REIP_REG_1__SCAN_IN, P3_U4320);
  nand ginst26619 (P3_U4444, P3_ADDRESS_REG_0__SCAN_IN, P3_U3077);
  not ginst26620 (P3_U4445, P3_U3087);
  nand ginst26621 (P3_U4446, P3_U2630, P3_U4445);
  nand ginst26622 (P3_U4447, NA, P3_U4346);
  not ginst26623 (P3_U4448, P3_U3088);
  nand ginst26624 (P3_U4449, P3_U2630, P3_U4448);
  or ginst26625 (P3_U4450, NA, P3_STATE_REG_0__SCAN_IN);
  nand ginst26626 (P3_U4451, P3_U4450, P3_U7912, P3_U7913);
  not ginst26627 (P3_U4452, P3_U3083);
  nand ginst26628 (P3_U4453, P3_U3088, P3_U4346, U209);
  nand ginst26629 (P3_U4454, HOLD, P3_U3075, P3_U4452);
  nand ginst26630 (P3_U4455, P3_U4453, P3_U4454);
  nand ginst26631 (P3_U4456, P3_U3309, P3_U4455);
  nand ginst26632 (P3_U4457, P3_STATE_REG_2__SCAN_IN, P3_U4451);
  nand ginst26633 (P3_U4458, P3_U4308, U209);
  nand ginst26634 (P3_U4459, P3_U3312, P3_U7915);
  nand ginst26635 (P3_U4460, P3_STATE_REG_2__SCAN_IN, P3_U3087);
  nand ginst26636 (P3_U4461, NA, P3_U3085);
  nand ginst26637 (P3_U4462, P3_U4460, P3_U4461);
  nand ginst26638 (P3_U4463, P3_U3076, P3_U4462);
  nand ginst26639 (P3_U4464, P3_U3083, P3_U4286);
  nand ginst26640 (P3_U4465, P3_STATE_REG_2__SCAN_IN, P3_U3076);
  nand ginst26641 (P3_U4466, P3_U3082, P3_U4465);
  not ginst26642 (P3_U4467, P3_U3091);
  not ginst26643 (P3_U4468, P3_U3096);
  not ginst26644 (P3_U4469, P3_U3092);
  not ginst26645 (P3_U4470, P3_U3098);
  not ginst26646 (P3_U4471, P3_U3099);
  nand ginst26647 (P3_U4472, P3_INSTQUEUE_REG_0__0__SCAN_IN, P3_U2484);
  nand ginst26648 (P3_U4473, P3_INSTQUEUE_REG_1__0__SCAN_IN, P3_U2483);
  nand ginst26649 (P3_U4474, P3_INSTQUEUE_REG_2__0__SCAN_IN, P3_U2482);
  nand ginst26650 (P3_U4475, P3_INSTQUEUE_REG_3__0__SCAN_IN, P3_U2480);
  nand ginst26651 (P3_U4476, P3_INSTQUEUE_REG_4__0__SCAN_IN, P3_U2479);
  nand ginst26652 (P3_U4477, P3_INSTQUEUE_REG_5__0__SCAN_IN, P3_U2478);
  nand ginst26653 (P3_U4478, P3_INSTQUEUE_REG_6__0__SCAN_IN, P3_U2477);
  nand ginst26654 (P3_U4479, P3_INSTQUEUE_REG_7__0__SCAN_IN, P3_U4471);
  nand ginst26655 (P3_U4480, P3_INSTQUEUE_REG_8__0__SCAN_IN, P3_U2476);
  nand ginst26656 (P3_U4481, P3_INSTQUEUE_REG_9__0__SCAN_IN, P3_U2475);
  nand ginst26657 (P3_U4482, P3_INSTQUEUE_REG_10__0__SCAN_IN, P3_U2473);
  nand ginst26658 (P3_U4483, P3_INSTQUEUE_REG_11__0__SCAN_IN, P3_U2471);
  nand ginst26659 (P3_U4484, P3_INSTQUEUE_REG_12__0__SCAN_IN, P3_U2470);
  nand ginst26660 (P3_U4485, P3_INSTQUEUE_REG_13__0__SCAN_IN, P3_U2469);
  nand ginst26661 (P3_U4486, P3_INSTQUEUE_REG_14__0__SCAN_IN, P3_U2467);
  nand ginst26662 (P3_U4487, P3_INSTQUEUE_REG_15__0__SCAN_IN, P3_U2465);
  not ginst26663 (P3_U4488, P3_U3108);
  nand ginst26664 (P3_U4489, P3_INSTQUEUE_REG_0__1__SCAN_IN, P3_U2484);
  nand ginst26665 (P3_U4490, P3_INSTQUEUE_REG_1__1__SCAN_IN, P3_U2483);
  nand ginst26666 (P3_U4491, P3_INSTQUEUE_REG_2__1__SCAN_IN, P3_U2482);
  nand ginst26667 (P3_U4492, P3_INSTQUEUE_REG_3__1__SCAN_IN, P3_U2480);
  nand ginst26668 (P3_U4493, P3_INSTQUEUE_REG_4__1__SCAN_IN, P3_U2479);
  nand ginst26669 (P3_U4494, P3_INSTQUEUE_REG_5__1__SCAN_IN, P3_U2478);
  nand ginst26670 (P3_U4495, P3_INSTQUEUE_REG_6__1__SCAN_IN, P3_U2477);
  nand ginst26671 (P3_U4496, P3_INSTQUEUE_REG_7__1__SCAN_IN, P3_U4471);
  nand ginst26672 (P3_U4497, P3_INSTQUEUE_REG_8__1__SCAN_IN, P3_U2476);
  nand ginst26673 (P3_U4498, P3_INSTQUEUE_REG_9__1__SCAN_IN, P3_U2475);
  nand ginst26674 (P3_U4499, P3_INSTQUEUE_REG_10__1__SCAN_IN, P3_U2473);
  nand ginst26675 (P3_U4500, P3_INSTQUEUE_REG_11__1__SCAN_IN, P3_U2471);
  nand ginst26676 (P3_U4501, P3_INSTQUEUE_REG_12__1__SCAN_IN, P3_U2470);
  nand ginst26677 (P3_U4502, P3_INSTQUEUE_REG_13__1__SCAN_IN, P3_U2469);
  nand ginst26678 (P3_U4503, P3_INSTQUEUE_REG_14__1__SCAN_IN, P3_U2467);
  nand ginst26679 (P3_U4504, P3_INSTQUEUE_REG_15__1__SCAN_IN, P3_U2465);
  not ginst26680 (P3_U4505, P3_U3104);
  nand ginst26681 (P3_U4506, P3_INSTQUEUE_REG_0__4__SCAN_IN, P3_U2484);
  nand ginst26682 (P3_U4507, P3_INSTQUEUE_REG_1__4__SCAN_IN, P3_U2483);
  nand ginst26683 (P3_U4508, P3_INSTQUEUE_REG_2__4__SCAN_IN, P3_U2482);
  nand ginst26684 (P3_U4509, P3_INSTQUEUE_REG_3__4__SCAN_IN, P3_U2480);
  nand ginst26685 (P3_U4510, P3_INSTQUEUE_REG_4__4__SCAN_IN, P3_U2479);
  nand ginst26686 (P3_U4511, P3_INSTQUEUE_REG_5__4__SCAN_IN, P3_U2478);
  nand ginst26687 (P3_U4512, P3_INSTQUEUE_REG_6__4__SCAN_IN, P3_U2477);
  nand ginst26688 (P3_U4513, P3_INSTQUEUE_REG_7__4__SCAN_IN, P3_U4471);
  nand ginst26689 (P3_U4514, P3_INSTQUEUE_REG_8__4__SCAN_IN, P3_U2476);
  nand ginst26690 (P3_U4515, P3_INSTQUEUE_REG_9__4__SCAN_IN, P3_U2475);
  nand ginst26691 (P3_U4516, P3_INSTQUEUE_REG_10__4__SCAN_IN, P3_U2473);
  nand ginst26692 (P3_U4517, P3_INSTQUEUE_REG_11__4__SCAN_IN, P3_U2471);
  nand ginst26693 (P3_U4518, P3_INSTQUEUE_REG_12__4__SCAN_IN, P3_U2470);
  nand ginst26694 (P3_U4519, P3_INSTQUEUE_REG_13__4__SCAN_IN, P3_U2469);
  nand ginst26695 (P3_U4520, P3_INSTQUEUE_REG_14__4__SCAN_IN, P3_U2467);
  nand ginst26696 (P3_U4521, P3_INSTQUEUE_REG_15__4__SCAN_IN, P3_U2465);
  not ginst26697 (P3_U4522, P3_U3102);
  nand ginst26698 (P3_U4523, P3_INSTQUEUE_REG_0__2__SCAN_IN, P3_U2484);
  nand ginst26699 (P3_U4524, P3_INSTQUEUE_REG_1__2__SCAN_IN, P3_U2483);
  nand ginst26700 (P3_U4525, P3_INSTQUEUE_REG_2__2__SCAN_IN, P3_U2482);
  nand ginst26701 (P3_U4526, P3_INSTQUEUE_REG_3__2__SCAN_IN, P3_U2480);
  nand ginst26702 (P3_U4527, P3_INSTQUEUE_REG_4__2__SCAN_IN, P3_U2479);
  nand ginst26703 (P3_U4528, P3_INSTQUEUE_REG_5__2__SCAN_IN, P3_U2478);
  nand ginst26704 (P3_U4529, P3_INSTQUEUE_REG_6__2__SCAN_IN, P3_U2477);
  nand ginst26705 (P3_U4530, P3_INSTQUEUE_REG_7__2__SCAN_IN, P3_U4471);
  nand ginst26706 (P3_U4531, P3_INSTQUEUE_REG_8__2__SCAN_IN, P3_U2476);
  nand ginst26707 (P3_U4532, P3_INSTQUEUE_REG_9__2__SCAN_IN, P3_U2475);
  nand ginst26708 (P3_U4533, P3_INSTQUEUE_REG_10__2__SCAN_IN, P3_U2473);
  nand ginst26709 (P3_U4534, P3_INSTQUEUE_REG_11__2__SCAN_IN, P3_U2471);
  nand ginst26710 (P3_U4535, P3_INSTQUEUE_REG_12__2__SCAN_IN, P3_U2470);
  nand ginst26711 (P3_U4536, P3_INSTQUEUE_REG_13__2__SCAN_IN, P3_U2469);
  nand ginst26712 (P3_U4537, P3_INSTQUEUE_REG_14__2__SCAN_IN, P3_U2467);
  nand ginst26713 (P3_U4538, P3_INSTQUEUE_REG_15__2__SCAN_IN, P3_U2465);
  not ginst26714 (P3_U4539, P3_U3101);
  nand ginst26715 (P3_U4540, P3_INSTQUEUE_REG_0__3__SCAN_IN, P3_U2484);
  nand ginst26716 (P3_U4541, P3_INSTQUEUE_REG_1__3__SCAN_IN, P3_U2483);
  nand ginst26717 (P3_U4542, P3_INSTQUEUE_REG_2__3__SCAN_IN, P3_U2482);
  nand ginst26718 (P3_U4543, P3_INSTQUEUE_REG_3__3__SCAN_IN, P3_U2480);
  nand ginst26719 (P3_U4544, P3_INSTQUEUE_REG_4__3__SCAN_IN, P3_U2479);
  nand ginst26720 (P3_U4545, P3_INSTQUEUE_REG_5__3__SCAN_IN, P3_U2478);
  nand ginst26721 (P3_U4546, P3_INSTQUEUE_REG_6__3__SCAN_IN, P3_U2477);
  nand ginst26722 (P3_U4547, P3_INSTQUEUE_REG_7__3__SCAN_IN, P3_U4471);
  nand ginst26723 (P3_U4548, P3_INSTQUEUE_REG_8__3__SCAN_IN, P3_U2476);
  nand ginst26724 (P3_U4549, P3_INSTQUEUE_REG_9__3__SCAN_IN, P3_U2475);
  nand ginst26725 (P3_U4550, P3_INSTQUEUE_REG_10__3__SCAN_IN, P3_U2473);
  nand ginst26726 (P3_U4551, P3_INSTQUEUE_REG_11__3__SCAN_IN, P3_U2471);
  nand ginst26727 (P3_U4552, P3_INSTQUEUE_REG_12__3__SCAN_IN, P3_U2470);
  nand ginst26728 (P3_U4553, P3_INSTQUEUE_REG_13__3__SCAN_IN, P3_U2469);
  nand ginst26729 (P3_U4554, P3_INSTQUEUE_REG_14__3__SCAN_IN, P3_U2467);
  nand ginst26730 (P3_U4555, P3_INSTQUEUE_REG_15__3__SCAN_IN, P3_U2465);
  not ginst26731 (P3_U4556, P3_U3107);
  nand ginst26732 (P3_U4557, P3_INSTQUEUE_REG_0__7__SCAN_IN, P3_U2484);
  nand ginst26733 (P3_U4558, P3_INSTQUEUE_REG_1__7__SCAN_IN, P3_U2483);
  nand ginst26734 (P3_U4559, P3_INSTQUEUE_REG_2__7__SCAN_IN, P3_U2482);
  nand ginst26735 (P3_U4560, P3_INSTQUEUE_REG_3__7__SCAN_IN, P3_U2480);
  nand ginst26736 (P3_U4561, P3_INSTQUEUE_REG_4__7__SCAN_IN, P3_U2479);
  nand ginst26737 (P3_U4562, P3_INSTQUEUE_REG_5__7__SCAN_IN, P3_U2478);
  nand ginst26738 (P3_U4563, P3_INSTQUEUE_REG_6__7__SCAN_IN, P3_U2477);
  nand ginst26739 (P3_U4564, P3_INSTQUEUE_REG_7__7__SCAN_IN, P3_U4471);
  nand ginst26740 (P3_U4565, P3_INSTQUEUE_REG_8__7__SCAN_IN, P3_U2476);
  nand ginst26741 (P3_U4566, P3_INSTQUEUE_REG_9__7__SCAN_IN, P3_U2475);
  nand ginst26742 (P3_U4567, P3_INSTQUEUE_REG_10__7__SCAN_IN, P3_U2473);
  nand ginst26743 (P3_U4568, P3_INSTQUEUE_REG_11__7__SCAN_IN, P3_U2471);
  nand ginst26744 (P3_U4569, P3_INSTQUEUE_REG_12__7__SCAN_IN, P3_U2470);
  nand ginst26745 (P3_U4570, P3_INSTQUEUE_REG_13__7__SCAN_IN, P3_U2469);
  nand ginst26746 (P3_U4571, P3_INSTQUEUE_REG_14__7__SCAN_IN, P3_U2467);
  nand ginst26747 (P3_U4572, P3_INSTQUEUE_REG_15__7__SCAN_IN, P3_U2465);
  not ginst26748 (P3_U4573, P3_U3218);
  nand ginst26749 (P3_U4574, P3_INSTQUEUE_REG_0__5__SCAN_IN, P3_U2484);
  nand ginst26750 (P3_U4575, P3_INSTQUEUE_REG_1__5__SCAN_IN, P3_U2483);
  nand ginst26751 (P3_U4576, P3_INSTQUEUE_REG_2__5__SCAN_IN, P3_U2482);
  nand ginst26752 (P3_U4577, P3_INSTQUEUE_REG_3__5__SCAN_IN, P3_U2480);
  nand ginst26753 (P3_U4578, P3_INSTQUEUE_REG_4__5__SCAN_IN, P3_U2479);
  nand ginst26754 (P3_U4579, P3_INSTQUEUE_REG_5__5__SCAN_IN, P3_U2478);
  nand ginst26755 (P3_U4580, P3_INSTQUEUE_REG_6__5__SCAN_IN, P3_U2477);
  nand ginst26756 (P3_U4581, P3_INSTQUEUE_REG_7__5__SCAN_IN, P3_U4471);
  nand ginst26757 (P3_U4582, P3_INSTQUEUE_REG_8__5__SCAN_IN, P3_U2476);
  nand ginst26758 (P3_U4583, P3_INSTQUEUE_REG_9__5__SCAN_IN, P3_U2475);
  nand ginst26759 (P3_U4584, P3_INSTQUEUE_REG_10__5__SCAN_IN, P3_U2473);
  nand ginst26760 (P3_U4585, P3_INSTQUEUE_REG_11__5__SCAN_IN, P3_U2471);
  nand ginst26761 (P3_U4586, P3_INSTQUEUE_REG_12__5__SCAN_IN, P3_U2470);
  nand ginst26762 (P3_U4587, P3_INSTQUEUE_REG_13__5__SCAN_IN, P3_U2469);
  nand ginst26763 (P3_U4588, P3_INSTQUEUE_REG_14__5__SCAN_IN, P3_U2467);
  nand ginst26764 (P3_U4589, P3_INSTQUEUE_REG_15__5__SCAN_IN, P3_U2465);
  not ginst26765 (P3_U4590, P3_U3110);
  nand ginst26766 (P3_U4591, P3_INSTQUEUE_REG_0__6__SCAN_IN, P3_U2484);
  nand ginst26767 (P3_U4592, P3_INSTQUEUE_REG_1__6__SCAN_IN, P3_U2483);
  nand ginst26768 (P3_U4593, P3_INSTQUEUE_REG_2__6__SCAN_IN, P3_U2482);
  nand ginst26769 (P3_U4594, P3_INSTQUEUE_REG_3__6__SCAN_IN, P3_U2480);
  nand ginst26770 (P3_U4595, P3_INSTQUEUE_REG_4__6__SCAN_IN, P3_U2479);
  nand ginst26771 (P3_U4596, P3_INSTQUEUE_REG_5__6__SCAN_IN, P3_U2478);
  nand ginst26772 (P3_U4597, P3_INSTQUEUE_REG_6__6__SCAN_IN, P3_U2477);
  nand ginst26773 (P3_U4598, P3_INSTQUEUE_REG_7__6__SCAN_IN, P3_U4471);
  nand ginst26774 (P3_U4599, P3_INSTQUEUE_REG_8__6__SCAN_IN, P3_U2476);
  nand ginst26775 (P3_U4600, P3_INSTQUEUE_REG_9__6__SCAN_IN, P3_U2475);
  nand ginst26776 (P3_U4601, P3_INSTQUEUE_REG_10__6__SCAN_IN, P3_U2473);
  nand ginst26777 (P3_U4602, P3_INSTQUEUE_REG_11__6__SCAN_IN, P3_U2471);
  nand ginst26778 (P3_U4603, P3_INSTQUEUE_REG_12__6__SCAN_IN, P3_U2470);
  nand ginst26779 (P3_U4604, P3_INSTQUEUE_REG_13__6__SCAN_IN, P3_U2469);
  nand ginst26780 (P3_U4605, P3_INSTQUEUE_REG_14__6__SCAN_IN, P3_U2467);
  nand ginst26781 (P3_U4606, P3_INSTQUEUE_REG_15__6__SCAN_IN, P3_U2465);
  not ginst26782 (P3_U4607, P3_U3074);
  not ginst26783 (P3_U4608, P3_U3113);
  nand ginst26784 (P3_U4609, P3_U2361, P3_U3238);
  nand ginst26785 (P3_U4610, P3_U2360, P3_U3237);
  nand ginst26786 (P3_U4611, P3_U2357, P3_U3212);
  nand ginst26787 (P3_U4612, P3_U3215, P3_U4305);
  nand ginst26788 (P3_U4613, P3_U3210, P3_U4304);
  nand ginst26789 (P3_U4614, P3_U3213, P3_U4303);
  nand ginst26790 (P3_U4615, P3_U2356, P3_U3211);
  nand ginst26791 (P3_U4616, P3_U3214, P3_U4302);
  nand ginst26792 (P3_U4617, P3_U3357, P3_U3358);
  nand ginst26793 (P3_U4618, P3_U2463, P3_U3360, P3_U4522, P3_U7944, P3_U7945);
  not ginst26794 (P3_U4619, P3_U3109);
  nand ginst26795 (P3_U4620, P3_U4280, P3_U4619);
  nand ginst26796 (P3_U4621, P3_U3359, P3_U7916);
  not ginst26797 (P3_U4622, P3_U4281);
  not ginst26798 (P3_U4623, P3_U3262);
  or ginst26799 (P3_U4624, P3_FLUSH_REG_SCAN_IN, P3_MORE_REG_SCAN_IN);
  not ginst26800 (P3_U4625, P3_U3120);
  nand ginst26801 (P3_U4626, P3_U3353, P3_U4303);
  nand ginst26802 (P3_U4627, P3_U3362, P3_U4625);
  nand ginst26803 (P3_U4628, P3_STATE2_REG_1__SCAN_IN, U209);
  nand ginst26804 (P3_U4629, P3_STATE2_REG_2__SCAN_IN, P3_U7952, P3_U7953);
  not ginst26805 (P3_U4630, P3_U3122);
  nand ginst26806 (P3_U4631, P3_STATE2_REG_1__SCAN_IN, P3_U7956, P3_U7957);
  nand ginst26807 (P3_U4632, P3_STATE2_REG_2__SCAN_IN, P3_U3122);
  nand ginst26808 (P3_U4633, P3_U4338, P3_U4629);
  nand ginst26809 (P3_U4634, P3_U3364, P3_U4630);
  nand ginst26810 (P3_U4635, P3_STATE2_REG_1__SCAN_IN, P3_U4633);
  nand ginst26811 (P3_U4636, P3_U2390, P3_U4629);
  nand ginst26812 (P3_U4637, P3_U4345, P3_U4354);
  nand ginst26813 (P3_U4638, P3_U4337, P3_U4629);
  nand ginst26814 (P3_U4639, P3_U2390, P3_U3120);
  not ginst26815 (P3_U4640, P3_U3153);
  nand ginst26816 (P3_U4641, P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN, P3_U3128);
  not ginst26817 (P3_U4642, P3_U3137);
  not ginst26818 (P3_U4643, P3_U3141);
  not ginst26819 (P3_U4644, P3_U3148);
  not ginst26820 (P3_U4645, P3_U3155);
  not ginst26821 (P3_U4646, P3_U3156);
  not ginst26822 (P3_U4647, P3_U3143);
  not ginst26823 (P3_U4648, P3_U3130);
  not ginst26824 (P3_U4649, P3_U3132);
  not ginst26825 (P3_U4650, P3_U3180);
  nand ginst26826 (P3_U4651, P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN, P3_U3132);
  not ginst26827 (P3_U4652, P3_U3139);
  not ginst26828 (P3_U4653, P3_U3138);
  nand ginst26829 (P3_U4654, P3_U3269, P3_U4653);
  nand ginst26830 (P3_U4655, P3_U3139, P3_U4654);
  not ginst26831 (P3_U4656, P3_U3142);
  not ginst26832 (P3_U4657, P3_U3140);
  not ginst26833 (P3_U4658, P3_U3165);
  nand ginst26834 (P3_U4659, P3_U3140, P3_U3142);
  not ginst26835 (P3_U4660, P3_U3182);
  not ginst26836 (P3_U4661, P3_U3144);
  not ginst26837 (P3_U4662, P3_U3134);
  nand ginst26838 (P3_U4663, P3_U2457, P3_U4653);
  not ginst26839 (P3_U4664, P3_U3146);
  nand ginst26840 (P3_U4665, P3_STATE2_REG_1__SCAN_IN, P3_U3090);
  nand ginst26841 (P3_U4666, P3_U3124, P3_U3126, P3_U4665);
  nand ginst26842 (P3_U4667, P3_U2487, P3_U4657);
  not ginst26843 (P3_U4668, P3_U3145);
  nand ginst26844 (P3_U4669, P3_U2489, P3_U3145);
  nand ginst26845 (P3_U4670, P3_U4664, P3_U4669);
  nand ginst26846 (P3_U4671, P3_STATE2_REG_3__SCAN_IN, P3_U3134);
  nand ginst26847 (P3_U4672, P3_U3369, P3_U4670);
  nand ginst26848 (P3_U4673, P3_U4322, P3_U4668);
  nand ginst26849 (P3_U4674, P3_U2489, P3_U4673);
  nand ginst26850 (P3_U4675, P3_U2445, P3_U4662);
  nand ginst26851 (P3_U4676, P3_U2436, P3_U2488);
  nand ginst26852 (P3_U4677, P3_U2435, P3_U4661);
  nand ginst26853 (P3_U4678, P3_U2378, P3_U2420);
  nand ginst26854 (P3_U4679, P3_INSTQUEUE_REG_15__7__SCAN_IN, P3_U4672);
  nand ginst26855 (P3_U4680, P3_U2443, P3_U4662);
  nand ginst26856 (P3_U4681, P3_U2434, P3_U2488);
  nand ginst26857 (P3_U4682, P3_U2433, P3_U4661);
  nand ginst26858 (P3_U4683, P3_U2378, P3_U2419);
  nand ginst26859 (P3_U4684, P3_INSTQUEUE_REG_15__6__SCAN_IN, P3_U4672);
  nand ginst26860 (P3_U4685, P3_U2442, P3_U4662);
  nand ginst26861 (P3_U4686, P3_U2432, P3_U2488);
  nand ginst26862 (P3_U4687, P3_U2431, P3_U4661);
  nand ginst26863 (P3_U4688, P3_U2378, P3_U2418);
  nand ginst26864 (P3_U4689, P3_INSTQUEUE_REG_15__5__SCAN_IN, P3_U4672);
  nand ginst26865 (P3_U4690, P3_U2441, P3_U4662);
  nand ginst26866 (P3_U4691, P3_U2430, P3_U2488);
  nand ginst26867 (P3_U4692, P3_U2429, P3_U4661);
  nand ginst26868 (P3_U4693, P3_U2378, P3_U2417);
  nand ginst26869 (P3_U4694, P3_INSTQUEUE_REG_15__4__SCAN_IN, P3_U4672);
  nand ginst26870 (P3_U4695, P3_U2440, P3_U4662);
  nand ginst26871 (P3_U4696, P3_U2428, P3_U2488);
  nand ginst26872 (P3_U4697, P3_U2427, P3_U4661);
  nand ginst26873 (P3_U4698, P3_U2378, P3_U2416);
  nand ginst26874 (P3_U4699, P3_INSTQUEUE_REG_15__3__SCAN_IN, P3_U4672);
  nand ginst26875 (P3_U4700, P3_U2439, P3_U4662);
  nand ginst26876 (P3_U4701, P3_U2426, P3_U2488);
  nand ginst26877 (P3_U4702, P3_U2425, P3_U4661);
  nand ginst26878 (P3_U4703, P3_U2378, P3_U2415);
  nand ginst26879 (P3_U4704, P3_INSTQUEUE_REG_15__2__SCAN_IN, P3_U4672);
  nand ginst26880 (P3_U4705, P3_U2438, P3_U4662);
  nand ginst26881 (P3_U4706, P3_U2424, P3_U2488);
  nand ginst26882 (P3_U4707, P3_U2423, P3_U4661);
  nand ginst26883 (P3_U4708, P3_U2378, P3_U2414);
  nand ginst26884 (P3_U4709, P3_INSTQUEUE_REG_15__1__SCAN_IN, P3_U4672);
  nand ginst26885 (P3_U4710, P3_U2437, P3_U4662);
  nand ginst26886 (P3_U4711, P3_U2422, P3_U2488);
  nand ginst26887 (P3_U4712, P3_U2421, P3_U4661);
  nand ginst26888 (P3_U4713, P3_U2378, P3_U2413);
  nand ginst26889 (P3_U4714, P3_INSTQUEUE_REG_15__0__SCAN_IN, P3_U4672);
  not ginst26890 (P3_U4715, P3_U3149);
  not ginst26891 (P3_U4716, P3_U3147);
  nand ginst26892 (P3_U4717, P3_U2457, P3_U4342);
  not ginst26893 (P3_U4718, P3_U3152);
  nand ginst26894 (P3_U4719, P3_U2487, P3_U4644);
  not ginst26895 (P3_U4720, P3_U3151);
  nand ginst26896 (P3_U4721, P3_U2489, P3_U3151);
  nand ginst26897 (P3_U4722, P3_U4718, P3_U4721);
  nand ginst26898 (P3_U4723, P3_STATE2_REG_3__SCAN_IN, P3_U3147);
  nand ginst26899 (P3_U4724, P3_U3387, P3_U4722);
  nand ginst26900 (P3_U4725, P3_U4322, P3_U4720);
  nand ginst26901 (P3_U4726, P3_U2489, P3_U4725);
  nand ginst26902 (P3_U4727, P3_U2445, P3_U4716);
  nand ginst26903 (P3_U4728, P3_U2436, P3_U2491);
  nand ginst26904 (P3_U4729, P3_U2435, P3_U4715);
  nand ginst26905 (P3_U4730, P3_U2377, P3_U2420);
  nand ginst26906 (P3_U4731, P3_INSTQUEUE_REG_14__7__SCAN_IN, P3_U4724);
  nand ginst26907 (P3_U4732, P3_U2443, P3_U4716);
  nand ginst26908 (P3_U4733, P3_U2434, P3_U2491);
  nand ginst26909 (P3_U4734, P3_U2433, P3_U4715);
  nand ginst26910 (P3_U4735, P3_U2377, P3_U2419);
  nand ginst26911 (P3_U4736, P3_INSTQUEUE_REG_14__6__SCAN_IN, P3_U4724);
  nand ginst26912 (P3_U4737, P3_U2442, P3_U4716);
  nand ginst26913 (P3_U4738, P3_U2432, P3_U2491);
  nand ginst26914 (P3_U4739, P3_U2431, P3_U4715);
  nand ginst26915 (P3_U4740, P3_U2377, P3_U2418);
  nand ginst26916 (P3_U4741, P3_INSTQUEUE_REG_14__5__SCAN_IN, P3_U4724);
  nand ginst26917 (P3_U4742, P3_U2441, P3_U4716);
  nand ginst26918 (P3_U4743, P3_U2430, P3_U2491);
  nand ginst26919 (P3_U4744, P3_U2429, P3_U4715);
  nand ginst26920 (P3_U4745, P3_U2377, P3_U2417);
  nand ginst26921 (P3_U4746, P3_INSTQUEUE_REG_14__4__SCAN_IN, P3_U4724);
  nand ginst26922 (P3_U4747, P3_U2440, P3_U4716);
  nand ginst26923 (P3_U4748, P3_U2428, P3_U2491);
  nand ginst26924 (P3_U4749, P3_U2427, P3_U4715);
  nand ginst26925 (P3_U4750, P3_U2377, P3_U2416);
  nand ginst26926 (P3_U4751, P3_INSTQUEUE_REG_14__3__SCAN_IN, P3_U4724);
  nand ginst26927 (P3_U4752, P3_U2439, P3_U4716);
  nand ginst26928 (P3_U4753, P3_U2426, P3_U2491);
  nand ginst26929 (P3_U4754, P3_U2425, P3_U4715);
  nand ginst26930 (P3_U4755, P3_U2377, P3_U2415);
  nand ginst26931 (P3_U4756, P3_INSTQUEUE_REG_14__2__SCAN_IN, P3_U4724);
  nand ginst26932 (P3_U4757, P3_U2438, P3_U4716);
  nand ginst26933 (P3_U4758, P3_U2424, P3_U2491);
  nand ginst26934 (P3_U4759, P3_U2423, P3_U4715);
  nand ginst26935 (P3_U4760, P3_U2377, P3_U2414);
  nand ginst26936 (P3_U4761, P3_INSTQUEUE_REG_14__1__SCAN_IN, P3_U4724);
  nand ginst26937 (P3_U4762, P3_U2437, P3_U4716);
  nand ginst26938 (P3_U4763, P3_U2422, P3_U2491);
  nand ginst26939 (P3_U4764, P3_U2421, P3_U4715);
  nand ginst26940 (P3_U4765, P3_U2377, P3_U2413);
  nand ginst26941 (P3_U4766, P3_INSTQUEUE_REG_14__0__SCAN_IN, P3_U4724);
  not ginst26942 (P3_U4767, P3_U3157);
  not ginst26943 (P3_U4768, P3_U3154);
  nand ginst26944 (P3_U4769, P3_U2457, P3_U4343);
  not ginst26945 (P3_U4770, P3_U3160);
  nand ginst26946 (P3_U4771, P3_U2487, P3_U4645);
  not ginst26947 (P3_U4772, P3_U3159);
  nand ginst26948 (P3_U4773, P3_U2489, P3_U3159);
  nand ginst26949 (P3_U4774, P3_U4770, P3_U4773);
  nand ginst26950 (P3_U4775, P3_STATE2_REG_3__SCAN_IN, P3_U3154);
  nand ginst26951 (P3_U4776, P3_U3405, P3_U4774);
  nand ginst26952 (P3_U4777, P3_U4322, P3_U4772);
  nand ginst26953 (P3_U4778, P3_U2489, P3_U4777);
  nand ginst26954 (P3_U4779, P3_U2445, P3_U4768);
  nand ginst26955 (P3_U4780, P3_U2436, P3_U2494);
  nand ginst26956 (P3_U4781, P3_U2435, P3_U4767);
  nand ginst26957 (P3_U4782, P3_U2376, P3_U2420);
  nand ginst26958 (P3_U4783, P3_INSTQUEUE_REG_13__7__SCAN_IN, P3_U4776);
  nand ginst26959 (P3_U4784, P3_U2443, P3_U4768);
  nand ginst26960 (P3_U4785, P3_U2434, P3_U2494);
  nand ginst26961 (P3_U4786, P3_U2433, P3_U4767);
  nand ginst26962 (P3_U4787, P3_U2376, P3_U2419);
  nand ginst26963 (P3_U4788, P3_INSTQUEUE_REG_13__6__SCAN_IN, P3_U4776);
  nand ginst26964 (P3_U4789, P3_U2442, P3_U4768);
  nand ginst26965 (P3_U4790, P3_U2432, P3_U2494);
  nand ginst26966 (P3_U4791, P3_U2431, P3_U4767);
  nand ginst26967 (P3_U4792, P3_U2376, P3_U2418);
  nand ginst26968 (P3_U4793, P3_INSTQUEUE_REG_13__5__SCAN_IN, P3_U4776);
  nand ginst26969 (P3_U4794, P3_U2441, P3_U4768);
  nand ginst26970 (P3_U4795, P3_U2430, P3_U2494);
  nand ginst26971 (P3_U4796, P3_U2429, P3_U4767);
  nand ginst26972 (P3_U4797, P3_U2376, P3_U2417);
  nand ginst26973 (P3_U4798, P3_INSTQUEUE_REG_13__4__SCAN_IN, P3_U4776);
  nand ginst26974 (P3_U4799, P3_U2440, P3_U4768);
  nand ginst26975 (P3_U4800, P3_U2428, P3_U2494);
  nand ginst26976 (P3_U4801, P3_U2427, P3_U4767);
  nand ginst26977 (P3_U4802, P3_U2376, P3_U2416);
  nand ginst26978 (P3_U4803, P3_INSTQUEUE_REG_13__3__SCAN_IN, P3_U4776);
  nand ginst26979 (P3_U4804, P3_U2439, P3_U4768);
  nand ginst26980 (P3_U4805, P3_U2426, P3_U2494);
  nand ginst26981 (P3_U4806, P3_U2425, P3_U4767);
  nand ginst26982 (P3_U4807, P3_U2376, P3_U2415);
  nand ginst26983 (P3_U4808, P3_INSTQUEUE_REG_13__2__SCAN_IN, P3_U4776);
  nand ginst26984 (P3_U4809, P3_U2438, P3_U4768);
  nand ginst26985 (P3_U4810, P3_U2424, P3_U2494);
  nand ginst26986 (P3_U4811, P3_U2423, P3_U4767);
  nand ginst26987 (P3_U4812, P3_U2376, P3_U2414);
  nand ginst26988 (P3_U4813, P3_INSTQUEUE_REG_13__1__SCAN_IN, P3_U4776);
  nand ginst26989 (P3_U4814, P3_U2437, P3_U4768);
  nand ginst26990 (P3_U4815, P3_U2422, P3_U2494);
  nand ginst26991 (P3_U4816, P3_U2421, P3_U4767);
  nand ginst26992 (P3_U4817, P3_U2376, P3_U2413);
  nand ginst26993 (P3_U4818, P3_INSTQUEUE_REG_13__0__SCAN_IN, P3_U4776);
  not ginst26994 (P3_U4819, P3_U3162);
  not ginst26995 (P3_U4820, P3_U3161);
  not ginst26996 (P3_U4821, P3_U3070);
  nand ginst26997 (P3_U4822, P3_U2487, P3_U2496);
  not ginst26998 (P3_U4823, P3_U3163);
  nand ginst26999 (P3_U4824, P3_U2489, P3_U3163);
  nand ginst27000 (P3_U4825, P3_U3070, P3_U4824);
  nand ginst27001 (P3_U4826, P3_STATE2_REG_3__SCAN_IN, P3_U3161);
  nand ginst27002 (P3_U4827, P3_U3423, P3_U4825);
  nand ginst27003 (P3_U4828, P3_U4322, P3_U4823);
  nand ginst27004 (P3_U4829, P3_U2489, P3_U4828);
  nand ginst27005 (P3_U4830, P3_U2445, P3_U4820);
  nand ginst27006 (P3_U4831, P3_U2436, P3_U2497);
  nand ginst27007 (P3_U4832, P3_U2435, P3_U4819);
  nand ginst27008 (P3_U4833, P3_U2375, P3_U2420);
  nand ginst27009 (P3_U4834, P3_INSTQUEUE_REG_12__7__SCAN_IN, P3_U4827);
  nand ginst27010 (P3_U4835, P3_U2443, P3_U4820);
  nand ginst27011 (P3_U4836, P3_U2434, P3_U2497);
  nand ginst27012 (P3_U4837, P3_U2433, P3_U4819);
  nand ginst27013 (P3_U4838, P3_U2375, P3_U2419);
  nand ginst27014 (P3_U4839, P3_INSTQUEUE_REG_12__6__SCAN_IN, P3_U4827);
  nand ginst27015 (P3_U4840, P3_U2442, P3_U4820);
  nand ginst27016 (P3_U4841, P3_U2432, P3_U2497);
  nand ginst27017 (P3_U4842, P3_U2431, P3_U4819);
  nand ginst27018 (P3_U4843, P3_U2375, P3_U2418);
  nand ginst27019 (P3_U4844, P3_INSTQUEUE_REG_12__5__SCAN_IN, P3_U4827);
  nand ginst27020 (P3_U4845, P3_U2441, P3_U4820);
  nand ginst27021 (P3_U4846, P3_U2430, P3_U2497);
  nand ginst27022 (P3_U4847, P3_U2429, P3_U4819);
  nand ginst27023 (P3_U4848, P3_U2375, P3_U2417);
  nand ginst27024 (P3_U4849, P3_INSTQUEUE_REG_12__4__SCAN_IN, P3_U4827);
  nand ginst27025 (P3_U4850, P3_U2440, P3_U4820);
  nand ginst27026 (P3_U4851, P3_U2428, P3_U2497);
  nand ginst27027 (P3_U4852, P3_U2427, P3_U4819);
  nand ginst27028 (P3_U4853, P3_U2375, P3_U2416);
  nand ginst27029 (P3_U4854, P3_INSTQUEUE_REG_12__3__SCAN_IN, P3_U4827);
  nand ginst27030 (P3_U4855, P3_U2439, P3_U4820);
  nand ginst27031 (P3_U4856, P3_U2426, P3_U2497);
  nand ginst27032 (P3_U4857, P3_U2425, P3_U4819);
  nand ginst27033 (P3_U4858, P3_U2375, P3_U2415);
  nand ginst27034 (P3_U4859, P3_INSTQUEUE_REG_12__2__SCAN_IN, P3_U4827);
  nand ginst27035 (P3_U4860, P3_U2438, P3_U4820);
  nand ginst27036 (P3_U4861, P3_U2424, P3_U2497);
  nand ginst27037 (P3_U4862, P3_U2423, P3_U4819);
  nand ginst27038 (P3_U4863, P3_U2375, P3_U2414);
  nand ginst27039 (P3_U4864, P3_INSTQUEUE_REG_12__1__SCAN_IN, P3_U4827);
  nand ginst27040 (P3_U4865, P3_U2437, P3_U4820);
  nand ginst27041 (P3_U4866, P3_U2422, P3_U2497);
  nand ginst27042 (P3_U4867, P3_U2421, P3_U4819);
  nand ginst27043 (P3_U4868, P3_U2375, P3_U2413);
  nand ginst27044 (P3_U4869, P3_INSTQUEUE_REG_12__0__SCAN_IN, P3_U4827);
  not ginst27045 (P3_U4870, P3_U3166);
  not ginst27046 (P3_U4871, P3_U3164);
  nand ginst27047 (P3_U4872, P3_U2459, P3_U4653);
  not ginst27048 (P3_U4873, P3_U3168);
  nand ginst27049 (P3_U4874, P3_U4657, P3_U4658);
  not ginst27050 (P3_U4875, P3_U3167);
  nand ginst27051 (P3_U4876, P3_U2489, P3_U3167);
  nand ginst27052 (P3_U4877, P3_U4873, P3_U4876);
  nand ginst27053 (P3_U4878, P3_STATE2_REG_3__SCAN_IN, P3_U3164);
  nand ginst27054 (P3_U4879, P3_U3440, P3_U4877);
  nand ginst27055 (P3_U4880, P3_U4322, P3_U4875);
  nand ginst27056 (P3_U4881, P3_U2489, P3_U4880);
  nand ginst27057 (P3_U4882, P3_U2445, P3_U4871);
  nand ginst27058 (P3_U4883, P3_U2436, P3_U2499);
  nand ginst27059 (P3_U4884, P3_U2435, P3_U4870);
  nand ginst27060 (P3_U4885, P3_U2374, P3_U2420);
  nand ginst27061 (P3_U4886, P3_INSTQUEUE_REG_11__7__SCAN_IN, P3_U4879);
  nand ginst27062 (P3_U4887, P3_U2443, P3_U4871);
  nand ginst27063 (P3_U4888, P3_U2434, P3_U2499);
  nand ginst27064 (P3_U4889, P3_U2433, P3_U4870);
  nand ginst27065 (P3_U4890, P3_U2374, P3_U2419);
  nand ginst27066 (P3_U4891, P3_INSTQUEUE_REG_11__6__SCAN_IN, P3_U4879);
  nand ginst27067 (P3_U4892, P3_U2442, P3_U4871);
  nand ginst27068 (P3_U4893, P3_U2432, P3_U2499);
  nand ginst27069 (P3_U4894, P3_U2431, P3_U4870);
  nand ginst27070 (P3_U4895, P3_U2374, P3_U2418);
  nand ginst27071 (P3_U4896, P3_INSTQUEUE_REG_11__5__SCAN_IN, P3_U4879);
  nand ginst27072 (P3_U4897, P3_U2441, P3_U4871);
  nand ginst27073 (P3_U4898, P3_U2430, P3_U2499);
  nand ginst27074 (P3_U4899, P3_U2429, P3_U4870);
  nand ginst27075 (P3_U4900, P3_U2374, P3_U2417);
  nand ginst27076 (P3_U4901, P3_INSTQUEUE_REG_11__4__SCAN_IN, P3_U4879);
  nand ginst27077 (P3_U4902, P3_U2440, P3_U4871);
  nand ginst27078 (P3_U4903, P3_U2428, P3_U2499);
  nand ginst27079 (P3_U4904, P3_U2427, P3_U4870);
  nand ginst27080 (P3_U4905, P3_U2374, P3_U2416);
  nand ginst27081 (P3_U4906, P3_INSTQUEUE_REG_11__3__SCAN_IN, P3_U4879);
  nand ginst27082 (P3_U4907, P3_U2439, P3_U4871);
  nand ginst27083 (P3_U4908, P3_U2426, P3_U2499);
  nand ginst27084 (P3_U4909, P3_U2425, P3_U4870);
  nand ginst27085 (P3_U4910, P3_U2374, P3_U2415);
  nand ginst27086 (P3_U4911, P3_INSTQUEUE_REG_11__2__SCAN_IN, P3_U4879);
  nand ginst27087 (P3_U4912, P3_U2438, P3_U4871);
  nand ginst27088 (P3_U4913, P3_U2424, P3_U2499);
  nand ginst27089 (P3_U4914, P3_U2423, P3_U4870);
  nand ginst27090 (P3_U4915, P3_U2374, P3_U2414);
  nand ginst27091 (P3_U4916, P3_INSTQUEUE_REG_11__1__SCAN_IN, P3_U4879);
  nand ginst27092 (P3_U4917, P3_U2437, P3_U4871);
  nand ginst27093 (P3_U4918, P3_U2422, P3_U2499);
  nand ginst27094 (P3_U4919, P3_U2421, P3_U4870);
  nand ginst27095 (P3_U4920, P3_U2374, P3_U2413);
  nand ginst27096 (P3_U4921, P3_INSTQUEUE_REG_11__0__SCAN_IN, P3_U4879);
  not ginst27097 (P3_U4922, P3_U3170);
  not ginst27098 (P3_U4923, P3_U3169);
  nand ginst27099 (P3_U4924, P3_U2459, P3_U4342);
  not ginst27100 (P3_U4925, P3_U3172);
  nand ginst27101 (P3_U4926, P3_U4644, P3_U4658);
  not ginst27102 (P3_U4927, P3_U3171);
  nand ginst27103 (P3_U4928, P3_U2489, P3_U3171);
  nand ginst27104 (P3_U4929, P3_U4925, P3_U4928);
  nand ginst27105 (P3_U4930, P3_STATE2_REG_3__SCAN_IN, P3_U3169);
  nand ginst27106 (P3_U4931, P3_U3458, P3_U4929);
  nand ginst27107 (P3_U4932, P3_U4322, P3_U4927);
  nand ginst27108 (P3_U4933, P3_U2489, P3_U4932);
  nand ginst27109 (P3_U4934, P3_U2445, P3_U4923);
  nand ginst27110 (P3_U4935, P3_U2436, P3_U2500);
  nand ginst27111 (P3_U4936, P3_U2435, P3_U4922);
  nand ginst27112 (P3_U4937, P3_U2373, P3_U2420);
  nand ginst27113 (P3_U4938, P3_INSTQUEUE_REG_10__7__SCAN_IN, P3_U4931);
  nand ginst27114 (P3_U4939, P3_U2443, P3_U4923);
  nand ginst27115 (P3_U4940, P3_U2434, P3_U2500);
  nand ginst27116 (P3_U4941, P3_U2433, P3_U4922);
  nand ginst27117 (P3_U4942, P3_U2373, P3_U2419);
  nand ginst27118 (P3_U4943, P3_INSTQUEUE_REG_10__6__SCAN_IN, P3_U4931);
  nand ginst27119 (P3_U4944, P3_U2442, P3_U4923);
  nand ginst27120 (P3_U4945, P3_U2432, P3_U2500);
  nand ginst27121 (P3_U4946, P3_U2431, P3_U4922);
  nand ginst27122 (P3_U4947, P3_U2373, P3_U2418);
  nand ginst27123 (P3_U4948, P3_INSTQUEUE_REG_10__5__SCAN_IN, P3_U4931);
  nand ginst27124 (P3_U4949, P3_U2441, P3_U4923);
  nand ginst27125 (P3_U4950, P3_U2430, P3_U2500);
  nand ginst27126 (P3_U4951, P3_U2429, P3_U4922);
  nand ginst27127 (P3_U4952, P3_U2373, P3_U2417);
  nand ginst27128 (P3_U4953, P3_INSTQUEUE_REG_10__4__SCAN_IN, P3_U4931);
  nand ginst27129 (P3_U4954, P3_U2440, P3_U4923);
  nand ginst27130 (P3_U4955, P3_U2428, P3_U2500);
  nand ginst27131 (P3_U4956, P3_U2427, P3_U4922);
  nand ginst27132 (P3_U4957, P3_U2373, P3_U2416);
  nand ginst27133 (P3_U4958, P3_INSTQUEUE_REG_10__3__SCAN_IN, P3_U4931);
  nand ginst27134 (P3_U4959, P3_U2439, P3_U4923);
  nand ginst27135 (P3_U4960, P3_U2426, P3_U2500);
  nand ginst27136 (P3_U4961, P3_U2425, P3_U4922);
  nand ginst27137 (P3_U4962, P3_U2373, P3_U2415);
  nand ginst27138 (P3_U4963, P3_INSTQUEUE_REG_10__2__SCAN_IN, P3_U4931);
  nand ginst27139 (P3_U4964, P3_U2438, P3_U4923);
  nand ginst27140 (P3_U4965, P3_U2424, P3_U2500);
  nand ginst27141 (P3_U4966, P3_U2423, P3_U4922);
  nand ginst27142 (P3_U4967, P3_U2373, P3_U2414);
  nand ginst27143 (P3_U4968, P3_INSTQUEUE_REG_10__1__SCAN_IN, P3_U4931);
  nand ginst27144 (P3_U4969, P3_U2437, P3_U4923);
  nand ginst27145 (P3_U4970, P3_U2422, P3_U2500);
  nand ginst27146 (P3_U4971, P3_U2421, P3_U4922);
  nand ginst27147 (P3_U4972, P3_U2373, P3_U2413);
  nand ginst27148 (P3_U4973, P3_INSTQUEUE_REG_10__0__SCAN_IN, P3_U4931);
  not ginst27149 (P3_U4974, P3_U3174);
  not ginst27150 (P3_U4975, P3_U3173);
  nand ginst27151 (P3_U4976, P3_U2459, P3_U4343);
  not ginst27152 (P3_U4977, P3_U3176);
  nand ginst27153 (P3_U4978, P3_U4645, P3_U4658);
  not ginst27154 (P3_U4979, P3_U3175);
  nand ginst27155 (P3_U4980, P3_U2489, P3_U3175);
  nand ginst27156 (P3_U4981, P3_U4977, P3_U4980);
  nand ginst27157 (P3_U4982, P3_STATE2_REG_3__SCAN_IN, P3_U3173);
  nand ginst27158 (P3_U4983, P3_U3476, P3_U4981);
  nand ginst27159 (P3_U4984, P3_U4322, P3_U4979);
  nand ginst27160 (P3_U4985, P3_U2489, P3_U4984);
  nand ginst27161 (P3_U4986, P3_U2445, P3_U4975);
  nand ginst27162 (P3_U4987, P3_U2436, P3_U2502);
  nand ginst27163 (P3_U4988, P3_U2435, P3_U4974);
  nand ginst27164 (P3_U4989, P3_U2372, P3_U2420);
  nand ginst27165 (P3_U4990, P3_INSTQUEUE_REG_9__7__SCAN_IN, P3_U4983);
  nand ginst27166 (P3_U4991, P3_U2443, P3_U4975);
  nand ginst27167 (P3_U4992, P3_U2434, P3_U2502);
  nand ginst27168 (P3_U4993, P3_U2433, P3_U4974);
  nand ginst27169 (P3_U4994, P3_U2372, P3_U2419);
  nand ginst27170 (P3_U4995, P3_INSTQUEUE_REG_9__6__SCAN_IN, P3_U4983);
  nand ginst27171 (P3_U4996, P3_U2442, P3_U4975);
  nand ginst27172 (P3_U4997, P3_U2432, P3_U2502);
  nand ginst27173 (P3_U4998, P3_U2431, P3_U4974);
  nand ginst27174 (P3_U4999, P3_U2372, P3_U2418);
  nand ginst27175 (P3_U5000, P3_INSTQUEUE_REG_9__5__SCAN_IN, P3_U4983);
  nand ginst27176 (P3_U5001, P3_U2441, P3_U4975);
  nand ginst27177 (P3_U5002, P3_U2430, P3_U2502);
  nand ginst27178 (P3_U5003, P3_U2429, P3_U4974);
  nand ginst27179 (P3_U5004, P3_U2372, P3_U2417);
  nand ginst27180 (P3_U5005, P3_INSTQUEUE_REG_9__4__SCAN_IN, P3_U4983);
  nand ginst27181 (P3_U5006, P3_U2440, P3_U4975);
  nand ginst27182 (P3_U5007, P3_U2428, P3_U2502);
  nand ginst27183 (P3_U5008, P3_U2427, P3_U4974);
  nand ginst27184 (P3_U5009, P3_U2372, P3_U2416);
  nand ginst27185 (P3_U5010, P3_INSTQUEUE_REG_9__3__SCAN_IN, P3_U4983);
  nand ginst27186 (P3_U5011, P3_U2439, P3_U4975);
  nand ginst27187 (P3_U5012, P3_U2426, P3_U2502);
  nand ginst27188 (P3_U5013, P3_U2425, P3_U4974);
  nand ginst27189 (P3_U5014, P3_U2372, P3_U2415);
  nand ginst27190 (P3_U5015, P3_INSTQUEUE_REG_9__2__SCAN_IN, P3_U4983);
  nand ginst27191 (P3_U5016, P3_U2438, P3_U4975);
  nand ginst27192 (P3_U5017, P3_U2424, P3_U2502);
  nand ginst27193 (P3_U5018, P3_U2423, P3_U4974);
  nand ginst27194 (P3_U5019, P3_U2372, P3_U2414);
  nand ginst27195 (P3_U5020, P3_INSTQUEUE_REG_9__1__SCAN_IN, P3_U4983);
  nand ginst27196 (P3_U5021, P3_U2437, P3_U4975);
  nand ginst27197 (P3_U5022, P3_U2422, P3_U2502);
  nand ginst27198 (P3_U5023, P3_U2421, P3_U4974);
  nand ginst27199 (P3_U5024, P3_U2372, P3_U2413);
  nand ginst27200 (P3_U5025, P3_INSTQUEUE_REG_9__0__SCAN_IN, P3_U4983);
  not ginst27201 (P3_U5026, P3_U3178);
  not ginst27202 (P3_U5027, P3_U3177);
  not ginst27203 (P3_U5028, P3_U3071);
  nand ginst27204 (P3_U5029, P3_U2496, P3_U4658);
  not ginst27205 (P3_U5030, P3_U3179);
  nand ginst27206 (P3_U5031, P3_U2489, P3_U3179);
  nand ginst27207 (P3_U5032, P3_U3071, P3_U5031);
  nand ginst27208 (P3_U5033, P3_STATE2_REG_3__SCAN_IN, P3_U3177);
  nand ginst27209 (P3_U5034, P3_U3493, P3_U5032);
  nand ginst27210 (P3_U5035, P3_U4322, P3_U5030);
  nand ginst27211 (P3_U5036, P3_U2489, P3_U5035);
  nand ginst27212 (P3_U5037, P3_U2445, P3_U5027);
  nand ginst27213 (P3_U5038, P3_U2436, P3_U2503);
  nand ginst27214 (P3_U5039, P3_U2435, P3_U5026);
  nand ginst27215 (P3_U5040, P3_U2371, P3_U2420);
  nand ginst27216 (P3_U5041, P3_INSTQUEUE_REG_8__7__SCAN_IN, P3_U5034);
  nand ginst27217 (P3_U5042, P3_U2443, P3_U5027);
  nand ginst27218 (P3_U5043, P3_U2434, P3_U2503);
  nand ginst27219 (P3_U5044, P3_U2433, P3_U5026);
  nand ginst27220 (P3_U5045, P3_U2371, P3_U2419);
  nand ginst27221 (P3_U5046, P3_INSTQUEUE_REG_8__6__SCAN_IN, P3_U5034);
  nand ginst27222 (P3_U5047, P3_U2442, P3_U5027);
  nand ginst27223 (P3_U5048, P3_U2432, P3_U2503);
  nand ginst27224 (P3_U5049, P3_U2431, P3_U5026);
  nand ginst27225 (P3_U5050, P3_U2371, P3_U2418);
  nand ginst27226 (P3_U5051, P3_INSTQUEUE_REG_8__5__SCAN_IN, P3_U5034);
  nand ginst27227 (P3_U5052, P3_U2441, P3_U5027);
  nand ginst27228 (P3_U5053, P3_U2430, P3_U2503);
  nand ginst27229 (P3_U5054, P3_U2429, P3_U5026);
  nand ginst27230 (P3_U5055, P3_U2371, P3_U2417);
  nand ginst27231 (P3_U5056, P3_INSTQUEUE_REG_8__4__SCAN_IN, P3_U5034);
  nand ginst27232 (P3_U5057, P3_U2440, P3_U5027);
  nand ginst27233 (P3_U5058, P3_U2428, P3_U2503);
  nand ginst27234 (P3_U5059, P3_U2427, P3_U5026);
  nand ginst27235 (P3_U5060, P3_U2371, P3_U2416);
  nand ginst27236 (P3_U5061, P3_INSTQUEUE_REG_8__3__SCAN_IN, P3_U5034);
  nand ginst27237 (P3_U5062, P3_U2439, P3_U5027);
  nand ginst27238 (P3_U5063, P3_U2426, P3_U2503);
  nand ginst27239 (P3_U5064, P3_U2425, P3_U5026);
  nand ginst27240 (P3_U5065, P3_U2371, P3_U2415);
  nand ginst27241 (P3_U5066, P3_INSTQUEUE_REG_8__2__SCAN_IN, P3_U5034);
  nand ginst27242 (P3_U5067, P3_U2438, P3_U5027);
  nand ginst27243 (P3_U5068, P3_U2424, P3_U2503);
  nand ginst27244 (P3_U5069, P3_U2423, P3_U5026);
  nand ginst27245 (P3_U5070, P3_U2371, P3_U2414);
  nand ginst27246 (P3_U5071, P3_INSTQUEUE_REG_8__1__SCAN_IN, P3_U5034);
  nand ginst27247 (P3_U5072, P3_U2437, P3_U5027);
  nand ginst27248 (P3_U5073, P3_U2422, P3_U2503);
  nand ginst27249 (P3_U5074, P3_U2421, P3_U5026);
  nand ginst27250 (P3_U5075, P3_U2371, P3_U2413);
  nand ginst27251 (P3_U5076, P3_INSTQUEUE_REG_8__0__SCAN_IN, P3_U5034);
  not ginst27252 (P3_U5077, P3_U3183);
  not ginst27253 (P3_U5078, P3_U3185);
  not ginst27254 (P3_U5079, P3_U3184);
  nand ginst27255 (P3_U5080, P3_U2489, P3_U3184);
  nand ginst27256 (P3_U5081, P3_U5078, P3_U5080);
  nand ginst27257 (P3_U5082, P3_STATE2_REG_3__SCAN_IN, P3_U3180);
  nand ginst27258 (P3_U5083, P3_U3510, P3_U5081);
  nand ginst27259 (P3_U5084, P3_U4322, P3_U5079);
  nand ginst27260 (P3_U5085, P3_U2489, P3_U5084);
  nand ginst27261 (P3_U5086, P3_U2445, P3_U4650);
  nand ginst27262 (P3_U5087, P3_U2436, P3_U4326);
  nand ginst27263 (P3_U5088, P3_U2435, P3_U5077);
  nand ginst27264 (P3_U5089, P3_U2370, P3_U2420);
  nand ginst27265 (P3_U5090, P3_INSTQUEUE_REG_7__7__SCAN_IN, P3_U5083);
  nand ginst27266 (P3_U5091, P3_U2443, P3_U4650);
  nand ginst27267 (P3_U5092, P3_U2434, P3_U4326);
  nand ginst27268 (P3_U5093, P3_U2433, P3_U5077);
  nand ginst27269 (P3_U5094, P3_U2370, P3_U2419);
  nand ginst27270 (P3_U5095, P3_INSTQUEUE_REG_7__6__SCAN_IN, P3_U5083);
  nand ginst27271 (P3_U5096, P3_U2442, P3_U4650);
  nand ginst27272 (P3_U5097, P3_U2432, P3_U4326);
  nand ginst27273 (P3_U5098, P3_U2431, P3_U5077);
  nand ginst27274 (P3_U5099, P3_U2370, P3_U2418);
  nand ginst27275 (P3_U5100, P3_INSTQUEUE_REG_7__5__SCAN_IN, P3_U5083);
  nand ginst27276 (P3_U5101, P3_U2441, P3_U4650);
  nand ginst27277 (P3_U5102, P3_U2430, P3_U4326);
  nand ginst27278 (P3_U5103, P3_U2429, P3_U5077);
  nand ginst27279 (P3_U5104, P3_U2370, P3_U2417);
  nand ginst27280 (P3_U5105, P3_INSTQUEUE_REG_7__4__SCAN_IN, P3_U5083);
  nand ginst27281 (P3_U5106, P3_U2440, P3_U4650);
  nand ginst27282 (P3_U5107, P3_U2428, P3_U4326);
  nand ginst27283 (P3_U5108, P3_U2427, P3_U5077);
  nand ginst27284 (P3_U5109, P3_U2370, P3_U2416);
  nand ginst27285 (P3_U5110, P3_INSTQUEUE_REG_7__3__SCAN_IN, P3_U5083);
  nand ginst27286 (P3_U5111, P3_U2439, P3_U4650);
  nand ginst27287 (P3_U5112, P3_U2426, P3_U4326);
  nand ginst27288 (P3_U5113, P3_U2425, P3_U5077);
  nand ginst27289 (P3_U5114, P3_U2370, P3_U2415);
  nand ginst27290 (P3_U5115, P3_INSTQUEUE_REG_7__2__SCAN_IN, P3_U5083);
  nand ginst27291 (P3_U5116, P3_U2438, P3_U4650);
  nand ginst27292 (P3_U5117, P3_U2424, P3_U4326);
  nand ginst27293 (P3_U5118, P3_U2423, P3_U5077);
  nand ginst27294 (P3_U5119, P3_U2370, P3_U2414);
  nand ginst27295 (P3_U5120, P3_INSTQUEUE_REG_7__1__SCAN_IN, P3_U5083);
  nand ginst27296 (P3_U5121, P3_U2437, P3_U4650);
  nand ginst27297 (P3_U5122, P3_U2422, P3_U4326);
  nand ginst27298 (P3_U5123, P3_U2421, P3_U5077);
  nand ginst27299 (P3_U5124, P3_U2370, P3_U2413);
  nand ginst27300 (P3_U5125, P3_INSTQUEUE_REG_7__0__SCAN_IN, P3_U5083);
  not ginst27301 (P3_U5126, P3_U3187);
  not ginst27302 (P3_U5127, P3_U3186);
  nand ginst27303 (P3_U5128, P3_U2458, P3_U4342);
  not ginst27304 (P3_U5129, P3_U3189);
  nand ginst27305 (P3_U5130, P3_U2485, P3_U4644);
  not ginst27306 (P3_U5131, P3_U3188);
  nand ginst27307 (P3_U5132, P3_U2489, P3_U3188);
  nand ginst27308 (P3_U5133, P3_U5129, P3_U5132);
  nand ginst27309 (P3_U5134, P3_STATE2_REG_3__SCAN_IN, P3_U3186);
  nand ginst27310 (P3_U5135, P3_U3528, P3_U5133);
  nand ginst27311 (P3_U5136, P3_U4322, P3_U5131);
  nand ginst27312 (P3_U5137, P3_U2489, P3_U5136);
  nand ginst27313 (P3_U5138, P3_U2445, P3_U5127);
  nand ginst27314 (P3_U5139, P3_U2436, P3_U2505);
  nand ginst27315 (P3_U5140, P3_U2435, P3_U5126);
  nand ginst27316 (P3_U5141, P3_U2369, P3_U2420);
  nand ginst27317 (P3_U5142, P3_INSTQUEUE_REG_6__7__SCAN_IN, P3_U5135);
  nand ginst27318 (P3_U5143, P3_U2443, P3_U5127);
  nand ginst27319 (P3_U5144, P3_U2434, P3_U2505);
  nand ginst27320 (P3_U5145, P3_U2433, P3_U5126);
  nand ginst27321 (P3_U5146, P3_U2369, P3_U2419);
  nand ginst27322 (P3_U5147, P3_INSTQUEUE_REG_6__6__SCAN_IN, P3_U5135);
  nand ginst27323 (P3_U5148, P3_U2442, P3_U5127);
  nand ginst27324 (P3_U5149, P3_U2432, P3_U2505);
  nand ginst27325 (P3_U5150, P3_U2431, P3_U5126);
  nand ginst27326 (P3_U5151, P3_U2369, P3_U2418);
  nand ginst27327 (P3_U5152, P3_INSTQUEUE_REG_6__5__SCAN_IN, P3_U5135);
  nand ginst27328 (P3_U5153, P3_U2441, P3_U5127);
  nand ginst27329 (P3_U5154, P3_U2430, P3_U2505);
  nand ginst27330 (P3_U5155, P3_U2429, P3_U5126);
  nand ginst27331 (P3_U5156, P3_U2369, P3_U2417);
  nand ginst27332 (P3_U5157, P3_INSTQUEUE_REG_6__4__SCAN_IN, P3_U5135);
  nand ginst27333 (P3_U5158, P3_U2440, P3_U5127);
  nand ginst27334 (P3_U5159, P3_U2428, P3_U2505);
  nand ginst27335 (P3_U5160, P3_U2427, P3_U5126);
  nand ginst27336 (P3_U5161, P3_U2369, P3_U2416);
  nand ginst27337 (P3_U5162, P3_INSTQUEUE_REG_6__3__SCAN_IN, P3_U5135);
  nand ginst27338 (P3_U5163, P3_U2439, P3_U5127);
  nand ginst27339 (P3_U5164, P3_U2426, P3_U2505);
  nand ginst27340 (P3_U5165, P3_U2425, P3_U5126);
  nand ginst27341 (P3_U5166, P3_U2369, P3_U2415);
  nand ginst27342 (P3_U5167, P3_INSTQUEUE_REG_6__2__SCAN_IN, P3_U5135);
  nand ginst27343 (P3_U5168, P3_U2438, P3_U5127);
  nand ginst27344 (P3_U5169, P3_U2424, P3_U2505);
  nand ginst27345 (P3_U5170, P3_U2423, P3_U5126);
  nand ginst27346 (P3_U5171, P3_U2369, P3_U2414);
  nand ginst27347 (P3_U5172, P3_INSTQUEUE_REG_6__1__SCAN_IN, P3_U5135);
  nand ginst27348 (P3_U5173, P3_U2437, P3_U5127);
  nand ginst27349 (P3_U5174, P3_U2422, P3_U2505);
  nand ginst27350 (P3_U5175, P3_U2421, P3_U5126);
  nand ginst27351 (P3_U5176, P3_U2369, P3_U2413);
  nand ginst27352 (P3_U5177, P3_INSTQUEUE_REG_6__0__SCAN_IN, P3_U5135);
  not ginst27353 (P3_U5178, P3_U3191);
  not ginst27354 (P3_U5179, P3_U3190);
  nand ginst27355 (P3_U5180, P3_U2458, P3_U4343);
  not ginst27356 (P3_U5181, P3_U3193);
  nand ginst27357 (P3_U5182, P3_U2485, P3_U4645);
  not ginst27358 (P3_U5183, P3_U3192);
  nand ginst27359 (P3_U5184, P3_U2489, P3_U3192);
  nand ginst27360 (P3_U5185, P3_U5181, P3_U5184);
  nand ginst27361 (P3_U5186, P3_STATE2_REG_3__SCAN_IN, P3_U3190);
  nand ginst27362 (P3_U5187, P3_U3546, P3_U5185);
  nand ginst27363 (P3_U5188, P3_U4322, P3_U5183);
  nand ginst27364 (P3_U5189, P3_U2489, P3_U5188);
  nand ginst27365 (P3_U5190, P3_U2445, P3_U5179);
  nand ginst27366 (P3_U5191, P3_U2436, P3_U2506);
  nand ginst27367 (P3_U5192, P3_U2435, P3_U5178);
  nand ginst27368 (P3_U5193, P3_U2368, P3_U2420);
  nand ginst27369 (P3_U5194, P3_INSTQUEUE_REG_5__7__SCAN_IN, P3_U5187);
  nand ginst27370 (P3_U5195, P3_U2443, P3_U5179);
  nand ginst27371 (P3_U5196, P3_U2434, P3_U2506);
  nand ginst27372 (P3_U5197, P3_U2433, P3_U5178);
  nand ginst27373 (P3_U5198, P3_U2368, P3_U2419);
  nand ginst27374 (P3_U5199, P3_INSTQUEUE_REG_5__6__SCAN_IN, P3_U5187);
  nand ginst27375 (P3_U5200, P3_U2442, P3_U5179);
  nand ginst27376 (P3_U5201, P3_U2432, P3_U2506);
  nand ginst27377 (P3_U5202, P3_U2431, P3_U5178);
  nand ginst27378 (P3_U5203, P3_U2368, P3_U2418);
  nand ginst27379 (P3_U5204, P3_INSTQUEUE_REG_5__5__SCAN_IN, P3_U5187);
  nand ginst27380 (P3_U5205, P3_U2441, P3_U5179);
  nand ginst27381 (P3_U5206, P3_U2430, P3_U2506);
  nand ginst27382 (P3_U5207, P3_U2429, P3_U5178);
  nand ginst27383 (P3_U5208, P3_U2368, P3_U2417);
  nand ginst27384 (P3_U5209, P3_INSTQUEUE_REG_5__4__SCAN_IN, P3_U5187);
  nand ginst27385 (P3_U5210, P3_U2440, P3_U5179);
  nand ginst27386 (P3_U5211, P3_U2428, P3_U2506);
  nand ginst27387 (P3_U5212, P3_U2427, P3_U5178);
  nand ginst27388 (P3_U5213, P3_U2368, P3_U2416);
  nand ginst27389 (P3_U5214, P3_INSTQUEUE_REG_5__3__SCAN_IN, P3_U5187);
  nand ginst27390 (P3_U5215, P3_U2439, P3_U5179);
  nand ginst27391 (P3_U5216, P3_U2426, P3_U2506);
  nand ginst27392 (P3_U5217, P3_U2425, P3_U5178);
  nand ginst27393 (P3_U5218, P3_U2368, P3_U2415);
  nand ginst27394 (P3_U5219, P3_INSTQUEUE_REG_5__2__SCAN_IN, P3_U5187);
  nand ginst27395 (P3_U5220, P3_U2438, P3_U5179);
  nand ginst27396 (P3_U5221, P3_U2424, P3_U2506);
  nand ginst27397 (P3_U5222, P3_U2423, P3_U5178);
  nand ginst27398 (P3_U5223, P3_U2368, P3_U2414);
  nand ginst27399 (P3_U5224, P3_INSTQUEUE_REG_5__1__SCAN_IN, P3_U5187);
  nand ginst27400 (P3_U5225, P3_U2437, P3_U5179);
  nand ginst27401 (P3_U5226, P3_U2422, P3_U2506);
  nand ginst27402 (P3_U5227, P3_U2421, P3_U5178);
  nand ginst27403 (P3_U5228, P3_U2368, P3_U2413);
  nand ginst27404 (P3_U5229, P3_INSTQUEUE_REG_5__0__SCAN_IN, P3_U5187);
  not ginst27405 (P3_U5230, P3_U3195);
  not ginst27406 (P3_U5231, P3_U3194);
  not ginst27407 (P3_U5232, P3_U3072);
  nand ginst27408 (P3_U5233, P3_U2485, P3_U2496);
  nand ginst27409 (P3_U5234, P3_U3195, P3_U5233);
  nand ginst27410 (P3_U5235, P3_U2489, P3_U5234);
  nand ginst27411 (P3_U5236, P3_U3072, P3_U5235);
  nand ginst27412 (P3_U5237, P3_STATE2_REG_3__SCAN_IN, P3_U3194);
  nand ginst27413 (P3_U5238, P3_U3564, P3_U5236);
  nand ginst27414 (P3_U5239, P3_U2489, P3_U3136);
  nand ginst27415 (P3_U5240, P3_U2445, P3_U5231);
  nand ginst27416 (P3_U5241, P3_U2436, P3_U2507);
  nand ginst27417 (P3_U5242, P3_U2435, P3_U5230);
  nand ginst27418 (P3_U5243, P3_U2367, P3_U2420);
  nand ginst27419 (P3_U5244, P3_INSTQUEUE_REG_4__7__SCAN_IN, P3_U5238);
  nand ginst27420 (P3_U5245, P3_U2443, P3_U5231);
  nand ginst27421 (P3_U5246, P3_U2434, P3_U2507);
  nand ginst27422 (P3_U5247, P3_U2433, P3_U5230);
  nand ginst27423 (P3_U5248, P3_U2367, P3_U2419);
  nand ginst27424 (P3_U5249, P3_INSTQUEUE_REG_4__6__SCAN_IN, P3_U5238);
  nand ginst27425 (P3_U5250, P3_U2442, P3_U5231);
  nand ginst27426 (P3_U5251, P3_U2432, P3_U2507);
  nand ginst27427 (P3_U5252, P3_U2431, P3_U5230);
  nand ginst27428 (P3_U5253, P3_U2367, P3_U2418);
  nand ginst27429 (P3_U5254, P3_INSTQUEUE_REG_4__5__SCAN_IN, P3_U5238);
  nand ginst27430 (P3_U5255, P3_U2441, P3_U5231);
  nand ginst27431 (P3_U5256, P3_U2430, P3_U2507);
  nand ginst27432 (P3_U5257, P3_U2429, P3_U5230);
  nand ginst27433 (P3_U5258, P3_U2367, P3_U2417);
  nand ginst27434 (P3_U5259, P3_INSTQUEUE_REG_4__4__SCAN_IN, P3_U5238);
  nand ginst27435 (P3_U5260, P3_U2440, P3_U5231);
  nand ginst27436 (P3_U5261, P3_U2428, P3_U2507);
  nand ginst27437 (P3_U5262, P3_U2427, P3_U5230);
  nand ginst27438 (P3_U5263, P3_U2367, P3_U2416);
  nand ginst27439 (P3_U5264, P3_INSTQUEUE_REG_4__3__SCAN_IN, P3_U5238);
  nand ginst27440 (P3_U5265, P3_U2439, P3_U5231);
  nand ginst27441 (P3_U5266, P3_U2426, P3_U2507);
  nand ginst27442 (P3_U5267, P3_U2425, P3_U5230);
  nand ginst27443 (P3_U5268, P3_U2367, P3_U2415);
  nand ginst27444 (P3_U5269, P3_INSTQUEUE_REG_4__2__SCAN_IN, P3_U5238);
  nand ginst27445 (P3_U5270, P3_U2438, P3_U5231);
  nand ginst27446 (P3_U5271, P3_U2424, P3_U2507);
  nand ginst27447 (P3_U5272, P3_U2423, P3_U5230);
  nand ginst27448 (P3_U5273, P3_U2367, P3_U2414);
  nand ginst27449 (P3_U5274, P3_INSTQUEUE_REG_4__1__SCAN_IN, P3_U5238);
  nand ginst27450 (P3_U5275, P3_U2437, P3_U5231);
  nand ginst27451 (P3_U5276, P3_U2422, P3_U2507);
  nand ginst27452 (P3_U5277, P3_U2421, P3_U5230);
  nand ginst27453 (P3_U5278, P3_U2367, P3_U2413);
  nand ginst27454 (P3_U5279, P3_INSTQUEUE_REG_4__0__SCAN_IN, P3_U5238);
  not ginst27455 (P3_U5280, P3_U3197);
  not ginst27456 (P3_U5281, P3_U3196);
  nand ginst27457 (P3_U5282, P3_U2460, P3_U4653);
  not ginst27458 (P3_U5283, P3_U3198);
  nand ginst27459 (P3_U5284, P3_U2509, P3_U4657);
  nand ginst27460 (P3_U5285, P3_U3197, P3_U5284);
  nand ginst27461 (P3_U5286, P3_U2489, P3_U5285);
  nand ginst27462 (P3_U5287, P3_U5283, P3_U5286);
  nand ginst27463 (P3_U5288, P3_STATE2_REG_3__SCAN_IN, P3_U3196);
  nand ginst27464 (P3_U5289, P3_U3582, P3_U5287);
  nand ginst27465 (P3_U5290, P3_U2489, P3_U3136);
  nand ginst27466 (P3_U5291, P3_U2445, P3_U5281);
  nand ginst27467 (P3_U5292, P3_U2436, P3_U2510);
  nand ginst27468 (P3_U5293, P3_U2435, P3_U5280);
  nand ginst27469 (P3_U5294, P3_U2366, P3_U2420);
  nand ginst27470 (P3_U5295, P3_INSTQUEUE_REG_3__7__SCAN_IN, P3_U5289);
  nand ginst27471 (P3_U5296, P3_U2443, P3_U5281);
  nand ginst27472 (P3_U5297, P3_U2434, P3_U2510);
  nand ginst27473 (P3_U5298, P3_U2433, P3_U5280);
  nand ginst27474 (P3_U5299, P3_U2366, P3_U2419);
  nand ginst27475 (P3_U5300, P3_INSTQUEUE_REG_3__6__SCAN_IN, P3_U5289);
  nand ginst27476 (P3_U5301, P3_U2442, P3_U5281);
  nand ginst27477 (P3_U5302, P3_U2432, P3_U2510);
  nand ginst27478 (P3_U5303, P3_U2431, P3_U5280);
  nand ginst27479 (P3_U5304, P3_U2366, P3_U2418);
  nand ginst27480 (P3_U5305, P3_INSTQUEUE_REG_3__5__SCAN_IN, P3_U5289);
  nand ginst27481 (P3_U5306, P3_U2441, P3_U5281);
  nand ginst27482 (P3_U5307, P3_U2430, P3_U2510);
  nand ginst27483 (P3_U5308, P3_U2429, P3_U5280);
  nand ginst27484 (P3_U5309, P3_U2366, P3_U2417);
  nand ginst27485 (P3_U5310, P3_INSTQUEUE_REG_3__4__SCAN_IN, P3_U5289);
  nand ginst27486 (P3_U5311, P3_U2440, P3_U5281);
  nand ginst27487 (P3_U5312, P3_U2428, P3_U2510);
  nand ginst27488 (P3_U5313, P3_U2427, P3_U5280);
  nand ginst27489 (P3_U5314, P3_U2366, P3_U2416);
  nand ginst27490 (P3_U5315, P3_INSTQUEUE_REG_3__3__SCAN_IN, P3_U5289);
  nand ginst27491 (P3_U5316, P3_U2439, P3_U5281);
  nand ginst27492 (P3_U5317, P3_U2426, P3_U2510);
  nand ginst27493 (P3_U5318, P3_U2425, P3_U5280);
  nand ginst27494 (P3_U5319, P3_U2366, P3_U2415);
  nand ginst27495 (P3_U5320, P3_INSTQUEUE_REG_3__2__SCAN_IN, P3_U5289);
  nand ginst27496 (P3_U5321, P3_U2438, P3_U5281);
  nand ginst27497 (P3_U5322, P3_U2424, P3_U2510);
  nand ginst27498 (P3_U5323, P3_U2423, P3_U5280);
  nand ginst27499 (P3_U5324, P3_U2366, P3_U2414);
  nand ginst27500 (P3_U5325, P3_INSTQUEUE_REG_3__1__SCAN_IN, P3_U5289);
  nand ginst27501 (P3_U5326, P3_U2437, P3_U5281);
  nand ginst27502 (P3_U5327, P3_U2422, P3_U2510);
  nand ginst27503 (P3_U5328, P3_U2421, P3_U5280);
  nand ginst27504 (P3_U5329, P3_U2366, P3_U2413);
  nand ginst27505 (P3_U5330, P3_INSTQUEUE_REG_3__0__SCAN_IN, P3_U5289);
  not ginst27506 (P3_U5331, P3_U3200);
  not ginst27507 (P3_U5332, P3_U3199);
  nand ginst27508 (P3_U5333, P3_U2460, P3_U4342);
  not ginst27509 (P3_U5334, P3_U3201);
  nand ginst27510 (P3_U5335, P3_U2509, P3_U4644);
  nand ginst27511 (P3_U5336, P3_U3200, P3_U5335);
  nand ginst27512 (P3_U5337, P3_U2489, P3_U5336);
  nand ginst27513 (P3_U5338, P3_U5334, P3_U5337);
  nand ginst27514 (P3_U5339, P3_STATE2_REG_3__SCAN_IN, P3_U3199);
  nand ginst27515 (P3_U5340, P3_U3599, P3_U5338);
  nand ginst27516 (P3_U5341, P3_U2489, P3_U3136);
  nand ginst27517 (P3_U5342, P3_U2445, P3_U5332);
  nand ginst27518 (P3_U5343, P3_U2436, P3_U2511);
  nand ginst27519 (P3_U5344, P3_U2435, P3_U5331);
  nand ginst27520 (P3_U5345, P3_U2365, P3_U2420);
  nand ginst27521 (P3_U5346, P3_INSTQUEUE_REG_2__7__SCAN_IN, P3_U5340);
  nand ginst27522 (P3_U5347, P3_U2443, P3_U5332);
  nand ginst27523 (P3_U5348, P3_U2434, P3_U2511);
  nand ginst27524 (P3_U5349, P3_U2433, P3_U5331);
  nand ginst27525 (P3_U5350, P3_U2365, P3_U2419);
  nand ginst27526 (P3_U5351, P3_INSTQUEUE_REG_2__6__SCAN_IN, P3_U5340);
  nand ginst27527 (P3_U5352, P3_U2442, P3_U5332);
  nand ginst27528 (P3_U5353, P3_U2432, P3_U2511);
  nand ginst27529 (P3_U5354, P3_U2431, P3_U5331);
  nand ginst27530 (P3_U5355, P3_U2365, P3_U2418);
  nand ginst27531 (P3_U5356, P3_INSTQUEUE_REG_2__5__SCAN_IN, P3_U5340);
  nand ginst27532 (P3_U5357, P3_U2441, P3_U5332);
  nand ginst27533 (P3_U5358, P3_U2430, P3_U2511);
  nand ginst27534 (P3_U5359, P3_U2429, P3_U5331);
  nand ginst27535 (P3_U5360, P3_U2365, P3_U2417);
  nand ginst27536 (P3_U5361, P3_INSTQUEUE_REG_2__4__SCAN_IN, P3_U5340);
  nand ginst27537 (P3_U5362, P3_U2440, P3_U5332);
  nand ginst27538 (P3_U5363, P3_U2428, P3_U2511);
  nand ginst27539 (P3_U5364, P3_U2427, P3_U5331);
  nand ginst27540 (P3_U5365, P3_U2365, P3_U2416);
  nand ginst27541 (P3_U5366, P3_INSTQUEUE_REG_2__3__SCAN_IN, P3_U5340);
  nand ginst27542 (P3_U5367, P3_U2439, P3_U5332);
  nand ginst27543 (P3_U5368, P3_U2426, P3_U2511);
  nand ginst27544 (P3_U5369, P3_U2425, P3_U5331);
  nand ginst27545 (P3_U5370, P3_U2365, P3_U2415);
  nand ginst27546 (P3_U5371, P3_INSTQUEUE_REG_2__2__SCAN_IN, P3_U5340);
  nand ginst27547 (P3_U5372, P3_U2438, P3_U5332);
  nand ginst27548 (P3_U5373, P3_U2424, P3_U2511);
  nand ginst27549 (P3_U5374, P3_U2423, P3_U5331);
  nand ginst27550 (P3_U5375, P3_U2365, P3_U2414);
  nand ginst27551 (P3_U5376, P3_INSTQUEUE_REG_2__1__SCAN_IN, P3_U5340);
  nand ginst27552 (P3_U5377, P3_U2437, P3_U5332);
  nand ginst27553 (P3_U5378, P3_U2422, P3_U2511);
  nand ginst27554 (P3_U5379, P3_U2421, P3_U5331);
  nand ginst27555 (P3_U5380, P3_U2365, P3_U2413);
  nand ginst27556 (P3_U5381, P3_INSTQUEUE_REG_2__0__SCAN_IN, P3_U5340);
  not ginst27557 (P3_U5382, P3_U3203);
  not ginst27558 (P3_U5383, P3_U3202);
  nand ginst27559 (P3_U5384, P3_U2460, P3_U4343);
  not ginst27560 (P3_U5385, P3_U3204);
  nand ginst27561 (P3_U5386, P3_U2509, P3_U4645);
  nand ginst27562 (P3_U5387, P3_U3203, P3_U5386);
  nand ginst27563 (P3_U5388, P3_U2489, P3_U5387);
  nand ginst27564 (P3_U5389, P3_U5385, P3_U5388);
  nand ginst27565 (P3_U5390, P3_STATE2_REG_3__SCAN_IN, P3_U3202);
  nand ginst27566 (P3_U5391, P3_U3617, P3_U5389);
  nand ginst27567 (P3_U5392, P3_U2489, P3_U3136);
  nand ginst27568 (P3_U5393, P3_U2445, P3_U5383);
  nand ginst27569 (P3_U5394, P3_U2436, P3_U2512);
  nand ginst27570 (P3_U5395, P3_U2435, P3_U5382);
  nand ginst27571 (P3_U5396, P3_U2364, P3_U2420);
  nand ginst27572 (P3_U5397, P3_INSTQUEUE_REG_1__7__SCAN_IN, P3_U5391);
  nand ginst27573 (P3_U5398, P3_U2443, P3_U5383);
  nand ginst27574 (P3_U5399, P3_U2434, P3_U2512);
  nand ginst27575 (P3_U5400, P3_U2433, P3_U5382);
  nand ginst27576 (P3_U5401, P3_U2364, P3_U2419);
  nand ginst27577 (P3_U5402, P3_INSTQUEUE_REG_1__6__SCAN_IN, P3_U5391);
  nand ginst27578 (P3_U5403, P3_U2442, P3_U5383);
  nand ginst27579 (P3_U5404, P3_U2432, P3_U2512);
  nand ginst27580 (P3_U5405, P3_U2431, P3_U5382);
  nand ginst27581 (P3_U5406, P3_U2364, P3_U2418);
  nand ginst27582 (P3_U5407, P3_INSTQUEUE_REG_1__5__SCAN_IN, P3_U5391);
  nand ginst27583 (P3_U5408, P3_U2441, P3_U5383);
  nand ginst27584 (P3_U5409, P3_U2430, P3_U2512);
  nand ginst27585 (P3_U5410, P3_U2429, P3_U5382);
  nand ginst27586 (P3_U5411, P3_U2364, P3_U2417);
  nand ginst27587 (P3_U5412, P3_INSTQUEUE_REG_1__4__SCAN_IN, P3_U5391);
  nand ginst27588 (P3_U5413, P3_U2440, P3_U5383);
  nand ginst27589 (P3_U5414, P3_U2428, P3_U2512);
  nand ginst27590 (P3_U5415, P3_U2427, P3_U5382);
  nand ginst27591 (P3_U5416, P3_U2364, P3_U2416);
  nand ginst27592 (P3_U5417, P3_INSTQUEUE_REG_1__3__SCAN_IN, P3_U5391);
  nand ginst27593 (P3_U5418, P3_U2439, P3_U5383);
  nand ginst27594 (P3_U5419, P3_U2426, P3_U2512);
  nand ginst27595 (P3_U5420, P3_U2425, P3_U5382);
  nand ginst27596 (P3_U5421, P3_U2364, P3_U2415);
  nand ginst27597 (P3_U5422, P3_INSTQUEUE_REG_1__2__SCAN_IN, P3_U5391);
  nand ginst27598 (P3_U5423, P3_U2438, P3_U5383);
  nand ginst27599 (P3_U5424, P3_U2424, P3_U2512);
  nand ginst27600 (P3_U5425, P3_U2423, P3_U5382);
  nand ginst27601 (P3_U5426, P3_U2364, P3_U2414);
  nand ginst27602 (P3_U5427, P3_INSTQUEUE_REG_1__1__SCAN_IN, P3_U5391);
  nand ginst27603 (P3_U5428, P3_U2437, P3_U5383);
  nand ginst27604 (P3_U5429, P3_U2422, P3_U2512);
  nand ginst27605 (P3_U5430, P3_U2421, P3_U5382);
  nand ginst27606 (P3_U5431, P3_U2364, P3_U2413);
  nand ginst27607 (P3_U5432, P3_INSTQUEUE_REG_1__0__SCAN_IN, P3_U5391);
  not ginst27608 (P3_U5433, P3_U3206);
  not ginst27609 (P3_U5434, P3_U3205);
  not ginst27610 (P3_U5435, P3_U3073);
  nand ginst27611 (P3_U5436, P3_U2496, P3_U2509);
  nand ginst27612 (P3_U5437, P3_U3206, P3_U5436);
  nand ginst27613 (P3_U5438, P3_U2489, P3_U5437);
  nand ginst27614 (P3_U5439, P3_U3073, P3_U5438);
  nand ginst27615 (P3_U5440, P3_STATE2_REG_3__SCAN_IN, P3_U3205);
  nand ginst27616 (P3_U5441, P3_U3635, P3_U5439);
  nand ginst27617 (P3_U5442, P3_U2489, P3_U3136);
  nand ginst27618 (P3_U5443, P3_U2445, P3_U5434);
  nand ginst27619 (P3_U5444, P3_U2436, P3_U2513);
  nand ginst27620 (P3_U5445, P3_U2435, P3_U5433);
  nand ginst27621 (P3_U5446, P3_U2363, P3_U2420);
  nand ginst27622 (P3_U5447, P3_INSTQUEUE_REG_0__7__SCAN_IN, P3_U5441);
  nand ginst27623 (P3_U5448, P3_U2443, P3_U5434);
  nand ginst27624 (P3_U5449, P3_U2434, P3_U2513);
  nand ginst27625 (P3_U5450, P3_U2433, P3_U5433);
  nand ginst27626 (P3_U5451, P3_U2363, P3_U2419);
  nand ginst27627 (P3_U5452, P3_INSTQUEUE_REG_0__6__SCAN_IN, P3_U5441);
  nand ginst27628 (P3_U5453, P3_U2442, P3_U5434);
  nand ginst27629 (P3_U5454, P3_U2432, P3_U2513);
  nand ginst27630 (P3_U5455, P3_U2431, P3_U5433);
  nand ginst27631 (P3_U5456, P3_U2363, P3_U2418);
  nand ginst27632 (P3_U5457, P3_INSTQUEUE_REG_0__5__SCAN_IN, P3_U5441);
  nand ginst27633 (P3_U5458, P3_U2441, P3_U5434);
  nand ginst27634 (P3_U5459, P3_U2430, P3_U2513);
  nand ginst27635 (P3_U5460, P3_U2429, P3_U5433);
  nand ginst27636 (P3_U5461, P3_U2363, P3_U2417);
  nand ginst27637 (P3_U5462, P3_INSTQUEUE_REG_0__4__SCAN_IN, P3_U5441);
  nand ginst27638 (P3_U5463, P3_U2440, P3_U5434);
  nand ginst27639 (P3_U5464, P3_U2428, P3_U2513);
  nand ginst27640 (P3_U5465, P3_U2427, P3_U5433);
  nand ginst27641 (P3_U5466, P3_U2363, P3_U2416);
  nand ginst27642 (P3_U5467, P3_INSTQUEUE_REG_0__3__SCAN_IN, P3_U5441);
  nand ginst27643 (P3_U5468, P3_U2439, P3_U5434);
  nand ginst27644 (P3_U5469, P3_U2426, P3_U2513);
  nand ginst27645 (P3_U5470, P3_U2425, P3_U5433);
  nand ginst27646 (P3_U5471, P3_U2363, P3_U2415);
  nand ginst27647 (P3_U5472, P3_INSTQUEUE_REG_0__2__SCAN_IN, P3_U5441);
  nand ginst27648 (P3_U5473, P3_U2438, P3_U5434);
  nand ginst27649 (P3_U5474, P3_U2424, P3_U2513);
  nand ginst27650 (P3_U5475, P3_U2423, P3_U5433);
  nand ginst27651 (P3_U5476, P3_U2363, P3_U2414);
  nand ginst27652 (P3_U5477, P3_INSTQUEUE_REG_0__1__SCAN_IN, P3_U5441);
  nand ginst27653 (P3_U5478, P3_U2437, P3_U5434);
  nand ginst27654 (P3_U5479, P3_U2422, P3_U2513);
  nand ginst27655 (P3_U5480, P3_U2421, P3_U5433);
  nand ginst27656 (P3_U5481, P3_U2363, P3_U2413);
  nand ginst27657 (P3_U5482, P3_INSTQUEUE_REG_0__0__SCAN_IN, P3_U5441);
  nand ginst27658 (P3_U5483, P3_U2514, P3_U3655, P3_U4339, P3_U7917);
  not ginst27659 (P3_U5484, P3_U3209);
  nand ginst27660 (P3_U5485, P3_U3209, P3_U4296);
  nand ginst27661 (P3_U5486, P3_GTE_450_U6, P3_U4303);
  nand ginst27662 (P3_U5487, P3_GTE_504_U6, P3_U4302);
  not ginst27663 (P3_U5488, P3_U3255);
  nand ginst27664 (P3_U5489, P3_GTE_412_U6, P3_U4304);
  nand ginst27665 (P3_U5490, P3_GTE_485_U6, P3_U2356);
  not ginst27666 (P3_U5491, P3_U3254);
  nand ginst27667 (P3_U5492, P3_U2630, P3_U3254);
  nand ginst27668 (P3_U5493, P3_GTE_390_U6, P3_U2357);
  nand ginst27669 (P3_U5494, P3_U3255, P3_U4294);
  nand ginst27670 (P3_U5495, P3_GTE_401_U6, P3_U4305);
  not ginst27671 (P3_U5496, P3_U4290);
  nand ginst27672 (P3_U5497, P3_U2390, P3_U4290);
  nand ginst27673 (P3_U5498, P3_STATE2_REG_3__SCAN_IN, P3_U3121);
  not ginst27674 (P3_U5499, P3_U4283);
  nand ginst27675 (P3_U5500, P3_U3095, P3_U3097);
  nand ginst27676 (P3_U5501, P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P3_U5500);
  nand ginst27677 (P3_U5502, P3_U2481, P3_U3095);
  nand ginst27678 (P3_U5503, P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN, P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN);
  not ginst27679 (P3_U5504, P3_U3223);
  nand ginst27680 (P3_U5505, P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN, P3_U4332);
  not ginst27681 (P3_U5506, P3_U3224);
  nand ginst27682 (P3_U5507, P3_U3107, P3_U5484);
  nand ginst27683 (P3_U5508, P3_U4488, P3_U4522, P3_U4607);
  nand ginst27684 (P3_U5509, P3_U4296, P3_U5507);
  nand ginst27685 (P3_U5510, P3_U3104, P3_U7973, P3_U7974);
  nand ginst27686 (P3_U5511, P3_U4323, P3_U4344);
  nand ginst27687 (P3_U5512, P3_U3665, P3_U5509);
  nand ginst27688 (P3_U5513, P3_U4522, P3_U4607);
  nand ginst27689 (P3_U5514, P3_U3218, P3_U4607);
  nand ginst27690 (P3_U5515, P3_U3216, P3_U4556, P3_U5514);
  nand ginst27691 (P3_U5516, P3_U4505, P3_U4573);
  nand ginst27692 (P3_U5517, P3_U4488, P3_U5516);
  nand ginst27693 (P3_U5518, P3_U3103, P3_U3112, P3_U3218);
  nand ginst27694 (P3_U5519, P3_U3104, P3_U4573, P3_U4607);
  nand ginst27695 (P3_U5520, P3_U3103, P3_U4324);
  nand ginst27696 (P3_U5521, P3_U3102, P3_U5518);
  not ginst27697 (P3_U5522, P3_U3220);
  nand ginst27698 (P3_U5523, P3_U3111, P3_U3114);
  nand ginst27699 (P3_U5524, P3_U2452, P3_U3108);
  not ginst27700 (P3_U5525, P3_U3221);
  nand ginst27701 (P3_U5526, P3_U2462, P3_U3104);
  nand ginst27702 (P3_U5527, P3_U3219, P3_U3229);
  nand ginst27703 (P3_U5528, P3_U2456, P3_U5527);
  nand ginst27704 (P3_U5529, P3_U2518, P3_U3217);
  nand ginst27705 (P3_U5530, P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN, P3_U5529);
  nand ginst27706 (P3_U5531, P3_U5525, P3_U5530);
  nand ginst27707 (P3_U5532, P3_U2450, P3_U2461, P3_U5523);
  nand ginst27708 (P3_U5533, P3_U3673, P3_U7918);
  not ginst27709 (P3_U5534, P3_U3226);
  nand ginst27710 (P3_U5535, P3_U3672, P3_U5522);
  nand ginst27711 (P3_U5536, P3_U2451, P3_U3659, P3_U5523);
  nand ginst27712 (P3_U5537, P3_U3669, P3_U5531);
  nand ginst27713 (P3_U5538, P3_U3220, P3_U3670);
  nand ginst27714 (P3_U5539, P3_U5504, P3_U5535);
  nand ginst27715 (P3_U5540, P3_U3226, P3_U5506);
  nand ginst27716 (P3_U5541, P3_ADD_495_U9, P3_U2356);
  nand ginst27717 (P3_U5542, P3_U3676, P3_U5537);
  not ginst27718 (P3_U5543, P3_U3265);
  nand ginst27719 (P3_U5544, P3_U3265, P3_U4345);
  nand ginst27720 (P3_U5545, P3_U4340, P3_U5542);
  nand ginst27721 (P3_U5546, P3_U5544, P3_U5545);
  not ginst27722 (P3_U5547, P3_U3227);
  not ginst27723 (P3_U5548, P3_U3225);
  nand ginst27724 (P3_U5549, P3_U5522, P3_U5534);
  nand ginst27725 (P3_U5550, P3_U2451, P3_U5523, P3_U5548);
  nand ginst27726 (P3_U5551, P3_U5547, P3_U5549);
  nand ginst27727 (P3_U5552, P3_ADD_495_U10, P3_U2356);
  nand ginst27728 (P3_U5553, P3_U3679, P3_U7981, P3_U7982);
  nand ginst27729 (P3_U5554, P3_STATE2_REG_1__SCAN_IN, P3_U3286, P3_U3287);
  nand ginst27730 (P3_U5555, P3_U3225, P3_U4345);
  nand ginst27731 (P3_U5556, P3_U4340, P3_U5553);
  nand ginst27732 (P3_U5557, P3_U3680, P3_U5556);
  not ginst27733 (P3_U5558, P3_U3228);
  nand ginst27734 (P3_U5559, P3_U4341, P3_U4608);
  not ginst27735 (P3_U5560, P3_U3231);
  not ginst27736 (P3_U5561, P3_U3230);
  nand ginst27737 (P3_U5562, P3_U2466, P3_U3230);
  nand ginst27738 (P3_U5563, P3_U3094, P3_U5531);
  nand ginst27739 (P3_U5564, P3_U3231, P3_U5558);
  nand ginst27740 (P3_U5565, P3_ADD_495_U4, P3_U2356);
  nand ginst27741 (P3_U5566, P3_U3681, P3_U5563);
  nand ginst27742 (P3_U5567, P3_STATE2_REG_1__SCAN_IN, P3_U3286, P3_U7985);
  nand ginst27743 (P3_U5568, P3_U4345, P3_U5558);
  nand ginst27744 (P3_U5569, P3_U4340, P3_U5566);
  nand ginst27745 (P3_U5570, P3_U3683, P3_U5569);
  nand ginst27746 (P3_U5571, P3_U5560, P3_U5561);
  nand ginst27747 (P3_U5572, P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN, P3_U2356);
  nand ginst27748 (P3_U5573, P3_U5572, P3_U7993, P3_U7994);
  nand ginst27749 (P3_U5574, P3_U3093, P3_U4345);
  nand ginst27750 (P3_U5575, P3_U4340, P3_U5573);
  nand ginst27751 (P3_U5576, P3_STATE2_REG_1__SCAN_IN, P3_U7988);
  nand ginst27752 (P3_U5577, P3_U3684, P3_U5575);
  nand ginst27753 (P3_U5578, P3_STATE2_REG_0__SCAN_IN, P3_LT_589_U6, P3_U2453);
  not ginst27754 (P3_U5579, P3_U3233);
  nand ginst27755 (P3_U5580, P3_STATE2_REG_3__SCAN_IN, P3_U3132);
  nand ginst27756 (P3_U5581, P3_U3233, P3_U5580);
  nand ginst27757 (P3_U5582, P3_U3123, P3_U4315);
  nand ginst27758 (P3_U5583, P3_U3271, P3_U4647);
  nand ginst27759 (P3_U5584, P3_U3182, P3_U5583);
  nand ginst27760 (P3_U5585, P3_U3183, P3_U5584);
  nand ginst27761 (P3_U5586, P3_U4322, P3_U5585);
  nand ginst27762 (P3_U5587, P3_U3142, P3_U5582);
  nand ginst27763 (P3_U5588, P3_STATE2_REG_3__SCAN_IN, P3_U4650);
  nand ginst27764 (P3_U5589, P3_U3685, P3_U5586);
  nand ginst27765 (P3_U5590, P3_U3233, P3_U5589);
  nand ginst27766 (P3_U5591, P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN, P3_U5581);
  nand ginst27767 (P3_U5592, P3_STATE2_REG_3__SCAN_IN, P3_U3131, P3_U4648);
  nand ginst27768 (P3_U5593, P3_U4322, P3_U7999);
  nand ginst27769 (P3_U5594, P3_U3270, P3_U5582);
  nand ginst27770 (P3_U5595, P3_U3686, P3_U5593);
  nand ginst27771 (P3_U5596, P3_STATE2_REG_3__SCAN_IN, P3_U3130);
  nand ginst27772 (P3_U5597, P3_U3233, P3_U5596);
  nand ginst27773 (P3_U5598, P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN, P3_U5597);
  nand ginst27774 (P3_U5599, P3_U3233, P3_U5595);
  nand ginst27775 (P3_U5600, P3_U3156, P3_U4322);
  nand ginst27776 (P3_U5601, P3_STATE2_REG_3__SCAN_IN, P3_U3129);
  nand ginst27777 (P3_U5602, P3_U5600, P3_U5601);
  nand ginst27778 (P3_U5603, P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P3_U5602);
  nand ginst27779 (P3_U5604, P3_U2493, P3_U4322);
  nand ginst27780 (P3_U5605, P3_U3141, P3_U5582);
  nand ginst27781 (P3_U5606, P3_U5603, P3_U5604, P3_U5605);
  nand ginst27782 (P3_U5607, P3_STATE2_REG_3__SCAN_IN, P3_U3128);
  nand ginst27783 (P3_U5608, P3_U3233, P3_U5607);
  nand ginst27784 (P3_U5609, P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN, P3_U5608);
  nand ginst27785 (P3_U5610, P3_U3233, P3_U5606);
  not ginst27786 (P3_U5611, P3_U3234);
  nand ginst27787 (P3_U5612, P3_U3233, P3_U5611);
  nand ginst27788 (P3_U5613, P3_STATE2_REG_3__SCAN_IN, P3_U3128);
  nand ginst27789 (P3_U5614, P3_U4337, P3_U5613);
  nand ginst27790 (P3_U5615, P3_U3233, P3_U5614);
  nand ginst27791 (P3_U5616, P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P3_U5612);
  nand ginst27792 (P3_U5617, P3_GTE_450_U6, P3_U2463, P3_U4294);
  nand ginst27793 (P3_U5618, P3_GTE_370_U6, P3_U4344);
  nand ginst27794 (P3_U5619, P3_U5617, P3_U5618);
  nand ginst27795 (P3_U5620, P3_GTE_412_U6, P3_U2630, P3_U4590);
  nand ginst27796 (P3_U5621, P3_GTE_355_U6, P3_U3074);
  nand ginst27797 (P3_U5622, P3_U5620, P3_U5621);
  nand ginst27798 (P3_U5623, P3_GTE_390_U6, P3_U4488);
  nand ginst27799 (P3_U5624, P3_U5623, P3_U8000, P3_U8001);
  nand ginst27800 (P3_U5625, P3_GTE_401_U6, P3_U3102, P3_U3108);
  nand ginst27801 (P3_U5626, P3_GTE_504_U6, P3_U4349);
  nand ginst27802 (P3_U5627, P3_GTE_485_U6, P3_U4348);
  nand ginst27803 (P3_U5628, P3_U4539, P3_U5624);
  nand ginst27804 (P3_U5629, P3_U2515, P3_U3687, P3_U5627, P3_U5628);
  nand ginst27805 (P3_U5630, P3_U2390, P3_U5629);
  not ginst27806 (P3_U5631, P3_U3248);
  nand ginst27807 (P3_U5632, P3_ADD_360_1242_U85, P3_U2395);
  nand ginst27808 (P3_U5633, P3_SUB_357_1258_U69, P3_U2393);
  nand ginst27809 (P3_U5634, P3_ADD_558_U5, P3_U3220);
  nand ginst27810 (P3_U5635, P3_ADD_553_U5, P3_U4298);
  nand ginst27811 (P3_U5636, P3_ADD_547_U5, P3_U4299);
  nand ginst27812 (P3_U5637, P3_INSTADDRPOINTER_REG_0__SCAN_IN, P3_U4300);
  nand ginst27813 (P3_U5638, P3_INSTADDRPOINTER_REG_0__SCAN_IN, P3_U4301);
  nand ginst27814 (P3_U5639, P3_ADD_531_U5, P3_U2354);
  nand ginst27815 (P3_U5640, P3_ADD_526_U5, P3_U2355);
  nand ginst27816 (P3_U5641, P3_INSTADDRPOINTER_REG_0__SCAN_IN, P3_U4302);
  nand ginst27817 (P3_U5642, P3_INSTADDRPOINTER_REG_0__SCAN_IN, P3_U2356);
  nand ginst27818 (P3_U5643, P3_INSTADDRPOINTER_REG_0__SCAN_IN, P3_U4303);
  nand ginst27819 (P3_U5644, P3_INSTADDRPOINTER_REG_0__SCAN_IN, P3_U4304);
  nand ginst27820 (P3_U5645, P3_ADD_405_U4, P3_U4305);
  nand ginst27821 (P3_U5646, P3_ADD_394_U4, P3_U2357);
  nand ginst27822 (P3_U5647, P3_ADD_385_U5, P3_U2358);
  nand ginst27823 (P3_U5648, P3_ADD_380_U5, P3_U2359);
  nand ginst27824 (P3_U5649, P3_ADD_349_U5, P3_U4306);
  nand ginst27825 (P3_U5650, P3_ADD_344_U5, P3_U2362);
  nand ginst27826 (P3_U5651, P3_ADD_371_1212_U87, P3_U2360);
  nand ginst27827 (P3_U5652, P3_U3692, P3_U3693, P3_U3698, P3_U5634);
  nand ginst27828 (P3_U5653, P3_REIP_REG_0__SCAN_IN, P3_U2402);
  nand ginst27829 (P3_U5654, P3_U4318, P3_U5652);
  nand ginst27830 (P3_U5655, P3_INSTADDRPOINTER_REG_0__SCAN_IN, P3_U5631);
  nand ginst27831 (P3_U5656, P3_ADD_360_1242_U19, P3_U2395);
  nand ginst27832 (P3_U5657, P3_SUB_357_1258_U21, P3_U2393);
  nand ginst27833 (P3_U5658, P3_ADD_558_U85, P3_U3220);
  nand ginst27834 (P3_U5659, P3_ADD_553_U85, P3_U4298);
  nand ginst27835 (P3_U5660, P3_ADD_547_U85, P3_U4299);
  nand ginst27836 (P3_U5661, P3_ADD_541_U4, P3_U4300);
  nand ginst27837 (P3_U5662, P3_ADD_536_U4, P3_U4301);
  nand ginst27838 (P3_U5663, P3_ADD_531_U85, P3_U2354);
  nand ginst27839 (P3_U5664, P3_ADD_526_U71, P3_U2355);
  nand ginst27840 (P3_U5665, P3_ADD_515_U4, P3_U4302);
  nand ginst27841 (P3_U5666, P3_ADD_494_U4, P3_U2356);
  nand ginst27842 (P3_U5667, P3_ADD_476_U4, P3_U4303);
  nand ginst27843 (P3_U5668, P3_ADD_441_U4, P3_U4304);
  nand ginst27844 (P3_U5669, P3_ADD_405_U81, P3_U4305);
  nand ginst27845 (P3_U5670, P3_ADD_394_U81, P3_U2357);
  nand ginst27846 (P3_U5671, P3_ADD_385_U85, P3_U2358);
  nand ginst27847 (P3_U5672, P3_ADD_380_U85, P3_U2359);
  nand ginst27848 (P3_U5673, P3_ADD_349_U85, P3_U4306);
  nand ginst27849 (P3_U5674, P3_ADD_344_U85, P3_U2362);
  nand ginst27850 (P3_U5675, P3_ADD_371_1212_U20, P3_U2360);
  nand ginst27851 (P3_U5676, P3_U3699, P3_U3700, P3_U3705, P3_U5656, P3_U5658);
  nand ginst27852 (P3_U5677, P3_REIP_REG_1__SCAN_IN, P3_U2402);
  nand ginst27853 (P3_U5678, P3_U4318, P3_U5676);
  nand ginst27854 (P3_U5679, P3_INSTADDRPOINTER_REG_1__SCAN_IN, P3_U5631);
  nand ginst27855 (P3_U5680, P3_ADD_360_1242_U91, P3_U2395);
  nand ginst27856 (P3_U5681, P3_SUB_357_1258_U78, P3_U2393);
  nand ginst27857 (P3_U5682, P3_ADD_558_U74, P3_U3220);
  nand ginst27858 (P3_U5683, P3_ADD_553_U74, P3_U4298);
  nand ginst27859 (P3_U5684, P3_ADD_547_U74, P3_U4299);
  nand ginst27860 (P3_U5685, P3_ADD_541_U71, P3_U4300);
  nand ginst27861 (P3_U5686, P3_ADD_536_U71, P3_U4301);
  nand ginst27862 (P3_U5687, P3_ADD_531_U74, P3_U2354);
  nand ginst27863 (P3_U5688, P3_ADD_526_U60, P3_U2355);
  nand ginst27864 (P3_U5689, P3_ADD_515_U71, P3_U4302);
  nand ginst27865 (P3_U5690, P3_ADD_494_U71, P3_U2356);
  nand ginst27866 (P3_U5691, P3_ADD_476_U71, P3_U4303);
  nand ginst27867 (P3_U5692, P3_ADD_441_U71, P3_U4304);
  nand ginst27868 (P3_U5693, P3_ADD_405_U5, P3_U4305);
  nand ginst27869 (P3_U5694, P3_ADD_394_U5, P3_U2357);
  nand ginst27870 (P3_U5695, P3_ADD_385_U74, P3_U2358);
  nand ginst27871 (P3_U5696, P3_ADD_380_U74, P3_U2359);
  nand ginst27872 (P3_U5697, P3_ADD_349_U74, P3_U4306);
  nand ginst27873 (P3_U5698, P3_ADD_344_U74, P3_U2362);
  nand ginst27874 (P3_U5699, P3_ADD_371_1212_U93, P3_U2360);
  nand ginst27875 (P3_U5700, P3_U3706, P3_U3710, P3_U3713, P3_U5680, P3_U5682);
  nand ginst27876 (P3_U5701, P3_REIP_REG_2__SCAN_IN, P3_U2402);
  nand ginst27877 (P3_U5702, P3_U4318, P3_U5700);
  nand ginst27878 (P3_U5703, P3_INSTADDRPOINTER_REG_2__SCAN_IN, P3_U5631);
  nand ginst27879 (P3_U5704, P3_ADD_360_1242_U17, P3_U2395);
  nand ginst27880 (P3_U5705, P3_SUB_357_1258_U76, P3_U2393);
  nand ginst27881 (P3_U5706, P3_ADD_558_U71, P3_U3220);
  nand ginst27882 (P3_U5707, P3_ADD_553_U71, P3_U4298);
  nand ginst27883 (P3_U5708, P3_ADD_547_U71, P3_U4299);
  nand ginst27884 (P3_U5709, P3_ADD_541_U68, P3_U4300);
  nand ginst27885 (P3_U5710, P3_ADD_536_U68, P3_U4301);
  nand ginst27886 (P3_U5711, P3_ADD_531_U71, P3_U2354);
  nand ginst27887 (P3_U5712, P3_ADD_526_U57, P3_U2355);
  nand ginst27888 (P3_U5713, P3_ADD_515_U68, P3_U4302);
  nand ginst27889 (P3_U5714, P3_ADD_494_U68, P3_U2356);
  nand ginst27890 (P3_U5715, P3_ADD_476_U68, P3_U4303);
  nand ginst27891 (P3_U5716, P3_ADD_441_U68, P3_U4304);
  nand ginst27892 (P3_U5717, P3_ADD_405_U93, P3_U4305);
  nand ginst27893 (P3_U5718, P3_ADD_394_U93, P3_U2357);
  nand ginst27894 (P3_U5719, P3_ADD_385_U71, P3_U2358);
  nand ginst27895 (P3_U5720, P3_ADD_380_U71, P3_U2359);
  nand ginst27896 (P3_U5721, P3_ADD_349_U71, P3_U4306);
  nand ginst27897 (P3_U5722, P3_ADD_344_U71, P3_U2362);
  nand ginst27898 (P3_U5723, P3_ADD_371_1212_U18, P3_U2360);
  nand ginst27899 (P3_U5724, P3_U3714, P3_U3715, P3_U3718, P3_U3721, P3_U5706);
  nand ginst27900 (P3_U5725, P3_REIP_REG_3__SCAN_IN, P3_U2402);
  nand ginst27901 (P3_U5726, P3_U4318, P3_U5724);
  nand ginst27902 (P3_U5727, P3_INSTADDRPOINTER_REG_3__SCAN_IN, P3_U5631);
  nand ginst27903 (P3_U5728, P3_ADD_360_1242_U18, P3_U2395);
  nand ginst27904 (P3_U5729, P3_SUB_357_1258_U75, P3_U2393);
  nand ginst27905 (P3_U5730, P3_ADD_558_U70, P3_U3220);
  nand ginst27906 (P3_U5731, P3_ADD_553_U70, P3_U4298);
  nand ginst27907 (P3_U5732, P3_ADD_547_U70, P3_U4299);
  nand ginst27908 (P3_U5733, P3_ADD_541_U67, P3_U4300);
  nand ginst27909 (P3_U5734, P3_ADD_536_U67, P3_U4301);
  nand ginst27910 (P3_U5735, P3_ADD_531_U70, P3_U2354);
  nand ginst27911 (P3_U5736, P3_ADD_526_U56, P3_U2355);
  nand ginst27912 (P3_U5737, P3_ADD_515_U67, P3_U4302);
  nand ginst27913 (P3_U5738, P3_ADD_494_U67, P3_U2356);
  nand ginst27914 (P3_U5739, P3_ADD_476_U67, P3_U4303);
  nand ginst27915 (P3_U5740, P3_ADD_441_U67, P3_U4304);
  nand ginst27916 (P3_U5741, P3_ADD_405_U68, P3_U4305);
  nand ginst27917 (P3_U5742, P3_ADD_394_U68, P3_U2357);
  nand ginst27918 (P3_U5743, P3_ADD_385_U70, P3_U2358);
  nand ginst27919 (P3_U5744, P3_ADD_380_U70, P3_U2359);
  nand ginst27920 (P3_U5745, P3_ADD_349_U70, P3_U4306);
  nand ginst27921 (P3_U5746, P3_ADD_344_U70, P3_U2362);
  nand ginst27922 (P3_U5747, P3_ADD_371_1212_U91, P3_U2360);
  nand ginst27923 (P3_U5748, P3_U3722, P3_U3726, P3_U3729, P3_U5728, P3_U5730);
  nand ginst27924 (P3_U5749, P3_REIP_REG_4__SCAN_IN, P3_U2402);
  nand ginst27925 (P3_U5750, P3_U4318, P3_U5748);
  nand ginst27926 (P3_U5751, P3_INSTADDRPOINTER_REG_4__SCAN_IN, P3_U5631);
  nand ginst27927 (P3_U5752, P3_ADD_360_1242_U89, P3_U2395);
  nand ginst27928 (P3_U5753, P3_SUB_357_1258_U74, P3_U2393);
  nand ginst27929 (P3_U5754, P3_ADD_558_U69, P3_U3220);
  nand ginst27930 (P3_U5755, P3_ADD_553_U69, P3_U4298);
  nand ginst27931 (P3_U5756, P3_ADD_547_U69, P3_U4299);
  nand ginst27932 (P3_U5757, P3_ADD_541_U66, P3_U4300);
  nand ginst27933 (P3_U5758, P3_ADD_536_U66, P3_U4301);
  nand ginst27934 (P3_U5759, P3_ADD_531_U69, P3_U2354);
  nand ginst27935 (P3_U5760, P3_ADD_526_U55, P3_U2355);
  nand ginst27936 (P3_U5761, P3_ADD_515_U66, P3_U4302);
  nand ginst27937 (P3_U5762, P3_ADD_494_U66, P3_U2356);
  nand ginst27938 (P3_U5763, P3_ADD_476_U66, P3_U4303);
  nand ginst27939 (P3_U5764, P3_ADD_441_U66, P3_U4304);
  nand ginst27940 (P3_U5765, P3_ADD_405_U67, P3_U4305);
  nand ginst27941 (P3_U5766, P3_ADD_394_U67, P3_U2357);
  nand ginst27942 (P3_U5767, P3_ADD_385_U69, P3_U2358);
  nand ginst27943 (P3_U5768, P3_ADD_380_U69, P3_U2359);
  nand ginst27944 (P3_U5769, P3_ADD_349_U69, P3_U4306);
  nand ginst27945 (P3_U5770, P3_ADD_344_U69, P3_U2362);
  nand ginst27946 (P3_U5771, P3_ADD_371_1212_U19, P3_U2360);
  nand ginst27947 (P3_U5772, P3_U3730, P3_U3734, P3_U3737, P3_U5753, P3_U5754);
  nand ginst27948 (P3_U5773, P3_REIP_REG_5__SCAN_IN, P3_U2402);
  nand ginst27949 (P3_U5774, P3_U4318, P3_U5772);
  nand ginst27950 (P3_U5775, P3_INSTADDRPOINTER_REG_5__SCAN_IN, P3_U5631);
  nand ginst27951 (P3_U5776, P3_ADD_360_1242_U88, P3_U2395);
  nand ginst27952 (P3_U5777, P3_SUB_357_1258_U73, P3_U2393);
  nand ginst27953 (P3_U5778, P3_ADD_558_U68, P3_U3220);
  nand ginst27954 (P3_U5779, P3_ADD_553_U68, P3_U4298);
  nand ginst27955 (P3_U5780, P3_ADD_547_U68, P3_U4299);
  nand ginst27956 (P3_U5781, P3_ADD_541_U65, P3_U4300);
  nand ginst27957 (P3_U5782, P3_ADD_536_U65, P3_U4301);
  nand ginst27958 (P3_U5783, P3_ADD_531_U68, P3_U2354);
  nand ginst27959 (P3_U5784, P3_ADD_526_U54, P3_U2355);
  nand ginst27960 (P3_U5785, P3_ADD_515_U65, P3_U4302);
  nand ginst27961 (P3_U5786, P3_ADD_494_U65, P3_U2356);
  nand ginst27962 (P3_U5787, P3_ADD_476_U65, P3_U4303);
  nand ginst27963 (P3_U5788, P3_ADD_441_U65, P3_U4304);
  nand ginst27964 (P3_U5789, P3_ADD_405_U66, P3_U4305);
  nand ginst27965 (P3_U5790, P3_ADD_394_U66, P3_U2357);
  nand ginst27966 (P3_U5791, P3_ADD_385_U68, P3_U2358);
  nand ginst27967 (P3_U5792, P3_ADD_380_U68, P3_U2359);
  nand ginst27968 (P3_U5793, P3_ADD_349_U68, P3_U4306);
  nand ginst27969 (P3_U5794, P3_ADD_344_U68, P3_U2362);
  nand ginst27970 (P3_U5795, P3_ADD_371_1212_U90, P3_U2360);
  nand ginst27971 (P3_U5796, P3_U3738, P3_U3742, P3_U3745, P3_U5777, P3_U5778);
  nand ginst27972 (P3_U5797, P3_REIP_REG_6__SCAN_IN, P3_U2402);
  nand ginst27973 (P3_U5798, P3_U4318, P3_U5796);
  nand ginst27974 (P3_U5799, P3_INSTADDRPOINTER_REG_6__SCAN_IN, P3_U5631);
  nand ginst27975 (P3_U5800, P3_ADD_360_1242_U87, P3_U2395);
  nand ginst27976 (P3_U5801, P3_SUB_357_1258_U72, P3_U2393);
  nand ginst27977 (P3_U5802, P3_ADD_558_U67, P3_U3220);
  nand ginst27978 (P3_U5803, P3_ADD_553_U67, P3_U4298);
  nand ginst27979 (P3_U5804, P3_ADD_547_U67, P3_U4299);
  nand ginst27980 (P3_U5805, P3_ADD_541_U64, P3_U4300);
  nand ginst27981 (P3_U5806, P3_ADD_536_U64, P3_U4301);
  nand ginst27982 (P3_U5807, P3_ADD_531_U67, P3_U2354);
  nand ginst27983 (P3_U5808, P3_ADD_526_U53, P3_U2355);
  nand ginst27984 (P3_U5809, P3_ADD_515_U64, P3_U4302);
  nand ginst27985 (P3_U5810, P3_ADD_494_U64, P3_U2356);
  nand ginst27986 (P3_U5811, P3_ADD_476_U64, P3_U4303);
  nand ginst27987 (P3_U5812, P3_ADD_441_U64, P3_U4304);
  nand ginst27988 (P3_U5813, P3_ADD_405_U65, P3_U4305);
  nand ginst27989 (P3_U5814, P3_ADD_394_U65, P3_U2357);
  nand ginst27990 (P3_U5815, P3_ADD_385_U67, P3_U2358);
  nand ginst27991 (P3_U5816, P3_ADD_380_U67, P3_U2359);
  nand ginst27992 (P3_U5817, P3_ADD_349_U67, P3_U4306);
  nand ginst27993 (P3_U5818, P3_ADD_344_U67, P3_U2362);
  nand ginst27994 (P3_U5819, P3_ADD_371_1212_U89, P3_U2360);
  nand ginst27995 (P3_U5820, P3_U3746, P3_U3750, P3_U3753, P3_U5801, P3_U5802);
  nand ginst27996 (P3_U5821, P3_REIP_REG_7__SCAN_IN, P3_U2402);
  nand ginst27997 (P3_U5822, P3_U4318, P3_U5820);
  nand ginst27998 (P3_U5823, P3_INSTADDRPOINTER_REG_7__SCAN_IN, P3_U5631);
  nand ginst27999 (P3_U5824, P3_ADD_360_1242_U86, P3_U2395);
  nand ginst28000 (P3_U5825, P3_SUB_357_1258_U71, P3_U2393);
  nand ginst28001 (P3_U5826, P3_ADD_558_U66, P3_U3220);
  nand ginst28002 (P3_U5827, P3_ADD_553_U66, P3_U4298);
  nand ginst28003 (P3_U5828, P3_ADD_547_U66, P3_U4299);
  nand ginst28004 (P3_U5829, P3_ADD_541_U63, P3_U4300);
  nand ginst28005 (P3_U5830, P3_ADD_536_U63, P3_U4301);
  nand ginst28006 (P3_U5831, P3_ADD_531_U66, P3_U2354);
  nand ginst28007 (P3_U5832, P3_ADD_526_U52, P3_U2355);
  nand ginst28008 (P3_U5833, P3_ADD_515_U63, P3_U4302);
  nand ginst28009 (P3_U5834, P3_ADD_494_U63, P3_U2356);
  nand ginst28010 (P3_U5835, P3_ADD_476_U63, P3_U4303);
  nand ginst28011 (P3_U5836, P3_ADD_441_U63, P3_U4304);
  nand ginst28012 (P3_U5837, P3_ADD_405_U64, P3_U4305);
  nand ginst28013 (P3_U5838, P3_ADD_394_U64, P3_U2357);
  nand ginst28014 (P3_U5839, P3_ADD_385_U66, P3_U2358);
  nand ginst28015 (P3_U5840, P3_ADD_380_U66, P3_U2359);
  nand ginst28016 (P3_U5841, P3_ADD_349_U66, P3_U4306);
  nand ginst28017 (P3_U5842, P3_ADD_344_U66, P3_U2362);
  nand ginst28018 (P3_U5843, P3_ADD_371_1212_U88, P3_U2360);
  nand ginst28019 (P3_U5844, P3_U3754, P3_U3757, P3_U3760, P3_U5825, P3_U5826);
  nand ginst28020 (P3_U5845, P3_REIP_REG_8__SCAN_IN, P3_U2402);
  nand ginst28021 (P3_U5846, P3_U4318, P3_U5844);
  nand ginst28022 (P3_U5847, P3_INSTADDRPOINTER_REG_8__SCAN_IN, P3_U5631);
  nand ginst28023 (P3_U5848, P3_ADD_360_1242_U106, P3_U2395);
  nand ginst28024 (P3_U5849, P3_SUB_357_1258_U70, P3_U2393);
  nand ginst28025 (P3_U5850, P3_ADD_558_U65, P3_U3220);
  nand ginst28026 (P3_U5851, P3_ADD_553_U65, P3_U4298);
  nand ginst28027 (P3_U5852, P3_ADD_547_U65, P3_U4299);
  nand ginst28028 (P3_U5853, P3_ADD_541_U62, P3_U4300);
  nand ginst28029 (P3_U5854, P3_ADD_536_U62, P3_U4301);
  nand ginst28030 (P3_U5855, P3_ADD_531_U65, P3_U2354);
  nand ginst28031 (P3_U5856, P3_ADD_526_U51, P3_U2355);
  nand ginst28032 (P3_U5857, P3_ADD_515_U62, P3_U4302);
  nand ginst28033 (P3_U5858, P3_ADD_494_U62, P3_U2356);
  nand ginst28034 (P3_U5859, P3_ADD_476_U62, P3_U4303);
  nand ginst28035 (P3_U5860, P3_ADD_441_U62, P3_U4304);
  nand ginst28036 (P3_U5861, P3_ADD_405_U63, P3_U4305);
  nand ginst28037 (P3_U5862, P3_ADD_394_U63, P3_U2357);
  nand ginst28038 (P3_U5863, P3_ADD_385_U65, P3_U2358);
  nand ginst28039 (P3_U5864, P3_ADD_380_U65, P3_U2359);
  nand ginst28040 (P3_U5865, P3_ADD_349_U65, P3_U4306);
  nand ginst28041 (P3_U5866, P3_ADD_344_U65, P3_U2362);
  nand ginst28042 (P3_U5867, P3_ADD_371_1212_U109, P3_U2360);
  nand ginst28043 (P3_U5868, P3_U3761, P3_U3764, P3_U3767, P3_U5849, P3_U5850);
  nand ginst28044 (P3_U5869, P3_REIP_REG_9__SCAN_IN, P3_U2402);
  nand ginst28045 (P3_U5870, P3_U4318, P3_U5868);
  nand ginst28046 (P3_U5871, P3_INSTADDRPOINTER_REG_9__SCAN_IN, P3_U5631);
  nand ginst28047 (P3_U5872, P3_ADD_360_1242_U4, P3_U2395);
  nand ginst28048 (P3_U5873, P3_SUB_357_1258_U93, P3_U2393);
  nand ginst28049 (P3_U5874, P3_ADD_558_U95, P3_U3220);
  nand ginst28050 (P3_U5875, P3_ADD_553_U95, P3_U4298);
  nand ginst28051 (P3_U5876, P3_ADD_547_U95, P3_U4299);
  nand ginst28052 (P3_U5877, P3_ADD_541_U91, P3_U4300);
  nand ginst28053 (P3_U5878, P3_ADD_536_U91, P3_U4301);
  nand ginst28054 (P3_U5879, P3_ADD_531_U95, P3_U2354);
  nand ginst28055 (P3_U5880, P3_ADD_526_U81, P3_U2355);
  nand ginst28056 (P3_U5881, P3_ADD_515_U91, P3_U4302);
  nand ginst28057 (P3_U5882, P3_ADD_494_U91, P3_U2356);
  nand ginst28058 (P3_U5883, P3_ADD_476_U91, P3_U4303);
  nand ginst28059 (P3_U5884, P3_ADD_441_U91, P3_U4304);
  nand ginst28060 (P3_U5885, P3_ADD_405_U91, P3_U4305);
  nand ginst28061 (P3_U5886, P3_ADD_394_U91, P3_U2357);
  nand ginst28062 (P3_U5887, P3_ADD_385_U95, P3_U2358);
  nand ginst28063 (P3_U5888, P3_ADD_380_U95, P3_U2359);
  nand ginst28064 (P3_U5889, P3_ADD_349_U95, P3_U4306);
  nand ginst28065 (P3_U5890, P3_ADD_344_U95, P3_U2362);
  nand ginst28066 (P3_U5891, P3_ADD_371_1212_U5, P3_U2360);
  nand ginst28067 (P3_U5892, P3_U3768, P3_U3771, P3_U3774, P3_U5872, P3_U5874);
  nand ginst28068 (P3_U5893, P3_REIP_REG_10__SCAN_IN, P3_U2402);
  nand ginst28069 (P3_U5894, P3_U4318, P3_U5892);
  nand ginst28070 (P3_U5895, P3_INSTADDRPOINTER_REG_10__SCAN_IN, P3_U5631);
  nand ginst28071 (P3_U5896, P3_ADD_360_1242_U84, P3_U2395);
  nand ginst28072 (P3_U5897, P3_SUB_357_1258_U92, P3_U2393);
  nand ginst28073 (P3_U5898, P3_ADD_558_U94, P3_U3220);
  nand ginst28074 (P3_U5899, P3_ADD_553_U94, P3_U4298);
  nand ginst28075 (P3_U5900, P3_ADD_547_U94, P3_U4299);
  nand ginst28076 (P3_U5901, P3_ADD_541_U90, P3_U4300);
  nand ginst28077 (P3_U5902, P3_ADD_536_U90, P3_U4301);
  nand ginst28078 (P3_U5903, P3_ADD_531_U94, P3_U2354);
  nand ginst28079 (P3_U5904, P3_ADD_526_U80, P3_U2355);
  nand ginst28080 (P3_U5905, P3_ADD_515_U90, P3_U4302);
  nand ginst28081 (P3_U5906, P3_ADD_494_U90, P3_U2356);
  nand ginst28082 (P3_U5907, P3_ADD_476_U90, P3_U4303);
  nand ginst28083 (P3_U5908, P3_ADD_441_U90, P3_U4304);
  nand ginst28084 (P3_U5909, P3_ADD_405_U90, P3_U4305);
  nand ginst28085 (P3_U5910, P3_ADD_394_U90, P3_U2357);
  nand ginst28086 (P3_U5911, P3_ADD_385_U94, P3_U2358);
  nand ginst28087 (P3_U5912, P3_ADD_380_U94, P3_U2359);
  nand ginst28088 (P3_U5913, P3_ADD_349_U94, P3_U4306);
  nand ginst28089 (P3_U5914, P3_ADD_344_U94, P3_U2362);
  nand ginst28090 (P3_U5915, P3_ADD_371_1212_U86, P3_U2360);
  nand ginst28091 (P3_U5916, P3_U3775, P3_U3778, P3_U3781, P3_U5896, P3_U5898);
  nand ginst28092 (P3_U5917, P3_REIP_REG_11__SCAN_IN, P3_U2402);
  nand ginst28093 (P3_U5918, P3_U4318, P3_U5916);
  nand ginst28094 (P3_U5919, P3_INSTADDRPOINTER_REG_11__SCAN_IN, P3_U5631);
  nand ginst28095 (P3_U5920, P3_ADD_360_1242_U5, P3_U2395);
  nand ginst28096 (P3_U5921, P3_SUB_357_1258_U91, P3_U2393);
  nand ginst28097 (P3_U5922, P3_ADD_558_U93, P3_U3220);
  nand ginst28098 (P3_U5923, P3_ADD_553_U93, P3_U4298);
  nand ginst28099 (P3_U5924, P3_ADD_547_U93, P3_U4299);
  nand ginst28100 (P3_U5925, P3_ADD_541_U89, P3_U4300);
  nand ginst28101 (P3_U5926, P3_ADD_536_U89, P3_U4301);
  nand ginst28102 (P3_U5927, P3_ADD_531_U93, P3_U2354);
  nand ginst28103 (P3_U5928, P3_ADD_526_U79, P3_U2355);
  nand ginst28104 (P3_U5929, P3_ADD_515_U89, P3_U4302);
  nand ginst28105 (P3_U5930, P3_ADD_494_U89, P3_U2356);
  nand ginst28106 (P3_U5931, P3_ADD_476_U89, P3_U4303);
  nand ginst28107 (P3_U5932, P3_ADD_441_U89, P3_U4304);
  nand ginst28108 (P3_U5933, P3_ADD_405_U89, P3_U4305);
  nand ginst28109 (P3_U5934, P3_ADD_394_U89, P3_U2357);
  nand ginst28110 (P3_U5935, P3_ADD_385_U93, P3_U2358);
  nand ginst28111 (P3_U5936, P3_ADD_380_U93, P3_U2359);
  nand ginst28112 (P3_U5937, P3_ADD_349_U93, P3_U4306);
  nand ginst28113 (P3_U5938, P3_ADD_344_U93, P3_U2362);
  nand ginst28114 (P3_U5939, P3_ADD_371_1212_U6, P3_U2360);
  nand ginst28115 (P3_U5940, P3_U3782, P3_U3785, P3_U3788, P3_U5921, P3_U5922);
  nand ginst28116 (P3_U5941, P3_REIP_REG_12__SCAN_IN, P3_U2402);
  nand ginst28117 (P3_U5942, P3_U4318, P3_U5940);
  nand ginst28118 (P3_U5943, P3_INSTADDRPOINTER_REG_12__SCAN_IN, P3_U5631);
  nand ginst28119 (P3_U5944, P3_ADD_360_1242_U6, P3_U2395);
  nand ginst28120 (P3_U5945, P3_SUB_357_1258_U15, P3_U2393);
  nand ginst28121 (P3_U5946, P3_ADD_558_U92, P3_U3220);
  nand ginst28122 (P3_U5947, P3_ADD_553_U92, P3_U4298);
  nand ginst28123 (P3_U5948, P3_ADD_547_U92, P3_U4299);
  nand ginst28124 (P3_U5949, P3_ADD_541_U88, P3_U4300);
  nand ginst28125 (P3_U5950, P3_ADD_536_U88, P3_U4301);
  nand ginst28126 (P3_U5951, P3_ADD_531_U92, P3_U2354);
  nand ginst28127 (P3_U5952, P3_ADD_526_U78, P3_U2355);
  nand ginst28128 (P3_U5953, P3_ADD_515_U88, P3_U4302);
  nand ginst28129 (P3_U5954, P3_ADD_494_U88, P3_U2356);
  nand ginst28130 (P3_U5955, P3_ADD_476_U88, P3_U4303);
  nand ginst28131 (P3_U5956, P3_ADD_441_U88, P3_U4304);
  nand ginst28132 (P3_U5957, P3_ADD_405_U88, P3_U4305);
  nand ginst28133 (P3_U5958, P3_ADD_394_U88, P3_U2357);
  nand ginst28134 (P3_U5959, P3_ADD_385_U92, P3_U2358);
  nand ginst28135 (P3_U5960, P3_ADD_380_U92, P3_U2359);
  nand ginst28136 (P3_U5961, P3_ADD_349_U92, P3_U4306);
  nand ginst28137 (P3_U5962, P3_ADD_344_U92, P3_U2362);
  nand ginst28138 (P3_U5963, P3_ADD_371_1212_U7, P3_U2360);
  nand ginst28139 (P3_U5964, P3_U3789, P3_U3792, P3_U3795, P3_U5945, P3_U5946);
  nand ginst28140 (P3_U5965, P3_REIP_REG_13__SCAN_IN, P3_U2402);
  nand ginst28141 (P3_U5966, P3_U4318, P3_U5964);
  nand ginst28142 (P3_U5967, P3_INSTADDRPOINTER_REG_13__SCAN_IN, P3_U5631);
  nand ginst28143 (P3_U5968, P3_ADD_360_1242_U83, P3_U2395);
  nand ginst28144 (P3_U5969, P3_SUB_357_1258_U90, P3_U2393);
  nand ginst28145 (P3_U5970, P3_ADD_558_U91, P3_U3220);
  nand ginst28146 (P3_U5971, P3_ADD_553_U91, P3_U4298);
  nand ginst28147 (P3_U5972, P3_ADD_547_U91, P3_U4299);
  nand ginst28148 (P3_U5973, P3_ADD_541_U87, P3_U4300);
  nand ginst28149 (P3_U5974, P3_ADD_536_U87, P3_U4301);
  nand ginst28150 (P3_U5975, P3_ADD_531_U91, P3_U2354);
  nand ginst28151 (P3_U5976, P3_ADD_526_U77, P3_U2355);
  nand ginst28152 (P3_U5977, P3_ADD_515_U87, P3_U4302);
  nand ginst28153 (P3_U5978, P3_ADD_494_U87, P3_U2356);
  nand ginst28154 (P3_U5979, P3_ADD_476_U87, P3_U4303);
  nand ginst28155 (P3_U5980, P3_ADD_441_U87, P3_U4304);
  nand ginst28156 (P3_U5981, P3_ADD_405_U87, P3_U4305);
  nand ginst28157 (P3_U5982, P3_ADD_394_U87, P3_U2357);
  nand ginst28158 (P3_U5983, P3_ADD_385_U91, P3_U2358);
  nand ginst28159 (P3_U5984, P3_ADD_380_U91, P3_U2359);
  nand ginst28160 (P3_U5985, P3_ADD_349_U91, P3_U4306);
  nand ginst28161 (P3_U5986, P3_ADD_344_U91, P3_U2362);
  nand ginst28162 (P3_U5987, P3_ADD_371_1212_U85, P3_U2360);
  nand ginst28163 (P3_U5988, P3_U3799, P3_U3802);
  nand ginst28164 (P3_U5989, P3_REIP_REG_14__SCAN_IN, P3_U2402);
  nand ginst28165 (P3_U5990, P3_U4318, P3_U5988);
  nand ginst28166 (P3_U5991, P3_INSTADDRPOINTER_REG_14__SCAN_IN, P3_U5631);
  nand ginst28167 (P3_U5992, P3_ADD_360_1242_U7, P3_U2395);
  nand ginst28168 (P3_U5993, P3_SUB_357_1258_U89, P3_U2393);
  nand ginst28169 (P3_U5994, P3_ADD_558_U90, P3_U3220);
  nand ginst28170 (P3_U5995, P3_ADD_553_U90, P3_U4298);
  nand ginst28171 (P3_U5996, P3_ADD_547_U90, P3_U4299);
  nand ginst28172 (P3_U5997, P3_ADD_541_U86, P3_U4300);
  nand ginst28173 (P3_U5998, P3_ADD_536_U86, P3_U4301);
  nand ginst28174 (P3_U5999, P3_ADD_531_U90, P3_U2354);
  nand ginst28175 (P3_U6000, P3_ADD_526_U76, P3_U2355);
  nand ginst28176 (P3_U6001, P3_ADD_515_U86, P3_U4302);
  nand ginst28177 (P3_U6002, P3_ADD_494_U86, P3_U2356);
  nand ginst28178 (P3_U6003, P3_ADD_476_U86, P3_U4303);
  nand ginst28179 (P3_U6004, P3_ADD_441_U86, P3_U4304);
  nand ginst28180 (P3_U6005, P3_ADD_405_U86, P3_U4305);
  nand ginst28181 (P3_U6006, P3_ADD_394_U86, P3_U2357);
  nand ginst28182 (P3_U6007, P3_ADD_385_U90, P3_U2358);
  nand ginst28183 (P3_U6008, P3_ADD_380_U90, P3_U2359);
  nand ginst28184 (P3_U6009, P3_ADD_349_U90, P3_U4306);
  nand ginst28185 (P3_U6010, P3_ADD_344_U90, P3_U2362);
  nand ginst28186 (P3_U6011, P3_ADD_371_1212_U8, P3_U2360);
  nand ginst28187 (P3_U6012, P3_U3807, P3_U3810);
  nand ginst28188 (P3_U6013, P3_REIP_REG_15__SCAN_IN, P3_U2402);
  nand ginst28189 (P3_U6014, P3_U4318, P3_U6012);
  nand ginst28190 (P3_U6015, P3_INSTADDRPOINTER_REG_15__SCAN_IN, P3_U5631);
  nand ginst28191 (P3_U6016, P3_ADD_360_1242_U82, P3_U2395);
  nand ginst28192 (P3_U6017, P3_SUB_357_1258_U88, P3_U2393);
  nand ginst28193 (P3_U6018, P3_ADD_558_U89, P3_U3220);
  nand ginst28194 (P3_U6019, P3_ADD_553_U89, P3_U4298);
  nand ginst28195 (P3_U6020, P3_ADD_547_U89, P3_U4299);
  nand ginst28196 (P3_U6021, P3_ADD_541_U85, P3_U4300);
  nand ginst28197 (P3_U6022, P3_ADD_536_U85, P3_U4301);
  nand ginst28198 (P3_U6023, P3_ADD_531_U89, P3_U2354);
  nand ginst28199 (P3_U6024, P3_ADD_526_U75, P3_U2355);
  nand ginst28200 (P3_U6025, P3_ADD_515_U85, P3_U4302);
  nand ginst28201 (P3_U6026, P3_ADD_494_U85, P3_U2356);
  nand ginst28202 (P3_U6027, P3_ADD_476_U85, P3_U4303);
  nand ginst28203 (P3_U6028, P3_ADD_441_U85, P3_U4304);
  nand ginst28204 (P3_U6029, P3_ADD_405_U85, P3_U4305);
  nand ginst28205 (P3_U6030, P3_ADD_394_U85, P3_U2357);
  nand ginst28206 (P3_U6031, P3_ADD_385_U89, P3_U2358);
  nand ginst28207 (P3_U6032, P3_ADD_380_U89, P3_U2359);
  nand ginst28208 (P3_U6033, P3_ADD_349_U89, P3_U4306);
  nand ginst28209 (P3_U6034, P3_ADD_344_U89, P3_U2362);
  nand ginst28210 (P3_U6035, P3_ADD_371_1212_U84, P3_U2360);
  nand ginst28211 (P3_U6036, P3_U3812, P3_U3815, P3_U3818, P3_U6016, P3_U6018);
  nand ginst28212 (P3_U6037, P3_REIP_REG_16__SCAN_IN, P3_U2402);
  nand ginst28213 (P3_U6038, P3_U4318, P3_U6036);
  nand ginst28214 (P3_U6039, P3_INSTADDRPOINTER_REG_16__SCAN_IN, P3_U5631);
  nand ginst28215 (P3_U6040, P3_ADD_360_1242_U8, P3_U2395);
  nand ginst28216 (P3_U6041, P3_SUB_357_1258_U16, P3_U2393);
  nand ginst28217 (P3_U6042, P3_ADD_558_U88, P3_U3220);
  nand ginst28218 (P3_U6043, P3_ADD_553_U88, P3_U4298);
  nand ginst28219 (P3_U6044, P3_ADD_547_U88, P3_U4299);
  nand ginst28220 (P3_U6045, P3_ADD_541_U84, P3_U4300);
  nand ginst28221 (P3_U6046, P3_ADD_536_U84, P3_U4301);
  nand ginst28222 (P3_U6047, P3_ADD_531_U88, P3_U2354);
  nand ginst28223 (P3_U6048, P3_ADD_526_U74, P3_U2355);
  nand ginst28224 (P3_U6049, P3_ADD_515_U84, P3_U4302);
  nand ginst28225 (P3_U6050, P3_ADD_494_U84, P3_U2356);
  nand ginst28226 (P3_U6051, P3_ADD_476_U84, P3_U4303);
  nand ginst28227 (P3_U6052, P3_ADD_441_U84, P3_U4304);
  nand ginst28228 (P3_U6053, P3_ADD_405_U84, P3_U4305);
  nand ginst28229 (P3_U6054, P3_ADD_394_U84, P3_U2357);
  nand ginst28230 (P3_U6055, P3_ADD_385_U88, P3_U2358);
  nand ginst28231 (P3_U6056, P3_ADD_380_U88, P3_U2359);
  nand ginst28232 (P3_U6057, P3_ADD_349_U88, P3_U4306);
  nand ginst28233 (P3_U6058, P3_ADD_344_U88, P3_U2362);
  nand ginst28234 (P3_U6059, P3_ADD_371_1212_U9, P3_U2360);
  nand ginst28235 (P3_U6060, P3_U3819, P3_U3820, P3_U3824, P3_U6040, P3_U6042);
  nand ginst28236 (P3_U6061, P3_REIP_REG_17__SCAN_IN, P3_U2402);
  nand ginst28237 (P3_U6062, P3_U4318, P3_U6060);
  nand ginst28238 (P3_U6063, P3_INSTADDRPOINTER_REG_17__SCAN_IN, P3_U5631);
  nand ginst28239 (P3_U6064, P3_ADD_360_1242_U81, P3_U2395);
  nand ginst28240 (P3_U6065, P3_SUB_357_1258_U87, P3_U2393);
  nand ginst28241 (P3_U6066, P3_ADD_558_U87, P3_U3220);
  nand ginst28242 (P3_U6067, P3_ADD_553_U87, P3_U4298);
  nand ginst28243 (P3_U6068, P3_ADD_547_U87, P3_U4299);
  nand ginst28244 (P3_U6069, P3_ADD_541_U83, P3_U4300);
  nand ginst28245 (P3_U6070, P3_ADD_536_U83, P3_U4301);
  nand ginst28246 (P3_U6071, P3_ADD_531_U87, P3_U2354);
  nand ginst28247 (P3_U6072, P3_ADD_526_U73, P3_U2355);
  nand ginst28248 (P3_U6073, P3_ADD_515_U83, P3_U4302);
  nand ginst28249 (P3_U6074, P3_ADD_494_U83, P3_U2356);
  nand ginst28250 (P3_U6075, P3_ADD_476_U83, P3_U4303);
  nand ginst28251 (P3_U6076, P3_ADD_441_U83, P3_U4304);
  nand ginst28252 (P3_U6077, P3_ADD_405_U83, P3_U4305);
  nand ginst28253 (P3_U6078, P3_ADD_394_U83, P3_U2357);
  nand ginst28254 (P3_U6079, P3_ADD_385_U87, P3_U2358);
  nand ginst28255 (P3_U6080, P3_ADD_380_U87, P3_U2359);
  nand ginst28256 (P3_U6081, P3_ADD_349_U87, P3_U4306);
  nand ginst28257 (P3_U6082, P3_ADD_344_U87, P3_U2362);
  nand ginst28258 (P3_U6083, P3_ADD_371_1212_U83, P3_U2360);
  nand ginst28259 (P3_U6084, P3_U3825, P3_U3828, P3_U3831, P3_U6064, P3_U6066);
  nand ginst28260 (P3_U6085, P3_REIP_REG_18__SCAN_IN, P3_U2402);
  nand ginst28261 (P3_U6086, P3_U4318, P3_U6084);
  nand ginst28262 (P3_U6087, P3_INSTADDRPOINTER_REG_18__SCAN_IN, P3_U5631);
  nand ginst28263 (P3_U6088, P3_ADD_360_1242_U9, P3_U2395);
  nand ginst28264 (P3_U6089, P3_SUB_357_1258_U86, P3_U2393);
  nand ginst28265 (P3_U6090, P3_ADD_558_U86, P3_U3220);
  nand ginst28266 (P3_U6091, P3_ADD_553_U86, P3_U4298);
  nand ginst28267 (P3_U6092, P3_ADD_547_U86, P3_U4299);
  nand ginst28268 (P3_U6093, P3_ADD_541_U82, P3_U4300);
  nand ginst28269 (P3_U6094, P3_ADD_536_U82, P3_U4301);
  nand ginst28270 (P3_U6095, P3_ADD_531_U86, P3_U2354);
  nand ginst28271 (P3_U6096, P3_ADD_526_U72, P3_U2355);
  nand ginst28272 (P3_U6097, P3_ADD_515_U82, P3_U4302);
  nand ginst28273 (P3_U6098, P3_ADD_494_U82, P3_U2356);
  nand ginst28274 (P3_U6099, P3_ADD_476_U82, P3_U4303);
  nand ginst28275 (P3_U6100, P3_ADD_441_U82, P3_U4304);
  nand ginst28276 (P3_U6101, P3_ADD_405_U82, P3_U4305);
  nand ginst28277 (P3_U6102, P3_ADD_394_U82, P3_U2357);
  nand ginst28278 (P3_U6103, P3_ADD_385_U86, P3_U2358);
  nand ginst28279 (P3_U6104, P3_ADD_380_U86, P3_U2359);
  nand ginst28280 (P3_U6105, P3_ADD_349_U86, P3_U4306);
  nand ginst28281 (P3_U6106, P3_ADD_344_U86, P3_U2362);
  nand ginst28282 (P3_U6107, P3_ADD_371_1212_U10, P3_U2360);
  nand ginst28283 (P3_U6108, P3_U3832, P3_U3833, P3_U3837, P3_U6088, P3_U6090);
  nand ginst28284 (P3_U6109, P3_REIP_REG_19__SCAN_IN, P3_U2402);
  nand ginst28285 (P3_U6110, P3_U4318, P3_U6108);
  nand ginst28286 (P3_U6111, P3_INSTADDRPOINTER_REG_19__SCAN_IN, P3_U5631);
  nand ginst28287 (P3_U6112, P3_ADD_360_1242_U10, P3_U2395);
  nand ginst28288 (P3_U6113, P3_SUB_357_1258_U17, P3_U2393);
  nand ginst28289 (P3_U6114, P3_ADD_558_U84, P3_U3220);
  nand ginst28290 (P3_U6115, P3_ADD_553_U84, P3_U4298);
  nand ginst28291 (P3_U6116, P3_ADD_547_U84, P3_U4299);
  nand ginst28292 (P3_U6117, P3_ADD_541_U81, P3_U4300);
  nand ginst28293 (P3_U6118, P3_ADD_536_U81, P3_U4301);
  nand ginst28294 (P3_U6119, P3_ADD_531_U84, P3_U2354);
  nand ginst28295 (P3_U6120, P3_ADD_526_U70, P3_U2355);
  nand ginst28296 (P3_U6121, P3_ADD_515_U81, P3_U4302);
  nand ginst28297 (P3_U6122, P3_ADD_494_U81, P3_U2356);
  nand ginst28298 (P3_U6123, P3_ADD_476_U81, P3_U4303);
  nand ginst28299 (P3_U6124, P3_ADD_441_U81, P3_U4304);
  nand ginst28300 (P3_U6125, P3_ADD_405_U80, P3_U4305);
  nand ginst28301 (P3_U6126, P3_ADD_394_U80, P3_U2357);
  nand ginst28302 (P3_U6127, P3_ADD_385_U84, P3_U2358);
  nand ginst28303 (P3_U6128, P3_ADD_380_U84, P3_U2359);
  nand ginst28304 (P3_U6129, P3_ADD_349_U84, P3_U4306);
  nand ginst28305 (P3_U6130, P3_ADD_344_U84, P3_U2362);
  nand ginst28306 (P3_U6131, P3_ADD_371_1212_U11, P3_U2360);
  nand ginst28307 (P3_U6132, P3_U3841, P3_U6113);
  nand ginst28308 (P3_U6133, P3_REIP_REG_20__SCAN_IN, P3_U2402);
  nand ginst28309 (P3_U6134, P3_U4318, P3_U6132);
  nand ginst28310 (P3_U6135, P3_INSTADDRPOINTER_REG_20__SCAN_IN, P3_U5631);
  nand ginst28311 (P3_U6136, P3_ADD_360_1242_U11, P3_U2395);
  nand ginst28312 (P3_U6137, P3_SUB_357_1258_U85, P3_U2393);
  nand ginst28313 (P3_U6138, P3_ADD_558_U83, P3_U3220);
  nand ginst28314 (P3_U6139, P3_ADD_553_U83, P3_U4298);
  nand ginst28315 (P3_U6140, P3_ADD_547_U83, P3_U4299);
  nand ginst28316 (P3_U6141, P3_ADD_541_U80, P3_U4300);
  nand ginst28317 (P3_U6142, P3_ADD_536_U80, P3_U4301);
  nand ginst28318 (P3_U6143, P3_ADD_531_U83, P3_U2354);
  nand ginst28319 (P3_U6144, P3_ADD_526_U69, P3_U2355);
  nand ginst28320 (P3_U6145, P3_ADD_515_U80, P3_U4302);
  nand ginst28321 (P3_U6146, P3_ADD_494_U80, P3_U2356);
  nand ginst28322 (P3_U6147, P3_ADD_476_U80, P3_U4303);
  nand ginst28323 (P3_U6148, P3_ADD_441_U80, P3_U4304);
  nand ginst28324 (P3_U6149, P3_ADD_405_U79, P3_U4305);
  nand ginst28325 (P3_U6150, P3_ADD_394_U79, P3_U2357);
  nand ginst28326 (P3_U6151, P3_ADD_385_U83, P3_U2358);
  nand ginst28327 (P3_U6152, P3_ADD_380_U83, P3_U2359);
  nand ginst28328 (P3_U6153, P3_ADD_349_U83, P3_U4306);
  nand ginst28329 (P3_U6154, P3_ADD_344_U83, P3_U2362);
  nand ginst28330 (P3_U6155, P3_ADD_371_1212_U12, P3_U2360);
  nand ginst28331 (P3_U6156, P3_U3849, P3_U6137);
  nand ginst28332 (P3_U6157, P3_REIP_REG_21__SCAN_IN, P3_U2402);
  nand ginst28333 (P3_U6158, P3_U4318, P3_U6156);
  nand ginst28334 (P3_U6159, P3_INSTADDRPOINTER_REG_21__SCAN_IN, P3_U5631);
  nand ginst28335 (P3_U6160, P3_ADD_360_1242_U80, P3_U2395);
  nand ginst28336 (P3_U6161, P3_SUB_357_1258_U84, P3_U2393);
  nand ginst28337 (P3_U6162, P3_ADD_558_U82, P3_U3220);
  nand ginst28338 (P3_U6163, P3_ADD_553_U82, P3_U4298);
  nand ginst28339 (P3_U6164, P3_ADD_547_U82, P3_U4299);
  nand ginst28340 (P3_U6165, P3_ADD_541_U79, P3_U4300);
  nand ginst28341 (P3_U6166, P3_ADD_536_U79, P3_U4301);
  nand ginst28342 (P3_U6167, P3_ADD_531_U82, P3_U2354);
  nand ginst28343 (P3_U6168, P3_ADD_526_U68, P3_U2355);
  nand ginst28344 (P3_U6169, P3_ADD_515_U79, P3_U4302);
  nand ginst28345 (P3_U6170, P3_ADD_494_U79, P3_U2356);
  nand ginst28346 (P3_U6171, P3_ADD_476_U79, P3_U4303);
  nand ginst28347 (P3_U6172, P3_ADD_441_U79, P3_U4304);
  nand ginst28348 (P3_U6173, P3_ADD_405_U78, P3_U4305);
  nand ginst28349 (P3_U6174, P3_ADD_394_U78, P3_U2357);
  nand ginst28350 (P3_U6175, P3_ADD_385_U82, P3_U2358);
  nand ginst28351 (P3_U6176, P3_ADD_380_U82, P3_U2359);
  nand ginst28352 (P3_U6177, P3_ADD_349_U82, P3_U4306);
  nand ginst28353 (P3_U6178, P3_ADD_344_U82, P3_U2362);
  nand ginst28354 (P3_U6179, P3_ADD_371_1212_U82, P3_U2360);
  nand ginst28355 (P3_U6180, P3_U3857, P3_U3862);
  nand ginst28356 (P3_U6181, P3_REIP_REG_22__SCAN_IN, P3_U2402);
  nand ginst28357 (P3_U6182, P3_U4318, P3_U6180);
  nand ginst28358 (P3_U6183, P3_INSTADDRPOINTER_REG_22__SCAN_IN, P3_U5631);
  nand ginst28359 (P3_U6184, P3_ADD_360_1242_U12, P3_U2395);
  nand ginst28360 (P3_U6185, P3_SUB_357_1258_U83, P3_U2393);
  nand ginst28361 (P3_U6186, P3_ADD_558_U81, P3_U3220);
  nand ginst28362 (P3_U6187, P3_ADD_553_U81, P3_U4298);
  nand ginst28363 (P3_U6188, P3_ADD_547_U81, P3_U4299);
  nand ginst28364 (P3_U6189, P3_ADD_541_U78, P3_U4300);
  nand ginst28365 (P3_U6190, P3_ADD_536_U78, P3_U4301);
  nand ginst28366 (P3_U6191, P3_ADD_531_U81, P3_U2354);
  nand ginst28367 (P3_U6192, P3_ADD_526_U67, P3_U2355);
  nand ginst28368 (P3_U6193, P3_ADD_515_U78, P3_U4302);
  nand ginst28369 (P3_U6194, P3_ADD_494_U78, P3_U2356);
  nand ginst28370 (P3_U6195, P3_ADD_476_U78, P3_U4303);
  nand ginst28371 (P3_U6196, P3_ADD_441_U78, P3_U4304);
  nand ginst28372 (P3_U6197, P3_ADD_405_U77, P3_U4305);
  nand ginst28373 (P3_U6198, P3_ADD_394_U77, P3_U2357);
  nand ginst28374 (P3_U6199, P3_ADD_385_U81, P3_U2358);
  nand ginst28375 (P3_U6200, P3_ADD_380_U81, P3_U2359);
  nand ginst28376 (P3_U6201, P3_ADD_349_U81, P3_U4306);
  nand ginst28377 (P3_U6202, P3_ADD_344_U81, P3_U2362);
  nand ginst28378 (P3_U6203, P3_ADD_371_1212_U13, P3_U2360);
  nand ginst28379 (P3_U6204, P3_U3867, P3_U3872);
  nand ginst28380 (P3_U6205, P3_REIP_REG_23__SCAN_IN, P3_U2402);
  nand ginst28381 (P3_U6206, P3_U4318, P3_U6204);
  nand ginst28382 (P3_U6207, P3_INSTADDRPOINTER_REG_23__SCAN_IN, P3_U5631);
  nand ginst28383 (P3_U6208, P3_ADD_360_1242_U79, P3_U2395);
  nand ginst28384 (P3_U6209, P3_SUB_357_1258_U82, P3_U2393);
  nand ginst28385 (P3_U6210, P3_ADD_558_U80, P3_U3220);
  nand ginst28386 (P3_U6211, P3_ADD_553_U80, P3_U4298);
  nand ginst28387 (P3_U6212, P3_ADD_547_U80, P3_U4299);
  nand ginst28388 (P3_U6213, P3_ADD_541_U77, P3_U4300);
  nand ginst28389 (P3_U6214, P3_ADD_536_U77, P3_U4301);
  nand ginst28390 (P3_U6215, P3_ADD_531_U80, P3_U2354);
  nand ginst28391 (P3_U6216, P3_ADD_526_U66, P3_U2355);
  nand ginst28392 (P3_U6217, P3_ADD_515_U77, P3_U4302);
  nand ginst28393 (P3_U6218, P3_ADD_494_U77, P3_U2356);
  nand ginst28394 (P3_U6219, P3_ADD_476_U77, P3_U4303);
  nand ginst28395 (P3_U6220, P3_ADD_441_U77, P3_U4304);
  nand ginst28396 (P3_U6221, P3_ADD_405_U76, P3_U4305);
  nand ginst28397 (P3_U6222, P3_ADD_394_U76, P3_U2357);
  nand ginst28398 (P3_U6223, P3_ADD_385_U80, P3_U2358);
  nand ginst28399 (P3_U6224, P3_ADD_380_U80, P3_U2359);
  nand ginst28400 (P3_U6225, P3_ADD_349_U80, P3_U4306);
  nand ginst28401 (P3_U6226, P3_ADD_344_U80, P3_U2362);
  nand ginst28402 (P3_U6227, P3_ADD_371_1212_U81, P3_U2360);
  nand ginst28403 (P3_U6228, P3_U3877, P3_U3882);
  nand ginst28404 (P3_U6229, P3_REIP_REG_24__SCAN_IN, P3_U2402);
  nand ginst28405 (P3_U6230, P3_U4318, P3_U6228);
  nand ginst28406 (P3_U6231, P3_INSTADDRPOINTER_REG_24__SCAN_IN, P3_U5631);
  nand ginst28407 (P3_U6232, P3_ADD_360_1242_U13, P3_U2395);
  nand ginst28408 (P3_U6233, P3_SUB_357_1258_U81, P3_U2393);
  nand ginst28409 (P3_U6234, P3_ADD_558_U79, P3_U3220);
  nand ginst28410 (P3_U6235, P3_ADD_553_U79, P3_U4298);
  nand ginst28411 (P3_U6236, P3_ADD_547_U79, P3_U4299);
  nand ginst28412 (P3_U6237, P3_ADD_541_U76, P3_U4300);
  nand ginst28413 (P3_U6238, P3_ADD_536_U76, P3_U4301);
  nand ginst28414 (P3_U6239, P3_ADD_531_U79, P3_U2354);
  nand ginst28415 (P3_U6240, P3_ADD_526_U65, P3_U2355);
  nand ginst28416 (P3_U6241, P3_ADD_515_U76, P3_U4302);
  nand ginst28417 (P3_U6242, P3_ADD_494_U76, P3_U2356);
  nand ginst28418 (P3_U6243, P3_ADD_476_U76, P3_U4303);
  nand ginst28419 (P3_U6244, P3_ADD_441_U76, P3_U4304);
  nand ginst28420 (P3_U6245, P3_ADD_405_U75, P3_U4305);
  nand ginst28421 (P3_U6246, P3_ADD_394_U75, P3_U2357);
  nand ginst28422 (P3_U6247, P3_ADD_385_U79, P3_U2358);
  nand ginst28423 (P3_U6248, P3_ADD_380_U79, P3_U2359);
  nand ginst28424 (P3_U6249, P3_ADD_349_U79, P3_U4306);
  nand ginst28425 (P3_U6250, P3_ADD_344_U79, P3_U2362);
  nand ginst28426 (P3_U6251, P3_ADD_371_1212_U14, P3_U2360);
  nand ginst28427 (P3_U6252, P3_U3887, P3_U3892);
  nand ginst28428 (P3_U6253, P3_REIP_REG_25__SCAN_IN, P3_U2402);
  nand ginst28429 (P3_U6254, P3_U4318, P3_U6252);
  nand ginst28430 (P3_U6255, P3_INSTADDRPOINTER_REG_25__SCAN_IN, P3_U5631);
  nand ginst28431 (P3_U6256, P3_ADD_360_1242_U14, P3_U2395);
  nand ginst28432 (P3_U6257, P3_SUB_357_1258_U18, P3_U2393);
  nand ginst28433 (P3_U6258, P3_ADD_558_U78, P3_U3220);
  nand ginst28434 (P3_U6259, P3_ADD_553_U78, P3_U4298);
  nand ginst28435 (P3_U6260, P3_ADD_547_U78, P3_U4299);
  nand ginst28436 (P3_U6261, P3_ADD_541_U75, P3_U4300);
  nand ginst28437 (P3_U6262, P3_ADD_536_U75, P3_U4301);
  nand ginst28438 (P3_U6263, P3_ADD_531_U78, P3_U2354);
  nand ginst28439 (P3_U6264, P3_ADD_526_U64, P3_U2355);
  nand ginst28440 (P3_U6265, P3_ADD_515_U75, P3_U4302);
  nand ginst28441 (P3_U6266, P3_ADD_494_U75, P3_U2356);
  nand ginst28442 (P3_U6267, P3_ADD_476_U75, P3_U4303);
  nand ginst28443 (P3_U6268, P3_ADD_441_U75, P3_U4304);
  nand ginst28444 (P3_U6269, P3_ADD_405_U74, P3_U4305);
  nand ginst28445 (P3_U6270, P3_ADD_394_U74, P3_U2357);
  nand ginst28446 (P3_U6271, P3_ADD_385_U78, P3_U2358);
  nand ginst28447 (P3_U6272, P3_ADD_380_U78, P3_U2359);
  nand ginst28448 (P3_U6273, P3_ADD_349_U78, P3_U4306);
  nand ginst28449 (P3_U6274, P3_ADD_344_U78, P3_U2362);
  nand ginst28450 (P3_U6275, P3_ADD_371_1212_U15, P3_U2360);
  nand ginst28451 (P3_U6276, P3_U3894, P3_U3895, P3_U3897, P3_U3902, P3_U6258);
  nand ginst28452 (P3_U6277, P3_REIP_REG_26__SCAN_IN, P3_U2402);
  nand ginst28453 (P3_U6278, P3_U4318, P3_U6276);
  nand ginst28454 (P3_U6279, P3_INSTADDRPOINTER_REG_26__SCAN_IN, P3_U5631);
  nand ginst28455 (P3_U6280, P3_ADD_360_1242_U78, P3_U2395);
  nand ginst28456 (P3_U6281, P3_SUB_357_1258_U80, P3_U2393);
  nand ginst28457 (P3_U6282, P3_ADD_558_U77, P3_U3220);
  nand ginst28458 (P3_U6283, P3_ADD_553_U77, P3_U4298);
  nand ginst28459 (P3_U6284, P3_ADD_547_U77, P3_U4299);
  nand ginst28460 (P3_U6285, P3_ADD_541_U74, P3_U4300);
  nand ginst28461 (P3_U6286, P3_ADD_536_U74, P3_U4301);
  nand ginst28462 (P3_U6287, P3_ADD_531_U77, P3_U2354);
  nand ginst28463 (P3_U6288, P3_ADD_526_U63, P3_U2355);
  nand ginst28464 (P3_U6289, P3_ADD_515_U74, P3_U4302);
  nand ginst28465 (P3_U6290, P3_ADD_494_U74, P3_U2356);
  nand ginst28466 (P3_U6291, P3_ADD_476_U74, P3_U4303);
  nand ginst28467 (P3_U6292, P3_ADD_441_U74, P3_U4304);
  nand ginst28468 (P3_U6293, P3_ADD_405_U73, P3_U4305);
  nand ginst28469 (P3_U6294, P3_ADD_394_U73, P3_U2357);
  nand ginst28470 (P3_U6295, P3_ADD_385_U77, P3_U2358);
  nand ginst28471 (P3_U6296, P3_ADD_380_U77, P3_U2359);
  nand ginst28472 (P3_U6297, P3_ADD_349_U77, P3_U4306);
  nand ginst28473 (P3_U6298, P3_ADD_344_U77, P3_U2362);
  nand ginst28474 (P3_U6299, P3_ADD_371_1212_U80, P3_U2360);
  nand ginst28475 (P3_U6300, P3_U3903, P3_U3904, P3_U3906, P3_U3911, P3_U6282);
  nand ginst28476 (P3_U6301, P3_REIP_REG_27__SCAN_IN, P3_U2402);
  nand ginst28477 (P3_U6302, P3_U4318, P3_U6300);
  nand ginst28478 (P3_U6303, P3_INSTADDRPOINTER_REG_27__SCAN_IN, P3_U5631);
  nand ginst28479 (P3_U6304, P3_ADD_360_1242_U15, P3_U2395);
  nand ginst28480 (P3_U6305, P3_SUB_357_1258_U19, P3_U2393);
  nand ginst28481 (P3_U6306, P3_ADD_558_U76, P3_U3220);
  nand ginst28482 (P3_U6307, P3_ADD_553_U76, P3_U4298);
  nand ginst28483 (P3_U6308, P3_ADD_547_U76, P3_U4299);
  nand ginst28484 (P3_U6309, P3_ADD_541_U73, P3_U4300);
  nand ginst28485 (P3_U6310, P3_ADD_536_U73, P3_U4301);
  nand ginst28486 (P3_U6311, P3_ADD_531_U76, P3_U2354);
  nand ginst28487 (P3_U6312, P3_ADD_526_U62, P3_U2355);
  nand ginst28488 (P3_U6313, P3_ADD_515_U73, P3_U4302);
  nand ginst28489 (P3_U6314, P3_ADD_494_U73, P3_U2356);
  nand ginst28490 (P3_U6315, P3_ADD_476_U73, P3_U4303);
  nand ginst28491 (P3_U6316, P3_ADD_441_U73, P3_U4304);
  nand ginst28492 (P3_U6317, P3_ADD_405_U72, P3_U4305);
  nand ginst28493 (P3_U6318, P3_ADD_394_U72, P3_U2357);
  nand ginst28494 (P3_U6319, P3_ADD_385_U76, P3_U2358);
  nand ginst28495 (P3_U6320, P3_ADD_380_U76, P3_U2359);
  nand ginst28496 (P3_U6321, P3_ADD_349_U76, P3_U4306);
  nand ginst28497 (P3_U6322, P3_ADD_344_U76, P3_U2362);
  nand ginst28498 (P3_U6323, P3_ADD_371_1212_U16, P3_U2360);
  nand ginst28499 (P3_U6324, P3_U3912, P3_U3913, P3_U3915, P3_U3920, P3_U6306);
  nand ginst28500 (P3_U6325, P3_REIP_REG_28__SCAN_IN, P3_U2402);
  nand ginst28501 (P3_U6326, P3_U4318, P3_U6324);
  nand ginst28502 (P3_U6327, P3_INSTADDRPOINTER_REG_28__SCAN_IN, P3_U5631);
  nand ginst28503 (P3_U6328, P3_ADD_360_1242_U16, P3_U2395);
  nand ginst28504 (P3_U6329, P3_SUB_357_1258_U79, P3_U2393);
  nand ginst28505 (P3_U6330, P3_ADD_558_U75, P3_U3220);
  nand ginst28506 (P3_U6331, P3_ADD_553_U75, P3_U4298);
  nand ginst28507 (P3_U6332, P3_ADD_547_U75, P3_U4299);
  nand ginst28508 (P3_U6333, P3_ADD_541_U72, P3_U4300);
  nand ginst28509 (P3_U6334, P3_ADD_536_U72, P3_U4301);
  nand ginst28510 (P3_U6335, P3_ADD_531_U75, P3_U2354);
  nand ginst28511 (P3_U6336, P3_ADD_526_U61, P3_U2355);
  nand ginst28512 (P3_U6337, P3_ADD_515_U72, P3_U4302);
  nand ginst28513 (P3_U6338, P3_ADD_494_U72, P3_U2356);
  nand ginst28514 (P3_U6339, P3_ADD_476_U72, P3_U4303);
  nand ginst28515 (P3_U6340, P3_ADD_441_U72, P3_U4304);
  nand ginst28516 (P3_U6341, P3_ADD_405_U71, P3_U4305);
  nand ginst28517 (P3_U6342, P3_ADD_394_U71, P3_U2357);
  nand ginst28518 (P3_U6343, P3_ADD_385_U75, P3_U2358);
  nand ginst28519 (P3_U6344, P3_ADD_380_U75, P3_U2359);
  nand ginst28520 (P3_U6345, P3_ADD_349_U75, P3_U4306);
  nand ginst28521 (P3_U6346, P3_ADD_344_U75, P3_U2362);
  nand ginst28522 (P3_U6347, P3_ADD_371_1212_U17, P3_U2360);
  nand ginst28523 (P3_U6348, P3_U3921, P3_U3922, P3_U3924, P3_U3929, P3_U6330);
  nand ginst28524 (P3_U6349, P3_REIP_REG_29__SCAN_IN, P3_U2402);
  nand ginst28525 (P3_U6350, P3_U4318, P3_U6348);
  nand ginst28526 (P3_U6351, P3_INSTADDRPOINTER_REG_29__SCAN_IN, P3_U5631);
  nand ginst28527 (P3_U6352, P3_ADD_360_1242_U77, P3_U2395);
  nand ginst28528 (P3_U6353, P3_SUB_357_1258_U77, P3_U2393);
  nand ginst28529 (P3_U6354, P3_ADD_558_U73, P3_U3220);
  nand ginst28530 (P3_U6355, P3_ADD_553_U73, P3_U4298);
  nand ginst28531 (P3_U6356, P3_ADD_547_U73, P3_U4299);
  nand ginst28532 (P3_U6357, P3_ADD_541_U70, P3_U4300);
  nand ginst28533 (P3_U6358, P3_ADD_536_U70, P3_U4301);
  nand ginst28534 (P3_U6359, P3_ADD_531_U73, P3_U2354);
  nand ginst28535 (P3_U6360, P3_ADD_526_U59, P3_U2355);
  nand ginst28536 (P3_U6361, P3_ADD_515_U70, P3_U4302);
  nand ginst28537 (P3_U6362, P3_ADD_494_U70, P3_U2356);
  nand ginst28538 (P3_U6363, P3_ADD_476_U70, P3_U4303);
  nand ginst28539 (P3_U6364, P3_ADD_441_U70, P3_U4304);
  nand ginst28540 (P3_U6365, P3_ADD_405_U70, P3_U4305);
  nand ginst28541 (P3_U6366, P3_ADD_394_U70, P3_U2357);
  nand ginst28542 (P3_U6367, P3_ADD_385_U73, P3_U2358);
  nand ginst28543 (P3_U6368, P3_ADD_380_U73, P3_U2359);
  nand ginst28544 (P3_U6369, P3_ADD_349_U73, P3_U4306);
  nand ginst28545 (P3_U6370, P3_ADD_344_U73, P3_U2362);
  nand ginst28546 (P3_U6371, P3_ADD_371_1212_U79, P3_U2360);
  nand ginst28547 (P3_U6372, P3_U3930, P3_U3931, P3_U3933, P3_U3938, P3_U6354);
  nand ginst28548 (P3_U6373, P3_REIP_REG_30__SCAN_IN, P3_U2402);
  nand ginst28549 (P3_U6374, P3_U4318, P3_U6372);
  nand ginst28550 (P3_U6375, P3_INSTADDRPOINTER_REG_30__SCAN_IN, P3_U5631);
  nand ginst28551 (P3_U6376, P3_ADD_360_1242_U90, P3_U2395);
  nand ginst28552 (P3_U6377, P3_SUB_357_1258_U20, P3_U2393);
  nand ginst28553 (P3_U6378, P3_ADD_558_U72, P3_U3220);
  nand ginst28554 (P3_U6379, P3_ADD_553_U72, P3_U4298);
  nand ginst28555 (P3_U6380, P3_ADD_547_U72, P3_U4299);
  nand ginst28556 (P3_U6381, P3_ADD_541_U69, P3_U4300);
  nand ginst28557 (P3_U6382, P3_ADD_536_U69, P3_U4301);
  nand ginst28558 (P3_U6383, P3_ADD_531_U72, P3_U2354);
  nand ginst28559 (P3_U6384, P3_ADD_526_U58, P3_U2355);
  nand ginst28560 (P3_U6385, P3_ADD_515_U69, P3_U4302);
  nand ginst28561 (P3_U6386, P3_ADD_494_U69, P3_U2356);
  nand ginst28562 (P3_U6387, P3_ADD_476_U69, P3_U4303);
  nand ginst28563 (P3_U6388, P3_ADD_441_U69, P3_U4304);
  nand ginst28564 (P3_U6389, P3_ADD_405_U69, P3_U4305);
  nand ginst28565 (P3_U6390, P3_ADD_394_U69, P3_U2357);
  nand ginst28566 (P3_U6391, P3_ADD_385_U72, P3_U2358);
  nand ginst28567 (P3_U6392, P3_ADD_380_U72, P3_U2359);
  nand ginst28568 (P3_U6393, P3_ADD_349_U72, P3_U4306);
  nand ginst28569 (P3_U6394, P3_ADD_344_U72, P3_U2362);
  nand ginst28570 (P3_U6395, P3_ADD_371_1212_U92, P3_U2360);
  nand ginst28571 (P3_U6396, P3_U3945, P3_U3950);
  nand ginst28572 (P3_U6397, P3_REIP_REG_31__SCAN_IN, P3_U2402);
  nand ginst28573 (P3_U6398, P3_INSTADDRPOINTER_REG_31__SCAN_IN, P3_U5631);
  nand ginst28574 (P3_U6399, P3_GTE_355_U6, P3_U2361);
  nand ginst28575 (P3_U6400, P3_GTE_370_U6, P3_U2360);
  nand ginst28576 (P3_U6401, P3_U6399, P3_U6400);
  nand ginst28577 (P3_U6402, P3_U2390, P3_U6401);
  nand ginst28578 (P3_U6403, P3_U3121, P3_U3234);
  not ginst28579 (P3_U6404, P3_U3249);
  nand ginst28580 (P3_U6405, P3_PHYADDRPOINTER_REG_0__SCAN_IN, P3_U2398);
  nand ginst28581 (P3_U6406, P3_PHYADDRPOINTER_REG_0__SCAN_IN, P3_U2397);
  nand ginst28582 (P3_U6407, P3_ADD_360_1242_U85, P3_U2396);
  nand ginst28583 (P3_U6408, P3_SUB_357_1258_U69, P3_U2394);
  nand ginst28584 (P3_U6409, P3_REIP_REG_0__SCAN_IN, P3_U2389);
  nand ginst28585 (P3_U6410, P3_PHYADDRPOINTER_REG_0__SCAN_IN, P3_U2388);
  nand ginst28586 (P3_U6411, P3_ADD_371_1212_U87, P3_U2387);
  nand ginst28587 (P3_U6412, P3_PHYADDRPOINTER_REG_0__SCAN_IN, P3_U6404);
  nand ginst28588 (P3_U6413, P3_ADD_318_U4, P3_U2398);
  nand ginst28589 (P3_U6414, P3_PHYADDRPOINTER_REG_1__SCAN_IN, P3_U2397);
  nand ginst28590 (P3_U6415, P3_ADD_360_1242_U19, P3_U2396);
  nand ginst28591 (P3_U6416, P3_SUB_357_1258_U21, P3_U2394);
  nand ginst28592 (P3_U6417, P3_REIP_REG_1__SCAN_IN, P3_U2389);
  nand ginst28593 (P3_U6418, P3_ADD_339_U4, P3_U2388);
  nand ginst28594 (P3_U6419, P3_ADD_371_1212_U20, P3_U2387);
  nand ginst28595 (P3_U6420, P3_PHYADDRPOINTER_REG_1__SCAN_IN, P3_U6404);
  nand ginst28596 (P3_U6421, P3_ADD_318_U71, P3_U2398);
  nand ginst28597 (P3_U6422, P3_ADD_315_U4, P3_U2397);
  nand ginst28598 (P3_U6423, P3_ADD_360_1242_U91, P3_U2396);
  nand ginst28599 (P3_U6424, P3_SUB_357_1258_U78, P3_U2394);
  nand ginst28600 (P3_U6425, P3_REIP_REG_2__SCAN_IN, P3_U2389);
  nand ginst28601 (P3_U6426, P3_ADD_339_U71, P3_U2388);
  nand ginst28602 (P3_U6427, P3_ADD_371_1212_U93, P3_U2387);
  nand ginst28603 (P3_U6428, P3_PHYADDRPOINTER_REG_2__SCAN_IN, P3_U6404);
  nand ginst28604 (P3_U6429, P3_ADD_318_U68, P3_U2398);
  nand ginst28605 (P3_U6430, P3_ADD_315_U66, P3_U2397);
  nand ginst28606 (P3_U6431, P3_ADD_360_1242_U17, P3_U2396);
  nand ginst28607 (P3_U6432, P3_SUB_357_1258_U76, P3_U2394);
  nand ginst28608 (P3_U6433, P3_REIP_REG_3__SCAN_IN, P3_U2389);
  nand ginst28609 (P3_U6434, P3_ADD_339_U68, P3_U2388);
  nand ginst28610 (P3_U6435, P3_ADD_371_1212_U18, P3_U2387);
  nand ginst28611 (P3_U6436, P3_PHYADDRPOINTER_REG_3__SCAN_IN, P3_U6404);
  nand ginst28612 (P3_U6437, P3_ADD_318_U67, P3_U2398);
  nand ginst28613 (P3_U6438, P3_ADD_315_U65, P3_U2397);
  nand ginst28614 (P3_U6439, P3_ADD_360_1242_U18, P3_U2396);
  nand ginst28615 (P3_U6440, P3_SUB_357_1258_U75, P3_U2394);
  nand ginst28616 (P3_U6441, P3_REIP_REG_4__SCAN_IN, P3_U2389);
  nand ginst28617 (P3_U6442, P3_ADD_339_U67, P3_U2388);
  nand ginst28618 (P3_U6443, P3_ADD_371_1212_U91, P3_U2387);
  nand ginst28619 (P3_U6444, P3_PHYADDRPOINTER_REG_4__SCAN_IN, P3_U6404);
  nand ginst28620 (P3_U6445, P3_ADD_318_U66, P3_U2398);
  nand ginst28621 (P3_U6446, P3_ADD_315_U64, P3_U2397);
  nand ginst28622 (P3_U6447, P3_ADD_360_1242_U89, P3_U2396);
  nand ginst28623 (P3_U6448, P3_SUB_357_1258_U74, P3_U2394);
  nand ginst28624 (P3_U6449, P3_REIP_REG_5__SCAN_IN, P3_U2389);
  nand ginst28625 (P3_U6450, P3_ADD_339_U66, P3_U2388);
  nand ginst28626 (P3_U6451, P3_ADD_371_1212_U19, P3_U2387);
  nand ginst28627 (P3_U6452, P3_PHYADDRPOINTER_REG_5__SCAN_IN, P3_U6404);
  nand ginst28628 (P3_U6453, P3_ADD_318_U65, P3_U2398);
  nand ginst28629 (P3_U6454, P3_ADD_315_U63, P3_U2397);
  nand ginst28630 (P3_U6455, P3_ADD_360_1242_U88, P3_U2396);
  nand ginst28631 (P3_U6456, P3_SUB_357_1258_U73, P3_U2394);
  nand ginst28632 (P3_U6457, P3_REIP_REG_6__SCAN_IN, P3_U2389);
  nand ginst28633 (P3_U6458, P3_ADD_339_U65, P3_U2388);
  nand ginst28634 (P3_U6459, P3_ADD_371_1212_U90, P3_U2387);
  nand ginst28635 (P3_U6460, P3_PHYADDRPOINTER_REG_6__SCAN_IN, P3_U6404);
  nand ginst28636 (P3_U6461, P3_ADD_318_U64, P3_U2398);
  nand ginst28637 (P3_U6462, P3_ADD_315_U62, P3_U2397);
  nand ginst28638 (P3_U6463, P3_ADD_360_1242_U87, P3_U2396);
  nand ginst28639 (P3_U6464, P3_SUB_357_1258_U72, P3_U2394);
  nand ginst28640 (P3_U6465, P3_REIP_REG_7__SCAN_IN, P3_U2389);
  nand ginst28641 (P3_U6466, P3_ADD_339_U64, P3_U2388);
  nand ginst28642 (P3_U6467, P3_ADD_371_1212_U89, P3_U2387);
  nand ginst28643 (P3_U6468, P3_PHYADDRPOINTER_REG_7__SCAN_IN, P3_U6404);
  nand ginst28644 (P3_U6469, P3_ADD_318_U63, P3_U2398);
  nand ginst28645 (P3_U6470, P3_ADD_315_U61, P3_U2397);
  nand ginst28646 (P3_U6471, P3_ADD_360_1242_U86, P3_U2396);
  nand ginst28647 (P3_U6472, P3_SUB_357_1258_U71, P3_U2394);
  nand ginst28648 (P3_U6473, P3_REIP_REG_8__SCAN_IN, P3_U2389);
  nand ginst28649 (P3_U6474, P3_ADD_339_U63, P3_U2388);
  nand ginst28650 (P3_U6475, P3_ADD_371_1212_U88, P3_U2387);
  nand ginst28651 (P3_U6476, P3_PHYADDRPOINTER_REG_8__SCAN_IN, P3_U6404);
  nand ginst28652 (P3_U6477, P3_ADD_318_U62, P3_U2398);
  nand ginst28653 (P3_U6478, P3_ADD_315_U60, P3_U2397);
  nand ginst28654 (P3_U6479, P3_ADD_360_1242_U106, P3_U2396);
  nand ginst28655 (P3_U6480, P3_SUB_357_1258_U70, P3_U2394);
  nand ginst28656 (P3_U6481, P3_REIP_REG_9__SCAN_IN, P3_U2389);
  nand ginst28657 (P3_U6482, P3_ADD_339_U62, P3_U2388);
  nand ginst28658 (P3_U6483, P3_ADD_371_1212_U109, P3_U2387);
  nand ginst28659 (P3_U6484, P3_PHYADDRPOINTER_REG_9__SCAN_IN, P3_U6404);
  nand ginst28660 (P3_U6485, P3_ADD_318_U91, P3_U2398);
  nand ginst28661 (P3_U6486, P3_ADD_315_U88, P3_U2397);
  nand ginst28662 (P3_U6487, P3_ADD_360_1242_U4, P3_U2396);
  nand ginst28663 (P3_U6488, P3_SUB_357_1258_U93, P3_U2394);
  nand ginst28664 (P3_U6489, P3_REIP_REG_10__SCAN_IN, P3_U2389);
  nand ginst28665 (P3_U6490, P3_ADD_339_U91, P3_U2388);
  nand ginst28666 (P3_U6491, P3_ADD_371_1212_U5, P3_U2387);
  nand ginst28667 (P3_U6492, P3_PHYADDRPOINTER_REG_10__SCAN_IN, P3_U6404);
  nand ginst28668 (P3_U6493, P3_ADD_318_U90, P3_U2398);
  nand ginst28669 (P3_U6494, P3_ADD_315_U87, P3_U2397);
  nand ginst28670 (P3_U6495, P3_ADD_360_1242_U84, P3_U2396);
  nand ginst28671 (P3_U6496, P3_SUB_357_1258_U92, P3_U2394);
  nand ginst28672 (P3_U6497, P3_REIP_REG_11__SCAN_IN, P3_U2389);
  nand ginst28673 (P3_U6498, P3_ADD_339_U90, P3_U2388);
  nand ginst28674 (P3_U6499, P3_ADD_371_1212_U86, P3_U2387);
  nand ginst28675 (P3_U6500, P3_PHYADDRPOINTER_REG_11__SCAN_IN, P3_U6404);
  nand ginst28676 (P3_U6501, P3_ADD_318_U89, P3_U2398);
  nand ginst28677 (P3_U6502, P3_ADD_315_U86, P3_U2397);
  nand ginst28678 (P3_U6503, P3_ADD_360_1242_U5, P3_U2396);
  nand ginst28679 (P3_U6504, P3_SUB_357_1258_U91, P3_U2394);
  nand ginst28680 (P3_U6505, P3_REIP_REG_12__SCAN_IN, P3_U2389);
  nand ginst28681 (P3_U6506, P3_ADD_339_U89, P3_U2388);
  nand ginst28682 (P3_U6507, P3_ADD_371_1212_U6, P3_U2387);
  nand ginst28683 (P3_U6508, P3_PHYADDRPOINTER_REG_12__SCAN_IN, P3_U6404);
  nand ginst28684 (P3_U6509, P3_ADD_318_U88, P3_U2398);
  nand ginst28685 (P3_U6510, P3_ADD_315_U85, P3_U2397);
  nand ginst28686 (P3_U6511, P3_ADD_360_1242_U6, P3_U2396);
  nand ginst28687 (P3_U6512, P3_SUB_357_1258_U15, P3_U2394);
  nand ginst28688 (P3_U6513, P3_REIP_REG_13__SCAN_IN, P3_U2389);
  nand ginst28689 (P3_U6514, P3_ADD_339_U88, P3_U2388);
  nand ginst28690 (P3_U6515, P3_ADD_371_1212_U7, P3_U2387);
  nand ginst28691 (P3_U6516, P3_PHYADDRPOINTER_REG_13__SCAN_IN, P3_U6404);
  nand ginst28692 (P3_U6517, P3_ADD_318_U87, P3_U2398);
  nand ginst28693 (P3_U6518, P3_ADD_315_U84, P3_U2397);
  nand ginst28694 (P3_U6519, P3_ADD_360_1242_U83, P3_U2396);
  nand ginst28695 (P3_U6520, P3_SUB_357_1258_U90, P3_U2394);
  nand ginst28696 (P3_U6521, P3_REIP_REG_14__SCAN_IN, P3_U2389);
  nand ginst28697 (P3_U6522, P3_ADD_339_U87, P3_U2388);
  nand ginst28698 (P3_U6523, P3_ADD_371_1212_U85, P3_U2387);
  nand ginst28699 (P3_U6524, P3_PHYADDRPOINTER_REG_14__SCAN_IN, P3_U6404);
  nand ginst28700 (P3_U6525, P3_ADD_318_U86, P3_U2398);
  nand ginst28701 (P3_U6526, P3_ADD_315_U83, P3_U2397);
  nand ginst28702 (P3_U6527, P3_ADD_360_1242_U7, P3_U2396);
  nand ginst28703 (P3_U6528, P3_SUB_357_1258_U89, P3_U2394);
  nand ginst28704 (P3_U6529, P3_REIP_REG_15__SCAN_IN, P3_U2389);
  nand ginst28705 (P3_U6530, P3_ADD_339_U86, P3_U2388);
  nand ginst28706 (P3_U6531, P3_ADD_371_1212_U8, P3_U2387);
  nand ginst28707 (P3_U6532, P3_PHYADDRPOINTER_REG_15__SCAN_IN, P3_U6404);
  nand ginst28708 (P3_U6533, P3_ADD_318_U85, P3_U2398);
  nand ginst28709 (P3_U6534, P3_ADD_315_U82, P3_U2397);
  nand ginst28710 (P3_U6535, P3_ADD_360_1242_U82, P3_U2396);
  nand ginst28711 (P3_U6536, P3_SUB_357_1258_U88, P3_U2394);
  nand ginst28712 (P3_U6537, P3_REIP_REG_16__SCAN_IN, P3_U2389);
  nand ginst28713 (P3_U6538, P3_ADD_339_U85, P3_U2388);
  nand ginst28714 (P3_U6539, P3_ADD_371_1212_U84, P3_U2387);
  nand ginst28715 (P3_U6540, P3_PHYADDRPOINTER_REG_16__SCAN_IN, P3_U6404);
  nand ginst28716 (P3_U6541, P3_ADD_318_U84, P3_U2398);
  nand ginst28717 (P3_U6542, P3_ADD_315_U81, P3_U2397);
  nand ginst28718 (P3_U6543, P3_ADD_360_1242_U8, P3_U2396);
  nand ginst28719 (P3_U6544, P3_SUB_357_1258_U16, P3_U2394);
  nand ginst28720 (P3_U6545, P3_REIP_REG_17__SCAN_IN, P3_U2389);
  nand ginst28721 (P3_U6546, P3_ADD_339_U84, P3_U2388);
  nand ginst28722 (P3_U6547, P3_ADD_371_1212_U9, P3_U2387);
  nand ginst28723 (P3_U6548, P3_PHYADDRPOINTER_REG_17__SCAN_IN, P3_U6404);
  nand ginst28724 (P3_U6549, P3_ADD_318_U83, P3_U2398);
  nand ginst28725 (P3_U6550, P3_ADD_315_U80, P3_U2397);
  nand ginst28726 (P3_U6551, P3_ADD_360_1242_U81, P3_U2396);
  nand ginst28727 (P3_U6552, P3_SUB_357_1258_U87, P3_U2394);
  nand ginst28728 (P3_U6553, P3_REIP_REG_18__SCAN_IN, P3_U2389);
  nand ginst28729 (P3_U6554, P3_ADD_339_U83, P3_U2388);
  nand ginst28730 (P3_U6555, P3_ADD_371_1212_U83, P3_U2387);
  nand ginst28731 (P3_U6556, P3_PHYADDRPOINTER_REG_18__SCAN_IN, P3_U6404);
  nand ginst28732 (P3_U6557, P3_ADD_318_U82, P3_U2398);
  nand ginst28733 (P3_U6558, P3_ADD_315_U79, P3_U2397);
  nand ginst28734 (P3_U6559, P3_ADD_360_1242_U9, P3_U2396);
  nand ginst28735 (P3_U6560, P3_SUB_357_1258_U86, P3_U2394);
  nand ginst28736 (P3_U6561, P3_REIP_REG_19__SCAN_IN, P3_U2389);
  nand ginst28737 (P3_U6562, P3_ADD_339_U82, P3_U2388);
  nand ginst28738 (P3_U6563, P3_ADD_371_1212_U10, P3_U2387);
  nand ginst28739 (P3_U6564, P3_PHYADDRPOINTER_REG_19__SCAN_IN, P3_U6404);
  nand ginst28740 (P3_U6565, P3_ADD_318_U81, P3_U2398);
  nand ginst28741 (P3_U6566, P3_ADD_315_U78, P3_U2397);
  nand ginst28742 (P3_U6567, P3_ADD_360_1242_U10, P3_U2396);
  nand ginst28743 (P3_U6568, P3_SUB_357_1258_U17, P3_U2394);
  nand ginst28744 (P3_U6569, P3_REIP_REG_20__SCAN_IN, P3_U2389);
  nand ginst28745 (P3_U6570, P3_ADD_339_U81, P3_U2388);
  nand ginst28746 (P3_U6571, P3_ADD_371_1212_U11, P3_U2387);
  nand ginst28747 (P3_U6572, P3_PHYADDRPOINTER_REG_20__SCAN_IN, P3_U6404);
  nand ginst28748 (P3_U6573, P3_ADD_318_U80, P3_U2398);
  nand ginst28749 (P3_U6574, P3_ADD_315_U77, P3_U2397);
  nand ginst28750 (P3_U6575, P3_ADD_360_1242_U11, P3_U2396);
  nand ginst28751 (P3_U6576, P3_SUB_357_1258_U85, P3_U2394);
  nand ginst28752 (P3_U6577, P3_REIP_REG_21__SCAN_IN, P3_U2389);
  nand ginst28753 (P3_U6578, P3_ADD_339_U80, P3_U2388);
  nand ginst28754 (P3_U6579, P3_ADD_371_1212_U12, P3_U2387);
  nand ginst28755 (P3_U6580, P3_PHYADDRPOINTER_REG_21__SCAN_IN, P3_U6404);
  nand ginst28756 (P3_U6581, P3_ADD_318_U79, P3_U2398);
  nand ginst28757 (P3_U6582, P3_ADD_315_U76, P3_U2397);
  nand ginst28758 (P3_U6583, P3_ADD_360_1242_U80, P3_U2396);
  nand ginst28759 (P3_U6584, P3_SUB_357_1258_U84, P3_U2394);
  nand ginst28760 (P3_U6585, P3_REIP_REG_22__SCAN_IN, P3_U2389);
  nand ginst28761 (P3_U6586, P3_ADD_339_U79, P3_U2388);
  nand ginst28762 (P3_U6587, P3_ADD_371_1212_U82, P3_U2387);
  nand ginst28763 (P3_U6588, P3_PHYADDRPOINTER_REG_22__SCAN_IN, P3_U6404);
  nand ginst28764 (P3_U6589, P3_ADD_318_U78, P3_U2398);
  nand ginst28765 (P3_U6590, P3_ADD_315_U75, P3_U2397);
  nand ginst28766 (P3_U6591, P3_ADD_360_1242_U12, P3_U2396);
  nand ginst28767 (P3_U6592, P3_SUB_357_1258_U83, P3_U2394);
  nand ginst28768 (P3_U6593, P3_REIP_REG_23__SCAN_IN, P3_U2389);
  nand ginst28769 (P3_U6594, P3_ADD_339_U78, P3_U2388);
  nand ginst28770 (P3_U6595, P3_ADD_371_1212_U13, P3_U2387);
  nand ginst28771 (P3_U6596, P3_PHYADDRPOINTER_REG_23__SCAN_IN, P3_U6404);
  nand ginst28772 (P3_U6597, P3_ADD_318_U77, P3_U2398);
  nand ginst28773 (P3_U6598, P3_ADD_315_U74, P3_U2397);
  nand ginst28774 (P3_U6599, P3_ADD_360_1242_U79, P3_U2396);
  nand ginst28775 (P3_U6600, P3_SUB_357_1258_U82, P3_U2394);
  nand ginst28776 (P3_U6601, P3_REIP_REG_24__SCAN_IN, P3_U2389);
  nand ginst28777 (P3_U6602, P3_ADD_339_U77, P3_U2388);
  nand ginst28778 (P3_U6603, P3_ADD_371_1212_U81, P3_U2387);
  nand ginst28779 (P3_U6604, P3_PHYADDRPOINTER_REG_24__SCAN_IN, P3_U6404);
  nand ginst28780 (P3_U6605, P3_ADD_318_U76, P3_U2398);
  nand ginst28781 (P3_U6606, P3_ADD_315_U73, P3_U2397);
  nand ginst28782 (P3_U6607, P3_ADD_360_1242_U13, P3_U2396);
  nand ginst28783 (P3_U6608, P3_SUB_357_1258_U81, P3_U2394);
  nand ginst28784 (P3_U6609, P3_REIP_REG_25__SCAN_IN, P3_U2389);
  nand ginst28785 (P3_U6610, P3_ADD_339_U76, P3_U2388);
  nand ginst28786 (P3_U6611, P3_ADD_371_1212_U14, P3_U2387);
  nand ginst28787 (P3_U6612, P3_PHYADDRPOINTER_REG_25__SCAN_IN, P3_U6404);
  nand ginst28788 (P3_U6613, P3_ADD_318_U75, P3_U2398);
  nand ginst28789 (P3_U6614, P3_ADD_315_U72, P3_U2397);
  nand ginst28790 (P3_U6615, P3_ADD_360_1242_U14, P3_U2396);
  nand ginst28791 (P3_U6616, P3_SUB_357_1258_U18, P3_U2394);
  nand ginst28792 (P3_U6617, P3_REIP_REG_26__SCAN_IN, P3_U2389);
  nand ginst28793 (P3_U6618, P3_ADD_339_U75, P3_U2388);
  nand ginst28794 (P3_U6619, P3_ADD_371_1212_U15, P3_U2387);
  nand ginst28795 (P3_U6620, P3_PHYADDRPOINTER_REG_26__SCAN_IN, P3_U6404);
  nand ginst28796 (P3_U6621, P3_ADD_318_U74, P3_U2398);
  nand ginst28797 (P3_U6622, P3_ADD_315_U71, P3_U2397);
  nand ginst28798 (P3_U6623, P3_ADD_360_1242_U78, P3_U2396);
  nand ginst28799 (P3_U6624, P3_SUB_357_1258_U80, P3_U2394);
  nand ginst28800 (P3_U6625, P3_REIP_REG_27__SCAN_IN, P3_U2389);
  nand ginst28801 (P3_U6626, P3_ADD_339_U74, P3_U2388);
  nand ginst28802 (P3_U6627, P3_ADD_371_1212_U80, P3_U2387);
  nand ginst28803 (P3_U6628, P3_PHYADDRPOINTER_REG_27__SCAN_IN, P3_U6404);
  nand ginst28804 (P3_U6629, P3_ADD_318_U73, P3_U2398);
  nand ginst28805 (P3_U6630, P3_ADD_315_U70, P3_U2397);
  nand ginst28806 (P3_U6631, P3_ADD_360_1242_U15, P3_U2396);
  nand ginst28807 (P3_U6632, P3_SUB_357_1258_U19, P3_U2394);
  nand ginst28808 (P3_U6633, P3_REIP_REG_28__SCAN_IN, P3_U2389);
  nand ginst28809 (P3_U6634, P3_ADD_339_U73, P3_U2388);
  nand ginst28810 (P3_U6635, P3_ADD_371_1212_U16, P3_U2387);
  nand ginst28811 (P3_U6636, P3_PHYADDRPOINTER_REG_28__SCAN_IN, P3_U6404);
  nand ginst28812 (P3_U6637, P3_ADD_318_U72, P3_U2398);
  nand ginst28813 (P3_U6638, P3_ADD_315_U69, P3_U2397);
  nand ginst28814 (P3_U6639, P3_ADD_360_1242_U16, P3_U2396);
  nand ginst28815 (P3_U6640, P3_SUB_357_1258_U79, P3_U2394);
  nand ginst28816 (P3_U6641, P3_REIP_REG_29__SCAN_IN, P3_U2389);
  nand ginst28817 (P3_U6642, P3_ADD_339_U72, P3_U2388);
  nand ginst28818 (P3_U6643, P3_ADD_371_1212_U17, P3_U2387);
  nand ginst28819 (P3_U6644, P3_PHYADDRPOINTER_REG_29__SCAN_IN, P3_U6404);
  nand ginst28820 (P3_U6645, P3_ADD_318_U70, P3_U2398);
  nand ginst28821 (P3_U6646, P3_ADD_315_U68, P3_U2397);
  nand ginst28822 (P3_U6647, P3_ADD_360_1242_U77, P3_U2396);
  nand ginst28823 (P3_U6648, P3_SUB_357_1258_U77, P3_U2394);
  nand ginst28824 (P3_U6649, P3_REIP_REG_30__SCAN_IN, P3_U2389);
  nand ginst28825 (P3_U6650, P3_ADD_339_U70, P3_U2388);
  nand ginst28826 (P3_U6651, P3_ADD_371_1212_U79, P3_U2387);
  nand ginst28827 (P3_U6652, P3_PHYADDRPOINTER_REG_30__SCAN_IN, P3_U6404);
  nand ginst28828 (P3_U6653, P3_ADD_318_U69, P3_U2398);
  nand ginst28829 (P3_U6654, P3_ADD_315_U67, P3_U2397);
  nand ginst28830 (P3_U6655, P3_ADD_360_1242_U90, P3_U2396);
  nand ginst28831 (P3_U6656, P3_SUB_357_1258_U20, P3_U2394);
  nand ginst28832 (P3_U6657, P3_REIP_REG_31__SCAN_IN, P3_U2389);
  nand ginst28833 (P3_U6658, P3_ADD_339_U69, P3_U2388);
  nand ginst28834 (P3_U6659, P3_ADD_371_1212_U92, P3_U2387);
  nand ginst28835 (P3_U6660, P3_PHYADDRPOINTER_REG_31__SCAN_IN, P3_U6404);
  nand ginst28836 (P3_U6661, P3_GTE_412_U6, P3_U2630, P3_U4304);
  nand ginst28837 (P3_U6662, P3_GTE_450_U6, P3_U4303);
  nand ginst28838 (P3_U6663, P3_U6661, P3_U6662);
  nand ginst28839 (P3_U6664, P3_EAX_REG_15__SCAN_IN, P3_U2407);
  nand ginst28840 (P3_U6665, BUF2_REG_15__SCAN_IN, P3_U2406);
  nand ginst28841 (P3_U6666, P3_LWORD_REG_15__SCAN_IN, P3_U3250);
  nand ginst28842 (P3_U6667, P3_EAX_REG_14__SCAN_IN, P3_U2407);
  nand ginst28843 (P3_U6668, BUF2_REG_14__SCAN_IN, P3_U2406);
  nand ginst28844 (P3_U6669, P3_LWORD_REG_14__SCAN_IN, P3_U3250);
  nand ginst28845 (P3_U6670, P3_EAX_REG_13__SCAN_IN, P3_U2407);
  nand ginst28846 (P3_U6671, BUF2_REG_13__SCAN_IN, P3_U2406);
  nand ginst28847 (P3_U6672, P3_LWORD_REG_13__SCAN_IN, P3_U3250);
  nand ginst28848 (P3_U6673, P3_EAX_REG_12__SCAN_IN, P3_U2407);
  nand ginst28849 (P3_U6674, BUF2_REG_12__SCAN_IN, P3_U2406);
  nand ginst28850 (P3_U6675, P3_LWORD_REG_12__SCAN_IN, P3_U3250);
  nand ginst28851 (P3_U6676, P3_EAX_REG_11__SCAN_IN, P3_U2407);
  nand ginst28852 (P3_U6677, BUF2_REG_11__SCAN_IN, P3_U2406);
  nand ginst28853 (P3_U6678, P3_LWORD_REG_11__SCAN_IN, P3_U3250);
  nand ginst28854 (P3_U6679, P3_EAX_REG_10__SCAN_IN, P3_U2407);
  nand ginst28855 (P3_U6680, BUF2_REG_10__SCAN_IN, P3_U2406);
  nand ginst28856 (P3_U6681, P3_LWORD_REG_10__SCAN_IN, P3_U3250);
  nand ginst28857 (P3_U6682, P3_EAX_REG_9__SCAN_IN, P3_U2407);
  nand ginst28858 (P3_U6683, BUF2_REG_9__SCAN_IN, P3_U2406);
  nand ginst28859 (P3_U6684, P3_LWORD_REG_9__SCAN_IN, P3_U3250);
  nand ginst28860 (P3_U6685, P3_EAX_REG_8__SCAN_IN, P3_U2407);
  nand ginst28861 (P3_U6686, BUF2_REG_8__SCAN_IN, P3_U2406);
  nand ginst28862 (P3_U6687, P3_LWORD_REG_8__SCAN_IN, P3_U3250);
  nand ginst28863 (P3_U6688, P3_EAX_REG_7__SCAN_IN, P3_U2407);
  nand ginst28864 (P3_U6689, BUF2_REG_7__SCAN_IN, P3_U2406);
  nand ginst28865 (P3_U6690, P3_LWORD_REG_7__SCAN_IN, P3_U3250);
  nand ginst28866 (P3_U6691, P3_EAX_REG_6__SCAN_IN, P3_U2407);
  nand ginst28867 (P3_U6692, BUF2_REG_6__SCAN_IN, P3_U2406);
  nand ginst28868 (P3_U6693, P3_LWORD_REG_6__SCAN_IN, P3_U3250);
  nand ginst28869 (P3_U6694, P3_EAX_REG_5__SCAN_IN, P3_U2407);
  nand ginst28870 (P3_U6695, BUF2_REG_5__SCAN_IN, P3_U2406);
  nand ginst28871 (P3_U6696, P3_LWORD_REG_5__SCAN_IN, P3_U3250);
  nand ginst28872 (P3_U6697, P3_EAX_REG_4__SCAN_IN, P3_U2407);
  nand ginst28873 (P3_U6698, BUF2_REG_4__SCAN_IN, P3_U2406);
  nand ginst28874 (P3_U6699, P3_LWORD_REG_4__SCAN_IN, P3_U3250);
  nand ginst28875 (P3_U6700, P3_EAX_REG_3__SCAN_IN, P3_U2407);
  nand ginst28876 (P3_U6701, BUF2_REG_3__SCAN_IN, P3_U2406);
  nand ginst28877 (P3_U6702, P3_LWORD_REG_3__SCAN_IN, P3_U3250);
  nand ginst28878 (P3_U6703, P3_EAX_REG_2__SCAN_IN, P3_U2407);
  nand ginst28879 (P3_U6704, BUF2_REG_2__SCAN_IN, P3_U2406);
  nand ginst28880 (P3_U6705, P3_LWORD_REG_2__SCAN_IN, P3_U3250);
  nand ginst28881 (P3_U6706, P3_EAX_REG_1__SCAN_IN, P3_U2407);
  nand ginst28882 (P3_U6707, BUF2_REG_1__SCAN_IN, P3_U2406);
  nand ginst28883 (P3_U6708, P3_LWORD_REG_1__SCAN_IN, P3_U3250);
  nand ginst28884 (P3_U6709, P3_EAX_REG_0__SCAN_IN, P3_U2407);
  nand ginst28885 (P3_U6710, BUF2_REG_0__SCAN_IN, P3_U2406);
  nand ginst28886 (P3_U6711, P3_LWORD_REG_0__SCAN_IN, P3_U3250);
  nand ginst28887 (P3_U6712, P3_EAX_REG_30__SCAN_IN, P3_U2407);
  nand ginst28888 (P3_U6713, BUF2_REG_14__SCAN_IN, P3_U2406);
  nand ginst28889 (P3_U6714, P3_UWORD_REG_14__SCAN_IN, P3_U3250);
  nand ginst28890 (P3_U6715, P3_EAX_REG_29__SCAN_IN, P3_U2407);
  nand ginst28891 (P3_U6716, BUF2_REG_13__SCAN_IN, P3_U2406);
  nand ginst28892 (P3_U6717, P3_UWORD_REG_13__SCAN_IN, P3_U3250);
  nand ginst28893 (P3_U6718, P3_EAX_REG_28__SCAN_IN, P3_U2407);
  nand ginst28894 (P3_U6719, BUF2_REG_12__SCAN_IN, P3_U2406);
  nand ginst28895 (P3_U6720, P3_UWORD_REG_12__SCAN_IN, P3_U3250);
  nand ginst28896 (P3_U6721, P3_EAX_REG_27__SCAN_IN, P3_U2407);
  nand ginst28897 (P3_U6722, BUF2_REG_11__SCAN_IN, P3_U2406);
  nand ginst28898 (P3_U6723, P3_UWORD_REG_11__SCAN_IN, P3_U3250);
  nand ginst28899 (P3_U6724, P3_EAX_REG_26__SCAN_IN, P3_U2407);
  nand ginst28900 (P3_U6725, BUF2_REG_10__SCAN_IN, P3_U2406);
  nand ginst28901 (P3_U6726, P3_UWORD_REG_10__SCAN_IN, P3_U3250);
  nand ginst28902 (P3_U6727, P3_EAX_REG_25__SCAN_IN, P3_U2407);
  nand ginst28903 (P3_U6728, BUF2_REG_9__SCAN_IN, P3_U2406);
  nand ginst28904 (P3_U6729, P3_UWORD_REG_9__SCAN_IN, P3_U3250);
  nand ginst28905 (P3_U6730, P3_EAX_REG_24__SCAN_IN, P3_U2407);
  nand ginst28906 (P3_U6731, BUF2_REG_8__SCAN_IN, P3_U2406);
  nand ginst28907 (P3_U6732, P3_UWORD_REG_8__SCAN_IN, P3_U3250);
  nand ginst28908 (P3_U6733, P3_EAX_REG_23__SCAN_IN, P3_U2407);
  nand ginst28909 (P3_U6734, BUF2_REG_7__SCAN_IN, P3_U2406);
  nand ginst28910 (P3_U6735, P3_UWORD_REG_7__SCAN_IN, P3_U3250);
  nand ginst28911 (P3_U6736, P3_EAX_REG_22__SCAN_IN, P3_U2407);
  nand ginst28912 (P3_U6737, BUF2_REG_6__SCAN_IN, P3_U2406);
  nand ginst28913 (P3_U6738, P3_UWORD_REG_6__SCAN_IN, P3_U3250);
  nand ginst28914 (P3_U6739, P3_EAX_REG_21__SCAN_IN, P3_U2407);
  nand ginst28915 (P3_U6740, BUF2_REG_5__SCAN_IN, P3_U2406);
  nand ginst28916 (P3_U6741, P3_UWORD_REG_5__SCAN_IN, P3_U3250);
  nand ginst28917 (P3_U6742, P3_EAX_REG_20__SCAN_IN, P3_U2407);
  nand ginst28918 (P3_U6743, BUF2_REG_4__SCAN_IN, P3_U2406);
  nand ginst28919 (P3_U6744, P3_UWORD_REG_4__SCAN_IN, P3_U3250);
  nand ginst28920 (P3_U6745, P3_EAX_REG_19__SCAN_IN, P3_U2407);
  nand ginst28921 (P3_U6746, BUF2_REG_3__SCAN_IN, P3_U2406);
  nand ginst28922 (P3_U6747, P3_UWORD_REG_3__SCAN_IN, P3_U3250);
  nand ginst28923 (P3_U6748, P3_EAX_REG_18__SCAN_IN, P3_U2407);
  nand ginst28924 (P3_U6749, BUF2_REG_2__SCAN_IN, P3_U2406);
  nand ginst28925 (P3_U6750, P3_UWORD_REG_2__SCAN_IN, P3_U3250);
  nand ginst28926 (P3_U6751, P3_EAX_REG_17__SCAN_IN, P3_U2407);
  nand ginst28927 (P3_U6752, BUF2_REG_1__SCAN_IN, P3_U2406);
  nand ginst28928 (P3_U6753, P3_UWORD_REG_1__SCAN_IN, P3_U3250);
  nand ginst28929 (P3_U6754, P3_EAX_REG_16__SCAN_IN, P3_U2407);
  nand ginst28930 (P3_U6755, BUF2_REG_0__SCAN_IN, P3_U2406);
  nand ginst28931 (P3_U6756, P3_UWORD_REG_0__SCAN_IN, P3_U3250);
  nand ginst28932 (P3_U6757, P3_U3255, P3_U3986);
  nand ginst28933 (P3_U6758, P3_U2453, P3_U3121);
  not ginst28934 (P3_U6759, P3_U3251);
  nand ginst28935 (P3_U6760, P3_LWORD_REG_0__SCAN_IN, P3_U2410);
  nand ginst28936 (P3_U6761, P3_EAX_REG_0__SCAN_IN, P3_U2409);
  nand ginst28937 (P3_U6762, P3_DATAO_REG_0__SCAN_IN, P3_U6759);
  nand ginst28938 (P3_U6763, P3_LWORD_REG_1__SCAN_IN, P3_U2410);
  nand ginst28939 (P3_U6764, P3_EAX_REG_1__SCAN_IN, P3_U2409);
  nand ginst28940 (P3_U6765, P3_DATAO_REG_1__SCAN_IN, P3_U6759);
  nand ginst28941 (P3_U6766, P3_LWORD_REG_2__SCAN_IN, P3_U2410);
  nand ginst28942 (P3_U6767, P3_EAX_REG_2__SCAN_IN, P3_U2409);
  nand ginst28943 (P3_U6768, P3_DATAO_REG_2__SCAN_IN, P3_U6759);
  nand ginst28944 (P3_U6769, P3_LWORD_REG_3__SCAN_IN, P3_U2410);
  nand ginst28945 (P3_U6770, P3_EAX_REG_3__SCAN_IN, P3_U2409);
  nand ginst28946 (P3_U6771, P3_DATAO_REG_3__SCAN_IN, P3_U6759);
  nand ginst28947 (P3_U6772, P3_LWORD_REG_4__SCAN_IN, P3_U2410);
  nand ginst28948 (P3_U6773, P3_EAX_REG_4__SCAN_IN, P3_U2409);
  nand ginst28949 (P3_U6774, P3_DATAO_REG_4__SCAN_IN, P3_U6759);
  nand ginst28950 (P3_U6775, P3_LWORD_REG_5__SCAN_IN, P3_U2410);
  nand ginst28951 (P3_U6776, P3_EAX_REG_5__SCAN_IN, P3_U2409);
  nand ginst28952 (P3_U6777, P3_DATAO_REG_5__SCAN_IN, P3_U6759);
  nand ginst28953 (P3_U6778, P3_LWORD_REG_6__SCAN_IN, P3_U2410);
  nand ginst28954 (P3_U6779, P3_EAX_REG_6__SCAN_IN, P3_U2409);
  nand ginst28955 (P3_U6780, P3_DATAO_REG_6__SCAN_IN, P3_U6759);
  nand ginst28956 (P3_U6781, P3_LWORD_REG_7__SCAN_IN, P3_U2410);
  nand ginst28957 (P3_U6782, P3_EAX_REG_7__SCAN_IN, P3_U2409);
  nand ginst28958 (P3_U6783, P3_DATAO_REG_7__SCAN_IN, P3_U6759);
  nand ginst28959 (P3_U6784, P3_LWORD_REG_8__SCAN_IN, P3_U2410);
  nand ginst28960 (P3_U6785, P3_EAX_REG_8__SCAN_IN, P3_U2409);
  nand ginst28961 (P3_U6786, P3_DATAO_REG_8__SCAN_IN, P3_U6759);
  nand ginst28962 (P3_U6787, P3_LWORD_REG_9__SCAN_IN, P3_U2410);
  nand ginst28963 (P3_U6788, P3_EAX_REG_9__SCAN_IN, P3_U2409);
  nand ginst28964 (P3_U6789, P3_DATAO_REG_9__SCAN_IN, P3_U6759);
  nand ginst28965 (P3_U6790, P3_LWORD_REG_10__SCAN_IN, P3_U2410);
  nand ginst28966 (P3_U6791, P3_EAX_REG_10__SCAN_IN, P3_U2409);
  nand ginst28967 (P3_U6792, P3_DATAO_REG_10__SCAN_IN, P3_U6759);
  nand ginst28968 (P3_U6793, P3_LWORD_REG_11__SCAN_IN, P3_U2410);
  nand ginst28969 (P3_U6794, P3_EAX_REG_11__SCAN_IN, P3_U2409);
  nand ginst28970 (P3_U6795, P3_DATAO_REG_11__SCAN_IN, P3_U6759);
  nand ginst28971 (P3_U6796, P3_LWORD_REG_12__SCAN_IN, P3_U2410);
  nand ginst28972 (P3_U6797, P3_EAX_REG_12__SCAN_IN, P3_U2409);
  nand ginst28973 (P3_U6798, P3_DATAO_REG_12__SCAN_IN, P3_U6759);
  nand ginst28974 (P3_U6799, P3_LWORD_REG_13__SCAN_IN, P3_U2410);
  nand ginst28975 (P3_U6800, P3_EAX_REG_13__SCAN_IN, P3_U2409);
  nand ginst28976 (P3_U6801, P3_DATAO_REG_13__SCAN_IN, P3_U6759);
  nand ginst28977 (P3_U6802, P3_LWORD_REG_14__SCAN_IN, P3_U2410);
  nand ginst28978 (P3_U6803, P3_EAX_REG_14__SCAN_IN, P3_U2409);
  nand ginst28979 (P3_U6804, P3_DATAO_REG_14__SCAN_IN, P3_U6759);
  nand ginst28980 (P3_U6805, P3_LWORD_REG_15__SCAN_IN, P3_U2410);
  nand ginst28981 (P3_U6806, P3_EAX_REG_15__SCAN_IN, P3_U2409);
  nand ginst28982 (P3_U6807, P3_DATAO_REG_15__SCAN_IN, P3_U6759);
  nand ginst28983 (P3_U6808, P3_EAX_REG_16__SCAN_IN, P3_U2447);
  nand ginst28984 (P3_U6809, P3_UWORD_REG_0__SCAN_IN, P3_U2410);
  nand ginst28985 (P3_U6810, P3_DATAO_REG_16__SCAN_IN, P3_U6759);
  nand ginst28986 (P3_U6811, P3_EAX_REG_17__SCAN_IN, P3_U2447);
  nand ginst28987 (P3_U6812, P3_UWORD_REG_1__SCAN_IN, P3_U2410);
  nand ginst28988 (P3_U6813, P3_DATAO_REG_17__SCAN_IN, P3_U6759);
  nand ginst28989 (P3_U6814, P3_EAX_REG_18__SCAN_IN, P3_U2447);
  nand ginst28990 (P3_U6815, P3_UWORD_REG_2__SCAN_IN, P3_U2410);
  nand ginst28991 (P3_U6816, P3_DATAO_REG_18__SCAN_IN, P3_U6759);
  nand ginst28992 (P3_U6817, P3_EAX_REG_19__SCAN_IN, P3_U2447);
  nand ginst28993 (P3_U6818, P3_UWORD_REG_3__SCAN_IN, P3_U2410);
  nand ginst28994 (P3_U6819, P3_DATAO_REG_19__SCAN_IN, P3_U6759);
  nand ginst28995 (P3_U6820, P3_EAX_REG_20__SCAN_IN, P3_U2447);
  nand ginst28996 (P3_U6821, P3_UWORD_REG_4__SCAN_IN, P3_U2410);
  nand ginst28997 (P3_U6822, P3_DATAO_REG_20__SCAN_IN, P3_U6759);
  nand ginst28998 (P3_U6823, P3_EAX_REG_21__SCAN_IN, P3_U2447);
  nand ginst28999 (P3_U6824, P3_UWORD_REG_5__SCAN_IN, P3_U2410);
  nand ginst29000 (P3_U6825, P3_DATAO_REG_21__SCAN_IN, P3_U6759);
  nand ginst29001 (P3_U6826, P3_EAX_REG_22__SCAN_IN, P3_U2447);
  nand ginst29002 (P3_U6827, P3_UWORD_REG_6__SCAN_IN, P3_U2410);
  nand ginst29003 (P3_U6828, P3_DATAO_REG_22__SCAN_IN, P3_U6759);
  nand ginst29004 (P3_U6829, P3_EAX_REG_23__SCAN_IN, P3_U2447);
  nand ginst29005 (P3_U6830, P3_UWORD_REG_7__SCAN_IN, P3_U2410);
  nand ginst29006 (P3_U6831, P3_DATAO_REG_23__SCAN_IN, P3_U6759);
  nand ginst29007 (P3_U6832, P3_EAX_REG_24__SCAN_IN, P3_U2447);
  nand ginst29008 (P3_U6833, P3_UWORD_REG_8__SCAN_IN, P3_U2410);
  nand ginst29009 (P3_U6834, P3_DATAO_REG_24__SCAN_IN, P3_U6759);
  nand ginst29010 (P3_U6835, P3_EAX_REG_25__SCAN_IN, P3_U2447);
  nand ginst29011 (P3_U6836, P3_UWORD_REG_9__SCAN_IN, P3_U2410);
  nand ginst29012 (P3_U6837, P3_DATAO_REG_25__SCAN_IN, P3_U6759);
  nand ginst29013 (P3_U6838, P3_EAX_REG_26__SCAN_IN, P3_U2447);
  nand ginst29014 (P3_U6839, P3_UWORD_REG_10__SCAN_IN, P3_U2410);
  nand ginst29015 (P3_U6840, P3_DATAO_REG_26__SCAN_IN, P3_U6759);
  nand ginst29016 (P3_U6841, P3_EAX_REG_27__SCAN_IN, P3_U2447);
  nand ginst29017 (P3_U6842, P3_UWORD_REG_11__SCAN_IN, P3_U2410);
  nand ginst29018 (P3_U6843, P3_DATAO_REG_27__SCAN_IN, P3_U6759);
  nand ginst29019 (P3_U6844, P3_EAX_REG_28__SCAN_IN, P3_U2447);
  nand ginst29020 (P3_U6845, P3_UWORD_REG_12__SCAN_IN, P3_U2410);
  nand ginst29021 (P3_U6846, P3_DATAO_REG_28__SCAN_IN, P3_U6759);
  nand ginst29022 (P3_U6847, P3_EAX_REG_29__SCAN_IN, P3_U2447);
  nand ginst29023 (P3_U6848, P3_UWORD_REG_13__SCAN_IN, P3_U2410);
  nand ginst29024 (P3_U6849, P3_DATAO_REG_29__SCAN_IN, P3_U6759);
  nand ginst29025 (P3_U6850, P3_EAX_REG_30__SCAN_IN, P3_U2447);
  nand ginst29026 (P3_U6851, P3_UWORD_REG_14__SCAN_IN, P3_U2410);
  nand ginst29027 (P3_U6852, P3_DATAO_REG_30__SCAN_IN, P3_U6759);
  nand ginst29028 (P3_U6853, P3_U2516, P3_U3243);
  nand ginst29029 (P3_U6854, BUF2_REG_0__SCAN_IN, P3_U2446);
  nand ginst29030 (P3_U6855, P3_U2411, P3_U2621);
  nand ginst29031 (P3_U6856, P3_ADD_546_U5, P3_U2400);
  nand ginst29032 (P3_U6857, P3_EAX_REG_0__SCAN_IN, P3_U3252);
  nand ginst29033 (P3_U6858, BUF2_REG_1__SCAN_IN, P3_U2446);
  nand ginst29034 (P3_U6859, P3_U2411, P3_U2622);
  nand ginst29035 (P3_U6860, P3_ADD_546_U71, P3_U2400);
  nand ginst29036 (P3_U6861, P3_EAX_REG_1__SCAN_IN, P3_U3252);
  nand ginst29037 (P3_U6862, BUF2_REG_2__SCAN_IN, P3_U2446);
  nand ginst29038 (P3_U6863, P3_U2411, P3_U2623);
  nand ginst29039 (P3_U6864, P3_ADD_546_U60, P3_U2400);
  nand ginst29040 (P3_U6865, P3_EAX_REG_2__SCAN_IN, P3_U3252);
  nand ginst29041 (P3_U6866, BUF2_REG_3__SCAN_IN, P3_U2446);
  nand ginst29042 (P3_U6867, P3_U2411, P3_U2624);
  nand ginst29043 (P3_U6868, P3_ADD_546_U57, P3_U2400);
  nand ginst29044 (P3_U6869, P3_EAX_REG_3__SCAN_IN, P3_U3252);
  nand ginst29045 (P3_U6870, BUF2_REG_4__SCAN_IN, P3_U2446);
  nand ginst29046 (P3_U6871, P3_U2411, P3_U2625);
  nand ginst29047 (P3_U6872, P3_ADD_546_U56, P3_U2400);
  nand ginst29048 (P3_U6873, P3_EAX_REG_4__SCAN_IN, P3_U3252);
  nand ginst29049 (P3_U6874, BUF2_REG_5__SCAN_IN, P3_U2446);
  nand ginst29050 (P3_U6875, P3_U2411, P3_U2626);
  nand ginst29051 (P3_U6876, P3_ADD_546_U55, P3_U2400);
  nand ginst29052 (P3_U6877, P3_EAX_REG_5__SCAN_IN, P3_U3252);
  nand ginst29053 (P3_U6878, BUF2_REG_6__SCAN_IN, P3_U2446);
  nand ginst29054 (P3_U6879, P3_U2411, P3_U2627);
  nand ginst29055 (P3_U6880, P3_ADD_546_U54, P3_U2400);
  nand ginst29056 (P3_U6881, P3_EAX_REG_6__SCAN_IN, P3_U3252);
  nand ginst29057 (P3_U6882, BUF2_REG_7__SCAN_IN, P3_U2446);
  nand ginst29058 (P3_U6883, P3_U2411, P3_U2628);
  nand ginst29059 (P3_U6884, P3_ADD_546_U53, P3_U2400);
  nand ginst29060 (P3_U6885, P3_EAX_REG_7__SCAN_IN, P3_U3252);
  nand ginst29061 (P3_U6886, BUF2_REG_8__SCAN_IN, P3_U2446);
  nand ginst29062 (P3_U6887, P3_U2411, P3_U2605);
  nand ginst29063 (P3_U6888, P3_ADD_546_U52, P3_U2400);
  nand ginst29064 (P3_U6889, P3_EAX_REG_8__SCAN_IN, P3_U3252);
  nand ginst29065 (P3_U6890, BUF2_REG_9__SCAN_IN, P3_U2446);
  nand ginst29066 (P3_U6891, P3_U2411, P3_U2606);
  nand ginst29067 (P3_U6892, P3_ADD_546_U51, P3_U2400);
  nand ginst29068 (P3_U6893, P3_EAX_REG_9__SCAN_IN, P3_U3252);
  nand ginst29069 (P3_U6894, BUF2_REG_10__SCAN_IN, P3_U2446);
  nand ginst29070 (P3_U6895, P3_U2411, P3_U2607);
  nand ginst29071 (P3_U6896, P3_ADD_546_U81, P3_U2400);
  nand ginst29072 (P3_U6897, P3_EAX_REG_10__SCAN_IN, P3_U3252);
  nand ginst29073 (P3_U6898, BUF2_REG_11__SCAN_IN, P3_U2446);
  nand ginst29074 (P3_U6899, P3_U2411, P3_U2608);
  nand ginst29075 (P3_U6900, P3_ADD_546_U80, P3_U2400);
  nand ginst29076 (P3_U6901, P3_EAX_REG_11__SCAN_IN, P3_U3252);
  nand ginst29077 (P3_U6902, BUF2_REG_12__SCAN_IN, P3_U2446);
  nand ginst29078 (P3_U6903, P3_U2411, P3_U2609);
  nand ginst29079 (P3_U6904, P3_ADD_546_U79, P3_U2400);
  nand ginst29080 (P3_U6905, P3_EAX_REG_12__SCAN_IN, P3_U3252);
  nand ginst29081 (P3_U6906, BUF2_REG_13__SCAN_IN, P3_U2446);
  nand ginst29082 (P3_U6907, P3_U2411, P3_U2610);
  nand ginst29083 (P3_U6908, P3_ADD_546_U78, P3_U2400);
  nand ginst29084 (P3_U6909, P3_EAX_REG_13__SCAN_IN, P3_U3252);
  nand ginst29085 (P3_U6910, BUF2_REG_14__SCAN_IN, P3_U2446);
  nand ginst29086 (P3_U6911, P3_U2411, P3_U2611);
  nand ginst29087 (P3_U6912, P3_ADD_546_U77, P3_U2400);
  nand ginst29088 (P3_U6913, P3_EAX_REG_14__SCAN_IN, P3_U3252);
  nand ginst29089 (P3_U6914, BUF2_REG_15__SCAN_IN, P3_U2446);
  nand ginst29090 (P3_U6915, P3_U2411, P3_U2612);
  nand ginst29091 (P3_U6916, P3_ADD_546_U76, P3_U2400);
  nand ginst29092 (P3_U6917, P3_EAX_REG_15__SCAN_IN, P3_U3252);
  nand ginst29093 (P3_U6918, BUF2_REG_0__SCAN_IN, P3_U2448);
  nand ginst29094 (P3_U6919, BUF2_REG_16__SCAN_IN, P3_U2444);
  nand ginst29095 (P3_U6920, P3_U2411, P3_U3062);
  nand ginst29096 (P3_U6921, P3_ADD_546_U75, P3_U2400);
  nand ginst29097 (P3_U6922, P3_EAX_REG_16__SCAN_IN, P3_U3252);
  nand ginst29098 (P3_U6923, BUF2_REG_1__SCAN_IN, P3_U2448);
  nand ginst29099 (P3_U6924, BUF2_REG_17__SCAN_IN, P3_U2444);
  nand ginst29100 (P3_U6925, P3_U2411, P3_U3063);
  nand ginst29101 (P3_U6926, P3_ADD_546_U74, P3_U2400);
  nand ginst29102 (P3_U6927, P3_EAX_REG_17__SCAN_IN, P3_U3252);
  nand ginst29103 (P3_U6928, BUF2_REG_2__SCAN_IN, P3_U2448);
  nand ginst29104 (P3_U6929, BUF2_REG_18__SCAN_IN, P3_U2444);
  nand ginst29105 (P3_U6930, P3_U2411, P3_U3064);
  nand ginst29106 (P3_U6931, P3_ADD_546_U73, P3_U2400);
  nand ginst29107 (P3_U6932, P3_EAX_REG_18__SCAN_IN, P3_U3252);
  nand ginst29108 (P3_U6933, BUF2_REG_3__SCAN_IN, P3_U2448);
  nand ginst29109 (P3_U6934, BUF2_REG_19__SCAN_IN, P3_U2444);
  nand ginst29110 (P3_U6935, P3_U2411, P3_U3065);
  nand ginst29111 (P3_U6936, P3_ADD_546_U72, P3_U2400);
  nand ginst29112 (P3_U6937, P3_EAX_REG_19__SCAN_IN, P3_U3252);
  nand ginst29113 (P3_U6938, BUF2_REG_4__SCAN_IN, P3_U2448);
  nand ginst29114 (P3_U6939, BUF2_REG_20__SCAN_IN, P3_U2444);
  nand ginst29115 (P3_U6940, P3_U2411, P3_U3066);
  nand ginst29116 (P3_U6941, P3_ADD_546_U70, P3_U2400);
  nand ginst29117 (P3_U6942, P3_EAX_REG_20__SCAN_IN, P3_U3252);
  nand ginst29118 (P3_U6943, BUF2_REG_5__SCAN_IN, P3_U2448);
  nand ginst29119 (P3_U6944, BUF2_REG_21__SCAN_IN, P3_U2444);
  nand ginst29120 (P3_U6945, P3_U2411, P3_U3067);
  nand ginst29121 (P3_U6946, P3_ADD_546_U69, P3_U2400);
  nand ginst29122 (P3_U6947, P3_EAX_REG_21__SCAN_IN, P3_U3252);
  nand ginst29123 (P3_U6948, BUF2_REG_6__SCAN_IN, P3_U2448);
  nand ginst29124 (P3_U6949, BUF2_REG_22__SCAN_IN, P3_U2444);
  nand ginst29125 (P3_U6950, P3_U2411, P3_U3068);
  nand ginst29126 (P3_U6951, P3_ADD_546_U68, P3_U2400);
  nand ginst29127 (P3_U6952, P3_EAX_REG_22__SCAN_IN, P3_U3252);
  nand ginst29128 (P3_U6953, BUF2_REG_7__SCAN_IN, P3_U2448);
  nand ginst29129 (P3_U6954, BUF2_REG_23__SCAN_IN, P3_U2444);
  nand ginst29130 (P3_U6955, P3_ADD_391_1180_U25, P3_U2411);
  nand ginst29131 (P3_U6956, P3_ADD_546_U67, P3_U2400);
  nand ginst29132 (P3_U6957, P3_EAX_REG_23__SCAN_IN, P3_U3252);
  nand ginst29133 (P3_U6958, BUF2_REG_8__SCAN_IN, P3_U2448);
  nand ginst29134 (P3_U6959, BUF2_REG_24__SCAN_IN, P3_U2444);
  nand ginst29135 (P3_U6960, P3_ADD_391_1180_U24, P3_U2411);
  nand ginst29136 (P3_U6961, P3_ADD_546_U66, P3_U2400);
  nand ginst29137 (P3_U6962, P3_EAX_REG_24__SCAN_IN, P3_U3252);
  nand ginst29138 (P3_U6963, BUF2_REG_9__SCAN_IN, P3_U2448);
  nand ginst29139 (P3_U6964, BUF2_REG_25__SCAN_IN, P3_U2444);
  nand ginst29140 (P3_U6965, P3_ADD_391_1180_U23, P3_U2411);
  nand ginst29141 (P3_U6966, P3_ADD_546_U65, P3_U2400);
  nand ginst29142 (P3_U6967, P3_EAX_REG_25__SCAN_IN, P3_U3252);
  nand ginst29143 (P3_U6968, BUF2_REG_10__SCAN_IN, P3_U2448);
  nand ginst29144 (P3_U6969, BUF2_REG_26__SCAN_IN, P3_U2444);
  nand ginst29145 (P3_U6970, P3_ADD_391_1180_U22, P3_U2411);
  nand ginst29146 (P3_U6971, P3_ADD_546_U64, P3_U2400);
  nand ginst29147 (P3_U6972, P3_EAX_REG_26__SCAN_IN, P3_U3252);
  nand ginst29148 (P3_U6973, BUF2_REG_11__SCAN_IN, P3_U2448);
  nand ginst29149 (P3_U6974, BUF2_REG_27__SCAN_IN, P3_U2444);
  nand ginst29150 (P3_U6975, P3_ADD_391_1180_U21, P3_U2411);
  nand ginst29151 (P3_U6976, P3_ADD_546_U63, P3_U2400);
  nand ginst29152 (P3_U6977, P3_EAX_REG_27__SCAN_IN, P3_U3252);
  nand ginst29153 (P3_U6978, BUF2_REG_12__SCAN_IN, P3_U2448);
  nand ginst29154 (P3_U6979, BUF2_REG_28__SCAN_IN, P3_U2444);
  nand ginst29155 (P3_U6980, P3_ADD_391_1180_U20, P3_U2411);
  nand ginst29156 (P3_U6981, P3_ADD_546_U62, P3_U2400);
  nand ginst29157 (P3_U6982, P3_EAX_REG_28__SCAN_IN, P3_U3252);
  nand ginst29158 (P3_U6983, BUF2_REG_13__SCAN_IN, P3_U2448);
  nand ginst29159 (P3_U6984, BUF2_REG_29__SCAN_IN, P3_U2444);
  nand ginst29160 (P3_U6985, P3_ADD_391_1180_U19, P3_U2411);
  nand ginst29161 (P3_U6986, P3_ADD_546_U61, P3_U2400);
  nand ginst29162 (P3_U6987, P3_EAX_REG_29__SCAN_IN, P3_U3252);
  nand ginst29163 (P3_U6988, BUF2_REG_14__SCAN_IN, P3_U2448);
  nand ginst29164 (P3_U6989, BUF2_REG_30__SCAN_IN, P3_U2444);
  nand ginst29165 (P3_U6990, P3_ADD_391_1180_U18, P3_U2411);
  nand ginst29166 (P3_U6991, P3_ADD_546_U59, P3_U2400);
  nand ginst29167 (P3_U6992, P3_EAX_REG_30__SCAN_IN, P3_U3252);
  nand ginst29168 (P3_U6993, BUF2_REG_31__SCAN_IN, P3_U2444);
  nand ginst29169 (P3_U6994, P3_ADD_546_U58, P3_U2400);
  nand ginst29170 (P3_U6995, P3_EAX_REG_31__SCAN_IN, P3_U3252);
  nand ginst29171 (P3_U6996, P3_GTE_401_U6, P3_U4305);
  nand ginst29172 (P3_U6997, P3_U3242, P3_U6996);
  nand ginst29173 (P3_U6998, P3_INSTQUEUE_REG_0__0__SCAN_IN, P3_U2408);
  nand ginst29174 (P3_U6999, P3_ADD_552_U5, P3_U2399);
  nand ginst29175 (P3_U7000, P3_EBX_REG_0__SCAN_IN, P3_U3253);
  nand ginst29176 (P3_U7001, P3_INSTQUEUE_REG_0__1__SCAN_IN, P3_U2408);
  nand ginst29177 (P3_U7002, P3_ADD_552_U71, P3_U2399);
  nand ginst29178 (P3_U7003, P3_EBX_REG_1__SCAN_IN, P3_U3253);
  nand ginst29179 (P3_U7004, P3_INSTQUEUE_REG_0__2__SCAN_IN, P3_U2408);
  nand ginst29180 (P3_U7005, P3_ADD_552_U60, P3_U2399);
  nand ginst29181 (P3_U7006, P3_EBX_REG_2__SCAN_IN, P3_U3253);
  nand ginst29182 (P3_U7007, P3_INSTQUEUE_REG_0__3__SCAN_IN, P3_U2408);
  nand ginst29183 (P3_U7008, P3_ADD_552_U57, P3_U2399);
  nand ginst29184 (P3_U7009, P3_EBX_REG_3__SCAN_IN, P3_U3253);
  nand ginst29185 (P3_U7010, P3_INSTQUEUE_REG_0__4__SCAN_IN, P3_U2408);
  nand ginst29186 (P3_U7011, P3_ADD_552_U56, P3_U2399);
  nand ginst29187 (P3_U7012, P3_EBX_REG_4__SCAN_IN, P3_U3253);
  nand ginst29188 (P3_U7013, P3_INSTQUEUE_REG_0__5__SCAN_IN, P3_U2408);
  nand ginst29189 (P3_U7014, P3_ADD_552_U55, P3_U2399);
  nand ginst29190 (P3_U7015, P3_EBX_REG_5__SCAN_IN, P3_U3253);
  nand ginst29191 (P3_U7016, P3_INSTQUEUE_REG_0__6__SCAN_IN, P3_U2408);
  nand ginst29192 (P3_U7017, P3_ADD_552_U54, P3_U2399);
  nand ginst29193 (P3_U7018, P3_EBX_REG_6__SCAN_IN, P3_U3253);
  nand ginst29194 (P3_U7019, P3_INSTQUEUE_REG_0__7__SCAN_IN, P3_U2408);
  nand ginst29195 (P3_U7020, P3_ADD_552_U53, P3_U2399);
  nand ginst29196 (P3_U7021, P3_EBX_REG_7__SCAN_IN, P3_U3253);
  nand ginst29197 (P3_U7022, P3_U2408, P3_U2605);
  nand ginst29198 (P3_U7023, P3_ADD_552_U52, P3_U2399);
  nand ginst29199 (P3_U7024, P3_EBX_REG_8__SCAN_IN, P3_U3253);
  nand ginst29200 (P3_U7025, P3_U2408, P3_U2606);
  nand ginst29201 (P3_U7026, P3_ADD_552_U51, P3_U2399);
  nand ginst29202 (P3_U7027, P3_EBX_REG_9__SCAN_IN, P3_U3253);
  nand ginst29203 (P3_U7028, P3_U2408, P3_U2607);
  nand ginst29204 (P3_U7029, P3_ADD_552_U81, P3_U2399);
  nand ginst29205 (P3_U7030, P3_EBX_REG_10__SCAN_IN, P3_U3253);
  nand ginst29206 (P3_U7031, P3_U2408, P3_U2608);
  nand ginst29207 (P3_U7032, P3_ADD_552_U80, P3_U2399);
  nand ginst29208 (P3_U7033, P3_EBX_REG_11__SCAN_IN, P3_U3253);
  nand ginst29209 (P3_U7034, P3_U2408, P3_U2609);
  nand ginst29210 (P3_U7035, P3_ADD_552_U79, P3_U2399);
  nand ginst29211 (P3_U7036, P3_EBX_REG_12__SCAN_IN, P3_U3253);
  nand ginst29212 (P3_U7037, P3_U2408, P3_U2610);
  nand ginst29213 (P3_U7038, P3_ADD_552_U78, P3_U2399);
  nand ginst29214 (P3_U7039, P3_EBX_REG_13__SCAN_IN, P3_U3253);
  nand ginst29215 (P3_U7040, P3_U2408, P3_U2611);
  nand ginst29216 (P3_U7041, P3_ADD_552_U77, P3_U2399);
  nand ginst29217 (P3_U7042, P3_EBX_REG_14__SCAN_IN, P3_U3253);
  nand ginst29218 (P3_U7043, P3_U2408, P3_U2612);
  nand ginst29219 (P3_U7044, P3_ADD_552_U76, P3_U2399);
  nand ginst29220 (P3_U7045, P3_EBX_REG_15__SCAN_IN, P3_U3253);
  nand ginst29221 (P3_U7046, P3_U2408, P3_U3062);
  nand ginst29222 (P3_U7047, P3_ADD_552_U75, P3_U2399);
  nand ginst29223 (P3_U7048, P3_EBX_REG_16__SCAN_IN, P3_U3253);
  nand ginst29224 (P3_U7049, P3_U2408, P3_U3063);
  nand ginst29225 (P3_U7050, P3_ADD_552_U74, P3_U2399);
  nand ginst29226 (P3_U7051, P3_EBX_REG_17__SCAN_IN, P3_U3253);
  nand ginst29227 (P3_U7052, P3_U2408, P3_U3064);
  nand ginst29228 (P3_U7053, P3_ADD_552_U73, P3_U2399);
  nand ginst29229 (P3_U7054, P3_EBX_REG_18__SCAN_IN, P3_U3253);
  nand ginst29230 (P3_U7055, P3_U2408, P3_U3065);
  nand ginst29231 (P3_U7056, P3_ADD_552_U72, P3_U2399);
  nand ginst29232 (P3_U7057, P3_EBX_REG_19__SCAN_IN, P3_U3253);
  nand ginst29233 (P3_U7058, P3_U2408, P3_U3066);
  nand ginst29234 (P3_U7059, P3_ADD_552_U70, P3_U2399);
  nand ginst29235 (P3_U7060, P3_EBX_REG_20__SCAN_IN, P3_U3253);
  nand ginst29236 (P3_U7061, P3_U2408, P3_U3067);
  nand ginst29237 (P3_U7062, P3_ADD_552_U69, P3_U2399);
  nand ginst29238 (P3_U7063, P3_EBX_REG_21__SCAN_IN, P3_U3253);
  nand ginst29239 (P3_U7064, P3_U2408, P3_U3068);
  nand ginst29240 (P3_U7065, P3_ADD_552_U68, P3_U2399);
  nand ginst29241 (P3_U7066, P3_EBX_REG_22__SCAN_IN, P3_U3253);
  nand ginst29242 (P3_U7067, P3_ADD_402_1132_U25, P3_U2408);
  nand ginst29243 (P3_U7068, P3_ADD_552_U67, P3_U2399);
  nand ginst29244 (P3_U7069, P3_EBX_REG_23__SCAN_IN, P3_U3253);
  nand ginst29245 (P3_U7070, P3_ADD_402_1132_U24, P3_U2408);
  nand ginst29246 (P3_U7071, P3_ADD_552_U66, P3_U2399);
  nand ginst29247 (P3_U7072, P3_EBX_REG_24__SCAN_IN, P3_U3253);
  nand ginst29248 (P3_U7073, P3_ADD_402_1132_U23, P3_U2408);
  nand ginst29249 (P3_U7074, P3_ADD_552_U65, P3_U2399);
  nand ginst29250 (P3_U7075, P3_EBX_REG_25__SCAN_IN, P3_U3253);
  nand ginst29251 (P3_U7076, P3_ADD_402_1132_U22, P3_U2408);
  nand ginst29252 (P3_U7077, P3_ADD_552_U64, P3_U2399);
  nand ginst29253 (P3_U7078, P3_EBX_REG_26__SCAN_IN, P3_U3253);
  nand ginst29254 (P3_U7079, P3_ADD_402_1132_U21, P3_U2408);
  nand ginst29255 (P3_U7080, P3_ADD_552_U63, P3_U2399);
  nand ginst29256 (P3_U7081, P3_EBX_REG_27__SCAN_IN, P3_U3253);
  nand ginst29257 (P3_U7082, P3_ADD_402_1132_U20, P3_U2408);
  nand ginst29258 (P3_U7083, P3_ADD_552_U62, P3_U2399);
  nand ginst29259 (P3_U7084, P3_EBX_REG_28__SCAN_IN, P3_U3253);
  nand ginst29260 (P3_U7085, P3_ADD_402_1132_U19, P3_U2408);
  nand ginst29261 (P3_U7086, P3_ADD_552_U61, P3_U2399);
  nand ginst29262 (P3_U7087, P3_EBX_REG_29__SCAN_IN, P3_U3253);
  nand ginst29263 (P3_U7088, P3_ADD_402_1132_U18, P3_U2408);
  nand ginst29264 (P3_U7089, P3_ADD_552_U59, P3_U2399);
  nand ginst29265 (P3_U7090, P3_EBX_REG_30__SCAN_IN, P3_U3253);
  nand ginst29266 (P3_U7091, P3_ADD_552_U58, P3_U2399);
  nand ginst29267 (P3_U7092, P3_EBX_REG_31__SCAN_IN, P3_U3253);
  nand ginst29268 (P3_U7093, P3_U5488, P3_U5491);
  not ginst29269 (P3_U7094, P3_U3260);
  not ginst29270 (P3_U7095, P3_U3257);
  or ginst29271 (P3_U7096, P3_STATEBS16_REG_SCAN_IN, U209);
  nand ginst29272 (P3_U7097, P3_EBX_REG_0__SCAN_IN, P3_U2602);
  nand ginst29273 (P3_U7098, P3_REIP_REG_0__SCAN_IN, P3_U2601);
  nand ginst29274 (P3_U7099, P3_EBX_REG_0__SCAN_IN, P3_U7910);
  nand ginst29275 (P3_U7100, P3_ADD_505_U5, P3_U2455);
  nand ginst29276 (P3_U7101, P3_ADD_486_U5, P3_U2454);
  nand ginst29277 (P3_U7102, P3_REIP_REG_0__SCAN_IN, P3_U2405);
  nand ginst29278 (P3_U7103, P3_PHYADDRPOINTER_REG_0__SCAN_IN, P3_U2403);
  nand ginst29279 (P3_U7104, P3_PHYADDRPOINTER_REG_0__SCAN_IN, P3_U4319);
  nand ginst29280 (P3_U7105, P3_PHYADDRPOINTER_REG_0__SCAN_IN, P3_U2401);
  nand ginst29281 (P3_U7106, P3_REIP_REG_0__SCAN_IN, P3_U7094);
  nand ginst29282 (P3_U7107, P3_SUB_414_U50, P3_U2602);
  nand ginst29283 (P3_U7108, P3_ADD_467_U4, P3_U2601);
  nand ginst29284 (P3_U7109, P3_EBX_REG_1__SCAN_IN, P3_U7910);
  nand ginst29285 (P3_U7110, P3_ADD_505_U17, P3_U2455);
  nand ginst29286 (P3_U7111, P3_ADD_486_U17, P3_U2454);
  nand ginst29287 (P3_U7112, P3_ADD_430_U4, P3_U2405);
  nand ginst29288 (P3_U7113, P3_ADD_318_U4, P3_U2403);
  nand ginst29289 (P3_U7114, P3_SUB_320_U50, P3_U4319);
  nand ginst29290 (P3_U7115, P3_PHYADDRPOINTER_REG_1__SCAN_IN, P3_U2401);
  nand ginst29291 (P3_U7116, P3_REIP_REG_1__SCAN_IN, P3_U7094);
  nand ginst29292 (P3_U7117, P3_SUB_414_U17, P3_U2602);
  nand ginst29293 (P3_U7118, P3_ADD_467_U71, P3_U2601);
  nand ginst29294 (P3_U7119, P3_EBX_REG_2__SCAN_IN, P3_U7910);
  nand ginst29295 (P3_U7120, P3_ADD_505_U16, P3_U2455);
  nand ginst29296 (P3_U7121, P3_ADD_486_U16, P3_U2454);
  nand ginst29297 (P3_U7122, P3_ADD_430_U71, P3_U2405);
  nand ginst29298 (P3_U7123, P3_ADD_318_U71, P3_U2403);
  nand ginst29299 (P3_U7124, P3_SUB_320_U17, P3_U4319);
  nand ginst29300 (P3_U7125, P3_PHYADDRPOINTER_REG_2__SCAN_IN, P3_U2401);
  nand ginst29301 (P3_U7126, P3_REIP_REG_2__SCAN_IN, P3_U7094);
  nand ginst29302 (P3_U7127, P3_SUB_414_U59, P3_U2602);
  nand ginst29303 (P3_U7128, P3_ADD_467_U68, P3_U2601);
  nand ginst29304 (P3_U7129, P3_EBX_REG_3__SCAN_IN, P3_U7910);
  nand ginst29305 (P3_U7130, P3_ADD_505_U15, P3_U2455);
  nand ginst29306 (P3_U7131, P3_ADD_486_U15, P3_U2454);
  nand ginst29307 (P3_U7132, P3_ADD_430_U68, P3_U2405);
  nand ginst29308 (P3_U7133, P3_ADD_318_U68, P3_U2403);
  nand ginst29309 (P3_U7134, P3_SUB_320_U59, P3_U4319);
  nand ginst29310 (P3_U7135, P3_PHYADDRPOINTER_REG_3__SCAN_IN, P3_U2401);
  nand ginst29311 (P3_U7136, P3_REIP_REG_3__SCAN_IN, P3_U7094);
  nand ginst29312 (P3_U7137, P3_SUB_414_U18, P3_U2602);
  nand ginst29313 (P3_U7138, P3_ADD_467_U67, P3_U2601);
  nand ginst29314 (P3_U7139, P3_EBX_REG_4__SCAN_IN, P3_U7910);
  nand ginst29315 (P3_U7140, P3_ADD_505_U14, P3_U2455);
  nand ginst29316 (P3_U7141, P3_ADD_486_U14, P3_U2454);
  nand ginst29317 (P3_U7142, P3_ADD_430_U67, P3_U2405);
  nand ginst29318 (P3_U7143, P3_ADD_318_U67, P3_U2403);
  nand ginst29319 (P3_U7144, P3_SUB_320_U18, P3_U4319);
  nand ginst29320 (P3_U7145, P3_PHYADDRPOINTER_REG_4__SCAN_IN, P3_U2401);
  nand ginst29321 (P3_U7146, P3_REIP_REG_4__SCAN_IN, P3_U7094);
  nand ginst29322 (P3_U7147, P3_SUB_414_U57, P3_U2602);
  nand ginst29323 (P3_U7148, P3_ADD_467_U66, P3_U2601);
  nand ginst29324 (P3_U7149, P3_EBX_REG_5__SCAN_IN, P3_U7910);
  nand ginst29325 (P3_U7150, P3_ADD_505_U6, P3_U2455);
  nand ginst29326 (P3_U7151, P3_ADD_486_U6, P3_U2454);
  nand ginst29327 (P3_U7152, P3_ADD_430_U66, P3_U2405);
  nand ginst29328 (P3_U7153, P3_ADD_318_U66, P3_U2403);
  nand ginst29329 (P3_U7154, P3_SUB_320_U57, P3_U4319);
  nand ginst29330 (P3_U7155, P3_PHYADDRPOINTER_REG_5__SCAN_IN, P3_U2401);
  nand ginst29331 (P3_U7156, P3_REIP_REG_5__SCAN_IN, P3_U7094);
  nand ginst29332 (P3_U7157, P3_SUB_414_U19, P3_U2602);
  nand ginst29333 (P3_U7158, P3_ADD_467_U65, P3_U2601);
  nand ginst29334 (P3_U7159, P3_EBX_REG_6__SCAN_IN, P3_U7910);
  nand ginst29335 (P3_U7160, P3_ADD_430_U65, P3_U2405);
  nand ginst29336 (P3_U7161, P3_ADD_318_U65, P3_U2403);
  nand ginst29337 (P3_U7162, P3_SUB_320_U19, P3_U4319);
  nand ginst29338 (P3_U7163, P3_PHYADDRPOINTER_REG_6__SCAN_IN, P3_U2401);
  nand ginst29339 (P3_U7164, P3_REIP_REG_6__SCAN_IN, P3_U7094);
  nand ginst29340 (P3_U7165, P3_SUB_414_U55, P3_U2602);
  nand ginst29341 (P3_U7166, P3_ADD_467_U64, P3_U2601);
  nand ginst29342 (P3_U7167, P3_EBX_REG_7__SCAN_IN, P3_U7910);
  nand ginst29343 (P3_U7168, P3_ADD_430_U64, P3_U2405);
  nand ginst29344 (P3_U7169, P3_ADD_318_U64, P3_U2403);
  nand ginst29345 (P3_U7170, P3_SUB_320_U55, P3_U4319);
  nand ginst29346 (P3_U7171, P3_PHYADDRPOINTER_REG_7__SCAN_IN, P3_U2401);
  nand ginst29347 (P3_U7172, P3_REIP_REG_7__SCAN_IN, P3_U7094);
  nand ginst29348 (P3_U7173, P3_SUB_414_U20, P3_U2602);
  nand ginst29349 (P3_U7174, P3_ADD_467_U63, P3_U2601);
  nand ginst29350 (P3_U7175, P3_EBX_REG_8__SCAN_IN, P3_U7910);
  nand ginst29351 (P3_U7176, P3_ADD_430_U63, P3_U2405);
  nand ginst29352 (P3_U7177, P3_ADD_318_U63, P3_U2403);
  nand ginst29353 (P3_U7178, P3_SUB_320_U20, P3_U4319);
  nand ginst29354 (P3_U7179, P3_PHYADDRPOINTER_REG_8__SCAN_IN, P3_U2401);
  nand ginst29355 (P3_U7180, P3_REIP_REG_8__SCAN_IN, P3_U7094);
  nand ginst29356 (P3_U7181, P3_SUB_414_U53, P3_U2602);
  nand ginst29357 (P3_U7182, P3_ADD_467_U62, P3_U2601);
  nand ginst29358 (P3_U7183, P3_EBX_REG_9__SCAN_IN, P3_U7910);
  nand ginst29359 (P3_U7184, P3_ADD_430_U62, P3_U2405);
  nand ginst29360 (P3_U7185, P3_ADD_318_U62, P3_U2403);
  nand ginst29361 (P3_U7186, P3_SUB_320_U53, P3_U4319);
  nand ginst29362 (P3_U7187, P3_PHYADDRPOINTER_REG_9__SCAN_IN, P3_U2401);
  nand ginst29363 (P3_U7188, P3_REIP_REG_9__SCAN_IN, P3_U7094);
  nand ginst29364 (P3_U7189, P3_SUB_414_U6, P3_U2602);
  nand ginst29365 (P3_U7190, P3_ADD_467_U91, P3_U2601);
  nand ginst29366 (P3_U7191, P3_EBX_REG_10__SCAN_IN, P3_U7910);
  nand ginst29367 (P3_U7192, P3_ADD_430_U91, P3_U2405);
  nand ginst29368 (P3_U7193, P3_ADD_318_U91, P3_U2403);
  nand ginst29369 (P3_U7194, P3_SUB_320_U6, P3_U4319);
  nand ginst29370 (P3_U7195, P3_PHYADDRPOINTER_REG_10__SCAN_IN, P3_U2401);
  nand ginst29371 (P3_U7196, P3_REIP_REG_10__SCAN_IN, P3_U7094);
  nand ginst29372 (P3_U7197, P3_SUB_414_U82, P3_U2602);
  nand ginst29373 (P3_U7198, P3_ADD_467_U90, P3_U2601);
  nand ginst29374 (P3_U7199, P3_EBX_REG_11__SCAN_IN, P3_U7910);
  nand ginst29375 (P3_U7200, P3_ADD_430_U90, P3_U2405);
  nand ginst29376 (P3_U7201, P3_ADD_318_U90, P3_U2403);
  nand ginst29377 (P3_U7202, P3_SUB_320_U82, P3_U4319);
  nand ginst29378 (P3_U7203, P3_PHYADDRPOINTER_REG_11__SCAN_IN, P3_U2401);
  nand ginst29379 (P3_U7204, P3_REIP_REG_11__SCAN_IN, P3_U7094);
  nand ginst29380 (P3_U7205, P3_SUB_414_U7, P3_U2602);
  nand ginst29381 (P3_U7206, P3_ADD_467_U89, P3_U2601);
  nand ginst29382 (P3_U7207, P3_EBX_REG_12__SCAN_IN, P3_U7910);
  nand ginst29383 (P3_U7208, P3_ADD_430_U89, P3_U2405);
  nand ginst29384 (P3_U7209, P3_ADD_318_U89, P3_U2403);
  nand ginst29385 (P3_U7210, P3_SUB_320_U7, P3_U4319);
  nand ginst29386 (P3_U7211, P3_PHYADDRPOINTER_REG_12__SCAN_IN, P3_U2401);
  nand ginst29387 (P3_U7212, P3_REIP_REG_12__SCAN_IN, P3_U7094);
  nand ginst29388 (P3_U7213, P3_SUB_414_U80, P3_U2602);
  nand ginst29389 (P3_U7214, P3_ADD_467_U88, P3_U2601);
  nand ginst29390 (P3_U7215, P3_EBX_REG_13__SCAN_IN, P3_U7910);
  nand ginst29391 (P3_U7216, P3_ADD_430_U88, P3_U2405);
  nand ginst29392 (P3_U7217, P3_ADD_318_U88, P3_U2403);
  nand ginst29393 (P3_U7218, P3_SUB_320_U80, P3_U4319);
  nand ginst29394 (P3_U7219, P3_PHYADDRPOINTER_REG_13__SCAN_IN, P3_U2401);
  nand ginst29395 (P3_U7220, P3_REIP_REG_13__SCAN_IN, P3_U7094);
  nand ginst29396 (P3_U7221, P3_SUB_414_U8, P3_U2602);
  nand ginst29397 (P3_U7222, P3_ADD_467_U87, P3_U2601);
  nand ginst29398 (P3_U7223, P3_EBX_REG_14__SCAN_IN, P3_U7910);
  nand ginst29399 (P3_U7224, P3_ADD_430_U87, P3_U2405);
  nand ginst29400 (P3_U7225, P3_ADD_318_U87, P3_U2403);
  nand ginst29401 (P3_U7226, P3_SUB_320_U8, P3_U4319);
  nand ginst29402 (P3_U7227, P3_PHYADDRPOINTER_REG_14__SCAN_IN, P3_U2401);
  nand ginst29403 (P3_U7228, P3_REIP_REG_14__SCAN_IN, P3_U7094);
  nand ginst29404 (P3_U7229, P3_SUB_414_U78, P3_U2602);
  nand ginst29405 (P3_U7230, P3_ADD_467_U86, P3_U2601);
  nand ginst29406 (P3_U7231, P3_EBX_REG_15__SCAN_IN, P3_U7910);
  nand ginst29407 (P3_U7232, P3_ADD_430_U86, P3_U2405);
  nand ginst29408 (P3_U7233, P3_ADD_318_U86, P3_U2403);
  nand ginst29409 (P3_U7234, P3_SUB_320_U78, P3_U4319);
  nand ginst29410 (P3_U7235, P3_PHYADDRPOINTER_REG_15__SCAN_IN, P3_U2401);
  nand ginst29411 (P3_U7236, P3_REIP_REG_15__SCAN_IN, P3_U7094);
  nand ginst29412 (P3_U7237, P3_SUB_414_U9, P3_U2602);
  nand ginst29413 (P3_U7238, P3_ADD_467_U85, P3_U2601);
  nand ginst29414 (P3_U7239, P3_EBX_REG_16__SCAN_IN, P3_U7910);
  nand ginst29415 (P3_U7240, P3_ADD_430_U85, P3_U2405);
  nand ginst29416 (P3_U7241, P3_ADD_318_U85, P3_U2403);
  nand ginst29417 (P3_U7242, P3_SUB_320_U9, P3_U4319);
  nand ginst29418 (P3_U7243, P3_PHYADDRPOINTER_REG_16__SCAN_IN, P3_U2401);
  nand ginst29419 (P3_U7244, P3_REIP_REG_16__SCAN_IN, P3_U7094);
  nand ginst29420 (P3_U7245, P3_SUB_414_U76, P3_U2602);
  nand ginst29421 (P3_U7246, P3_ADD_467_U84, P3_U2601);
  nand ginst29422 (P3_U7247, P3_EBX_REG_17__SCAN_IN, P3_U7910);
  nand ginst29423 (P3_U7248, P3_ADD_430_U84, P3_U2405);
  nand ginst29424 (P3_U7249, P3_ADD_318_U84, P3_U2403);
  nand ginst29425 (P3_U7250, P3_SUB_320_U76, P3_U4319);
  nand ginst29426 (P3_U7251, P3_PHYADDRPOINTER_REG_17__SCAN_IN, P3_U2401);
  nand ginst29427 (P3_U7252, P3_REIP_REG_17__SCAN_IN, P3_U7094);
  nand ginst29428 (P3_U7253, P3_SUB_414_U10, P3_U2602);
  nand ginst29429 (P3_U7254, P3_ADD_467_U83, P3_U2601);
  nand ginst29430 (P3_U7255, P3_EBX_REG_18__SCAN_IN, P3_U7910);
  nand ginst29431 (P3_U7256, P3_ADD_430_U83, P3_U2405);
  nand ginst29432 (P3_U7257, P3_ADD_318_U83, P3_U2403);
  nand ginst29433 (P3_U7258, P3_SUB_320_U10, P3_U4319);
  nand ginst29434 (P3_U7259, P3_PHYADDRPOINTER_REG_18__SCAN_IN, P3_U2401);
  nand ginst29435 (P3_U7260, P3_REIP_REG_18__SCAN_IN, P3_U7094);
  nand ginst29436 (P3_U7261, P3_SUB_414_U74, P3_U2602);
  nand ginst29437 (P3_U7262, P3_ADD_467_U82, P3_U2601);
  nand ginst29438 (P3_U7263, P3_EBX_REG_19__SCAN_IN, P3_U7910);
  nand ginst29439 (P3_U7264, P3_ADD_430_U82, P3_U2405);
  nand ginst29440 (P3_U7265, P3_ADD_318_U82, P3_U2403);
  nand ginst29441 (P3_U7266, P3_SUB_320_U74, P3_U4319);
  nand ginst29442 (P3_U7267, P3_PHYADDRPOINTER_REG_19__SCAN_IN, P3_U2401);
  nand ginst29443 (P3_U7268, P3_REIP_REG_19__SCAN_IN, P3_U7094);
  nand ginst29444 (P3_U7269, P3_SUB_414_U11, P3_U2602);
  nand ginst29445 (P3_U7270, P3_ADD_467_U81, P3_U2601);
  nand ginst29446 (P3_U7271, P3_EBX_REG_20__SCAN_IN, P3_U7910);
  nand ginst29447 (P3_U7272, P3_ADD_430_U81, P3_U2405);
  nand ginst29448 (P3_U7273, P3_ADD_318_U81, P3_U2403);
  nand ginst29449 (P3_U7274, P3_SUB_320_U11, P3_U4319);
  nand ginst29450 (P3_U7275, P3_PHYADDRPOINTER_REG_20__SCAN_IN, P3_U2401);
  nand ginst29451 (P3_U7276, P3_REIP_REG_20__SCAN_IN, P3_U7094);
  nand ginst29452 (P3_U7277, P3_SUB_414_U70, P3_U2602);
  nand ginst29453 (P3_U7278, P3_ADD_467_U80, P3_U2601);
  nand ginst29454 (P3_U7279, P3_EBX_REG_21__SCAN_IN, P3_U7910);
  nand ginst29455 (P3_U7280, P3_ADD_430_U80, P3_U2405);
  nand ginst29456 (P3_U7281, P3_ADD_318_U80, P3_U2403);
  nand ginst29457 (P3_U7282, P3_SUB_320_U70, P3_U4319);
  nand ginst29458 (P3_U7283, P3_PHYADDRPOINTER_REG_21__SCAN_IN, P3_U2401);
  nand ginst29459 (P3_U7284, P3_REIP_REG_21__SCAN_IN, P3_U7094);
  nand ginst29460 (P3_U7285, P3_SUB_414_U12, P3_U2602);
  nand ginst29461 (P3_U7286, P3_ADD_467_U79, P3_U2601);
  nand ginst29462 (P3_U7287, P3_EBX_REG_22__SCAN_IN, P3_U7910);
  nand ginst29463 (P3_U7288, P3_ADD_430_U79, P3_U2405);
  nand ginst29464 (P3_U7289, P3_ADD_318_U79, P3_U2403);
  nand ginst29465 (P3_U7290, P3_SUB_320_U12, P3_U4319);
  nand ginst29466 (P3_U7291, P3_PHYADDRPOINTER_REG_22__SCAN_IN, P3_U2401);
  nand ginst29467 (P3_U7292, P3_REIP_REG_22__SCAN_IN, P3_U7094);
  nand ginst29468 (P3_U7293, P3_SUB_414_U68, P3_U2602);
  nand ginst29469 (P3_U7294, P3_ADD_467_U78, P3_U2601);
  nand ginst29470 (P3_U7295, P3_EBX_REG_23__SCAN_IN, P3_U7910);
  nand ginst29471 (P3_U7296, P3_ADD_430_U78, P3_U2405);
  nand ginst29472 (P3_U7297, P3_ADD_318_U78, P3_U2403);
  nand ginst29473 (P3_U7298, P3_SUB_320_U68, P3_U4319);
  nand ginst29474 (P3_U7299, P3_PHYADDRPOINTER_REG_23__SCAN_IN, P3_U2401);
  nand ginst29475 (P3_U7300, P3_REIP_REG_23__SCAN_IN, P3_U7094);
  nand ginst29476 (P3_U7301, P3_SUB_414_U13, P3_U2602);
  nand ginst29477 (P3_U7302, P3_ADD_467_U77, P3_U2601);
  nand ginst29478 (P3_U7303, P3_EBX_REG_24__SCAN_IN, P3_U7910);
  nand ginst29479 (P3_U7304, P3_ADD_430_U77, P3_U2405);
  nand ginst29480 (P3_U7305, P3_ADD_318_U77, P3_U2403);
  nand ginst29481 (P3_U7306, P3_SUB_320_U13, P3_U4319);
  nand ginst29482 (P3_U7307, P3_PHYADDRPOINTER_REG_24__SCAN_IN, P3_U2401);
  nand ginst29483 (P3_U7308, P3_REIP_REG_24__SCAN_IN, P3_U7094);
  nand ginst29484 (P3_U7309, P3_SUB_414_U66, P3_U2602);
  nand ginst29485 (P3_U7310, P3_ADD_467_U76, P3_U2601);
  nand ginst29486 (P3_U7311, P3_EBX_REG_25__SCAN_IN, P3_U7910);
  nand ginst29487 (P3_U7312, P3_ADD_430_U76, P3_U2405);
  nand ginst29488 (P3_U7313, P3_ADD_318_U76, P3_U2403);
  nand ginst29489 (P3_U7314, P3_SUB_320_U66, P3_U4319);
  nand ginst29490 (P3_U7315, P3_PHYADDRPOINTER_REG_25__SCAN_IN, P3_U2401);
  nand ginst29491 (P3_U7316, P3_REIP_REG_25__SCAN_IN, P3_U7094);
  nand ginst29492 (P3_U7317, P3_SUB_414_U14, P3_U2602);
  nand ginst29493 (P3_U7318, P3_ADD_467_U75, P3_U2601);
  nand ginst29494 (P3_U7319, P3_EBX_REG_26__SCAN_IN, P3_U7910);
  nand ginst29495 (P3_U7320, P3_ADD_430_U75, P3_U2405);
  nand ginst29496 (P3_U7321, P3_ADD_318_U75, P3_U2403);
  nand ginst29497 (P3_U7322, P3_SUB_320_U14, P3_U4319);
  nand ginst29498 (P3_U7323, P3_PHYADDRPOINTER_REG_26__SCAN_IN, P3_U2401);
  nand ginst29499 (P3_U7324, P3_REIP_REG_26__SCAN_IN, P3_U7094);
  nand ginst29500 (P3_U7325, P3_SUB_414_U64, P3_U2602);
  nand ginst29501 (P3_U7326, P3_ADD_467_U74, P3_U2601);
  nand ginst29502 (P3_U7327, P3_EBX_REG_27__SCAN_IN, P3_U7910);
  nand ginst29503 (P3_U7328, P3_ADD_430_U74, P3_U2405);
  nand ginst29504 (P3_U7329, P3_ADD_318_U74, P3_U2403);
  nand ginst29505 (P3_U7330, P3_SUB_320_U64, P3_U4319);
  nand ginst29506 (P3_U7331, P3_PHYADDRPOINTER_REG_27__SCAN_IN, P3_U2401);
  nand ginst29507 (P3_U7332, P3_REIP_REG_27__SCAN_IN, P3_U7094);
  nand ginst29508 (P3_U7333, P3_SUB_414_U15, P3_U2602);
  nand ginst29509 (P3_U7334, P3_ADD_467_U73, P3_U2601);
  nand ginst29510 (P3_U7335, P3_EBX_REG_28__SCAN_IN, P3_U7910);
  nand ginst29511 (P3_U7336, P3_ADD_430_U73, P3_U2405);
  nand ginst29512 (P3_U7337, P3_ADD_318_U73, P3_U2403);
  nand ginst29513 (P3_U7338, P3_SUB_320_U15, P3_U4319);
  nand ginst29514 (P3_U7339, P3_PHYADDRPOINTER_REG_28__SCAN_IN, P3_U2401);
  nand ginst29515 (P3_U7340, P3_REIP_REG_28__SCAN_IN, P3_U7094);
  nand ginst29516 (P3_U7341, P3_SUB_414_U16, P3_U2602);
  nand ginst29517 (P3_U7342, P3_ADD_467_U72, P3_U2601);
  nand ginst29518 (P3_U7343, P3_EBX_REG_29__SCAN_IN, P3_U7910);
  nand ginst29519 (P3_U7344, P3_ADD_430_U72, P3_U2405);
  nand ginst29520 (P3_U7345, P3_ADD_318_U72, P3_U2403);
  nand ginst29521 (P3_U7346, P3_SUB_320_U16, P3_U4319);
  nand ginst29522 (P3_U7347, P3_PHYADDRPOINTER_REG_29__SCAN_IN, P3_U2401);
  nand ginst29523 (P3_U7348, P3_REIP_REG_29__SCAN_IN, P3_U7094);
  nand ginst29524 (P3_U7349, P3_SUB_414_U62, P3_U2602);
  nand ginst29525 (P3_U7350, P3_ADD_467_U70, P3_U2601);
  nand ginst29526 (P3_U7351, P3_EBX_REG_30__SCAN_IN, P3_U7910);
  nand ginst29527 (P3_U7352, P3_ADD_430_U70, P3_U2405);
  nand ginst29528 (P3_U7353, P3_ADD_318_U70, P3_U2403);
  nand ginst29529 (P3_U7354, P3_SUB_320_U62, P3_U4319);
  nand ginst29530 (P3_U7355, P3_PHYADDRPOINTER_REG_30__SCAN_IN, P3_U2401);
  nand ginst29531 (P3_U7356, P3_REIP_REG_30__SCAN_IN, P3_U7094);
  nand ginst29532 (P3_U7357, P3_U2603, P3_U4135);
  nand ginst29533 (P3_U7358, P3_SUB_414_U51, P3_U2602);
  nand ginst29534 (P3_U7359, P3_ADD_467_U69, P3_U2601);
  nand ginst29535 (P3_U7360, P3_EBX_REG_31__SCAN_IN, P3_U7910);
  nand ginst29536 (P3_U7361, P3_ADD_430_U69, P3_U2405);
  nand ginst29537 (P3_U7362, P3_ADD_318_U69, P3_U2403);
  not ginst29538 (P3_U7363, P3_U7362);
  nand ginst29539 (P3_U7364, P3_PHYADDRPOINTER_REG_31__SCAN_IN, P3_U2401);
  nand ginst29540 (P3_U7365, P3_REIP_REG_31__SCAN_IN, P3_U7094);
  nand ginst29541 (P3_U7366, P3_DATAWIDTH_REG_0__SCAN_IN, P3_DATAWIDTH_REG_1__SCAN_IN);
  or ginst29542 (P3_U7367, P3_REIP_REG_0__SCAN_IN, P3_REIP_REG_1__SCAN_IN);
  not ginst29543 (P3_U7368, P3_U4285);
  nand ginst29544 (P3_U7369, P3_FLUSH_REG_SCAN_IN, P3_U4285);
  nand ginst29545 (P3_U7370, P3_U2390, P3_U4623);
  nand ginst29546 (P3_U7371, P3_U2453, P3_U2630);
  nand ginst29547 (P3_U7372, P3_U3123, P3_U7371);
  nand ginst29548 (P3_U7373, P3_U3121, P3_U7372);
  not ginst29549 (P3_U7374, P3_U4287);
  nand ginst29550 (P3_U7375, P3_U2631, P3_U4296);
  nand ginst29551 (P3_U7376, P3_U3112, P3_U3118);
  nand ginst29552 (P3_U7377, P3_STATE2_REG_2__SCAN_IN, P3_U4150, P3_U7919);
  nand ginst29553 (P3_U7378, P3_STATE2_REG_0__SCAN_IN, P3_U7377);
  nand ginst29554 (P3_U7379, P3_U3125, P3_U7378);
  nand ginst29555 (P3_U7380, P3_U2390, P3_U2604);
  nand ginst29556 (P3_U7381, P3_CODEFETCH_REG_SCAN_IN, P3_U7380);
  nand ginst29557 (P3_U7382, P3_STATE2_REG_0__SCAN_IN, P3_U4347);
  nand ginst29558 (P3_U7383, P3_STATE_REG_0__SCAN_IN, P3_ADS_N_REG_SCAN_IN);
  not ginst29559 (P3_U7384, P3_U4288);
  nand ginst29560 (P3_U7385, P3_STATE2_REG_2__SCAN_IN, P3_U3111, P3_U3114);
  nand ginst29561 (P3_U7386, P3_STATE2_REG_2__SCAN_IN, P3_U4488);
  nand ginst29562 (P3_U7387, P3_INSTQUEUE_REG_15__7__SCAN_IN, P3_U2542);
  nand ginst29563 (P3_U7388, P3_INSTQUEUE_REG_14__7__SCAN_IN, P3_U2541);
  nand ginst29564 (P3_U7389, P3_INSTQUEUE_REG_13__7__SCAN_IN, P3_U2540);
  nand ginst29565 (P3_U7390, P3_INSTQUEUE_REG_12__7__SCAN_IN, P3_U2539);
  nand ginst29566 (P3_U7391, P3_INSTQUEUE_REG_11__7__SCAN_IN, P3_U2537);
  nand ginst29567 (P3_U7392, P3_INSTQUEUE_REG_10__7__SCAN_IN, P3_U2536);
  nand ginst29568 (P3_U7393, P3_INSTQUEUE_REG_9__7__SCAN_IN, P3_U2535);
  nand ginst29569 (P3_U7394, P3_INSTQUEUE_REG_8__7__SCAN_IN, P3_U2534);
  nand ginst29570 (P3_U7395, P3_INSTQUEUE_REG_7__7__SCAN_IN, P3_U2532);
  nand ginst29571 (P3_U7396, P3_INSTQUEUE_REG_6__7__SCAN_IN, P3_U2531);
  nand ginst29572 (P3_U7397, P3_INSTQUEUE_REG_5__7__SCAN_IN, P3_U2530);
  nand ginst29573 (P3_U7398, P3_INSTQUEUE_REG_4__7__SCAN_IN, P3_U2529);
  nand ginst29574 (P3_U7399, P3_INSTQUEUE_REG_3__7__SCAN_IN, P3_U2527);
  nand ginst29575 (P3_U7400, P3_INSTQUEUE_REG_2__7__SCAN_IN, P3_U2525);
  nand ginst29576 (P3_U7401, P3_INSTQUEUE_REG_1__7__SCAN_IN, P3_U2523);
  nand ginst29577 (P3_U7402, P3_INSTQUEUE_REG_0__7__SCAN_IN, P3_U2521);
  nand ginst29578 (P3_U7403, P3_INSTQUEUE_REG_15__6__SCAN_IN, P3_U2542);
  nand ginst29579 (P3_U7404, P3_INSTQUEUE_REG_14__6__SCAN_IN, P3_U2541);
  nand ginst29580 (P3_U7405, P3_INSTQUEUE_REG_13__6__SCAN_IN, P3_U2540);
  nand ginst29581 (P3_U7406, P3_INSTQUEUE_REG_12__6__SCAN_IN, P3_U2539);
  nand ginst29582 (P3_U7407, P3_INSTQUEUE_REG_11__6__SCAN_IN, P3_U2537);
  nand ginst29583 (P3_U7408, P3_INSTQUEUE_REG_10__6__SCAN_IN, P3_U2536);
  nand ginst29584 (P3_U7409, P3_INSTQUEUE_REG_9__6__SCAN_IN, P3_U2535);
  nand ginst29585 (P3_U7410, P3_INSTQUEUE_REG_8__6__SCAN_IN, P3_U2534);
  nand ginst29586 (P3_U7411, P3_INSTQUEUE_REG_7__6__SCAN_IN, P3_U2532);
  nand ginst29587 (P3_U7412, P3_INSTQUEUE_REG_6__6__SCAN_IN, P3_U2531);
  nand ginst29588 (P3_U7413, P3_INSTQUEUE_REG_5__6__SCAN_IN, P3_U2530);
  nand ginst29589 (P3_U7414, P3_INSTQUEUE_REG_4__6__SCAN_IN, P3_U2529);
  nand ginst29590 (P3_U7415, P3_INSTQUEUE_REG_3__6__SCAN_IN, P3_U2527);
  nand ginst29591 (P3_U7416, P3_INSTQUEUE_REG_2__6__SCAN_IN, P3_U2525);
  nand ginst29592 (P3_U7417, P3_INSTQUEUE_REG_1__6__SCAN_IN, P3_U2523);
  nand ginst29593 (P3_U7418, P3_INSTQUEUE_REG_0__6__SCAN_IN, P3_U2521);
  nand ginst29594 (P3_U7419, P3_INSTQUEUE_REG_15__5__SCAN_IN, P3_U2542);
  nand ginst29595 (P3_U7420, P3_INSTQUEUE_REG_14__5__SCAN_IN, P3_U2541);
  nand ginst29596 (P3_U7421, P3_INSTQUEUE_REG_13__5__SCAN_IN, P3_U2540);
  nand ginst29597 (P3_U7422, P3_INSTQUEUE_REG_12__5__SCAN_IN, P3_U2539);
  nand ginst29598 (P3_U7423, P3_INSTQUEUE_REG_11__5__SCAN_IN, P3_U2537);
  nand ginst29599 (P3_U7424, P3_INSTQUEUE_REG_10__5__SCAN_IN, P3_U2536);
  nand ginst29600 (P3_U7425, P3_INSTQUEUE_REG_9__5__SCAN_IN, P3_U2535);
  nand ginst29601 (P3_U7426, P3_INSTQUEUE_REG_8__5__SCAN_IN, P3_U2534);
  nand ginst29602 (P3_U7427, P3_INSTQUEUE_REG_7__5__SCAN_IN, P3_U2532);
  nand ginst29603 (P3_U7428, P3_INSTQUEUE_REG_6__5__SCAN_IN, P3_U2531);
  nand ginst29604 (P3_U7429, P3_INSTQUEUE_REG_5__5__SCAN_IN, P3_U2530);
  nand ginst29605 (P3_U7430, P3_INSTQUEUE_REG_4__5__SCAN_IN, P3_U2529);
  nand ginst29606 (P3_U7431, P3_INSTQUEUE_REG_3__5__SCAN_IN, P3_U2527);
  nand ginst29607 (P3_U7432, P3_INSTQUEUE_REG_2__5__SCAN_IN, P3_U2525);
  nand ginst29608 (P3_U7433, P3_INSTQUEUE_REG_1__5__SCAN_IN, P3_U2523);
  nand ginst29609 (P3_U7434, P3_INSTQUEUE_REG_0__5__SCAN_IN, P3_U2521);
  nand ginst29610 (P3_U7435, P3_INSTQUEUE_REG_15__4__SCAN_IN, P3_U2542);
  nand ginst29611 (P3_U7436, P3_INSTQUEUE_REG_14__4__SCAN_IN, P3_U2541);
  nand ginst29612 (P3_U7437, P3_INSTQUEUE_REG_13__4__SCAN_IN, P3_U2540);
  nand ginst29613 (P3_U7438, P3_INSTQUEUE_REG_12__4__SCAN_IN, P3_U2539);
  nand ginst29614 (P3_U7439, P3_INSTQUEUE_REG_11__4__SCAN_IN, P3_U2537);
  nand ginst29615 (P3_U7440, P3_INSTQUEUE_REG_10__4__SCAN_IN, P3_U2536);
  nand ginst29616 (P3_U7441, P3_INSTQUEUE_REG_9__4__SCAN_IN, P3_U2535);
  nand ginst29617 (P3_U7442, P3_INSTQUEUE_REG_8__4__SCAN_IN, P3_U2534);
  nand ginst29618 (P3_U7443, P3_INSTQUEUE_REG_7__4__SCAN_IN, P3_U2532);
  nand ginst29619 (P3_U7444, P3_INSTQUEUE_REG_6__4__SCAN_IN, P3_U2531);
  nand ginst29620 (P3_U7445, P3_INSTQUEUE_REG_5__4__SCAN_IN, P3_U2530);
  nand ginst29621 (P3_U7446, P3_INSTQUEUE_REG_4__4__SCAN_IN, P3_U2529);
  nand ginst29622 (P3_U7447, P3_INSTQUEUE_REG_3__4__SCAN_IN, P3_U2527);
  nand ginst29623 (P3_U7448, P3_INSTQUEUE_REG_2__4__SCAN_IN, P3_U2525);
  nand ginst29624 (P3_U7449, P3_INSTQUEUE_REG_1__4__SCAN_IN, P3_U2523);
  nand ginst29625 (P3_U7450, P3_INSTQUEUE_REG_0__4__SCAN_IN, P3_U2521);
  nand ginst29626 (P3_U7451, P3_INSTQUEUE_REG_15__3__SCAN_IN, P3_U2542);
  nand ginst29627 (P3_U7452, P3_INSTQUEUE_REG_14__3__SCAN_IN, P3_U2541);
  nand ginst29628 (P3_U7453, P3_INSTQUEUE_REG_13__3__SCAN_IN, P3_U2540);
  nand ginst29629 (P3_U7454, P3_INSTQUEUE_REG_12__3__SCAN_IN, P3_U2539);
  nand ginst29630 (P3_U7455, P3_INSTQUEUE_REG_11__3__SCAN_IN, P3_U2537);
  nand ginst29631 (P3_U7456, P3_INSTQUEUE_REG_10__3__SCAN_IN, P3_U2536);
  nand ginst29632 (P3_U7457, P3_INSTQUEUE_REG_9__3__SCAN_IN, P3_U2535);
  nand ginst29633 (P3_U7458, P3_INSTQUEUE_REG_8__3__SCAN_IN, P3_U2534);
  nand ginst29634 (P3_U7459, P3_INSTQUEUE_REG_7__3__SCAN_IN, P3_U2532);
  nand ginst29635 (P3_U7460, P3_INSTQUEUE_REG_6__3__SCAN_IN, P3_U2531);
  nand ginst29636 (P3_U7461, P3_INSTQUEUE_REG_5__3__SCAN_IN, P3_U2530);
  nand ginst29637 (P3_U7462, P3_INSTQUEUE_REG_4__3__SCAN_IN, P3_U2529);
  nand ginst29638 (P3_U7463, P3_INSTQUEUE_REG_3__3__SCAN_IN, P3_U2527);
  nand ginst29639 (P3_U7464, P3_INSTQUEUE_REG_2__3__SCAN_IN, P3_U2525);
  nand ginst29640 (P3_U7465, P3_INSTQUEUE_REG_1__3__SCAN_IN, P3_U2523);
  nand ginst29641 (P3_U7466, P3_INSTQUEUE_REG_0__3__SCAN_IN, P3_U2521);
  nand ginst29642 (P3_U7467, P3_INSTQUEUE_REG_15__2__SCAN_IN, P3_U2542);
  nand ginst29643 (P3_U7468, P3_INSTQUEUE_REG_14__2__SCAN_IN, P3_U2541);
  nand ginst29644 (P3_U7469, P3_INSTQUEUE_REG_13__2__SCAN_IN, P3_U2540);
  nand ginst29645 (P3_U7470, P3_INSTQUEUE_REG_12__2__SCAN_IN, P3_U2539);
  nand ginst29646 (P3_U7471, P3_INSTQUEUE_REG_11__2__SCAN_IN, P3_U2537);
  nand ginst29647 (P3_U7472, P3_INSTQUEUE_REG_10__2__SCAN_IN, P3_U2536);
  nand ginst29648 (P3_U7473, P3_INSTQUEUE_REG_9__2__SCAN_IN, P3_U2535);
  nand ginst29649 (P3_U7474, P3_INSTQUEUE_REG_8__2__SCAN_IN, P3_U2534);
  nand ginst29650 (P3_U7475, P3_INSTQUEUE_REG_7__2__SCAN_IN, P3_U2532);
  nand ginst29651 (P3_U7476, P3_INSTQUEUE_REG_6__2__SCAN_IN, P3_U2531);
  nand ginst29652 (P3_U7477, P3_INSTQUEUE_REG_5__2__SCAN_IN, P3_U2530);
  nand ginst29653 (P3_U7478, P3_INSTQUEUE_REG_4__2__SCAN_IN, P3_U2529);
  nand ginst29654 (P3_U7479, P3_INSTQUEUE_REG_3__2__SCAN_IN, P3_U2527);
  nand ginst29655 (P3_U7480, P3_INSTQUEUE_REG_2__2__SCAN_IN, P3_U2525);
  nand ginst29656 (P3_U7481, P3_INSTQUEUE_REG_1__2__SCAN_IN, P3_U2523);
  nand ginst29657 (P3_U7482, P3_INSTQUEUE_REG_0__2__SCAN_IN, P3_U2521);
  nand ginst29658 (P3_U7483, P3_INSTQUEUE_REG_15__1__SCAN_IN, P3_U2542);
  nand ginst29659 (P3_U7484, P3_INSTQUEUE_REG_14__1__SCAN_IN, P3_U2541);
  nand ginst29660 (P3_U7485, P3_INSTQUEUE_REG_13__1__SCAN_IN, P3_U2540);
  nand ginst29661 (P3_U7486, P3_INSTQUEUE_REG_12__1__SCAN_IN, P3_U2539);
  nand ginst29662 (P3_U7487, P3_INSTQUEUE_REG_11__1__SCAN_IN, P3_U2537);
  nand ginst29663 (P3_U7488, P3_INSTQUEUE_REG_10__1__SCAN_IN, P3_U2536);
  nand ginst29664 (P3_U7489, P3_INSTQUEUE_REG_9__1__SCAN_IN, P3_U2535);
  nand ginst29665 (P3_U7490, P3_INSTQUEUE_REG_8__1__SCAN_IN, P3_U2534);
  nand ginst29666 (P3_U7491, P3_INSTQUEUE_REG_7__1__SCAN_IN, P3_U2532);
  nand ginst29667 (P3_U7492, P3_INSTQUEUE_REG_6__1__SCAN_IN, P3_U2531);
  nand ginst29668 (P3_U7493, P3_INSTQUEUE_REG_5__1__SCAN_IN, P3_U2530);
  nand ginst29669 (P3_U7494, P3_INSTQUEUE_REG_4__1__SCAN_IN, P3_U2529);
  nand ginst29670 (P3_U7495, P3_INSTQUEUE_REG_3__1__SCAN_IN, P3_U2527);
  nand ginst29671 (P3_U7496, P3_INSTQUEUE_REG_2__1__SCAN_IN, P3_U2525);
  nand ginst29672 (P3_U7497, P3_INSTQUEUE_REG_1__1__SCAN_IN, P3_U2523);
  nand ginst29673 (P3_U7498, P3_INSTQUEUE_REG_0__1__SCAN_IN, P3_U2521);
  nand ginst29674 (P3_U7499, P3_INSTQUEUE_REG_15__0__SCAN_IN, P3_U2542);
  nand ginst29675 (P3_U7500, P3_INSTQUEUE_REG_14__0__SCAN_IN, P3_U2541);
  nand ginst29676 (P3_U7501, P3_INSTQUEUE_REG_13__0__SCAN_IN, P3_U2540);
  nand ginst29677 (P3_U7502, P3_INSTQUEUE_REG_12__0__SCAN_IN, P3_U2539);
  nand ginst29678 (P3_U7503, P3_INSTQUEUE_REG_11__0__SCAN_IN, P3_U2537);
  nand ginst29679 (P3_U7504, P3_INSTQUEUE_REG_10__0__SCAN_IN, P3_U2536);
  nand ginst29680 (P3_U7505, P3_INSTQUEUE_REG_9__0__SCAN_IN, P3_U2535);
  nand ginst29681 (P3_U7506, P3_INSTQUEUE_REG_8__0__SCAN_IN, P3_U2534);
  nand ginst29682 (P3_U7507, P3_INSTQUEUE_REG_7__0__SCAN_IN, P3_U2532);
  nand ginst29683 (P3_U7508, P3_INSTQUEUE_REG_6__0__SCAN_IN, P3_U2531);
  nand ginst29684 (P3_U7509, P3_INSTQUEUE_REG_5__0__SCAN_IN, P3_U2530);
  nand ginst29685 (P3_U7510, P3_INSTQUEUE_REG_4__0__SCAN_IN, P3_U2529);
  nand ginst29686 (P3_U7511, P3_INSTQUEUE_REG_3__0__SCAN_IN, P3_U2527);
  nand ginst29687 (P3_U7512, P3_INSTQUEUE_REG_2__0__SCAN_IN, P3_U2525);
  nand ginst29688 (P3_U7513, P3_INSTQUEUE_REG_1__0__SCAN_IN, P3_U2523);
  nand ginst29689 (P3_U7514, P3_INSTQUEUE_REG_0__0__SCAN_IN, P3_U2521);
  nand ginst29690 (P3_U7515, P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P3_U4470);
  not ginst29691 (P3_U7516, P3_U3266);
  nand ginst29692 (P3_U7517, P3_INSTQUEUE_REG_0__7__SCAN_IN, P3_U2562);
  nand ginst29693 (P3_U7518, P3_INSTQUEUE_REG_1__7__SCAN_IN, P3_U2561);
  nand ginst29694 (P3_U7519, P3_INSTQUEUE_REG_2__7__SCAN_IN, P3_U2560);
  nand ginst29695 (P3_U7520, P3_INSTQUEUE_REG_3__7__SCAN_IN, P3_U2559);
  nand ginst29696 (P3_U7521, P3_INSTQUEUE_REG_4__7__SCAN_IN, P3_U2557);
  nand ginst29697 (P3_U7522, P3_INSTQUEUE_REG_5__7__SCAN_IN, P3_U2556);
  nand ginst29698 (P3_U7523, P3_INSTQUEUE_REG_6__7__SCAN_IN, P3_U2555);
  nand ginst29699 (P3_U7524, P3_INSTQUEUE_REG_7__7__SCAN_IN, P3_U2554);
  nand ginst29700 (P3_U7525, P3_INSTQUEUE_REG_8__7__SCAN_IN, P3_U2552);
  nand ginst29701 (P3_U7526, P3_INSTQUEUE_REG_9__7__SCAN_IN, P3_U2551);
  nand ginst29702 (P3_U7527, P3_INSTQUEUE_REG_10__7__SCAN_IN, P3_U2550);
  nand ginst29703 (P3_U7528, P3_INSTQUEUE_REG_11__7__SCAN_IN, P3_U2549);
  nand ginst29704 (P3_U7529, P3_INSTQUEUE_REG_12__7__SCAN_IN, P3_U2547);
  nand ginst29705 (P3_U7530, P3_INSTQUEUE_REG_13__7__SCAN_IN, P3_U2546);
  nand ginst29706 (P3_U7531, P3_INSTQUEUE_REG_14__7__SCAN_IN, P3_U2545);
  nand ginst29707 (P3_U7532, P3_INSTQUEUE_REG_15__7__SCAN_IN, P3_U2544);
  nand ginst29708 (P3_U7533, P3_INSTQUEUE_REG_0__6__SCAN_IN, P3_U2562);
  nand ginst29709 (P3_U7534, P3_INSTQUEUE_REG_1__6__SCAN_IN, P3_U2561);
  nand ginst29710 (P3_U7535, P3_INSTQUEUE_REG_2__6__SCAN_IN, P3_U2560);
  nand ginst29711 (P3_U7536, P3_INSTQUEUE_REG_3__6__SCAN_IN, P3_U2559);
  nand ginst29712 (P3_U7537, P3_INSTQUEUE_REG_4__6__SCAN_IN, P3_U2557);
  nand ginst29713 (P3_U7538, P3_INSTQUEUE_REG_5__6__SCAN_IN, P3_U2556);
  nand ginst29714 (P3_U7539, P3_INSTQUEUE_REG_6__6__SCAN_IN, P3_U2555);
  nand ginst29715 (P3_U7540, P3_INSTQUEUE_REG_7__6__SCAN_IN, P3_U2554);
  nand ginst29716 (P3_U7541, P3_INSTQUEUE_REG_8__6__SCAN_IN, P3_U2552);
  nand ginst29717 (P3_U7542, P3_INSTQUEUE_REG_9__6__SCAN_IN, P3_U2551);
  nand ginst29718 (P3_U7543, P3_INSTQUEUE_REG_10__6__SCAN_IN, P3_U2550);
  nand ginst29719 (P3_U7544, P3_INSTQUEUE_REG_11__6__SCAN_IN, P3_U2549);
  nand ginst29720 (P3_U7545, P3_INSTQUEUE_REG_12__6__SCAN_IN, P3_U2547);
  nand ginst29721 (P3_U7546, P3_INSTQUEUE_REG_13__6__SCAN_IN, P3_U2546);
  nand ginst29722 (P3_U7547, P3_INSTQUEUE_REG_14__6__SCAN_IN, P3_U2545);
  nand ginst29723 (P3_U7548, P3_INSTQUEUE_REG_15__6__SCAN_IN, P3_U2544);
  nand ginst29724 (P3_U7549, P3_INSTQUEUE_REG_0__5__SCAN_IN, P3_U2562);
  nand ginst29725 (P3_U7550, P3_INSTQUEUE_REG_1__5__SCAN_IN, P3_U2561);
  nand ginst29726 (P3_U7551, P3_INSTQUEUE_REG_2__5__SCAN_IN, P3_U2560);
  nand ginst29727 (P3_U7552, P3_INSTQUEUE_REG_3__5__SCAN_IN, P3_U2559);
  nand ginst29728 (P3_U7553, P3_INSTQUEUE_REG_4__5__SCAN_IN, P3_U2557);
  nand ginst29729 (P3_U7554, P3_INSTQUEUE_REG_5__5__SCAN_IN, P3_U2556);
  nand ginst29730 (P3_U7555, P3_INSTQUEUE_REG_6__5__SCAN_IN, P3_U2555);
  nand ginst29731 (P3_U7556, P3_INSTQUEUE_REG_7__5__SCAN_IN, P3_U2554);
  nand ginst29732 (P3_U7557, P3_INSTQUEUE_REG_8__5__SCAN_IN, P3_U2552);
  nand ginst29733 (P3_U7558, P3_INSTQUEUE_REG_9__5__SCAN_IN, P3_U2551);
  nand ginst29734 (P3_U7559, P3_INSTQUEUE_REG_10__5__SCAN_IN, P3_U2550);
  nand ginst29735 (P3_U7560, P3_INSTQUEUE_REG_11__5__SCAN_IN, P3_U2549);
  nand ginst29736 (P3_U7561, P3_INSTQUEUE_REG_12__5__SCAN_IN, P3_U2547);
  nand ginst29737 (P3_U7562, P3_INSTQUEUE_REG_13__5__SCAN_IN, P3_U2546);
  nand ginst29738 (P3_U7563, P3_INSTQUEUE_REG_14__5__SCAN_IN, P3_U2545);
  nand ginst29739 (P3_U7564, P3_INSTQUEUE_REG_15__5__SCAN_IN, P3_U2544);
  nand ginst29740 (P3_U7565, P3_INSTQUEUE_REG_0__4__SCAN_IN, P3_U2562);
  nand ginst29741 (P3_U7566, P3_INSTQUEUE_REG_1__4__SCAN_IN, P3_U2561);
  nand ginst29742 (P3_U7567, P3_INSTQUEUE_REG_2__4__SCAN_IN, P3_U2560);
  nand ginst29743 (P3_U7568, P3_INSTQUEUE_REG_3__4__SCAN_IN, P3_U2559);
  nand ginst29744 (P3_U7569, P3_INSTQUEUE_REG_4__4__SCAN_IN, P3_U2557);
  nand ginst29745 (P3_U7570, P3_INSTQUEUE_REG_5__4__SCAN_IN, P3_U2556);
  nand ginst29746 (P3_U7571, P3_INSTQUEUE_REG_6__4__SCAN_IN, P3_U2555);
  nand ginst29747 (P3_U7572, P3_INSTQUEUE_REG_7__4__SCAN_IN, P3_U2554);
  nand ginst29748 (P3_U7573, P3_INSTQUEUE_REG_8__4__SCAN_IN, P3_U2552);
  nand ginst29749 (P3_U7574, P3_INSTQUEUE_REG_9__4__SCAN_IN, P3_U2551);
  nand ginst29750 (P3_U7575, P3_INSTQUEUE_REG_10__4__SCAN_IN, P3_U2550);
  nand ginst29751 (P3_U7576, P3_INSTQUEUE_REG_11__4__SCAN_IN, P3_U2549);
  nand ginst29752 (P3_U7577, P3_INSTQUEUE_REG_12__4__SCAN_IN, P3_U2547);
  nand ginst29753 (P3_U7578, P3_INSTQUEUE_REG_13__4__SCAN_IN, P3_U2546);
  nand ginst29754 (P3_U7579, P3_INSTQUEUE_REG_14__4__SCAN_IN, P3_U2545);
  nand ginst29755 (P3_U7580, P3_INSTQUEUE_REG_15__4__SCAN_IN, P3_U2544);
  nand ginst29756 (P3_U7581, P3_INSTQUEUE_REG_0__3__SCAN_IN, P3_U2562);
  nand ginst29757 (P3_U7582, P3_INSTQUEUE_REG_1__3__SCAN_IN, P3_U2561);
  nand ginst29758 (P3_U7583, P3_INSTQUEUE_REG_2__3__SCAN_IN, P3_U2560);
  nand ginst29759 (P3_U7584, P3_INSTQUEUE_REG_3__3__SCAN_IN, P3_U2559);
  nand ginst29760 (P3_U7585, P3_INSTQUEUE_REG_4__3__SCAN_IN, P3_U2557);
  nand ginst29761 (P3_U7586, P3_INSTQUEUE_REG_5__3__SCAN_IN, P3_U2556);
  nand ginst29762 (P3_U7587, P3_INSTQUEUE_REG_6__3__SCAN_IN, P3_U2555);
  nand ginst29763 (P3_U7588, P3_INSTQUEUE_REG_7__3__SCAN_IN, P3_U2554);
  nand ginst29764 (P3_U7589, P3_INSTQUEUE_REG_8__3__SCAN_IN, P3_U2552);
  nand ginst29765 (P3_U7590, P3_INSTQUEUE_REG_9__3__SCAN_IN, P3_U2551);
  nand ginst29766 (P3_U7591, P3_INSTQUEUE_REG_10__3__SCAN_IN, P3_U2550);
  nand ginst29767 (P3_U7592, P3_INSTQUEUE_REG_11__3__SCAN_IN, P3_U2549);
  nand ginst29768 (P3_U7593, P3_INSTQUEUE_REG_12__3__SCAN_IN, P3_U2547);
  nand ginst29769 (P3_U7594, P3_INSTQUEUE_REG_13__3__SCAN_IN, P3_U2546);
  nand ginst29770 (P3_U7595, P3_INSTQUEUE_REG_14__3__SCAN_IN, P3_U2545);
  nand ginst29771 (P3_U7596, P3_INSTQUEUE_REG_15__3__SCAN_IN, P3_U2544);
  nand ginst29772 (P3_U7597, P3_INSTQUEUE_REG_0__2__SCAN_IN, P3_U2562);
  nand ginst29773 (P3_U7598, P3_INSTQUEUE_REG_1__2__SCAN_IN, P3_U2561);
  nand ginst29774 (P3_U7599, P3_INSTQUEUE_REG_2__2__SCAN_IN, P3_U2560);
  nand ginst29775 (P3_U7600, P3_INSTQUEUE_REG_3__2__SCAN_IN, P3_U2559);
  nand ginst29776 (P3_U7601, P3_INSTQUEUE_REG_4__2__SCAN_IN, P3_U2557);
  nand ginst29777 (P3_U7602, P3_INSTQUEUE_REG_5__2__SCAN_IN, P3_U2556);
  nand ginst29778 (P3_U7603, P3_INSTQUEUE_REG_6__2__SCAN_IN, P3_U2555);
  nand ginst29779 (P3_U7604, P3_INSTQUEUE_REG_7__2__SCAN_IN, P3_U2554);
  nand ginst29780 (P3_U7605, P3_INSTQUEUE_REG_8__2__SCAN_IN, P3_U2552);
  nand ginst29781 (P3_U7606, P3_INSTQUEUE_REG_9__2__SCAN_IN, P3_U2551);
  nand ginst29782 (P3_U7607, P3_INSTQUEUE_REG_10__2__SCAN_IN, P3_U2550);
  nand ginst29783 (P3_U7608, P3_INSTQUEUE_REG_11__2__SCAN_IN, P3_U2549);
  nand ginst29784 (P3_U7609, P3_INSTQUEUE_REG_12__2__SCAN_IN, P3_U2547);
  nand ginst29785 (P3_U7610, P3_INSTQUEUE_REG_13__2__SCAN_IN, P3_U2546);
  nand ginst29786 (P3_U7611, P3_INSTQUEUE_REG_14__2__SCAN_IN, P3_U2545);
  nand ginst29787 (P3_U7612, P3_INSTQUEUE_REG_15__2__SCAN_IN, P3_U2544);
  nand ginst29788 (P3_U7613, P3_INSTQUEUE_REG_0__1__SCAN_IN, P3_U2562);
  nand ginst29789 (P3_U7614, P3_INSTQUEUE_REG_1__1__SCAN_IN, P3_U2561);
  nand ginst29790 (P3_U7615, P3_INSTQUEUE_REG_2__1__SCAN_IN, P3_U2560);
  nand ginst29791 (P3_U7616, P3_INSTQUEUE_REG_3__1__SCAN_IN, P3_U2559);
  nand ginst29792 (P3_U7617, P3_INSTQUEUE_REG_4__1__SCAN_IN, P3_U2557);
  nand ginst29793 (P3_U7618, P3_INSTQUEUE_REG_5__1__SCAN_IN, P3_U2556);
  nand ginst29794 (P3_U7619, P3_INSTQUEUE_REG_6__1__SCAN_IN, P3_U2555);
  nand ginst29795 (P3_U7620, P3_INSTQUEUE_REG_7__1__SCAN_IN, P3_U2554);
  nand ginst29796 (P3_U7621, P3_INSTQUEUE_REG_8__1__SCAN_IN, P3_U2552);
  nand ginst29797 (P3_U7622, P3_INSTQUEUE_REG_9__1__SCAN_IN, P3_U2551);
  nand ginst29798 (P3_U7623, P3_INSTQUEUE_REG_10__1__SCAN_IN, P3_U2550);
  nand ginst29799 (P3_U7624, P3_INSTQUEUE_REG_11__1__SCAN_IN, P3_U2549);
  nand ginst29800 (P3_U7625, P3_INSTQUEUE_REG_12__1__SCAN_IN, P3_U2547);
  nand ginst29801 (P3_U7626, P3_INSTQUEUE_REG_13__1__SCAN_IN, P3_U2546);
  nand ginst29802 (P3_U7627, P3_INSTQUEUE_REG_14__1__SCAN_IN, P3_U2545);
  nand ginst29803 (P3_U7628, P3_INSTQUEUE_REG_15__1__SCAN_IN, P3_U2544);
  nand ginst29804 (P3_U7629, P3_INSTQUEUE_REG_0__0__SCAN_IN, P3_U2562);
  nand ginst29805 (P3_U7630, P3_INSTQUEUE_REG_1__0__SCAN_IN, P3_U2561);
  nand ginst29806 (P3_U7631, P3_INSTQUEUE_REG_2__0__SCAN_IN, P3_U2560);
  nand ginst29807 (P3_U7632, P3_INSTQUEUE_REG_3__0__SCAN_IN, P3_U2559);
  nand ginst29808 (P3_U7633, P3_INSTQUEUE_REG_4__0__SCAN_IN, P3_U2557);
  nand ginst29809 (P3_U7634, P3_INSTQUEUE_REG_5__0__SCAN_IN, P3_U2556);
  nand ginst29810 (P3_U7635, P3_INSTQUEUE_REG_6__0__SCAN_IN, P3_U2555);
  nand ginst29811 (P3_U7636, P3_INSTQUEUE_REG_7__0__SCAN_IN, P3_U2554);
  nand ginst29812 (P3_U7637, P3_INSTQUEUE_REG_8__0__SCAN_IN, P3_U2552);
  nand ginst29813 (P3_U7638, P3_INSTQUEUE_REG_9__0__SCAN_IN, P3_U2551);
  nand ginst29814 (P3_U7639, P3_INSTQUEUE_REG_10__0__SCAN_IN, P3_U2550);
  nand ginst29815 (P3_U7640, P3_INSTQUEUE_REG_11__0__SCAN_IN, P3_U2549);
  nand ginst29816 (P3_U7641, P3_INSTQUEUE_REG_12__0__SCAN_IN, P3_U2547);
  nand ginst29817 (P3_U7642, P3_INSTQUEUE_REG_13__0__SCAN_IN, P3_U2546);
  nand ginst29818 (P3_U7643, P3_INSTQUEUE_REG_14__0__SCAN_IN, P3_U2545);
  nand ginst29819 (P3_U7644, P3_INSTQUEUE_REG_15__0__SCAN_IN, P3_U2544);
  not ginst29820 (P3_U7645, P3_U4289);
  nand ginst29821 (P3_U7646, P3_INSTQUEUE_REG_8__7__SCAN_IN, P3_U2582);
  nand ginst29822 (P3_U7647, P3_INSTQUEUE_REG_9__7__SCAN_IN, P3_U2581);
  nand ginst29823 (P3_U7648, P3_INSTQUEUE_REG_10__7__SCAN_IN, P3_U2580);
  nand ginst29824 (P3_U7649, P3_INSTQUEUE_REG_11__7__SCAN_IN, P3_U2579);
  nand ginst29825 (P3_U7650, P3_INSTQUEUE_REG_12__7__SCAN_IN, P3_U2577);
  nand ginst29826 (P3_U7651, P3_INSTQUEUE_REG_13__7__SCAN_IN, P3_U2576);
  nand ginst29827 (P3_U7652, P3_INSTQUEUE_REG_14__7__SCAN_IN, P3_U2575);
  nand ginst29828 (P3_U7653, P3_INSTQUEUE_REG_15__7__SCAN_IN, P3_U2574);
  nand ginst29829 (P3_U7654, P3_INSTQUEUE_REG_0__7__SCAN_IN, P3_U2572);
  nand ginst29830 (P3_U7655, P3_INSTQUEUE_REG_1__7__SCAN_IN, P3_U2571);
  nand ginst29831 (P3_U7656, P3_INSTQUEUE_REG_2__7__SCAN_IN, P3_U2570);
  nand ginst29832 (P3_U7657, P3_INSTQUEUE_REG_3__7__SCAN_IN, P3_U2569);
  nand ginst29833 (P3_U7658, P3_INSTQUEUE_REG_4__7__SCAN_IN, P3_U2567);
  nand ginst29834 (P3_U7659, P3_INSTQUEUE_REG_5__7__SCAN_IN, P3_U2566);
  nand ginst29835 (P3_U7660, P3_INSTQUEUE_REG_6__7__SCAN_IN, P3_U2565);
  nand ginst29836 (P3_U7661, P3_INSTQUEUE_REG_7__7__SCAN_IN, P3_U2564);
  nand ginst29837 (P3_U7662, P3_INSTQUEUE_REG_8__6__SCAN_IN, P3_U2582);
  nand ginst29838 (P3_U7663, P3_INSTQUEUE_REG_9__6__SCAN_IN, P3_U2581);
  nand ginst29839 (P3_U7664, P3_INSTQUEUE_REG_10__6__SCAN_IN, P3_U2580);
  nand ginst29840 (P3_U7665, P3_INSTQUEUE_REG_11__6__SCAN_IN, P3_U2579);
  nand ginst29841 (P3_U7666, P3_INSTQUEUE_REG_12__6__SCAN_IN, P3_U2577);
  nand ginst29842 (P3_U7667, P3_INSTQUEUE_REG_13__6__SCAN_IN, P3_U2576);
  nand ginst29843 (P3_U7668, P3_INSTQUEUE_REG_14__6__SCAN_IN, P3_U2575);
  nand ginst29844 (P3_U7669, P3_INSTQUEUE_REG_15__6__SCAN_IN, P3_U2574);
  nand ginst29845 (P3_U7670, P3_INSTQUEUE_REG_0__6__SCAN_IN, P3_U2572);
  nand ginst29846 (P3_U7671, P3_INSTQUEUE_REG_1__6__SCAN_IN, P3_U2571);
  nand ginst29847 (P3_U7672, P3_INSTQUEUE_REG_2__6__SCAN_IN, P3_U2570);
  nand ginst29848 (P3_U7673, P3_INSTQUEUE_REG_3__6__SCAN_IN, P3_U2569);
  nand ginst29849 (P3_U7674, P3_INSTQUEUE_REG_4__6__SCAN_IN, P3_U2567);
  nand ginst29850 (P3_U7675, P3_INSTQUEUE_REG_5__6__SCAN_IN, P3_U2566);
  nand ginst29851 (P3_U7676, P3_INSTQUEUE_REG_6__6__SCAN_IN, P3_U2565);
  nand ginst29852 (P3_U7677, P3_INSTQUEUE_REG_7__6__SCAN_IN, P3_U2564);
  nand ginst29853 (P3_U7678, P3_INSTQUEUE_REG_8__5__SCAN_IN, P3_U2582);
  nand ginst29854 (P3_U7679, P3_INSTQUEUE_REG_9__5__SCAN_IN, P3_U2581);
  nand ginst29855 (P3_U7680, P3_INSTQUEUE_REG_10__5__SCAN_IN, P3_U2580);
  nand ginst29856 (P3_U7681, P3_INSTQUEUE_REG_11__5__SCAN_IN, P3_U2579);
  nand ginst29857 (P3_U7682, P3_INSTQUEUE_REG_12__5__SCAN_IN, P3_U2577);
  nand ginst29858 (P3_U7683, P3_INSTQUEUE_REG_13__5__SCAN_IN, P3_U2576);
  nand ginst29859 (P3_U7684, P3_INSTQUEUE_REG_14__5__SCAN_IN, P3_U2575);
  nand ginst29860 (P3_U7685, P3_INSTQUEUE_REG_15__5__SCAN_IN, P3_U2574);
  nand ginst29861 (P3_U7686, P3_INSTQUEUE_REG_0__5__SCAN_IN, P3_U2572);
  nand ginst29862 (P3_U7687, P3_INSTQUEUE_REG_1__5__SCAN_IN, P3_U2571);
  nand ginst29863 (P3_U7688, P3_INSTQUEUE_REG_2__5__SCAN_IN, P3_U2570);
  nand ginst29864 (P3_U7689, P3_INSTQUEUE_REG_3__5__SCAN_IN, P3_U2569);
  nand ginst29865 (P3_U7690, P3_INSTQUEUE_REG_4__5__SCAN_IN, P3_U2567);
  nand ginst29866 (P3_U7691, P3_INSTQUEUE_REG_5__5__SCAN_IN, P3_U2566);
  nand ginst29867 (P3_U7692, P3_INSTQUEUE_REG_6__5__SCAN_IN, P3_U2565);
  nand ginst29868 (P3_U7693, P3_INSTQUEUE_REG_7__5__SCAN_IN, P3_U2564);
  nand ginst29869 (P3_U7694, P3_INSTQUEUE_REG_8__4__SCAN_IN, P3_U2582);
  nand ginst29870 (P3_U7695, P3_INSTQUEUE_REG_9__4__SCAN_IN, P3_U2581);
  nand ginst29871 (P3_U7696, P3_INSTQUEUE_REG_10__4__SCAN_IN, P3_U2580);
  nand ginst29872 (P3_U7697, P3_INSTQUEUE_REG_11__4__SCAN_IN, P3_U2579);
  nand ginst29873 (P3_U7698, P3_INSTQUEUE_REG_12__4__SCAN_IN, P3_U2577);
  nand ginst29874 (P3_U7699, P3_INSTQUEUE_REG_13__4__SCAN_IN, P3_U2576);
  nand ginst29875 (P3_U7700, P3_INSTQUEUE_REG_14__4__SCAN_IN, P3_U2575);
  nand ginst29876 (P3_U7701, P3_INSTQUEUE_REG_15__4__SCAN_IN, P3_U2574);
  nand ginst29877 (P3_U7702, P3_INSTQUEUE_REG_0__4__SCAN_IN, P3_U2572);
  nand ginst29878 (P3_U7703, P3_INSTQUEUE_REG_1__4__SCAN_IN, P3_U2571);
  nand ginst29879 (P3_U7704, P3_INSTQUEUE_REG_2__4__SCAN_IN, P3_U2570);
  nand ginst29880 (P3_U7705, P3_INSTQUEUE_REG_3__4__SCAN_IN, P3_U2569);
  nand ginst29881 (P3_U7706, P3_INSTQUEUE_REG_4__4__SCAN_IN, P3_U2567);
  nand ginst29882 (P3_U7707, P3_INSTQUEUE_REG_5__4__SCAN_IN, P3_U2566);
  nand ginst29883 (P3_U7708, P3_INSTQUEUE_REG_6__4__SCAN_IN, P3_U2565);
  nand ginst29884 (P3_U7709, P3_INSTQUEUE_REG_7__4__SCAN_IN, P3_U2564);
  nand ginst29885 (P3_U7710, P3_INSTQUEUE_REG_8__3__SCAN_IN, P3_U2582);
  nand ginst29886 (P3_U7711, P3_INSTQUEUE_REG_9__3__SCAN_IN, P3_U2581);
  nand ginst29887 (P3_U7712, P3_INSTQUEUE_REG_10__3__SCAN_IN, P3_U2580);
  nand ginst29888 (P3_U7713, P3_INSTQUEUE_REG_11__3__SCAN_IN, P3_U2579);
  nand ginst29889 (P3_U7714, P3_INSTQUEUE_REG_12__3__SCAN_IN, P3_U2577);
  nand ginst29890 (P3_U7715, P3_INSTQUEUE_REG_13__3__SCAN_IN, P3_U2576);
  nand ginst29891 (P3_U7716, P3_INSTQUEUE_REG_14__3__SCAN_IN, P3_U2575);
  nand ginst29892 (P3_U7717, P3_INSTQUEUE_REG_15__3__SCAN_IN, P3_U2574);
  nand ginst29893 (P3_U7718, P3_INSTQUEUE_REG_0__3__SCAN_IN, P3_U2572);
  nand ginst29894 (P3_U7719, P3_INSTQUEUE_REG_1__3__SCAN_IN, P3_U2571);
  nand ginst29895 (P3_U7720, P3_INSTQUEUE_REG_2__3__SCAN_IN, P3_U2570);
  nand ginst29896 (P3_U7721, P3_INSTQUEUE_REG_3__3__SCAN_IN, P3_U2569);
  nand ginst29897 (P3_U7722, P3_INSTQUEUE_REG_4__3__SCAN_IN, P3_U2567);
  nand ginst29898 (P3_U7723, P3_INSTQUEUE_REG_5__3__SCAN_IN, P3_U2566);
  nand ginst29899 (P3_U7724, P3_INSTQUEUE_REG_6__3__SCAN_IN, P3_U2565);
  nand ginst29900 (P3_U7725, P3_INSTQUEUE_REG_7__3__SCAN_IN, P3_U2564);
  nand ginst29901 (P3_U7726, P3_INSTQUEUE_REG_8__2__SCAN_IN, P3_U2582);
  nand ginst29902 (P3_U7727, P3_INSTQUEUE_REG_9__2__SCAN_IN, P3_U2581);
  nand ginst29903 (P3_U7728, P3_INSTQUEUE_REG_10__2__SCAN_IN, P3_U2580);
  nand ginst29904 (P3_U7729, P3_INSTQUEUE_REG_11__2__SCAN_IN, P3_U2579);
  nand ginst29905 (P3_U7730, P3_INSTQUEUE_REG_12__2__SCAN_IN, P3_U2577);
  nand ginst29906 (P3_U7731, P3_INSTQUEUE_REG_13__2__SCAN_IN, P3_U2576);
  nand ginst29907 (P3_U7732, P3_INSTQUEUE_REG_14__2__SCAN_IN, P3_U2575);
  nand ginst29908 (P3_U7733, P3_INSTQUEUE_REG_15__2__SCAN_IN, P3_U2574);
  nand ginst29909 (P3_U7734, P3_INSTQUEUE_REG_0__2__SCAN_IN, P3_U2572);
  nand ginst29910 (P3_U7735, P3_INSTQUEUE_REG_1__2__SCAN_IN, P3_U2571);
  nand ginst29911 (P3_U7736, P3_INSTQUEUE_REG_2__2__SCAN_IN, P3_U2570);
  nand ginst29912 (P3_U7737, P3_INSTQUEUE_REG_3__2__SCAN_IN, P3_U2569);
  nand ginst29913 (P3_U7738, P3_INSTQUEUE_REG_4__2__SCAN_IN, P3_U2567);
  nand ginst29914 (P3_U7739, P3_INSTQUEUE_REG_5__2__SCAN_IN, P3_U2566);
  nand ginst29915 (P3_U7740, P3_INSTQUEUE_REG_6__2__SCAN_IN, P3_U2565);
  nand ginst29916 (P3_U7741, P3_INSTQUEUE_REG_7__2__SCAN_IN, P3_U2564);
  nand ginst29917 (P3_U7742, P3_INSTQUEUE_REG_8__1__SCAN_IN, P3_U2582);
  nand ginst29918 (P3_U7743, P3_INSTQUEUE_REG_9__1__SCAN_IN, P3_U2581);
  nand ginst29919 (P3_U7744, P3_INSTQUEUE_REG_10__1__SCAN_IN, P3_U2580);
  nand ginst29920 (P3_U7745, P3_INSTQUEUE_REG_11__1__SCAN_IN, P3_U2579);
  nand ginst29921 (P3_U7746, P3_INSTQUEUE_REG_12__1__SCAN_IN, P3_U2577);
  nand ginst29922 (P3_U7747, P3_INSTQUEUE_REG_13__1__SCAN_IN, P3_U2576);
  nand ginst29923 (P3_U7748, P3_INSTQUEUE_REG_14__1__SCAN_IN, P3_U2575);
  nand ginst29924 (P3_U7749, P3_INSTQUEUE_REG_15__1__SCAN_IN, P3_U2574);
  nand ginst29925 (P3_U7750, P3_INSTQUEUE_REG_0__1__SCAN_IN, P3_U2572);
  nand ginst29926 (P3_U7751, P3_INSTQUEUE_REG_1__1__SCAN_IN, P3_U2571);
  nand ginst29927 (P3_U7752, P3_INSTQUEUE_REG_2__1__SCAN_IN, P3_U2570);
  nand ginst29928 (P3_U7753, P3_INSTQUEUE_REG_3__1__SCAN_IN, P3_U2569);
  nand ginst29929 (P3_U7754, P3_INSTQUEUE_REG_4__1__SCAN_IN, P3_U2567);
  nand ginst29930 (P3_U7755, P3_INSTQUEUE_REG_5__1__SCAN_IN, P3_U2566);
  nand ginst29931 (P3_U7756, P3_INSTQUEUE_REG_6__1__SCAN_IN, P3_U2565);
  nand ginst29932 (P3_U7757, P3_INSTQUEUE_REG_7__1__SCAN_IN, P3_U2564);
  nand ginst29933 (P3_U7758, P3_INSTQUEUE_REG_8__0__SCAN_IN, P3_U2582);
  nand ginst29934 (P3_U7759, P3_INSTQUEUE_REG_9__0__SCAN_IN, P3_U2581);
  nand ginst29935 (P3_U7760, P3_INSTQUEUE_REG_10__0__SCAN_IN, P3_U2580);
  nand ginst29936 (P3_U7761, P3_INSTQUEUE_REG_11__0__SCAN_IN, P3_U2579);
  nand ginst29937 (P3_U7762, P3_INSTQUEUE_REG_12__0__SCAN_IN, P3_U2577);
  nand ginst29938 (P3_U7763, P3_INSTQUEUE_REG_13__0__SCAN_IN, P3_U2576);
  nand ginst29939 (P3_U7764, P3_INSTQUEUE_REG_14__0__SCAN_IN, P3_U2575);
  nand ginst29940 (P3_U7765, P3_INSTQUEUE_REG_15__0__SCAN_IN, P3_U2574);
  nand ginst29941 (P3_U7766, P3_INSTQUEUE_REG_0__0__SCAN_IN, P3_U2572);
  nand ginst29942 (P3_U7767, P3_INSTQUEUE_REG_1__0__SCAN_IN, P3_U2571);
  nand ginst29943 (P3_U7768, P3_INSTQUEUE_REG_2__0__SCAN_IN, P3_U2570);
  nand ginst29944 (P3_U7769, P3_INSTQUEUE_REG_3__0__SCAN_IN, P3_U2569);
  nand ginst29945 (P3_U7770, P3_INSTQUEUE_REG_4__0__SCAN_IN, P3_U2567);
  nand ginst29946 (P3_U7771, P3_INSTQUEUE_REG_5__0__SCAN_IN, P3_U2566);
  nand ginst29947 (P3_U7772, P3_INSTQUEUE_REG_6__0__SCAN_IN, P3_U2565);
  nand ginst29948 (P3_U7773, P3_INSTQUEUE_REG_7__0__SCAN_IN, P3_U2564);
  nand ginst29949 (P3_U7774, P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P3_U3097);
  not ginst29950 (P3_U7775, P3_U3268);
  nand ginst29951 (P3_U7776, P3_INSTQUEUE_REG_8__7__SCAN_IN, P3_U2600);
  nand ginst29952 (P3_U7777, P3_INSTQUEUE_REG_9__7__SCAN_IN, P3_U2599);
  nand ginst29953 (P3_U7778, P3_INSTQUEUE_REG_10__7__SCAN_IN, P3_U2598);
  nand ginst29954 (P3_U7779, P3_INSTQUEUE_REG_11__7__SCAN_IN, P3_U2597);
  nand ginst29955 (P3_U7780, P3_INSTQUEUE_REG_12__7__SCAN_IN, P3_U2595);
  nand ginst29956 (P3_U7781, P3_INSTQUEUE_REG_13__7__SCAN_IN, P3_U2594);
  nand ginst29957 (P3_U7782, P3_INSTQUEUE_REG_14__7__SCAN_IN, P3_U2593);
  nand ginst29958 (P3_U7783, P3_INSTQUEUE_REG_15__7__SCAN_IN, P3_U2592);
  nand ginst29959 (P3_U7784, P3_INSTQUEUE_REG_0__7__SCAN_IN, P3_U2591);
  nand ginst29960 (P3_U7785, P3_INSTQUEUE_REG_1__7__SCAN_IN, P3_U2590);
  nand ginst29961 (P3_U7786, P3_INSTQUEUE_REG_2__7__SCAN_IN, P3_U2589);
  nand ginst29962 (P3_U7787, P3_INSTQUEUE_REG_3__7__SCAN_IN, P3_U2588);
  nand ginst29963 (P3_U7788, P3_INSTQUEUE_REG_4__7__SCAN_IN, P3_U2586);
  nand ginst29964 (P3_U7789, P3_INSTQUEUE_REG_5__7__SCAN_IN, P3_U2585);
  nand ginst29965 (P3_U7790, P3_INSTQUEUE_REG_6__7__SCAN_IN, P3_U2584);
  nand ginst29966 (P3_U7791, P3_INSTQUEUE_REG_7__7__SCAN_IN, P3_U2583);
  nand ginst29967 (P3_U7792, P3_INSTQUEUE_REG_8__6__SCAN_IN, P3_U2600);
  nand ginst29968 (P3_U7793, P3_INSTQUEUE_REG_9__6__SCAN_IN, P3_U2599);
  nand ginst29969 (P3_U7794, P3_INSTQUEUE_REG_10__6__SCAN_IN, P3_U2598);
  nand ginst29970 (P3_U7795, P3_INSTQUEUE_REG_11__6__SCAN_IN, P3_U2597);
  nand ginst29971 (P3_U7796, P3_INSTQUEUE_REG_12__6__SCAN_IN, P3_U2595);
  nand ginst29972 (P3_U7797, P3_INSTQUEUE_REG_13__6__SCAN_IN, P3_U2594);
  nand ginst29973 (P3_U7798, P3_INSTQUEUE_REG_14__6__SCAN_IN, P3_U2593);
  nand ginst29974 (P3_U7799, P3_INSTQUEUE_REG_15__6__SCAN_IN, P3_U2592);
  nand ginst29975 (P3_U7800, P3_INSTQUEUE_REG_0__6__SCAN_IN, P3_U2591);
  nand ginst29976 (P3_U7801, P3_INSTQUEUE_REG_1__6__SCAN_IN, P3_U2590);
  nand ginst29977 (P3_U7802, P3_INSTQUEUE_REG_2__6__SCAN_IN, P3_U2589);
  nand ginst29978 (P3_U7803, P3_INSTQUEUE_REG_3__6__SCAN_IN, P3_U2588);
  nand ginst29979 (P3_U7804, P3_INSTQUEUE_REG_4__6__SCAN_IN, P3_U2586);
  nand ginst29980 (P3_U7805, P3_INSTQUEUE_REG_5__6__SCAN_IN, P3_U2585);
  nand ginst29981 (P3_U7806, P3_INSTQUEUE_REG_6__6__SCAN_IN, P3_U2584);
  nand ginst29982 (P3_U7807, P3_INSTQUEUE_REG_7__6__SCAN_IN, P3_U2583);
  nand ginst29983 (P3_U7808, P3_INSTQUEUE_REG_8__5__SCAN_IN, P3_U2600);
  nand ginst29984 (P3_U7809, P3_INSTQUEUE_REG_9__5__SCAN_IN, P3_U2599);
  nand ginst29985 (P3_U7810, P3_INSTQUEUE_REG_10__5__SCAN_IN, P3_U2598);
  nand ginst29986 (P3_U7811, P3_INSTQUEUE_REG_11__5__SCAN_IN, P3_U2597);
  nand ginst29987 (P3_U7812, P3_INSTQUEUE_REG_12__5__SCAN_IN, P3_U2595);
  nand ginst29988 (P3_U7813, P3_INSTQUEUE_REG_13__5__SCAN_IN, P3_U2594);
  nand ginst29989 (P3_U7814, P3_INSTQUEUE_REG_14__5__SCAN_IN, P3_U2593);
  nand ginst29990 (P3_U7815, P3_INSTQUEUE_REG_15__5__SCAN_IN, P3_U2592);
  nand ginst29991 (P3_U7816, P3_INSTQUEUE_REG_0__5__SCAN_IN, P3_U2591);
  nand ginst29992 (P3_U7817, P3_INSTQUEUE_REG_1__5__SCAN_IN, P3_U2590);
  nand ginst29993 (P3_U7818, P3_INSTQUEUE_REG_2__5__SCAN_IN, P3_U2589);
  nand ginst29994 (P3_U7819, P3_INSTQUEUE_REG_3__5__SCAN_IN, P3_U2588);
  nand ginst29995 (P3_U7820, P3_INSTQUEUE_REG_4__5__SCAN_IN, P3_U2586);
  nand ginst29996 (P3_U7821, P3_INSTQUEUE_REG_5__5__SCAN_IN, P3_U2585);
  nand ginst29997 (P3_U7822, P3_INSTQUEUE_REG_6__5__SCAN_IN, P3_U2584);
  nand ginst29998 (P3_U7823, P3_INSTQUEUE_REG_7__5__SCAN_IN, P3_U2583);
  nand ginst29999 (P3_U7824, P3_INSTQUEUE_REG_8__4__SCAN_IN, P3_U2600);
  nand ginst30000 (P3_U7825, P3_INSTQUEUE_REG_9__4__SCAN_IN, P3_U2599);
  nand ginst30001 (P3_U7826, P3_INSTQUEUE_REG_10__4__SCAN_IN, P3_U2598);
  nand ginst30002 (P3_U7827, P3_INSTQUEUE_REG_11__4__SCAN_IN, P3_U2597);
  nand ginst30003 (P3_U7828, P3_INSTQUEUE_REG_12__4__SCAN_IN, P3_U2595);
  nand ginst30004 (P3_U7829, P3_INSTQUEUE_REG_13__4__SCAN_IN, P3_U2594);
  nand ginst30005 (P3_U7830, P3_INSTQUEUE_REG_14__4__SCAN_IN, P3_U2593);
  nand ginst30006 (P3_U7831, P3_INSTQUEUE_REG_15__4__SCAN_IN, P3_U2592);
  nand ginst30007 (P3_U7832, P3_INSTQUEUE_REG_0__4__SCAN_IN, P3_U2591);
  nand ginst30008 (P3_U7833, P3_INSTQUEUE_REG_1__4__SCAN_IN, P3_U2590);
  nand ginst30009 (P3_U7834, P3_INSTQUEUE_REG_2__4__SCAN_IN, P3_U2589);
  nand ginst30010 (P3_U7835, P3_INSTQUEUE_REG_3__4__SCAN_IN, P3_U2588);
  nand ginst30011 (P3_U7836, P3_INSTQUEUE_REG_4__4__SCAN_IN, P3_U2586);
  nand ginst30012 (P3_U7837, P3_INSTQUEUE_REG_5__4__SCAN_IN, P3_U2585);
  nand ginst30013 (P3_U7838, P3_INSTQUEUE_REG_6__4__SCAN_IN, P3_U2584);
  nand ginst30014 (P3_U7839, P3_INSTQUEUE_REG_7__4__SCAN_IN, P3_U2583);
  nand ginst30015 (P3_U7840, P3_INSTQUEUE_REG_8__3__SCAN_IN, P3_U2600);
  nand ginst30016 (P3_U7841, P3_INSTQUEUE_REG_9__3__SCAN_IN, P3_U2599);
  nand ginst30017 (P3_U7842, P3_INSTQUEUE_REG_10__3__SCAN_IN, P3_U2598);
  nand ginst30018 (P3_U7843, P3_INSTQUEUE_REG_11__3__SCAN_IN, P3_U2597);
  nand ginst30019 (P3_U7844, P3_INSTQUEUE_REG_12__3__SCAN_IN, P3_U2595);
  nand ginst30020 (P3_U7845, P3_INSTQUEUE_REG_13__3__SCAN_IN, P3_U2594);
  nand ginst30021 (P3_U7846, P3_INSTQUEUE_REG_14__3__SCAN_IN, P3_U2593);
  nand ginst30022 (P3_U7847, P3_INSTQUEUE_REG_15__3__SCAN_IN, P3_U2592);
  nand ginst30023 (P3_U7848, P3_INSTQUEUE_REG_0__3__SCAN_IN, P3_U2591);
  nand ginst30024 (P3_U7849, P3_INSTQUEUE_REG_1__3__SCAN_IN, P3_U2590);
  nand ginst30025 (P3_U7850, P3_INSTQUEUE_REG_2__3__SCAN_IN, P3_U2589);
  nand ginst30026 (P3_U7851, P3_INSTQUEUE_REG_3__3__SCAN_IN, P3_U2588);
  nand ginst30027 (P3_U7852, P3_INSTQUEUE_REG_4__3__SCAN_IN, P3_U2586);
  nand ginst30028 (P3_U7853, P3_INSTQUEUE_REG_5__3__SCAN_IN, P3_U2585);
  nand ginst30029 (P3_U7854, P3_INSTQUEUE_REG_6__3__SCAN_IN, P3_U2584);
  nand ginst30030 (P3_U7855, P3_INSTQUEUE_REG_7__3__SCAN_IN, P3_U2583);
  nand ginst30031 (P3_U7856, P3_INSTQUEUE_REG_8__2__SCAN_IN, P3_U2600);
  nand ginst30032 (P3_U7857, P3_INSTQUEUE_REG_9__2__SCAN_IN, P3_U2599);
  nand ginst30033 (P3_U7858, P3_INSTQUEUE_REG_10__2__SCAN_IN, P3_U2598);
  nand ginst30034 (P3_U7859, P3_INSTQUEUE_REG_11__2__SCAN_IN, P3_U2597);
  nand ginst30035 (P3_U7860, P3_INSTQUEUE_REG_12__2__SCAN_IN, P3_U2595);
  nand ginst30036 (P3_U7861, P3_INSTQUEUE_REG_13__2__SCAN_IN, P3_U2594);
  nand ginst30037 (P3_U7862, P3_INSTQUEUE_REG_14__2__SCAN_IN, P3_U2593);
  nand ginst30038 (P3_U7863, P3_INSTQUEUE_REG_15__2__SCAN_IN, P3_U2592);
  nand ginst30039 (P3_U7864, P3_INSTQUEUE_REG_0__2__SCAN_IN, P3_U2591);
  nand ginst30040 (P3_U7865, P3_INSTQUEUE_REG_1__2__SCAN_IN, P3_U2590);
  nand ginst30041 (P3_U7866, P3_INSTQUEUE_REG_2__2__SCAN_IN, P3_U2589);
  nand ginst30042 (P3_U7867, P3_INSTQUEUE_REG_3__2__SCAN_IN, P3_U2588);
  nand ginst30043 (P3_U7868, P3_INSTQUEUE_REG_4__2__SCAN_IN, P3_U2586);
  nand ginst30044 (P3_U7869, P3_INSTQUEUE_REG_5__2__SCAN_IN, P3_U2585);
  nand ginst30045 (P3_U7870, P3_INSTQUEUE_REG_6__2__SCAN_IN, P3_U2584);
  nand ginst30046 (P3_U7871, P3_INSTQUEUE_REG_7__2__SCAN_IN, P3_U2583);
  nand ginst30047 (P3_U7872, P3_INSTQUEUE_REG_8__1__SCAN_IN, P3_U2600);
  nand ginst30048 (P3_U7873, P3_INSTQUEUE_REG_9__1__SCAN_IN, P3_U2599);
  nand ginst30049 (P3_U7874, P3_INSTQUEUE_REG_10__1__SCAN_IN, P3_U2598);
  nand ginst30050 (P3_U7875, P3_INSTQUEUE_REG_11__1__SCAN_IN, P3_U2597);
  nand ginst30051 (P3_U7876, P3_INSTQUEUE_REG_12__1__SCAN_IN, P3_U2595);
  nand ginst30052 (P3_U7877, P3_INSTQUEUE_REG_13__1__SCAN_IN, P3_U2594);
  nand ginst30053 (P3_U7878, P3_INSTQUEUE_REG_14__1__SCAN_IN, P3_U2593);
  nand ginst30054 (P3_U7879, P3_INSTQUEUE_REG_15__1__SCAN_IN, P3_U2592);
  nand ginst30055 (P3_U7880, P3_INSTQUEUE_REG_0__1__SCAN_IN, P3_U2591);
  nand ginst30056 (P3_U7881, P3_INSTQUEUE_REG_1__1__SCAN_IN, P3_U2590);
  nand ginst30057 (P3_U7882, P3_INSTQUEUE_REG_2__1__SCAN_IN, P3_U2589);
  nand ginst30058 (P3_U7883, P3_INSTQUEUE_REG_3__1__SCAN_IN, P3_U2588);
  nand ginst30059 (P3_U7884, P3_INSTQUEUE_REG_4__1__SCAN_IN, P3_U2586);
  nand ginst30060 (P3_U7885, P3_INSTQUEUE_REG_5__1__SCAN_IN, P3_U2585);
  nand ginst30061 (P3_U7886, P3_INSTQUEUE_REG_6__1__SCAN_IN, P3_U2584);
  nand ginst30062 (P3_U7887, P3_INSTQUEUE_REG_7__1__SCAN_IN, P3_U2583);
  nand ginst30063 (P3_U7888, P3_INSTQUEUE_REG_8__0__SCAN_IN, P3_U2600);
  nand ginst30064 (P3_U7889, P3_INSTQUEUE_REG_9__0__SCAN_IN, P3_U2599);
  nand ginst30065 (P3_U7890, P3_INSTQUEUE_REG_10__0__SCAN_IN, P3_U2598);
  nand ginst30066 (P3_U7891, P3_INSTQUEUE_REG_11__0__SCAN_IN, P3_U2597);
  nand ginst30067 (P3_U7892, P3_INSTQUEUE_REG_12__0__SCAN_IN, P3_U2595);
  nand ginst30068 (P3_U7893, P3_INSTQUEUE_REG_13__0__SCAN_IN, P3_U2594);
  nand ginst30069 (P3_U7894, P3_INSTQUEUE_REG_14__0__SCAN_IN, P3_U2593);
  nand ginst30070 (P3_U7895, P3_INSTQUEUE_REG_15__0__SCAN_IN, P3_U2592);
  nand ginst30071 (P3_U7896, P3_INSTQUEUE_REG_0__0__SCAN_IN, P3_U2591);
  nand ginst30072 (P3_U7897, P3_INSTQUEUE_REG_1__0__SCAN_IN, P3_U2590);
  nand ginst30073 (P3_U7898, P3_INSTQUEUE_REG_2__0__SCAN_IN, P3_U2589);
  nand ginst30074 (P3_U7899, P3_INSTQUEUE_REG_3__0__SCAN_IN, P3_U2588);
  nand ginst30075 (P3_U7900, P3_INSTQUEUE_REG_4__0__SCAN_IN, P3_U2586);
  nand ginst30076 (P3_U7901, P3_INSTQUEUE_REG_5__0__SCAN_IN, P3_U2585);
  nand ginst30077 (P3_U7902, P3_INSTQUEUE_REG_6__0__SCAN_IN, P3_U2584);
  nand ginst30078 (P3_U7903, P3_INSTQUEUE_REG_7__0__SCAN_IN, P3_U2583);
  nand ginst30079 (P3_U7904, P3_STATE_REG_0__SCAN_IN, P3_U4292);
  or ginst30080 (P3_U7905, P3_STATE2_REG_2__SCAN_IN, U209);
  nand ginst30081 (P3_U7906, P3_U3939, P3_U6397);
  nand ginst30082 (P3_U7907, P3_U2603, P3_U4134);
  nand ginst30083 (P3_U7908, P3_U2404, P3_U3256);
  nand ginst30084 (P3_U7909, P3_U2392, P3_U7096);
  nand ginst30085 (P3_U7910, P3_U4317, P3_U7908, P3_U7909);
  not ginst30086 (P3_U7911, P3_U3086);
  nand ginst30087 (P3_U7912, P3_U3088, P3_U7911);
  nand ginst30088 (P3_U7913, P3_STATE_REG_1__SCAN_IN, P3_U4446, P3_U4449);
  nand ginst30089 (P3_U7914, P3_STATE_REG_2__SCAN_IN, P3_U7904);
  nand ginst30090 (P3_U7915, P3_STATE_REG_1__SCAN_IN, P3_U4446);
  nand ginst30091 (P3_U7916, P3_U3106, P3_U4505);
  nand ginst30092 (P3_U7917, P3_U4488, P3_U4522);
  nand ginst30093 (P3_U7918, P3_U3208, P3_U3219);
  nand ginst30094 (P3_U7919, P3_U3105, P3_U7376);
  nand ginst30095 (P3_U7920, P3_BE_N_REG_3__SCAN_IN, P3_U3077);
  nand ginst30096 (P3_U7921, P3_BYTEENABLE_REG_3__SCAN_IN, P3_U4308);
  nand ginst30097 (P3_U7922, P3_BE_N_REG_2__SCAN_IN, P3_U3077);
  nand ginst30098 (P3_U7923, P3_BYTEENABLE_REG_2__SCAN_IN, P3_U4308);
  nand ginst30099 (P3_U7924, P3_BE_N_REG_1__SCAN_IN, P3_U3077);
  nand ginst30100 (P3_U7925, P3_BYTEENABLE_REG_1__SCAN_IN, P3_U4308);
  nand ginst30101 (P3_U7926, P3_BE_N_REG_0__SCAN_IN, P3_U3077);
  nand ginst30102 (P3_U7927, P3_BYTEENABLE_REG_0__SCAN_IN, P3_U4308);
  nand ginst30103 (P3_U7928, P3_STATE_REG_0__SCAN_IN, P3_REQUESTPENDING_REG_SCAN_IN, P3_U3079);
  nand ginst30104 (P3_U7929, P3_STATE_REG_2__SCAN_IN, P3_U3086);
  nand ginst30105 (P3_U7930, P3_U7928, P3_U7929);
  nand ginst30106 (P3_U7931, P3_STATE_REG_1__SCAN_IN, P3_U4449, P3_U7914);
  nand ginst30107 (P3_U7932, P3_U3076, P3_U7930);
  nand ginst30108 (P3_U7933, P3_STATE_REG_2__SCAN_IN, P3_STATE_REG_0__SCAN_IN, P3_U3087);
  nand ginst30109 (P3_U7934, P3_U3079, P3_U4459);
  or ginst30110 (P3_U7935, P3_STATE_REG_1__SCAN_IN, P3_STATE_REG_0__SCAN_IN);
  nand ginst30111 (P3_U7936, P3_STATE_REG_0__SCAN_IN, P3_U4346);
  not ginst30112 (P3_U7937, P3_U3278);
  nand ginst30113 (P3_U7938, P3_DATAWIDTH_REG_0__SCAN_IN, P3_U7937);
  nand ginst30114 (P3_U7939, P3_U3278, P3_U3279);
  nand ginst30115 (P3_U7940, P3_U3278, P3_U4464);
  nand ginst30116 (P3_U7941, P3_DATAWIDTH_REG_1__SCAN_IN, P3_U7937);
  nand ginst30117 (P3_U7942, P3_U3211, P3_U4505);
  nand ginst30118 (P3_U7943, P3_U3104, P3_U3214);
  nand ginst30119 (P3_U7944, P3_U3213, P3_U4505);
  nand ginst30120 (P3_U7945, P3_U3104, P3_U3210);
  nand ginst30121 (P3_U7946, P3_U4539, P3_U4618);
  nand ginst30122 (P3_U7947, P3_U3101, P3_U4620);
  nand ginst30123 (P3_U7948, P3_U4281, P3_U4617);
  nand ginst30124 (P3_U7949, P3_U4622, P3_U4624);
  nand ginst30125 (P3_U7950, P3_U3237, P3_U4505);
  nand ginst30126 (P3_U7951, P3_U3104, P3_U3238);
  nand ginst30127 (P3_U7952, P3_STATE2_REG_0__SCAN_IN, P3_U4627);
  nand ginst30128 (P3_U7953, P3_U3121, P3_U4628);
  nand ginst30129 (P3_U7954, P3_STATE2_REG_3__SCAN_IN, P3_U3122);
  nand ginst30130 (P3_U7955, P3_U2453, P3_U4630);
  or ginst30131 (P3_U7956, P3_STATE2_REG_0__SCAN_IN, P3_STATEBS16_REG_SCAN_IN);
  nand ginst30132 (P3_U7957, P3_STATE2_REG_0__SCAN_IN, P3_U7905);
  nand ginst30133 (P3_U7958, P3_STATE2_REG_0__SCAN_IN, P3_U4638);
  nand ginst30134 (P3_U7959, P3_U3121, P3_U4629, P3_U4637);
  nand ginst30135 (P3_U7960, P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN, P3_U3130);
  nand ginst30136 (P3_U7961, P3_U3131, P3_U4648);
  not ginst30137 (P3_U7962, P3_U3269);
  nand ginst30138 (P3_U7963, P3_U4653, P3_U7962);
  nand ginst30139 (P3_U7964, P3_U3138, P3_U3269);
  not ginst30140 (P3_U7965, P3_U3270);
  nand ginst30141 (P3_U7966, P3_U4657, P3_U7965);
  nand ginst30142 (P3_U7967, P3_U3140, P3_U3270);
  not ginst30143 (P3_U7968, P3_U3271);
  nand ginst30144 (P3_U7969, P3_U3101, P3_U3109);
  nand ginst30145 (P3_U7970, P3_U4539, P3_U5483);
  nand ginst30146 (P3_U7971, P3_U3283, P3_U4283);
  nand ginst30147 (P3_U7972, P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN, P3_U5499);
  nand ginst30148 (P3_U7973, P3_U3107, P3_U3218);
  nand ginst30149 (P3_U7974, P3_U4573, P3_U4590);
  nand ginst30150 (P3_U7975, P3_U4539, P3_U5512);
  nand ginst30151 (P3_U7976, P3_U3101, P3_U5515);
  nand ginst30152 (P3_U7977, P3_U3110, P3_U4556, P3_U5517);
  nand ginst30153 (P3_U7978, P3_U3107, P3_U4590, P3_U5513);
  nand ginst30154 (P3_U7979, P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P3_U5499);
  nand ginst30155 (P3_U7980, P3_U4283, P3_U5546);
  nand ginst30156 (P3_U7981, P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN, P3_U3094, P3_U3221);
  nand ginst30157 (P3_U7982, P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P3_U3097, P3_U5531);
  nand ginst30158 (P3_U7983, P3_INSTADDRPOINTER_REG_1__SCAN_IN, P3_U4284);
  nand ginst30159 (P3_U7984, P3_INSTADDRPOINTER_REG_31__SCAN_IN, P3_SUB_580_U6);
  not ginst30160 (P3_U7985, P3_U3287);
  nand ginst30161 (P3_U7986, P3_INSTADDRPOINTER_REG_0__SCAN_IN, P3_U4284);
  nand ginst30162 (P3_U7987, P3_INSTADDRPOINTER_REG_0__SCAN_IN, P3_INSTADDRPOINTER_REG_31__SCAN_IN);
  not ginst30163 (P3_U7988, P3_U3286);
  nand ginst30164 (P3_U7989, P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN, P3_U5499);
  nand ginst30165 (P3_U7990, P3_U4283, P3_U5557);
  nand ginst30166 (P3_U7991, P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P3_U5499);
  nand ginst30167 (P3_U7992, P3_U4283, P3_U5570);
  nand ginst30168 (P3_U7993, P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN, P3_U3221);
  nand ginst30169 (P3_U7994, P3_U3093, P3_U5571);
  nand ginst30170 (P3_U7995, P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN, P3_U5499);
  nand ginst30171 (P3_U7996, P3_U4283, P3_U5577);
  nand ginst30172 (P3_U7997, P3_U4647, P3_U7968);
  nand ginst30173 (P3_U7998, P3_U3143, P3_U3271);
  nand ginst30174 (P3_U7999, P3_U7997, P3_U7998);
  nand ginst30175 (P3_U8000, P3_U3104, P3_U5622);
  nand ginst30176 (P3_U8001, P3_U4505, P3_U5619);
  nand ginst30177 (P3_U8002, P3_BYTEENABLE_REG_3__SCAN_IN, P3_U3261);
  nand ginst30178 (P3_U8003, P3_U3291, P3_U4307);
  or ginst30179 (P3_U8004, P3_DATAWIDTH_REG_0__SCAN_IN, P3_DATAWIDTH_REG_1__SCAN_IN);
  nand ginst30180 (P3_U8005, P3_DATAWIDTH_REG_0__SCAN_IN, P3_U3240);
  nand ginst30181 (P3_U8006, P3_U8004, P3_U8005);
  nand ginst30182 (P3_U8007, P3_U3081, P3_U8006);
  nand ginst30183 (P3_U8008, P3_REIP_REG_0__SCAN_IN, P3_REIP_REG_1__SCAN_IN);
  nand ginst30184 (P3_U8009, P3_U8007, P3_U8008);
  nand ginst30185 (P3_U8010, P3_BYTEENABLE_REG_2__SCAN_IN, P3_U3261);
  nand ginst30186 (P3_U8011, P3_U4307, P3_U8009);
  nand ginst30187 (P3_U8012, P3_BYTEENABLE_REG_1__SCAN_IN, P3_U3261);
  nand ginst30188 (P3_U8013, P3_REIP_REG_1__SCAN_IN, P3_U4307);
  nand ginst30189 (P3_U8014, P3_BYTEENABLE_REG_0__SCAN_IN, P3_U3261);
  nand ginst30190 (P3_U8015, P3_U4307, P3_U7367);
  nand ginst30191 (P3_U8016, P3_U3264, P3_U4308);
  nand ginst30192 (P3_U8017, P3_W_R_N_REG_SCAN_IN, P3_U3077);
  nand ginst30193 (P3_U8018, P3_U4617, P3_U7368);
  nand ginst30194 (P3_U8019, P3_MORE_REG_SCAN_IN, P3_U4285);
  nand ginst30195 (P3_U8020, P3_STATEBS16_REG_SCAN_IN, P3_U7937);
  nand ginst30196 (P3_U8021, BS16, P3_U3278);
  nand ginst30197 (P3_U8022, P3_REQUESTPENDING_REG_SCAN_IN, P3_U7374);
  nand ginst30198 (P3_U8023, P3_U4287, P3_U7379);
  nand ginst30199 (P3_U8024, P3_U3263, P3_U4308);
  nand ginst30200 (P3_U8025, P3_D_C_N_REG_SCAN_IN, P3_U3077);
  nand ginst30201 (P3_U8026, P3_M_IO_N_REG_SCAN_IN, P3_U3077);
  nand ginst30202 (P3_U8027, P3_MEMORYFETCH_REG_SCAN_IN, P3_U4308);
  nand ginst30203 (P3_U8028, P3_READREQUEST_REG_SCAN_IN, P3_U7384);
  nand ginst30204 (P3_U8029, P3_U4288, P3_U7385);
  nand ginst30205 (P3_U8030, P3_MEMORYFETCH_REG_SCAN_IN, P3_U7384);
  nand ginst30206 (P3_U8031, P3_U4288, P3_U7386);
  nand ginst30207 (P3_U8032, P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P3_U3097);
  nand ginst30208 (P3_U8033, P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN, P3_U3094);
  not ginst30209 (P3_U8034, P3_U3272);
  nand ginst30210 (P3_U8035, P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P3_U4289);
  nand ginst30211 (P3_U8036, P3_U3100, P3_U7645);
  not ginst30212 (P3_U8037, P3_U3273);
  nand ginst30213 (P3_U8038, P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN, P3_U3207);
  nand ginst30214 (P3_U8039, P3_FLUSH_REG_SCAN_IN, P3_U3286, P3_U3287);
  nand ginst30215 (P3_U8040, P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P3_U3207);
  nand ginst30216 (P3_U8041, P3_FLUSH_REG_SCAN_IN, P3_U3286, P3_U7985);
  nand ginst30217 (P3_U8042, P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN, P3_U3207);
  nand ginst30218 (P3_U8043, P3_FLUSH_REG_SCAN_IN, P3_U7988);
  nand ginst30219 (P3_U8044, P3_U3303, P3_U4290);
  nand ginst30220 (P3_U8045, P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN, P3_U5496);
  nand ginst30221 (P3_U8046, P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P3_U5496);
  nand ginst30222 (P3_U8047, P3_U4290, P3_U5542);
  nand ginst30223 (P3_U8048, P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN, P3_U5496);
  nand ginst30224 (P3_U8049, P3_U4290, P3_U5553);
  nand ginst30225 (P3_U8050, P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P3_U5496);
  nand ginst30226 (P3_U8051, P3_U4290, P3_U5566);
  nand ginst30227 (P3_U8052, P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN, P3_U5496);
  nand ginst30228 (P3_U8053, P3_U4290, P3_U5573);
  nor ginst30229 (R165_U10, P1_ADDRESS_REG_23__SCAN_IN, P1_ADDRESS_REG_11__SCAN_IN, P1_ADDRESS_REG_1__SCAN_IN, R165_U9);
  or ginst30230 (R165_U11, P1_ADDRESS_REG_28__SCAN_IN, P1_ADDRESS_REG_26__SCAN_IN, P1_ADDRESS_REG_21__SCAN_IN, P1_ADDRESS_REG_6__SCAN_IN);
  nor ginst30231 (R165_U12, P1_ADDRESS_REG_14__SCAN_IN, P1_ADDRESS_REG_12__SCAN_IN, P1_ADDRESS_REG_4__SCAN_IN, R165_U11);
  or ginst30232 (R165_U13, P1_ADDRESS_REG_27__SCAN_IN, P1_ADDRESS_REG_20__SCAN_IN, P1_ADDRESS_REG_13__SCAN_IN, P1_ADDRESS_REG_3__SCAN_IN);
  nor ginst30233 (R165_U14, P1_ADDRESS_REG_15__SCAN_IN, P1_ADDRESS_REG_5__SCAN_IN, P1_ADDRESS_REG_2__SCAN_IN, R165_U13);
  nand ginst30234 (R165_U15, R165_U10, R165_U12, R165_U14, R165_U8);
  and ginst30235 (R165_U6, P1_ADDRESS_REG_29__SCAN_IN, R165_U15);
  or ginst30236 (R165_U7, P1_ADDRESS_REG_22__SCAN_IN, P1_ADDRESS_REG_17__SCAN_IN, P1_ADDRESS_REG_9__SCAN_IN, P1_ADDRESS_REG_7__SCAN_IN);
  nor ginst30237 (R165_U8, P1_ADDRESS_REG_25__SCAN_IN, P1_ADDRESS_REG_24__SCAN_IN, P1_ADDRESS_REG_19__SCAN_IN, P1_ADDRESS_REG_10__SCAN_IN, R165_U7);
  or ginst30238 (R165_U9, P1_ADDRESS_REG_18__SCAN_IN, P1_ADDRESS_REG_16__SCAN_IN, P1_ADDRESS_REG_8__SCAN_IN, P1_ADDRESS_REG_0__SCAN_IN);
  nor ginst30239 (R170_U10, P2_ADDRESS_REG_23__SCAN_IN, P2_ADDRESS_REG_11__SCAN_IN, P2_ADDRESS_REG_1__SCAN_IN, R170_U9);
  or ginst30240 (R170_U11, P2_ADDRESS_REG_28__SCAN_IN, P2_ADDRESS_REG_26__SCAN_IN, P2_ADDRESS_REG_21__SCAN_IN, P2_ADDRESS_REG_6__SCAN_IN);
  nor ginst30241 (R170_U12, P2_ADDRESS_REG_14__SCAN_IN, P2_ADDRESS_REG_12__SCAN_IN, P2_ADDRESS_REG_4__SCAN_IN, R170_U11);
  or ginst30242 (R170_U13, P2_ADDRESS_REG_27__SCAN_IN, P2_ADDRESS_REG_20__SCAN_IN, P2_ADDRESS_REG_13__SCAN_IN, P2_ADDRESS_REG_3__SCAN_IN);
  nor ginst30243 (R170_U14, P2_ADDRESS_REG_15__SCAN_IN, P2_ADDRESS_REG_5__SCAN_IN, P2_ADDRESS_REG_2__SCAN_IN, R170_U13);
  nand ginst30244 (R170_U15, R170_U10, R170_U12, R170_U14, R170_U8);
  and ginst30245 (R170_U6, P2_ADDRESS_REG_29__SCAN_IN, R170_U15);
  or ginst30246 (R170_U7, P2_ADDRESS_REG_22__SCAN_IN, P2_ADDRESS_REG_17__SCAN_IN, P2_ADDRESS_REG_9__SCAN_IN, P2_ADDRESS_REG_7__SCAN_IN);
  nor ginst30247 (R170_U8, P2_ADDRESS_REG_25__SCAN_IN, P2_ADDRESS_REG_24__SCAN_IN, P2_ADDRESS_REG_19__SCAN_IN, P2_ADDRESS_REG_10__SCAN_IN, R170_U7);
  or ginst30248 (R170_U9, P2_ADDRESS_REG_18__SCAN_IN, P2_ADDRESS_REG_16__SCAN_IN, P2_ADDRESS_REG_8__SCAN_IN, P2_ADDRESS_REG_0__SCAN_IN);
  and ginst30249 (U207, U214, U250);
  and ginst30250 (U208, P2_W_R_N_REG_SCAN_IN, P2_M_IO_N_REG_SCAN_IN, U377, U378);
  and ginst30251 (U209, READY2, READY22_REG_SCAN_IN);
  and ginst30252 (U210, READY1, READY11_REG_SCAN_IN);
  and ginst30253 (U211, READY12_REG_SCAN_IN, READY21_REG_SCAN_IN);
  nand ginst30254 (U212, R170_U6, U208, U214);
  nand ginst30255 (U213, P3_M_IO_N_REG_SCAN_IN, U215, U379, U380);
  nand ginst30256 (U214, P1_M_IO_N_REG_SCAN_IN, P1_W_R_N_REG_SCAN_IN, R165_U6, U381, U383);
  nand ginst30257 (U215, LT_748_U6, U208);
  nand ginst30258 (U216, U482, U483, U484);
  nand ginst30259 (U217, U479, U480, U481);
  nand ginst30260 (U218, U476, U477, U478);
  nand ginst30261 (U219, U473, U474, U475);
  nand ginst30262 (U220, U470, U471, U472);
  nand ginst30263 (U221, U467, U468, U469);
  nand ginst30264 (U222, U464, U465, U466);
  nand ginst30265 (U223, U461, U462, U463);
  nand ginst30266 (U224, U458, U459, U460);
  nand ginst30267 (U225, U455, U456, U457);
  nand ginst30268 (U226, U452, U453, U454);
  nand ginst30269 (U227, U449, U450, U451);
  nand ginst30270 (U228, U446, U447, U448);
  nand ginst30271 (U229, U443, U444, U445);
  nand ginst30272 (U230, U440, U441, U442);
  nand ginst30273 (U231, U437, U438, U439);
  nand ginst30274 (U232, U434, U435, U436);
  nand ginst30275 (U233, U431, U432, U433);
  nand ginst30276 (U234, U428, U429, U430);
  nand ginst30277 (U235, U425, U426, U427);
  nand ginst30278 (U236, U422, U423, U424);
  nand ginst30279 (U237, U419, U420, U421);
  nand ginst30280 (U238, U416, U417, U418);
  nand ginst30281 (U239, U413, U414, U415);
  nand ginst30282 (U240, U410, U411, U412);
  nand ginst30283 (U241, U407, U408, U409);
  nand ginst30284 (U242, U404, U405, U406);
  nand ginst30285 (U243, U401, U402, U403);
  nand ginst30286 (U244, U398, U399, U400);
  nand ginst30287 (U245, U395, U396, U397);
  nand ginst30288 (U246, U392, U393, U394);
  nand ginst30289 (U247, U389, U390, U391);
  not ginst30290 (U248, R165_U6);
  not ginst30291 (U249, R170_U6);
  nand ginst30292 (U250, U214, U387);
  nand ginst30293 (U251, U485, U486);
  nand ginst30294 (U252, U487, U488);
  nand ginst30295 (U253, U489, U490);
  nand ginst30296 (U254, U491, U492);
  nand ginst30297 (U255, U493, U494);
  nand ginst30298 (U256, U495, U496);
  nand ginst30299 (U257, U497, U498);
  nand ginst30300 (U258, U499, U500);
  nand ginst30301 (U259, U501, U502);
  nand ginst30302 (U260, U503, U504);
  nand ginst30303 (U261, U505, U506);
  nand ginst30304 (U262, U507, U508);
  nand ginst30305 (U263, U509, U510);
  nand ginst30306 (U264, U511, U512);
  nand ginst30307 (U265, U513, U514);
  nand ginst30308 (U266, U515, U516);
  nand ginst30309 (U267, U517, U518);
  nand ginst30310 (U268, U519, U520);
  nand ginst30311 (U269, U521, U522);
  nand ginst30312 (U270, U523, U524);
  nand ginst30313 (U271, U525, U526);
  nand ginst30314 (U272, U527, U528);
  nand ginst30315 (U273, U529, U530);
  nand ginst30316 (U274, U531, U532);
  nand ginst30317 (U275, U533, U534);
  nand ginst30318 (U276, U535, U536);
  nand ginst30319 (U277, U537, U538);
  nand ginst30320 (U278, U539, U540);
  nand ginst30321 (U279, U541, U542);
  nand ginst30322 (U280, U543, U544);
  nand ginst30323 (U281, U545, U546);
  nand ginst30324 (U282, U547, U548);
  nand ginst30325 (U283, U549, U550);
  nand ginst30326 (U284, U551, U552);
  nand ginst30327 (U285, U553, U554);
  nand ginst30328 (U286, U555, U556);
  nand ginst30329 (U287, U557, U558);
  nand ginst30330 (U288, U559, U560);
  nand ginst30331 (U289, U561, U562);
  nand ginst30332 (U290, U563, U564);
  nand ginst30333 (U291, U565, U566);
  nand ginst30334 (U292, U567, U568);
  nand ginst30335 (U293, U569, U570);
  nand ginst30336 (U294, U571, U572);
  nand ginst30337 (U295, U573, U574);
  nand ginst30338 (U296, U575, U576);
  nand ginst30339 (U297, U577, U578);
  nand ginst30340 (U298, U579, U580);
  nand ginst30341 (U299, U581, U582);
  nand ginst30342 (U300, U583, U584);
  nand ginst30343 (U301, U585, U586);
  nand ginst30344 (U302, U587, U588);
  nand ginst30345 (U303, U589, U590);
  nand ginst30346 (U304, U591, U592);
  nand ginst30347 (U305, U593, U594);
  nand ginst30348 (U306, U595, U596);
  nand ginst30349 (U307, U597, U598);
  nand ginst30350 (U308, U599, U600);
  nand ginst30351 (U309, U601, U602);
  nand ginst30352 (U310, U603, U604);
  nand ginst30353 (U311, U605, U606);
  nand ginst30354 (U312, U607, U608);
  nand ginst30355 (U313, U609, U610);
  nand ginst30356 (U314, U611, U612);
  nand ginst30357 (U315, U613, U614);
  nand ginst30358 (U316, U615, U616);
  nand ginst30359 (U317, U617, U618);
  nand ginst30360 (U318, U619, U620);
  nand ginst30361 (U319, U621, U622);
  nand ginst30362 (U320, U623, U624);
  nand ginst30363 (U321, U625, U626);
  nand ginst30364 (U322, U627, U628);
  nand ginst30365 (U323, U629, U630);
  nand ginst30366 (U324, U631, U632);
  nand ginst30367 (U325, U633, U634);
  nand ginst30368 (U326, U635, U636);
  nand ginst30369 (U327, U637, U638);
  nand ginst30370 (U328, U639, U640);
  nand ginst30371 (U329, U641, U642);
  nand ginst30372 (U330, U643, U644);
  nand ginst30373 (U331, U645, U646);
  nand ginst30374 (U332, U647, U648);
  nand ginst30375 (U333, U649, U650);
  nand ginst30376 (U334, U651, U652);
  nand ginst30377 (U335, U653, U654);
  nand ginst30378 (U336, U655, U656);
  nand ginst30379 (U337, U657, U658);
  nand ginst30380 (U338, U659, U660);
  nand ginst30381 (U339, U661, U662);
  nand ginst30382 (U340, U663, U664);
  nand ginst30383 (U341, U665, U666);
  nand ginst30384 (U342, U667, U668);
  nand ginst30385 (U343, U669, U670);
  nand ginst30386 (U344, U671, U672);
  nand ginst30387 (U345, U673, U674);
  nand ginst30388 (U346, U675, U676);
  nand ginst30389 (U347, U677, U678);
  nand ginst30390 (U348, U679, U680);
  nand ginst30391 (U349, U681, U682);
  nand ginst30392 (U350, U683, U684);
  nand ginst30393 (U351, U685, U686);
  nand ginst30394 (U352, U687, U688);
  nand ginst30395 (U353, U689, U690);
  nand ginst30396 (U354, U691, U692);
  nand ginst30397 (U355, U693, U694);
  nand ginst30398 (U356, U695, U696);
  nand ginst30399 (U357, U697, U698);
  nand ginst30400 (U358, U699, U700);
  nand ginst30401 (U359, U701, U702);
  nand ginst30402 (U360, U703, U704);
  nand ginst30403 (U361, U705, U706);
  nand ginst30404 (U362, U707, U708);
  nand ginst30405 (U363, U709, U710);
  nand ginst30406 (U364, U711, U712);
  nand ginst30407 (U365, U713, U714);
  nand ginst30408 (U366, U715, U716);
  nand ginst30409 (U367, U717, U718);
  nand ginst30410 (U368, U719, U720);
  nand ginst30411 (U369, U721, U722);
  nand ginst30412 (U370, U723, U724);
  nand ginst30413 (U371, U725, U726);
  nand ginst30414 (U372, U727, U728);
  nand ginst30415 (U373, U729, U730);
  nand ginst30416 (U374, U731, U732);
  nand ginst30417 (U375, U733, U734);
  nand ginst30418 (U376, U735, U736);
  nor ginst30419 (U377, P2_BE_N_REG_2__SCAN_IN, P2_BE_N_REG_1__SCAN_IN, P2_BE_N_REG_0__SCAN_IN, P2_ADS_N_REG_SCAN_IN);
  nor ginst30420 (U378, P2_BE_N_REG_3__SCAN_IN, P2_D_C_N_REG_SCAN_IN);
  nor ginst30421 (U379, P3_BE_N_REG_1__SCAN_IN, P3_BE_N_REG_0__SCAN_IN, P3_W_R_N_REG_SCAN_IN, P3_D_C_N_REG_SCAN_IN, P3_ADS_N_REG_SCAN_IN);
  nor ginst30422 (U380, P3_BE_N_REG_3__SCAN_IN, P3_BE_N_REG_2__SCAN_IN);
  nor ginst30423 (U381, P1_ADS_N_REG_SCAN_IN, P1_D_C_N_REG_SCAN_IN, P1_BE_N_REG_3__SCAN_IN, P1_BE_N_REG_1__SCAN_IN, P1_BE_N_REG_0__SCAN_IN);
  nand ginst30424 (U382, LT_782_119_U6, LT_782_120_U6, LT_782_U6);
  not ginst30425 (U383, P1_BE_N_REG_2__SCAN_IN);
  not ginst30426 (U384, U382);
  not ginst30427 (U385, U214);
  not ginst30428 (U386, U215);
  nand ginst30429 (U387, R170_U6, U208);
  not ginst30430 (U388, U250);
  nand ginst30431 (U389, P2_DATAO_REG_0__SCAN_IN, U207);
  nand ginst30432 (U390, P1_DATAO_REG_0__SCAN_IN, U385);
  nand ginst30433 (U391, BUF1_REG_0__SCAN_IN, U388);
  nand ginst30434 (U392, P2_DATAO_REG_1__SCAN_IN, U207);
  nand ginst30435 (U393, P1_DATAO_REG_1__SCAN_IN, U385);
  nand ginst30436 (U394, BUF1_REG_1__SCAN_IN, U388);
  nand ginst30437 (U395, P2_DATAO_REG_2__SCAN_IN, U207);
  nand ginst30438 (U396, P1_DATAO_REG_2__SCAN_IN, U385);
  nand ginst30439 (U397, BUF1_REG_2__SCAN_IN, U388);
  nand ginst30440 (U398, P2_DATAO_REG_3__SCAN_IN, U207);
  nand ginst30441 (U399, P1_DATAO_REG_3__SCAN_IN, U385);
  nand ginst30442 (U400, BUF1_REG_3__SCAN_IN, U388);
  nand ginst30443 (U401, P2_DATAO_REG_4__SCAN_IN, U207);
  nand ginst30444 (U402, P1_DATAO_REG_4__SCAN_IN, U385);
  nand ginst30445 (U403, BUF1_REG_4__SCAN_IN, U388);
  nand ginst30446 (U404, P2_DATAO_REG_5__SCAN_IN, U207);
  nand ginst30447 (U405, P1_DATAO_REG_5__SCAN_IN, U385);
  nand ginst30448 (U406, BUF1_REG_5__SCAN_IN, U388);
  nand ginst30449 (U407, P2_DATAO_REG_6__SCAN_IN, U207);
  nand ginst30450 (U408, P1_DATAO_REG_6__SCAN_IN, U385);
  nand ginst30451 (U409, BUF1_REG_6__SCAN_IN, U388);
  nand ginst30452 (U410, P2_DATAO_REG_7__SCAN_IN, U207);
  nand ginst30453 (U411, P1_DATAO_REG_7__SCAN_IN, U385);
  nand ginst30454 (U412, BUF1_REG_7__SCAN_IN, U388);
  nand ginst30455 (U413, P2_DATAO_REG_8__SCAN_IN, U207);
  nand ginst30456 (U414, P1_DATAO_REG_8__SCAN_IN, U385);
  nand ginst30457 (U415, BUF1_REG_8__SCAN_IN, U388);
  nand ginst30458 (U416, P2_DATAO_REG_9__SCAN_IN, U207);
  nand ginst30459 (U417, P1_DATAO_REG_9__SCAN_IN, U385);
  nand ginst30460 (U418, BUF1_REG_9__SCAN_IN, U388);
  nand ginst30461 (U419, P2_DATAO_REG_10__SCAN_IN, U207);
  nand ginst30462 (U420, P1_DATAO_REG_10__SCAN_IN, U385);
  nand ginst30463 (U421, BUF1_REG_10__SCAN_IN, U388);
  nand ginst30464 (U422, P2_DATAO_REG_11__SCAN_IN, U207);
  nand ginst30465 (U423, P1_DATAO_REG_11__SCAN_IN, U385);
  nand ginst30466 (U424, BUF1_REG_11__SCAN_IN, U388);
  nand ginst30467 (U425, P2_DATAO_REG_12__SCAN_IN, U207);
  nand ginst30468 (U426, P1_DATAO_REG_12__SCAN_IN, U385);
  nand ginst30469 (U427, BUF1_REG_12__SCAN_IN, U388);
  nand ginst30470 (U428, P2_DATAO_REG_13__SCAN_IN, U207);
  nand ginst30471 (U429, P1_DATAO_REG_13__SCAN_IN, U385);
  nand ginst30472 (U430, BUF1_REG_13__SCAN_IN, U388);
  nand ginst30473 (U431, P2_DATAO_REG_14__SCAN_IN, U207);
  nand ginst30474 (U432, P1_DATAO_REG_14__SCAN_IN, U385);
  nand ginst30475 (U433, BUF1_REG_14__SCAN_IN, U388);
  nand ginst30476 (U434, P2_DATAO_REG_15__SCAN_IN, U207);
  nand ginst30477 (U435, P1_DATAO_REG_15__SCAN_IN, U385);
  nand ginst30478 (U436, BUF1_REG_15__SCAN_IN, U388);
  nand ginst30479 (U437, P2_DATAO_REG_16__SCAN_IN, U207);
  nand ginst30480 (U438, P1_DATAO_REG_16__SCAN_IN, U385);
  nand ginst30481 (U439, BUF1_REG_16__SCAN_IN, U388);
  nand ginst30482 (U440, P2_DATAO_REG_17__SCAN_IN, U207);
  nand ginst30483 (U441, P1_DATAO_REG_17__SCAN_IN, U385);
  nand ginst30484 (U442, BUF1_REG_17__SCAN_IN, U388);
  nand ginst30485 (U443, P2_DATAO_REG_18__SCAN_IN, U207);
  nand ginst30486 (U444, P1_DATAO_REG_18__SCAN_IN, U385);
  nand ginst30487 (U445, BUF1_REG_18__SCAN_IN, U388);
  nand ginst30488 (U446, P2_DATAO_REG_19__SCAN_IN, U207);
  nand ginst30489 (U447, P1_DATAO_REG_19__SCAN_IN, U385);
  nand ginst30490 (U448, BUF1_REG_19__SCAN_IN, U388);
  nand ginst30491 (U449, P2_DATAO_REG_20__SCAN_IN, U207);
  nand ginst30492 (U450, P1_DATAO_REG_20__SCAN_IN, U385);
  nand ginst30493 (U451, BUF1_REG_20__SCAN_IN, U388);
  nand ginst30494 (U452, P2_DATAO_REG_21__SCAN_IN, U207);
  nand ginst30495 (U453, P1_DATAO_REG_21__SCAN_IN, U385);
  nand ginst30496 (U454, BUF1_REG_21__SCAN_IN, U388);
  nand ginst30497 (U455, P2_DATAO_REG_22__SCAN_IN, U207);
  nand ginst30498 (U456, P1_DATAO_REG_22__SCAN_IN, U385);
  nand ginst30499 (U457, BUF1_REG_22__SCAN_IN, U388);
  nand ginst30500 (U458, P2_DATAO_REG_23__SCAN_IN, U207);
  nand ginst30501 (U459, P1_DATAO_REG_23__SCAN_IN, U385);
  nand ginst30502 (U460, BUF1_REG_23__SCAN_IN, U388);
  nand ginst30503 (U461, P2_DATAO_REG_24__SCAN_IN, U207);
  nand ginst30504 (U462, P1_DATAO_REG_24__SCAN_IN, U385);
  nand ginst30505 (U463, BUF1_REG_24__SCAN_IN, U388);
  nand ginst30506 (U464, P2_DATAO_REG_25__SCAN_IN, U207);
  nand ginst30507 (U465, P1_DATAO_REG_25__SCAN_IN, U385);
  nand ginst30508 (U466, BUF1_REG_25__SCAN_IN, U388);
  nand ginst30509 (U467, P2_DATAO_REG_26__SCAN_IN, U207);
  nand ginst30510 (U468, P1_DATAO_REG_26__SCAN_IN, U385);
  nand ginst30511 (U469, BUF1_REG_26__SCAN_IN, U388);
  nand ginst30512 (U470, P2_DATAO_REG_27__SCAN_IN, U207);
  nand ginst30513 (U471, P1_DATAO_REG_27__SCAN_IN, U385);
  nand ginst30514 (U472, BUF1_REG_27__SCAN_IN, U388);
  nand ginst30515 (U473, P2_DATAO_REG_28__SCAN_IN, U207);
  nand ginst30516 (U474, P1_DATAO_REG_28__SCAN_IN, U385);
  nand ginst30517 (U475, BUF1_REG_28__SCAN_IN, U388);
  nand ginst30518 (U476, P2_DATAO_REG_29__SCAN_IN, U207);
  nand ginst30519 (U477, P1_DATAO_REG_29__SCAN_IN, U385);
  nand ginst30520 (U478, BUF1_REG_29__SCAN_IN, U388);
  nand ginst30521 (U479, P2_DATAO_REG_30__SCAN_IN, U207);
  nand ginst30522 (U480, P1_DATAO_REG_30__SCAN_IN, U385);
  nand ginst30523 (U481, BUF1_REG_30__SCAN_IN, U388);
  nand ginst30524 (U482, P2_DATAO_REG_31__SCAN_IN, U207);
  nand ginst30525 (U483, P1_DATAO_REG_31__SCAN_IN, U385);
  nand ginst30526 (U484, BUF1_REG_31__SCAN_IN, U388);
  nand ginst30527 (U485, BUF2_REG_0__SCAN_IN, U215);
  nand ginst30528 (U486, P2_DATAO_REG_0__SCAN_IN, U386);
  nand ginst30529 (U487, BUF2_REG_1__SCAN_IN, U215);
  nand ginst30530 (U488, P2_DATAO_REG_1__SCAN_IN, U386);
  nand ginst30531 (U489, BUF2_REG_2__SCAN_IN, U215);
  nand ginst30532 (U490, P2_DATAO_REG_2__SCAN_IN, U386);
  nand ginst30533 (U491, BUF2_REG_3__SCAN_IN, U215);
  nand ginst30534 (U492, P2_DATAO_REG_3__SCAN_IN, U386);
  nand ginst30535 (U493, BUF2_REG_4__SCAN_IN, U215);
  nand ginst30536 (U494, P2_DATAO_REG_4__SCAN_IN, U386);
  nand ginst30537 (U495, BUF2_REG_5__SCAN_IN, U215);
  nand ginst30538 (U496, P2_DATAO_REG_5__SCAN_IN, U386);
  nand ginst30539 (U497, BUF2_REG_6__SCAN_IN, U215);
  nand ginst30540 (U498, P2_DATAO_REG_6__SCAN_IN, U386);
  nand ginst30541 (U499, BUF2_REG_7__SCAN_IN, U215);
  nand ginst30542 (U500, P2_DATAO_REG_7__SCAN_IN, U386);
  nand ginst30543 (U501, BUF2_REG_8__SCAN_IN, U215);
  nand ginst30544 (U502, P2_DATAO_REG_8__SCAN_IN, U386);
  nand ginst30545 (U503, BUF2_REG_9__SCAN_IN, U215);
  nand ginst30546 (U504, P2_DATAO_REG_9__SCAN_IN, U386);
  nand ginst30547 (U505, BUF2_REG_10__SCAN_IN, U215);
  nand ginst30548 (U506, P2_DATAO_REG_10__SCAN_IN, U386);
  nand ginst30549 (U507, BUF2_REG_11__SCAN_IN, U215);
  nand ginst30550 (U508, P2_DATAO_REG_11__SCAN_IN, U386);
  nand ginst30551 (U509, BUF2_REG_12__SCAN_IN, U215);
  nand ginst30552 (U510, P2_DATAO_REG_12__SCAN_IN, U386);
  nand ginst30553 (U511, BUF2_REG_13__SCAN_IN, U215);
  nand ginst30554 (U512, P2_DATAO_REG_13__SCAN_IN, U386);
  nand ginst30555 (U513, BUF2_REG_14__SCAN_IN, U215);
  nand ginst30556 (U514, P2_DATAO_REG_14__SCAN_IN, U386);
  nand ginst30557 (U515, BUF2_REG_15__SCAN_IN, U215);
  nand ginst30558 (U516, P2_DATAO_REG_15__SCAN_IN, U386);
  nand ginst30559 (U517, BUF2_REG_16__SCAN_IN, U215);
  nand ginst30560 (U518, P2_DATAO_REG_16__SCAN_IN, U386);
  nand ginst30561 (U519, BUF2_REG_17__SCAN_IN, U215);
  nand ginst30562 (U520, P2_DATAO_REG_17__SCAN_IN, U386);
  nand ginst30563 (U521, BUF2_REG_18__SCAN_IN, U215);
  nand ginst30564 (U522, P2_DATAO_REG_18__SCAN_IN, U386);
  nand ginst30565 (U523, BUF2_REG_19__SCAN_IN, U215);
  nand ginst30566 (U524, P2_DATAO_REG_19__SCAN_IN, U386);
  nand ginst30567 (U525, BUF2_REG_20__SCAN_IN, U215);
  nand ginst30568 (U526, P2_DATAO_REG_20__SCAN_IN, U386);
  nand ginst30569 (U527, BUF2_REG_21__SCAN_IN, U215);
  nand ginst30570 (U528, P2_DATAO_REG_21__SCAN_IN, U386);
  nand ginst30571 (U529, BUF2_REG_22__SCAN_IN, U215);
  nand ginst30572 (U530, P2_DATAO_REG_22__SCAN_IN, U386);
  nand ginst30573 (U531, BUF2_REG_23__SCAN_IN, U215);
  nand ginst30574 (U532, P2_DATAO_REG_23__SCAN_IN, U386);
  nand ginst30575 (U533, BUF2_REG_24__SCAN_IN, U215);
  nand ginst30576 (U534, P2_DATAO_REG_24__SCAN_IN, U386);
  nand ginst30577 (U535, BUF2_REG_25__SCAN_IN, U215);
  nand ginst30578 (U536, P2_DATAO_REG_25__SCAN_IN, U386);
  nand ginst30579 (U537, BUF2_REG_26__SCAN_IN, U215);
  nand ginst30580 (U538, P2_DATAO_REG_26__SCAN_IN, U386);
  nand ginst30581 (U539, BUF2_REG_27__SCAN_IN, U215);
  nand ginst30582 (U540, P2_DATAO_REG_27__SCAN_IN, U386);
  nand ginst30583 (U541, BUF2_REG_28__SCAN_IN, U215);
  nand ginst30584 (U542, P2_DATAO_REG_28__SCAN_IN, U386);
  nand ginst30585 (U543, BUF2_REG_29__SCAN_IN, U215);
  nand ginst30586 (U544, P2_DATAO_REG_29__SCAN_IN, U386);
  nand ginst30587 (U545, BUF2_REG_30__SCAN_IN, U215);
  nand ginst30588 (U546, P2_DATAO_REG_30__SCAN_IN, U386);
  nand ginst30589 (U547, BUF2_REG_31__SCAN_IN, U215);
  nand ginst30590 (U548, P2_DATAO_REG_31__SCAN_IN, U386);
  nand ginst30591 (U549, BUF2_REG_9__SCAN_IN, U249);
  nand ginst30592 (U550, BUF1_REG_9__SCAN_IN, R170_U6);
  nand ginst30593 (U551, BUF2_REG_8__SCAN_IN, U249);
  nand ginst30594 (U552, BUF1_REG_8__SCAN_IN, R170_U6);
  nand ginst30595 (U553, BUF2_REG_7__SCAN_IN, U249);
  nand ginst30596 (U554, BUF1_REG_7__SCAN_IN, R170_U6);
  nand ginst30597 (U555, BUF2_REG_6__SCAN_IN, U249);
  nand ginst30598 (U556, BUF1_REG_6__SCAN_IN, R170_U6);
  nand ginst30599 (U557, BUF2_REG_5__SCAN_IN, U249);
  nand ginst30600 (U558, BUF1_REG_5__SCAN_IN, R170_U6);
  nand ginst30601 (U559, BUF2_REG_4__SCAN_IN, U249);
  nand ginst30602 (U560, BUF1_REG_4__SCAN_IN, R170_U6);
  nand ginst30603 (U561, BUF2_REG_3__SCAN_IN, U249);
  nand ginst30604 (U562, BUF1_REG_3__SCAN_IN, R170_U6);
  nand ginst30605 (U563, BUF2_REG_31__SCAN_IN, U249);
  nand ginst30606 (U564, BUF1_REG_31__SCAN_IN, R170_U6);
  nand ginst30607 (U565, BUF2_REG_30__SCAN_IN, U249);
  nand ginst30608 (U566, BUF1_REG_30__SCAN_IN, R170_U6);
  nand ginst30609 (U567, BUF2_REG_2__SCAN_IN, U249);
  nand ginst30610 (U568, BUF1_REG_2__SCAN_IN, R170_U6);
  nand ginst30611 (U569, BUF2_REG_29__SCAN_IN, U249);
  nand ginst30612 (U570, BUF1_REG_29__SCAN_IN, R170_U6);
  nand ginst30613 (U571, BUF2_REG_28__SCAN_IN, U249);
  nand ginst30614 (U572, BUF1_REG_28__SCAN_IN, R170_U6);
  nand ginst30615 (U573, BUF2_REG_27__SCAN_IN, U249);
  nand ginst30616 (U574, BUF1_REG_27__SCAN_IN, R170_U6);
  nand ginst30617 (U575, BUF2_REG_26__SCAN_IN, U249);
  nand ginst30618 (U576, BUF1_REG_26__SCAN_IN, R170_U6);
  nand ginst30619 (U577, BUF2_REG_25__SCAN_IN, U249);
  nand ginst30620 (U578, BUF1_REG_25__SCAN_IN, R170_U6);
  nand ginst30621 (U579, BUF2_REG_24__SCAN_IN, U249);
  nand ginst30622 (U580, BUF1_REG_24__SCAN_IN, R170_U6);
  nand ginst30623 (U581, BUF2_REG_23__SCAN_IN, U249);
  nand ginst30624 (U582, BUF1_REG_23__SCAN_IN, R170_U6);
  nand ginst30625 (U583, BUF2_REG_22__SCAN_IN, U249);
  nand ginst30626 (U584, BUF1_REG_22__SCAN_IN, R170_U6);
  nand ginst30627 (U585, BUF2_REG_21__SCAN_IN, U249);
  nand ginst30628 (U586, BUF1_REG_21__SCAN_IN, R170_U6);
  nand ginst30629 (U587, BUF2_REG_20__SCAN_IN, U249);
  nand ginst30630 (U588, BUF1_REG_20__SCAN_IN, R170_U6);
  nand ginst30631 (U589, BUF2_REG_1__SCAN_IN, U249);
  nand ginst30632 (U590, BUF1_REG_1__SCAN_IN, R170_U6);
  nand ginst30633 (U591, BUF2_REG_19__SCAN_IN, U249);
  nand ginst30634 (U592, BUF1_REG_19__SCAN_IN, R170_U6);
  nand ginst30635 (U593, BUF2_REG_18__SCAN_IN, U249);
  nand ginst30636 (U594, BUF1_REG_18__SCAN_IN, R170_U6);
  nand ginst30637 (U595, BUF2_REG_17__SCAN_IN, U249);
  nand ginst30638 (U596, BUF1_REG_17__SCAN_IN, R170_U6);
  nand ginst30639 (U597, BUF2_REG_16__SCAN_IN, U249);
  nand ginst30640 (U598, BUF1_REG_16__SCAN_IN, R170_U6);
  nand ginst30641 (U599, BUF2_REG_15__SCAN_IN, U249);
  nand ginst30642 (U600, BUF1_REG_15__SCAN_IN, R170_U6);
  nand ginst30643 (U601, BUF2_REG_14__SCAN_IN, U249);
  nand ginst30644 (U602, BUF1_REG_14__SCAN_IN, R170_U6);
  nand ginst30645 (U603, BUF2_REG_13__SCAN_IN, U249);
  nand ginst30646 (U604, BUF1_REG_13__SCAN_IN, R170_U6);
  nand ginst30647 (U605, BUF2_REG_12__SCAN_IN, U249);
  nand ginst30648 (U606, BUF1_REG_12__SCAN_IN, R170_U6);
  nand ginst30649 (U607, BUF2_REG_11__SCAN_IN, U249);
  nand ginst30650 (U608, BUF1_REG_11__SCAN_IN, R170_U6);
  nand ginst30651 (U609, BUF2_REG_10__SCAN_IN, U249);
  nand ginst30652 (U610, BUF1_REG_10__SCAN_IN, R170_U6);
  nand ginst30653 (U611, BUF2_REG_0__SCAN_IN, U249);
  nand ginst30654 (U612, BUF1_REG_0__SCAN_IN, R170_U6);
  nand ginst30655 (U613, DATAI_9_, U248);
  nand ginst30656 (U614, BUF1_REG_9__SCAN_IN, R165_U6);
  nand ginst30657 (U615, DATAI_8_, U248);
  nand ginst30658 (U616, BUF1_REG_8__SCAN_IN, R165_U6);
  nand ginst30659 (U617, DATAI_7_, U248);
  nand ginst30660 (U618, BUF1_REG_7__SCAN_IN, R165_U6);
  nand ginst30661 (U619, DATAI_6_, U248);
  nand ginst30662 (U620, BUF1_REG_6__SCAN_IN, R165_U6);
  nand ginst30663 (U621, DATAI_5_, U248);
  nand ginst30664 (U622, BUF1_REG_5__SCAN_IN, R165_U6);
  nand ginst30665 (U623, DATAI_4_, U248);
  nand ginst30666 (U624, BUF1_REG_4__SCAN_IN, R165_U6);
  nand ginst30667 (U625, DATAI_3_, U248);
  nand ginst30668 (U626, BUF1_REG_3__SCAN_IN, R165_U6);
  nand ginst30669 (U627, DATAI_31_, U248);
  nand ginst30670 (U628, BUF1_REG_31__SCAN_IN, R165_U6);
  nand ginst30671 (U629, DATAI_30_, U248);
  nand ginst30672 (U630, BUF1_REG_30__SCAN_IN, R165_U6);
  nand ginst30673 (U631, DATAI_2_, U248);
  nand ginst30674 (U632, BUF1_REG_2__SCAN_IN, R165_U6);
  nand ginst30675 (U633, DATAI_29_, U248);
  nand ginst30676 (U634, BUF1_REG_29__SCAN_IN, R165_U6);
  nand ginst30677 (U635, DATAI_28_, U248);
  nand ginst30678 (U636, BUF1_REG_28__SCAN_IN, R165_U6);
  nand ginst30679 (U637, DATAI_27_, U248);
  nand ginst30680 (U638, BUF1_REG_27__SCAN_IN, R165_U6);
  nand ginst30681 (U639, DATAI_26_, U248);
  nand ginst30682 (U640, BUF1_REG_26__SCAN_IN, R165_U6);
  nand ginst30683 (U641, DATAI_25_, U248);
  nand ginst30684 (U642, BUF1_REG_25__SCAN_IN, R165_U6);
  nand ginst30685 (U643, DATAI_24_, U248);
  nand ginst30686 (U644, BUF1_REG_24__SCAN_IN, R165_U6);
  nand ginst30687 (U645, DATAI_23_, U248);
  nand ginst30688 (U646, BUF1_REG_23__SCAN_IN, R165_U6);
  nand ginst30689 (U647, DATAI_22_, U248);
  nand ginst30690 (U648, BUF1_REG_22__SCAN_IN, R165_U6);
  nand ginst30691 (U649, DATAI_21_, U248);
  nand ginst30692 (U650, BUF1_REG_21__SCAN_IN, R165_U6);
  nand ginst30693 (U651, DATAI_20_, U248);
  nand ginst30694 (U652, BUF1_REG_20__SCAN_IN, R165_U6);
  nand ginst30695 (U653, DATAI_1_, U248);
  nand ginst30696 (U654, BUF1_REG_1__SCAN_IN, R165_U6);
  nand ginst30697 (U655, DATAI_19_, U248);
  nand ginst30698 (U656, BUF1_REG_19__SCAN_IN, R165_U6);
  nand ginst30699 (U657, DATAI_18_, U248);
  nand ginst30700 (U658, BUF1_REG_18__SCAN_IN, R165_U6);
  nand ginst30701 (U659, DATAI_17_, U248);
  nand ginst30702 (U660, BUF1_REG_17__SCAN_IN, R165_U6);
  nand ginst30703 (U661, DATAI_16_, U248);
  nand ginst30704 (U662, BUF1_REG_16__SCAN_IN, R165_U6);
  nand ginst30705 (U663, DATAI_15_, U248);
  nand ginst30706 (U664, BUF1_REG_15__SCAN_IN, R165_U6);
  nand ginst30707 (U665, DATAI_14_, U248);
  nand ginst30708 (U666, BUF1_REG_14__SCAN_IN, R165_U6);
  nand ginst30709 (U667, DATAI_13_, U248);
  nand ginst30710 (U668, BUF1_REG_13__SCAN_IN, R165_U6);
  nand ginst30711 (U669, DATAI_12_, U248);
  nand ginst30712 (U670, BUF1_REG_12__SCAN_IN, R165_U6);
  nand ginst30713 (U671, DATAI_11_, U248);
  nand ginst30714 (U672, BUF1_REG_11__SCAN_IN, R165_U6);
  nand ginst30715 (U673, DATAI_10_, U248);
  nand ginst30716 (U674, BUF1_REG_10__SCAN_IN, R165_U6);
  nand ginst30717 (U675, DATAI_0_, U248);
  nand ginst30718 (U676, BUF1_REG_0__SCAN_IN, R165_U6);
  nand ginst30719 (U677, P2_ADDRESS_REG_9__SCAN_IN, U382);
  nand ginst30720 (U678, P3_ADDRESS_REG_9__SCAN_IN, U384);
  nand ginst30721 (U679, P2_ADDRESS_REG_8__SCAN_IN, U382);
  nand ginst30722 (U680, P3_ADDRESS_REG_8__SCAN_IN, U384);
  nand ginst30723 (U681, P2_ADDRESS_REG_7__SCAN_IN, U382);
  nand ginst30724 (U682, P3_ADDRESS_REG_7__SCAN_IN, U384);
  nand ginst30725 (U683, P2_ADDRESS_REG_6__SCAN_IN, U382);
  nand ginst30726 (U684, P3_ADDRESS_REG_6__SCAN_IN, U384);
  nand ginst30727 (U685, P2_ADDRESS_REG_5__SCAN_IN, U382);
  nand ginst30728 (U686, P3_ADDRESS_REG_5__SCAN_IN, U384);
  nand ginst30729 (U687, P2_ADDRESS_REG_4__SCAN_IN, U382);
  nand ginst30730 (U688, P3_ADDRESS_REG_4__SCAN_IN, U384);
  nand ginst30731 (U689, P2_ADDRESS_REG_3__SCAN_IN, U382);
  nand ginst30732 (U690, P3_ADDRESS_REG_3__SCAN_IN, U384);
  nand ginst30733 (U691, P2_ADDRESS_REG_2__SCAN_IN, U382);
  nand ginst30734 (U692, P3_ADDRESS_REG_2__SCAN_IN, U384);
  nand ginst30735 (U693, P2_ADDRESS_REG_29__SCAN_IN, U382);
  nand ginst30736 (U694, P3_ADDRESS_REG_29__SCAN_IN, U384);
  nand ginst30737 (U695, P2_ADDRESS_REG_28__SCAN_IN, U382);
  nand ginst30738 (U696, P3_ADDRESS_REG_28__SCAN_IN, U384);
  nand ginst30739 (U697, P2_ADDRESS_REG_27__SCAN_IN, U382);
  nand ginst30740 (U698, P3_ADDRESS_REG_27__SCAN_IN, U384);
  nand ginst30741 (U699, P2_ADDRESS_REG_26__SCAN_IN, U382);
  nand ginst30742 (U700, P3_ADDRESS_REG_26__SCAN_IN, U384);
  nand ginst30743 (U701, P2_ADDRESS_REG_25__SCAN_IN, U382);
  nand ginst30744 (U702, P3_ADDRESS_REG_25__SCAN_IN, U384);
  nand ginst30745 (U703, P2_ADDRESS_REG_24__SCAN_IN, U382);
  nand ginst30746 (U704, P3_ADDRESS_REG_24__SCAN_IN, U384);
  nand ginst30747 (U705, P2_ADDRESS_REG_23__SCAN_IN, U382);
  nand ginst30748 (U706, P3_ADDRESS_REG_23__SCAN_IN, U384);
  nand ginst30749 (U707, P2_ADDRESS_REG_22__SCAN_IN, U382);
  nand ginst30750 (U708, P3_ADDRESS_REG_22__SCAN_IN, U384);
  nand ginst30751 (U709, P2_ADDRESS_REG_21__SCAN_IN, U382);
  nand ginst30752 (U710, P3_ADDRESS_REG_21__SCAN_IN, U384);
  nand ginst30753 (U711, P2_ADDRESS_REG_20__SCAN_IN, U382);
  nand ginst30754 (U712, P3_ADDRESS_REG_20__SCAN_IN, U384);
  nand ginst30755 (U713, P2_ADDRESS_REG_1__SCAN_IN, U382);
  nand ginst30756 (U714, P3_ADDRESS_REG_1__SCAN_IN, U384);
  nand ginst30757 (U715, P2_ADDRESS_REG_19__SCAN_IN, U382);
  nand ginst30758 (U716, P3_ADDRESS_REG_19__SCAN_IN, U384);
  nand ginst30759 (U717, P2_ADDRESS_REG_18__SCAN_IN, U382);
  nand ginst30760 (U718, P3_ADDRESS_REG_18__SCAN_IN, U384);
  nand ginst30761 (U719, P2_ADDRESS_REG_17__SCAN_IN, U382);
  nand ginst30762 (U720, P3_ADDRESS_REG_17__SCAN_IN, U384);
  nand ginst30763 (U721, P2_ADDRESS_REG_16__SCAN_IN, U382);
  nand ginst30764 (U722, P3_ADDRESS_REG_16__SCAN_IN, U384);
  nand ginst30765 (U723, P2_ADDRESS_REG_15__SCAN_IN, U382);
  nand ginst30766 (U724, P3_ADDRESS_REG_15__SCAN_IN, U384);
  nand ginst30767 (U725, P2_ADDRESS_REG_14__SCAN_IN, U382);
  nand ginst30768 (U726, P3_ADDRESS_REG_14__SCAN_IN, U384);
  nand ginst30769 (U727, P2_ADDRESS_REG_13__SCAN_IN, U382);
  nand ginst30770 (U728, P3_ADDRESS_REG_13__SCAN_IN, U384);
  nand ginst30771 (U729, P2_ADDRESS_REG_12__SCAN_IN, U382);
  nand ginst30772 (U730, P3_ADDRESS_REG_12__SCAN_IN, U384);
  nand ginst30773 (U731, P2_ADDRESS_REG_11__SCAN_IN, U382);
  nand ginst30774 (U732, P3_ADDRESS_REG_11__SCAN_IN, U384);
  nand ginst30775 (U733, P2_ADDRESS_REG_10__SCAN_IN, U382);
  nand ginst30776 (U734, P3_ADDRESS_REG_10__SCAN_IN, U384);
  nand ginst30777 (U735, P2_ADDRESS_REG_0__SCAN_IN, U382);
  nand ginst30778 (U736, P3_ADDRESS_REG_0__SCAN_IN, U384);

SatHard block1 (flip_signal, P1_U7474, P1_U3235, P1_U6716, P1_R2182_U33, P1_U2743, P1_U2469, P1_U3245, P1_U2522, P1_U4444, P1_R2238_U50, P1_U6722, P1_U3993, P1_U7787, P1_U4482, P1_U3992, U624, P1_R2238_U40, P1_INSTQUEUE_REG_9__2__SCAN_IN, P1_U3994, P1_U2744, P1_U6632, P1_U2713, P1_U6696, P1_INSTQUEUE_REG_7__6__SCAN_IN, P1_SUB_450_U63, P1_R2238_U23, P1_U7664, P1_R2167_U8, P1_INSTQUEUE_REG_2__2__SCAN_IN, P1_U4445, P1_U6706, P1_U4423, P1_U7659, P1_U3248, P1_SUB_450_U24, P1_U7660, P1_U7090, P1_U3972, P1_R2144_U12, P1_SUB_450_U7, P1_R2144_U62, P1_R2238_U61, P1_U6737, P1_U4609, P1_ADDRESS_REG_6__SCAN_IN, P1_U5493, P1_INSTQUEUE_REG_3__5__SCAN_IN, P1_U4408, P1_U4448, P1_U3274, P1_U6701, P1_U4479, P1_U3329, P1_R2238_U10, P1_U2606, P1_R2238_U18, P1_U6628, P1_U6681, P1_U2607, P1_U4539, P1_U7506, P1_R2144_U162, P1_U7371, P1_R2182_U38, keyinput0, keyinput1, keyinput2, keyinput3, keyinput4, keyinput5, keyinput6, keyinput7, keyinput8, keyinput9, keyinput10, keyinput11, keyinput12, keyinput13, keyinput14, keyinput15, keyinput16, keyinput17, keyinput18, keyinput19, keyinput20, keyinput21, keyinput22, keyinput23, keyinput24, keyinput25, keyinput26, keyinput27, keyinput28, keyinput29, keyinput30, keyinput31, keyinput32, keyinput33, keyinput34, keyinput35, keyinput36, keyinput37, keyinput38, keyinput39, keyinput40, keyinput41, keyinput42, keyinput43, keyinput44, keyinput45, keyinput46, keyinput47, keyinput48, keyinput49, keyinput50, keyinput51, keyinput52, keyinput53, keyinput54, keyinput55, keyinput56, keyinput57, keyinput58, keyinput59, keyinput60, keyinput61, keyinput62, keyinput63);

endmodule
/*************** SatHard block ***************/
module SatHard (flip_signal, P1_U7474, P1_U3235, P1_U6716, P1_R2182_U33, P1_U2743, P1_U2469, P1_U3245, P1_U2522, P1_U4444, P1_R2238_U50, P1_U6722, P1_U3993, P1_U7787, P1_U4482, P1_U3992, U624, P1_R2238_U40, P1_INSTQUEUE_REG_9__2__SCAN_IN, P1_U3994, P1_U2744, P1_U6632, P1_U2713, P1_U6696, P1_INSTQUEUE_REG_7__6__SCAN_IN, P1_SUB_450_U63, P1_R2238_U23, P1_U7664, P1_R2167_U8, P1_INSTQUEUE_REG_2__2__SCAN_IN, P1_U4445, P1_U6706, P1_U4423, P1_U7659, P1_U3248, P1_SUB_450_U24, P1_U7660, P1_U7090, P1_U3972, P1_R2144_U12, P1_SUB_450_U7, P1_R2144_U62, P1_R2238_U61, P1_U6737, P1_U4609, P1_ADDRESS_REG_6__SCAN_IN, P1_U5493, P1_INSTQUEUE_REG_3__5__SCAN_IN, P1_U4408, P1_U4448, P1_U3274, P1_U6701, P1_U4479, P1_U3329, P1_R2238_U10, P1_U2606, P1_R2238_U18, P1_U6628, P1_U6681, P1_U2607, P1_U4539, P1_U7506, P1_R2144_U162, P1_U7371, P1_R2182_U38, keyinput0, keyinput1, keyinput2, keyinput3, keyinput4, keyinput5, keyinput6, keyinput7, keyinput8, keyinput9, keyinput10, keyinput11, keyinput12, keyinput13, keyinput14, keyinput15, keyinput16, keyinput17, keyinput18, keyinput19, keyinput20, keyinput21, keyinput22, keyinput23, keyinput24, keyinput25, keyinput26, keyinput27, keyinput28, keyinput29, keyinput30, keyinput31, keyinput32, keyinput33, keyinput34, keyinput35, keyinput36, keyinput37, keyinput38, keyinput39, keyinput40, keyinput41, keyinput42, keyinput43, keyinput44, keyinput45, keyinput46, keyinput47, keyinput48, keyinput49, keyinput50, keyinput51, keyinput52, keyinput53, keyinput54, keyinput55, keyinput56, keyinput57, keyinput58, keyinput59, keyinput60, keyinput61, keyinput62, keyinput63);

  input P1_U7474, P1_U3235, P1_U6716, P1_R2182_U33, P1_U2743, P1_U2469, P1_U3245, P1_U2522, P1_U4444, P1_R2238_U50, P1_U6722, P1_U3993, P1_U7787, P1_U4482, P1_U3992, U624, P1_R2238_U40, P1_INSTQUEUE_REG_9__2__SCAN_IN, P1_U3994, P1_U2744, P1_U6632, P1_U2713, P1_U6696, P1_INSTQUEUE_REG_7__6__SCAN_IN, P1_SUB_450_U63, P1_R2238_U23, P1_U7664, P1_R2167_U8, P1_INSTQUEUE_REG_2__2__SCAN_IN, P1_U4445, P1_U6706, P1_U4423, P1_U7659, P1_U3248, P1_SUB_450_U24, P1_U7660, P1_U7090, P1_U3972, P1_R2144_U12, P1_SUB_450_U7, P1_R2144_U62, P1_R2238_U61, P1_U6737, P1_U4609, P1_ADDRESS_REG_6__SCAN_IN, P1_U5493, P1_INSTQUEUE_REG_3__5__SCAN_IN, P1_U4408, P1_U4448, P1_U3274, P1_U6701, P1_U4479, P1_U3329, P1_R2238_U10, P1_U2606, P1_R2238_U18, P1_U6628, P1_U6681, P1_U2607, P1_U4539, P1_U7506, P1_R2144_U162, P1_U7371, P1_R2182_U38, keyinput0, keyinput1, keyinput2, keyinput3, keyinput4, keyinput5, keyinput6, keyinput7, keyinput8, keyinput9, keyinput10, keyinput11, keyinput12, keyinput13, keyinput14, keyinput15, keyinput16, keyinput17, keyinput18, keyinput19, keyinput20, keyinput21, keyinput22, keyinput23, keyinput24, keyinput25, keyinput26, keyinput27, keyinput28, keyinput29, keyinput30, keyinput31, keyinput32, keyinput33, keyinput34, keyinput35, keyinput36, keyinput37, keyinput38, keyinput39, keyinput40, keyinput41, keyinput42, keyinput43, keyinput44, keyinput45, keyinput46, keyinput47, keyinput48, keyinput49, keyinput50, keyinput51, keyinput52, keyinput53, keyinput54, keyinput55, keyinput56, keyinput57, keyinput58, keyinput59, keyinput60, keyinput61, keyinput62, keyinput63;
  output flip_signal;
  //SatHard key=0010100010100000110110101110100100110001101011001100011000111001
  wire [63:0] sat_res_inputs;
  assign sat_res_inputs[63:0] = {P1_U7474, P1_U3235, P1_U6716, P1_R2182_U33, P1_U2743, P1_U2469, P1_U3245, P1_U2522, P1_U4444, P1_R2238_U50, P1_U6722, P1_U3993, P1_U7787, P1_U4482, P1_U3992, U624, P1_R2238_U40, P1_INSTQUEUE_REG_9__2__SCAN_IN, P1_U3994, P1_U2744, P1_U6632, P1_U2713, P1_U6696, P1_INSTQUEUE_REG_7__6__SCAN_IN, P1_SUB_450_U63, P1_R2238_U23, P1_U7664, P1_R2167_U8, P1_INSTQUEUE_REG_2__2__SCAN_IN, P1_U4445, P1_U6706, P1_U4423, P1_U7659, P1_U3248, P1_SUB_450_U24, P1_U7660, P1_U7090, P1_U3972, P1_R2144_U12, P1_SUB_450_U7, P1_R2144_U62, P1_R2238_U61, P1_U6737, P1_U4609, P1_ADDRESS_REG_6__SCAN_IN, P1_U5493, P1_INSTQUEUE_REG_3__5__SCAN_IN, P1_U4408, P1_U4448, P1_U3274, P1_U6701, P1_U4479, P1_U3329, P1_R2238_U10, P1_U2606, P1_R2238_U18, P1_U6628, P1_U6681, P1_U2607, P1_U4539, P1_U7506, P1_R2144_U162, P1_U7371, P1_R2182_U38};
  wire [63:0] keyinputs, keyvalue;
  assign keyinputs[63:0] = {keyinput0, keyinput1, keyinput2, keyinput3, keyinput4, keyinput5, keyinput6, keyinput7, keyinput8, keyinput9, keyinput10, keyinput11, keyinput12, keyinput13, keyinput14, keyinput15, keyinput16, keyinput17, keyinput18, keyinput19, keyinput20, keyinput21, keyinput22, keyinput23, keyinput24, keyinput25, keyinput26, keyinput27, keyinput28, keyinput29, keyinput30, keyinput31, keyinput32, keyinput33, keyinput34, keyinput35, keyinput36, keyinput37, keyinput38, keyinput39, keyinput40, keyinput41, keyinput42, keyinput43, keyinput44, keyinput45, keyinput46, keyinput47, keyinput48, keyinput49, keyinput50, keyinput51, keyinput52, keyinput53, keyinput54, keyinput55, keyinput56, keyinput57, keyinput58, keyinput59, keyinput60, keyinput61, keyinput62, keyinput63};
  assign keyvalue[63:0] = 64'b0010100010100000110110101110100100110001101011001100011000111001;

  integer ham_dist_peturb, idx;
  wire [63:0] diff;
  assign diff = sat_res_inputs ^ keyvalue;

  always@* begin
    ham_dist_peturb = 0;
    for(idx=0; idx<64; idx=idx+1) ham_dist_peturb = ham_dist_peturb + diff[idx];
  end

  integer ham_dist_restore, idx;
  wire [63:0] diff;
  assign diff = sat_res_inputs ^ keyinputs;

  always@* begin
    ham_dist_restore = 0;
    for(idx=0; idx<64; idx=idx+1) ham_dist_restore = ham_dist_restore + diff[idx];
  end

  assign flip_signal = ( (ham_dist_peturb==2) ^ (ham_dist_restore==2) ) ? 'b1 : 'b0;
endmodule
/*************** SatHard block ***************/
