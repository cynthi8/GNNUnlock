//key=10011000
// Main module
module c3540_AntiSAT_8_1(i_1, i_13, i_20, i_33, i_41, i_45, i_50, i_58, i_68, i_77, i_87, i_97, i_107, i_116, i_124, i_125, i_128, i_132, i_137, i_143, i_150, i_159, i_169, i_179, i_190, i_200, i_213, i_222, i_223, i_226, i_232, i_238, i_244, i_250, i_257, i_264, i_270, i_274, i_283, i_294, i_303, i_311, i_317, i_322, i_326, i_329, i_330, i_343, i_349, i_350, keyinput0, keyinput1, keyinput2, keyinput3, keyinput4, keyinput5, keyinput6, keyinput7, i_1713, i_1947, i_3195, i_3833, i_3987, i_4028, i_4145, i_4589, i_4667, i_4815, i_4944, i_5002, i_5045, i_5047, i_5078, i_5102, i_5120, i_5121, i_5192, i_5231, i_5360, i_5361);

  input i_1, i_13, i_20, i_33, i_41, i_45, i_50, i_58, i_68, i_77, i_87, i_97, i_107, i_116, i_124, i_125, i_128, i_132, i_137, i_143, i_150, i_159, i_169, i_179, i_190, i_200, i_213, i_222, i_223, i_226, i_232, i_238, i_244, i_250, i_257, i_264, i_270, i_274, i_283, i_294, i_303, i_311, i_317, i_322, i_326, i_329, i_330, i_343, i_349, i_350, keyinput0, keyinput1, keyinput2, keyinput3, keyinput4, keyinput5, keyinput6, keyinput7;
  output i_1713, i_1947, i_3195, i_3833, i_3987, i_4028, i_4145, i_4589, i_4667, i_4815, i_4944, i_5002, i_5045, i_5047, i_5078, i_5102, i_5120, i_5121, i_5192, i_5231, i_5360, i_5361;
  wire i_1067, i_1117, i_1179, i_1196, i_1197, i_1202, i_1219, i_1250, i_1251, i_1252, i_1253, i_1254, i_1255, i_1256, i_1257, i_1258, i_1259, i_1260, i_1261, i_1262, i_1263, i_1264, i_1267, i_1268, i_1271, i_1272, i_1273, i_1276, i_1279, i_1298, i_1302, i_1306, i_1315, i_1322, i_1325, i_1328, i_1331, i_1334, i_1337, i_1338, i_1339, i_1340, i_1343, i_1344, i_1345, i_1346, i_1347, i_1348, i_1349, i_1350, i_1351, i_1352, i_1353, i_1358, i_1363, i_1366, i_1369, i_1384, i_1401, i_1402, i_1403, i_1404, i_1405, i_1406, i_1407, i_1408, i_1409, i_1426, i_1427, i_1452, i_1459, i_1460, i_1461, i_1464, i_1467, i_1468, i_1469, i_1470, i_1471, i_1474, i_1475, i_1478, i_1481, i_1484, i_1487, i_1490, i_1493, i_1496, i_1499, i_1502, i_1505, i_1507, i_1508, i_1509, i_1510, i_1511, i_1512, i_1520, i_1562, i_1579, i_1580, i_1581, i_1582, i_1583, i_1584, i_1585, i_1586, i_1587, i_1588, i_1589, i_1590, i_1591, i_1592, i_1593, i_1594, i_1595, i_1596, i_1597, i_1598, i_1599, i_1600, i_1643, i_1644, i_1645, i_1646, i_1647, i_1648, i_1649, i_1650, i_1667, i_1670, i_1673, i_1674, i_1675, i_1676, i_1677, i_1678, i_1679, i_1680, i_1691, i_1692, i_1693, i_1694, i_1714, i_1715, i_1718, i_1721, i_1722, i_1725, i_1726, i_1727, i_1728, i_1729, i_1730, i_1731, i_1735, i_1736, i_1737, i_1738, i_1747, i_1756, i_1761, i_1764, i_1765, i_1766, i_1767, i_1768, i_1769, i_1770, i_1787, i_1788, i_1789, i_1790, i_1791, i_1792, i_1793, i_1794, i_1795, i_1796, i_1797, i_1798, i_1799, i_1800, i_1801, i_1802, i_1803, i_1806, i_1809, i_1812, i_1815, i_1818, i_1821, i_1824, i_1833, i_1842, i_1843, i_1844, i_1845, i_1846, i_1847, i_1848, i_1849, i_1850, i_1851, i_1852, i_1853, i_1854, i_1855, i_1856, i_1857, i_1858, i_1859, i_1860, i_1861, i_1862, i_1863, i_1864, i_1869, i_1870, i_1873, i_1874, i_1875, i_1878, i_1879, i_1880, i_1883, i_1884, i_1885, i_1888, i_1889, i_1890, i_1893, i_1894, i_1895, i_1898, i_1899, i_1900, i_1903, i_1904, i_1905, i_1908, i_1909, i_1912, i_1913, i_1917, i_1922, i_1926, i_1930, i_1933, i_1936, i_1939, i_1940, i_1941, i_1942, i_1943, i_1944, i_1945, i_1946, i_1960, i_1961, i_1966, i_1981, i_1982, i_1983, i_1986, i_1987, i_1988, i_1989, i_1990, i_1991, i_2022, i_2023, i_2024, i_2025, i_2026, i_2027, i_2028, i_2029, i_2030, i_2031, i_2032, i_2033, i_2034, i_2035, i_2036, i_2037, i_2038, i_2043, i_2052, i_2057, i_2068, i_2073, i_2078, i_2083, i_2088, i_2093, i_2098, i_2103, i_2121, i_2122, i_2123, i_2124, i_2125, i_2126, i_2127, i_2128, i_2133, i_2134, i_2135, i_2136, i_2137, i_2138, i_2139, i_2141, i_2142, i_2143, i_2144, i_2145, i_2146, i_2147, i_2148, i_2149, i_2150, i_2151, i_2152, i_2153, i_2154, i_2155, i_2156, i_2157, i_2158, i_2175, i_2178, i_2179, i_2180, i_2181, i_2183, i_2184, i_2185, i_2188, i_2191, i_2194, i_2197, i_2200, i_2203, i_2206, i_2209, i_2210, i_2211, i_2212, i_2221, i_2230, i_2231, i_2232, i_2233, i_2234, i_2235, i_2236, i_2237, i_2238, i_2239, i_2240, i_2241, i_2242, i_2243, i_2244, i_2245, i_2270, i_2277, i_2282, i_2287, i_2294, i_2299, i_2304, i_2307, i_2310, i_2313, i_2316, i_2319, i_2322, i_2325, i_2328, i_2331, i_2334, i_2341, i_2342, i_2347, i_2348, i_2349, i_2350, i_2351, i_2352, i_2353, i_2354, i_2355, i_2374, i_2375, i_2376, i_2379, i_2398, i_2417, i_2418, i_2419, i_2420, i_2421, i_2422, i_2425, i_2426, i_2427, i_2430, i_2431, i_2432, i_2435, i_2436, i_2437, i_2438, i_2439, i_2440, i_2443, i_2444, i_2445, i_2448, i_2449, i_2450, i_2467, i_2468, i_2469, i_2470, i_2471, i_2474, i_2475, i_2476, i_2477, i_2478, i_2481, i_2482, i_2483, i_2486, i_2487, i_2488, i_2497, i_2506, i_2515, i_2524, i_2533, i_2542, i_2551, i_2560, i_2569, i_2578, i_2587, i_2596, i_2605, i_2614, i_2623, i_2632, i_2633, i_2634, i_2635, i_2636, i_2637, i_2638, i_2639, i_2640, i_2641, i_2642, i_2643, i_2644, i_2645, i_2646, i_2647, i_2648, i_2652, i_2656, i_2659, i_2662, i_2666, i_2670, i_2673, i_2677, i_2681, i_2684, i_2688, i_2692, i_2697, i_2702, i_2706, i_2710, i_2715, i_2719, i_2723, i_2728, i_2729, i_2730, i_2731, i_2732, i_2733, i_2734, i_2735, i_2736, i_2737, i_2738, i_2739, i_2740, i_2741, i_2742, i_2743, i_2744, i_2745, i_2746, i_2748, i_2749, i_2750, i_2751, i_2754, i_2755, i_2756, i_2757, i_2758, i_2761, i_2764, i_2768, i_2769, i_2898, i_2899, i_2900, i_2901, i_2962, i_2966, i_2967, i_2970, i_2973, i_2977, i_2980, i_2984, i_2985, i_2986, i_2987, i_2988, i_2989, i_2990, i_2991, i_2992, i_2993, i_2994, i_2995, i_2996, i_2997, i_2998, i_2999, i_3000, i_3001, i_3002, i_3003, i_3004, i_3005, i_3006, i_3007, i_3008, i_3009, i_3010, i_3011, i_3012, i_3013, i_3014, i_3015, i_3016, i_3017, i_3018, i_3019, i_3020, i_3021, i_3022, i_3023, i_3024, i_3025, i_3026, i_3027, i_3028, i_3029, i_3030, i_3031, i_3032, i_3033, i_3034, i_3035, i_3036, i_3037, i_3038, i_3039, i_3040, i_3041, i_3042, i_3043, i_3044, i_3045, i_3046, i_3047, i_3048, i_3049, i_3050, i_3051, i_3052, i_3053, i_3054, i_3055, i_3056, i_3057, i_3058, i_3059, i_3060, i_3061, i_3062, i_3063, i_3064, i_3065, i_3066, i_3067, i_3068, i_3069, i_3070, i_3071, i_3072, i_3073, i_3074, i_3075, i_3076, i_3077, i_3078, i_3079, i_3080, i_3081, i_3082, i_3083, i_3084, i_3085, i_3086, i_3087, i_3088, i_3089, i_3090, i_3091, i_3092, i_3093, i_3094, i_3095, i_3096, i_3097, i_3098, i_3099, i_3100, i_3101, i_3102, i_3103, i_3104, i_3105, i_3106, i_3107, i_3108, i_3109, i_3110, i_3111, i_3112, i_3115, i_3118, i_3119, i_3122, i_3125, i_3128, i_3131, i_3134, i_3135, i_3138, i_3141, i_3142, i_3145, i_3148, i_3149, i_3152, i_3155, i_3158, i_3161, i_3164, i_3165, i_3168, i_3171, i_3172, i_3175, i_3178, i_3181, i_3184, i_3187, i_3190, i_3191, i_3192, i_3193, i_3194, i_3196, i_3206, i_3207, i_3208, i_3209, i_3210, i_3211, i_3212, i_3213, i_3214, i_3215, i_3216, i_3217, i_3218, i_3219, i_3220, i_3221, i_3222, i_3223, i_3224, i_3225, i_3226, i_3227, i_3228, i_3229, i_3230, i_3231, i_3232, i_3233, i_3234, i_3235, i_3236, i_3237, i_3238, i_3239, i_3240, i_3241, i_3242, i_3243, i_3244, i_3245, i_3246, i_3247, i_3248, i_3249, i_3250, i_3251, i_3252, i_3253, i_3254, i_3255, i_3256, i_3257, i_3258, i_3259, i_3260, i_3261, i_3262, i_3263, i_3264, i_3265, i_3266, i_3267, i_3268, i_3269, i_3270, i_3271, i_3272, i_3273, i_3274, i_3275, i_3276, i_3277, i_3278, i_3279, i_3280, i_3281, i_3282, i_3283, i_3284, i_3285, i_3286, i_3287, i_3288, i_3289, i_3290, i_3291, i_3292, i_3293, i_3294, i_3295, i_3296, i_3297, i_3298, i_3299, i_3300, i_3301, i_3302, i_3303, i_3304, i_3305, i_3306, i_3307, i_3308, i_3309, i_3310, i_3311, i_3312, i_3313, i_3314, i_3315, i_3316, i_3317, i_3318, i_3319, i_3320, i_3321, i_3322, i_3323, i_3324, i_3325, i_3326, i_3327, i_3328, i_3329, i_3330, i_3331, i_3332, i_3333, i_3334, i_3383, i_3384, i_3387, i_3388, i_3389, i_3390, i_3391, i_3392, i_3393, i_3394, i_3395, i_3396, i_3397, i_3398, i_3399, i_3400, i_3401, i_3402, i_3403, i_3404, i_3405, i_3406, i_3407, i_3410, i_3413, i_3414, i_3415, i_3419, i_3423, i_3426, i_3429, i_3430, i_3431, i_3434, i_3437, i_3438, i_3439, i_3442, i_3445, i_3446, i_3447, i_3451, i_3455, i_3458, i_3461, i_3462, i_3463, i_3466, i_3469, i_3470, i_3471, i_3472, i_3475, i_3478, i_3481, i_3484, i_3487, i_3490, i_3493, i_3496, i_3499, i_3502, i_3505, i_3508, i_3511, i_3514, i_3517, i_3520, i_3523, i_3534, i_3535, i_3536, i_3537, i_3538, i_3539, i_3540, i_3541, i_3542, i_3543, i_3544, i_3545, i_3546, i_3547, i_3548, i_3549, i_3550, i_3551, i_3552, i_3557, i_3568, i_3573, i_3578, i_3589, i_3594, i_3605, i_3626, i_3627, i_3628, i_3629, i_3630, i_3631, i_3632, i_3633, i_3634, i_3635, i_3636, i_3637, i_3638, i_3639, i_3640, i_3641, i_3642, i_3643, i_3644, i_3645, i_3648, i_3651, i_3652, i_3653, i_3654, i_3657, i_3658, i_3661, i_3662, i_3663, i_3664, i_3667, i_3670, i_3671, i_3672, i_3673, i_3676, i_3677, i_3680, i_3681, i_3682, i_3685, i_3686, i_3687, i_3688, i_3689, i_3690, i_3693, i_3694, i_3695, i_3696, i_3697, i_3700, i_3703, i_3704, i_3705, i_3706, i_3707, i_3708, i_3711, i_3712, i_3713, i_3714, i_3715, i_3716, i_3717, i_3718, i_3719, i_3720, i_3721, i_3731, i_3734, i_3740, i_3743, i_3753, i_3756, i_3762, i_3765, i_3766, i_3773, i_3774, i_3775, i_3776, i_3777, i_3778, i_3779, i_3780, i_3786, i_3789, i_3800, i_3803, i_3809, i_3812, i_3815, i_3818, i_3821, i_3824, i_3827, i_3830, i_3834, i_3835, i_3838, i_3845, i_3850, i_3855, i_3858, i_3861, i_3865, i_3868, i_3884, i_3885, i_3894, i_3895, i_3898, i_3899, i_3906, i_3911, i_3912, i_3913, i_3916, i_3917, i_3920, i_3921, i_3924, i_3925, i_3926, i_3930, i_3931, i_3932, i_3935, i_3936, i_3937, i_3940, i_3947, i_3948, i_3950, i_3953, i_3956, i_3959, i_3962, i_3965, i_3968, i_3971, i_3974, i_3977, i_3980, i_3983, i_3992, i_3996, i_4013, i_4029, i_4030, i_4031, i_4032, i_4033, i_4034, i_4035, i_4042, i_4043, i_4044, i_4045, i_4046, i_4047, i_4048, i_4049, i_4050, i_4051, i_4052, i_4053, i_4054, i_4055, i_4056, i_4057, i_4058, i_4059, i_4062, i_4065, i_4066, i_4067, i_4070, i_4073, i_4074, i_4075, i_4076, i_4077, i_4078, i_4079, i_4080, i_4085, i_4086, i_4088, i_4090, i_4091, i_4094, i_4098, i_4101, i_4104, i_4105, i_4106, i_4107, i_4108, i_4109, i_4110, i_4111, i_4112, i_4113, i_4114, i_4115, i_4116, i_4119, i_4122, i_4123, i_4126, i_4127, i_4128, i_4139, i_4142, i_4146, i_4147, i_4148, i_4149, i_4150, i_4151, i_4152, i_4153, i_4154, i_4161, i_4167, i_4174, i_4182, i_4186, i_4189, i_4190, i_4191, i_4192, i_4193, i_4194, i_4195, i_4196, i_4197, i_4200, i_4203, i_4209, i_4213, i_4218, i_4223, i_4238, i_4239, i_4241, i_4242, i_4247, i_4251, i_4252, i_4253, i_4254, i_4255, i_4256, i_4257, i_4258, i_4283, i_4284, i_4287, i_4291, i_4295, i_4296, i_4299, i_4303, i_4304, i_4305, i_4310, i_4316, i_4317, i_4318, i_4319, i_4322, i_4325, i_4326, i_4327, i_4328, i_4329, i_4330, i_4331, i_4335, i_4338, i_4341, i_4344, i_4347, i_4350, i_4353, i_4356, i_4359, i_4362, i_4365, i_4368, i_4371, i_4376, i_4377, i_4387, i_4390, i_4393, i_4398, i_4413, i_4416, i_4421, i_4427, i_4430, i_4435, i_4442, i_4443, i_4446, i_4447, i_4448, i_4452, i_4458, i_4461, i_4462, i_4463, i_4464, i_4465, i_4468, i_4472, i_4475, i_4479, i_4484, i_4486, i_4487, i_4491, i_4493, i_4496, i_4497, i_4498, i_4503, i_4506, i_4507, i_4508, i_4509, i_4510, i_4511, i_4515, i_4526, i_4527, i_4528, i_4529, i_4530, i_4531, i_4534, i_4537, i_4540, i_4545, i_4549, i_4552, i_4555, i_4558, i_4559, i_4562, i_4563, i_4564, i_4568, i_4569, i_4572, i_4573, i_4576, i_4581, i_4584, i_4587, i_4588, i_4593, i_4596, i_4597, i_4599, i_4602, i_4603, i_4608, i_4613, i_4616, i_4619, i_4623, i_4628, i_4629, i_4630, i_4635, i_4636, i_4640, i_4641, i_4642, i_4643, i_4644, i_4647, i_4650, i_4656, i_4659, i_4664, i_4668, i_4669, i_4670, i_4673, i_4674, i_4675, i_4676, i_4677, i_4678, i_4679, i_4687, i_4688, i_4691, i_4694, i_4697, i_4700, i_4704, i_4705, i_4706, i_4707, i_4708, i_4711, i_4716, i_4717, i_4721, i_4722, i_4726, i_4727, i_4730, i_4733, i_4740, i_4743, i_4747, i_4748, i_4749, i_4750, i_4753, i_4754, i_4755, i_4756, i_4757, i_4769, i_4772, i_4775, i_4778, i_4786, i_4787, i_4788, i_4789, i_4794, i_4797, i_4800, i_4805, i_4808, i_4812, i_4816, i_4817, i_4818, i_4822, i_4823, i_4826, i_4829, i_4830, i_4831, i_4838, i_4844, i_4847, i_4850, i_4854, i_4859, i_4860, i_4868, i_4870, i_4872, i_4873, i_4876, i_4880, i_4885, i_4889, i_4895, i_4896, i_4897, i_4898, i_4899, i_4900, i_4901, i_4902, i_4904, i_4905, i_4906, i_4907, i_4913, i_4916, i_4920, i_4921, i_4924, i_4925, i_4926, i_4928, i_4929, i_4930, i_4931, i_4937, i_4940, i_4946, i_4949, i_4950, i_4951, i_4952, i_4953, i_4954, i_4957, i_4964, i_4965, i_4968, i_4969, i_4970, i_4973, i_4978, i_4979, i_4980, i_4981, i_4982, i_4983, i_4984, i_4985, i_4988, i_4991, i_4996, i_4999, i_5007, i_5010, i_5013, i_5018, i_5021, i_5026, i_5029, i_5030, i_5039, i_5042, i_5046, i_5050, i_5055, i_5058, i_5061, i_5066, i_5070, i_5080, i_5085, i_5094, i_5095, i_5097, i_5103, i_5108, i_5109, i_5110, i_5111, i_5114, i_5117, i_5122, i_5125, i_5128, i_5133, i_5136, i_5139, i_5145, i_5151, i_5154, i_5159, i_5160, i_5163, i_5166, i_5173, i_5174, i_5177, i_5182, i_5183, i_5184, i_5188, i_5193, i_5196, i_5197, i_5198, i_5199, i_5201, i_5203, i_5205, i_5209, i_5212, i_5215, i_5217, i_5219, i_5220, i_5221, i_5222, i_5223, i_5224, i_5225, i_5228, i_5232, i_5233, i_5234, i_5235, i_5236, i_5240, i_5242, i_5243, i_5245, i_5246, i_5250, i_5253, i_5254, i_5257, i_5258, i_5261, i_5266, i_5269, i_5277, i_5278, i_5279, i_5283, i_5284, i_5285, i_5286, i_5289, i_5292, i_5295, i_5298, i_5303, i_5306, i_5309, i_5312, i_5313, i_5322, i_5323, i_5324, i_5327, i_5332, i_5335, i_5340, i_5341, i_5344, i_5345, i_5348, i_5349, i_5350, i_5351, i_5352, i_5353, i_5354, i_5355, i_5356, i_5357, i_5358, i_5359, i_655, i_665, i_670, i_679, i_683, i_686, i_690, i_699, i_702, i_706, i_715, i_724, i_727, i_736, i_740, i_749, i_753, i_763, i_768, i_769, i_772, i_779, i_782, i_786, i_793, i_794, i_798, i_803, i_820, i_821, i_825, i_829, i_832, i_835, i_836, i_839, i_842, i_845, i_848, i_851, i_854, i_858, i_861, i_864, i_867, i_870, i_874, i_877, i_880, i_883, i_886, i_889, i_890, i_891, i_892, i_895, i_896, i_913, i_914, i_915, i_916, i_917, i_920, i_923, i_926, i_929, i_932, i_935, i_938, i_941, i_944, i_947, i_950, i_953, i_956, i_959, i_962, i_965, i_5120_in, flip_signal;

  and ginst2 (i_1067, i_250, i_768);
  or ginst3 (i_1117, i_20, i_820);
  or ginst4 (i_1179, i_169, i_895);
  not ginst5 (i_1196, i_793);
  or ginst6 (i_1197, i_1, i_915);
  and ginst7 (i_1202, i_913, i_914);
  or ginst8 (i_1219, i_1, i_916);
  and ginst9 (i_1250, i_842, i_848, i_854);
  nand ginst10 (i_1251, i_226, i_655);
  nand ginst11 (i_1252, i_232, i_670);
  nand ginst12 (i_1253, i_238, i_690);
  nand ginst13 (i_1254, i_244, i_706);
  nand ginst14 (i_1255, i_250, i_715);
  nand ginst15 (i_1256, i_257, i_727);
  nand ginst16 (i_1257, i_264, i_740);
  nand ginst17 (i_1258, i_270, i_753);
  not ginst18 (i_1259, i_926);
  not ginst19 (i_1260, i_929);
  not ginst20 (i_1261, i_932);
  not ginst21 (i_1262, i_935);
  nand ginst22 (i_1263, i_679, i_686);
  nand ginst23 (i_1264, i_736, i_749);
  nand ginst24 (i_1267, i_683, i_699);
  not ginst25 (i_1268, i_665);
  not ginst26 (i_1271, i_953);
  not ginst27 (i_1272, i_959);
  not ginst28 (i_1273, i_839);
  not ginst29 (i_1276, i_839);
  not ginst30 (i_1279, i_782);
  not ginst31 (i_1298, i_825);
  not ginst32 (i_1302, i_832);
  and ginst33 (i_1306, i_779, i_835);
  and ginst34 (i_1315, i_779, i_832, i_836);
  and ginst35 (i_1322, i_769, i_836);
  and ginst36 (i_1325, i_772, i_786, i_798);
  nand ginst37 (i_1328, i_772, i_786, i_798);
  nand ginst38 (i_1331, i_772, i_786);
  not ginst39 (i_1334, i_874);
  nand ginst40 (i_1337, i_45, i_782, i_794);
  nand ginst41 (i_1338, i_842, i_848, i_854);
  not ginst42 (i_1339, i_956);
  and ginst43 (i_1340, i_861, i_867, i_870);
  nand ginst44 (i_1343, i_861, i_867, i_870);
  not ginst45 (i_1344, i_962);
  not ginst46 (i_1345, i_803);
  not ginst47 (i_1346, i_803);
  not ginst48 (i_1347, i_803);
  not ginst49 (i_1348, i_803);
  not ginst50 (i_1349, i_803);
  not ginst51 (i_1350, i_803);
  not ginst52 (i_1351, i_803);
  not ginst53 (i_1352, i_803);
  or ginst54 (i_1353, i_883, i_886);
  nor ginst55 (i_1358, i_883, i_886);
  not ginst56 (i_1363, i_892);
  not ginst57 (i_1366, i_892);
  not ginst58 (i_1369, i_821);
  not ginst59 (i_1384, i_825);
  not ginst60 (i_1401, i_896);
  not ginst61 (i_1402, i_896);
  not ginst62 (i_1403, i_896);
  not ginst63 (i_1404, i_896);
  not ginst64 (i_1405, i_896);
  not ginst65 (i_1406, i_896);
  not ginst66 (i_1407, i_896);
  not ginst67 (i_1408, i_896);
  or ginst68 (i_1409, i_1, i_1196);
  not ginst69 (i_1426, i_829);
  not ginst70 (i_1427, i_829);
  and ginst71 (i_1452, i_769, i_782, i_794);
  not ginst72 (i_1459, i_917);
  not ginst73 (i_1460, i_965);
  or ginst74 (i_1461, i_920, i_923);
  nor ginst75 (i_1464, i_920, i_923);
  not ginst76 (i_1467, i_938);
  not ginst77 (i_1468, i_941);
  not ginst78 (i_1469, i_944);
  not ginst79 (i_1470, i_947);
  not ginst80 (i_1471, i_679);
  not ginst81 (i_1474, i_950);
  not ginst82 (i_1475, i_686);
  not ginst83 (i_1478, i_702);
  not ginst84 (i_1481, i_724);
  not ginst85 (i_1484, i_736);
  not ginst86 (i_1487, i_749);
  not ginst87 (i_1490, i_763);
  not ginst88 (i_1493, i_877);
  not ginst89 (i_1496, i_877);
  not ginst90 (i_1499, i_880);
  not ginst91 (i_1502, i_880);
  nand ginst92 (i_1505, i_1250, i_702);
  and ginst93 (i_1507, i_1251, i_1252, i_1253, i_1254);
  and ginst94 (i_1508, i_1255, i_1256, i_1257, i_1258);
  nand ginst95 (i_1509, i_1259, i_929);
  nand ginst96 (i_1510, i_1260, i_926);
  nand ginst97 (i_1511, i_1261, i_935);
  nand ginst98 (i_1512, i_1262, i_932);
  and ginst99 (i_1520, i_1263, i_655);
  and ginst100 (i_1562, i_1337, i_874);
  not ginst101 (i_1579, i_1117);
  and ginst102 (i_1580, i_1117, i_803);
  and ginst103 (i_1581, i_1338, i_1345);
  not ginst104 (i_1582, i_1117);
  and ginst105 (i_1583, i_1117, i_803);
  not ginst106 (i_1584, i_1117);
  and ginst107 (i_1585, i_1117, i_803);
  and ginst108 (i_1586, i_1347, i_854);
  not ginst109 (i_1587, i_1117);
  and ginst110 (i_1588, i_1117, i_803);
  and ginst111 (i_1589, i_77, i_1348);
  not ginst112 (i_1590, i_1117);
  and ginst113 (i_1591, i_1117, i_803);
  and ginst114 (i_1592, i_1343, i_1349);
  not ginst115 (i_1593, i_1117);
  and ginst116 (i_1594, i_1117, i_803);
  not ginst117 (i_1595, i_1117);
  and ginst118 (i_1596, i_1117, i_803);
  and ginst119 (i_1597, i_1351, i_870);
  not ginst120 (i_1598, i_1117);
  and ginst121 (i_1599, i_1117, i_803);
  and ginst122 (i_1600, i_116, i_1352);
  and ginst123 (i_1643, i_222, i_1401);
  and ginst124 (i_1644, i_223, i_1402);
  and ginst125 (i_1645, i_226, i_1403);
  and ginst126 (i_1646, i_232, i_1404);
  and ginst127 (i_1647, i_238, i_1405);
  and ginst128 (i_1648, i_244, i_1406);
  and ginst129 (i_1649, i_250, i_1407);
  and ginst130 (i_1650, i_257, i_1408);
  and ginst131 (i_1667, i_1, i_13, i_1426);
  and ginst132 (i_1670, i_1, i_13, i_1427);
  not ginst133 (i_1673, i_1202);
  not ginst134 (i_1674, i_1202);
  not ginst135 (i_1675, i_1202);
  not ginst136 (i_1676, i_1202);
  not ginst137 (i_1677, i_1202);
  not ginst138 (i_1678, i_1202);
  not ginst139 (i_1679, i_1202);
  not ginst140 (i_1680, i_1202);
  nand ginst141 (i_1691, i_1467, i_941);
  nand ginst142 (i_1692, i_1468, i_938);
  nand ginst143 (i_1693, i_1469, i_947);
  nand ginst144 (i_1694, i_1470, i_944);
  not ginst145 (i_1713, i_1505);
  and ginst146 (i_1714, i_87, i_1264);
  nand ginst147 (i_1715, i_1509, i_1510);
  nand ginst148 (i_1718, i_1511, i_1512);
  nand ginst149 (i_1721, i_1507, i_1508);
  and ginst150 (i_1722, i_1340, i_763);
  nand ginst151 (i_1725, i_1340, i_763);
  not ginst152 (i_1726, i_1268);
  nand ginst153 (i_1727, i_1271, i_1493);
  not ginst154 (i_1728, i_1493);
  and ginst155 (i_1729, i_1268, i_683);
  nand ginst156 (i_1730, i_1272, i_1499);
  not ginst157 (i_1731, i_1499);
  nand ginst158 (i_1735, i_87, i_1264);
  not ginst159 (i_1736, i_1273);
  not ginst160 (i_1737, i_1276);
  nand ginst161 (i_1738, i_1325, i_821);
  nand ginst162 (i_1747, i_1325, i_825);
  nand ginst163 (i_1756, i_1279, i_772, i_798);
  nand ginst164 (i_1761, i_1302, i_772, i_786, i_798);
  nand ginst165 (i_1764, i_1339, i_1496);
  not ginst166 (i_1765, i_1496);
  nand ginst167 (i_1766, i_1344, i_1502);
  not ginst168 (i_1767, i_1502);
  not ginst169 (i_1768, i_1328);
  not ginst170 (i_1769, i_1334);
  not ginst171 (i_1770, i_1331);
  and ginst172 (i_1787, i_1579, i_845);
  and ginst173 (i_1788, i_150, i_1580);
  and ginst174 (i_1789, i_1582, i_851);
  and ginst175 (i_1790, i_159, i_1583);
  and ginst176 (i_1791, i_77, i_1584);
  and ginst177 (i_1792, i_50, i_1585);
  and ginst178 (i_1793, i_1587, i_858);
  and ginst179 (i_1794, i_1588, i_845);
  and ginst180 (i_1795, i_1590, i_864);
  and ginst181 (i_1796, i_1591, i_851);
  and ginst182 (i_1797, i_107, i_1593);
  and ginst183 (i_1798, i_77, i_1594);
  and ginst184 (i_1799, i_116, i_1595);
  and ginst185 (i_1800, i_1596, i_858);
  and ginst186 (i_1801, i_283, i_1598);
  and ginst187 (i_1802, i_1599, i_864);
  and ginst188 (i_1803, i_200, i_1363);
  and ginst189 (i_1806, i_1363, i_889);
  and ginst190 (i_1809, i_1366, i_890);
  and ginst191 (i_1812, i_1366, i_891);
  nand ginst192 (i_1815, i_1298, i_1302);
  nand ginst193 (i_1818, i_1302, i_821);
  nand ginst194 (i_1821, i_1179, i_1279, i_772);
  nand ginst195 (i_1824, i_1298, i_786, i_794);
  nand ginst196 (i_1833, i_1298, i_786);
  not ginst197 (i_1842, i_1369);
  not ginst198 (i_1843, i_1369);
  not ginst199 (i_1844, i_1369);
  not ginst200 (i_1845, i_1369);
  not ginst201 (i_1846, i_1369);
  not ginst202 (i_1847, i_1369);
  not ginst203 (i_1848, i_1369);
  not ginst204 (i_1849, i_1384);
  and ginst205 (i_1850, i_1384, i_896);
  not ginst206 (i_1851, i_1384);
  and ginst207 (i_1852, i_1384, i_896);
  not ginst208 (i_1853, i_1384);
  and ginst209 (i_1854, i_1384, i_896);
  not ginst210 (i_1855, i_1384);
  and ginst211 (i_1856, i_1384, i_896);
  not ginst212 (i_1857, i_1384);
  and ginst213 (i_1858, i_1384, i_896);
  not ginst214 (i_1859, i_1384);
  and ginst215 (i_1860, i_1384, i_896);
  not ginst216 (i_1861, i_1384);
  and ginst217 (i_1862, i_1384, i_896);
  not ginst218 (i_1863, i_1384);
  and ginst219 (i_1864, i_1384, i_896);
  and ginst220 (i_1869, i_1202, i_1409);
  nor ginst221 (i_1870, i_50, i_1409);
  not ginst222 (i_1873, i_1306);
  and ginst223 (i_1874, i_1202, i_1409);
  nor ginst224 (i_1875, i_58, i_1409);
  not ginst225 (i_1878, i_1306);
  and ginst226 (i_1879, i_1202, i_1409);
  nor ginst227 (i_1880, i_68, i_1409);
  not ginst228 (i_1883, i_1306);
  and ginst229 (i_1884, i_1202, i_1409);
  nor ginst230 (i_1885, i_77, i_1409);
  not ginst231 (i_1888, i_1306);
  and ginst232 (i_1889, i_1202, i_1409);
  nor ginst233 (i_1890, i_87, i_1409);
  not ginst234 (i_1893, i_1322);
  and ginst235 (i_1894, i_1202, i_1409);
  nor ginst236 (i_1895, i_97, i_1409);
  not ginst237 (i_1898, i_1315);
  and ginst238 (i_1899, i_1202, i_1409);
  nor ginst239 (i_1900, i_107, i_1409);
  not ginst240 (i_1903, i_1315);
  and ginst241 (i_1904, i_1202, i_1409);
  nor ginst242 (i_1905, i_116, i_1409);
  not ginst243 (i_1908, i_1315);
  and ginst244 (i_1909, i_213, i_1452);
  nand ginst245 (i_1912, i_213, i_1452);
  and ginst246 (i_1913, i_213, i_343, i_1452);
  nand ginst247 (i_1917, i_213, i_343, i_1452);
  and ginst248 (i_1922, i_213, i_343, i_1452);
  nand ginst249 (i_1926, i_213, i_343, i_1452);
  not ginst250 (i_1930, i_1464);
  nand ginst251 (i_1933, i_1691, i_1692);
  nand ginst252 (i_1936, i_1693, i_1694);
  not ginst253 (i_1939, i_1471);
  nand ginst254 (i_1940, i_1471, i_1474);
  not ginst255 (i_1941, i_1475);
  not ginst256 (i_1942, i_1478);
  not ginst257 (i_1943, i_1481);
  not ginst258 (i_1944, i_1484);
  not ginst259 (i_1945, i_1487);
  not ginst260 (i_1946, i_1490);
  not ginst261 (i_1947, i_1714);
  nand ginst262 (i_1960, i_1728, i_953);
  nand ginst263 (i_1961, i_1731, i_959);
  and ginst264 (i_1966, i_1276, i_1520);
  nand ginst265 (i_1981, i_1765, i_956);
  nand ginst266 (i_1982, i_1767, i_962);
  and ginst267 (i_1983, i_1067, i_1768);
  or ginst268 (i_1986, i_1581, i_1787, i_1788);
  or ginst269 (i_1987, i_1586, i_1791, i_1792);
  or ginst270 (i_1988, i_1589, i_1793, i_1794);
  or ginst271 (i_1989, i_1592, i_1795, i_1796);
  or ginst272 (i_1990, i_1597, i_1799, i_1800);
  or ginst273 (i_1991, i_1600, i_1801, i_1802);
  and ginst274 (i_2022, i_77, i_1849);
  and ginst275 (i_2023, i_223, i_1850);
  and ginst276 (i_2024, i_87, i_1851);
  and ginst277 (i_2025, i_226, i_1852);
  and ginst278 (i_2026, i_97, i_1853);
  and ginst279 (i_2027, i_232, i_1854);
  and ginst280 (i_2028, i_107, i_1855);
  and ginst281 (i_2029, i_238, i_1856);
  and ginst282 (i_2030, i_116, i_1857);
  and ginst283 (i_2031, i_244, i_1858);
  and ginst284 (i_2032, i_283, i_1859);
  and ginst285 (i_2033, i_250, i_1860);
  and ginst286 (i_2034, i_294, i_1861);
  and ginst287 (i_2035, i_257, i_1862);
  and ginst288 (i_2036, i_303, i_1863);
  and ginst289 (i_2037, i_264, i_1864);
  not ginst290 (i_2038, i_1667);
  not ginst291 (i_2043, i_1667);
  not ginst292 (i_2052, i_1670);
  not ginst293 (i_2057, i_1670);
  and ginst294 (i_2068, i_50, i_1197, i_1869);
  and ginst295 (i_2073, i_58, i_1197, i_1874);
  and ginst296 (i_2078, i_68, i_1197, i_1879);
  and ginst297 (i_2083, i_77, i_1197, i_1884);
  and ginst298 (i_2088, i_87, i_1219, i_1889);
  and ginst299 (i_2093, i_97, i_1219, i_1894);
  and ginst300 (i_2098, i_107, i_1219, i_1899);
  and ginst301 (i_2103, i_116, i_1219, i_1904);
  not ginst302 (i_2121, i_1562);
  not ginst303 (i_2122, i_1562);
  not ginst304 (i_2123, i_1562);
  not ginst305 (i_2124, i_1562);
  not ginst306 (i_2125, i_1562);
  not ginst307 (i_2126, i_1562);
  not ginst308 (i_2127, i_1562);
  not ginst309 (i_2128, i_1562);
  nand ginst310 (i_2133, i_1939, i_950);
  nand ginst311 (i_2134, i_1478, i_1941);
  nand ginst312 (i_2135, i_1475, i_1942);
  nand ginst313 (i_2136, i_1484, i_1943);
  nand ginst314 (i_2137, i_1481, i_1944);
  nand ginst315 (i_2138, i_1490, i_1945);
  nand ginst316 (i_2139, i_1487, i_1946);
  not ginst317 (i_2141, i_1933);
  not ginst318 (i_2142, i_1936);
  not ginst319 (i_2143, i_1738);
  and ginst320 (i_2144, i_1738, i_1747);
  not ginst321 (i_2145, i_1747);
  nand ginst322 (i_2146, i_1727, i_1960);
  nand ginst323 (i_2147, i_1730, i_1961);
  and ginst324 (i_2148, i_58, i_1267, i_1722, i_665);
  not ginst325 (i_2149, i_1738);
  and ginst326 (i_2150, i_1738, i_1747);
  not ginst327 (i_2151, i_1747);
  not ginst328 (i_2152, i_1738);
  not ginst329 (i_2153, i_1747);
  and ginst330 (i_2154, i_1738, i_1747);
  not ginst331 (i_2155, i_1738);
  not ginst332 (i_2156, i_1747);
  and ginst333 (i_2157, i_1738, i_1747);
  not ginst334 (i_2158, i_1761);
  not ginst335 (i_2175, i_1761);
  nand ginst336 (i_2178, i_1764, i_1981);
  nand ginst337 (i_2179, i_1766, i_1982);
  not ginst338 (i_2180, i_1756);
  and ginst339 (i_2181, i_1328, i_1756);
  not ginst340 (i_2183, i_1756);
  and ginst341 (i_2184, i_1331, i_1756);
  nand ginst342 (i_2185, i_1358, i_1812);
  nand ginst343 (i_2188, i_1358, i_1809);
  nand ginst344 (i_2191, i_1353, i_1812);
  nand ginst345 (i_2194, i_1353, i_1809);
  nand ginst346 (i_2197, i_1358, i_1806);
  nand ginst347 (i_2200, i_1358, i_1803);
  nand ginst348 (i_2203, i_1353, i_1806);
  nand ginst349 (i_2206, i_1353, i_1803);
  not ginst350 (i_2209, i_1815);
  not ginst351 (i_2210, i_1818);
  and ginst352 (i_2211, i_1815, i_1818);
  not ginst353 (i_2212, i_1821);
  not ginst354 (i_2221, i_1821);
  not ginst355 (i_2230, i_1833);
  not ginst356 (i_2231, i_1833);
  not ginst357 (i_2232, i_1833);
  not ginst358 (i_2233, i_1833);
  not ginst359 (i_2234, i_1824);
  not ginst360 (i_2235, i_1824);
  not ginst361 (i_2236, i_1824);
  not ginst362 (i_2237, i_1824);
  or ginst363 (i_2238, i_1643, i_2022, i_2023);
  or ginst364 (i_2239, i_1644, i_2024, i_2025);
  or ginst365 (i_2240, i_1645, i_2026, i_2027);
  or ginst366 (i_2241, i_1646, i_2028, i_2029);
  or ginst367 (i_2242, i_1647, i_2030, i_2031);
  or ginst368 (i_2243, i_1648, i_2032, i_2033);
  or ginst369 (i_2244, i_1649, i_2034, i_2035);
  or ginst370 (i_2245, i_1650, i_2036, i_2037);
  and ginst371 (i_2270, i_1673, i_1986);
  and ginst372 (i_2277, i_1675, i_1987);
  and ginst373 (i_2282, i_1676, i_1988);
  and ginst374 (i_2287, i_1677, i_1989);
  and ginst375 (i_2294, i_1679, i_1990);
  and ginst376 (i_2299, i_1680, i_1991);
  not ginst377 (i_2304, i_1917);
  and ginst378 (i_2307, i_350, i_1930);
  nand ginst379 (i_2310, i_350, i_1930);
  not ginst380 (i_2313, i_1715);
  not ginst381 (i_2316, i_1718);
  not ginst382 (i_2319, i_1715);
  not ginst383 (i_2322, i_1718);
  nand ginst384 (i_2325, i_1940, i_2133);
  nand ginst385 (i_2328, i_2134, i_2135);
  nand ginst386 (i_2331, i_2136, i_2137);
  nand ginst387 (i_2334, i_2138, i_2139);
  nand ginst388 (i_2341, i_1936, i_2141);
  nand ginst389 (i_2342, i_1933, i_2142);
  and ginst390 (i_2347, i_2144, i_724);
  and ginst391 (i_2348, i_1726, i_2146, i_699);
  and ginst392 (i_2349, i_2147, i_753);
  and ginst393 (i_2350, i_1273, i_2148);
  and ginst394 (i_2351, i_2150, i_736);
  and ginst395 (i_2352, i_1735, i_2153);
  and ginst396 (i_2353, i_2154, i_763);
  and ginst397 (i_2354, i_1725, i_2156);
  and ginst398 (i_2355, i_2157, i_749);
  not ginst399 (i_2374, i_2178);
  not ginst400 (i_2375, i_2179);
  and ginst401 (i_2376, i_1520, i_2180);
  and ginst402 (i_2379, i_1721, i_2181);
  and ginst403 (i_2398, i_2211, i_665);
  and ginst404 (i_2417, i_226, i_1873, i_2057);
  and ginst405 (i_2418, i_274, i_1306, i_2057);
  and ginst406 (i_2419, i_2052, i_2238);
  and ginst407 (i_2420, i_232, i_1878, i_2057);
  and ginst408 (i_2421, i_274, i_1306, i_2057);
  and ginst409 (i_2422, i_2052, i_2239);
  and ginst410 (i_2425, i_238, i_1883, i_2057);
  and ginst411 (i_2426, i_274, i_1306, i_2057);
  and ginst412 (i_2427, i_2052, i_2240);
  and ginst413 (i_2430, i_244, i_1888, i_2057);
  and ginst414 (i_2431, i_274, i_1306, i_2057);
  and ginst415 (i_2432, i_2052, i_2241);
  and ginst416 (i_2435, i_250, i_1893, i_2043);
  and ginst417 (i_2436, i_274, i_1322, i_2043);
  and ginst418 (i_2437, i_2038, i_2242);
  and ginst419 (i_2438, i_257, i_1898, i_2043);
  and ginst420 (i_2439, i_274, i_1315, i_2043);
  and ginst421 (i_2440, i_2038, i_2243);
  and ginst422 (i_2443, i_264, i_1903, i_2043);
  and ginst423 (i_2444, i_274, i_1315, i_2043);
  and ginst424 (i_2445, i_2038, i_2244);
  and ginst425 (i_2448, i_270, i_1908, i_2043);
  and ginst426 (i_2449, i_274, i_1315, i_2043);
  and ginst427 (i_2450, i_2038, i_2245);
  not ginst428 (i_2467, i_2313);
  not ginst429 (i_2468, i_2316);
  not ginst430 (i_2469, i_2319);
  not ginst431 (i_2470, i_2322);
  nand ginst432 (i_2471, i_2341, i_2342);
  not ginst433 (i_2474, i_2325);
  not ginst434 (i_2475, i_2328);
  not ginst435 (i_2476, i_2331);
  not ginst436 (i_2477, i_2334);
  or ginst437 (i_2478, i_1729, i_2348);
  not ginst438 (i_2481, i_2175);
  and ginst439 (i_2482, i_1334, i_2175);
  and ginst440 (i_2483, i_2183, i_2349);
  and ginst441 (i_2486, i_1346, i_2374);
  and ginst442 (i_2487, i_1350, i_2375);
  not ginst443 (i_2488, i_2185);
  not ginst444 (i_2497, i_2188);
  not ginst445 (i_2506, i_2191);
  not ginst446 (i_2515, i_2194);
  not ginst447 (i_2524, i_2197);
  not ginst448 (i_2533, i_2200);
  not ginst449 (i_2542, i_2203);
  not ginst450 (i_2551, i_2206);
  not ginst451 (i_2560, i_2185);
  not ginst452 (i_2569, i_2188);
  not ginst453 (i_2578, i_2191);
  not ginst454 (i_2587, i_2194);
  not ginst455 (i_2596, i_2197);
  not ginst456 (i_2605, i_2200);
  not ginst457 (i_2614, i_2203);
  not ginst458 (i_2623, i_2206);
  not ginst459 (i_2632, i_2212);
  and ginst460 (i_2633, i_1833, i_2212);
  not ginst461 (i_2634, i_2212);
  and ginst462 (i_2635, i_1833, i_2212);
  not ginst463 (i_2636, i_2212);
  and ginst464 (i_2637, i_1833, i_2212);
  not ginst465 (i_2638, i_2212);
  and ginst466 (i_2639, i_1833, i_2212);
  not ginst467 (i_2640, i_2221);
  and ginst468 (i_2641, i_1824, i_2221);
  not ginst469 (i_2642, i_2221);
  and ginst470 (i_2643, i_1824, i_2221);
  not ginst471 (i_2644, i_2221);
  and ginst472 (i_2645, i_1824, i_2221);
  not ginst473 (i_2646, i_2221);
  and ginst474 (i_2647, i_1824, i_2221);
  or ginst475 (i_2648, i_1870, i_2068, i_2270);
  nor ginst476 (i_2652, i_1870, i_2068, i_2270);
  or ginst477 (i_2656, i_2417, i_2418, i_2419);
  or ginst478 (i_2659, i_2420, i_2421, i_2422);
  or ginst479 (i_2662, i_1880, i_2078, i_2277);
  nor ginst480 (i_2666, i_1880, i_2078, i_2277);
  or ginst481 (i_2670, i_2425, i_2426, i_2427);
  or ginst482 (i_2673, i_1885, i_2083, i_2282);
  nor ginst483 (i_2677, i_1885, i_2083, i_2282);
  or ginst484 (i_2681, i_2430, i_2431, i_2432);
  or ginst485 (i_2684, i_1890, i_2088, i_2287);
  nor ginst486 (i_2688, i_1890, i_2088, i_2287);
  or ginst487 (i_2692, i_2435, i_2436, i_2437);
  or ginst488 (i_2697, i_2438, i_2439, i_2440);
  or ginst489 (i_2702, i_1900, i_2098, i_2294);
  nor ginst490 (i_2706, i_1900, i_2098, i_2294);
  or ginst491 (i_2710, i_2443, i_2444, i_2445);
  or ginst492 (i_2715, i_1905, i_2103, i_2299);
  nor ginst493 (i_2719, i_1905, i_2103, i_2299);
  or ginst494 (i_2723, i_2448, i_2449, i_2450);
  not ginst495 (i_2728, i_2304);
  not ginst496 (i_2729, i_2158);
  and ginst497 (i_2730, i_1562, i_2158);
  not ginst498 (i_2731, i_2158);
  and ginst499 (i_2732, i_1562, i_2158);
  not ginst500 (i_2733, i_2158);
  and ginst501 (i_2734, i_1562, i_2158);
  not ginst502 (i_2735, i_2158);
  and ginst503 (i_2736, i_1562, i_2158);
  not ginst504 (i_2737, i_2158);
  and ginst505 (i_2738, i_1562, i_2158);
  not ginst506 (i_2739, i_2158);
  and ginst507 (i_2740, i_1562, i_2158);
  not ginst508 (i_2741, i_2158);
  and ginst509 (i_2742, i_1562, i_2158);
  not ginst510 (i_2743, i_2158);
  and ginst511 (i_2744, i_1562, i_2158);
  or ginst512 (i_2745, i_1983, i_2376, i_2379);
  nor ginst513 (i_2746, i_1983, i_2376, i_2379);
  nand ginst514 (i_2748, i_2316, i_2467);
  nand ginst515 (i_2749, i_2313, i_2468);
  nand ginst516 (i_2750, i_2322, i_2469);
  nand ginst517 (i_2751, i_2319, i_2470);
  nand ginst518 (i_2754, i_2328, i_2474);
  nand ginst519 (i_2755, i_2325, i_2475);
  nand ginst520 (i_2756, i_2334, i_2476);
  nand ginst521 (i_2757, i_2331, i_2477);
  and ginst522 (i_2758, i_1520, i_2481);
  and ginst523 (i_2761, i_1722, i_2482);
  and ginst524 (i_2764, i_1770, i_2478);
  or ginst525 (i_2768, i_1789, i_1790, i_2486);
  or ginst526 (i_2769, i_1797, i_1798, i_2487);
  and ginst527 (i_2898, i_2633, i_665);
  and ginst528 (i_2899, i_2635, i_679);
  and ginst529 (i_2900, i_2637, i_686);
  and ginst530 (i_2901, i_2639, i_702);
  not ginst531 (i_2962, i_2746);
  nand ginst532 (i_2966, i_2748, i_2749);
  nand ginst533 (i_2967, i_2750, i_2751);
  not ginst534 (i_2970, i_2471);
  nand ginst535 (i_2973, i_2754, i_2755);
  nand ginst536 (i_2977, i_2756, i_2757);
  and ginst537 (i_2980, i_2143, i_2471);
  not ginst538 (i_2984, i_2488);
  not ginst539 (i_2985, i_2497);
  not ginst540 (i_2986, i_2506);
  not ginst541 (i_2987, i_2515);
  not ginst542 (i_2988, i_2524);
  not ginst543 (i_2989, i_2533);
  not ginst544 (i_2990, i_2542);
  not ginst545 (i_2991, i_2551);
  not ginst546 (i_2992, i_2488);
  not ginst547 (i_2993, i_2497);
  not ginst548 (i_2994, i_2506);
  not ginst549 (i_2995, i_2515);
  not ginst550 (i_2996, i_2524);
  not ginst551 (i_2997, i_2533);
  not ginst552 (i_2998, i_2542);
  not ginst553 (i_2999, i_2551);
  not ginst554 (i_3000, i_2488);
  not ginst555 (i_3001, i_2497);
  not ginst556 (i_3002, i_2506);
  not ginst557 (i_3003, i_2515);
  not ginst558 (i_3004, i_2524);
  not ginst559 (i_3005, i_2533);
  not ginst560 (i_3006, i_2542);
  not ginst561 (i_3007, i_2551);
  not ginst562 (i_3008, i_2488);
  not ginst563 (i_3009, i_2497);
  not ginst564 (i_3010, i_2506);
  not ginst565 (i_3011, i_2515);
  not ginst566 (i_3012, i_2524);
  not ginst567 (i_3013, i_2533);
  not ginst568 (i_3014, i_2542);
  not ginst569 (i_3015, i_2551);
  not ginst570 (i_3016, i_2488);
  not ginst571 (i_3017, i_2497);
  not ginst572 (i_3018, i_2506);
  not ginst573 (i_3019, i_2515);
  not ginst574 (i_3020, i_2524);
  not ginst575 (i_3021, i_2533);
  not ginst576 (i_3022, i_2542);
  not ginst577 (i_3023, i_2551);
  not ginst578 (i_3024, i_2488);
  not ginst579 (i_3025, i_2497);
  not ginst580 (i_3026, i_2506);
  not ginst581 (i_3027, i_2515);
  not ginst582 (i_3028, i_2524);
  not ginst583 (i_3029, i_2533);
  not ginst584 (i_3030, i_2542);
  not ginst585 (i_3031, i_2551);
  not ginst586 (i_3032, i_2488);
  not ginst587 (i_3033, i_2497);
  not ginst588 (i_3034, i_2506);
  not ginst589 (i_3035, i_2515);
  not ginst590 (i_3036, i_2524);
  not ginst591 (i_3037, i_2533);
  not ginst592 (i_3038, i_2542);
  not ginst593 (i_3039, i_2551);
  not ginst594 (i_3040, i_2488);
  not ginst595 (i_3041, i_2497);
  not ginst596 (i_3042, i_2506);
  not ginst597 (i_3043, i_2515);
  not ginst598 (i_3044, i_2524);
  not ginst599 (i_3045, i_2533);
  not ginst600 (i_3046, i_2542);
  not ginst601 (i_3047, i_2551);
  not ginst602 (i_3048, i_2560);
  not ginst603 (i_3049, i_2569);
  not ginst604 (i_3050, i_2578);
  not ginst605 (i_3051, i_2587);
  not ginst606 (i_3052, i_2596);
  not ginst607 (i_3053, i_2605);
  not ginst608 (i_3054, i_2614);
  not ginst609 (i_3055, i_2623);
  not ginst610 (i_3056, i_2560);
  not ginst611 (i_3057, i_2569);
  not ginst612 (i_3058, i_2578);
  not ginst613 (i_3059, i_2587);
  not ginst614 (i_3060, i_2596);
  not ginst615 (i_3061, i_2605);
  not ginst616 (i_3062, i_2614);
  not ginst617 (i_3063, i_2623);
  not ginst618 (i_3064, i_2560);
  not ginst619 (i_3065, i_2569);
  not ginst620 (i_3066, i_2578);
  not ginst621 (i_3067, i_2587);
  not ginst622 (i_3068, i_2596);
  not ginst623 (i_3069, i_2605);
  not ginst624 (i_3070, i_2614);
  not ginst625 (i_3071, i_2623);
  not ginst626 (i_3072, i_2560);
  not ginst627 (i_3073, i_2569);
  not ginst628 (i_3074, i_2578);
  not ginst629 (i_3075, i_2587);
  not ginst630 (i_3076, i_2596);
  not ginst631 (i_3077, i_2605);
  not ginst632 (i_3078, i_2614);
  not ginst633 (i_3079, i_2623);
  not ginst634 (i_3080, i_2560);
  not ginst635 (i_3081, i_2569);
  not ginst636 (i_3082, i_2578);
  not ginst637 (i_3083, i_2587);
  not ginst638 (i_3084, i_2596);
  not ginst639 (i_3085, i_2605);
  not ginst640 (i_3086, i_2614);
  not ginst641 (i_3087, i_2623);
  not ginst642 (i_3088, i_2560);
  not ginst643 (i_3089, i_2569);
  not ginst644 (i_3090, i_2578);
  not ginst645 (i_3091, i_2587);
  not ginst646 (i_3092, i_2596);
  not ginst647 (i_3093, i_2605);
  not ginst648 (i_3094, i_2614);
  not ginst649 (i_3095, i_2623);
  not ginst650 (i_3096, i_2560);
  not ginst651 (i_3097, i_2569);
  not ginst652 (i_3098, i_2578);
  not ginst653 (i_3099, i_2587);
  not ginst654 (i_3100, i_2596);
  not ginst655 (i_3101, i_2605);
  not ginst656 (i_3102, i_2614);
  not ginst657 (i_3103, i_2623);
  not ginst658 (i_3104, i_2560);
  not ginst659 (i_3105, i_2569);
  not ginst660 (i_3106, i_2578);
  not ginst661 (i_3107, i_2587);
  not ginst662 (i_3108, i_2596);
  not ginst663 (i_3109, i_2605);
  not ginst664 (i_3110, i_2614);
  not ginst665 (i_3111, i_2623);
  not ginst666 (i_3112, i_2656);
  not ginst667 (i_3115, i_2656);
  not ginst668 (i_3118, i_2652);
  and ginst669 (i_3119, i_1674, i_2768);
  not ginst670 (i_3122, i_2659);
  not ginst671 (i_3125, i_2659);
  not ginst672 (i_3128, i_2670);
  not ginst673 (i_3131, i_2670);
  not ginst674 (i_3134, i_2666);
  not ginst675 (i_3135, i_2681);
  not ginst676 (i_3138, i_2681);
  not ginst677 (i_3141, i_2677);
  not ginst678 (i_3142, i_2692);
  not ginst679 (i_3145, i_2692);
  not ginst680 (i_3148, i_2688);
  and ginst681 (i_3149, i_1678, i_2769);
  not ginst682 (i_3152, i_2697);
  not ginst683 (i_3155, i_2697);
  not ginst684 (i_3158, i_2710);
  not ginst685 (i_3161, i_2710);
  not ginst686 (i_3164, i_2706);
  not ginst687 (i_3165, i_2723);
  not ginst688 (i_3168, i_2723);
  not ginst689 (i_3171, i_2719);
  and ginst690 (i_3172, i_1909, i_2648);
  and ginst691 (i_3175, i_1913, i_2662);
  and ginst692 (i_3178, i_1913, i_2673);
  and ginst693 (i_3181, i_1913, i_2684);
  and ginst694 (i_3184, i_1922, i_2702);
  and ginst695 (i_3187, i_1922, i_2715);
  not ginst696 (i_3190, i_2692);
  not ginst697 (i_3191, i_2697);
  not ginst698 (i_3192, i_2710);
  not ginst699 (i_3193, i_2723);
  and ginst700 (i_3194, i_1459, i_2692, i_2697, i_2710, i_2723);
  nand ginst701 (i_3195, i_2745, i_2962);
  not ginst702 (i_3196, i_2966);
  or ginst703 (i_3206, i_2145, i_2347, i_2980);
  and ginst704 (i_3207, i_124, i_2984);
  and ginst705 (i_3208, i_159, i_2985);
  and ginst706 (i_3209, i_150, i_2986);
  and ginst707 (i_3210, i_143, i_2987);
  and ginst708 (i_3211, i_137, i_2988);
  and ginst709 (i_3212, i_132, i_2989);
  and ginst710 (i_3213, i_128, i_2990);
  and ginst711 (i_3214, i_125, i_2991);
  and ginst712 (i_3215, i_125, i_2992);
  and ginst713 (i_3216, i_2993, i_655);
  and ginst714 (i_3217, i_159, i_2994);
  and ginst715 (i_3218, i_150, i_2995);
  and ginst716 (i_3219, i_143, i_2996);
  and ginst717 (i_3220, i_137, i_2997);
  and ginst718 (i_3221, i_132, i_2998);
  and ginst719 (i_3222, i_128, i_2999);
  and ginst720 (i_3223, i_128, i_3000);
  and ginst721 (i_3224, i_3001, i_670);
  and ginst722 (i_3225, i_3002, i_655);
  and ginst723 (i_3226, i_159, i_3003);
  and ginst724 (i_3227, i_150, i_3004);
  and ginst725 (i_3228, i_143, i_3005);
  and ginst726 (i_3229, i_137, i_3006);
  and ginst727 (i_3230, i_132, i_3007);
  and ginst728 (i_3231, i_132, i_3008);
  and ginst729 (i_3232, i_3009, i_690);
  and ginst730 (i_3233, i_3010, i_670);
  and ginst731 (i_3234, i_3011, i_655);
  and ginst732 (i_3235, i_159, i_3012);
  and ginst733 (i_3236, i_150, i_3013);
  and ginst734 (i_3237, i_143, i_3014);
  and ginst735 (i_3238, i_137, i_3015);
  and ginst736 (i_3239, i_137, i_3016);
  and ginst737 (i_3240, i_3017, i_706);
  and ginst738 (i_3241, i_3018, i_690);
  and ginst739 (i_3242, i_3019, i_670);
  and ginst740 (i_3243, i_3020, i_655);
  and ginst741 (i_3244, i_159, i_3021);
  and ginst742 (i_3245, i_150, i_3022);
  and ginst743 (i_3246, i_143, i_3023);
  and ginst744 (i_3247, i_143, i_3024);
  and ginst745 (i_3248, i_3025, i_715);
  and ginst746 (i_3249, i_3026, i_706);
  and ginst747 (i_3250, i_3027, i_690);
  and ginst748 (i_3251, i_3028, i_670);
  and ginst749 (i_3252, i_3029, i_655);
  and ginst750 (i_3253, i_159, i_3030);
  and ginst751 (i_3254, i_150, i_3031);
  and ginst752 (i_3255, i_150, i_3032);
  and ginst753 (i_3256, i_3033, i_727);
  and ginst754 (i_3257, i_3034, i_715);
  and ginst755 (i_3258, i_3035, i_706);
  and ginst756 (i_3259, i_3036, i_690);
  and ginst757 (i_3260, i_3037, i_670);
  and ginst758 (i_3261, i_3038, i_655);
  and ginst759 (i_3262, i_159, i_3039);
  and ginst760 (i_3263, i_159, i_3040);
  and ginst761 (i_3264, i_3041, i_740);
  and ginst762 (i_3265, i_3042, i_727);
  and ginst763 (i_3266, i_3043, i_715);
  and ginst764 (i_3267, i_3044, i_706);
  and ginst765 (i_3268, i_3045, i_690);
  and ginst766 (i_3269, i_3046, i_670);
  and ginst767 (i_3270, i_3047, i_655);
  and ginst768 (i_3271, i_283, i_3048);
  and ginst769 (i_3272, i_3049, i_670);
  and ginst770 (i_3273, i_3050, i_690);
  and ginst771 (i_3274, i_3051, i_706);
  and ginst772 (i_3275, i_3052, i_715);
  and ginst773 (i_3276, i_3053, i_727);
  and ginst774 (i_3277, i_3054, i_740);
  and ginst775 (i_3278, i_3055, i_753);
  and ginst776 (i_3279, i_294, i_3056);
  and ginst777 (i_3280, i_3057, i_690);
  and ginst778 (i_3281, i_3058, i_706);
  and ginst779 (i_3282, i_3059, i_715);
  and ginst780 (i_3283, i_3060, i_727);
  and ginst781 (i_3284, i_3061, i_740);
  and ginst782 (i_3285, i_3062, i_753);
  and ginst783 (i_3286, i_283, i_3063);
  and ginst784 (i_3287, i_303, i_3064);
  and ginst785 (i_3288, i_3065, i_706);
  and ginst786 (i_3289, i_3066, i_715);
  and ginst787 (i_3290, i_3067, i_727);
  and ginst788 (i_3291, i_3068, i_740);
  and ginst789 (i_3292, i_3069, i_753);
  and ginst790 (i_3293, i_283, i_3070);
  and ginst791 (i_3294, i_294, i_3071);
  and ginst792 (i_3295, i_311, i_3072);
  and ginst793 (i_3296, i_3073, i_715);
  and ginst794 (i_3297, i_3074, i_727);
  and ginst795 (i_3298, i_3075, i_740);
  and ginst796 (i_3299, i_3076, i_753);
  and ginst797 (i_3300, i_283, i_3077);
  and ginst798 (i_3301, i_294, i_3078);
  and ginst799 (i_3302, i_303, i_3079);
  and ginst800 (i_3303, i_317, i_3080);
  and ginst801 (i_3304, i_3081, i_727);
  and ginst802 (i_3305, i_3082, i_740);
  and ginst803 (i_3306, i_3083, i_753);
  and ginst804 (i_3307, i_283, i_3084);
  and ginst805 (i_3308, i_294, i_3085);
  and ginst806 (i_3309, i_303, i_3086);
  and ginst807 (i_3310, i_311, i_3087);
  and ginst808 (i_3311, i_322, i_3088);
  and ginst809 (i_3312, i_3089, i_740);
  and ginst810 (i_3313, i_3090, i_753);
  and ginst811 (i_3314, i_283, i_3091);
  and ginst812 (i_3315, i_294, i_3092);
  and ginst813 (i_3316, i_303, i_3093);
  and ginst814 (i_3317, i_311, i_3094);
  and ginst815 (i_3318, i_317, i_3095);
  and ginst816 (i_3319, i_326, i_3096);
  and ginst817 (i_3320, i_3097, i_753);
  and ginst818 (i_3321, i_283, i_3098);
  and ginst819 (i_3322, i_294, i_3099);
  and ginst820 (i_3323, i_303, i_3100);
  and ginst821 (i_3324, i_311, i_3101);
  and ginst822 (i_3325, i_317, i_3102);
  and ginst823 (i_3326, i_322, i_3103);
  and ginst824 (i_3327, i_329, i_3104);
  and ginst825 (i_3328, i_283, i_3105);
  and ginst826 (i_3329, i_294, i_3106);
  and ginst827 (i_3330, i_303, i_3107);
  and ginst828 (i_3331, i_311, i_3108);
  and ginst829 (i_3332, i_317, i_3109);
  and ginst830 (i_3333, i_322, i_3110);
  and ginst831 (i_3334, i_326, i_3111);
  and ginst832 (i_3383, i_3190, i_3191, i_3192, i_3193, i_917);
  not ginst833 (i_3384, i_2977);
  and ginst834 (i_3387, i_1736, i_3196);
  and ginst835 (i_3388, i_2149, i_2977);
  and ginst836 (i_3389, i_1737, i_2973);
  nor ginst837 (i_3390, i_3207, i_3208, i_3209, i_3210, i_3211, i_3212, i_3213, i_3214);
  nor ginst838 (i_3391, i_3215, i_3216, i_3217, i_3218, i_3219, i_3220, i_3221, i_3222);
  nor ginst839 (i_3392, i_3223, i_3224, i_3225, i_3226, i_3227, i_3228, i_3229, i_3230);
  nor ginst840 (i_3393, i_3231, i_3232, i_3233, i_3234, i_3235, i_3236, i_3237, i_3238);
  nor ginst841 (i_3394, i_3239, i_3240, i_3241, i_3242, i_3243, i_3244, i_3245, i_3246);
  nor ginst842 (i_3395, i_3247, i_3248, i_3249, i_3250, i_3251, i_3252, i_3253, i_3254);
  nor ginst843 (i_3396, i_3255, i_3256, i_3257, i_3258, i_3259, i_3260, i_3261, i_3262);
  nor ginst844 (i_3397, i_3263, i_3264, i_3265, i_3266, i_3267, i_3268, i_3269, i_3270);
  nor ginst845 (i_3398, i_3271, i_3272, i_3273, i_3274, i_3275, i_3276, i_3277, i_3278);
  nor ginst846 (i_3399, i_3279, i_3280, i_3281, i_3282, i_3283, i_3284, i_3285, i_3286);
  nor ginst847 (i_3400, i_3287, i_3288, i_3289, i_3290, i_3291, i_3292, i_3293, i_3294);
  nor ginst848 (i_3401, i_3295, i_3296, i_3297, i_3298, i_3299, i_3300, i_3301, i_3302);
  nor ginst849 (i_3402, i_3303, i_3304, i_3305, i_3306, i_3307, i_3308, i_3309, i_3310);
  nor ginst850 (i_3403, i_3311, i_3312, i_3313, i_3314, i_3315, i_3316, i_3317, i_3318);
  nor ginst851 (i_3404, i_3319, i_3320, i_3321, i_3322, i_3323, i_3324, i_3325, i_3326);
  nor ginst852 (i_3405, i_3327, i_3328, i_3329, i_3330, i_3331, i_3332, i_3333, i_3334);
  and ginst853 (i_3406, i_2641, i_3206);
  and ginst854 (i_3407, i_169, i_2648, i_3112);
  and ginst855 (i_3410, i_179, i_2648, i_3115);
  and ginst856 (i_3413, i_190, i_2652, i_3115);
  and ginst857 (i_3414, i_200, i_2652, i_3112);
  or ginst858 (i_3415, i_1875, i_2073, i_3119);
  nor ginst859 (i_3419, i_1875, i_2073, i_3119);
  and ginst860 (i_3423, i_169, i_2662, i_3128);
  and ginst861 (i_3426, i_179, i_2662, i_3131);
  and ginst862 (i_3429, i_190, i_2666, i_3131);
  and ginst863 (i_3430, i_200, i_2666, i_3128);
  and ginst864 (i_3431, i_169, i_2673, i_3135);
  and ginst865 (i_3434, i_179, i_2673, i_3138);
  and ginst866 (i_3437, i_190, i_2677, i_3138);
  and ginst867 (i_3438, i_200, i_2677, i_3135);
  and ginst868 (i_3439, i_169, i_2684, i_3142);
  and ginst869 (i_3442, i_179, i_2684, i_3145);
  and ginst870 (i_3445, i_190, i_2688, i_3145);
  and ginst871 (i_3446, i_200, i_2688, i_3142);
  or ginst872 (i_3447, i_1895, i_2093, i_3149);
  nor ginst873 (i_3451, i_1895, i_2093, i_3149);
  and ginst874 (i_3455, i_169, i_2702, i_3158);
  and ginst875 (i_3458, i_179, i_2702, i_3161);
  and ginst876 (i_3461, i_190, i_2706, i_3161);
  and ginst877 (i_3462, i_200, i_2706, i_3158);
  and ginst878 (i_3463, i_169, i_2715, i_3165);
  and ginst879 (i_3466, i_179, i_2715, i_3168);
  and ginst880 (i_3469, i_190, i_2719, i_3168);
  and ginst881 (i_3470, i_200, i_2719, i_3165);
  or ginst882 (i_3471, i_3194, i_3383);
  not ginst883 (i_3472, i_2967);
  not ginst884 (i_3475, i_2970);
  not ginst885 (i_3478, i_2967);
  not ginst886 (i_3481, i_2970);
  not ginst887 (i_3484, i_2973);
  not ginst888 (i_3487, i_2973);
  not ginst889 (i_3490, i_3172);
  not ginst890 (i_3493, i_3172);
  not ginst891 (i_3496, i_3175);
  not ginst892 (i_3499, i_3175);
  not ginst893 (i_3502, i_3178);
  not ginst894 (i_3505, i_3178);
  not ginst895 (i_3508, i_3181);
  not ginst896 (i_3511, i_3181);
  not ginst897 (i_3514, i_3184);
  not ginst898 (i_3517, i_3184);
  not ginst899 (i_3520, i_3187);
  not ginst900 (i_3523, i_3187);
  nor ginst901 (i_3534, i_2350, i_3387);
  or ginst902 (i_3535, i_2151, i_2351, i_3388);
  nor ginst903 (i_3536, i_1966, i_3389);
  and ginst904 (i_3537, i_2209, i_3390);
  and ginst905 (i_3538, i_2210, i_3398);
  and ginst906 (i_3539, i_1842, i_3391);
  and ginst907 (i_3540, i_1369, i_3399);
  and ginst908 (i_3541, i_1843, i_3392);
  and ginst909 (i_3542, i_1369, i_3400);
  and ginst910 (i_3543, i_1844, i_3393);
  and ginst911 (i_3544, i_1369, i_3401);
  and ginst912 (i_3545, i_1845, i_3394);
  and ginst913 (i_3546, i_1369, i_3402);
  and ginst914 (i_3547, i_1846, i_3395);
  and ginst915 (i_3548, i_1369, i_3403);
  and ginst916 (i_3549, i_1847, i_3396);
  and ginst917 (i_3550, i_1369, i_3404);
  and ginst918 (i_3551, i_1848, i_3397);
  and ginst919 (i_3552, i_1369, i_3405);
  or ginst920 (i_3557, i_3118, i_3413, i_3414);
  or ginst921 (i_3568, i_3134, i_3429, i_3430);
  or ginst922 (i_3573, i_3141, i_3437, i_3438);
  or ginst923 (i_3578, i_3148, i_3445, i_3446);
  or ginst924 (i_3589, i_3164, i_3461, i_3462);
  or ginst925 (i_3594, i_3171, i_3469, i_3470);
  and ginst926 (i_3605, i_2728, i_3471);
  not ginst927 (i_3626, i_3478);
  not ginst928 (i_3627, i_3481);
  not ginst929 (i_3628, i_3487);
  not ginst930 (i_3629, i_3484);
  not ginst931 (i_3630, i_3472);
  not ginst932 (i_3631, i_3475);
  and ginst933 (i_3632, i_2152, i_3536);
  and ginst934 (i_3633, i_2155, i_3534);
  or ginst935 (i_3634, i_2398, i_3537, i_3538);
  or ginst936 (i_3635, i_3539, i_3540);
  or ginst937 (i_3636, i_3541, i_3542);
  or ginst938 (i_3637, i_3543, i_3544);
  or ginst939 (i_3638, i_3545, i_3546);
  or ginst940 (i_3639, i_3547, i_3548);
  or ginst941 (i_3640, i_3549, i_3550);
  or ginst942 (i_3641, i_3551, i_3552);
  and ginst943 (i_3642, i_2643, i_3535);
  or ginst944 (i_3643, i_3407, i_3410);
  nor ginst945 (i_3644, i_3407, i_3410);
  and ginst946 (i_3645, i_169, i_3122, i_3415);
  and ginst947 (i_3648, i_179, i_3125, i_3415);
  and ginst948 (i_3651, i_190, i_3125, i_3419);
  and ginst949 (i_3652, i_200, i_3122, i_3419);
  not ginst950 (i_3653, i_3419);
  or ginst951 (i_3654, i_3423, i_3426);
  nor ginst952 (i_3657, i_3423, i_3426);
  or ginst953 (i_3658, i_3431, i_3434);
  nor ginst954 (i_3661, i_3431, i_3434);
  or ginst955 (i_3662, i_3439, i_3442);
  nor ginst956 (i_3663, i_3439, i_3442);
  and ginst957 (i_3664, i_169, i_3152, i_3447);
  and ginst958 (i_3667, i_179, i_3155, i_3447);
  and ginst959 (i_3670, i_190, i_3155, i_3451);
  and ginst960 (i_3671, i_200, i_3152, i_3451);
  not ginst961 (i_3672, i_3451);
  or ginst962 (i_3673, i_3455, i_3458);
  nor ginst963 (i_3676, i_3455, i_3458);
  or ginst964 (i_3677, i_3463, i_3466);
  nor ginst965 (i_3680, i_3463, i_3466);
  not ginst966 (i_3681, i_3493);
  and ginst967 (i_3682, i_1909, i_3415);
  not ginst968 (i_3685, i_3496);
  not ginst969 (i_3686, i_3499);
  not ginst970 (i_3687, i_3502);
  not ginst971 (i_3688, i_3505);
  not ginst972 (i_3689, i_3511);
  and ginst973 (i_3690, i_1922, i_3447);
  not ginst974 (i_3693, i_3517);
  not ginst975 (i_3694, i_3520);
  not ginst976 (i_3695, i_3523);
  not ginst977 (i_3696, i_3514);
  not ginst978 (i_3697, i_3384);
  not ginst979 (i_3700, i_3384);
  not ginst980 (i_3703, i_3490);
  not ginst981 (i_3704, i_3508);
  nand ginst982 (i_3705, i_3475, i_3630);
  nand ginst983 (i_3706, i_3472, i_3631);
  nand ginst984 (i_3707, i_3481, i_3626);
  nand ginst985 (i_3708, i_3478, i_3627);
  or ginst986 (i_3711, i_2352, i_2353, i_3632);
  or ginst987 (i_3712, i_2354, i_2355, i_3633);
  and ginst988 (i_3713, i_2632, i_3634);
  and ginst989 (i_3714, i_2634, i_3635);
  and ginst990 (i_3715, i_2636, i_3636);
  and ginst991 (i_3716, i_2638, i_3637);
  and ginst992 (i_3717, i_2640, i_3638);
  and ginst993 (i_3718, i_2642, i_3639);
  and ginst994 (i_3719, i_2644, i_3640);
  and ginst995 (i_3720, i_2646, i_3641);
  and ginst996 (i_3721, i_3557, i_3644);
  or ginst997 (i_3731, i_3651, i_3652, i_3653);
  and ginst998 (i_3734, i_3568, i_3657);
  and ginst999 (i_3740, i_3573, i_3661);
  and ginst1000 (i_3743, i_3578, i_3663);
  or ginst1001 (i_3753, i_3670, i_3671, i_3672);
  and ginst1002 (i_3756, i_3589, i_3676);
  and ginst1003 (i_3762, i_3594, i_3680);
  not ginst1004 (i_3765, i_3643);
  not ginst1005 (i_3766, i_3662);
  nand ginst1006 (i_3773, i_3705, i_3706);
  nand ginst1007 (i_3774, i_3707, i_3708);
  nand ginst1008 (i_3775, i_3628, i_3700);
  not ginst1009 (i_3776, i_3700);
  nand ginst1010 (i_3777, i_3629, i_3697);
  not ginst1011 (i_3778, i_3697);
  and ginst1012 (i_3779, i_2645, i_3712);
  and ginst1013 (i_3780, i_2647, i_3711);
  or ginst1014 (i_3786, i_3645, i_3648);
  nor ginst1015 (i_3789, i_3645, i_3648);
  or ginst1016 (i_3800, i_3664, i_3667);
  nor ginst1017 (i_3803, i_3664, i_3667);
  and ginst1018 (i_3809, i_1917, i_3654);
  and ginst1019 (i_3812, i_1917, i_3658);
  and ginst1020 (i_3815, i_1926, i_3673);
  and ginst1021 (i_3818, i_1926, i_3677);
  not ginst1022 (i_3821, i_3682);
  not ginst1023 (i_3824, i_3682);
  not ginst1024 (i_3827, i_3690);
  not ginst1025 (i_3830, i_3690);
  nand ginst1026 (i_3833, i_3773, i_3774);
  nand ginst1027 (i_3834, i_3487, i_3776);
  nand ginst1028 (i_3835, i_3484, i_3778);
  and ginst1029 (i_3838, i_3731, i_3789);
  and ginst1030 (i_3845, i_3753, i_3803);
  not ginst1031 (i_3850, i_3721);
  not ginst1032 (i_3855, i_3734);
  not ginst1033 (i_3858, i_3740);
  not ginst1034 (i_3861, i_3743);
  not ginst1035 (i_3865, i_3756);
  not ginst1036 (i_3868, i_3762);
  nand ginst1037 (i_3884, i_3775, i_3834);
  nand ginst1038 (i_3885, i_3777, i_3835);
  nand ginst1039 (i_3894, i_3721, i_3786);
  nand ginst1040 (i_3895, i_3743, i_3800);
  not ginst1041 (i_3898, i_3821);
  not ginst1042 (i_3899, i_3824);
  not ginst1043 (i_3906, i_3830);
  not ginst1044 (i_3911, i_3827);
  and ginst1045 (i_3912, i_1912, i_3786);
  not ginst1046 (i_3913, i_3812);
  and ginst1047 (i_3916, i_1917, i_3800);
  not ginst1048 (i_3917, i_3818);
  not ginst1049 (i_3920, i_3809);
  not ginst1050 (i_3921, i_3818);
  not ginst1051 (i_3924, i_3884);
  not ginst1052 (i_3925, i_3885);
  and ginst1053 (i_3926, i_3721, i_3734, i_3740, i_3838);
  nand ginst1054 (i_3930, i_3654, i_3721, i_3838);
  nand ginst1055 (i_3931, i_3658, i_3721, i_3734, i_3838);
  and ginst1056 (i_3932, i_3743, i_3756, i_3762, i_3845);
  nand ginst1057 (i_3935, i_3673, i_3743, i_3845);
  nand ginst1058 (i_3936, i_3677, i_3743, i_3756, i_3845);
  not ginst1059 (i_3937, i_3838);
  not ginst1060 (i_3940, i_3845);
  not ginst1061 (i_3947, i_3912);
  not ginst1062 (i_3948, i_3916);
  not ginst1063 (i_3950, i_3850);
  not ginst1064 (i_3953, i_3850);
  not ginst1065 (i_3956, i_3855);
  not ginst1066 (i_3959, i_3855);
  not ginst1067 (i_3962, i_3858);
  not ginst1068 (i_3965, i_3858);
  not ginst1069 (i_3968, i_3861);
  not ginst1070 (i_3971, i_3861);
  not ginst1071 (i_3974, i_3865);
  not ginst1072 (i_3977, i_3865);
  not ginst1073 (i_3980, i_3868);
  not ginst1074 (i_3983, i_3868);
  nand ginst1075 (i_3987, i_3924, i_3925);
  nand ginst1076 (i_3992, i_3765, i_3894, i_3930, i_3931);
  nand ginst1077 (i_3996, i_3766, i_3895, i_3935, i_3936);
  not ginst1078 (i_4013, i_3921);
  and ginst1079 (i_4028, i_3926, i_3932);
  nand ginst1080 (i_4029, i_3681, i_3953);
  nand ginst1081 (i_4030, i_3686, i_3959);
  nand ginst1082 (i_4031, i_3688, i_3965);
  nand ginst1083 (i_4032, i_3689, i_3971);
  nand ginst1084 (i_4033, i_3693, i_3977);
  nand ginst1085 (i_4034, i_3695, i_3983);
  not ginst1086 (i_4035, i_3926);
  not ginst1087 (i_4042, i_3953);
  not ginst1088 (i_4043, i_3956);
  nand ginst1089 (i_4044, i_3685, i_3956);
  not ginst1090 (i_4045, i_3959);
  not ginst1091 (i_4046, i_3962);
  nand ginst1092 (i_4047, i_3687, i_3962);
  not ginst1093 (i_4048, i_3965);
  not ginst1094 (i_4049, i_3971);
  not ginst1095 (i_4050, i_3977);
  not ginst1096 (i_4051, i_3980);
  nand ginst1097 (i_4052, i_3694, i_3980);
  not ginst1098 (i_4053, i_3983);
  not ginst1099 (i_4054, i_3974);
  nand ginst1100 (i_4055, i_3696, i_3974);
  and ginst1101 (i_4056, i_2304, i_3932);
  not ginst1102 (i_4057, i_3950);
  nand ginst1103 (i_4058, i_3703, i_3950);
  not ginst1104 (i_4059, i_3937);
  not ginst1105 (i_4062, i_3937);
  not ginst1106 (i_4065, i_3968);
  nand ginst1107 (i_4066, i_3704, i_3968);
  not ginst1108 (i_4067, i_3940);
  not ginst1109 (i_4070, i_3940);
  nand ginst1110 (i_4073, i_3926, i_3996);
  not ginst1111 (i_4074, i_3992);
  nand ginst1112 (i_4075, i_3493, i_4042);
  nand ginst1113 (i_4076, i_3499, i_4045);
  nand ginst1114 (i_4077, i_3505, i_4048);
  nand ginst1115 (i_4078, i_3511, i_4049);
  nand ginst1116 (i_4079, i_3517, i_4050);
  nand ginst1117 (i_4080, i_3523, i_4053);
  nand ginst1118 (i_4085, i_3496, i_4043);
  nand ginst1119 (i_4086, i_3502, i_4046);
  nand ginst1120 (i_4088, i_3520, i_4051);
  nand ginst1121 (i_4090, i_3514, i_4054);
  and ginst1122 (i_4091, i_1926, i_3996);
  or ginst1123 (i_4094, i_3605, i_4056);
  nand ginst1124 (i_4098, i_3490, i_4057);
  nand ginst1125 (i_4101, i_3508, i_4065);
  and ginst1126 (i_4104, i_4073, i_4074);
  nand ginst1127 (i_4105, i_4029, i_4075);
  nand ginst1128 (i_4106, i_3899, i_4062);
  nand ginst1129 (i_4107, i_4030, i_4076);
  nand ginst1130 (i_4108, i_4031, i_4077);
  nand ginst1131 (i_4109, i_4032, i_4078);
  nand ginst1132 (i_4110, i_3906, i_4070);
  nand ginst1133 (i_4111, i_4033, i_4079);
  nand ginst1134 (i_4112, i_4034, i_4080);
  not ginst1135 (i_4113, i_4059);
  nand ginst1136 (i_4114, i_3898, i_4059);
  not ginst1137 (i_4115, i_4062);
  nand ginst1138 (i_4116, i_4044, i_4085);
  nand ginst1139 (i_4119, i_4047, i_4086);
  not ginst1140 (i_4122, i_4070);
  nand ginst1141 (i_4123, i_4052, i_4088);
  not ginst1142 (i_4126, i_4067);
  nand ginst1143 (i_4127, i_3911, i_4067);
  nand ginst1144 (i_4128, i_4055, i_4090);
  nand ginst1145 (i_4139, i_4058, i_4098);
  nand ginst1146 (i_4142, i_4066, i_4101);
  not ginst1147 (i_4145, i_4104);
  not ginst1148 (i_4146, i_4105);
  nand ginst1149 (i_4147, i_3824, i_4115);
  not ginst1150 (i_4148, i_4107);
  not ginst1151 (i_4149, i_4108);
  not ginst1152 (i_4150, i_4109);
  nand ginst1153 (i_4151, i_3830, i_4122);
  not ginst1154 (i_4152, i_4111);
  not ginst1155 (i_4153, i_4112);
  nand ginst1156 (i_4154, i_3821, i_4113);
  nand ginst1157 (i_4161, i_3827, i_4126);
  not ginst1158 (i_4167, i_4091);
  not ginst1159 (i_4174, i_4094);
  not ginst1160 (i_4182, i_4091);
  and ginst1161 (i_4186, i_330, i_4094);
  and ginst1162 (i_4189, i_2230, i_4146);
  nand ginst1163 (i_4190, i_4106, i_4147);
  and ginst1164 (i_4191, i_2232, i_4148);
  and ginst1165 (i_4192, i_2233, i_4149);
  and ginst1166 (i_4193, i_2234, i_4150);
  nand ginst1167 (i_4194, i_4110, i_4151);
  and ginst1168 (i_4195, i_2236, i_4152);
  and ginst1169 (i_4196, i_2237, i_4153);
  nand ginst1170 (i_4197, i_4114, i_4154);
  not ginst1171 (i_4200, i_4116);
  not ginst1172 (i_4203, i_4116);
  not ginst1173 (i_4209, i_4119);
  not ginst1174 (i_4213, i_4119);
  nand ginst1175 (i_4218, i_4127, i_4161);
  not ginst1176 (i_4223, i_4123);
  and ginst1177 (i_4238, i_3917, i_4128);
  not ginst1178 (i_4239, i_4139);
  not ginst1179 (i_4241, i_4142);
  and ginst1180 (i_4242, i_330, i_4123);
  not ginst1181 (i_4247, i_4128);
  nor ginst1182 (i_4251, i_2898, i_3713, i_4189);
  not ginst1183 (i_4252, i_4190);
  nor ginst1184 (i_4253, i_2900, i_3715, i_4191);
  nor ginst1185 (i_4254, i_2901, i_3716, i_4192);
  nor ginst1186 (i_4255, i_3406, i_3717, i_4193);
  not ginst1187 (i_4256, i_4194);
  nor ginst1188 (i_4257, i_3719, i_3779, i_4195);
  nor ginst1189 (i_4258, i_3720, i_3780, i_4196);
  and ginst1190 (i_4283, i_4035, i_4167);
  and ginst1191 (i_4284, i_4035, i_4174);
  or ginst1192 (i_4287, i_3815, i_4238);
  not ginst1193 (i_4291, i_4186);
  not ginst1194 (i_4295, i_4167);
  not ginst1195 (i_4296, i_4167);
  not ginst1196 (i_4299, i_4182);
  and ginst1197 (i_4303, i_2231, i_4252);
  and ginst1198 (i_4304, i_2235, i_4256);
  not ginst1199 (i_4305, i_4197);
  or ginst1200 (i_4310, i_3992, i_4283);
  and ginst1201 (i_4316, i_4174, i_4203, i_4213);
  and ginst1202 (i_4317, i_4174, i_4209);
  and ginst1203 (i_4318, i_4128, i_4218, i_4223);
  and ginst1204 (i_4319, i_4128, i_4223);
  and ginst1205 (i_4322, i_4167, i_4209);
  nand ginst1206 (i_4325, i_3913, i_4203);
  nand ginst1207 (i_4326, i_4167, i_4203, i_4213);
  nand ginst1208 (i_4327, i_3815, i_4218);
  nand ginst1209 (i_4328, i_3917, i_4128, i_4218);
  nand ginst1210 (i_4329, i_4013, i_4247);
  not ginst1211 (i_4330, i_4247);
  and ginst1212 (i_4331, i_330, i_4094, i_4295);
  and ginst1213 (i_4335, i_2730, i_4251);
  and ginst1214 (i_4338, i_2734, i_4253);
  and ginst1215 (i_4341, i_2736, i_4254);
  and ginst1216 (i_4344, i_2738, i_4255);
  and ginst1217 (i_4347, i_2742, i_4257);
  and ginst1218 (i_4350, i_2744, i_4258);
  not ginst1219 (i_4353, i_4197);
  not ginst1220 (i_4356, i_4203);
  not ginst1221 (i_4359, i_4209);
  not ginst1222 (i_4362, i_4218);
  not ginst1223 (i_4365, i_4242);
  not ginst1224 (i_4368, i_4242);
  and ginst1225 (i_4371, i_4223, i_4223);
  nor ginst1226 (i_4376, i_2899, i_3714, i_4303);
  nor ginst1227 (i_4377, i_3642, i_3718, i_4304);
  and ginst1228 (i_4387, i_330, i_4317);
  and ginst1229 (i_4390, i_330, i_4318);
  nand ginst1230 (i_4393, i_3921, i_4330);
  not ginst1231 (i_4398, i_4287);
  not ginst1232 (i_4413, i_4284);
  nand ginst1233 (i_4416, i_3920, i_4325, i_4326);
  or ginst1234 (i_4421, i_3812, i_4322);
  nand ginst1235 (i_4427, i_3948, i_4327, i_4328);
  not ginst1236 (i_4430, i_4287);
  and ginst1237 (i_4435, i_330, i_4316);
  or ginst1238 (i_4442, i_4296, i_4331);
  and ginst1239 (i_4443, i_4174, i_4203, i_4213, i_4305);
  nand ginst1240 (i_4446, i_3809, i_4305);
  nand ginst1241 (i_4447, i_3913, i_4200, i_4305);
  nand ginst1242 (i_4448, i_4167, i_4200, i_4213, i_4305);
  not ginst1243 (i_4452, i_4356);
  nand ginst1244 (i_4458, i_4329, i_4393);
  not ginst1245 (i_4461, i_4365);
  not ginst1246 (i_4462, i_4368);
  nand ginst1247 (i_4463, i_1460, i_4371);
  not ginst1248 (i_4464, i_4371);
  not ginst1249 (i_4465, i_4310);
  nor ginst1250 (i_4468, i_4296, i_4331);
  and ginst1251 (i_4472, i_2732, i_4376);
  and ginst1252 (i_4475, i_2740, i_4377);
  not ginst1253 (i_4479, i_4310);
  not ginst1254 (i_4484, i_4353);
  not ginst1255 (i_4486, i_4359);
  nand ginst1256 (i_4487, i_4299, i_4359);
  not ginst1257 (i_4491, i_4362);
  and ginst1258 (i_4493, i_330, i_4319);
  not ginst1259 (i_4496, i_4398);
  and ginst1260 (i_4497, i_4287, i_4398);
  and ginst1261 (i_4498, i_1769, i_4442);
  nand ginst1262 (i_4503, i_3947, i_4446, i_4447, i_4448);
  not ginst1263 (i_4506, i_4413);
  not ginst1264 (i_4507, i_4435);
  not ginst1265 (i_4508, i_4421);
  nand ginst1266 (i_4509, i_4421, i_4452);
  not ginst1267 (i_4510, i_4427);
  nand ginst1268 (i_4511, i_4241, i_4427);
  nand ginst1269 (i_4515, i_4464, i_965);
  not ginst1270 (i_4526, i_4416);
  nand ginst1271 (i_4527, i_4416, i_4484);
  nand ginst1272 (i_4528, i_4182, i_4486);
  not ginst1273 (i_4529, i_4430);
  nand ginst1274 (i_4530, i_4430, i_4491);
  not ginst1275 (i_4531, i_4387);
  not ginst1276 (i_4534, i_4387);
  not ginst1277 (i_4537, i_4390);
  not ginst1278 (i_4540, i_4390);
  and ginst1279 (i_4545, i_330, i_4319, i_4496);
  and ginst1280 (i_4549, i_330, i_4443);
  nand ginst1281 (i_4552, i_4356, i_4508);
  nand ginst1282 (i_4555, i_4142, i_4510);
  not ginst1283 (i_4558, i_4493);
  nand ginst1284 (i_4559, i_4463, i_4515);
  not ginst1285 (i_4562, i_4465);
  and ginst1286 (i_4563, i_4310, i_4465);
  not ginst1287 (i_4564, i_4468);
  not ginst1288 (i_4568, i_4479);
  not ginst1289 (i_4569, i_4443);
  nand ginst1290 (i_4572, i_4353, i_4526);
  nand ginst1291 (i_4573, i_4362, i_4529);
  nand ginst1292 (i_4576, i_4487, i_4528);
  not ginst1293 (i_4581, i_4458);
  not ginst1294 (i_4584, i_4458);
  or ginst1295 (i_4587, i_2758, i_2761, i_4498);
  nor ginst1296 (i_4588, i_2758, i_2761, i_4498);
  or ginst1297 (i_4589, i_4497, i_4545);
  nand ginst1298 (i_4593, i_4509, i_4552);
  not ginst1299 (i_4596, i_4531);
  not ginst1300 (i_4597, i_4534);
  nand ginst1301 (i_4599, i_4511, i_4555);
  not ginst1302 (i_4602, i_4537);
  not ginst1303 (i_4603, i_4540);
  and ginst1304 (i_4608, i_330, i_4284, i_4562);
  not ginst1305 (i_4613, i_4503);
  not ginst1306 (i_4616, i_4503);
  nand ginst1307 (i_4619, i_4527, i_4572);
  nand ginst1308 (i_4623, i_4530, i_4573);
  not ginst1309 (i_4628, i_4588);
  nand ginst1310 (i_4629, i_4506, i_4569);
  not ginst1311 (i_4630, i_4569);
  not ginst1312 (i_4635, i_4576);
  nand ginst1313 (i_4636, i_4291, i_4576);
  not ginst1314 (i_4640, i_4581);
  nand ginst1315 (i_4641, i_4461, i_4581);
  not ginst1316 (i_4642, i_4584);
  nand ginst1317 (i_4643, i_4462, i_4584);
  nor ginst1318 (i_4644, i_4563, i_4608);
  and ginst1319 (i_4647, i_2128, i_4559);
  and ginst1320 (i_4650, i_2743, i_4559);
  not ginst1321 (i_4656, i_4549);
  not ginst1322 (i_4659, i_4549);
  not ginst1323 (i_4664, i_4564);
  and ginst1324 (i_4667, i_4587, i_4628);
  nand ginst1325 (i_4668, i_4413, i_4630);
  not ginst1326 (i_4669, i_4616);
  nand ginst1327 (i_4670, i_4239, i_4616);
  not ginst1328 (i_4673, i_4619);
  nand ginst1329 (i_4674, i_4507, i_4619);
  nand ginst1330 (i_4675, i_4186, i_4635);
  not ginst1331 (i_4676, i_4623);
  nand ginst1332 (i_4677, i_4558, i_4623);
  nand ginst1333 (i_4678, i_4365, i_4640);
  nand ginst1334 (i_4679, i_4368, i_4642);
  not ginst1335 (i_4687, i_4613);
  nand ginst1336 (i_4688, i_4568, i_4613);
  not ginst1337 (i_4691, i_4593);
  not ginst1338 (i_4694, i_4593);
  not ginst1339 (i_4697, i_4599);
  not ginst1340 (i_4700, i_4599);
  nand ginst1341 (i_4704, i_4629, i_4668);
  nand ginst1342 (i_4705, i_4139, i_4669);
  not ginst1343 (i_4706, i_4656);
  not ginst1344 (i_4707, i_4659);
  nand ginst1345 (i_4708, i_4435, i_4673);
  nand ginst1346 (i_4711, i_4636, i_4675);
  nand ginst1347 (i_4716, i_4493, i_4676);
  nand ginst1348 (i_4717, i_4641, i_4678);
  nand ginst1349 (i_4721, i_4643, i_4679);
  not ginst1350 (i_4722, i_4644);
  not ginst1351 (i_4726, i_4664);
  or ginst1352 (i_4727, i_4350, i_4647, i_4650);
  nor ginst1353 (i_4730, i_4350, i_4647, i_4650);
  nand ginst1354 (i_4733, i_4479, i_4687);
  nand ginst1355 (i_4740, i_4670, i_4705);
  nand ginst1356 (i_4743, i_4674, i_4708);
  not ginst1357 (i_4747, i_4691);
  nand ginst1358 (i_4748, i_4596, i_4691);
  not ginst1359 (i_4749, i_4694);
  nand ginst1360 (i_4750, i_4597, i_4694);
  not ginst1361 (i_4753, i_4697);
  nand ginst1362 (i_4754, i_4602, i_4697);
  not ginst1363 (i_4755, i_4700);
  nand ginst1364 (i_4756, i_4603, i_4700);
  nand ginst1365 (i_4757, i_4677, i_4716);
  nand ginst1366 (i_4769, i_4688, i_4733);
  and ginst1367 (i_4772, i_330, i_4704);
  not ginst1368 (i_4775, i_4721);
  not ginst1369 (i_4778, i_4730);
  nand ginst1370 (i_4786, i_4531, i_4747);
  nand ginst1371 (i_4787, i_4534, i_4749);
  nand ginst1372 (i_4788, i_4537, i_4753);
  nand ginst1373 (i_4789, i_4540, i_4755);
  and ginst1374 (i_4794, i_2124, i_4711);
  and ginst1375 (i_4797, i_2735, i_4711);
  and ginst1376 (i_4800, i_2127, i_4717);
  not ginst1377 (i_4805, i_4722);
  and ginst1378 (i_4808, i_4468, i_4717);
  not ginst1379 (i_4812, i_4727);
  and ginst1380 (i_4815, i_4727, i_4778);
  not ginst1381 (i_4816, i_4769);
  not ginst1382 (i_4817, i_4772);
  nand ginst1383 (i_4818, i_4748, i_4786);
  nand ginst1384 (i_4822, i_4750, i_4787);
  nand ginst1385 (i_4823, i_4754, i_4788);
  nand ginst1386 (i_4826, i_4756, i_4789);
  nand ginst1387 (i_4829, i_4726, i_4775);
  not ginst1388 (i_4830, i_4775);
  and ginst1389 (i_4831, i_2122, i_4743);
  and ginst1390 (i_4838, i_2126, i_4757);
  not ginst1391 (i_4844, i_4740);
  not ginst1392 (i_4847, i_4740);
  not ginst1393 (i_4850, i_4743);
  not ginst1394 (i_4854, i_4757);
  nand ginst1395 (i_4859, i_4772, i_4816);
  nand ginst1396 (i_4860, i_4769, i_4817);
  not ginst1397 (i_4868, i_4826);
  not ginst1398 (i_4870, i_4805);
  not ginst1399 (i_4872, i_4808);
  nand ginst1400 (i_4873, i_4664, i_4830);
  or ginst1401 (i_4876, i_4341, i_4794, i_4797);
  nor ginst1402 (i_4880, i_4341, i_4794, i_4797);
  not ginst1403 (i_4885, i_4812);
  not ginst1404 (i_4889, i_4822);
  nand ginst1405 (i_4895, i_4859, i_4860);
  not ginst1406 (i_4896, i_4844);
  nand ginst1407 (i_4897, i_4706, i_4844);
  not ginst1408 (i_4898, i_4847);
  nand ginst1409 (i_4899, i_4707, i_4847);
  nor ginst1410 (i_4900, i_4564, i_4868);
  and ginst1411 (i_4901, i_4564, i_4717, i_4757, i_4823);
  not ginst1412 (i_4902, i_4850);
  not ginst1413 (i_4904, i_4854);
  nand ginst1414 (i_4905, i_4854, i_4872);
  nand ginst1415 (i_4906, i_4829, i_4873);
  and ginst1416 (i_4907, i_2123, i_4818);
  and ginst1417 (i_4913, i_2125, i_4823);
  and ginst1418 (i_4916, i_4644, i_4818);
  not ginst1419 (i_4920, i_4880);
  and ginst1420 (i_4921, i_2184, i_4895);
  nand ginst1421 (i_4924, i_4656, i_4896);
  nand ginst1422 (i_4925, i_4659, i_4898);
  or ginst1423 (i_4926, i_4900, i_4901);
  nand ginst1424 (i_4928, i_4870, i_4889);
  not ginst1425 (i_4929, i_4889);
  nand ginst1426 (i_4930, i_4808, i_4904);
  not ginst1427 (i_4931, i_4906);
  not ginst1428 (i_4937, i_4876);
  not ginst1429 (i_4940, i_4876);
  and ginst1430 (i_4944, i_4876, i_4920);
  nand ginst1431 (i_4946, i_4897, i_4924);
  nand ginst1432 (i_4949, i_4899, i_4925);
  nand ginst1433 (i_4950, i_4902, i_4916);
  not ginst1434 (i_4951, i_4916);
  nand ginst1435 (i_4952, i_4805, i_4929);
  nand ginst1436 (i_4953, i_4905, i_4930);
  and ginst1437 (i_4954, i_2737, i_4926);
  and ginst1438 (i_4957, i_2741, i_4931);
  or ginst1439 (i_4964, i_2483, i_2764, i_4921);
  nor ginst1440 (i_4965, i_2483, i_2764, i_4921);
  not ginst1441 (i_4968, i_4949);
  nand ginst1442 (i_4969, i_4850, i_4951);
  nand ginst1443 (i_4970, i_4928, i_4952);
  and ginst1444 (i_4973, i_2739, i_4953);
  not ginst1445 (i_4978, i_4937);
  not ginst1446 (i_4979, i_4940);
  not ginst1447 (i_4980, i_4965);
  nor ginst1448 (i_4981, i_4722, i_4968);
  and ginst1449 (i_4982, i_4722, i_4743, i_4818, i_4946);
  nand ginst1450 (i_4983, i_4950, i_4969);
  not ginst1451 (i_4984, i_4970);
  and ginst1452 (i_4985, i_2121, i_4946);
  or ginst1453 (i_4988, i_4344, i_4913, i_4954);
  nor ginst1454 (i_4991, i_4344, i_4913, i_4954);
  or ginst1455 (i_4996, i_4347, i_4800, i_4957);
  nor ginst1456 (i_4999, i_4347, i_4800, i_4957);
  and ginst1457 (i_5002, i_4964, i_4980);
  or ginst1458 (i_5007, i_4981, i_4982);
  and ginst1459 (i_5010, i_2731, i_4983);
  and ginst1460 (i_5013, i_2733, i_4984);
  or ginst1461 (i_5018, i_4475, i_4838, i_4973);
  nor ginst1462 (i_5021, i_4475, i_4838, i_4973);
  not ginst1463 (i_5026, i_4991);
  not ginst1464 (i_5029, i_4999);
  and ginst1465 (i_5030, i_2729, i_5007);
  not ginst1466 (i_5039, i_4996);
  not ginst1467 (i_5042, i_4988);
  and ginst1468 (i_5045, i_4988, i_5026);
  not ginst1469 (i_5046, i_5021);
  and ginst1470 (i_5047, i_4996, i_5029);
  or ginst1471 (i_5050, i_4472, i_4831, i_5010);
  nor ginst1472 (i_5055, i_4472, i_4831, i_5010);
  or ginst1473 (i_5058, i_4338, i_4907, i_5013);
  nor ginst1474 (i_5061, i_4338, i_4907, i_5013);
  and ginst1475 (i_5066, i_4730, i_4991, i_4999, i_5021);
  not ginst1476 (i_5070, i_5018);
  and ginst1477 (i_5078, i_5018, i_5046);
  or ginst1478 (i_5080, i_4335, i_4985, i_5030);
  nor ginst1479 (i_5085, i_4335, i_4985, i_5030);
  nand ginst1480 (i_5094, i_4885, i_5039);
  not ginst1481 (i_5095, i_5039);
  not ginst1482 (i_5097, i_5042);
  and ginst1483 (i_5102, i_5050, i_5050);
  not ginst1484 (i_5103, i_5061);
  nand ginst1485 (i_5108, i_4812, i_5095);
  not ginst1486 (i_5109, i_5070);
  nand ginst1487 (i_5110, i_5070, i_5097);
  not ginst1488 (i_5111, i_5058);
  and ginst1489 (i_5114, i_1461, i_5050);
  not ginst1490 (i_5117, i_5050);
  xor ginst1491 (i_5120, i_5120_in, flip_signal);
  and ginst1492 (i_5120_in, i_5080, i_5080);
  and ginst1493 (i_5121, i_5058, i_5103);
  nand ginst1494 (i_5122, i_5094, i_5108);
  nand ginst1495 (i_5125, i_5042, i_5109);
  and ginst1496 (i_5128, i_1461, i_5080);
  and ginst1497 (i_5133, i_4880, i_5055, i_5061, i_5085);
  and ginst1498 (i_5136, i_1464, i_5055, i_5085);
  not ginst1499 (i_5139, i_5080);
  nand ginst1500 (i_5145, i_5110, i_5125);
  not ginst1501 (i_5151, i_5111);
  not ginst1502 (i_5154, i_5111);
  not ginst1503 (i_5159, i_5117);
  not ginst1504 (i_5160, i_5114);
  not ginst1505 (i_5163, i_5114);
  and ginst1506 (i_5166, i_5066, i_5133);
  and ginst1507 (i_5173, i_5066, i_5133);
  not ginst1508 (i_5174, i_5122);
  not ginst1509 (i_5177, i_5122);
  not ginst1510 (i_5182, i_5139);
  nand ginst1511 (i_5183, i_5139, i_5159);
  not ginst1512 (i_5184, i_5128);
  not ginst1513 (i_5188, i_5128);
  not ginst1514 (i_5192, i_5166);
  nor ginst1515 (i_5193, i_5136, i_5173);
  nand ginst1516 (i_5196, i_4978, i_5151);
  not ginst1517 (i_5197, i_5151);
  nand ginst1518 (i_5198, i_4979, i_5154);
  not ginst1519 (i_5199, i_5154);
  not ginst1520 (i_5201, i_5160);
  not ginst1521 (i_5203, i_5163);
  not ginst1522 (i_5205, i_5145);
  not ginst1523 (i_5209, i_5145);
  nand ginst1524 (i_5212, i_5117, i_5182);
  and ginst1525 (i_5215, i_213, i_5193);
  not ginst1526 (i_5217, i_5174);
  not ginst1527 (i_5219, i_5177);
  nand ginst1528 (i_5220, i_4937, i_5197);
  nand ginst1529 (i_5221, i_4940, i_5199);
  not ginst1530 (i_5222, i_5184);
  nand ginst1531 (i_5223, i_5184, i_5201);
  nand ginst1532 (i_5224, i_5188, i_5203);
  not ginst1533 (i_5225, i_5188);
  nand ginst1534 (i_5228, i_5183, i_5212);
  not ginst1535 (i_5231, i_5215);
  nand ginst1536 (i_5232, i_5205, i_5217);
  not ginst1537 (i_5233, i_5205);
  nand ginst1538 (i_5234, i_5209, i_5219);
  not ginst1539 (i_5235, i_5209);
  nand ginst1540 (i_5236, i_5196, i_5220);
  nand ginst1541 (i_5240, i_5198, i_5221);
  nand ginst1542 (i_5242, i_5160, i_5222);
  nand ginst1543 (i_5243, i_5163, i_5225);
  nand ginst1544 (i_5245, i_5174, i_5233);
  nand ginst1545 (i_5246, i_5177, i_5235);
  not ginst1546 (i_5250, i_5240);
  not ginst1547 (i_5253, i_5228);
  nand ginst1548 (i_5254, i_5223, i_5242);
  nand ginst1549 (i_5257, i_5224, i_5243);
  nand ginst1550 (i_5258, i_5232, i_5245);
  nand ginst1551 (i_5261, i_5234, i_5246);
  not ginst1552 (i_5266, i_5257);
  not ginst1553 (i_5269, i_5236);
  and ginst1554 (i_5277, i_2307, i_5236, i_5254);
  and ginst1555 (i_5278, i_2310, i_5250, i_5254);
  not ginst1556 (i_5279, i_5261);
  not ginst1557 (i_5283, i_5269);
  nand ginst1558 (i_5284, i_5253, i_5269);
  and ginst1559 (i_5285, i_2310, i_5236, i_5266);
  and ginst1560 (i_5286, i_2307, i_5250, i_5266);
  not ginst1561 (i_5289, i_5258);
  not ginst1562 (i_5292, i_5258);
  nand ginst1563 (i_5295, i_5228, i_5283);
  or ginst1564 (i_5298, i_5277, i_5278, i_5285, i_5286);
  not ginst1565 (i_5303, i_5279);
  not ginst1566 (i_5306, i_5279);
  nand ginst1567 (i_5309, i_5284, i_5295);
  not ginst1568 (i_5312, i_5292);
  not ginst1569 (i_5313, i_5289);
  not ginst1570 (i_5322, i_5306);
  not ginst1571 (i_5323, i_5303);
  not ginst1572 (i_5324, i_5298);
  not ginst1573 (i_5327, i_5298);
  not ginst1574 (i_5332, i_5309);
  not ginst1575 (i_5335, i_5309);
  nand ginst1576 (i_5340, i_5323, i_5324);
  nand ginst1577 (i_5341, i_5322, i_5327);
  not ginst1578 (i_5344, i_5327);
  not ginst1579 (i_5345, i_5324);
  nand ginst1580 (i_5348, i_5313, i_5332);
  nand ginst1581 (i_5349, i_5312, i_5335);
  nand ginst1582 (i_5350, i_5303, i_5345);
  nand ginst1583 (i_5351, i_5306, i_5344);
  not ginst1584 (i_5352, i_5335);
  not ginst1585 (i_5353, i_5332);
  nand ginst1586 (i_5354, i_5289, i_5353);
  nand ginst1587 (i_5355, i_5292, i_5352);
  nand ginst1588 (i_5356, i_5340, i_5350);
  nand ginst1589 (i_5357, i_5341, i_5351);
  nand ginst1590 (i_5358, i_5348, i_5354);
  nand ginst1591 (i_5359, i_5349, i_5355);
  and ginst1592 (i_5360, i_5356, i_5357);
  nand ginst1593 (i_5361, i_5358, i_5359);
  not ginst1594 (i_655, i_50);
  not ginst1595 (i_665, i_50);
  not ginst1596 (i_670, i_58);
  not ginst1597 (i_679, i_58);
  not ginst1598 (i_683, i_68);
  not ginst1599 (i_686, i_68);
  not ginst1600 (i_690, i_68);
  not ginst1601 (i_699, i_77);
  not ginst1602 (i_702, i_77);
  not ginst1603 (i_706, i_77);
  not ginst1604 (i_715, i_87);
  not ginst1605 (i_724, i_87);
  not ginst1606 (i_727, i_97);
  not ginst1607 (i_736, i_97);
  not ginst1608 (i_740, i_107);
  not ginst1609 (i_749, i_107);
  not ginst1610 (i_753, i_116);
  not ginst1611 (i_763, i_116);
  or ginst1612 (i_768, i_257, i_264);
  not ginst1613 (i_769, i_1);
  not ginst1614 (i_772, i_1);
  not ginst1615 (i_779, i_1);
  not ginst1616 (i_782, i_13);
  not ginst1617 (i_786, i_13);
  and ginst1618 (i_793, i_13, i_20);
  not ginst1619 (i_794, i_20);
  not ginst1620 (i_798, i_20);
  not ginst1621 (i_803, i_20);
  not ginst1622 (i_820, i_33);
  not ginst1623 (i_821, i_33);
  not ginst1624 (i_825, i_33);
  and ginst1625 (i_829, i_33, i_41);
  not ginst1626 (i_832, i_41);
  or ginst1627 (i_835, i_41, i_45);
  not ginst1628 (i_836, i_45);
  not ginst1629 (i_839, i_45);
  not ginst1630 (i_842, i_50);
  not ginst1631 (i_845, i_58);
  not ginst1632 (i_848, i_58);
  not ginst1633 (i_851, i_68);
  not ginst1634 (i_854, i_68);
  not ginst1635 (i_858, i_87);
  not ginst1636 (i_861, i_87);
  not ginst1637 (i_864, i_97);
  not ginst1638 (i_867, i_97);
  not ginst1639 (i_870, i_107);
  not ginst1640 (i_874, i_1);
  not ginst1641 (i_877, i_68);
  not ginst1642 (i_880, i_107);
  not ginst1643 (i_883, i_20);
  not ginst1644 (i_886, i_190);
  not ginst1645 (i_889, i_200);
  and ginst1646 (i_890, i_20, i_200);
  nand ginst1647 (i_891, i_20, i_200);
  and ginst1648 (i_892, i_20, i_179);
  not ginst1649 (i_895, i_20);
  or ginst1650 (i_896, i_33, i_349);
  nand ginst1651 (i_913, i_1, i_13);
  nand ginst1652 (i_914, i_1, i_20, i_33);
  not ginst1653 (i_915, i_20);
  not ginst1654 (i_916, i_33);
  not ginst1655 (i_917, i_179);
  not ginst1656 (i_920, i_213);
  not ginst1657 (i_923, i_343);
  not ginst1658 (i_926, i_226);
  not ginst1659 (i_929, i_232);
  not ginst1660 (i_932, i_238);
  not ginst1661 (i_935, i_244);
  not ginst1662 (i_938, i_250);
  not ginst1663 (i_941, i_257);
  not ginst1664 (i_944, i_264);
  not ginst1665 (i_947, i_270);
  not ginst1666 (i_950, i_50);
  not ginst1667 (i_953, i_58);
  not ginst1668 (i_956, i_58);
  not ginst1669 (i_959, i_97);
  not ginst1670 (i_962, i_97);
  not ginst1671 (i_965, i_330);

SatHard block1 (flip_signal, i_2243, i_150, i_4707, i_1, keyinput0, keyinput1, keyinput2, keyinput3, keyinput4, keyinput5, keyinput6, keyinput7);

endmodule
/*************** SatHard block ***************/
module SatHard (flip_signal, i_2243, i_150, i_4707, i_1, keyinput0, keyinput1, keyinput2, keyinput3, keyinput4, keyinput5, keyinput6, keyinput7);

  input i_2243, i_150, i_4707, i_1, keyinput0, keyinput1, keyinput2, keyinput3, keyinput4, keyinput5, keyinput6, keyinput7;
  output flip_signal;
  //SatHard key=10011000
  wire [3:0] sat_res_inputs;
  assign sat_res_inputs[3:0] = {i_2243, i_150, i_4707, i_1};
  wire [7:0] keyinputs, keyvalue;
  assign keyinputs[7:0] = {keyinput0, keyinput1, keyinput2, keyinput3, keyinput4, keyinput5, keyinput6, keyinput7};
  assign keyvalue[7:0] = 8'b10011000;

  wire g, g_bar;
  assign g = &(keyinputs[3:0] ^ sat_res_inputs ^ keyvalue[3:0]);
  assign g_bar = ~&(keyinputs[7:4] ^ sat_res_inputs ^ keyvalue[7:4]);
  assign flip_signal = g & g_bar;

endmodule
/*************** SatHard block ***************/
