/*************** Top Level ***************/
module c7552_AntiSAT_16_0_top (N241, N1, N5, N9, N12, N15, N18, N23, N26, N29, N32, N35, N38, N41, N44, N47, N50, N53, N54, N55, N56, N57, N58, N59, N60, N61, N62, N63, N64, N65, N66, N69, N70, N73, N74, N75, N76, N77, N78, N79, N80, N81, N82, N83, N84, N85, N86, N87, N88, N89, N94, N97, N100, N103, N106, N109, N110, N111, N112, N113, N114, N115, N118, N121, N124, N127, N130, N133, N134, N135, N138, N141, N144, N147, N150, N151, N152, N153, N154, N155, N156, N157, N158, N159, N160, N161, N162, N163, N164, N165, N166, N167, N168, N169, N170, N171, N172, N173, N174, N175, N176, N177, N178, N179, N180, N181, N182, N183, N184, N185, N186, N187, N188, N189, N190, N191, N192, N193, N194, N195, N196, N197, N198, N199, N200, N201, N202, N203, N204, N205, N206, N207, N208, N209, N210, N211, N212, N213, N214, N215, N216, N217, N218, N219, N220, N221, N222, N223, N224, N225, N226, N227, N228, N229, N230, N231, N232, N233, N234, N235, N236, N237, N238, N239, N240, N242, N245, N248, N251, N254, N257, N260, N263, N267, N271, N274, N277, N280, N283, N286, N289, N293, N296, N299, N303, N307, N310, N313, N316, N319, N322, N325, N328, N331, N334, N337, N340, N343, N346, N349, N352, N355, N358, N361, N364, N367, N382, keyinput0, keyinput1, keyinput2, keyinput3, keyinput4, keyinput5, keyinput6, keyinput7, keyinput8, keyinput9, keyinput10, keyinput11, keyinput12, keyinput13, keyinput14, keyinput15, N884, N535, N10759, N539, N10869, N10714, N10763, N515, N813, N486, N241_BUFF, N519, N556, N10760, N1110, N10351, N889, N10641, N1489, N573, N537, N10112, N10837, N553, N11333, N11342, N10870, N10706, N492, N11340, N482, N945, N10716, N505, N489, N10353, N10718, N567, N10827, N10871, N543, N10103, N1781, N1111, N509, N565, N582, N10352, N10838, N10908, N501, N545, N10905, N883, N10906, N707, N387, N511, N10025, N10109, N643, N10104, N10704, N10907, N10711, N885, N571, N551, N10350, N10102, N10632, N10111, N541, N549, N388, N11334, N547, N10713, N569, N10717, N559, N517, N10712, N10729, N1113, N10715, N513, N10839, N478, N10101, N10761, N10762, N507, N882, N10628, N10575, N10110, N1112, N10840, N10868, N881, N1490, N10574, N10576, N484, N1114, N563, N561);

  input N241, N1, N5, N9, N12, N15, N18, N23, N26, N29, N32, N35, N38, N41, N44, N47, N50, N53, N54, N55, N56, N57, N58, N59, N60, N61, N62, N63, N64, N65, N66, N69, N70, N73, N74, N75, N76, N77, N78, N79, N80, N81, N82, N83, N84, N85, N86, N87, N88, N89, N94, N97, N100, N103, N106, N109, N110, N111, N112, N113, N114, N115, N118, N121, N124, N127, N130, N133, N134, N135, N138, N141, N144, N147, N150, N151, N152, N153, N154, N155, N156, N157, N158, N159, N160, N161, N162, N163, N164, N165, N166, N167, N168, N169, N170, N171, N172, N173, N174, N175, N176, N177, N178, N179, N180, N181, N182, N183, N184, N185, N186, N187, N188, N189, N190, N191, N192, N193, N194, N195, N196, N197, N198, N199, N200, N201, N202, N203, N204, N205, N206, N207, N208, N209, N210, N211, N212, N213, N214, N215, N216, N217, N218, N219, N220, N221, N222, N223, N224, N225, N226, N227, N228, N229, N230, N231, N232, N233, N234, N235, N236, N237, N238, N239, N240, N242, N245, N248, N251, N254, N257, N260, N263, N267, N271, N274, N277, N280, N283, N286, N289, N293, N296, N299, N303, N307, N310, N313, N316, N319, N322, N325, N328, N331, N334, N337, N340, N343, N346, N349, N352, N355, N358, N361, N364, N367, N382, keyinput0, keyinput1, keyinput2, keyinput3, keyinput4, keyinput5, keyinput6, keyinput7, keyinput8, keyinput9, keyinput10, keyinput11, keyinput12, keyinput13, keyinput14, keyinput15;
  output N884, N535, N10759, N539, N10869, N10714, N10763, N515, N813, N486, N241_BUFF, N519, N556, N10760, N1110, N10351, N889, N10641, N1489, N573, N537, N10112, N10837, N553, N11333, N11342, N10870, N10706, N492, N11340, N482, N945, N10716, N505, N489, N10353, N10718, N567, N10827, N10871, N543, N10103, N1781, N1111, N509, N565, N582, N10352, N10838, N10908, N501, N545, N10905, N883, N10906, N707, N387, N511, N10025, N10109, N643, N10104, N10704, N10907, N10711, N885, N571, N551, N10350, N10102, N10632, N10111, N541, N549, N388, N11334, N547, N10713, N569, N10717, N559, N517, N10712, N10729, N1113, N10715, N513, N10839, N478, N10101, N10761, N10762, N507, N882, N10628, N10575, N10110, N1112, N10840, N10868, N881, N1490, N10574, N10576, N484, N1114, N563, N561;
  wire flip_signal;

  c7552_AntiSAT_16_0 main (N241, N1, N5, N9, N12, N15, N18, N23, N26, N29, N32, N35, N38, N41, N44, N47, N50, N53, N54, N55, N56, N57, N58, N59, N60, N61, N62, N63, N64, N65, N66, N69, N70, N73, N74, N75, N76, N77, N78, N79, N80, N81, N82, N83, N84, N85, N86, N87, N88, N89, N94, N97, N100, N103, N106, N109, N110, N111, N112, N113, N114, N115, N118, N121, N124, N127, N130, N133, N134, N135, N138, N141, N144, N147, N150, N151, N152, N153, N154, N155, N156, N157, N158, N159, N160, N161, N162, N163, N164, N165, N166, N167, N168, N169, N170, N171, N172, N173, N174, N175, N176, N177, N178, N179, N180, N181, N182, N183, N184, N185, N186, N187, N188, N189, N190, N191, N192, N193, N194, N195, N196, N197, N198, N199, N200, N201, N202, N203, N204, N205, N206, N207, N208, N209, N210, N211, N212, N213, N214, N215, N216, N217, N218, N219, N220, N221, N222, N223, N224, N225, N226, N227, N228, N229, N230, N231, N232, N233, N234, N235, N236, N237, N238, N239, N240, N242, N245, N248, N251, N254, N257, N260, N263, N267, N271, N274, N277, N280, N283, N286, N289, N293, N296, N299, N303, N307, N310, N313, N316, N319, N322, N325, N328, N331, N334, N337, N340, N343, N346, N349, N352, N355, N358, N361, N364, N367, N382, flip_signal, N241_BUFF, N387, N388, N478, N482, N484, N486, N489, N492, N501, N505, N507, N509, N511, N513, N515, N517, N519, N535, N537, N539, N541, N543, N545, N547, N549, N551, N553, N556, N559, N561, N563, N565, N567, N569, N571, N573, N582, N643, N707, N813, N881, N882, N883, N884, N885, N889, N945, N1110, N1111, N1112, N1113, N1114, N1489, N1490, N1781, N10025, N10101, N10102, N10103, N10104, N10109, N10110, N10111, N10112, N10350, N10351, N10352, N10353, N10574, N10575, N10576, N10628, N10632, N10641, N10704, N10706, N10711, N10712, N10713, N10714, N10715, N10716, N10717, N10718, N10729, N10759, N10760, N10761, N10762, N10763, N10827, N10837, N10838, N10839, N10840, N10868, N10869, N10870, N10871, N10905, N10906, N10907, N10908, N11333, N11334, N11340, N11342);
  SatHard flip (N29, N159, N325, N331, N158, N277, N299, N303, keyinput0, keyinput1, keyinput2, keyinput3, keyinput4, keyinput5, keyinput6, keyinput7, keyinput8, keyinput9, keyinput10, keyinput11, keyinput12, keyinput13, keyinput14, keyinput15, flip_signal);
endmodule
/*************** Top Level ***************/

// Main module
module c7552_AntiSAT_16_0(N241, N1, N5, N9, N12, N15, N18, N23, N26, N29, N32, N35, N38, N41, N44, N47, N50, N53, N54, N55, N56, N57, N58, N59, N60, N61, N62, N63, N64, N65, N66, N69, N70, N73, N74, N75, N76, N77, N78, N79, N80, N81, N82, N83, N84, N85, N86, N87, N88, N89, N94, N97, N100, N103, N106, N109, N110, N111, N112, N113, N114, N115, N118, N121, N124, N127, N130, N133, N134, N135, N138, N141, N144, N147, N150, N151, N152, N153, N154, N155, N156, N157, N158, N159, N160, N161, N162, N163, N164, N165, N166, N167, N168, N169, N170, N171, N172, N173, N174, N175, N176, N177, N178, N179, N180, N181, N182, N183, N184, N185, N186, N187, N188, N189, N190, N191, N192, N193, N194, N195, N196, N197, N198, N199, N200, N201, N202, N203, N204, N205, N206, N207, N208, N209, N210, N211, N212, N213, N214, N215, N216, N217, N218, N219, N220, N221, N222, N223, N224, N225, N226, N227, N228, N229, N230, N231, N232, N233, N234, N235, N236, N237, N238, N239, N240, N242, N245, N248, N251, N254, N257, N260, N263, N267, N271, N274, N277, N280, N283, N286, N289, N293, N296, N299, N303, N307, N310, N313, N316, N319, N322, N325, N328, N331, N334, N337, N340, N343, N346, N349, N352, N355, N358, N361, N364, N367, N382, flip_signal, N241_BUFF, N387, N388, N478, N482, N484, N486, N489, N492, N501, N505, N507, N509, N511, N513, N515, N517, N519, N535, N537, N539, N541, N543, N545, N547, N549, N551, N553, N556, N559, N561, N563, N565, N567, N569, N571, N573, N582, N643, N707, N813, N881, N882, N883, N884, N885, N889, N945, N1110, N1111, N1112, N1113, N1114, N1489, N1490, N1781, N10025, N10101, N10102, N10103, N10104, N10109, N10110, N10111, N10112, N10350, N10351, N10352, N10353, N10574, N10575, N10576, N10628, N10632, N10641, N10704, N10706, N10711, N10712, N10713, N10714, N10715, N10716, N10717, N10718, N10729, N10759, N10760, N10761, N10762, N10763, N10827, N10837, N10838, N10839, N10840, N10868, N10869, N10870, N10871, N10905, N10906, N10907, N10908, N11333, N11334, N11340, N11342);

  input N241, N1, N5, N9, N12, N15, N18, N23, N26, N29, N32, N35, N38, N41, N44, N47, N50, N53, N54, N55, N56, N57, N58, N59, N60, N61, N62, N63, N64, N65, N66, N69, N70, N73, N74, N75, N76, N77, N78, N79, N80, N81, N82, N83, N84, N85, N86, N87, N88, N89, N94, N97, N100, N103, N106, N109, N110, N111, N112, N113, N114, N115, N118, N121, N124, N127, N130, N133, N134, N135, N138, N141, N144, N147, N150, N151, N152, N153, N154, N155, N156, N157, N158, N159, N160, N161, N162, N163, N164, N165, N166, N167, N168, N169, N170, N171, N172, N173, N174, N175, N176, N177, N178, N179, N180, N181, N182, N183, N184, N185, N186, N187, N188, N189, N190, N191, N192, N193, N194, N195, N196, N197, N198, N199, N200, N201, N202, N203, N204, N205, N206, N207, N208, N209, N210, N211, N212, N213, N214, N215, N216, N217, N218, N219, N220, N221, N222, N223, N224, N225, N226, N227, N228, N229, N230, N231, N232, N233, N234, N235, N236, N237, N238, N239, N240, N242, N245, N248, N251, N254, N257, N260, N263, N267, N271, N274, N277, N280, N283, N286, N289, N293, N296, N299, N303, N307, N310, N313, N316, N319, N322, N325, N328, N331, N334, N337, N340, N343, N346, N349, N352, N355, N358, N361, N364, N367, N382, flip_signal;
  output N241_BUFF, N387, N388, N478, N482, N484, N486, N489, N492, N501, N505, N507, N509, N511, N513, N515, N517, N519, N535, N537, N539, N541, N543, N545, N547, N549, N551, N553, N556, N559, N561, N563, N565, N567, N569, N571, N573, N582, N643, N707, N813, N881, N882, N883, N884, N885, N889, N945, N1110, N1111, N1112, N1113, N1114, N1489, N1490, N1781, N10025, N10101, N10102, N10103, N10104, N10109, N10110, N10111, N10112, N10350, N10351, N10352, N10353, N10574, N10575, N10576, N10628, N10632, N10641, N10704, N10706, N10711, N10712, N10713, N10714, N10715, N10716, N10717, N10718, N10729, N10759, N10760, N10761, N10762, N10763, N10827, N10837, N10838, N10839, N10840, N10868, N10869, N10870, N10871, N10905, N10906, N10907, N10908, N11333, N11334, N11340, N11342;
  wire N10002, N10003, N10006, N10007, N10010, N10013, N10014, N10015, N10016, N10017, N10018, N10019, N10020, N10021, N10022, N10023, N10024, N10026, N10028, N10032, N10033, N10034, N10035, N10036, N10037, N10038, N10039, N10040, N10041, N10042, N10043, N10050, N10053, N10054, N10055, N10056, N10057, N10058, N10059, N10060, N10061, N10062, N10067, N10070, N10073, N10076, N10077, N10082, N10083, N10084, N10085, N10086, N10093, N10094, N10105, N10106, N10107, N10108, N10113, N10114, N10115, N10116, N10119, N10124, N10130, N10131, N10132, N10133, N10134, N10135, N10136, N10137, N10138, N10139, N10140, N10141, N10148, N10155, N10156, N10157, N10158, N10159, N10160, N10161, N10162, N10163, N10164, N10165, N10170, N10173, N10176, N10177, N10178, N10179, N10180, N10183, N10186, N10189, N10192, N10195, N10196, N10197, N10200, N10203, N10204, N10205, N10206, N10212, N10213, N10230, N10231, N10232, N10233, N10234, N10237, N10238, N10239, N10240, N10241, N10242, N10247, N10248, N10259, N10264, N10265, N10266, N10267, N10268, N10269, N10270, N10271, N10272, N10273, N10278, N10279, N1028, N10280, N10281, N10282, N10283, N10287, N10288, N10289, N1029, N10290, N10291, N10292, N10293, N10294, N10295, N10296, N10299, N10300, N10301, N10306, N10307, N10308, N10311, N10314, N10315, N10316, N10317, N10318, N10321, N10324, N10325, N10326, N10327, N10328, N10329, N10330, N10331, N10332, N10333, N10334, N10337, N10338, N10339, N10340, N10341, N10344, N10354, N10357, N10360, N10367, N10375, N10381, N10388, N10391, N10399, N10402, N10406, N10409, N10412, N10415, N10419, N10422, N10425, N10428, N10431, N10432, N10437, N10438, N10439, N10440, N10441, N10444, N10445, N10450, N10451, N10455, N10456, N10465, N10466, N10479, N10497, N10509, N10512, N10515, N10516, N10517, N10518, N10519, N10522, N10525, N10528, N10531, N10534, N10535, N10536, N10539, N10542, N10543, N10544, N10545, N10546, N10547, N10548, N10549, N10550, N10551, N10552, N10553, N10554, N10555, N10556, N10557, N10558, N10559, N10560, N10561, N10562, N10563, N10564, N10565, N10566, N10567, N10568, N10569, N10570, N10571, N10572, N10573, N10577, N10581, N10582, N10583, N10587, N10588, N10589, N10594, N10595, N10596, N10597, N10598, N10602, N10609, N10610, N10621, N10626, N10627, N10629, N10631, N10637, N10638, N10639, N10640, N10642, N10643, N10644, N10645, N10647, N10648, N10649, N10652, N10659, N10662, N10665, N10668, N10671, N10672, N10673, N10674, N10675, N10678, N10681, N10682, N10683, N10684, N10685, N10686, N10687, N10688, N10689, N10690, N10691, N10694, N10695, N10696, N10697, N10698, N10701, N10705, N10707, N10708, N10709, N10710, N10719, N10720, N10730, N10731, N10737, N10738, N10739, N10746, N10747, N10748, N10749, N10750, N10753, N10754, N10764, N10765, N10766, N10767, N10768, N10769, N10770, N10771, N10772, N10773, N10774, N10775, N10776, N10778, N10781, N10784, N10789, N10792, N10796, N10797, N10798, N10799, N10800, N10803, N10806, N10809, N10812, N10815, N10816, N10817, N10820, N10823, N10824, N10825, N10826, N10832, N10833, N10834, N10835, N10836, N10845, N10846, N10857, N10862, N10863, N10864, N10865, N10866, N10867, N10872, N10873, N10874, N10875, N10876, N10879, N10882, N10883, N10884, N10885, N10886, N10887, N10888, N10889, N10890, N10891, N10892, N10895, N10896, N10897, N10898, N10899, N10902, N10909, N10910, N10915, N10916, N10917, N10918, N10919, N10922, N10923, N10928, N10931, N10934, N10935, N10936, N10937, N10938, N10941, N10944, N10947, N10950, N10953, N10954, N10955, N10958, N10961, N10962, N10963, N10964, N10969, N10970, N10981, N10986, N10987, N10988, N10989, N10990, N10991, N10992, N10995, N10998, N10999, N11000, N11001, N11002, N11003, N11004, N11005, N11006, N11007, N11008, N11011, N11012, N11013, N11014, N11015, N11018, N11023, N11024, N11027, N11028, N11029, N11030, N11031, N11034, N11035, N11040, N11041, N11042, N11043, N11044, N11047, N11050, N11053, N11056, N11059, N11062, N11065, N11066, N11067, N11070, N11073, N11074, N11075, N11076, N11077, N11078, N1109, N11095, N11098, N11099, N11100, N11103, N11106, N11107, N11108, N11109, N11110, N11111, N11112, N11113, N11114, N11115, N11116, N11117, N11118, N11119, N11120, N11121, N11122, N11123, N11124, N11127, N11130, N11137, N11138, N11139, N11140, N11141, N11142, N11143, N11144, N11145, N1115, N11152, N11153, N11154, N11155, N11156, N11159, N1116, N11162, N11165, N11168, N11171, N11174, N11177, N11180, N11183, N11184, N11185, N11186, N11187, N11188, N1119, N11205, N11210, N11211, N11212, N11213, N11214, N11215, N11216, N11217, N11218, N11219, N11220, N11222, N11223, N11224, N11225, N11226, N11227, N11228, N11229, N11231, N11232, N11233, N11236, N11239, N11242, N11243, N11244, N11245, N11246, N1125, N11250, N11252, N11257, N11260, N11261, N11262, N11263, N11264, N11265, N11267, N11268, N11269, N11270, N11272, N11277, N11278, N11279, N11280, N11282, N11283, N11284, N11285, N11286, N11288, N11289, N11290, N11291, N11292, N11293, N11294, N11295, N11296, N11297, N11298, N11299, N11302, N11307, N11308, N11309, N11312, N11313, N11314, N11315, N11316, N11317, N1132, N11320, N11321, N11323, N11327, N11328, N11329, N11331, N11335, N11336, N11337, N11338, N11339, N11341, N1136, N1141, N1147, N1154, N1160, N1167, N1174, N1175, N1182, N1189, N1194, N1199, N1206, N1211, N1218, N1222, N1227, N1233, N1240, N1244, N1249, N1256, N1263, N1270, N1277, N1284, N1287, N1290, N1293, N1296, N1299, N1302, N1305, N1308, N1311, N1314, N1317, N1320, N1323, N1326, N1329, N1332, N1335, N1338, N1341, N1344, N1347, N1350, N1353, N1356, N1359, N1362, N1365, N1368, N1371, N1374, N1377, N1380, N1383, N1386, N1389, N1392, N1395, N1398, N1401, N1404, N1407, N1410, N1413, N1416, N1419, N1422, N1425, N1428, N1431, N1434, N1437, N1440, N1443, N1446, N1449, N1452, N1455, N1458, N1461, N1464, N1467, N1470, N1473, N1476, N1479, N1482, N1485, N1537, N1551, N1649, N1703, N1708, N1713, N1721, N1758, N1782, N1783, N1789, N1793, N1794, N1795, N1796, N1797, N1798, N1799, N1805, N1811, N1812, N1813, N1814, N1815, N1816, N1817, N1818, N1819, N1820, N1821, N1822, N1828, N1829, N1830, N1832, N1833, N1834, N1835, N1839, N1840, N1841, N1842, N1843, N1845, N1851, N1857, N1858, N1859, N1860, N1861, N1862, N1863, N1864, N1865, N1866, N1867, N1868, N1869, N1870, N1871, N1872, N1873, N1874, N1875, N1876, N1877, N1878, N1879, N1880, N1881, N1882, N1883, N1884, N1885, N1892, N1899, N1906, N1913, N1919, N1926, N1927, N1928, N1929, N1930, N1931, N1932, N1933, N1934, N1935, N1936, N1937, N1938, N1939, N1940, N1941, N1942, N1943, N1944, N1945, N1946, N1947, N1953, N1957, N1958, N1959, N1960, N1961, N1962, N1963, N1965, N1966, N1967, N1968, N1969, N1970, N1971, N1972, N1973, N1974, N1975, N1976, N1977, N1983, N1989, N1990, N1991, N1992, N1993, N1994, N1995, N1996, N1997, N2003, N2010, N2011, N2012, N2013, N2014, N2015, N2016, N2017, N2018, N2019, N2020, N2021, N2022, N2023, N2024, N2031, N2038, N2045, N2052, N2058, N2064, N2065, N2066, N2067, N2068, N2069, N2070, N2071, N2072, N2073, N2074, N2081, N2086, N2107, N2108, N2110, N2111, N2112, N2113, N2114, N2115, N2117, N2171, N2172, N2230, N2231, N2235, N2239, N2240, N2241, N2242, N2243, N2244, N2245, N2246, N2247, N2248, N2249, N2250, N2251, N2252, N2253, N2254, N2255, N2256, N2257, N2267, N2268, N2269, N2274, N2275, N2277, N2278, N2279, N2280, N2281, N2282, N2283, N2284, N2285, N2286, N2287, N2293, N2299, N2300, N2301, N2302, N2303, N2304, N2305, N2306, N2307, N2308, N2309, N2315, N2321, N2322, N2323, N2324, N2325, N2326, N2327, N2328, N2329, N2330, N2331, N2337, N2338, N2339, N2340, N2341, N2342, N2343, N2344, N2345, N2346, N2347, N2348, N2349, N2350, N2351, N2352, N2353, N2354, N2355, N2356, N2357, N2358, N2359, N2360, N2361, N2362, N2363, N2364, N2365, N2366, N2367, N2368, N2374, N2375, N2376, N2377, N2378, N2379, N2380, N2381, N2382, N2383, N2384, N2390, N2396, N2397, N2398, N2399, N2400, N2401, N2402, N2403, N2404, N2405, N2406, N2412, N2418, N2419, N2420, N2421, N2422, N2423, N2424, N2425, N2426, N2427, N2428, N2429, N2430, N2431, N2432, N2433, N2434, N2435, N2436, N2437, N2441, N2442, N2446, N2450, N2454, N2458, N2462, N2466, N2470, N2474, N2478, N2482, N2488, N2496, N2502, N2508, N2523, N2533, N2537, N2538, N2542, N2546, N2550, N2554, N2561, N2567, N2573, N2604, N2607, N2611, N2615, N2619, N2626, N2632, N2638, N2644, N2650, N2653, N2654, N2658, N2662, N2666, N2670, N2674, N2680, N2688, N2692, N2696, N2700, N2704, N2728, N2729, N2733, N2737, N2741, N2745, N2749, N2753, N2757, N2761, N2765, N2766, N2769, N2772, N2775, N2778, N2781, N2784, N2787, N2790, N2793, N2796, N2866, N2867, N2868, N2869, N2878, N2913, N2914, N2915, N2916, N2917, N2918, N2919, N2920, N2921, N2922, N2923, N2924, N2925, N2926, N2927, N2928, N2929, N2930, N2931, N2932, N2933, N2934, N2935, N2936, N2937, N2988, N3005, N3006, N3007, N3008, N3009, N3020, N3021, N3022, N3023, N3024, N3025, N3026, N3027, N3028, N3029, N3032, N3033, N3034, N3035, N3036, N3037, N3038, N3039, N3040, N3041, N3061, N3064, N3067, N3070, N3073, N3080, N3096, N3097, N3101, N3107, N3114, N3122, N3126, N3130, N3131, N3134, N3135, N3136, N3137, N3140, N3144, N3149, N3155, N3159, N3167, N3168, N3169, N3173, N3178, N3184, N3185, N3189, N3195, N3202, N3210, N3211, N3215, N3221, N3228, N3229, N3232, N3236, N3241, N3247, N3251, N3255, N3259, N3263, N3267, N3273, N3281, N3287, N3293, N3299, N3303, N3307, N3311, N3315, N3322, N3328, N3334, N3340, N3343, N3349, N3355, N3361, N3362, N3363, N3364, N3365, N3366, N3367, N3368, N3369, N3370, N3371, N3372, N3373, N3374, N3375, N3379, N3380, N3381, N3384, N3390, N3398, N3404, N3410, N3416, N3420, N3424, N3428, N3432, N3436, N3440, N3444, N3448, N3452, N3453, N3454, N3458, N3462, N3466, N3470, N3474, N3478, N3482, N3486, N3487, N3490, N3493, N3496, N3499, N3502, N3507, N3510, N3515, N3518, N3521, N3524, N3527, N3530, N3535, N3539, N3542, N3545, N3548, N3551, N3552, N3553, N3557, N3560, N3563, N3566, N3569, N3570, N3571, N3574, N3577, N3580, N3583, N3586, N3589, N3592, N3595, N3598, N3601, N3604, N3607, N3610, N3613, N3616, N3619, N3622, N3625, N3628, N3631, N3634, N3637, N3640, N3643, N3646, N3649, N3652, N3655, N3658, N3661, N3664, N3667, N3670, N3673, N3676, N3679, N3682, N3685, N3688, N3691, N3694, N3697, N3700, N3703, N3706, N3709, N3712, N3715, N3718, N3721, N3724, N3727, N3730, N3733, N3736, N3739, N3742, N3745, N3748, N3751, N3754, N3757, N3760, N3763, N3766, N3769, N3772, N3775, N3778, N3781, N3782, N3783, N3786, N3789, N3792, N3795, N3798, N3801, N3804, N3807, N3810, N3813, N3816, N3819, N3822, N3825, N3828, N3831, N3834, N3837, N3840, N3843, N3846, N3849, N3852, N3855, N3858, N3861, N3864, N3867, N3870, N3873, N3876, N3879, N3882, N3885, N3888, N3891, N3953, N3954, N3955, N3956, N3958, N3964, N4193, N4303, N4308, N4313, N4326, N4327, N4333, N4334, N4411, N4412, N4463, N4464, N4465, N4466, N4467, N4468, N4469, N4470, N4471, N4472, N4473, N4474, N4475, N4476, N4477, N4478, N4479, N4480, N4481, N4482, N4483, N4484, N4485, N4486, N4487, N4488, N4489, N4490, N4491, N4492, N4493, N4494, N4495, N4496, N4497, N4498, N4499, N4500, N4501, N4502, N4503, N4504, N4505, N4506, N4507, N4508, N4509, N4510, N4511, N4512, N4513, N4514, N4515, N4516, N4517, N4518, N4519, N4520, N4521, N4522, N4523, N4524, N4525, N4526, N4527, N4528, N4529, N4530, N4531, N4532, N4533, N4534, N4535, N4536, N4537, N4538, N4539, N4540, N4541, N4542, N4543, N4544, N4545, N4549, N4555, N4562, N4563, N4566, N4570, N4575, N4576, N4577, N4581, N4586, N4592, N4593, N4597, N4603, N4610, N4611, N4612, N4613, N4614, N4615, N4616, N4617, N4618, N4619, N4620, N4621, N4622, N4623, N4624, N4625, N4626, N4627, N4628, N4629, N4630, N4631, N4632, N4633, N4634, N4635, N4636, N4637, N4638, N4639, N4640, N4641, N4642, N4643, N4644, N4645, N4646, N4647, N4648, N4649, N4650, N4651, N4652, N4653, N4656, N4657, N4661, N4667, N467, N4674, N4675, N4678, N4682, N4687, N469, N4693, N4694, N4695, N4696, N4697, N4698, N4699, N4700, N4701, N4702, N4706, N4711, N4717, N4718, N4722, N4728, N4735, N4743, N4744, N4745, N4746, N4747, N4748, N4749, N4750, N4751, N4752, N4753, N4754, N4755, N4756, N4757, N4758, N4759, N4760, N4761, N4762, N4763, N4764, N4765, N4766, N4767, N4768, N4769, N4775, N4776, N4777, N4778, N4779, N4780, N4781, N4782, N4783, N4784, N4789, N4790, N4793, N4794, N4795, N4796, N4799, N4800, N4801, N4802, N4803, N4806, N4809, N4810, N4813, N4814, N4817, N4820, N4823, N4826, N4829, N4832, N4835, N4838, N4841, N4844, N4847, N4850, N4853, N4856, N4859, N4862, N4865, N4868, N4871, N4874, N4877, N4880, N4883, N4886, N4889, N4892, N4895, N4898, N4901, N4904, N4907, N4910, N4913, N4916, N4919, N4922, N4925, N4928, N4931, N4934, N4937, N494, N4940, N4943, N4946, N4949, N4952, N4955, N4958, N4961, N4964, N4967, N4970, N4973, N4976, N4979, N4982, N4985, N4988, N4991, N4994, N4997, N5000, N5003, N5006, N5009, N5012, N5015, N5018, N5021, N5024, N5027, N5030, N5033, N5036, N5039, N5042, N5045, N5046, N5047, N5048, N5049, N5052, N5055, N5058, N5061, N5064, N5065, N5066, N5067, N5068, N5071, N5074, N5077, N5080, N5083, N5086, N5089, N5092, N5095, N5098, N5101, N5104, N5107, N5110, N5111, N5112, N5113, N5114, N5117, N5120, N5123, N5126, N5129, N5132, N5135, N5138, N5141, N5144, N5147, N5150, N5153, N5156, N5159, N5162, N5165, N5166, N5167, N5168, N5169, N5170, N5171, N5172, N5173, N5174, N5175, N5176, N5177, N5178, N5179, N5180, N5181, N5182, N5183, N5184, N5185, N5186, N5187, N5188, N5189, N5190, N5191, N5192, N5193, N5196, N5197, N5198, N5199, N5200, N5201, N5202, N5203, N5204, N5205, N5206, N5207, N5208, N5209, N5210, N5211, N5212, N5213, N528, N5283, N5284, N5285, N5286, N5287, N5288, N5289, N5290, N5291, N5292, N5293, N5294, N5295, N5296, N5297, N5298, N5299, N5300, N5314, N5315, N5316, N5317, N5318, N5319, N5320, N5321, N5322, N5323, N5324, N5363, N5364, N5365, N5366, N5367, N5425, N5426, N5427, N5429, N5430, N5431, N5432, N5433, N5451, N5452, N5453, N5454, N5455, N5456, N5457, N5469, N5474, N5475, N5476, N5477, N5571, N5572, N5573, N5574, N5584, N5585, N5586, N5587, N5602, N5603, N5604, N5605, N5631, N5632, N5640, N5654, N5670, N5683, N5690, N5697, N5707, N5718, N5728, N5735, N5736, N5740, N5744, N5747, N575, N5751, N5755, N5758, N5762, N5766, N5769, N5770, N5771, N5778, N578, N5789, N5799, N5807, N5821, N5837, N585, N5850, N5856, N5863, N5870, N5881, N5892, N5898, N590, N5905, N5915, N5926, N593, N5936, N5943, N5944, N5945, N5946, N5947, N5948, N5949, N5950, N5951, N5952, N5953, N5954, N5955, N5956, N5957, N5958, N5959, N596, N5960, N5966, N5967, N5968, N5969, N5970, N5971, N5972, N5973, N5974, N5975, N5976, N5977, N5978, N5979, N5980, N5981, N5989, N599, N5990, N5991, N5996, N6000, N6003, N6009, N6014, N6018, N6021, N6022, N6023, N6024, N6025, N6026, N6027, N6028, N6029, N6030, N6031, N6032, N6033, N6034, N6035, N6036, N6037, N6038, N6039, N604, N6040, N6041, N6047, N6052, N6056, N6059, N6060, N6061, N6062, N6063, N6064, N6065, N6066, N6067, N6068, N6069, N6070, N6071, N6072, N6073, N6074, N6075, N6076, N6077, N6078, N6079, N6083, N6087, N609, N6090, N6091, N6092, N6093, N6094, N6095, N6096, N6097, N6098, N6099, N6100, N6101, N6102, N6103, N6104, N6105, N6106, N6107, N6108, N6109, N6110, N6111, N6112, N6113, N6114, N6115, N6116, N6117, N6118, N6119, N6120, N6121, N6122, N6123, N6124, N6125, N6126, N6127, N6131, N6135, N6136, N6137, N614, N6141, N6145, N6148, N6149, N6150, N6151, N6152, N6153, N6154, N6155, N6156, N6157, N6158, N6159, N6160, N6161, N6162, N6163, N6164, N6165, N6166, N6170, N6174, N6177, N6181, N6182, N6183, N6184, N6185, N6186, N6187, N6188, N6189, N6190, N6191, N6192, N6193, N6194, N6195, N6196, N6199, N6202, N6203, N6204, N6207, N6210, N6213, N6214, N6217, N6220, N6223, N6224, N6225, N6226, N6227, N6228, N6229, N6230, N6231, N6232, N6235, N6236, N6239, N6240, N6241, N6242, N6243, N6246, N6249, N625, N6252, N6255, N6256, N6257, N6258, N6259, N6260, N6261, N6262, N6263, N6266, N628, N632, N636, N641, N642, N644, N651, N6540, N6541, N6542, N6543, N6544, N6545, N6546, N6547, N6555, N6556, N6557, N6558, N6559, N6560, N6561, N6569, N657, N6594, N6595, N6596, N6597, N6598, N6599, N660, N6600, N6601, N6602, N6603, N6604, N6605, N6606, N6621, N6622, N6623, N6624, N6625, N6626, N6627, N6628, N6629, N6639, N6640, N6641, N6642, N6643, N6644, N6645, N6646, N6647, N6648, N6649, N6650, N6651, N6652, N6653, N6654, N6655, N6656, N6657, N6658, N6659, N666, N6660, N6661, N6668, N6677, N6678, N6679, N6680, N6681, N6682, N6683, N6684, N6685, N6686, N6687, N6688, N6689, N6690, N6702, N6703, N6704, N6705, N6706, N6707, N6708, N6709, N6710, N6711, N6712, N672, N6729, N673, N6730, N6731, N6732, N6733, N6734, N6735, N6736, N674, N6741, N6742, N6743, N6744, N6751, N6752, N6753, N6754, N6755, N6756, N6757, N6758, N676, N6761, N6762, N6766, N6767, N6768, N6769, N6770, N6771, N6772, N6773, N6774, N6775, N6776, N6777, N6778, N6779, N6780, N6781, N6782, N6783, N6784, N6787, N6788, N6789, N6790, N6791, N6792, N6793, N6794, N6795, N6796, N6797, N6800, N6803, N6806, N6809, N6812, N6815, N6818, N682, N6821, N6824, N6827, N6830, N6833, N6836, N6837, N6838, N6839, N6840, N6841, N6842, N6843, N6844, N6845, N6848, N6849, N6850, N6851, N6852, N6853, N6854, N6855, N6856, N6857, N6858, N6859, N6860, N6861, N6862, N6863, N6864, N6865, N6866, N6867, N6870, N6871, N6872, N6873, N6874, N6875, N6876, N6877, N6878, N6879, N688, N6880, N6881, N6884, N6885, N6886, N6887, N6888, N6889, N689, N6890, N6891, N6892, N6893, N6894, N6901, N6912, N6923, N6929, N6936, N6946, N695, N6957, N6967, N6968, N6969, N6970, N6977, N6988, N6998, N700, N7006, N7020, N7036, N7049, N705, N7055, N7056, N7057, N706, N7060, N7061, N7062, N7063, N7064, N7065, N7066, N7067, N7068, N7073, N7077, N708, N7080, N7086, N7091, N7095, N7098, N7099, N7100, N7103, N7104, N7105, N7106, N7107, N7114, N7125, N7136, N7142, N7149, N715, N7159, N7170, N7180, N7187, N7188, N7191, N7194, N7198, N7202, N7205, N7209, N721, N7213, N7216, N7219, N7222, N7229, N7240, N7250, N7258, N727, N7272, N7288, N7301, N7307, N7314, N7318, N7322, N7325, N7328, N733, N7331, N7334, N7337, N734, N7340, N7343, N7346, N7351, N7355, N7358, N7364, N7369, N7373, N7376, N7377, N7378, N7381, N7384, N7387, N7391, N7394, N7398, N7402, N7405, N7408, N7411, N7414, N7417, N742, N7420, N7423, N7426, N7429, N7432, N7435, N7438, N7441, N7444, N7447, N7450, N7453, N7456, N7459, N7462, N7465, N7468, N7471, N7474, N7477, N7478, N7479, N748, N7482, N7485, N7488, N749, N7491, N7494, N7497, N750, N7500, N7503, N7506, N7509, N7512, N7515, N7518, N7521, N7524, N7527, N7530, N7533, N7536, N7539, N7542, N7545, N7548, N7551, N7552, N7553, N7556, N7557, N7558, N7559, N7560, N7563, N7566, N7569, N7572, N7573, N7574, N7577, N758, N7580, N7581, N7582, N7585, N7588, N759, N7591, N7609, N7613, N762, N7620, N7649, N7650, N7655, N7659, N7668, N7671, N768, N774, N7744, N780, N7822, N7825, N7826, N7852, N786, N794, N800, N806, N8114, N8117, N812, N8131, N8134, N814, N8144, N8145, N8146, N8156, N8166, N8169, N8183, N8186, N8196, N8200, N8204, N8208, N821, N8216, N8217, N8218, N8219, N8232, N8233, N8242, N8243, N8244, N8245, N8246, N8247, N8248, N8249, N8250, N8251, N8252, N8253, N8254, N8260, N8261, N8262, N8269, N827, N8274, N8275, N8276, N8277, N8278, N8279, N8280, N8281, N8282, N8283, N8284, N8285, N8288, N8294, N8295, N8296, N8297, N8298, N8307, N8315, N8317, N8319, N8321, N8322, N8323, N8324, N8325, N8326, N833, N8333, N8337, N8338, N8339, N8340, N8341, N8342, N8343, N8344, N8345, N8346, N8347, N8348, N8349, N8350, N8351, N8352, N8353, N8354, N8355, N8356, N8357, N8358, N8365, N8369, N8370, N8371, N8372, N8373, N8374, N8375, N8376, N8377, N8378, N8379, N8380, N8381, N8382, N8383, N8384, N8385, N8386, N8387, N8388, N8389, N839, N8390, N8391, N8392, N8393, N8394, N8404, N8405, N8409, N8410, N8411, N8412, N8415, N8416, N8417, N8418, N8421, N8430, N8433, N8434, N8435, N8436, N8437, N8438, N8439, N8440, N8441, N8442, N8443, N8444, N8447, N8448, N8449, N845, N8450, N8451, N8452, N8453, N8454, N8455, N8456, N8457, N8460, N8463, N8466, N8469, N8470, N8471, N8474, N8477, N8480, N8483, N8484, N8485, N8488, N8489, N8490, N8491, N8492, N8493, N8494, N8495, N8496, N8497, N8500, N8501, N8502, N8503, N8504, N8505, N8506, N8507, N8508, N8509, N8510, N8511, N8512, N8513, N8514, N8515, N8516, N8517, N8518, N8519, N8522, N8525, N8528, N853, N8531, N8534, N8537, N8538, N8539, N8540, N8541, N8545, N8546, N8547, N8548, N8551, N8552, N8553, N8554, N8555, N8558, N8561, N8564, N8565, N8566, N8569, N8572, N8575, N8578, N8579, N8580, N8583, N8586, N8589, N859, N8592, N8595, N8598, N8601, N8604, N8607, N8608, N8609, N8610, N8615, N8616, N8617, N8618, N8619, N8624, N8625, N8626, N8627, N8632, N8633, N8634, N8637, N8638, N8639, N8644, N8645, N8646, N8647, N8648, N865, N8653, N8654, N8655, N8660, N8663, N8666, N8669, N8672, N8675, N8678, N8681, N8684, N8687, N8690, N8693, N8696, N8699, N8702, N8705, N8708, N871, N8711, N8714, N8717, N8718, N8721, N8724, N8727, N8730, N8733, N8734, N8735, N8738, N8741, N8744, N8747, N8750, N8753, N8754, N8755, N8756, N8757, N8760, N8763, N8766, N8769, N8772, N8775, N8778, N8781, N8784, N8787, N8790, N8793, N8796, N8799, N8802, N8805, N8808, N8811, N8814, N8815, N8816, N8817, N8818, N8840, N8857, N886, N8861, N8862, N8863, N8864, N8865, N8866, N887, N8871, N8874, N8878, N8879, N8880, N8881, N8882, N8883, N8884, N8885, N8886, N8887, N8888, N8898, N8902, N8920, N8924, N8927, N8931, N8943, N8950, N8956, N8959, N8960, N8963, N8966, N8991, N8992, N8995, N8996, N9001, N9005, N9024, N9025, N9029, N9035, N9053, N9054, N9064, N9065, N9066, N9067, N9068, N9071, N9072, N9073, N9074, N9077, N9079, N9082, N9083, N9086, N9087, N9088, N9089, N9092, N9093, N9094, N9095, N9098, N9099, N9103, N9107, N9111, N9117, N9127, N9146, N9149, N9159, N9160, N9161, N9165, N9169, N9173, N9179, N9180, N9181, N9182, N9183, N9193, N9203, N9206, N9220, N9223, N9234, N9235, N9236, N9237, N9238, N9242, N9243, N9244, N9245, N9246, N9247, N9248, N9249, N9250, N9251, N9252, N9256, N9257, N9258, N9259, N9260, N9261, N9262, N9265, N9268, N9271, N9272, N9273, N9274, N9275, N9276, N9280, N9285, N9286, N9287, N9288, N9290, N9292, N9294, N9296, N9297, N9298, N9299, N9300, N9301, N9307, N9314, N9315, N9318, N9319, N9320, N9321, N9322, N9323, N9324, N9326, N9332, N9339, N9344, N9352, N9354, N9356, N9358, N9359, N9360, N9361, N9362, N9363, N9364, N9365, N9366, N9367, N9368, N9369, N9370, N9371, N9372, N9375, N9381, N9382, N9383, N9384, N9385, N9392, N9393, N9394, N9395, N9396, N9397, N9398, N9399, N9400, N9401, N9402, N9407, N9408, N9412, N9413, N9414, N9415, N9416, N9417, N9418, N9419, N9420, N9421, N9422, N9423, N9426, N9429, N9432, N9435, N9442, N9445, N9454, N9455, N9456, N9459, N9460, N9461, N9462, N9465, N9466, N9467, N9468, N9473, N9476, N9477, N9478, N9485, N9488, N9493, N9494, N9495, N9498, N9499, N9500, N9505, N9506, N9507, N9508, N9509, N9514, N9515, N9516, N9517, N9520, N9526, N9531, N9539, N9540, N9541, N9543, N9551, N9555, N9556, N9557, N9560, N9561, N9562, N9563, N9564, N9565, N9566, N9567, N9568, N9569, N957, N9570, N9571, N9575, N9579, N9581, N9582, N9585, N9591, N9592, N9593, N9594, N9595, N9596, N9597, N9598, N9599, N9600, N9601, N9602, N9603, N9604, N9605, N9608, N9611, N9612, N9613, N9614, N9615, N9616, N9617, N9618, N9621, N9622, N9623, N9624, N9626, N9629, N9632, N9635, N9642, N9645, N9646, N9649, N9650, N9653, N9656, N9659, N9660, N9661, N9662, N9663, N9666, N9667, N9670, N9671, N9674, N9675, N9678, N9679, N9682, N9685, N9690, N9691, N9692, N9695, N9698, N9702, N9707, N9710, N9711, N9714, N9715, N9716, N9717, N9720, N9721, N9722, N9723, N9726, N9727, N9732, N9733, N9734, N9735, N9736, N9737, N9738, N9739, N9740, N9741, N9742, N9754, N9758, N9762, N9763, N9764, N9765, N9766, N9767, N9768, N9769, N9773, N9774, N9775, N9779, N9784, N9785, N9786, N9790, N9791, N9795, N9796, N9797, N9798, N9799, N9800, N9801, N9802, N9803, N9805, N9806, N9809, N9813, N9814, N9815, N9816, N9817, N9820, N9825, N9826, N9827, N9828, N9829, N9830, N9835, N9836, N9837, N9838, N9846, N9847, N9862, N9863, N9866, N9873, N9876, N9890, N9891, N9892, N9893, N9894, N9895, N9896, N9897, N9898, N9899, N9900, N9901, N9902, N9903, N9904, N9905, N9906, N9907, N9908, N9909, N9910, N9911, N9917, N9923, N9924, N9925, N9932, N9935, N9938, N9939, N9945, N9946, N9947, N9948, N9949, N9953, N9954, N9955, N9956, N9957, N9958, N9959, N9960, N9961, N9964, N9967, N9968, N9969, N9970, N9971, N9972, N9973, N9974, N9975, N9976, N9977, N9978, N9979, N9982, N9983, N9986, N9989, N9992, N9995, N9996, N9997, N9998, N9999, N10104_in;

  not ginst1 (N10002, N9717);
  nand ginst2 (N10003, N9722, N9876);
  not ginst3 (N10006, N9723);
  nand ginst4 (N10007, N9829, N9830);
  nand ginst5 (N10010, N9827, N9828);
  and ginst6 (N10013, N8269, N8307, N9791);
  and ginst7 (N10014, N8269, N8307, N9344, N9758);
  and ginst8 (N10015, N367, N8269, N8307, N9344, N9754);
  and ginst9 (N10016, N8394, N8421, N9786);
  and ginst10 (N10017, N8394, N8421, N9332, N9820);
  and ginst11 (N10018, N8394, N8421, N9786);
  and ginst12 (N10019, N8394, N8421, N9332, N9820);
  and ginst13 (N10020, N8262, N8298, N9809);
  and ginst14 (N10021, N8262, N8298, N9385, N9779);
  and ginst15 (N10022, N367, N8262, N8298, N9385, N9775);
  not ginst16 (N10023, N9945);
  not ginst17 (N10024, N9946);
  nand ginst18 (N10025, N9740, N9893);
  not ginst19 (N10026, N9923);
  not ginst20 (N10028, N9924);
  nand ginst21 (N10032, N8595, N9897);
  nand ginst22 (N10033, N8598, N9899);
  nand ginst23 (N10034, N8601, N9901);
  nand ginst24 (N10035, N8604, N9903);
  nand ginst25 (N10036, N4803, N9906);
  nand ginst26 (N10037, N4806, N9908);
  nand ginst27 (N10038, N8627, N9910);
  and ginst28 (N10039, N8298, N9809);
  and ginst29 (N10040, N8298, N9385, N9779);
  and ginst30 (N10041, N367, N8298, N9385, N9775);
  and ginst31 (N10042, N9385, N9779);
  and ginst32 (N10043, N367, N9385, N9775);
  nand ginst33 (N10050, N8727, N9938);
  not ginst34 (N10053, N9817);
  and ginst35 (N10054, N9029, N9817);
  and ginst36 (N10055, N8394, N9786);
  and ginst37 (N10056, N8394, N9332, N9820);
  and ginst38 (N10057, N8307, N9791);
  and ginst39 (N10058, N8307, N9344, N9758);
  and ginst40 (N10059, N367, N8307, N9344, N9754);
  and ginst41 (N10060, N9344, N9758);
  and ginst42 (N10061, N367, N9344, N9754);
  nand ginst43 (N10062, N4997, N9947);
  nand ginst44 (N10067, N8811, N9953);
  nand ginst45 (N10070, N9836, N9955);
  nand ginst46 (N10073, N9838, N9956);
  nand ginst47 (N10076, N9068, N9957);
  nand ginst48 (N10077, N9074, N9959);
  nand ginst49 (N10082, N9089, N9967);
  nand ginst50 (N10083, N9095, N9969);
  nand ginst51 (N10084, N4871, N9971);
  nand ginst52 (N10085, N6214, N9973);
  nand ginst53 (N10086, N6217, N9975);
  nand ginst54 (N10093, N5027, N9995);
  nand ginst55 (N10094, N6232, N9997);
  or ginst56 (N10101, N10013, N10014, N10015, N9238, N9732);
  or ginst57 (N10102, N10016, N10017, N9339, N9526, N9734);
  or ginst58 (N10103, N10018, N10019, N9339, N9531, N9735);
  xor ginst59 (N10104, N10104_in, flip_signal);
  or ginst60 (N10104_in, N10020, N10021, N10022, N9242, N9736);
  and ginst61 (N10105, N9894, N9925);
  and ginst62 (N10106, N9895, N9925);
  and ginst63 (N10107, N9896, N9925);
  and ginst64 (N10108, N8253, N9925);
  nand ginst65 (N10109, N10032, N9898);
  nand ginst66 (N10110, N10033, N9900);
  nand ginst67 (N10111, N10034, N9902);
  nand ginst68 (N10112, N10035, N9904);
  nand ginst69 (N10113, N10036, N9907);
  nand ginst70 (N10114, N10037, N9909);
  nand ginst71 (N10115, N10038, N9911);
  or ginst72 (N10116, N10039, N10040, N10041, N9265);
  or ginst73 (N10119, N10042, N10043, N9809);
  not ginst74 (N10124, N9925);
  and ginst75 (N10130, N9768, N9925);
  not ginst76 (N10131, N9932);
  not ginst77 (N10132, N9935);
  and ginst78 (N10133, N8920, N9932);
  nand ginst79 (N10134, N10050, N9939);
  not ginst80 (N10135, N9983);
  nand ginst81 (N10136, N9324, N9983);
  not ginst82 (N10137, N9986);
  nand ginst83 (N10138, N9784, N9986);
  and ginst84 (N10139, N10053, N9785);
  or ginst85 (N10140, N10055, N10056, N8943, N9790);
  or ginst86 (N10141, N10057, N10058, N10059, N9268);
  or ginst87 (N10148, N10060, N10061, N9791);
  nand ginst88 (N10155, N10062, N9948);
  not ginst89 (N10156, N9989);
  nand ginst90 (N10157, N9805, N9989);
  not ginst91 (N10158, N9992);
  nand ginst92 (N10159, N9806, N9992);
  not ginst93 (N10160, N9949);
  nand ginst94 (N10161, N10067, N9954);
  not ginst95 (N10162, N10007);
  nand ginst96 (N10163, N10007, N9825);
  not ginst97 (N10164, N10010);
  nand ginst98 (N10165, N10010, N9826);
  nand ginst99 (N10170, N10076, N9958);
  nand ginst100 (N10173, N10077, N9960);
  not ginst101 (N10176, N9961);
  nand ginst102 (N10177, N9082, N9961);
  not ginst103 (N10178, N9964);
  nand ginst104 (N10179, N9086, N9964);
  nand ginst105 (N10180, N10082, N9968);
  nand ginst106 (N10183, N10083, N9970);
  nand ginst107 (N10186, N10084, N9972);
  nand ginst108 (N10189, N10085, N9974);
  nand ginst109 (N10192, N10086, N9976);
  not ginst110 (N10195, N9979);
  nand ginst111 (N10196, N9979, N9982);
  nand ginst112 (N10197, N10093, N9996);
  nand ginst113 (N10200, N10094, N9998);
  not ginst114 (N10203, N9999);
  nand ginst115 (N10204, N10002, N9999);
  not ginst116 (N10205, N10003);
  nand ginst117 (N10206, N10003, N10006);
  nand ginst118 (N10212, N10070, N4308);
  nand ginst119 (N10213, N10073, N4313);
  and ginst120 (N10230, N10131, N9774);
  nand ginst121 (N10231, N10135, N8730);
  nand ginst122 (N10232, N10137, N9478);
  or ginst123 (N10233, N10054, N10139);
  nand ginst124 (N10234, N10140, N7100);
  nand ginst125 (N10237, N10156, N9485);
  nand ginst126 (N10238, N10158, N9488);
  nand ginst127 (N10239, N10162, N9517);
  nand ginst128 (N10240, N10164, N9520);
  not ginst129 (N10241, N10070);
  not ginst130 (N10242, N10073);
  nand ginst131 (N10247, N10176, N8146);
  nand ginst132 (N10248, N10178, N8156);
  nand ginst133 (N10259, N10195, N9692);
  nand ginst134 (N10264, N10203, N9717);
  nand ginst135 (N10265, N10205, N9723);
  and ginst136 (N10266, N10026, N10124);
  and ginst137 (N10267, N10028, N10124);
  and ginst138 (N10268, N10124, N9742);
  and ginst139 (N10269, N10124, N6923);
  nand ginst140 (N10270, N10116, N6762);
  nand ginst141 (N10271, N10241, N3061);
  nand ginst142 (N10272, N10242, N3064);
  buf ginst143 (N10273, N10116);
  and ginst144 (N10278, N10141, N5697, N5707, N5718, N5728);
  and ginst145 (N10279, N10141, N5707, N5718, N5728);
  and ginst146 (N1028, N382, N641);
  and ginst147 (N10280, N10141, N5718, N5728);
  and ginst148 (N10281, N10141, N5728);
  and ginst149 (N10282, N10141, N6784);
  not ginst150 (N10283, N10119);
  and ginst151 (N10287, N10148, N5905, N5915, N5926, N5936);
  and ginst152 (N10288, N10148, N5915, N5926, N5936);
  and ginst153 (N10289, N10148, N5926, N5936);
  nand ginst154 (N1029, N382, N705);
  and ginst155 (N10290, N10148, N5936);
  and ginst156 (N10291, N10148, N6881);
  and ginst157 (N10292, N10124, N8898);
  nand ginst158 (N10293, N10136, N10231);
  nand ginst159 (N10294, N10138, N10232);
  nand ginst160 (N10295, N10233, N8412);
  and ginst161 (N10296, N10234, N8959);
  nand ginst162 (N10299, N10157, N10237);
  nand ginst163 (N10300, N10159, N10238);
  or ginst164 (N10301, N10133, N10230);
  nand ginst165 (N10306, N10163, N10239);
  nand ginst166 (N10307, N10165, N10240);
  buf ginst167 (N10308, N10148);
  buf ginst168 (N10311, N10141);
  not ginst169 (N10314, N10170);
  nand ginst170 (N10315, N10170, N9071);
  not ginst171 (N10316, N10173);
  nand ginst172 (N10317, N10173, N9077);
  nand ginst173 (N10318, N10177, N10247);
  nand ginst174 (N10321, N10179, N10248);
  not ginst175 (N10324, N10180);
  nand ginst176 (N10325, N10180, N9092);
  not ginst177 (N10326, N10183);
  nand ginst178 (N10327, N10183, N9098);
  not ginst179 (N10328, N10186);
  nand ginst180 (N10329, N10186, N9674);
  not ginst181 (N10330, N10189);
  nand ginst182 (N10331, N10189, N9678);
  not ginst183 (N10332, N10192);
  nand ginst184 (N10333, N10192, N9977);
  nand ginst185 (N10334, N10196, N10259);
  not ginst186 (N10337, N10197);
  nand ginst187 (N10338, N10197, N9710);
  not ginst188 (N10339, N10200);
  nand ginst189 (N10340, N10200, N9714);
  nand ginst190 (N10341, N10204, N10264);
  nand ginst191 (N10344, N10206, N10265);
  or ginst192 (N10350, N10105, N10266);
  or ginst193 (N10351, N10106, N10267);
  or ginst194 (N10352, N10107, N10268);
  or ginst195 (N10353, N10108, N10269);
  and ginst196 (N10354, N10270, N8857);
  nand ginst197 (N10357, N10212, N10271);
  nand ginst198 (N10360, N10213, N10272);
  or ginst199 (N10367, N10282, N7620);
  or ginst200 (N10375, N10291, N7671);
  or ginst201 (N10381, N10130, N10292);
  and ginst202 (N10388, N10114, N10134, N10293, N10294);
  and ginst203 (N10391, N10295, N9582);
  and ginst204 (N10399, N10113, N10115, N10299, N10300);
  and ginst205 (N10402, N10155, N10161, N10306, N10307);
  or ginst206 (N10406, N10287, N3229, N6888, N6889, N6890);
  or ginst207 (N10409, N10288, N3232, N6891, N6892);
  or ginst208 (N10412, N10289, N3236, N6893);
  or ginst209 (N10415, N10290, N3241);
  or ginst210 (N10419, N10278, N3137, N6791, N6792, N6793);
  or ginst211 (N10422, N10279, N3140, N6794, N6795);
  or ginst212 (N10425, N10280, N3144, N6796);
  or ginst213 (N10428, N10281, N3149);
  nand ginst214 (N10431, N10314, N8117);
  nand ginst215 (N10432, N10316, N8134);
  nand ginst216 (N10437, N10324, N8169);
  nand ginst217 (N10438, N10326, N8186);
  nand ginst218 (N10439, N10328, N9117);
  nand ginst219 (N10440, N10330, N9127);
  nand ginst220 (N10441, N10332, N9682);
  nand ginst221 (N10444, N10337, N9183);
  nand ginst222 (N10445, N10339, N9193);
  not ginst223 (N10450, N10296);
  and ginst224 (N10451, N10296, N4193);
  not ginst225 (N10455, N10308);
  nand ginst226 (N10456, N10308, N8242);
  not ginst227 (N10465, N10311);
  nand ginst228 (N10466, N10311, N8247);
  not ginst229 (N10479, N10273);
  not ginst230 (N10497, N10301);
  nand ginst231 (N10509, N10315, N10431);
  nand ginst232 (N10512, N10317, N10432);
  not ginst233 (N10515, N10318);
  nand ginst234 (N10516, N10318, N8632);
  not ginst235 (N10517, N10321);
  nand ginst236 (N10518, N10321, N8637);
  nand ginst237 (N10519, N10325, N10437);
  nand ginst238 (N10522, N10327, N10438);
  nand ginst239 (N10525, N10329, N10439);
  nand ginst240 (N10528, N10331, N10440);
  nand ginst241 (N10531, N10333, N10441);
  not ginst242 (N10534, N10334);
  nand ginst243 (N10535, N10334, N9695);
  nand ginst244 (N10536, N10338, N10444);
  nand ginst245 (N10539, N10340, N10445);
  not ginst246 (N10542, N10341);
  nand ginst247 (N10543, N10341, N9720);
  not ginst248 (N10544, N10344);
  nand ginst249 (N10545, N10344, N9726);
  and ginst250 (N10546, N10450, N5631);
  not ginst251 (N10547, N10391);
  and ginst252 (N10548, N10391, N8950);
  and ginst253 (N10549, N10367, N5165);
  not ginst254 (N10550, N10354);
  and ginst255 (N10551, N10354, N3126);
  nand ginst256 (N10552, N10455, N7411);
  and ginst257 (N10553, N10375, N9539);
  and ginst258 (N10554, N10375, N9540);
  and ginst259 (N10555, N10375, N9541);
  and ginst260 (N10556, N10375, N6761);
  not ginst261 (N10557, N10406);
  nand ginst262 (N10558, N10406, N8243);
  not ginst263 (N10559, N10409);
  nand ginst264 (N10560, N10409, N8244);
  not ginst265 (N10561, N10412);
  nand ginst266 (N10562, N10412, N8245);
  not ginst267 (N10563, N10415);
  nand ginst268 (N10564, N10415, N8246);
  nand ginst269 (N10565, N10465, N7426);
  not ginst270 (N10566, N10419);
  nand ginst271 (N10567, N10419, N8248);
  not ginst272 (N10568, N10422);
  nand ginst273 (N10569, N10422, N8249);
  not ginst274 (N10570, N10425);
  nand ginst275 (N10571, N10425, N8250);
  not ginst276 (N10572, N10428);
  nand ginst277 (N10573, N10428, N8251);
  not ginst278 (N10574, N10399);
  not ginst279 (N10575, N10402);
  not ginst280 (N10576, N10388);
  and ginst281 (N10577, N10388, N10399, N10402);
  and ginst282 (N10581, N10273, N10360, N9543);
  and ginst283 (N10582, N10273, N10357, N9905);
  not ginst284 (N10583, N10367);
  and ginst285 (N10587, N10367, N5735);
  and ginst286 (N10588, N10367, N3135);
  not ginst287 (N10589, N10375);
  and ginst288 (N10594, N10381, N7149, N7159, N7170, N7180);
  and ginst289 (N10595, N10381, N7159, N7170, N7180);
  and ginst290 (N10596, N10381, N7170, N7180);
  and ginst291 (N10597, N10381, N7180);
  and ginst292 (N10598, N10381, N8444);
  buf ginst293 (N10602, N10381);
  nand ginst294 (N10609, N10515, N7479);
  nand ginst295 (N10610, N10517, N7491);
  nand ginst296 (N10621, N10534, N9149);
  nand ginst297 (N10626, N10542, N9206);
  nand ginst298 (N10627, N10544, N9223);
  or ginst299 (N10628, N10451, N10546);
  and ginst300 (N10629, N10547, N9733);
  and ginst301 (N10631, N10550, N5166);
  nand ginst302 (N10632, N10456, N10552);
  nand ginst303 (N10637, N10557, N7414);
  nand ginst304 (N10638, N10559, N7417);
  nand ginst305 (N10639, N10561, N7420);
  nand ginst306 (N10640, N10563, N7423);
  nand ginst307 (N10641, N10466, N10565);
  nand ginst308 (N10642, N10566, N7429);
  nand ginst309 (N10643, N10568, N7432);
  nand ginst310 (N10644, N10570, N7435);
  nand ginst311 (N10645, N10572, N7438);
  and ginst312 (N10647, N10577, N886, N887);
  and ginst313 (N10648, N10360, N10479, N8857);
  and ginst314 (N10649, N10357, N10479, N7609);
  or ginst315 (N10652, N10598, N8966);
  or ginst316 (N10659, N10594, N4675, N8451, N8452, N8453);
  or ginst317 (N10662, N10595, N4678, N8454, N8455);
  or ginst318 (N10665, N10596, N4682, N8456);
  or ginst319 (N10668, N10597, N4687);
  not ginst320 (N10671, N10509);
  nand ginst321 (N10672, N10509, N8615);
  not ginst322 (N10673, N10512);
  nand ginst323 (N10674, N10512, N8624);
  nand ginst324 (N10675, N10516, N10609);
  nand ginst325 (N10678, N10518, N10610);
  not ginst326 (N10681, N10519);
  nand ginst327 (N10682, N10519, N8644);
  not ginst328 (N10683, N10522);
  nand ginst329 (N10684, N10522, N8653);
  not ginst330 (N10685, N10525);
  nand ginst331 (N10686, N10525, N9454);
  not ginst332 (N10687, N10528);
  nand ginst333 (N10688, N10528, N9459);
  not ginst334 (N10689, N10531);
  nand ginst335 (N10690, N10531, N9978);
  nand ginst336 (N10691, N10535, N10621);
  not ginst337 (N10694, N10536);
  nand ginst338 (N10695, N10536, N9493);
  not ginst339 (N10696, N10539);
  nand ginst340 (N10697, N10539, N9498);
  nand ginst341 (N10698, N10543, N10626);
  nand ginst342 (N10701, N10545, N10627);
  or ginst343 (N10704, N10548, N10629);
  and ginst344 (N10705, N10583, N3159);
  or ginst345 (N10706, N10551, N10631);
  and ginst346 (N10707, N10589, N9737);
  and ginst347 (N10708, N10589, N9738);
  and ginst348 (N10709, N10589, N9243);
  and ginst349 (N10710, N10589, N5892);
  nand ginst350 (N10711, N10558, N10637);
  nand ginst351 (N10712, N10560, N10638);
  nand ginst352 (N10713, N10562, N10639);
  nand ginst353 (N10714, N10564, N10640);
  nand ginst354 (N10715, N10567, N10642);
  nand ginst355 (N10716, N10569, N10643);
  nand ginst356 (N10717, N10571, N10644);
  nand ginst357 (N10718, N10573, N10645);
  not ginst358 (N10719, N10602);
  nand ginst359 (N10720, N10602, N9244);
  not ginst360 (N10729, N10647);
  and ginst361 (N10730, N10583, N5178);
  and ginst362 (N10731, N10583, N2533);
  nand ginst363 (N10737, N10671, N7447);
  nand ginst364 (N10738, N10673, N7465);
  or ginst365 (N10739, N10581, N10582, N10648, N10649);
  nand ginst366 (N10746, N10681, N7503);
  nand ginst367 (N10747, N10683, N7521);
  nand ginst368 (N10748, N10685, N8678);
  nand ginst369 (N10749, N10687, N8690);
  nand ginst370 (N10750, N10689, N9685);
  nand ginst371 (N10753, N10694, N8757);
  nand ginst372 (N10754, N10696, N8769);
  or ginst373 (N10759, N10549, N10705);
  or ginst374 (N10760, N10553, N10707);
  or ginst375 (N10761, N10554, N10708);
  or ginst376 (N10762, N10555, N10709);
  or ginst377 (N10763, N10556, N10710);
  nand ginst378 (N10764, N10719, N8580);
  and ginst379 (N10765, N10652, N9890);
  and ginst380 (N10766, N10652, N9891);
  and ginst381 (N10767, N10652, N9892);
  and ginst382 (N10768, N10652, N8252);
  not ginst383 (N10769, N10659);
  nand ginst384 (N10770, N10659, N9245);
  not ginst385 (N10771, N10662);
  nand ginst386 (N10772, N10662, N9246);
  not ginst387 (N10773, N10665);
  nand ginst388 (N10774, N10665, N9247);
  not ginst389 (N10775, N10668);
  nand ginst390 (N10776, N10668, N9248);
  or ginst391 (N10778, N10587, N10730);
  or ginst392 (N10781, N10588, N10731);
  not ginst393 (N10784, N10652);
  nand ginst394 (N10789, N10672, N10737);
  nand ginst395 (N10792, N10674, N10738);
  not ginst396 (N10796, N10675);
  nand ginst397 (N10797, N10675, N8633);
  not ginst398 (N10798, N10678);
  nand ginst399 (N10799, N10678, N8638);
  nand ginst400 (N10800, N10682, N10746);
  nand ginst401 (N10803, N10684, N10747);
  nand ginst402 (N10806, N10686, N10748);
  nand ginst403 (N10809, N10688, N10749);
  nand ginst404 (N10812, N10690, N10750);
  not ginst405 (N10815, N10691);
  nand ginst406 (N10816, N10691, N9866);
  nand ginst407 (N10817, N10695, N10753);
  nand ginst408 (N10820, N10697, N10754);
  not ginst409 (N10823, N10698);
  nand ginst410 (N10824, N10698, N9505);
  not ginst411 (N10825, N10701);
  nand ginst412 (N10826, N10701, N9514);
  nand ginst413 (N10827, N10720, N10764);
  nand ginst414 (N10832, N10769, N8583);
  nand ginst415 (N10833, N10771, N8586);
  nand ginst416 (N10834, N10773, N8589);
  nand ginst417 (N10835, N10775, N8592);
  not ginst418 (N10836, N10739);
  buf ginst419 (N10837, N10778);
  buf ginst420 (N10838, N10778);
  buf ginst421 (N10839, N10781);
  buf ginst422 (N10840, N10781);
  nand ginst423 (N10845, N10796, N7482);
  nand ginst424 (N10846, N10798, N7494);
  nand ginst425 (N10857, N10815, N9473);
  nand ginst426 (N10862, N10823, N8781);
  nand ginst427 (N10863, N10825, N8799);
  and ginst428 (N10864, N10023, N10784);
  and ginst429 (N10865, N10024, N10784);
  and ginst430 (N10866, N10784, N9739);
  and ginst431 (N10867, N10784, N7136);
  nand ginst432 (N10868, N10770, N10832);
  nand ginst433 (N10869, N10772, N10833);
  nand ginst434 (N10870, N10774, N10834);
  nand ginst435 (N10871, N10776, N10835);
  not ginst436 (N10872, N10789);
  nand ginst437 (N10873, N10789, N8616);
  not ginst438 (N10874, N10792);
  nand ginst439 (N10875, N10792, N8625);
  nand ginst440 (N10876, N10797, N10845);
  nand ginst441 (N10879, N10799, N10846);
  not ginst442 (N10882, N10800);
  nand ginst443 (N10883, N10800, N8645);
  not ginst444 (N10884, N10803);
  nand ginst445 (N10885, N10803, N8654);
  not ginst446 (N10886, N10806);
  nand ginst447 (N10887, N10806, N9455);
  not ginst448 (N10888, N10809);
  nand ginst449 (N10889, N10809, N9460);
  not ginst450 (N10890, N10812);
  nand ginst451 (N10891, N10812, N9862);
  nand ginst452 (N10892, N10816, N10857);
  not ginst453 (N10895, N10817);
  nand ginst454 (N10896, N10817, N9494);
  not ginst455 (N10897, N10820);
  nand ginst456 (N10898, N10820, N9499);
  nand ginst457 (N10899, N10824, N10862);
  nand ginst458 (N10902, N10826, N10863);
  or ginst459 (N10905, N10765, N10864);
  or ginst460 (N10906, N10766, N10865);
  or ginst461 (N10907, N10767, N10866);
  or ginst462 (N10908, N10768, N10867);
  nand ginst463 (N10909, N10872, N7450);
  nand ginst464 (N10910, N10874, N7468);
  nand ginst465 (N10915, N10882, N7506);
  nand ginst466 (N10916, N10884, N7524);
  nand ginst467 (N10917, N10886, N8681);
  nand ginst468 (N10918, N10888, N8693);
  nand ginst469 (N10919, N10890, N9462);
  nand ginst470 (N10922, N10895, N8760);
  nand ginst471 (N10923, N10897, N8772);
  nand ginst472 (N10928, N10873, N10909);
  nand ginst473 (N10931, N10875, N10910);
  not ginst474 (N10934, N10876);
  nand ginst475 (N10935, N10876, N8634);
  not ginst476 (N10936, N10879);
  nand ginst477 (N10937, N10879, N8639);
  nand ginst478 (N10938, N10883, N10915);
  nand ginst479 (N10941, N10885, N10916);
  nand ginst480 (N10944, N10887, N10917);
  nand ginst481 (N10947, N10889, N10918);
  nand ginst482 (N10950, N10891, N10919);
  not ginst483 (N10953, N10892);
  nand ginst484 (N10954, N10892, N9476);
  nand ginst485 (N10955, N10896, N10922);
  nand ginst486 (N10958, N10898, N10923);
  not ginst487 (N10961, N10899);
  nand ginst488 (N10962, N10899, N9506);
  not ginst489 (N10963, N10902);
  nand ginst490 (N10964, N10902, N9515);
  nand ginst491 (N10969, N10934, N7485);
  nand ginst492 (N10970, N10936, N7497);
  nand ginst493 (N10981, N10953, N8718);
  nand ginst494 (N10986, N10961, N8784);
  nand ginst495 (N10987, N10963, N8802);
  not ginst496 (N10988, N10928);
  nand ginst497 (N10989, N10928, N8617);
  not ginst498 (N10990, N10931);
  nand ginst499 (N10991, N10931, N8626);
  nand ginst500 (N10992, N10935, N10969);
  nand ginst501 (N10995, N10937, N10970);
  not ginst502 (N10998, N10938);
  nand ginst503 (N10999, N10938, N8646);
  not ginst504 (N11000, N10941);
  nand ginst505 (N11001, N10941, N8655);
  not ginst506 (N11002, N10944);
  nand ginst507 (N11003, N10944, N9456);
  not ginst508 (N11004, N10947);
  nand ginst509 (N11005, N10947, N9461);
  not ginst510 (N11006, N10950);
  nand ginst511 (N11007, N10950, N9465);
  nand ginst512 (N11008, N10954, N10981);
  not ginst513 (N11011, N10955);
  nand ginst514 (N11012, N10955, N9495);
  not ginst515 (N11013, N10958);
  nand ginst516 (N11014, N10958, N9500);
  nand ginst517 (N11015, N10962, N10986);
  nand ginst518 (N11018, N10964, N10987);
  nand ginst519 (N11023, N10988, N7453);
  nand ginst520 (N11024, N10990, N7471);
  nand ginst521 (N11027, N10998, N7509);
  nand ginst522 (N11028, N11000, N7527);
  nand ginst523 (N11029, N11002, N8684);
  nand ginst524 (N11030, N11004, N8696);
  nand ginst525 (N11031, N11006, N8702);
  nand ginst526 (N11034, N11011, N8763);
  nand ginst527 (N11035, N11013, N8775);
  not ginst528 (N11040, N10992);
  nand ginst529 (N11041, N10992, N8294);
  not ginst530 (N11042, N10995);
  nand ginst531 (N11043, N10995, N8295);
  nand ginst532 (N11044, N10989, N11023);
  nand ginst533 (N11047, N10991, N11024);
  nand ginst534 (N11050, N10999, N11027);
  nand ginst535 (N11053, N11001, N11028);
  nand ginst536 (N11056, N11003, N11029);
  nand ginst537 (N11059, N11005, N11030);
  nand ginst538 (N11062, N11007, N11031);
  not ginst539 (N11065, N11008);
  nand ginst540 (N11066, N11008, N9477);
  nand ginst541 (N11067, N11012, N11034);
  nand ginst542 (N11070, N11014, N11035);
  not ginst543 (N11073, N11015);
  nand ginst544 (N11074, N11015, N9507);
  not ginst545 (N11075, N11018);
  nand ginst546 (N11076, N11018, N9516);
  nand ginst547 (N11077, N11040, N7488);
  nand ginst548 (N11078, N11042, N7500);
  and ginst549 (N1109, N469, N596);
  nand ginst550 (N11095, N11065, N8721);
  nand ginst551 (N11098, N11073, N8787);
  nand ginst552 (N11099, N11075, N8805);
  nand ginst553 (N1110, N242, N593);
  nand ginst554 (N11100, N11041, N11077);
  nand ginst555 (N11103, N11043, N11078);
  not ginst556 (N11106, N11056);
  nand ginst557 (N11107, N11056, N9319);
  not ginst558 (N11108, N11059);
  nand ginst559 (N11109, N11059, N9320);
  not ginst560 (N1111, N625);
  not ginst561 (N11110, N11067);
  nand ginst562 (N11111, N11067, N9381);
  not ginst563 (N11112, N11070);
  nand ginst564 (N11113, N11070, N9382);
  not ginst565 (N11114, N11044);
  nand ginst566 (N11115, N11044, N8618);
  not ginst567 (N11116, N11047);
  nand ginst568 (N11117, N11047, N8619);
  not ginst569 (N11118, N11050);
  nand ginst570 (N11119, N11050, N8647);
  nand ginst571 (N1112, N242, N593);
  not ginst572 (N11120, N11053);
  nand ginst573 (N11121, N11053, N8648);
  not ginst574 (N11122, N11062);
  nand ginst575 (N11123, N11062, N9466);
  nand ginst576 (N11124, N11066, N11095);
  nand ginst577 (N11127, N11074, N11098);
  nand ginst578 (N1113, N469, N596);
  nand ginst579 (N11130, N11076, N11099);
  nand ginst580 (N11137, N11106, N8687);
  nand ginst581 (N11138, N11108, N8699);
  nand ginst582 (N11139, N11110, N8766);
  not ginst583 (N1114, N625);
  nand ginst584 (N11140, N11112, N8778);
  nand ginst585 (N11141, N11114, N7456);
  nand ginst586 (N11142, N11116, N7474);
  nand ginst587 (N11143, N11118, N7512);
  nand ginst588 (N11144, N11120, N7530);
  nand ginst589 (N11145, N11122, N8705);
  not ginst590 (N1115, N871);
  and ginst591 (N11152, N10283, N11103, N8871);
  and ginst592 (N11153, N10283, N11100, N7655);
  and ginst593 (N11154, N10119, N11103, N9551);
  and ginst594 (N11155, N10119, N11100, N9917);
  nand ginst595 (N11156, N11107, N11137);
  nand ginst596 (N11159, N11109, N11138);
  buf ginst597 (N1116, N590);
  nand ginst598 (N11162, N11111, N11139);
  nand ginst599 (N11165, N11113, N11140);
  nand ginst600 (N11168, N11115, N11141);
  nand ginst601 (N11171, N11117, N11142);
  nand ginst602 (N11174, N11119, N11143);
  nand ginst603 (N11177, N11121, N11144);
  nand ginst604 (N11180, N11123, N11145);
  not ginst605 (N11183, N11124);
  nand ginst606 (N11184, N11124, N9468);
  not ginst607 (N11185, N11127);
  nand ginst608 (N11186, N11127, N9508);
  not ginst609 (N11187, N11130);
  nand ginst610 (N11188, N11130, N9509);
  buf ginst611 (N1119, N628);
  or ginst612 (N11205, N11152, N11153, N11154, N11155);
  nand ginst613 (N11210, N11183, N8724);
  nand ginst614 (N11211, N11185, N8790);
  nand ginst615 (N11212, N11187, N8808);
  not ginst616 (N11213, N11168);
  nand ginst617 (N11214, N11168, N8260);
  not ginst618 (N11215, N11171);
  nand ginst619 (N11216, N11171, N8261);
  not ginst620 (N11217, N11174);
  nand ginst621 (N11218, N11174, N8296);
  not ginst622 (N11219, N11177);
  nand ginst623 (N11220, N11177, N8297);
  and ginst624 (N11222, N11159, N1218, N9575);
  and ginst625 (N11223, N11156, N1218, N8927);
  and ginst626 (N11224, N11159, N750, N9935);
  and ginst627 (N11225, N10132, N11156, N750);
  and ginst628 (N11226, N10497, N11165, N9608);
  and ginst629 (N11227, N10497, N11162, N9001);
  and ginst630 (N11228, N10301, N11165, N9949);
  and ginst631 (N11229, N10160, N10301, N11162);
  not ginst632 (N11231, N11180);
  nand ginst633 (N11232, N11180, N9467);
  nand ginst634 (N11233, N11184, N11210);
  nand ginst635 (N11236, N11186, N11211);
  nand ginst636 (N11239, N11188, N11212);
  nand ginst637 (N11242, N11213, N7459);
  nand ginst638 (N11243, N11215, N7462);
  nand ginst639 (N11244, N11217, N7515);
  nand ginst640 (N11245, N11219, N7518);
  not ginst641 (N11246, N11205);
  buf ginst642 (N1125, N682);
  nand ginst643 (N11250, N11231, N8708);
  or ginst644 (N11252, N11222, N11223, N11224, N11225);
  or ginst645 (N11257, N11226, N11227, N11228, N11229);
  nand ginst646 (N11260, N11214, N11242);
  nand ginst647 (N11261, N11216, N11243);
  nand ginst648 (N11262, N11218, N11244);
  nand ginst649 (N11263, N11220, N11245);
  not ginst650 (N11264, N11233);
  nand ginst651 (N11265, N11233, N9322);
  not ginst652 (N11267, N11236);
  nand ginst653 (N11268, N11236, N9383);
  not ginst654 (N11269, N11239);
  nand ginst655 (N11270, N11239, N9384);
  nand ginst656 (N11272, N11232, N11250);
  not ginst657 (N11277, N11261);
  and ginst658 (N11278, N10273, N11260);
  not ginst659 (N11279, N11263);
  and ginst660 (N11280, N10119, N11262);
  nand ginst661 (N11282, N11264, N8714);
  not ginst662 (N11283, N11252);
  nand ginst663 (N11284, N11267, N8793);
  nand ginst664 (N11285, N11269, N8796);
  not ginst665 (N11286, N11257);
  and ginst666 (N11288, N10479, N11277);
  and ginst667 (N11289, N10283, N11279);
  not ginst668 (N11290, N11272);
  nand ginst669 (N11291, N11272, N9321);
  nand ginst670 (N11292, N11265, N11282);
  nand ginst671 (N11293, N11268, N11284);
  nand ginst672 (N11294, N11270, N11285);
  nand ginst673 (N11295, N11290, N8711);
  not ginst674 (N11296, N11292);
  not ginst675 (N11297, N11294);
  and ginst676 (N11298, N10301, N11293);
  or ginst677 (N11299, N11278, N11288);
  or ginst678 (N11302, N11280, N11289);
  nand ginst679 (N11307, N11291, N11295);
  and ginst680 (N11308, N11296, N1218);
  and ginst681 (N11309, N10497, N11297);
  nand ginst682 (N11312, N11246, N11302);
  nand ginst683 (N11313, N10836, N11299);
  not ginst684 (N11314, N11299);
  not ginst685 (N11315, N11302);
  and ginst686 (N11316, N11307, N750);
  or ginst687 (N11317, N11298, N11309);
  buf ginst688 (N1132, N628);
  nand ginst689 (N11320, N11205, N11315);
  nand ginst690 (N11321, N10739, N11314);
  or ginst691 (N11323, N11308, N11316);
  nand ginst692 (N11327, N11312, N11320);
  nand ginst693 (N11328, N11313, N11321);
  nand ginst694 (N11329, N11286, N11317);
  not ginst695 (N11331, N11317);
  not ginst696 (N11333, N11327);
  not ginst697 (N11334, N11328);
  nand ginst698 (N11335, N11257, N11331);
  nand ginst699 (N11336, N11283, N11323);
  not ginst700 (N11337, N11323);
  nand ginst701 (N11338, N11329, N11335);
  nand ginst702 (N11339, N11252, N11337);
  not ginst703 (N11340, N11338);
  nand ginst704 (N11341, N11336, N11339);
  not ginst705 (N11342, N11341);
  buf ginst706 (N1136, N682);
  buf ginst707 (N1141, N628);
  buf ginst708 (N1147, N682);
  buf ginst709 (N1154, N632);
  buf ginst710 (N1160, N676);
  and ginst711 (N1167, N614, N700);
  and ginst712 (N1174, N614, N700);
  buf ginst713 (N1175, N682);
  buf ginst714 (N1182, N676);
  not ginst715 (N1189, N657);
  not ginst716 (N1194, N676);
  not ginst717 (N1199, N682);
  not ginst718 (N1206, N689);
  buf ginst719 (N1211, N695);
  not ginst720 (N1218, N750);
  not ginst721 (N1222, N1028);
  buf ginst722 (N1227, N632);
  buf ginst723 (N1233, N676);
  buf ginst724 (N1240, N632);
  buf ginst725 (N1244, N676);
  buf ginst726 (N1249, N689);
  buf ginst727 (N1256, N689);
  buf ginst728 (N1263, N695);
  buf ginst729 (N1270, N689);
  buf ginst730 (N1277, N689);
  buf ginst731 (N1284, N700);
  buf ginst732 (N1287, N614);
  buf ginst733 (N1290, N666);
  buf ginst734 (N1293, N660);
  buf ginst735 (N1296, N651);
  buf ginst736 (N1299, N614);
  buf ginst737 (N1302, N644);
  buf ginst738 (N1305, N700);
  buf ginst739 (N1308, N614);
  buf ginst740 (N1311, N614);
  buf ginst741 (N1314, N666);
  buf ginst742 (N1317, N660);
  buf ginst743 (N1320, N651);
  buf ginst744 (N1323, N644);
  buf ginst745 (N1326, N609);
  buf ginst746 (N1329, N604);
  buf ginst747 (N1332, N742);
  buf ginst748 (N1335, N599);
  buf ginst749 (N1338, N727);
  buf ginst750 (N1341, N721);
  buf ginst751 (N1344, N715);
  buf ginst752 (N1347, N734);
  buf ginst753 (N1350, N708);
  buf ginst754 (N1353, N609);
  buf ginst755 (N1356, N604);
  buf ginst756 (N1359, N742);
  buf ginst757 (N1362, N734);
  buf ginst758 (N1365, N599);
  buf ginst759 (N1368, N727);
  buf ginst760 (N1371, N721);
  buf ginst761 (N1374, N715);
  buf ginst762 (N1377, N708);
  buf ginst763 (N1380, N806);
  buf ginst764 (N1383, N800);
  buf ginst765 (N1386, N794);
  buf ginst766 (N1389, N786);
  buf ginst767 (N1392, N780);
  buf ginst768 (N1395, N774);
  buf ginst769 (N1398, N768);
  buf ginst770 (N1401, N762);
  buf ginst771 (N1404, N806);
  buf ginst772 (N1407, N800);
  buf ginst773 (N1410, N794);
  buf ginst774 (N1413, N780);
  buf ginst775 (N1416, N774);
  buf ginst776 (N1419, N768);
  buf ginst777 (N1422, N762);
  buf ginst778 (N1425, N786);
  buf ginst779 (N1428, N636);
  buf ginst780 (N1431, N636);
  buf ginst781 (N1434, N865);
  buf ginst782 (N1437, N859);
  buf ginst783 (N1440, N853);
  buf ginst784 (N1443, N845);
  buf ginst785 (N1446, N839);
  buf ginst786 (N1449, N833);
  buf ginst787 (N1452, N827);
  buf ginst788 (N1455, N821);
  buf ginst789 (N1458, N814);
  buf ginst790 (N1461, N865);
  buf ginst791 (N1464, N859);
  buf ginst792 (N1467, N853);
  buf ginst793 (N1470, N839);
  buf ginst794 (N1473, N833);
  buf ginst795 (N1476, N827);
  buf ginst796 (N1479, N821);
  buf ginst797 (N1482, N845);
  buf ginst798 (N1485, N814);
  not ginst799 (N1489, N1109);
  buf ginst800 (N1490, N1116);
  and ginst801 (N1537, N614, N957);
  and ginst802 (N1551, N614, N957);
  and ginst803 (N1649, N1029, N636);
  buf ginst804 (N1703, N957);
  nor ginst805 (N1708, N614, N957);
  buf ginst806 (N1713, N957);
  nor ginst807 (N1721, N614, N957);
  buf ginst808 (N1758, N1029);
  and ginst809 (N1781, N163, N1116);
  and ginst810 (N1782, N170, N1125);
  not ginst811 (N1783, N1125);
  not ginst812 (N1789, N1136);
  and ginst813 (N1793, N169, N1125);
  and ginst814 (N1794, N168, N1125);
  and ginst815 (N1795, N167, N1125);
  and ginst816 (N1796, N166, N1136);
  and ginst817 (N1797, N165, N1136);
  and ginst818 (N1798, N164, N1136);
  not ginst819 (N1799, N1147);
  not ginst820 (N1805, N1160);
  and ginst821 (N1811, N177, N1147);
  and ginst822 (N1812, N176, N1147);
  and ginst823 (N1813, N175, N1147);
  and ginst824 (N1814, N174, N1147);
  and ginst825 (N1815, N173, N1147);
  and ginst826 (N1816, N157, N1160);
  and ginst827 (N1817, N156, N1160);
  and ginst828 (N1818, N155, N1160);
  and ginst829 (N1819, N154, N1160);
  and ginst830 (N1820, N153, N1160);
  not ginst831 (N1821, N1284);
  not ginst832 (N1822, N1287);
  not ginst833 (N1828, N1290);
  not ginst834 (N1829, N1293);
  not ginst835 (N1830, N1296);
  not ginst836 (N1832, N1299);
  not ginst837 (N1833, N1302);
  not ginst838 (N1834, N1305);
  not ginst839 (N1835, N1308);
  not ginst840 (N1839, N1311);
  not ginst841 (N1840, N1314);
  not ginst842 (N1841, N1317);
  not ginst843 (N1842, N1320);
  not ginst844 (N1843, N1323);
  not ginst845 (N1845, N1175);
  not ginst846 (N1851, N1182);
  and ginst847 (N1857, N181, N1175);
  and ginst848 (N1858, N171, N1175);
  and ginst849 (N1859, N180, N1175);
  and ginst850 (N1860, N179, N1175);
  and ginst851 (N1861, N178, N1175);
  and ginst852 (N1862, N161, N1182);
  and ginst853 (N1863, N151, N1182);
  and ginst854 (N1864, N160, N1182);
  and ginst855 (N1865, N159, N1182);
  and ginst856 (N1866, N158, N1182);
  not ginst857 (N1867, N1326);
  not ginst858 (N1868, N1329);
  not ginst859 (N1869, N1332);
  not ginst860 (N1870, N1335);
  not ginst861 (N1871, N1338);
  not ginst862 (N1872, N1341);
  not ginst863 (N1873, N1344);
  not ginst864 (N1874, N1347);
  not ginst865 (N1875, N1350);
  not ginst866 (N1876, N1353);
  not ginst867 (N1877, N1356);
  not ginst868 (N1878, N1359);
  not ginst869 (N1879, N1362);
  not ginst870 (N1880, N1365);
  not ginst871 (N1881, N1368);
  not ginst872 (N1882, N1371);
  not ginst873 (N1883, N1374);
  not ginst874 (N1884, N1377);
  buf ginst875 (N1885, N1199);
  buf ginst876 (N1892, N1194);
  buf ginst877 (N1899, N1199);
  buf ginst878 (N1906, N1194);
  not ginst879 (N1913, N1211);
  buf ginst880 (N1919, N1194);
  and ginst881 (N1926, N44, N1211);
  and ginst882 (N1927, N41, N1211);
  and ginst883 (N1928, N29, N1211);
  and ginst884 (N1929, N26, N1211);
  and ginst885 (N1930, N23, N1211);
  not ginst886 (N1931, N1380);
  not ginst887 (N1932, N1383);
  not ginst888 (N1933, N1386);
  not ginst889 (N1934, N1389);
  not ginst890 (N1935, N1392);
  not ginst891 (N1936, N1395);
  not ginst892 (N1937, N1398);
  not ginst893 (N1938, N1401);
  not ginst894 (N1939, N1404);
  not ginst895 (N1940, N1407);
  not ginst896 (N1941, N1410);
  not ginst897 (N1942, N1413);
  not ginst898 (N1943, N1416);
  not ginst899 (N1944, N1419);
  not ginst900 (N1945, N1422);
  not ginst901 (N1946, N1425);
  not ginst902 (N1947, N1233);
  not ginst903 (N1953, N1244);
  and ginst904 (N1957, N209, N1233);
  and ginst905 (N1958, N216, N1233);
  and ginst906 (N1959, N215, N1233);
  and ginst907 (N1960, N214, N1233);
  and ginst908 (N1961, N213, N1244);
  and ginst909 (N1962, N212, N1244);
  and ginst910 (N1963, N211, N1244);
  not ginst911 (N1965, N1428);
  and ginst912 (N1966, N1222, N636);
  not ginst913 (N1967, N1431);
  not ginst914 (N1968, N1434);
  not ginst915 (N1969, N1437);
  not ginst916 (N1970, N1440);
  not ginst917 (N1971, N1443);
  not ginst918 (N1972, N1446);
  not ginst919 (N1973, N1449);
  not ginst920 (N1974, N1452);
  not ginst921 (N1975, N1455);
  not ginst922 (N1976, N1458);
  not ginst923 (N1977, N1249);
  not ginst924 (N1983, N1256);
  and ginst925 (N1989, N1249, N642);
  and ginst926 (N1990, N1249, N644);
  and ginst927 (N1991, N1249, N651);
  and ginst928 (N1992, N1249, N674);
  and ginst929 (N1993, N1249, N660);
  and ginst930 (N1994, N1256, N666);
  and ginst931 (N1995, N1256, N672);
  and ginst932 (N1996, N1256, N673);
  not ginst933 (N1997, N1263);
  buf ginst934 (N2003, N1194);
  and ginst935 (N2010, N47, N1263);
  and ginst936 (N2011, N35, N1263);
  and ginst937 (N2012, N32, N1263);
  and ginst938 (N2013, N50, N1263);
  and ginst939 (N2014, N66, N1263);
  not ginst940 (N2015, N1461);
  not ginst941 (N2016, N1464);
  not ginst942 (N2017, N1467);
  not ginst943 (N2018, N1470);
  not ginst944 (N2019, N1473);
  not ginst945 (N2020, N1476);
  not ginst946 (N2021, N1479);
  not ginst947 (N2022, N1482);
  not ginst948 (N2023, N1485);
  buf ginst949 (N2024, N1206);
  buf ginst950 (N2031, N1206);
  buf ginst951 (N2038, N1206);
  buf ginst952 (N2045, N1206);
  not ginst953 (N2052, N1270);
  not ginst954 (N2058, N1277);
  and ginst955 (N2064, N1270, N706);
  and ginst956 (N2065, N1270, N708);
  and ginst957 (N2066, N1270, N715);
  and ginst958 (N2067, N1270, N721);
  and ginst959 (N2068, N1270, N727);
  and ginst960 (N2069, N1277, N733);
  and ginst961 (N2070, N1277, N734);
  and ginst962 (N2071, N1277, N742);
  and ginst963 (N2072, N1277, N748);
  and ginst964 (N2073, N1277, N749);
  buf ginst965 (N2074, N1189);
  buf ginst966 (N2081, N1189);
  buf ginst967 (N2086, N1222);
  nand ginst968 (N2107, N1287, N1821);
  nand ginst969 (N2108, N1284, N1822);
  not ginst970 (N2110, N1703);
  nand ginst971 (N2111, N1703, N1832);
  nand ginst972 (N2112, N1308, N1834);
  nand ginst973 (N2113, N1305, N1835);
  not ginst974 (N2114, N1713);
  nand ginst975 (N2115, N1713, N1839);
  not ginst976 (N2117, N1721);
  not ginst977 (N2171, N1758);
  nand ginst978 (N2172, N1758, N1965);
  not ginst979 (N2230, N1708);
  buf ginst980 (N2231, N1537);
  buf ginst981 (N2235, N1551);
  or ginst982 (N2239, N1782, N1783);
  or ginst983 (N2240, N1125, N1783);
  or ginst984 (N2241, N1783, N1793);
  or ginst985 (N2242, N1783, N1794);
  or ginst986 (N2243, N1783, N1795);
  or ginst987 (N2244, N1789, N1796);
  or ginst988 (N2245, N1789, N1797);
  or ginst989 (N2246, N1789, N1798);
  or ginst990 (N2247, N1799, N1811);
  or ginst991 (N2248, N1799, N1812);
  or ginst992 (N2249, N1799, N1813);
  or ginst993 (N2250, N1799, N1814);
  or ginst994 (N2251, N1799, N1815);
  or ginst995 (N2252, N1805, N1816);
  or ginst996 (N2253, N1805, N1817);
  or ginst997 (N2254, N1805, N1818);
  or ginst998 (N2255, N1805, N1819);
  or ginst999 (N2256, N1805, N1820);
  nand ginst1000 (N2257, N2107, N2108);
  not ginst1001 (N2267, N2074);
  nand ginst1002 (N2268, N1299, N2110);
  nand ginst1003 (N2269, N2112, N2113);
  nand ginst1004 (N2274, N1311, N2114);
  not ginst1005 (N2275, N2081);
  and ginst1006 (N2277, N141, N1845);
  and ginst1007 (N2278, N147, N1845);
  and ginst1008 (N2279, N138, N1845);
  and ginst1009 (N2280, N144, N1845);
  and ginst1010 (N2281, N135, N1845);
  and ginst1011 (N2282, N141, N1851);
  and ginst1012 (N2283, N147, N1851);
  and ginst1013 (N2284, N138, N1851);
  and ginst1014 (N2285, N144, N1851);
  and ginst1015 (N2286, N135, N1851);
  not ginst1016 (N2287, N1885);
  not ginst1017 (N2293, N1892);
  and ginst1018 (N2299, N103, N1885);
  and ginst1019 (N2300, N130, N1885);
  and ginst1020 (N2301, N127, N1885);
  and ginst1021 (N2302, N124, N1885);
  and ginst1022 (N2303, N100, N1885);
  and ginst1023 (N2304, N103, N1892);
  and ginst1024 (N2305, N130, N1892);
  and ginst1025 (N2306, N127, N1892);
  and ginst1026 (N2307, N124, N1892);
  and ginst1027 (N2308, N100, N1892);
  not ginst1028 (N2309, N1899);
  not ginst1029 (N2315, N1906);
  and ginst1030 (N2321, N115, N1899);
  and ginst1031 (N2322, N118, N1899);
  and ginst1032 (N2323, N97, N1899);
  and ginst1033 (N2324, N94, N1899);
  and ginst1034 (N2325, N121, N1899);
  and ginst1035 (N2326, N115, N1906);
  and ginst1036 (N2327, N118, N1906);
  and ginst1037 (N2328, N97, N1906);
  and ginst1038 (N2329, N94, N1906);
  and ginst1039 (N2330, N121, N1906);
  not ginst1040 (N2331, N1919);
  and ginst1041 (N2337, N208, N1913);
  and ginst1042 (N2338, N198, N1913);
  and ginst1043 (N2339, N207, N1913);
  and ginst1044 (N2340, N206, N1913);
  and ginst1045 (N2341, N205, N1913);
  and ginst1046 (N2342, N44, N1919);
  and ginst1047 (N2343, N41, N1919);
  and ginst1048 (N2344, N29, N1919);
  and ginst1049 (N2345, N26, N1919);
  and ginst1050 (N2346, N23, N1919);
  or ginst1051 (N2347, N1233, N1947);
  or ginst1052 (N2348, N1947, N1957);
  or ginst1053 (N2349, N1947, N1958);
  or ginst1054 (N2350, N1947, N1959);
  or ginst1055 (N2351, N1947, N1960);
  or ginst1056 (N2352, N1953, N1961);
  or ginst1057 (N2353, N1953, N1962);
  or ginst1058 (N2354, N1953, N1963);
  nand ginst1059 (N2355, N1428, N2171);
  not ginst1060 (N2356, N2086);
  nand ginst1061 (N2357, N1967, N2086);
  and ginst1062 (N2358, N114, N1977);
  and ginst1063 (N2359, N113, N1977);
  and ginst1064 (N2360, N111, N1977);
  and ginst1065 (N2361, N87, N1977);
  and ginst1066 (N2362, N112, N1977);
  and ginst1067 (N2363, N88, N1983);
  and ginst1068 (N2364, N245, N1983);
  and ginst1069 (N2365, N271, N1983);
  and ginst1070 (N2366, N1983, N759);
  and ginst1071 (N2367, N70, N1983);
  not ginst1072 (N2368, N2003);
  and ginst1073 (N2374, N193, N1997);
  and ginst1074 (N2375, N192, N1997);
  and ginst1075 (N2376, N191, N1997);
  and ginst1076 (N2377, N190, N1997);
  and ginst1077 (N2378, N189, N1997);
  and ginst1078 (N2379, N47, N2003);
  and ginst1079 (N2380, N35, N2003);
  and ginst1080 (N2381, N32, N2003);
  and ginst1081 (N2382, N50, N2003);
  and ginst1082 (N2383, N66, N2003);
  not ginst1083 (N2384, N2024);
  not ginst1084 (N2390, N2031);
  and ginst1085 (N2396, N58, N2024);
  and ginst1086 (N2397, N77, N2024);
  and ginst1087 (N2398, N78, N2024);
  and ginst1088 (N2399, N59, N2024);
  and ginst1089 (N2400, N81, N2024);
  and ginst1090 (N2401, N80, N2031);
  and ginst1091 (N2402, N79, N2031);
  and ginst1092 (N2403, N60, N2031);
  and ginst1093 (N2404, N61, N2031);
  and ginst1094 (N2405, N62, N2031);
  not ginst1095 (N2406, N2038);
  not ginst1096 (N2412, N2045);
  and ginst1097 (N2418, N69, N2038);
  and ginst1098 (N2419, N70, N2038);
  buf ginst1099 (N241_BUFF, N241);
  and ginst1100 (N2420, N74, N2038);
  and ginst1101 (N2421, N76, N2038);
  and ginst1102 (N2422, N75, N2038);
  and ginst1103 (N2423, N73, N2045);
  and ginst1104 (N2424, N53, N2045);
  and ginst1105 (N2425, N54, N2045);
  and ginst1106 (N2426, N55, N2045);
  and ginst1107 (N2427, N56, N2045);
  and ginst1108 (N2428, N82, N2052);
  and ginst1109 (N2429, N65, N2052);
  and ginst1110 (N2430, N83, N2052);
  and ginst1111 (N2431, N84, N2052);
  and ginst1112 (N2432, N85, N2052);
  and ginst1113 (N2433, N64, N2058);
  and ginst1114 (N2434, N63, N2058);
  and ginst1115 (N2435, N86, N2058);
  and ginst1116 (N2436, N109, N2058);
  and ginst1117 (N2437, N110, N2058);
  and ginst1118 (N2441, N1119, N2239);
  and ginst1119 (N2442, N1119, N2240);
  and ginst1120 (N2446, N1119, N2241);
  and ginst1121 (N2450, N1119, N2242);
  and ginst1122 (N2454, N1119, N2243);
  and ginst1123 (N2458, N1132, N2244);
  and ginst1124 (N2462, N1141, N2247);
  and ginst1125 (N2466, N1141, N2248);
  and ginst1126 (N2470, N1141, N2249);
  and ginst1127 (N2474, N1141, N2250);
  and ginst1128 (N2478, N1141, N2251);
  and ginst1129 (N2482, N1154, N2252);
  and ginst1130 (N2488, N1154, N2253);
  and ginst1131 (N2496, N1154, N2254);
  and ginst1132 (N2502, N1154, N2255);
  and ginst1133 (N2508, N1154, N2256);
  nand ginst1134 (N2523, N2111, N2268);
  nand ginst1135 (N2533, N2115, N2274);
  not ginst1136 (N2537, N2235);
  or ginst1137 (N2538, N1858, N2278);
  or ginst1138 (N2542, N1859, N2279);
  or ginst1139 (N2546, N1860, N2280);
  or ginst1140 (N2550, N1861, N2281);
  or ginst1141 (N2554, N1863, N2283);
  or ginst1142 (N2561, N1864, N2284);
  or ginst1143 (N2567, N1865, N2285);
  or ginst1144 (N2573, N1866, N2286);
  or ginst1145 (N2604, N1927, N2338);
  or ginst1146 (N2607, N1928, N2339);
  or ginst1147 (N2611, N1929, N2340);
  or ginst1148 (N2615, N1930, N2341);
  and ginst1149 (N2619, N1227, N2348);
  and ginst1150 (N2626, N1227, N2349);
  and ginst1151 (N2632, N1227, N2350);
  and ginst1152 (N2638, N1227, N2351);
  and ginst1153 (N2644, N1240, N2352);
  nand ginst1154 (N2650, N2172, N2355);
  nand ginst1155 (N2653, N1431, N2356);
  or ginst1156 (N2654, N1990, N2359);
  or ginst1157 (N2658, N1991, N2360);
  or ginst1158 (N2662, N1992, N2361);
  or ginst1159 (N2666, N1993, N2362);
  or ginst1160 (N2670, N1994, N2363);
  or ginst1161 (N2674, N1256, N2366);
  or ginst1162 (N2680, N1256, N2367);
  or ginst1163 (N2688, N2010, N2374);
  or ginst1164 (N2692, N2011, N2375);
  or ginst1165 (N2696, N2012, N2376);
  or ginst1166 (N2700, N2013, N2377);
  or ginst1167 (N2704, N2014, N2378);
  and ginst1168 (N2728, N1227, N2347);
  or ginst1169 (N2729, N2065, N2429);
  or ginst1170 (N2733, N2066, N2430);
  or ginst1171 (N2737, N2067, N2431);
  or ginst1172 (N2741, N2068, N2432);
  or ginst1173 (N2745, N2069, N2433);
  or ginst1174 (N2749, N2070, N2434);
  or ginst1175 (N2753, N2071, N2435);
  or ginst1176 (N2757, N2072, N2436);
  or ginst1177 (N2761, N2073, N2437);
  not ginst1178 (N2765, N2231);
  and ginst1179 (N2766, N1240, N2354);
  and ginst1180 (N2769, N1240, N2353);
  and ginst1181 (N2772, N1132, N2246);
  and ginst1182 (N2775, N1132, N2245);
  or ginst1183 (N2778, N1862, N2282);
  or ginst1184 (N2781, N1989, N2358);
  or ginst1185 (N2784, N1996, N2365);
  or ginst1186 (N2787, N1995, N2364);
  or ginst1187 (N2790, N1926, N2337);
  or ginst1188 (N2793, N1857, N2277);
  or ginst1189 (N2796, N2064, N2428);
  and ginst1190 (N2866, N1537, N2257);
  and ginst1191 (N2867, N1537, N2257);
  and ginst1192 (N2868, N1537, N2257);
  and ginst1193 (N2869, N1537, N2257);
  and ginst1194 (N2878, N1551, N2269);
  and ginst1195 (N2913, N204, N2287);
  and ginst1196 (N2914, N203, N2287);
  and ginst1197 (N2915, N202, N2287);
  and ginst1198 (N2916, N201, N2287);
  and ginst1199 (N2917, N200, N2287);
  and ginst1200 (N2918, N235, N2293);
  and ginst1201 (N2919, N234, N2293);
  and ginst1202 (N2920, N233, N2293);
  and ginst1203 (N2921, N232, N2293);
  and ginst1204 (N2922, N231, N2293);
  and ginst1205 (N2923, N197, N2309);
  and ginst1206 (N2924, N187, N2309);
  and ginst1207 (N2925, N196, N2309);
  and ginst1208 (N2926, N195, N2309);
  and ginst1209 (N2927, N194, N2309);
  and ginst1210 (N2928, N227, N2315);
  and ginst1211 (N2929, N217, N2315);
  and ginst1212 (N2930, N226, N2315);
  and ginst1213 (N2931, N225, N2315);
  and ginst1214 (N2932, N224, N2315);
  and ginst1215 (N2933, N239, N2331);
  and ginst1216 (N2934, N229, N2331);
  and ginst1217 (N2935, N238, N2331);
  and ginst1218 (N2936, N237, N2331);
  and ginst1219 (N2937, N236, N2331);
  nand ginst1220 (N2988, N2357, N2653);
  and ginst1221 (N3005, N223, N2368);
  and ginst1222 (N3006, N222, N2368);
  and ginst1223 (N3007, N221, N2368);
  and ginst1224 (N3008, N220, N2368);
  and ginst1225 (N3009, N219, N2368);
  and ginst1226 (N3020, N2384, N812);
  and ginst1227 (N3021, N2384, N814);
  and ginst1228 (N3022, N2384, N821);
  and ginst1229 (N3023, N2384, N827);
  and ginst1230 (N3024, N2384, N833);
  and ginst1231 (N3025, N2390, N839);
  and ginst1232 (N3026, N2390, N845);
  and ginst1233 (N3027, N2390, N853);
  and ginst1234 (N3028, N2390, N859);
  and ginst1235 (N3029, N2390, N865);
  and ginst1236 (N3032, N2406, N758);
  and ginst1237 (N3033, N2406, N759);
  and ginst1238 (N3034, N2406, N762);
  and ginst1239 (N3035, N2406, N768);
  and ginst1240 (N3036, N2406, N774);
  and ginst1241 (N3037, N2412, N780);
  and ginst1242 (N3038, N2412, N786);
  and ginst1243 (N3039, N2412, N794);
  and ginst1244 (N3040, N2412, N800);
  and ginst1245 (N3041, N2412, N806);
  buf ginst1246 (N3061, N2257);
  buf ginst1247 (N3064, N2257);
  buf ginst1248 (N3067, N2269);
  buf ginst1249 (N3070, N2269);
  not ginst1250 (N3073, N2728);
  not ginst1251 (N3080, N2441);
  and ginst1252 (N3096, N2644, N666);
  and ginst1253 (N3097, N2638, N660);
  and ginst1254 (N3101, N1189, N2632);
  and ginst1255 (N3107, N2626, N651);
  and ginst1256 (N3114, N2619, N644);
  and ginst1257 (N3122, N2257, N2523);
  or ginst1258 (N3126, N1167, N2866);
  and ginst1259 (N3130, N2257, N2523);
  or ginst1260 (N3131, N1167, N2869);
  and ginst1261 (N3134, N2257, N2523);
  not ginst1262 (N3135, N2533);
  and ginst1263 (N3136, N2644, N666);
  and ginst1264 (N3137, N2638, N660);
  and ginst1265 (N3140, N1189, N2632);
  and ginst1266 (N3144, N2626, N651);
  and ginst1267 (N3149, N2619, N644);
  and ginst1268 (N3155, N2269, N2533);
  or ginst1269 (N3159, N1174, N2878);
  not ginst1270 (N3167, N2778);
  and ginst1271 (N3168, N2508, N609);
  and ginst1272 (N3169, N2502, N604);
  and ginst1273 (N3173, N2496, N742);
  and ginst1274 (N3178, N2488, N734);
  and ginst1275 (N3184, N2482, N599);
  and ginst1276 (N3185, N2573, N727);
  and ginst1277 (N3189, N2567, N721);
  and ginst1278 (N3195, N2561, N715);
  and ginst1279 (N3202, N2554, N708);
  and ginst1280 (N3210, N2508, N609);
  and ginst1281 (N3211, N2502, N604);
  and ginst1282 (N3215, N2496, N742);
  and ginst1283 (N3221, N2488, N734);
  and ginst1284 (N3228, N2482, N599);
  and ginst1285 (N3229, N2573, N727);
  and ginst1286 (N3232, N2567, N721);
  and ginst1287 (N3236, N2561, N715);
  and ginst1288 (N3241, N2554, N708);
  or ginst1289 (N3247, N2299, N2913);
  or ginst1290 (N3251, N2300, N2914);
  or ginst1291 (N3255, N2301, N2915);
  or ginst1292 (N3259, N2302, N2916);
  or ginst1293 (N3263, N2303, N2917);
  or ginst1294 (N3267, N2304, N2918);
  or ginst1295 (N3273, N2305, N2919);
  or ginst1296 (N3281, N2306, N2920);
  or ginst1297 (N3287, N2307, N2921);
  or ginst1298 (N3293, N2308, N2922);
  or ginst1299 (N3299, N2322, N2924);
  or ginst1300 (N3303, N2323, N2925);
  or ginst1301 (N3307, N2324, N2926);
  or ginst1302 (N3311, N2325, N2927);
  or ginst1303 (N3315, N2327, N2929);
  or ginst1304 (N3322, N2328, N2930);
  or ginst1305 (N3328, N2329, N2931);
  or ginst1306 (N3334, N2330, N2932);
  or ginst1307 (N3340, N2343, N2934);
  or ginst1308 (N3343, N2344, N2935);
  or ginst1309 (N3349, N2345, N2936);
  or ginst1310 (N3355, N2346, N2937);
  and ginst1311 (N3361, N2478, N2761);
  and ginst1312 (N3362, N2474, N2757);
  and ginst1313 (N3363, N2470, N2753);
  and ginst1314 (N3364, N2466, N2749);
  and ginst1315 (N3365, N2462, N2745);
  and ginst1316 (N3366, N2550, N2741);
  and ginst1317 (N3367, N2546, N2737);
  and ginst1318 (N3368, N2542, N2733);
  and ginst1319 (N3369, N2538, N2729);
  and ginst1320 (N3370, N2458, N2670);
  and ginst1321 (N3371, N2454, N2666);
  and ginst1322 (N3372, N2450, N2662);
  and ginst1323 (N3373, N2446, N2658);
  and ginst1324 (N3374, N2442, N2654);
  and ginst1325 (N3375, N2650, N2988);
  and ginst1326 (N3379, N1966, N2650);
  not ginst1327 (N3380, N2781);
  and ginst1328 (N3381, N2604, N695);
  or ginst1329 (N3384, N2379, N3005);
  or ginst1330 (N3390, N2380, N3006);
  or ginst1331 (N3398, N2381, N3007);
  or ginst1332 (N3404, N2382, N3008);
  or ginst1333 (N3410, N2383, N3009);
  or ginst1334 (N3416, N2397, N3021);
  or ginst1335 (N3420, N2398, N3022);
  or ginst1336 (N3424, N2399, N3023);
  or ginst1337 (N3428, N2400, N3024);
  or ginst1338 (N3432, N2401, N3025);
  or ginst1339 (N3436, N2402, N3026);
  or ginst1340 (N3440, N2403, N3027);
  or ginst1341 (N3444, N2404, N3028);
  or ginst1342 (N3448, N2405, N3029);
  not ginst1343 (N3452, N2790);
  not ginst1344 (N3453, N2793);
  or ginst1345 (N3454, N2420, N3034);
  or ginst1346 (N3458, N2421, N3035);
  or ginst1347 (N3462, N2422, N3036);
  or ginst1348 (N3466, N2423, N3037);
  or ginst1349 (N3470, N2424, N3038);
  or ginst1350 (N3474, N2425, N3039);
  or ginst1351 (N3478, N2426, N3040);
  or ginst1352 (N3482, N2427, N3041);
  not ginst1353 (N3486, N2796);
  buf ginst1354 (N3487, N2644);
  buf ginst1355 (N3490, N2638);
  buf ginst1356 (N3493, N2632);
  buf ginst1357 (N3496, N2626);
  buf ginst1358 (N3499, N2619);
  buf ginst1359 (N3502, N2523);
  nor ginst1360 (N3507, N1167, N2868);
  buf ginst1361 (N3510, N2523);
  nor ginst1362 (N3515, N2619, N644);
  buf ginst1363 (N3518, N2644);
  buf ginst1364 (N3521, N2638);
  buf ginst1365 (N3524, N2632);
  buf ginst1366 (N3527, N2626);
  buf ginst1367 (N3530, N2619);
  buf ginst1368 (N3535, N2619);
  buf ginst1369 (N3539, N2632);
  buf ginst1370 (N3542, N2626);
  buf ginst1371 (N3545, N2644);
  buf ginst1372 (N3548, N2638);
  not ginst1373 (N3551, N2766);
  not ginst1374 (N3552, N2769);
  buf ginst1375 (N3553, N2442);
  buf ginst1376 (N3557, N2450);
  buf ginst1377 (N3560, N2446);
  buf ginst1378 (N3563, N2458);
  buf ginst1379 (N3566, N2454);
  not ginst1380 (N3569, N2772);
  not ginst1381 (N3570, N2775);
  buf ginst1382 (N3571, N2554);
  buf ginst1383 (N3574, N2567);
  buf ginst1384 (N3577, N2561);
  buf ginst1385 (N3580, N2482);
  buf ginst1386 (N3583, N2573);
  buf ginst1387 (N3586, N2496);
  buf ginst1388 (N3589, N2488);
  buf ginst1389 (N3592, N2508);
  buf ginst1390 (N3595, N2502);
  buf ginst1391 (N3598, N2508);
  buf ginst1392 (N3601, N2502);
  buf ginst1393 (N3604, N2496);
  buf ginst1394 (N3607, N2482);
  buf ginst1395 (N3610, N2573);
  buf ginst1396 (N3613, N2567);
  buf ginst1397 (N3616, N2561);
  buf ginst1398 (N3619, N2488);
  buf ginst1399 (N3622, N2554);
  nor ginst1400 (N3625, N2488, N734);
  nor ginst1401 (N3628, N2554, N708);
  buf ginst1402 (N3631, N2508);
  buf ginst1403 (N3634, N2502);
  buf ginst1404 (N3637, N2496);
  buf ginst1405 (N3640, N2488);
  buf ginst1406 (N3643, N2482);
  buf ginst1407 (N3646, N2573);
  buf ginst1408 (N3649, N2567);
  buf ginst1409 (N3652, N2561);
  buf ginst1410 (N3655, N2554);
  nor ginst1411 (N3658, N2488, N734);
  buf ginst1412 (N3661, N2674);
  buf ginst1413 (N3664, N2674);
  buf ginst1414 (N3667, N2761);
  buf ginst1415 (N3670, N2478);
  buf ginst1416 (N3673, N2757);
  buf ginst1417 (N3676, N2474);
  buf ginst1418 (N3679, N2753);
  buf ginst1419 (N3682, N2470);
  buf ginst1420 (N3685, N2745);
  buf ginst1421 (N3688, N2462);
  buf ginst1422 (N3691, N2741);
  buf ginst1423 (N3694, N2550);
  buf ginst1424 (N3697, N2737);
  buf ginst1425 (N3700, N2546);
  buf ginst1426 (N3703, N2733);
  buf ginst1427 (N3706, N2542);
  buf ginst1428 (N3709, N2749);
  buf ginst1429 (N3712, N2466);
  buf ginst1430 (N3715, N2729);
  buf ginst1431 (N3718, N2538);
  buf ginst1432 (N3721, N2704);
  buf ginst1433 (N3724, N2700);
  buf ginst1434 (N3727, N2696);
  buf ginst1435 (N3730, N2688);
  buf ginst1436 (N3733, N2692);
  buf ginst1437 (N3736, N2670);
  buf ginst1438 (N3739, N2458);
  buf ginst1439 (N3742, N2666);
  buf ginst1440 (N3745, N2454);
  buf ginst1441 (N3748, N2662);
  buf ginst1442 (N3751, N2450);
  buf ginst1443 (N3754, N2658);
  buf ginst1444 (N3757, N2446);
  buf ginst1445 (N3760, N2654);
  buf ginst1446 (N3763, N2442);
  buf ginst1447 (N3766, N2654);
  buf ginst1448 (N3769, N2662);
  buf ginst1449 (N3772, N2658);
  buf ginst1450 (N3775, N2670);
  buf ginst1451 (N3778, N2666);
  not ginst1452 (N3781, N2784);
  not ginst1453 (N3782, N2787);
  or ginst1454 (N3783, N2326, N2928);
  or ginst1455 (N3786, N2342, N2933);
  or ginst1456 (N3789, N2321, N2923);
  buf ginst1457 (N3792, N2688);
  buf ginst1458 (N3795, N2696);
  buf ginst1459 (N3798, N2692);
  buf ginst1460 (N3801, N2704);
  buf ginst1461 (N3804, N2700);
  buf ginst1462 (N3807, N2604);
  buf ginst1463 (N3810, N2611);
  buf ginst1464 (N3813, N2607);
  buf ginst1465 (N3816, N2615);
  buf ginst1466 (N3819, N2538);
  buf ginst1467 (N3822, N2546);
  buf ginst1468 (N3825, N2542);
  buf ginst1469 (N3828, N2462);
  buf ginst1470 (N3831, N2550);
  buf ginst1471 (N3834, N2470);
  buf ginst1472 (N3837, N2466);
  buf ginst1473 (N3840, N2478);
  buf ginst1474 (N3843, N2474);
  buf ginst1475 (N3846, N2615);
  buf ginst1476 (N3849, N2611);
  buf ginst1477 (N3852, N2607);
  buf ginst1478 (N3855, N2680);
  buf ginst1479 (N3858, N2729);
  buf ginst1480 (N3861, N2737);
  buf ginst1481 (N3864, N2733);
  buf ginst1482 (N3867, N2745);
  buf ginst1483 (N387, N1);
  buf ginst1484 (N3870, N2741);
  buf ginst1485 (N3873, N2753);
  buf ginst1486 (N3876, N2749);
  buf ginst1487 (N3879, N2761);
  buf ginst1488 (N388, N1);
  buf ginst1489 (N3882, N2757);
  or ginst1490 (N3885, N2419, N3033);
  or ginst1491 (N3888, N2418, N3032);
  or ginst1492 (N3891, N2396, N3020);
  nand ginst1493 (N3953, N2117, N3067);
  not ginst1494 (N3954, N3067);
  nand ginst1495 (N3955, N2537, N3070);
  not ginst1496 (N3956, N3070);
  not ginst1497 (N3958, N3073);
  not ginst1498 (N3964, N3080);
  or ginst1499 (N4193, N1649, N3379);
  or ginst1500 (N4303, N1167, N2867, N3130);
  not ginst1501 (N4308, N3061);
  not ginst1502 (N4313, N3064);
  nand ginst1503 (N4326, N2769, N3551);
  nand ginst1504 (N4327, N2766, N3552);
  nand ginst1505 (N4333, N2775, N3569);
  nand ginst1506 (N4334, N2772, N3570);
  nand ginst1507 (N4411, N2787, N3781);
  nand ginst1508 (N4412, N2784, N3782);
  nand ginst1509 (N4463, N1828, N3487);
  not ginst1510 (N4464, N3487);
  nand ginst1511 (N4465, N1829, N3490);
  not ginst1512 (N4466, N3490);
  nand ginst1513 (N4467, N2267, N3493);
  not ginst1514 (N4468, N3493);
  nand ginst1515 (N4469, N1830, N3496);
  not ginst1516 (N4470, N3496);
  nand ginst1517 (N4471, N1833, N3499);
  not ginst1518 (N4472, N3499);
  not ginst1519 (N4473, N3122);
  not ginst1520 (N4474, N3126);
  nand ginst1521 (N4475, N1840, N3518);
  not ginst1522 (N4476, N3518);
  nand ginst1523 (N4477, N1841, N3521);
  not ginst1524 (N4478, N3521);
  nand ginst1525 (N4479, N2275, N3524);
  not ginst1526 (N4480, N3524);
  nand ginst1527 (N4481, N1842, N3527);
  not ginst1528 (N4482, N3527);
  nand ginst1529 (N4483, N1843, N3530);
  not ginst1530 (N4484, N3530);
  not ginst1531 (N4485, N3155);
  not ginst1532 (N4486, N3159);
  nand ginst1533 (N4487, N1721, N3954);
  nand ginst1534 (N4488, N2235, N3956);
  not ginst1535 (N4489, N3535);
  nand ginst1536 (N4490, N3535, N3958);
  not ginst1537 (N4491, N3539);
  not ginst1538 (N4492, N3542);
  not ginst1539 (N4493, N3545);
  not ginst1540 (N4494, N3548);
  not ginst1541 (N4495, N3553);
  nand ginst1542 (N4496, N3553, N3964);
  not ginst1543 (N4497, N3557);
  not ginst1544 (N4498, N3560);
  not ginst1545 (N4499, N3563);
  not ginst1546 (N4500, N3566);
  not ginst1547 (N4501, N3571);
  nand ginst1548 (N4502, N3167, N3571);
  not ginst1549 (N4503, N3574);
  not ginst1550 (N4504, N3577);
  not ginst1551 (N4505, N3580);
  not ginst1552 (N4506, N3583);
  nand ginst1553 (N4507, N1867, N3598);
  not ginst1554 (N4508, N3598);
  nand ginst1555 (N4509, N1868, N3601);
  not ginst1556 (N4510, N3601);
  nand ginst1557 (N4511, N1869, N3604);
  not ginst1558 (N4512, N3604);
  nand ginst1559 (N4513, N1870, N3607);
  not ginst1560 (N4514, N3607);
  nand ginst1561 (N4515, N1871, N3610);
  not ginst1562 (N4516, N3610);
  nand ginst1563 (N4517, N1872, N3613);
  not ginst1564 (N4518, N3613);
  nand ginst1565 (N4519, N1873, N3616);
  not ginst1566 (N4520, N3616);
  nand ginst1567 (N4521, N1874, N3619);
  not ginst1568 (N4522, N3619);
  nand ginst1569 (N4523, N1875, N3622);
  not ginst1570 (N4524, N3622);
  nand ginst1571 (N4525, N1876, N3631);
  not ginst1572 (N4526, N3631);
  nand ginst1573 (N4527, N1877, N3634);
  not ginst1574 (N4528, N3634);
  nand ginst1575 (N4529, N1878, N3637);
  not ginst1576 (N4530, N3637);
  nand ginst1577 (N4531, N1879, N3640);
  not ginst1578 (N4532, N3640);
  nand ginst1579 (N4533, N1880, N3643);
  not ginst1580 (N4534, N3643);
  nand ginst1581 (N4535, N1881, N3646);
  not ginst1582 (N4536, N3646);
  nand ginst1583 (N4537, N1882, N3649);
  not ginst1584 (N4538, N3649);
  nand ginst1585 (N4539, N1883, N3652);
  not ginst1586 (N4540, N3652);
  nand ginst1587 (N4541, N1884, N3655);
  not ginst1588 (N4542, N3655);
  not ginst1589 (N4543, N3658);
  and ginst1590 (N4544, N3293, N806);
  and ginst1591 (N4545, N3287, N800);
  and ginst1592 (N4549, N3281, N794);
  and ginst1593 (N4555, N3273, N786);
  and ginst1594 (N4562, N3267, N780);
  and ginst1595 (N4563, N3355, N774);
  and ginst1596 (N4566, N3349, N768);
  and ginst1597 (N4570, N3343, N762);
  not ginst1598 (N4575, N3661);
  and ginst1599 (N4576, N3293, N806);
  and ginst1600 (N4577, N3287, N800);
  and ginst1601 (N4581, N3281, N794);
  and ginst1602 (N4586, N3273, N786);
  and ginst1603 (N4592, N3267, N780);
  and ginst1604 (N4593, N3355, N774);
  and ginst1605 (N4597, N3349, N768);
  and ginst1606 (N4603, N3343, N762);
  not ginst1607 (N4610, N3664);
  not ginst1608 (N4611, N3667);
  not ginst1609 (N4612, N3670);
  not ginst1610 (N4613, N3673);
  not ginst1611 (N4614, N3676);
  not ginst1612 (N4615, N3679);
  not ginst1613 (N4616, N3682);
  not ginst1614 (N4617, N3685);
  not ginst1615 (N4618, N3688);
  not ginst1616 (N4619, N3691);
  not ginst1617 (N4620, N3694);
  not ginst1618 (N4621, N3697);
  not ginst1619 (N4622, N3700);
  not ginst1620 (N4623, N3703);
  not ginst1621 (N4624, N3706);
  not ginst1622 (N4625, N3709);
  not ginst1623 (N4626, N3712);
  not ginst1624 (N4627, N3715);
  not ginst1625 (N4628, N3718);
  not ginst1626 (N4629, N3721);
  and ginst1627 (N4630, N2704, N3448);
  not ginst1628 (N4631, N3724);
  and ginst1629 (N4632, N2700, N3444);
  not ginst1630 (N4633, N3727);
  and ginst1631 (N4634, N2696, N3440);
  and ginst1632 (N4635, N2692, N3436);
  not ginst1633 (N4636, N3730);
  and ginst1634 (N4637, N2688, N3432);
  and ginst1635 (N4638, N3311, N3428);
  and ginst1636 (N4639, N3307, N3424);
  and ginst1637 (N4640, N3303, N3420);
  and ginst1638 (N4641, N3299, N3416);
  not ginst1639 (N4642, N3733);
  not ginst1640 (N4643, N3736);
  not ginst1641 (N4644, N3739);
  not ginst1642 (N4645, N3742);
  not ginst1643 (N4646, N3745);
  not ginst1644 (N4647, N3748);
  not ginst1645 (N4648, N3751);
  not ginst1646 (N4649, N3754);
  not ginst1647 (N4650, N3757);
  not ginst1648 (N4651, N3760);
  not ginst1649 (N4652, N3763);
  not ginst1650 (N4653, N3375);
  and ginst1651 (N4656, N3410, N865);
  and ginst1652 (N4657, N3404, N859);
  and ginst1653 (N4661, N3398, N853);
  and ginst1654 (N4667, N3390, N845);
  not ginst1655 (N467, N57);
  and ginst1656 (N4674, N3384, N839);
  and ginst1657 (N4675, N3334, N833);
  and ginst1658 (N4678, N3328, N827);
  and ginst1659 (N4682, N3322, N821);
  and ginst1660 (N4687, N3315, N814);
  and ginst1661 (N469, N133, N134);
  not ginst1662 (N4693, N3766);
  nand ginst1663 (N4694, N3380, N3766);
  not ginst1664 (N4695, N3769);
  not ginst1665 (N4696, N3772);
  not ginst1666 (N4697, N3775);
  not ginst1667 (N4698, N3778);
  not ginst1668 (N4699, N3783);
  not ginst1669 (N4700, N3786);
  and ginst1670 (N4701, N3410, N865);
  and ginst1671 (N4702, N3404, N859);
  and ginst1672 (N4706, N3398, N853);
  and ginst1673 (N4711, N3390, N845);
  and ginst1674 (N4717, N3384, N839);
  and ginst1675 (N4718, N3334, N833);
  and ginst1676 (N4722, N3328, N827);
  and ginst1677 (N4728, N3322, N821);
  and ginst1678 (N4735, N3315, N814);
  not ginst1679 (N4743, N3789);
  not ginst1680 (N4744, N3792);
  not ginst1681 (N4745, N3807);
  nand ginst1682 (N4746, N3452, N3807);
  not ginst1683 (N4747, N3810);
  not ginst1684 (N4748, N3813);
  not ginst1685 (N4749, N3816);
  not ginst1686 (N4750, N3819);
  nand ginst1687 (N4751, N3453, N3819);
  not ginst1688 (N4752, N3822);
  not ginst1689 (N4753, N3825);
  not ginst1690 (N4754, N3828);
  not ginst1691 (N4755, N3831);
  and ginst1692 (N4756, N3263, N3482);
  and ginst1693 (N4757, N3259, N3478);
  and ginst1694 (N4758, N3255, N3474);
  and ginst1695 (N4759, N3251, N3470);
  and ginst1696 (N4760, N3247, N3466);
  not ginst1697 (N4761, N3846);
  and ginst1698 (N4762, N2615, N3462);
  not ginst1699 (N4763, N3849);
  and ginst1700 (N4764, N2611, N3458);
  not ginst1701 (N4765, N3852);
  and ginst1702 (N4766, N2607, N3454);
  and ginst1703 (N4767, N2680, N3381);
  not ginst1704 (N4768, N3855);
  and ginst1705 (N4769, N3340, N695);
  not ginst1706 (N4775, N3858);
  nand ginst1707 (N4776, N3486, N3858);
  not ginst1708 (N4777, N3861);
  not ginst1709 (N4778, N3864);
  not ginst1710 (N4779, N3867);
  buf ginst1711 (N478, N248);
  not ginst1712 (N4780, N3870);
  not ginst1713 (N4781, N3885);
  not ginst1714 (N4782, N3888);
  not ginst1715 (N4783, N3891);
  or ginst1716 (N4784, N3131, N3134);
  not ginst1717 (N4789, N3502);
  not ginst1718 (N4790, N3131);
  not ginst1719 (N4793, N3507);
  not ginst1720 (N4794, N3510);
  not ginst1721 (N4795, N3515);
  buf ginst1722 (N4796, N3114);
  not ginst1723 (N4799, N3586);
  not ginst1724 (N4800, N3589);
  not ginst1725 (N4801, N3592);
  not ginst1726 (N4802, N3595);
  nand ginst1727 (N4803, N4326, N4327);
  nand ginst1728 (N4806, N4333, N4334);
  not ginst1729 (N4809, N3625);
  buf ginst1730 (N4810, N3178);
  not ginst1731 (N4813, N3628);
  buf ginst1732 (N4814, N3202);
  buf ginst1733 (N4817, N3221);
  buf ginst1734 (N482, N254);
  buf ginst1735 (N4820, N3293);
  buf ginst1736 (N4823, N3287);
  buf ginst1737 (N4826, N3281);
  buf ginst1738 (N4829, N3273);
  buf ginst1739 (N4832, N3267);
  buf ginst1740 (N4835, N3355);
  buf ginst1741 (N4838, N3349);
  buf ginst1742 (N484, N257);
  buf ginst1743 (N4841, N3343);
  nor ginst1744 (N4844, N3273, N786);
  buf ginst1745 (N4847, N3293);
  buf ginst1746 (N4850, N3287);
  buf ginst1747 (N4853, N3281);
  buf ginst1748 (N4856, N3267);
  buf ginst1749 (N4859, N3355);
  buf ginst1750 (N486, N260);
  buf ginst1751 (N4862, N3349);
  buf ginst1752 (N4865, N3343);
  buf ginst1753 (N4868, N3273);
  nor ginst1754 (N4871, N3273, N786);
  buf ginst1755 (N4874, N3448);
  buf ginst1756 (N4877, N3444);
  buf ginst1757 (N4880, N3440);
  buf ginst1758 (N4883, N3432);
  buf ginst1759 (N4886, N3428);
  buf ginst1760 (N4889, N3311);
  buf ginst1761 (N489, N263);
  buf ginst1762 (N4892, N3424);
  buf ginst1763 (N4895, N3307);
  buf ginst1764 (N4898, N3420);
  buf ginst1765 (N4901, N3303);
  buf ginst1766 (N4904, N3436);
  buf ginst1767 (N4907, N3416);
  buf ginst1768 (N4910, N3299);
  buf ginst1769 (N4913, N3410);
  buf ginst1770 (N4916, N3404);
  buf ginst1771 (N4919, N3398);
  buf ginst1772 (N492, N267);
  buf ginst1773 (N4922, N3390);
  buf ginst1774 (N4925, N3384);
  buf ginst1775 (N4928, N3334);
  buf ginst1776 (N4931, N3328);
  buf ginst1777 (N4934, N3322);
  buf ginst1778 (N4937, N3315);
  and ginst1779 (N494, N162, N172, N188, N199);
  nor ginst1780 (N4940, N3390, N845);
  buf ginst1781 (N4943, N3315);
  buf ginst1782 (N4946, N3328);
  buf ginst1783 (N4949, N3322);
  buf ginst1784 (N4952, N3384);
  buf ginst1785 (N4955, N3334);
  buf ginst1786 (N4958, N3398);
  buf ginst1787 (N4961, N3390);
  buf ginst1788 (N4964, N3410);
  buf ginst1789 (N4967, N3404);
  buf ginst1790 (N4970, N3340);
  buf ginst1791 (N4973, N3349);
  buf ginst1792 (N4976, N3343);
  buf ginst1793 (N4979, N3267);
  buf ginst1794 (N4982, N3355);
  buf ginst1795 (N4985, N3281);
  buf ginst1796 (N4988, N3273);
  buf ginst1797 (N4991, N3293);
  buf ginst1798 (N4994, N3287);
  nand ginst1799 (N4997, N4411, N4412);
  buf ginst1800 (N5000, N3410);
  buf ginst1801 (N5003, N3404);
  buf ginst1802 (N5006, N3398);
  buf ginst1803 (N5009, N3384);
  buf ginst1804 (N501, N274);
  buf ginst1805 (N5012, N3334);
  buf ginst1806 (N5015, N3328);
  buf ginst1807 (N5018, N3322);
  buf ginst1808 (N5021, N3390);
  buf ginst1809 (N5024, N3315);
  nor ginst1810 (N5027, N3390, N845);
  nor ginst1811 (N5030, N3315, N814);
  buf ginst1812 (N5033, N3299);
  buf ginst1813 (N5036, N3307);
  buf ginst1814 (N5039, N3303);
  buf ginst1815 (N5042, N3311);
  not ginst1816 (N5045, N3795);
  not ginst1817 (N5046, N3798);
  not ginst1818 (N5047, N3801);
  not ginst1819 (N5048, N3804);
  buf ginst1820 (N5049, N3247);
  buf ginst1821 (N505, N280);
  buf ginst1822 (N5052, N3255);
  buf ginst1823 (N5055, N3251);
  buf ginst1824 (N5058, N3263);
  buf ginst1825 (N5061, N3259);
  not ginst1826 (N5064, N3834);
  not ginst1827 (N5065, N3837);
  not ginst1828 (N5066, N3840);
  not ginst1829 (N5067, N3843);
  buf ginst1830 (N5068, N3482);
  buf ginst1831 (N507, N283);
  buf ginst1832 (N5071, N3263);
  buf ginst1833 (N5074, N3478);
  buf ginst1834 (N5077, N3259);
  buf ginst1835 (N5080, N3474);
  buf ginst1836 (N5083, N3255);
  buf ginst1837 (N5086, N3466);
  buf ginst1838 (N5089, N3247);
  buf ginst1839 (N509, N286);
  buf ginst1840 (N5092, N3462);
  buf ginst1841 (N5095, N3458);
  buf ginst1842 (N5098, N3454);
  buf ginst1843 (N5101, N3470);
  buf ginst1844 (N5104, N3251);
  buf ginst1845 (N5107, N3381);
  buf ginst1846 (N511, N289);
  not ginst1847 (N5110, N3873);
  not ginst1848 (N5111, N3876);
  not ginst1849 (N5112, N3879);
  not ginst1850 (N5113, N3882);
  buf ginst1851 (N5114, N3458);
  buf ginst1852 (N5117, N3454);
  buf ginst1853 (N5120, N3466);
  buf ginst1854 (N5123, N3462);
  buf ginst1855 (N5126, N3474);
  buf ginst1856 (N5129, N3470);
  buf ginst1857 (N513, N293);
  buf ginst1858 (N5132, N3482);
  buf ginst1859 (N5135, N3478);
  buf ginst1860 (N5138, N3416);
  buf ginst1861 (N5141, N3424);
  buf ginst1862 (N5144, N3420);
  buf ginst1863 (N5147, N3432);
  buf ginst1864 (N515, N296);
  buf ginst1865 (N5150, N3428);
  buf ginst1866 (N5153, N3440);
  buf ginst1867 (N5156, N3436);
  buf ginst1868 (N5159, N3448);
  buf ginst1869 (N5162, N3444);
  nand ginst1870 (N5165, N4485, N4486);
  nand ginst1871 (N5166, N4473, N4474);
  nand ginst1872 (N5167, N1290, N4464);
  nand ginst1873 (N5168, N1293, N4466);
  nand ginst1874 (N5169, N2074, N4468);
  buf ginst1875 (N517, N299);
  nand ginst1876 (N5170, N1296, N4470);
  nand ginst1877 (N5171, N1302, N4472);
  nand ginst1878 (N5172, N1314, N4476);
  nand ginst1879 (N5173, N1317, N4478);
  nand ginst1880 (N5174, N2081, N4480);
  nand ginst1881 (N5175, N1320, N4482);
  nand ginst1882 (N5176, N1323, N4484);
  nand ginst1883 (N5177, N3953, N4487);
  nand ginst1884 (N5178, N3955, N4488);
  nand ginst1885 (N5179, N3073, N4489);
  nand ginst1886 (N5180, N3542, N4491);
  nand ginst1887 (N5181, N3539, N4492);
  nand ginst1888 (N5182, N3548, N4493);
  nand ginst1889 (N5183, N3545, N4494);
  nand ginst1890 (N5184, N3080, N4495);
  nand ginst1891 (N5185, N3560, N4497);
  nand ginst1892 (N5186, N3557, N4498);
  nand ginst1893 (N5187, N3566, N4499);
  nand ginst1894 (N5188, N3563, N4500);
  nand ginst1895 (N5189, N2778, N4501);
  buf ginst1896 (N519, N303);
  nand ginst1897 (N5190, N3577, N4503);
  nand ginst1898 (N5191, N3574, N4504);
  nand ginst1899 (N5192, N3583, N4505);
  nand ginst1900 (N5193, N3580, N4506);
  nand ginst1901 (N5196, N1326, N4508);
  nand ginst1902 (N5197, N1329, N4510);
  nand ginst1903 (N5198, N1332, N4512);
  nand ginst1904 (N5199, N1335, N4514);
  nand ginst1905 (N5200, N1338, N4516);
  nand ginst1906 (N5201, N1341, N4518);
  nand ginst1907 (N5202, N1344, N4520);
  nand ginst1908 (N5203, N1347, N4522);
  nand ginst1909 (N5204, N1350, N4524);
  nand ginst1910 (N5205, N1353, N4526);
  nand ginst1911 (N5206, N1356, N4528);
  nand ginst1912 (N5207, N1359, N4530);
  nand ginst1913 (N5208, N1362, N4532);
  nand ginst1914 (N5209, N1365, N4534);
  nand ginst1915 (N5210, N1368, N4536);
  nand ginst1916 (N5211, N1371, N4538);
  nand ginst1917 (N5212, N1374, N4540);
  nand ginst1918 (N5213, N1377, N4542);
  and ginst1919 (N528, N150, N184, N228, N240);
  nand ginst1920 (N5283, N3670, N4611);
  nand ginst1921 (N5284, N3667, N4612);
  nand ginst1922 (N5285, N3676, N4613);
  nand ginst1923 (N5286, N3673, N4614);
  nand ginst1924 (N5287, N3682, N4615);
  nand ginst1925 (N5288, N3679, N4616);
  nand ginst1926 (N5289, N3688, N4617);
  nand ginst1927 (N5290, N3685, N4618);
  nand ginst1928 (N5291, N3694, N4619);
  nand ginst1929 (N5292, N3691, N4620);
  nand ginst1930 (N5293, N3700, N4621);
  nand ginst1931 (N5294, N3697, N4622);
  nand ginst1932 (N5295, N3706, N4623);
  nand ginst1933 (N5296, N3703, N4624);
  nand ginst1934 (N5297, N3712, N4625);
  nand ginst1935 (N5298, N3709, N4626);
  nand ginst1936 (N5299, N3718, N4627);
  nand ginst1937 (N5300, N3715, N4628);
  nand ginst1938 (N5314, N3739, N4643);
  nand ginst1939 (N5315, N3736, N4644);
  nand ginst1940 (N5316, N3745, N4645);
  nand ginst1941 (N5317, N3742, N4646);
  nand ginst1942 (N5318, N3751, N4647);
  nand ginst1943 (N5319, N3748, N4648);
  nand ginst1944 (N5320, N3757, N4649);
  nand ginst1945 (N5321, N3754, N4650);
  nand ginst1946 (N5322, N3763, N4651);
  nand ginst1947 (N5323, N3760, N4652);
  not ginst1948 (N5324, N4193);
  buf ginst1949 (N535, N307);
  nand ginst1950 (N5363, N2781, N4693);
  nand ginst1951 (N5364, N3772, N4695);
  nand ginst1952 (N5365, N3769, N4696);
  nand ginst1953 (N5366, N3778, N4697);
  nand ginst1954 (N5367, N3775, N4698);
  buf ginst1955 (N537, N310);
  buf ginst1956 (N539, N313);
  buf ginst1957 (N541, N316);
  nand ginst1958 (N5425, N2790, N4745);
  nand ginst1959 (N5426, N3813, N4747);
  nand ginst1960 (N5427, N3810, N4748);
  nand ginst1961 (N5429, N2793, N4750);
  buf ginst1962 (N543, N319);
  nand ginst1963 (N5430, N3825, N4752);
  nand ginst1964 (N5431, N3822, N4753);
  nand ginst1965 (N5432, N3831, N4754);
  nand ginst1966 (N5433, N3828, N4755);
  buf ginst1967 (N545, N322);
  nand ginst1968 (N5451, N2796, N4775);
  nand ginst1969 (N5452, N3864, N4777);
  nand ginst1970 (N5453, N3861, N4778);
  nand ginst1971 (N5454, N3870, N4779);
  nand ginst1972 (N5455, N3867, N4780);
  nand ginst1973 (N5456, N3888, N4781);
  nand ginst1974 (N5457, N3885, N4782);
  not ginst1975 (N5469, N4303);
  buf ginst1976 (N547, N325);
  nand ginst1977 (N5474, N3589, N4799);
  nand ginst1978 (N5475, N3586, N4800);
  nand ginst1979 (N5476, N3595, N4801);
  nand ginst1980 (N5477, N3592, N4802);
  buf ginst1981 (N549, N328);
  buf ginst1982 (N551, N331);
  buf ginst1983 (N553, N334);
  buf ginst1984 (N556, N337);
  nand ginst1985 (N5571, N3798, N5045);
  nand ginst1986 (N5572, N3795, N5046);
  nand ginst1987 (N5573, N3804, N5047);
  nand ginst1988 (N5574, N3801, N5048);
  nand ginst1989 (N5584, N3837, N5064);
  nand ginst1990 (N5585, N3834, N5065);
  nand ginst1991 (N5586, N3843, N5066);
  nand ginst1992 (N5587, N3840, N5067);
  buf ginst1993 (N559, N343);
  nand ginst1994 (N5602, N3876, N5110);
  nand ginst1995 (N5603, N3873, N5111);
  nand ginst1996 (N5604, N3882, N5112);
  nand ginst1997 (N5605, N3879, N5113);
  buf ginst1998 (N561, N346);
  buf ginst1999 (N563, N349);
  nand ginst2000 (N5631, N4653, N5324);
  nand ginst2001 (N5632, N4463, N5167);
  nand ginst2002 (N5640, N4465, N5168);
  buf ginst2003 (N565, N352);
  nand ginst2004 (N5654, N4467, N5169);
  buf ginst2005 (N567, N355);
  nand ginst2006 (N5670, N4469, N5170);
  nand ginst2007 (N5683, N4471, N5171);
  buf ginst2008 (N569, N358);
  nand ginst2009 (N5690, N4475, N5172);
  nand ginst2010 (N5697, N4477, N5173);
  nand ginst2011 (N5707, N4479, N5174);
  buf ginst2012 (N571, N361);
  nand ginst2013 (N5718, N4481, N5175);
  nand ginst2014 (N5728, N4483, N5176);
  buf ginst2015 (N573, N364);
  not ginst2016 (N5735, N5177);
  nand ginst2017 (N5736, N4490, N5179);
  nand ginst2018 (N5740, N5180, N5181);
  nand ginst2019 (N5744, N5182, N5183);
  nand ginst2020 (N5747, N4496, N5184);
  and ginst2021 (N575, N182, N183, N185, N186);
  nand ginst2022 (N5751, N5185, N5186);
  nand ginst2023 (N5755, N5187, N5188);
  nand ginst2024 (N5758, N4502, N5189);
  nand ginst2025 (N5762, N5190, N5191);
  nand ginst2026 (N5766, N5192, N5193);
  not ginst2027 (N5769, N4803);
  not ginst2028 (N5770, N4806);
  nand ginst2029 (N5771, N4507, N5196);
  nand ginst2030 (N5778, N4509, N5197);
  and ginst2031 (N578, N152, N210, N218, N230);
  nand ginst2032 (N5789, N4511, N5198);
  nand ginst2033 (N5799, N4513, N5199);
  nand ginst2034 (N5807, N4515, N5200);
  not ginst2035 (N582, N15);
  nand ginst2036 (N5821, N4517, N5201);
  nand ginst2037 (N5837, N4519, N5202);
  not ginst2038 (N585, N5);
  nand ginst2039 (N5850, N4521, N5203);
  nand ginst2040 (N5856, N4523, N5204);
  nand ginst2041 (N5863, N4525, N5205);
  nand ginst2042 (N5870, N4527, N5206);
  nand ginst2043 (N5881, N4529, N5207);
  nand ginst2044 (N5892, N4531, N5208);
  nand ginst2045 (N5898, N4533, N5209);
  buf ginst2046 (N590, N1);
  nand ginst2047 (N5905, N4535, N5210);
  nand ginst2048 (N5915, N4537, N5211);
  nand ginst2049 (N5926, N4539, N5212);
  not ginst2050 (N593, N5);
  nand ginst2051 (N5936, N4541, N5213);
  not ginst2052 (N5943, N4817);
  nand ginst2053 (N5944, N1931, N4820);
  not ginst2054 (N5945, N4820);
  nand ginst2055 (N5946, N1932, N4823);
  not ginst2056 (N5947, N4823);
  nand ginst2057 (N5948, N1933, N4826);
  not ginst2058 (N5949, N4826);
  nand ginst2059 (N5950, N1934, N4829);
  not ginst2060 (N5951, N4829);
  nand ginst2061 (N5952, N1935, N4832);
  not ginst2062 (N5953, N4832);
  nand ginst2063 (N5954, N1936, N4835);
  not ginst2064 (N5955, N4835);
  nand ginst2065 (N5956, N1937, N4838);
  not ginst2066 (N5957, N4838);
  nand ginst2067 (N5958, N1938, N4841);
  not ginst2068 (N5959, N4841);
  not ginst2069 (N596, N5);
  and ginst2070 (N5960, N2674, N4769);
  not ginst2071 (N5966, N4844);
  nand ginst2072 (N5967, N1939, N4847);
  not ginst2073 (N5968, N4847);
  nand ginst2074 (N5969, N1940, N4850);
  not ginst2075 (N5970, N4850);
  nand ginst2076 (N5971, N1941, N4853);
  not ginst2077 (N5972, N4853);
  nand ginst2078 (N5973, N1942, N4856);
  not ginst2079 (N5974, N4856);
  nand ginst2080 (N5975, N1943, N4859);
  not ginst2081 (N5976, N4859);
  nand ginst2082 (N5977, N1944, N4862);
  not ginst2083 (N5978, N4862);
  nand ginst2084 (N5979, N1945, N4865);
  not ginst2085 (N5980, N4865);
  and ginst2086 (N5981, N2674, N4769);
  nand ginst2087 (N5989, N1946, N4868);
  not ginst2088 (N599, N289);
  not ginst2089 (N5990, N4868);
  nand ginst2090 (N5991, N5283, N5284);
  nand ginst2091 (N5996, N5285, N5286);
  nand ginst2092 (N6000, N5287, N5288);
  nand ginst2093 (N6003, N5289, N5290);
  nand ginst2094 (N6009, N5291, N5292);
  nand ginst2095 (N6014, N5293, N5294);
  nand ginst2096 (N6018, N5295, N5296);
  nand ginst2097 (N6021, N5297, N5298);
  nand ginst2098 (N6022, N5299, N5300);
  not ginst2099 (N6023, N4874);
  nand ginst2100 (N6024, N4629, N4874);
  not ginst2101 (N6025, N4877);
  nand ginst2102 (N6026, N4631, N4877);
  not ginst2103 (N6027, N4880);
  nand ginst2104 (N6028, N4633, N4880);
  not ginst2105 (N6029, N4883);
  nand ginst2106 (N6030, N4636, N4883);
  not ginst2107 (N6031, N4886);
  not ginst2108 (N6032, N4889);
  not ginst2109 (N6033, N4892);
  not ginst2110 (N6034, N4895);
  not ginst2111 (N6035, N4898);
  not ginst2112 (N6036, N4901);
  not ginst2113 (N6037, N4904);
  nand ginst2114 (N6038, N4642, N4904);
  not ginst2115 (N6039, N4907);
  not ginst2116 (N604, N299);
  not ginst2117 (N6040, N4910);
  nand ginst2118 (N6041, N5314, N5315);
  nand ginst2119 (N6047, N5316, N5317);
  nand ginst2120 (N6052, N5318, N5319);
  nand ginst2121 (N6056, N5320, N5321);
  nand ginst2122 (N6059, N5322, N5323);
  nand ginst2123 (N6060, N1968, N4913);
  not ginst2124 (N6061, N4913);
  nand ginst2125 (N6062, N1969, N4916);
  not ginst2126 (N6063, N4916);
  nand ginst2127 (N6064, N1970, N4919);
  not ginst2128 (N6065, N4919);
  nand ginst2129 (N6066, N1971, N4922);
  not ginst2130 (N6067, N4922);
  nand ginst2131 (N6068, N1972, N4925);
  not ginst2132 (N6069, N4925);
  nand ginst2133 (N6070, N1973, N4928);
  not ginst2134 (N6071, N4928);
  nand ginst2135 (N6072, N1974, N4931);
  not ginst2136 (N6073, N4931);
  nand ginst2137 (N6074, N1975, N4934);
  not ginst2138 (N6075, N4934);
  nand ginst2139 (N6076, N1976, N4937);
  not ginst2140 (N6077, N4937);
  not ginst2141 (N6078, N4940);
  nand ginst2142 (N6079, N4694, N5363);
  nand ginst2143 (N6083, N5364, N5365);
  nand ginst2144 (N6087, N5366, N5367);
  not ginst2145 (N609, N303);
  not ginst2146 (N6090, N4943);
  nand ginst2147 (N6091, N4699, N4943);
  not ginst2148 (N6092, N4946);
  not ginst2149 (N6093, N4949);
  not ginst2150 (N6094, N4952);
  not ginst2151 (N6095, N4955);
  not ginst2152 (N6096, N4970);
  nand ginst2153 (N6097, N4700, N4970);
  not ginst2154 (N6098, N4973);
  not ginst2155 (N6099, N4976);
  not ginst2156 (N6100, N4979);
  not ginst2157 (N6101, N4982);
  not ginst2158 (N6102, N4997);
  nand ginst2159 (N6103, N2015, N5000);
  not ginst2160 (N6104, N5000);
  nand ginst2161 (N6105, N2016, N5003);
  not ginst2162 (N6106, N5003);
  nand ginst2163 (N6107, N2017, N5006);
  not ginst2164 (N6108, N5006);
  nand ginst2165 (N6109, N2018, N5009);
  not ginst2166 (N6110, N5009);
  nand ginst2167 (N6111, N2019, N5012);
  not ginst2168 (N6112, N5012);
  nand ginst2169 (N6113, N2020, N5015);
  not ginst2170 (N6114, N5015);
  nand ginst2171 (N6115, N2021, N5018);
  not ginst2172 (N6116, N5018);
  nand ginst2173 (N6117, N2022, N5021);
  not ginst2174 (N6118, N5021);
  nand ginst2175 (N6119, N2023, N5024);
  not ginst2176 (N6120, N5024);
  not ginst2177 (N6121, N5033);
  nand ginst2178 (N6122, N4743, N5033);
  not ginst2179 (N6123, N5036);
  not ginst2180 (N6124, N5039);
  nand ginst2181 (N6125, N4744, N5042);
  not ginst2182 (N6126, N5042);
  nand ginst2183 (N6127, N4746, N5425);
  nand ginst2184 (N6131, N5426, N5427);
  not ginst2185 (N6135, N5049);
  nand ginst2186 (N6136, N4749, N5049);
  nand ginst2187 (N6137, N4751, N5429);
  buf ginst2188 (N614, N38);
  nand ginst2189 (N6141, N5430, N5431);
  nand ginst2190 (N6145, N5432, N5433);
  not ginst2191 (N6148, N5068);
  not ginst2192 (N6149, N5071);
  not ginst2193 (N6150, N5074);
  not ginst2194 (N6151, N5077);
  not ginst2195 (N6152, N5080);
  not ginst2196 (N6153, N5083);
  not ginst2197 (N6154, N5086);
  not ginst2198 (N6155, N5089);
  not ginst2199 (N6156, N5092);
  nand ginst2200 (N6157, N4761, N5092);
  not ginst2201 (N6158, N5095);
  nand ginst2202 (N6159, N4763, N5095);
  not ginst2203 (N6160, N5098);
  nand ginst2204 (N6161, N4765, N5098);
  not ginst2205 (N6162, N5101);
  not ginst2206 (N6163, N5104);
  nand ginst2207 (N6164, N4768, N5107);
  not ginst2208 (N6165, N5107);
  nand ginst2209 (N6166, N4776, N5451);
  nand ginst2210 (N6170, N5452, N5453);
  nand ginst2211 (N6174, N5454, N5455);
  nand ginst2212 (N6177, N5456, N5457);
  not ginst2213 (N6181, N5114);
  not ginst2214 (N6182, N5117);
  not ginst2215 (N6183, N5120);
  not ginst2216 (N6184, N5123);
  not ginst2217 (N6185, N5138);
  nand ginst2218 (N6186, N4783, N5138);
  not ginst2219 (N6187, N5141);
  not ginst2220 (N6188, N5144);
  not ginst2221 (N6189, N5147);
  not ginst2222 (N6190, N5150);
  not ginst2223 (N6191, N4784);
  nand ginst2224 (N6192, N2230, N4784);
  not ginst2225 (N6193, N4790);
  nand ginst2226 (N6194, N2765, N4790);
  not ginst2227 (N6195, N4796);
  nand ginst2228 (N6196, N5476, N5477);
  nand ginst2229 (N6199, N5474, N5475);
  not ginst2230 (N6202, N4810);
  not ginst2231 (N6203, N4814);
  buf ginst2232 (N6204, N4769);
  buf ginst2233 (N6207, N4555);
  buf ginst2234 (N6210, N4769);
  not ginst2235 (N6213, N4871);
  buf ginst2236 (N6214, N4586);
  nor ginst2237 (N6217, N2674, N4769);
  buf ginst2238 (N6220, N4667);
  not ginst2239 (N6223, N4958);
  not ginst2240 (N6224, N4961);
  not ginst2241 (N6225, N4964);
  not ginst2242 (N6226, N4967);
  not ginst2243 (N6227, N4985);
  not ginst2244 (N6228, N4988);
  not ginst2245 (N6229, N4991);
  not ginst2246 (N6230, N4994);
  not ginst2247 (N6231, N5027);
  buf ginst2248 (N6232, N4711);
  not ginst2249 (N6235, N5030);
  buf ginst2250 (N6236, N4735);
  not ginst2251 (N6239, N5052);
  not ginst2252 (N6240, N5055);
  not ginst2253 (N6241, N5058);
  not ginst2254 (N6242, N5061);
  nand ginst2255 (N6243, N5573, N5574);
  nand ginst2256 (N6246, N5571, N5572);
  nand ginst2257 (N6249, N5586, N5587);
  buf ginst2258 (N625, N15);
  nand ginst2259 (N6252, N5584, N5585);
  not ginst2260 (N6255, N5126);
  not ginst2261 (N6256, N5129);
  not ginst2262 (N6257, N5132);
  not ginst2263 (N6258, N5135);
  not ginst2264 (N6259, N5153);
  not ginst2265 (N6260, N5156);
  not ginst2266 (N6261, N5159);
  not ginst2267 (N6262, N5162);
  nand ginst2268 (N6263, N5604, N5605);
  nand ginst2269 (N6266, N5602, N5603);
  nand ginst2270 (N628, N9, N12);
  nand ginst2271 (N632, N9, N12);
  buf ginst2272 (N636, N38);
  not ginst2273 (N641, N245);
  not ginst2274 (N642, N248);
  buf ginst2275 (N643, N251);
  not ginst2276 (N644, N251);
  not ginst2277 (N651, N254);
  nand ginst2278 (N6540, N1380, N5945);
  nand ginst2279 (N6541, N1383, N5947);
  nand ginst2280 (N6542, N1386, N5949);
  nand ginst2281 (N6543, N1389, N5951);
  nand ginst2282 (N6544, N1392, N5953);
  nand ginst2283 (N6545, N1395, N5955);
  nand ginst2284 (N6546, N1398, N5957);
  nand ginst2285 (N6547, N1401, N5959);
  nand ginst2286 (N6555, N1404, N5968);
  nand ginst2287 (N6556, N1407, N5970);
  nand ginst2288 (N6557, N1410, N5972);
  nand ginst2289 (N6558, N1413, N5974);
  nand ginst2290 (N6559, N1416, N5976);
  nand ginst2291 (N6560, N1419, N5978);
  nand ginst2292 (N6561, N1422, N5980);
  nand ginst2293 (N6569, N1425, N5990);
  buf ginst2294 (N657, N106);
  nand ginst2295 (N6594, N3721, N6023);
  nand ginst2296 (N6595, N3724, N6025);
  nand ginst2297 (N6596, N3727, N6027);
  nand ginst2298 (N6597, N3730, N6029);
  nand ginst2299 (N6598, N4889, N6031);
  nand ginst2300 (N6599, N4886, N6032);
  not ginst2301 (N660, N257);
  nand ginst2302 (N6600, N4895, N6033);
  nand ginst2303 (N6601, N4892, N6034);
  nand ginst2304 (N6602, N4901, N6035);
  nand ginst2305 (N6603, N4898, N6036);
  nand ginst2306 (N6604, N3733, N6037);
  nand ginst2307 (N6605, N4910, N6039);
  nand ginst2308 (N6606, N4907, N6040);
  nand ginst2309 (N6621, N1434, N6061);
  nand ginst2310 (N6622, N1437, N6063);
  nand ginst2311 (N6623, N1440, N6065);
  nand ginst2312 (N6624, N1443, N6067);
  nand ginst2313 (N6625, N1446, N6069);
  nand ginst2314 (N6626, N1449, N6071);
  nand ginst2315 (N6627, N1452, N6073);
  nand ginst2316 (N6628, N1455, N6075);
  nand ginst2317 (N6629, N1458, N6077);
  nand ginst2318 (N6639, N3783, N6090);
  nand ginst2319 (N6640, N4949, N6092);
  nand ginst2320 (N6641, N4946, N6093);
  nand ginst2321 (N6642, N4955, N6094);
  nand ginst2322 (N6643, N4952, N6095);
  nand ginst2323 (N6644, N3786, N6096);
  nand ginst2324 (N6645, N4976, N6098);
  nand ginst2325 (N6646, N4973, N6099);
  nand ginst2326 (N6647, N4982, N6100);
  nand ginst2327 (N6648, N4979, N6101);
  nand ginst2328 (N6649, N1461, N6104);
  nand ginst2329 (N6650, N1464, N6106);
  nand ginst2330 (N6651, N1467, N6108);
  nand ginst2331 (N6652, N1470, N6110);
  nand ginst2332 (N6653, N1473, N6112);
  nand ginst2333 (N6654, N1476, N6114);
  nand ginst2334 (N6655, N1479, N6116);
  nand ginst2335 (N6656, N1482, N6118);
  nand ginst2336 (N6657, N1485, N6120);
  nand ginst2337 (N6658, N3789, N6121);
  nand ginst2338 (N6659, N5039, N6123);
  not ginst2339 (N666, N260);
  nand ginst2340 (N6660, N5036, N6124);
  nand ginst2341 (N6661, N3792, N6126);
  nand ginst2342 (N6668, N3816, N6135);
  nand ginst2343 (N6677, N5071, N6148);
  nand ginst2344 (N6678, N5068, N6149);
  nand ginst2345 (N6679, N5077, N6150);
  nand ginst2346 (N6680, N5074, N6151);
  nand ginst2347 (N6681, N5083, N6152);
  nand ginst2348 (N6682, N5080, N6153);
  nand ginst2349 (N6683, N5089, N6154);
  nand ginst2350 (N6684, N5086, N6155);
  nand ginst2351 (N6685, N3846, N6156);
  nand ginst2352 (N6686, N3849, N6158);
  nand ginst2353 (N6687, N3852, N6160);
  nand ginst2354 (N6688, N5104, N6162);
  nand ginst2355 (N6689, N5101, N6163);
  nand ginst2356 (N6690, N3855, N6165);
  nand ginst2357 (N6702, N5117, N6181);
  nand ginst2358 (N6703, N5114, N6182);
  nand ginst2359 (N6704, N5123, N6183);
  nand ginst2360 (N6705, N5120, N6184);
  nand ginst2361 (N6706, N3891, N6185);
  nand ginst2362 (N6707, N5144, N6187);
  nand ginst2363 (N6708, N5141, N6188);
  nand ginst2364 (N6709, N5150, N6189);
  nand ginst2365 (N6710, N5147, N6190);
  nand ginst2366 (N6711, N1708, N6191);
  nand ginst2367 (N6712, N2231, N6193);
  not ginst2368 (N672, N263);
  nand ginst2369 (N6729, N4961, N6223);
  not ginst2370 (N673, N267);
  nand ginst2371 (N6730, N4958, N6224);
  nand ginst2372 (N6731, N4967, N6225);
  nand ginst2373 (N6732, N4964, N6226);
  nand ginst2374 (N6733, N4988, N6227);
  nand ginst2375 (N6734, N4985, N6228);
  nand ginst2376 (N6735, N4994, N6229);
  nand ginst2377 (N6736, N4991, N6230);
  not ginst2378 (N674, N106);
  nand ginst2379 (N6741, N5055, N6239);
  nand ginst2380 (N6742, N5052, N6240);
  nand ginst2381 (N6743, N5061, N6241);
  nand ginst2382 (N6744, N5058, N6242);
  nand ginst2383 (N6751, N5129, N6255);
  nand ginst2384 (N6752, N5126, N6256);
  nand ginst2385 (N6753, N5135, N6257);
  nand ginst2386 (N6754, N5132, N6258);
  nand ginst2387 (N6755, N5156, N6259);
  nand ginst2388 (N6756, N5153, N6260);
  nand ginst2389 (N6757, N5162, N6261);
  nand ginst2390 (N6758, N5159, N6262);
  buf ginst2391 (N676, N18);
  not ginst2392 (N6761, N5892);
  and ginst2393 (N6762, N5632, N5640, N5654, N5670, N5683);
  and ginst2394 (N6766, N3097, N5632);
  and ginst2395 (N6767, N3101, N5632, N5640);
  and ginst2396 (N6768, N3107, N5632, N5640, N5654);
  and ginst2397 (N6769, N3114, N5632, N5640, N5654, N5670);
  and ginst2398 (N6770, N3101, N5640);
  and ginst2399 (N6771, N3107, N5640, N5654);
  and ginst2400 (N6772, N3114, N5640, N5654, N5670);
  and ginst2401 (N6773, N5640, N5654, N5670, N5683);
  and ginst2402 (N6774, N3101, N5640);
  and ginst2403 (N6775, N3107, N5640, N5654);
  and ginst2404 (N6776, N3114, N5640, N5654, N5670);
  and ginst2405 (N6777, N3107, N5654);
  and ginst2406 (N6778, N3114, N5654, N5670);
  and ginst2407 (N6779, N5654, N5670, N5683);
  and ginst2408 (N6780, N3107, N5654);
  and ginst2409 (N6781, N3114, N5654, N5670);
  and ginst2410 (N6782, N3114, N5670);
  and ginst2411 (N6783, N5670, N5683);
  and ginst2412 (N6784, N5690, N5697, N5707, N5718, N5728);
  and ginst2413 (N6787, N3137, N5690);
  and ginst2414 (N6788, N3140, N5690, N5697);
  and ginst2415 (N6789, N3144, N5690, N5697, N5707);
  and ginst2416 (N6790, N3149, N5690, N5697, N5707, N5718);
  and ginst2417 (N6791, N3140, N5697);
  and ginst2418 (N6792, N3144, N5697, N5707);
  and ginst2419 (N6793, N3149, N5697, N5707, N5718);
  and ginst2420 (N6794, N3144, N5707);
  and ginst2421 (N6795, N3149, N5707, N5718);
  and ginst2422 (N6796, N3149, N5718);
  not ginst2423 (N6797, N5736);
  not ginst2424 (N6800, N5740);
  not ginst2425 (N6803, N5747);
  not ginst2426 (N6806, N5751);
  not ginst2427 (N6809, N5758);
  not ginst2428 (N6812, N5762);
  buf ginst2429 (N6815, N5744);
  buf ginst2430 (N6818, N5744);
  buf ginst2431 (N682, N18);
  buf ginst2432 (N6821, N5755);
  buf ginst2433 (N6824, N5755);
  buf ginst2434 (N6827, N5766);
  buf ginst2435 (N6830, N5766);
  and ginst2436 (N6833, N5771, N5778, N5789, N5850);
  and ginst2437 (N6836, N3169, N5771);
  and ginst2438 (N6837, N3173, N5771, N5778);
  and ginst2439 (N6838, N3178, N5771, N5778, N5789);
  and ginst2440 (N6839, N3173, N5778);
  and ginst2441 (N6840, N3178, N5778, N5789);
  and ginst2442 (N6841, N5778, N5789, N5850);
  and ginst2443 (N6842, N3173, N5778);
  and ginst2444 (N6843, N3178, N5778, N5789);
  and ginst2445 (N6844, N3178, N5789);
  and ginst2446 (N6845, N5799, N5807, N5821, N5837, N5856);
  and ginst2447 (N6848, N3185, N5799);
  and ginst2448 (N6849, N3189, N5799, N5807);
  and ginst2449 (N6850, N3195, N5799, N5807, N5821);
  and ginst2450 (N6851, N3202, N5799, N5807, N5821, N5837);
  and ginst2451 (N6852, N3189, N5807);
  and ginst2452 (N6853, N3195, N5807, N5821);
  and ginst2453 (N6854, N3202, N5807, N5821, N5837);
  and ginst2454 (N6855, N5807, N5821, N5837, N5856);
  and ginst2455 (N6856, N3189, N5807);
  and ginst2456 (N6857, N3195, N5807, N5821);
  and ginst2457 (N6858, N3202, N5807, N5821, N5837);
  and ginst2458 (N6859, N3195, N5821);
  and ginst2459 (N6860, N3202, N5821, N5837);
  and ginst2460 (N6861, N5821, N5837, N5856);
  and ginst2461 (N6862, N3195, N5821);
  and ginst2462 (N6863, N3202, N5821, N5837);
  and ginst2463 (N6864, N3202, N5837);
  and ginst2464 (N6865, N5789, N5850);
  and ginst2465 (N6866, N5837, N5856);
  and ginst2466 (N6867, N5863, N5870, N5881, N5892);
  and ginst2467 (N6870, N3211, N5863);
  and ginst2468 (N6871, N3215, N5863, N5870);
  and ginst2469 (N6872, N3221, N5863, N5870, N5881);
  and ginst2470 (N6873, N3215, N5870);
  and ginst2471 (N6874, N3221, N5870, N5881);
  and ginst2472 (N6875, N5870, N5881, N5892);
  and ginst2473 (N6876, N3215, N5870);
  and ginst2474 (N6877, N3221, N5870, N5881);
  and ginst2475 (N6878, N3221, N5881);
  and ginst2476 (N6879, N5881, N5892);
  and ginst2477 (N688, N263, N382);
  and ginst2478 (N6880, N3221, N5881);
  and ginst2479 (N6881, N5898, N5905, N5915, N5926, N5936);
  and ginst2480 (N6884, N3229, N5898);
  and ginst2481 (N6885, N3232, N5898, N5905);
  and ginst2482 (N6886, N3236, N5898, N5905, N5915);
  and ginst2483 (N6887, N3241, N5898, N5905, N5915, N5926);
  and ginst2484 (N6888, N3232, N5905);
  and ginst2485 (N6889, N3236, N5905, N5915);
  buf ginst2486 (N689, N18);
  and ginst2487 (N6890, N3241, N5905, N5915, N5926);
  and ginst2488 (N6891, N3236, N5915);
  and ginst2489 (N6892, N3241, N5915, N5926);
  and ginst2490 (N6893, N3241, N5926);
  nand ginst2491 (N6894, N5944, N6540);
  nand ginst2492 (N6901, N5946, N6541);
  nand ginst2493 (N6912, N5948, N6542);
  nand ginst2494 (N6923, N5950, N6543);
  nand ginst2495 (N6929, N5952, N6544);
  nand ginst2496 (N6936, N5954, N6545);
  nand ginst2497 (N6946, N5956, N6546);
  not ginst2498 (N695, N18);
  nand ginst2499 (N6957, N5958, N6547);
  nand ginst2500 (N6967, N4575, N6204);
  not ginst2501 (N6968, N6204);
  not ginst2502 (N6969, N6207);
  nand ginst2503 (N6970, N5967, N6555);
  nand ginst2504 (N6977, N5969, N6556);
  nand ginst2505 (N6988, N5971, N6557);
  nand ginst2506 (N6998, N5973, N6558);
  nand ginst2507 (N700, N267, N382);
  nand ginst2508 (N7006, N5975, N6559);
  nand ginst2509 (N7020, N5977, N6560);
  nand ginst2510 (N7036, N5979, N6561);
  nand ginst2511 (N7049, N5989, N6569);
  not ginst2512 (N705, N271);
  nand ginst2513 (N7055, N4610, N6210);
  not ginst2514 (N7056, N6210);
  and ginst2515 (N7057, N5991, N5996, N6000, N6021);
  not ginst2516 (N706, N274);
  and ginst2517 (N7060, N3362, N5991);
  and ginst2518 (N7061, N3363, N5991, N5996);
  and ginst2519 (N7062, N3364, N5991, N5996, N6000);
  and ginst2520 (N7063, N6003, N6009, N6014, N6018, N6022);
  and ginst2521 (N7064, N3366, N6003);
  and ginst2522 (N7065, N3367, N6003, N6009);
  and ginst2523 (N7066, N3368, N6003, N6009, N6014);
  and ginst2524 (N7067, N3369, N6003, N6009, N6014, N6018);
  nand ginst2525 (N7068, N6024, N6594);
  buf ginst2526 (N707, N277);
  nand ginst2527 (N7073, N6026, N6595);
  nand ginst2528 (N7077, N6028, N6596);
  not ginst2529 (N708, N277);
  nand ginst2530 (N7080, N6030, N6597);
  nand ginst2531 (N7086, N6598, N6599);
  nand ginst2532 (N7091, N6600, N6601);
  nand ginst2533 (N7095, N6602, N6603);
  nand ginst2534 (N7098, N6038, N6604);
  nand ginst2535 (N7099, N6605, N6606);
  and ginst2536 (N7100, N6041, N6047, N6052, N6056, N6059);
  and ginst2537 (N7103, N3371, N6041);
  and ginst2538 (N7104, N3372, N6041, N6047);
  and ginst2539 (N7105, N3373, N6041, N6047, N6052);
  and ginst2540 (N7106, N3374, N6041, N6047, N6052, N6056);
  nand ginst2541 (N7107, N6060, N6621);
  nand ginst2542 (N7114, N6062, N6622);
  nand ginst2543 (N7125, N6064, N6623);
  nand ginst2544 (N7136, N6066, N6624);
  nand ginst2545 (N7142, N6068, N6625);
  nand ginst2546 (N7149, N6070, N6626);
  not ginst2547 (N715, N280);
  nand ginst2548 (N7159, N6072, N6627);
  nand ginst2549 (N7170, N6074, N6628);
  nand ginst2550 (N7180, N6076, N6629);
  not ginst2551 (N7187, N6220);
  not ginst2552 (N7188, N6079);
  not ginst2553 (N7191, N6083);
  nand ginst2554 (N7194, N6091, N6639);
  nand ginst2555 (N7198, N6640, N6641);
  nand ginst2556 (N7202, N6642, N6643);
  nand ginst2557 (N7205, N6097, N6644);
  nand ginst2558 (N7209, N6645, N6646);
  not ginst2559 (N721, N283);
  nand ginst2560 (N7213, N6647, N6648);
  buf ginst2561 (N7216, N6087);
  buf ginst2562 (N7219, N6087);
  nand ginst2563 (N7222, N6103, N6649);
  nand ginst2564 (N7229, N6105, N6650);
  nand ginst2565 (N7240, N6107, N6651);
  nand ginst2566 (N7250, N6109, N6652);
  nand ginst2567 (N7258, N6111, N6653);
  not ginst2568 (N727, N286);
  nand ginst2569 (N7272, N6113, N6654);
  nand ginst2570 (N7288, N6115, N6655);
  nand ginst2571 (N7301, N6117, N6656);
  nand ginst2572 (N7307, N6119, N6657);
  nand ginst2573 (N7314, N6122, N6658);
  nand ginst2574 (N7318, N6659, N6660);
  nand ginst2575 (N7322, N6125, N6661);
  not ginst2576 (N7325, N6127);
  not ginst2577 (N7328, N6131);
  not ginst2578 (N733, N289);
  nand ginst2579 (N7331, N6136, N6668);
  not ginst2580 (N7334, N6137);
  not ginst2581 (N7337, N6141);
  not ginst2582 (N734, N293);
  buf ginst2583 (N7340, N6145);
  buf ginst2584 (N7343, N6145);
  nand ginst2585 (N7346, N6677, N6678);
  nand ginst2586 (N7351, N6679, N6680);
  nand ginst2587 (N7355, N6681, N6682);
  nand ginst2588 (N7358, N6683, N6684);
  nand ginst2589 (N7364, N6157, N6685);
  nand ginst2590 (N7369, N6159, N6686);
  nand ginst2591 (N7373, N6161, N6687);
  nand ginst2592 (N7376, N6688, N6689);
  nand ginst2593 (N7377, N6164, N6690);
  not ginst2594 (N7378, N6166);
  not ginst2595 (N7381, N6170);
  not ginst2596 (N7384, N6177);
  nand ginst2597 (N7387, N6702, N6703);
  nand ginst2598 (N7391, N6704, N6705);
  nand ginst2599 (N7394, N6186, N6706);
  nand ginst2600 (N7398, N6707, N6708);
  nand ginst2601 (N7402, N6709, N6710);
  buf ginst2602 (N7405, N6174);
  buf ginst2603 (N7408, N6174);
  buf ginst2604 (N7411, N5936);
  buf ginst2605 (N7414, N5898);
  buf ginst2606 (N7417, N5905);
  not ginst2607 (N742, N296);
  buf ginst2608 (N7420, N5915);
  buf ginst2609 (N7423, N5926);
  buf ginst2610 (N7426, N5728);
  buf ginst2611 (N7429, N5690);
  buf ginst2612 (N7432, N5697);
  buf ginst2613 (N7435, N5707);
  buf ginst2614 (N7438, N5718);
  nand ginst2615 (N7441, N6192, N6711);
  nand ginst2616 (N7444, N6194, N6712);
  buf ginst2617 (N7447, N5683);
  buf ginst2618 (N7450, N5670);
  buf ginst2619 (N7453, N5632);
  buf ginst2620 (N7456, N5654);
  buf ginst2621 (N7459, N5640);
  buf ginst2622 (N7462, N5640);
  buf ginst2623 (N7465, N5683);
  buf ginst2624 (N7468, N5670);
  buf ginst2625 (N7471, N5632);
  buf ginst2626 (N7474, N5654);
  not ginst2627 (N7477, N6196);
  not ginst2628 (N7478, N6199);
  buf ginst2629 (N7479, N5850);
  not ginst2630 (N748, N299);
  buf ginst2631 (N7482, N5789);
  buf ginst2632 (N7485, N5771);
  buf ginst2633 (N7488, N5778);
  not ginst2634 (N749, N303);
  buf ginst2635 (N7491, N5850);
  buf ginst2636 (N7494, N5789);
  buf ginst2637 (N7497, N5771);
  buf ginst2638 (N750, N367);
  buf ginst2639 (N7500, N5778);
  buf ginst2640 (N7503, N5856);
  buf ginst2641 (N7506, N5837);
  buf ginst2642 (N7509, N5799);
  buf ginst2643 (N7512, N5821);
  buf ginst2644 (N7515, N5807);
  buf ginst2645 (N7518, N5807);
  buf ginst2646 (N7521, N5856);
  buf ginst2647 (N7524, N5837);
  buf ginst2648 (N7527, N5799);
  buf ginst2649 (N7530, N5821);
  buf ginst2650 (N7533, N5863);
  buf ginst2651 (N7536, N5863);
  buf ginst2652 (N7539, N5870);
  buf ginst2653 (N7542, N5870);
  buf ginst2654 (N7545, N5881);
  buf ginst2655 (N7548, N5881);
  not ginst2656 (N7551, N6214);
  not ginst2657 (N7552, N6217);
  buf ginst2658 (N7553, N5981);
  not ginst2659 (N7556, N6249);
  not ginst2660 (N7557, N6252);
  not ginst2661 (N7558, N6243);
  not ginst2662 (N7559, N6246);
  nand ginst2663 (N7560, N6731, N6732);
  nand ginst2664 (N7563, N6729, N6730);
  nand ginst2665 (N7566, N6735, N6736);
  nand ginst2666 (N7569, N6733, N6734);
  not ginst2667 (N7572, N6232);
  not ginst2668 (N7573, N6236);
  nand ginst2669 (N7574, N6743, N6744);
  nand ginst2670 (N7577, N6741, N6742);
  not ginst2671 (N758, N307);
  not ginst2672 (N7580, N6263);
  not ginst2673 (N7581, N6266);
  nand ginst2674 (N7582, N6753, N6754);
  nand ginst2675 (N7585, N6751, N6752);
  nand ginst2676 (N7588, N6757, N6758);
  not ginst2677 (N759, N310);
  nand ginst2678 (N7591, N6755, N6756);
  or ginst2679 (N7609, N3096, N6766, N6767, N6768, N6769);
  or ginst2680 (N7613, N3107, N6782);
  not ginst2681 (N762, N313);
  or ginst2682 (N7620, N3136, N6787, N6788, N6789, N6790);
  or ginst2683 (N7649, N3168, N6836, N6837, N6838);
  or ginst2684 (N7650, N3173, N6844);
  or ginst2685 (N7655, N3184, N6848, N6849, N6850, N6851);
  or ginst2686 (N7659, N3195, N6864);
  or ginst2687 (N7668, N3210, N6870, N6871, N6872);
  or ginst2688 (N7671, N3228, N6884, N6885, N6886, N6887);
  not ginst2689 (N768, N316);
  not ginst2690 (N774, N319);
  nand ginst2691 (N7744, N3661, N6968);
  not ginst2692 (N780, N322);
  nand ginst2693 (N7822, N3664, N7056);
  or ginst2694 (N7825, N3361, N7060, N7061, N7062);
  or ginst2695 (N7826, N3365, N7064, N7065, N7066, N7067);
  or ginst2696 (N7852, N3370, N7103, N7104, N7105, N7106);
  not ginst2697 (N786, N325);
  not ginst2698 (N794, N328);
  not ginst2699 (N800, N331);
  not ginst2700 (N806, N334);
  or ginst2701 (N8114, N3101, N6777, N6778, N6779);
  or ginst2702 (N8117, N3097, N6770, N6771, N6772, N6773);
  not ginst2703 (N812, N337);
  buf ginst2704 (N813, N340);
  nor ginst2705 (N8131, N3101, N6780, N6781);
  nor ginst2706 (N8134, N3097, N6774, N6775, N6776);
  not ginst2707 (N814, N340);
  nand ginst2708 (N8144, N6199, N7477);
  nand ginst2709 (N8145, N6196, N7478);
  or ginst2710 (N8146, N3169, N6839, N6840, N6841);
  nor ginst2711 (N8156, N3169, N6842, N6843);
  or ginst2712 (N8166, N3189, N6859, N6860, N6861);
  or ginst2713 (N8169, N3185, N6852, N6853, N6854, N6855);
  nor ginst2714 (N8183, N3189, N6862, N6863);
  nor ginst2715 (N8186, N3185, N6856, N6857, N6858);
  or ginst2716 (N8196, N3211, N6873, N6874, N6875);
  nor ginst2717 (N8200, N3211, N6876, N6877);
  or ginst2718 (N8204, N3215, N6878, N6879);
  nor ginst2719 (N8208, N3215, N6880);
  not ginst2720 (N821, N343);
  nand ginst2721 (N8216, N6252, N7556);
  nand ginst2722 (N8217, N6249, N7557);
  nand ginst2723 (N8218, N6246, N7558);
  nand ginst2724 (N8219, N6243, N7559);
  nand ginst2725 (N8232, N6266, N7580);
  nand ginst2726 (N8233, N6263, N7581);
  not ginst2727 (N8242, N7411);
  not ginst2728 (N8243, N7414);
  not ginst2729 (N8244, N7417);
  not ginst2730 (N8245, N7420);
  not ginst2731 (N8246, N7423);
  not ginst2732 (N8247, N7426);
  not ginst2733 (N8248, N7429);
  not ginst2734 (N8249, N7432);
  not ginst2735 (N8250, N7435);
  not ginst2736 (N8251, N7438);
  not ginst2737 (N8252, N7136);
  not ginst2738 (N8253, N6923);
  not ginst2739 (N8254, N6762);
  not ginst2740 (N8260, N7459);
  not ginst2741 (N8261, N7462);
  and ginst2742 (N8262, N3122, N6762);
  and ginst2743 (N8269, N3155, N6784);
  not ginst2744 (N827, N346);
  not ginst2745 (N8274, N6815);
  not ginst2746 (N8275, N6818);
  not ginst2747 (N8276, N6821);
  not ginst2748 (N8277, N6824);
  not ginst2749 (N8278, N6827);
  not ginst2750 (N8279, N6830);
  and ginst2751 (N8280, N5736, N5740, N6815);
  and ginst2752 (N8281, N6797, N6800, N6818);
  and ginst2753 (N8282, N5747, N5751, N6821);
  and ginst2754 (N8283, N6803, N6806, N6824);
  and ginst2755 (N8284, N5758, N5762, N6827);
  and ginst2756 (N8285, N6809, N6812, N6830);
  not ginst2757 (N8288, N6845);
  not ginst2758 (N8294, N7488);
  not ginst2759 (N8295, N7500);
  not ginst2760 (N8296, N7515);
  not ginst2761 (N8297, N7518);
  and ginst2762 (N8298, N6833, N6845);
  and ginst2763 (N8307, N6867, N6881);
  not ginst2764 (N8315, N7533);
  not ginst2765 (N8317, N7536);
  not ginst2766 (N8319, N7539);
  not ginst2767 (N8321, N7542);
  nand ginst2768 (N8322, N4543, N7545);
  not ginst2769 (N8323, N7545);
  nand ginst2770 (N8324, N5943, N7548);
  not ginst2771 (N8325, N7548);
  nand ginst2772 (N8326, N6967, N7744);
  not ginst2773 (N833, N349);
  and ginst2774 (N8333, N6894, N6901, N6912, N6923);
  and ginst2775 (N8337, N4545, N6894);
  and ginst2776 (N8338, N4549, N6894, N6901);
  and ginst2777 (N8339, N4555, N6894, N6901, N6912);
  and ginst2778 (N8340, N4549, N6901);
  and ginst2779 (N8341, N4555, N6901, N6912);
  and ginst2780 (N8342, N6901, N6912, N6923);
  and ginst2781 (N8343, N4549, N6901);
  and ginst2782 (N8344, N4555, N6901, N6912);
  and ginst2783 (N8345, N4555, N6912);
  and ginst2784 (N8346, N6912, N6923);
  and ginst2785 (N8347, N4555, N6912);
  and ginst2786 (N8348, N4563, N6929);
  and ginst2787 (N8349, N4566, N6929, N6936);
  and ginst2788 (N8350, N4570, N6929, N6936, N6946);
  and ginst2789 (N8351, N5960, N6929, N6936, N6946, N6957);
  and ginst2790 (N8352, N4566, N6936);
  and ginst2791 (N8353, N4570, N6936, N6946);
  and ginst2792 (N8354, N5960, N6936, N6946, N6957);
  and ginst2793 (N8355, N4570, N6946);
  and ginst2794 (N8356, N5960, N6946, N6957);
  and ginst2795 (N8357, N5960, N6957);
  nand ginst2796 (N8358, N7055, N7822);
  and ginst2797 (N8365, N6970, N6977, N6988, N7049);
  and ginst2798 (N8369, N4577, N6970);
  and ginst2799 (N8370, N4581, N6970, N6977);
  and ginst2800 (N8371, N4586, N6970, N6977, N6988);
  and ginst2801 (N8372, N4581, N6977);
  and ginst2802 (N8373, N4586, N6977, N6988);
  and ginst2803 (N8374, N6977, N6988, N7049);
  and ginst2804 (N8375, N4581, N6977);
  and ginst2805 (N8376, N4586, N6977, N6988);
  and ginst2806 (N8377, N4586, N6988);
  and ginst2807 (N8378, N4593, N6998);
  and ginst2808 (N8379, N4597, N6998, N7006);
  and ginst2809 (N8380, N4603, N6998, N7006, N7020);
  and ginst2810 (N8381, N5981, N6998, N7006, N7020, N7036);
  and ginst2811 (N8382, N4597, N7006);
  and ginst2812 (N8383, N4603, N7006, N7020);
  and ginst2813 (N8384, N5981, N7006, N7020, N7036);
  and ginst2814 (N8385, N4597, N7006);
  and ginst2815 (N8386, N4603, N7006, N7020);
  and ginst2816 (N8387, N5981, N7006, N7020, N7036);
  and ginst2817 (N8388, N4603, N7020);
  and ginst2818 (N8389, N5981, N7020, N7036);
  not ginst2819 (N839, N352);
  and ginst2820 (N8390, N4603, N7020);
  and ginst2821 (N8391, N5981, N7020, N7036);
  and ginst2822 (N8392, N5981, N7036);
  and ginst2823 (N8393, N6988, N7049);
  and ginst2824 (N8394, N7057, N7063);
  and ginst2825 (N8404, N7057, N7826);
  and ginst2826 (N8405, N7068, N7073, N7077, N7098);
  and ginst2827 (N8409, N4632, N7068);
  and ginst2828 (N8410, N4634, N7068, N7073);
  and ginst2829 (N8411, N4635, N7068, N7073, N7077);
  and ginst2830 (N8412, N7080, N7086, N7091, N7095, N7099);
  and ginst2831 (N8415, N4638, N7080);
  and ginst2832 (N8416, N4639, N7080, N7086);
  and ginst2833 (N8417, N4640, N7080, N7086, N7091);
  and ginst2834 (N8418, N4641, N7080, N7086, N7091, N7095);
  and ginst2835 (N8421, N3375, N7100);
  and ginst2836 (N8430, N7107, N7114, N7125, N7136);
  and ginst2837 (N8433, N4657, N7107);
  and ginst2838 (N8434, N4661, N7107, N7114);
  and ginst2839 (N8435, N4667, N7107, N7114, N7125);
  and ginst2840 (N8436, N4661, N7114);
  and ginst2841 (N8437, N4667, N7114, N7125);
  and ginst2842 (N8438, N7114, N7125, N7136);
  and ginst2843 (N8439, N4661, N7114);
  and ginst2844 (N8440, N4667, N7114, N7125);
  and ginst2845 (N8441, N4667, N7125);
  and ginst2846 (N8442, N7125, N7136);
  and ginst2847 (N8443, N4667, N7125);
  and ginst2848 (N8444, N7142, N7149, N7159, N7170, N7180);
  and ginst2849 (N8447, N4675, N7142);
  and ginst2850 (N8448, N4678, N7142, N7149);
  and ginst2851 (N8449, N4682, N7142, N7149, N7159);
  not ginst2852 (N845, N355);
  and ginst2853 (N8450, N4687, N7142, N7149, N7159, N7170);
  and ginst2854 (N8451, N4678, N7149);
  and ginst2855 (N8452, N4682, N7149, N7159);
  and ginst2856 (N8453, N4687, N7149, N7159, N7170);
  and ginst2857 (N8454, N4682, N7159);
  and ginst2858 (N8455, N4687, N7159, N7170);
  and ginst2859 (N8456, N4687, N7170);
  not ginst2860 (N8457, N7194);
  not ginst2861 (N8460, N7198);
  not ginst2862 (N8463, N7205);
  not ginst2863 (N8466, N7209);
  not ginst2864 (N8469, N7216);
  not ginst2865 (N8470, N7219);
  buf ginst2866 (N8471, N7202);
  buf ginst2867 (N8474, N7202);
  buf ginst2868 (N8477, N7213);
  buf ginst2869 (N8480, N7213);
  and ginst2870 (N8483, N6079, N6083, N7216);
  and ginst2871 (N8484, N7188, N7191, N7219);
  and ginst2872 (N8485, N7222, N7229, N7240, N7301);
  and ginst2873 (N8488, N4702, N7222);
  and ginst2874 (N8489, N4706, N7222, N7229);
  and ginst2875 (N8490, N4711, N7222, N7229, N7240);
  and ginst2876 (N8491, N4706, N7229);
  and ginst2877 (N8492, N4711, N7229, N7240);
  and ginst2878 (N8493, N7229, N7240, N7301);
  and ginst2879 (N8494, N4706, N7229);
  and ginst2880 (N8495, N4711, N7229, N7240);
  and ginst2881 (N8496, N4711, N7240);
  and ginst2882 (N8497, N7250, N7258, N7272, N7288, N7307);
  and ginst2883 (N8500, N4718, N7250);
  and ginst2884 (N8501, N4722, N7250, N7258);
  and ginst2885 (N8502, N4728, N7250, N7258, N7272);
  and ginst2886 (N8503, N4735, N7250, N7258, N7272, N7288);
  and ginst2887 (N8504, N4722, N7258);
  and ginst2888 (N8505, N4728, N7258, N7272);
  and ginst2889 (N8506, N4735, N7258, N7272, N7288);
  and ginst2890 (N8507, N7258, N7272, N7288, N7307);
  and ginst2891 (N8508, N4722, N7258);
  and ginst2892 (N8509, N4728, N7258, N7272);
  and ginst2893 (N8510, N4735, N7258, N7272, N7288);
  and ginst2894 (N8511, N4728, N7272);
  and ginst2895 (N8512, N4735, N7272, N7288);
  and ginst2896 (N8513, N7272, N7288, N7307);
  and ginst2897 (N8514, N4728, N7272);
  and ginst2898 (N8515, N4735, N7272, N7288);
  and ginst2899 (N8516, N4735, N7288);
  and ginst2900 (N8517, N7240, N7301);
  and ginst2901 (N8518, N7288, N7307);
  not ginst2902 (N8519, N7314);
  not ginst2903 (N8522, N7318);
  buf ginst2904 (N8525, N7322);
  buf ginst2905 (N8528, N7322);
  not ginst2906 (N853, N358);
  buf ginst2907 (N8531, N7331);
  buf ginst2908 (N8534, N7331);
  not ginst2909 (N8537, N7340);
  not ginst2910 (N8538, N7343);
  and ginst2911 (N8539, N6137, N6141, N7340);
  and ginst2912 (N8540, N7334, N7337, N7343);
  and ginst2913 (N8541, N7346, N7351, N7355, N7376);
  and ginst2914 (N8545, N4757, N7346);
  and ginst2915 (N8546, N4758, N7346, N7351);
  and ginst2916 (N8547, N4759, N7346, N7351, N7355);
  and ginst2917 (N8548, N7358, N7364, N7369, N7373, N7377);
  and ginst2918 (N8551, N4762, N7358);
  and ginst2919 (N8552, N4764, N7358, N7364);
  and ginst2920 (N8553, N4766, N7358, N7364, N7369);
  and ginst2921 (N8554, N4767, N7358, N7364, N7369, N7373);
  not ginst2922 (N8555, N7387);
  not ginst2923 (N8558, N7394);
  not ginst2924 (N8561, N7398);
  not ginst2925 (N8564, N7405);
  not ginst2926 (N8565, N7408);
  buf ginst2927 (N8566, N7391);
  buf ginst2928 (N8569, N7391);
  buf ginst2929 (N8572, N7402);
  buf ginst2930 (N8575, N7402);
  and ginst2931 (N8578, N6166, N6170, N7405);
  and ginst2932 (N8579, N7378, N7381, N7408);
  buf ginst2933 (N8580, N7180);
  buf ginst2934 (N8583, N7142);
  buf ginst2935 (N8586, N7149);
  buf ginst2936 (N8589, N7159);
  not ginst2937 (N859, N361);
  buf ginst2938 (N8592, N7170);
  buf ginst2939 (N8595, N6929);
  buf ginst2940 (N8598, N6936);
  buf ginst2941 (N8601, N6946);
  buf ginst2942 (N8604, N6957);
  not ginst2943 (N8607, N7441);
  nand ginst2944 (N8608, N5469, N7441);
  not ginst2945 (N8609, N7444);
  nand ginst2946 (N8610, N4793, N7444);
  not ginst2947 (N8615, N7447);
  not ginst2948 (N8616, N7450);
  not ginst2949 (N8617, N7453);
  not ginst2950 (N8618, N7456);
  not ginst2951 (N8619, N7474);
  not ginst2952 (N8624, N7465);
  not ginst2953 (N8625, N7468);
  not ginst2954 (N8626, N7471);
  nand ginst2955 (N8627, N8144, N8145);
  not ginst2956 (N8632, N7479);
  not ginst2957 (N8633, N7482);
  not ginst2958 (N8634, N7485);
  not ginst2959 (N8637, N7491);
  not ginst2960 (N8638, N7494);
  not ginst2961 (N8639, N7497);
  not ginst2962 (N8644, N7503);
  not ginst2963 (N8645, N7506);
  not ginst2964 (N8646, N7509);
  not ginst2965 (N8647, N7512);
  not ginst2966 (N8648, N7530);
  not ginst2967 (N865, N364);
  not ginst2968 (N8653, N7521);
  not ginst2969 (N8654, N7524);
  not ginst2970 (N8655, N7527);
  buf ginst2971 (N8660, N6894);
  buf ginst2972 (N8663, N6894);
  buf ginst2973 (N8666, N6901);
  buf ginst2974 (N8669, N6901);
  buf ginst2975 (N8672, N6912);
  buf ginst2976 (N8675, N6912);
  buf ginst2977 (N8678, N7049);
  buf ginst2978 (N8681, N6988);
  buf ginst2979 (N8684, N6970);
  buf ginst2980 (N8687, N6977);
  buf ginst2981 (N8690, N7049);
  buf ginst2982 (N8693, N6988);
  buf ginst2983 (N8696, N6970);
  buf ginst2984 (N8699, N6977);
  buf ginst2985 (N8702, N7036);
  buf ginst2986 (N8705, N6998);
  buf ginst2987 (N8708, N7020);
  buf ginst2988 (N871, N367);
  buf ginst2989 (N8711, N7006);
  buf ginst2990 (N8714, N7006);
  not ginst2991 (N8717, N7553);
  buf ginst2992 (N8718, N7036);
  buf ginst2993 (N8721, N6998);
  buf ginst2994 (N8724, N7020);
  nand ginst2995 (N8727, N8216, N8217);
  nand ginst2996 (N8730, N8218, N8219);
  not ginst2997 (N8733, N7574);
  not ginst2998 (N8734, N7577);
  buf ginst2999 (N8735, N7107);
  buf ginst3000 (N8738, N7107);
  buf ginst3001 (N8741, N7114);
  buf ginst3002 (N8744, N7114);
  buf ginst3003 (N8747, N7125);
  buf ginst3004 (N8750, N7125);
  not ginst3005 (N8753, N7560);
  not ginst3006 (N8754, N7563);
  not ginst3007 (N8755, N7566);
  not ginst3008 (N8756, N7569);
  buf ginst3009 (N8757, N7301);
  buf ginst3010 (N8760, N7240);
  buf ginst3011 (N8763, N7222);
  buf ginst3012 (N8766, N7229);
  buf ginst3013 (N8769, N7301);
  buf ginst3014 (N8772, N7240);
  buf ginst3015 (N8775, N7222);
  buf ginst3016 (N8778, N7229);
  buf ginst3017 (N8781, N7307);
  buf ginst3018 (N8784, N7288);
  buf ginst3019 (N8787, N7250);
  buf ginst3020 (N8790, N7272);
  buf ginst3021 (N8793, N7258);
  buf ginst3022 (N8796, N7258);
  buf ginst3023 (N8799, N7307);
  buf ginst3024 (N8802, N7288);
  buf ginst3025 (N8805, N7250);
  buf ginst3026 (N8808, N7272);
  nand ginst3027 (N881, N467, N585);
  nand ginst3028 (N8811, N8232, N8233);
  not ginst3029 (N8814, N7588);
  not ginst3030 (N8815, N7591);
  not ginst3031 (N8816, N7582);
  not ginst3032 (N8817, N7585);
  and ginst3033 (N8818, N3155, N7620);
  not ginst3034 (N882, N528);
  not ginst3035 (N883, N578);
  not ginst3036 (N884, N575);
  and ginst3037 (N8840, N3122, N7609);
  not ginst3038 (N885, N494);
  not ginst3039 (N8857, N7609);
  and ginst3040 (N886, N528, N578);
  and ginst3041 (N8861, N5740, N6797, N8274);
  and ginst3042 (N8862, N5736, N6800, N8275);
  and ginst3043 (N8863, N5751, N6803, N8276);
  and ginst3044 (N8864, N5747, N6806, N8277);
  and ginst3045 (N8865, N5762, N6809, N8278);
  and ginst3046 (N8866, N5758, N6812, N8279);
  and ginst3047 (N887, N494, N575);
  not ginst3048 (N8871, N7655);
  and ginst3049 (N8874, N6833, N7655);
  and ginst3050 (N8878, N6867, N7671);
  not ginst3051 (N8879, N8196);
  nand ginst3052 (N8880, N8196, N8315);
  not ginst3053 (N8881, N8200);
  nand ginst3054 (N8882, N8200, N8317);
  not ginst3055 (N8883, N8204);
  nand ginst3056 (N8884, N8204, N8319);
  not ginst3057 (N8885, N8208);
  nand ginst3058 (N8886, N8208, N8321);
  nand ginst3059 (N8887, N3658, N8323);
  nand ginst3060 (N8888, N4817, N8325);
  buf ginst3061 (N889, N590);
  or ginst3062 (N8898, N4544, N8337, N8338, N8339);
  or ginst3063 (N8902, N4562, N8348, N8349, N8350, N8351);
  or ginst3064 (N8920, N4576, N8369, N8370, N8371);
  or ginst3065 (N8924, N4581, N8377);
  or ginst3066 (N8927, N4592, N8378, N8379, N8380, N8381);
  or ginst3067 (N8931, N4603, N8392);
  or ginst3068 (N8943, N7825, N8404);
  or ginst3069 (N8950, N4630, N8409, N8410, N8411);
  or ginst3070 (N8956, N4637, N8415, N8416, N8417, N8418);
  not ginst3071 (N8959, N7852);
  and ginst3072 (N8960, N3375, N7852);
  or ginst3073 (N8963, N4656, N8433, N8434, N8435);
  or ginst3074 (N8966, N4674, N8447, N8448, N8449, N8450);
  and ginst3075 (N8991, N6083, N7188, N8469);
  and ginst3076 (N8992, N6079, N7191, N8470);
  or ginst3077 (N8995, N4701, N8488, N8489, N8490);
  or ginst3078 (N8996, N4706, N8496);
  or ginst3079 (N9001, N4717, N8500, N8501, N8502, N8503);
  or ginst3080 (N9005, N4728, N8516);
  and ginst3081 (N9024, N6141, N7334, N8537);
  and ginst3082 (N9025, N6137, N7337, N8538);
  or ginst3083 (N9029, N4756, N8545, N8546, N8547);
  or ginst3084 (N9035, N4760, N8551, N8552, N8553, N8554);
  and ginst3085 (N9053, N6170, N7378, N8564);
  and ginst3086 (N9054, N6166, N7381, N8565);
  nand ginst3087 (N9064, N4303, N8607);
  nand ginst3088 (N9065, N3507, N8609);
  not ginst3089 (N9066, N8114);
  nand ginst3090 (N9067, N4795, N8114);
  or ginst3091 (N9068, N6783, N7613);
  not ginst3092 (N9071, N8117);
  not ginst3093 (N9072, N8131);
  nand ginst3094 (N9073, N6195, N8131);
  not ginst3095 (N9074, N7613);
  not ginst3096 (N9077, N8134);
  or ginst3097 (N9079, N6865, N7650);
  not ginst3098 (N9082, N8146);
  not ginst3099 (N9083, N7650);
  not ginst3100 (N9086, N8156);
  not ginst3101 (N9087, N8166);
  nand ginst3102 (N9088, N4813, N8166);
  or ginst3103 (N9089, N6866, N7659);
  not ginst3104 (N9092, N8169);
  not ginst3105 (N9093, N8183);
  nand ginst3106 (N9094, N6203, N8183);
  not ginst3107 (N9095, N7659);
  not ginst3108 (N9098, N8186);
  or ginst3109 (N9099, N4545, N8340, N8341, N8342);
  nor ginst3110 (N9103, N4545, N8343, N8344);
  or ginst3111 (N9107, N4549, N8345, N8346);
  nor ginst3112 (N9111, N4549, N8347);
  or ginst3113 (N9117, N4577, N8372, N8373, N8374);
  nor ginst3114 (N9127, N4577, N8375, N8376);
  nor ginst3115 (N9146, N4597, N8390, N8391);
  nor ginst3116 (N9149, N4593, N8385, N8386, N8387);
  nand ginst3117 (N9159, N7577, N8733);
  nand ginst3118 (N9160, N7574, N8734);
  or ginst3119 (N9161, N4657, N8436, N8437, N8438);
  nor ginst3120 (N9165, N4657, N8439, N8440);
  or ginst3121 (N9169, N4661, N8441, N8442);
  nor ginst3122 (N9173, N4661, N8443);
  nand ginst3123 (N9179, N7563, N8753);
  nand ginst3124 (N9180, N7560, N8754);
  nand ginst3125 (N9181, N7569, N8755);
  nand ginst3126 (N9182, N7566, N8756);
  or ginst3127 (N9183, N4702, N8491, N8492, N8493);
  nor ginst3128 (N9193, N4702, N8494, N8495);
  or ginst3129 (N9203, N4722, N8511, N8512, N8513);
  or ginst3130 (N9206, N4718, N8504, N8505, N8506, N8507);
  nor ginst3131 (N9220, N4722, N8514, N8515);
  nor ginst3132 (N9223, N4718, N8508, N8509, N8510);
  nand ginst3133 (N9234, N7591, N8814);
  nand ginst3134 (N9235, N7588, N8815);
  nand ginst3135 (N9236, N7585, N8816);
  nand ginst3136 (N9237, N7582, N8817);
  or ginst3137 (N9238, N3159, N8818);
  or ginst3138 (N9242, N3126, N8840);
  nand ginst3139 (N9243, N8324, N8888);
  not ginst3140 (N9244, N8580);
  not ginst3141 (N9245, N8583);
  not ginst3142 (N9246, N8586);
  not ginst3143 (N9247, N8589);
  not ginst3144 (N9248, N8592);
  not ginst3145 (N9249, N8595);
  not ginst3146 (N9250, N8598);
  not ginst3147 (N9251, N8601);
  not ginst3148 (N9252, N8604);
  nor ginst3149 (N9256, N8280, N8861);
  nor ginst3150 (N9257, N8281, N8862);
  nor ginst3151 (N9258, N8282, N8863);
  nor ginst3152 (N9259, N8283, N8864);
  nor ginst3153 (N9260, N8284, N8865);
  nor ginst3154 (N9261, N8285, N8866);
  not ginst3155 (N9262, N8627);
  or ginst3156 (N9265, N7649, N8874);
  or ginst3157 (N9268, N7668, N8878);
  nand ginst3158 (N9271, N7533, N8879);
  nand ginst3159 (N9272, N7536, N8881);
  nand ginst3160 (N9273, N7539, N8883);
  nand ginst3161 (N9274, N7542, N8885);
  nand ginst3162 (N9275, N8322, N8887);
  not ginst3163 (N9276, N8333);
  and ginst3164 (N9280, N6929, N6936, N6946, N6957, N8326);
  and ginst3165 (N9285, N367, N6936, N6946, N6957, N8326);
  and ginst3166 (N9286, N367, N6946, N6957, N8326);
  and ginst3167 (N9287, N367, N6957, N8326);
  and ginst3168 (N9288, N367, N8326);
  not ginst3169 (N9290, N8660);
  not ginst3170 (N9292, N8663);
  not ginst3171 (N9294, N8666);
  not ginst3172 (N9296, N8669);
  nand ginst3173 (N9297, N5966, N8672);
  not ginst3174 (N9298, N8672);
  nand ginst3175 (N9299, N6969, N8675);
  not ginst3176 (N9300, N8675);
  not ginst3177 (N9301, N8365);
  and ginst3178 (N9307, N6998, N7006, N7020, N7036, N8358);
  and ginst3179 (N9314, N7006, N7020, N7036, N8358);
  and ginst3180 (N9315, N7020, N7036, N8358);
  and ginst3181 (N9318, N7036, N8358);
  not ginst3182 (N9319, N8687);
  not ginst3183 (N9320, N8699);
  not ginst3184 (N9321, N8711);
  not ginst3185 (N9322, N8714);
  not ginst3186 (N9323, N8727);
  not ginst3187 (N9324, N8730);
  not ginst3188 (N9326, N8405);
  and ginst3189 (N9332, N8405, N8412);
  or ginst3190 (N9339, N4193, N8960);
  and ginst3191 (N9344, N8430, N8444);
  not ginst3192 (N9352, N8735);
  not ginst3193 (N9354, N8738);
  not ginst3194 (N9356, N8741);
  not ginst3195 (N9358, N8744);
  nand ginst3196 (N9359, N6078, N8747);
  not ginst3197 (N9360, N8747);
  nand ginst3198 (N9361, N7187, N8750);
  not ginst3199 (N9362, N8750);
  not ginst3200 (N9363, N8471);
  not ginst3201 (N9364, N8474);
  not ginst3202 (N9365, N8477);
  not ginst3203 (N9366, N8480);
  nor ginst3204 (N9367, N8483, N8991);
  nor ginst3205 (N9368, N8484, N8992);
  and ginst3206 (N9369, N7194, N7198, N8471);
  and ginst3207 (N9370, N8457, N8460, N8474);
  and ginst3208 (N9371, N7205, N7209, N8477);
  and ginst3209 (N9372, N8463, N8466, N8480);
  not ginst3210 (N9375, N8497);
  not ginst3211 (N9381, N8766);
  not ginst3212 (N9382, N8778);
  not ginst3213 (N9383, N8793);
  not ginst3214 (N9384, N8796);
  and ginst3215 (N9385, N8485, N8497);
  not ginst3216 (N9392, N8525);
  not ginst3217 (N9393, N8528);
  not ginst3218 (N9394, N8531);
  not ginst3219 (N9395, N8534);
  and ginst3220 (N9396, N7314, N7318, N8525);
  and ginst3221 (N9397, N8519, N8522, N8528);
  and ginst3222 (N9398, N6127, N6131, N8531);
  and ginst3223 (N9399, N7325, N7328, N8534);
  nor ginst3224 (N9400, N8539, N9024);
  nor ginst3225 (N9401, N8540, N9025);
  not ginst3226 (N9402, N8541);
  nand ginst3227 (N9407, N89, N8548);
  and ginst3228 (N9408, N8541, N8548);
  not ginst3229 (N9412, N8811);
  not ginst3230 (N9413, N8566);
  not ginst3231 (N9414, N8569);
  not ginst3232 (N9415, N8572);
  not ginst3233 (N9416, N8575);
  nor ginst3234 (N9417, N8578, N9053);
  nor ginst3235 (N9418, N8579, N9054);
  and ginst3236 (N9419, N6177, N7387, N8566);
  and ginst3237 (N9420, N7384, N8555, N8569);
  and ginst3238 (N9421, N7394, N7398, N8572);
  and ginst3239 (N9422, N8558, N8561, N8575);
  buf ginst3240 (N9423, N8326);
  nand ginst3241 (N9426, N8608, N9064);
  nand ginst3242 (N9429, N8610, N9065);
  nand ginst3243 (N9432, N3515, N9066);
  nand ginst3244 (N9435, N4796, N9072);
  nand ginst3245 (N9442, N3628, N9087);
  nand ginst3246 (N9445, N4814, N9093);
  buf ginst3247 (N945, N657);
  not ginst3248 (N9454, N8678);
  not ginst3249 (N9455, N8681);
  not ginst3250 (N9456, N8684);
  not ginst3251 (N9459, N8690);
  not ginst3252 (N9460, N8693);
  not ginst3253 (N9461, N8696);
  buf ginst3254 (N9462, N8358);
  not ginst3255 (N9465, N8702);
  not ginst3256 (N9466, N8705);
  not ginst3257 (N9467, N8708);
  not ginst3258 (N9468, N8724);
  buf ginst3259 (N9473, N8358);
  not ginst3260 (N9476, N8718);
  not ginst3261 (N9477, N8721);
  nand ginst3262 (N9478, N9159, N9160);
  nand ginst3263 (N9485, N9179, N9180);
  nand ginst3264 (N9488, N9181, N9182);
  not ginst3265 (N9493, N8757);
  not ginst3266 (N9494, N8760);
  not ginst3267 (N9495, N8763);
  not ginst3268 (N9498, N8769);
  not ginst3269 (N9499, N8772);
  not ginst3270 (N9500, N8775);
  not ginst3271 (N9505, N8781);
  not ginst3272 (N9506, N8784);
  not ginst3273 (N9507, N8787);
  not ginst3274 (N9508, N8790);
  not ginst3275 (N9509, N8808);
  not ginst3276 (N9514, N8799);
  not ginst3277 (N9515, N8802);
  not ginst3278 (N9516, N8805);
  nand ginst3279 (N9517, N9234, N9235);
  nand ginst3280 (N9520, N9236, N9237);
  and ginst3281 (N9526, N8421, N8943);
  and ginst3282 (N9531, N8421, N8943);
  nand ginst3283 (N9539, N8880, N9271);
  nand ginst3284 (N9540, N8884, N9273);
  not ginst3285 (N9541, N9275);
  and ginst3286 (N9543, N8254, N8857);
  and ginst3287 (N9551, N8288, N8871);
  nand ginst3288 (N9555, N8882, N9272);
  nand ginst3289 (N9556, N8886, N9274);
  not ginst3290 (N9557, N8898);
  and ginst3291 (N9560, N8333, N8902);
  not ginst3292 (N9561, N9099);
  nand ginst3293 (N9562, N9099, N9290);
  not ginst3294 (N9563, N9103);
  nand ginst3295 (N9564, N9103, N9292);
  not ginst3296 (N9565, N9107);
  nand ginst3297 (N9566, N9107, N9294);
  not ginst3298 (N9567, N9111);
  nand ginst3299 (N9568, N9111, N9296);
  nand ginst3300 (N9569, N4844, N9298);
  not ginst3301 (N957, N688);
  nand ginst3302 (N9570, N6207, N9300);
  not ginst3303 (N9571, N8920);
  not ginst3304 (N9575, N8927);
  and ginst3305 (N9579, N8365, N8927);
  not ginst3306 (N9581, N8950);
  not ginst3307 (N9582, N8956);
  and ginst3308 (N9585, N8405, N8956);
  and ginst3309 (N9591, N8430, N8966);
  not ginst3310 (N9592, N9161);
  nand ginst3311 (N9593, N9161, N9352);
  not ginst3312 (N9594, N9165);
  nand ginst3313 (N9595, N9165, N9354);
  not ginst3314 (N9596, N9169);
  nand ginst3315 (N9597, N9169, N9356);
  not ginst3316 (N9598, N9173);
  nand ginst3317 (N9599, N9173, N9358);
  nand ginst3318 (N9600, N4940, N9360);
  nand ginst3319 (N9601, N6220, N9362);
  and ginst3320 (N9602, N7198, N8457, N9363);
  and ginst3321 (N9603, N7194, N8460, N9364);
  and ginst3322 (N9604, N7209, N8463, N9365);
  and ginst3323 (N9605, N7205, N8466, N9366);
  not ginst3324 (N9608, N9001);
  and ginst3325 (N9611, N8485, N9001);
  and ginst3326 (N9612, N7318, N8519, N9392);
  and ginst3327 (N9613, N7314, N8522, N9393);
  and ginst3328 (N9614, N6131, N7325, N9394);
  and ginst3329 (N9615, N6127, N7328, N9395);
  not ginst3330 (N9616, N9029);
  not ginst3331 (N9617, N9035);
  and ginst3332 (N9618, N8541, N9035);
  and ginst3333 (N9621, N7384, N7387, N9413);
  and ginst3334 (N9622, N6177, N8555, N9414);
  and ginst3335 (N9623, N7398, N8558, N9415);
  and ginst3336 (N9624, N7394, N8561, N9416);
  or ginst3337 (N9626, N4563, N8352, N8353, N8354, N9285);
  or ginst3338 (N9629, N4566, N8355, N8356, N9286);
  or ginst3339 (N9632, N4570, N8357, N9287);
  or ginst3340 (N9635, N5960, N9288);
  nand ginst3341 (N9642, N9067, N9432);
  not ginst3342 (N9645, N9068);
  nand ginst3343 (N9646, N9073, N9435);
  not ginst3344 (N9649, N9074);
  nand ginst3345 (N9650, N9256, N9257);
  nand ginst3346 (N9653, N9258, N9259);
  nand ginst3347 (N9656, N9260, N9261);
  not ginst3348 (N9659, N9079);
  nand ginst3349 (N9660, N4809, N9079);
  not ginst3350 (N9661, N9083);
  nand ginst3351 (N9662, N6202, N9083);
  nand ginst3352 (N9663, N9088, N9442);
  not ginst3353 (N9666, N9089);
  nand ginst3354 (N9667, N9094, N9445);
  not ginst3355 (N9670, N9095);
  or ginst3356 (N9671, N8393, N8924);
  not ginst3357 (N9674, N9117);
  not ginst3358 (N9675, N8924);
  not ginst3359 (N9678, N9127);
  or ginst3360 (N9679, N4597, N8388, N8389, N9315);
  or ginst3361 (N9682, N8931, N9318);
  or ginst3362 (N9685, N4593, N8382, N8383, N8384, N9314);
  not ginst3363 (N9690, N9146);
  nand ginst3364 (N9691, N8717, N9146);
  not ginst3365 (N9692, N8931);
  not ginst3366 (N9695, N9149);
  nand ginst3367 (N9698, N9400, N9401);
  nand ginst3368 (N9702, N9367, N9368);
  or ginst3369 (N9707, N8517, N8996);
  not ginst3370 (N9710, N9183);
  not ginst3371 (N9711, N8996);
  not ginst3372 (N9714, N9193);
  not ginst3373 (N9715, N9203);
  nand ginst3374 (N9716, N6235, N9203);
  or ginst3375 (N9717, N8518, N9005);
  not ginst3376 (N9720, N9206);
  not ginst3377 (N9721, N9220);
  nand ginst3378 (N9722, N7573, N9220);
  not ginst3379 (N9723, N9005);
  not ginst3380 (N9726, N9223);
  nand ginst3381 (N9727, N9417, N9418);
  and ginst3382 (N9732, N8269, N9268);
  nand ginst3383 (N9733, N9326, N9581);
  and ginst3384 (N9734, N89, N8394, N8421, N9332, N9408);
  and ginst3385 (N9735, N89, N8394, N8421, N9332, N9408);
  and ginst3386 (N9736, N8262, N9265);
  not ginst3387 (N9737, N9555);
  not ginst3388 (N9738, N9556);
  nand ginst3389 (N9739, N9361, N9601);
  nand ginst3390 (N9740, N1115, N9423);
  not ginst3391 (N9741, N9423);
  nand ginst3392 (N9742, N9299, N9570);
  and ginst3393 (N9754, N8333, N9280);
  or ginst3394 (N9758, N8898, N9560);
  nand ginst3395 (N9762, N8660, N9561);
  nand ginst3396 (N9763, N8663, N9563);
  nand ginst3397 (N9764, N8666, N9565);
  nand ginst3398 (N9765, N8669, N9567);
  nand ginst3399 (N9766, N9297, N9569);
  and ginst3400 (N9767, N367, N9280);
  nand ginst3401 (N9768, N9276, N9557);
  not ginst3402 (N9769, N9307);
  nand ginst3403 (N9773, N367, N9307);
  nand ginst3404 (N9774, N9301, N9571);
  and ginst3405 (N9775, N8365, N9307);
  or ginst3406 (N9779, N8920, N9579);
  not ginst3407 (N9784, N9478);
  nand ginst3408 (N9785, N9402, N9616);
  or ginst3409 (N9786, N8950, N9585);
  and ginst3410 (N9790, N89, N8394, N9332, N9408);
  or ginst3411 (N9791, N8963, N9591);
  nand ginst3412 (N9795, N8735, N9592);
  nand ginst3413 (N9796, N8738, N9594);
  nand ginst3414 (N9797, N8741, N9596);
  nand ginst3415 (N9798, N8744, N9598);
  nand ginst3416 (N9799, N9359, N9600);
  nor ginst3417 (N9800, N9369, N9602);
  nor ginst3418 (N9801, N9370, N9603);
  nor ginst3419 (N9802, N9371, N9604);
  nor ginst3420 (N9803, N9372, N9605);
  not ginst3421 (N9805, N9485);
  not ginst3422 (N9806, N9488);
  or ginst3423 (N9809, N8995, N9611);
  nor ginst3424 (N9813, N9396, N9612);
  nor ginst3425 (N9814, N9397, N9613);
  nor ginst3426 (N9815, N9398, N9614);
  nor ginst3427 (N9816, N9399, N9615);
  and ginst3428 (N9817, N9407, N9617);
  or ginst3429 (N9820, N9029, N9618);
  not ginst3430 (N9825, N9517);
  not ginst3431 (N9826, N9520);
  nor ginst3432 (N9827, N9419, N9621);
  nor ginst3433 (N9828, N9420, N9622);
  nor ginst3434 (N9829, N9421, N9623);
  nor ginst3435 (N9830, N9422, N9624);
  not ginst3436 (N9835, N9426);
  nand ginst3437 (N9836, N4789, N9426);
  not ginst3438 (N9837, N9429);
  nand ginst3439 (N9838, N4794, N9429);
  nand ginst3440 (N9846, N3625, N9659);
  nand ginst3441 (N9847, N4810, N9661);
  not ginst3442 (N9862, N9462);
  nand ginst3443 (N9863, N7553, N9690);
  not ginst3444 (N9866, N9473);
  nand ginst3445 (N9873, N5030, N9715);
  nand ginst3446 (N9876, N6236, N9721);
  nand ginst3447 (N9890, N9593, N9795);
  nand ginst3448 (N9891, N9597, N9797);
  not ginst3449 (N9892, N9799);
  nand ginst3450 (N9893, N871, N9741);
  nand ginst3451 (N9894, N9562, N9762);
  nand ginst3452 (N9895, N9566, N9764);
  not ginst3453 (N9896, N9766);
  not ginst3454 (N9897, N9626);
  nand ginst3455 (N9898, N9249, N9626);
  not ginst3456 (N9899, N9629);
  nand ginst3457 (N9900, N9250, N9629);
  not ginst3458 (N9901, N9632);
  nand ginst3459 (N9902, N9251, N9632);
  not ginst3460 (N9903, N9635);
  nand ginst3461 (N9904, N9252, N9635);
  not ginst3462 (N9905, N9543);
  not ginst3463 (N9906, N9650);
  nand ginst3464 (N9907, N5769, N9650);
  not ginst3465 (N9908, N9653);
  nand ginst3466 (N9909, N5770, N9653);
  not ginst3467 (N9910, N9656);
  nand ginst3468 (N9911, N9262, N9656);
  not ginst3469 (N9917, N9551);
  nand ginst3470 (N9923, N9564, N9763);
  nand ginst3471 (N9924, N9568, N9765);
  or ginst3472 (N9925, N8902, N9767);
  and ginst3473 (N9932, N9575, N9773);
  and ginst3474 (N9935, N9575, N9769);
  not ginst3475 (N9938, N9698);
  nand ginst3476 (N9939, N9323, N9698);
  nand ginst3477 (N9945, N9595, N9796);
  nand ginst3478 (N9946, N9599, N9798);
  not ginst3479 (N9947, N9702);
  nand ginst3480 (N9948, N6102, N9702);
  and ginst3481 (N9949, N9375, N9608);
  not ginst3482 (N9953, N9727);
  nand ginst3483 (N9954, N9412, N9727);
  nand ginst3484 (N9955, N3502, N9835);
  nand ginst3485 (N9956, N3510, N9837);
  not ginst3486 (N9957, N9642);
  nand ginst3487 (N9958, N9642, N9645);
  not ginst3488 (N9959, N9646);
  nand ginst3489 (N9960, N9646, N9649);
  nand ginst3490 (N9961, N9660, N9846);
  nand ginst3491 (N9964, N9662, N9847);
  not ginst3492 (N9967, N9663);
  nand ginst3493 (N9968, N9663, N9666);
  not ginst3494 (N9969, N9667);
  nand ginst3495 (N9970, N9667, N9670);
  not ginst3496 (N9971, N9671);
  nand ginst3497 (N9972, N6213, N9671);
  not ginst3498 (N9973, N9675);
  nand ginst3499 (N9974, N7551, N9675);
  not ginst3500 (N9975, N9679);
  nand ginst3501 (N9976, N7552, N9679);
  not ginst3502 (N9977, N9682);
  not ginst3503 (N9978, N9685);
  nand ginst3504 (N9979, N9691, N9863);
  not ginst3505 (N9982, N9692);
  nand ginst3506 (N9983, N9813, N9814);
  nand ginst3507 (N9986, N9815, N9816);
  nand ginst3508 (N9989, N9800, N9801);
  nand ginst3509 (N9992, N9802, N9803);
  not ginst3510 (N9995, N9707);
  nand ginst3511 (N9996, N6231, N9707);
  not ginst3512 (N9997, N9711);
  nand ginst3513 (N9998, N7572, N9711);
  nand ginst3514 (N9999, N9716, N9873);

endmodule

/*************** SatHard block ***************/
module SatHard (N29, N159, N325, N331, N158, N277, N299, N303, keyinput0, keyinput1, keyinput2, keyinput3, keyinput4, keyinput5, keyinput6, keyinput7, keyinput8, keyinput9, keyinput10, keyinput11, keyinput12, keyinput13, keyinput14, keyinput15, flip_signal);

  input N29, N159, N325, N331, N158, N277, N299, N303, keyinput0, keyinput1, keyinput2, keyinput3, keyinput4, keyinput5, keyinput6, keyinput7, keyinput8, keyinput9, keyinput10, keyinput11, keyinput12, keyinput13, keyinput14, keyinput15;
  output flip_signal;
  //SatHard key=1001100010101011
  wire [7:0] sat_res_inputs;
  wire [15:0] keyinputs, keyvalue;
  assign sat_res_inputs[7:0] = {N29, N159, N325, N331, N158, N277, N299, N303};
  assign keyinputs[15:0] = {keyinput0, keyinput1, keyinput2, keyinput3, keyinput4, keyinput5, keyinput6, keyinput7, keyinput8, keyinput9, keyinput10, keyinput11, keyinput12, keyinput13, keyinput14, keyinput15};
  assign keyvalue[15:0] = 16'b1001100010101011;

  wire g, g_bar;
  assign g = &(keyinputs[7:0] ^ sat_res_inputs ^ keyvalue[7:0]);
  assign g_bar = ~&(keyinputs[15:8] ^ sat_res_inputs ^ keyvalue[15:8]);
  assign flip_signal = g & g_bar;

endmodule
/*************** SatHard block ***************/
