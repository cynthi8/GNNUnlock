//key=0110110100101000
// Main module
module c5315_AntiSAT_16_0(i_1, i_4, i_11, i_14, i_17, i_20, i_23, i_24, i_25, i_26, i_27, i_31, i_34, i_37, i_40, i_43, i_46, i_49, i_52, i_53, i_54, i_61, i_64, i_67, i_70, i_73, i_76, i_79, i_80, i_81, i_82, i_83, i_86, i_87, i_88, i_91, i_94, i_97, i_100, i_103, i_106, i_109, i_112, i_113, i_114, i_115, i_116, i_117, i_118, i_119, i_120, i_121, i_122, i_123, i_126, i_127, i_128, i_129, i_130, i_131, i_132, i_135, i_136, i_137, i_140, i_141, i_145, i_146, i_149, i_152, i_155, i_158, i_161, i_164, i_167, i_170, i_173, i_176, i_179, i_182, i_185, i_188, i_191, i_194, i_197, i_200, i_203, i_206, i_209, i_210, i_217, i_218, i_225, i_226, i_233, i_234, i_241, i_242, i_245, i_248, i_251, i_254, i_257, i_264, i_265, i_272, i_273, i_280, i_281, i_288, i_289, i_292, i_293, i_299, i_302, i_307, i_308, i_315, i_316, i_323, i_324, i_331, i_332, i_335, i_338, i_341, i_348, i_351, i_358, i_361, i_366, i_369, i_372, i_373, i_374, i_386, i_389, i_400, i_411, i_422, i_435, i_446, i_457, i_468, i_479, i_490, i_503, i_514, i_523, i_534, i_545, i_549, i_552, i_556, i_559, i_562, i_566, i_571, i_574, i_577, i_580, i_583, i_588, i_591, i_592, i_595, i_596, i_597, i_598, i_599, i_603, i_607, i_610, i_613, i_616, i_619, i_625, i_631, keyinput0, keyinput1, keyinput2, keyinput3, keyinput4, keyinput5, keyinput6, keyinput7, keyinput8, keyinput9, keyinput10, keyinput11, keyinput12, keyinput13, keyinput14, keyinput15, i_709, i_816, i_1066, i_1137, i_1138, i_1139, i_1140, i_1141, i_1142, i_1143, i_1144, i_1145, i_1147, i_1152, i_1153, i_1154, i_1155, i_1972, i_2054, i_2060, i_2061, i_2139, i_2142, i_2309, i_2387, i_2527, i_2584, i_2590, i_2623, i_3357, i_3358, i_3359, i_3360, i_3604, i_3613, i_4272, i_4275, i_4278, i_4279, i_4737, i_4738, i_4739, i_4740, i_5240, i_5388, i_6641, i_6643, i_6646, i_6648, i_6716, i_6877, i_6924, i_6925, i_6926, i_6927, i_7015, i_7363, i_7365, i_7432, i_7449, i_7465, i_7466, i_7467, i_7469, i_7470, i_7471, i_7472, i_7473, i_7474, i_7476, i_7503, i_7504, i_7506, i_7511, i_7515, i_7516, i_7517, i_7518, i_7519, i_7520, i_7521, i_7522, i_7600, i_7601, i_7602, i_7603, i_7604, i_7605, i_7606, i_7607, i_7626, i_7698, i_7699, i_7700, i_7701, i_7702, i_7703, i_7704, i_7705, i_7706, i_7707, i_7735, i_7736, i_7737, i_7738, i_7739, i_7740, i_7741, i_7742, i_7754, i_7755, i_7756, i_7757, i_7758, i_7759, i_7760, i_7761, i_8075, i_8076, i_8123, i_8124, i_8127, i_8128);

  input i_1, i_4, i_11, i_14, i_17, i_20, i_23, i_24, i_25, i_26, i_27, i_31, i_34, i_37, i_40, i_43, i_46, i_49, i_52, i_53, i_54, i_61, i_64, i_67, i_70, i_73, i_76, i_79, i_80, i_81, i_82, i_83, i_86, i_87, i_88, i_91, i_94, i_97, i_100, i_103, i_106, i_109, i_112, i_113, i_114, i_115, i_116, i_117, i_118, i_119, i_120, i_121, i_122, i_123, i_126, i_127, i_128, i_129, i_130, i_131, i_132, i_135, i_136, i_137, i_140, i_141, i_145, i_146, i_149, i_152, i_155, i_158, i_161, i_164, i_167, i_170, i_173, i_176, i_179, i_182, i_185, i_188, i_191, i_194, i_197, i_200, i_203, i_206, i_209, i_210, i_217, i_218, i_225, i_226, i_233, i_234, i_241, i_242, i_245, i_248, i_251, i_254, i_257, i_264, i_265, i_272, i_273, i_280, i_281, i_288, i_289, i_292, i_293, i_299, i_302, i_307, i_308, i_315, i_316, i_323, i_324, i_331, i_332, i_335, i_338, i_341, i_348, i_351, i_358, i_361, i_366, i_369, i_372, i_373, i_374, i_386, i_389, i_400, i_411, i_422, i_435, i_446, i_457, i_468, i_479, i_490, i_503, i_514, i_523, i_534, i_545, i_549, i_552, i_556, i_559, i_562, i_566, i_571, i_574, i_577, i_580, i_583, i_588, i_591, i_592, i_595, i_596, i_597, i_598, i_599, i_603, i_607, i_610, i_613, i_616, i_619, i_625, i_631, keyinput0, keyinput1, keyinput2, keyinput3, keyinput4, keyinput5, keyinput6, keyinput7, keyinput8, keyinput9, keyinput10, keyinput11, keyinput12, keyinput13, keyinput14, keyinput15;
  output i_709, i_816, i_1066, i_1137, i_1138, i_1139, i_1140, i_1141, i_1142, i_1143, i_1144, i_1145, i_1147, i_1152, i_1153, i_1154, i_1155, i_1972, i_2054, i_2060, i_2061, i_2139, i_2142, i_2309, i_2387, i_2527, i_2584, i_2590, i_2623, i_3357, i_3358, i_3359, i_3360, i_3604, i_3613, i_4272, i_4275, i_4278, i_4279, i_4737, i_4738, i_4739, i_4740, i_5240, i_5388, i_6641, i_6643, i_6646, i_6648, i_6716, i_6877, i_6924, i_6925, i_6926, i_6927, i_7015, i_7363, i_7365, i_7432, i_7449, i_7465, i_7466, i_7467, i_7469, i_7470, i_7471, i_7472, i_7473, i_7474, i_7476, i_7503, i_7504, i_7506, i_7511, i_7515, i_7516, i_7517, i_7518, i_7519, i_7520, i_7521, i_7522, i_7600, i_7601, i_7602, i_7603, i_7604, i_7605, i_7606, i_7607, i_7626, i_7698, i_7699, i_7700, i_7701, i_7702, i_7703, i_7704, i_7705, i_7706, i_7707, i_7735, i_7736, i_7737, i_7738, i_7739, i_7740, i_7741, i_7742, i_7754, i_7755, i_7756, i_7757, i_7758, i_7759, i_7760, i_7761, i_8075, i_8076, i_8123, i_8124, i_8127, i_8128;
  wire i_1042, i_1043, i_1067, i_1080, i_1092, i_1104, i_1146, i_1148, i_1149, i_1150, i_1151, i_1156, i_1157, i_1161, i_1173, i_1185, i_1197, i_1209, i_1213, i_1216, i_1219, i_1223, i_1235, i_1247, i_1259, i_1271, i_1280, i_1292, i_1303, i_1315, i_1327, i_1339, i_1351, i_1363, i_1375, i_1378, i_1381, i_1384, i_1387, i_1390, i_1393, i_1396, i_1415, i_1418, i_1421, i_1424, i_1427, i_1430, i_1433, i_1436, i_1455, i_1462, i_1469, i_1475, i_1479, i_1482, i_1492, i_1495, i_1498, i_1501, i_1504, i_1507, i_1510, i_1513, i_1516, i_1519, i_1522, i_1525, i_1542, i_1545, i_1548, i_1551, i_1554, i_1557, i_1560, i_1563, i_1566, i_1573, i_1580, i_1583, i_1588, i_1594, i_1597, i_1600, i_1603, i_1606, i_1609, i_1612, i_1615, i_1618, i_1621, i_1624, i_1627, i_1630, i_1633, i_1636, i_1639, i_1642, i_1645, i_1648, i_1651, i_1654, i_1657, i_1660, i_1663, i_1675, i_1685, i_1697, i_1709, i_1721, i_1727, i_1731, i_1743, i_1755, i_1758, i_1761, i_1769, i_1777, i_1785, i_1793, i_1800, i_1807, i_1814, i_1821, i_1824, i_1827, i_1830, i_1833, i_1836, i_1839, i_1842, i_1845, i_1848, i_1851, i_1854, i_1857, i_1860, i_1863, i_1866, i_1869, i_1872, i_1875, i_1878, i_1881, i_1884, i_1887, i_1890, i_1893, i_1896, i_1899, i_1902, i_1905, i_1908, i_1911, i_1914, i_1917, i_1920, i_1923, i_1926, i_1929, i_1932, i_1935, i_1938, i_1941, i_1944, i_1947, i_1950, i_1953, i_1956, i_1959, i_1962, i_1965, i_1968, i_2349, i_2350, i_2585, i_2586, i_2587, i_2588, i_2589, i_2591, i_2592, i_2593, i_2594, i_2595, i_2596, i_2597, i_2598, i_2599, i_2600, i_2601, i_2602, i_2603, i_2604, i_2605, i_2606, i_2607, i_2608, i_2609, i_2610, i_2611, i_2612, i_2613, i_2614, i_2615, i_2616, i_2617, i_2618, i_2619, i_2620, i_2621, i_2622, i_2624, i_2625, i_2626, i_2627, i_2628, i_2629, i_2630, i_2631, i_2632, i_2633, i_2634, i_2635, i_2636, i_2637, i_2638, i_2639, i_2640, i_2641, i_2642, i_2643, i_2644, i_2645, i_2646, i_2647, i_2653, i_2664, i_2675, i_2681, i_2692, i_2703, i_2704, i_2709, i_2710, i_2711, i_2712, i_2713, i_2714, i_2715, i_2716, i_2717, i_2718, i_2719, i_2720, i_2721, i_2722, i_2728, i_2739, i_2750, i_2756, i_2767, i_2778, i_2779, i_2790, i_2801, i_2812, i_2823, i_2824, i_2825, i_2826, i_2827, i_2828, i_2829, i_2830, i_2831, i_2832, i_2833, i_2834, i_2835, i_2836, i_2837, i_2838, i_2839, i_2840, i_2841, i_2842, i_2843, i_2844, i_2845, i_2846, i_2847, i_2848, i_2849, i_2850, i_2851, i_2852, i_2853, i_2854, i_2855, i_2861, i_2867, i_2868, i_2869, i_2870, i_2871, i_2872, i_2873, i_2874, i_2875, i_2876, i_2877, i_2882, i_2891, i_2901, i_2902, i_2903, i_2904, i_2905, i_2906, i_2907, i_2908, i_2909, i_2910, i_2911, i_2912, i_2913, i_2914, i_2915, i_2916, i_2917, i_2918, i_2919, i_2920, i_2921, i_2922, i_2923, i_2924, i_2925, i_2926, i_2927, i_2928, i_2929, i_2930, i_2931, i_2932, i_2933, i_2934, i_2935, i_2936, i_2937, i_2938, i_2939, i_2940, i_2941, i_2942, i_2948, i_2954, i_2955, i_2956, i_2957, i_2958, i_2959, i_2960, i_2961, i_2962, i_2963, i_2964, i_2969, i_2970, i_2971, i_2972, i_2973, i_2974, i_2975, i_2976, i_2977, i_2978, i_2979, i_2980, i_2981, i_2982, i_2983, i_2984, i_2985, i_2986, i_2987, i_2988, i_2989, i_2990, i_2991, i_2992, i_2993, i_2994, i_2995, i_2996, i_2997, i_2998, i_2999, i_3000, i_3003, i_3006, i_3007, i_3010, i_3013, i_3014, i_3015, i_3016, i_3017, i_3018, i_3019, i_3020, i_3021, i_3022, i_3023, i_3024, i_3025, i_3026, i_3027, i_3028, i_3029, i_3030, i_3031, i_3032, i_3033, i_3034, i_3035, i_3038, i_3041, i_3052, i_3063, i_3068, i_3071, i_3072, i_3073, i_3074, i_3075, i_3086, i_3097, i_3108, i_3119, i_3130, i_3141, i_3142, i_3143, i_3144, i_3145, i_3146, i_3147, i_3158, i_3169, i_3180, i_3191, i_3194, i_3195, i_3196, i_3197, i_3198, i_3199, i_3200, i_3203, i_3401, i_3402, i_3403, i_3404, i_3405, i_3406, i_3407, i_3408, i_3409, i_3410, i_3411, i_3412, i_3413, i_3414, i_3415, i_3416, i_3444, i_3445, i_3446, i_3447, i_3448, i_3449, i_3450, i_3451, i_3452, i_3453, i_3454, i_3455, i_3456, i_3459, i_3460, i_3461, i_3462, i_3463, i_3464, i_3465, i_3466, i_3481, i_3482, i_3483, i_3484, i_3485, i_3486, i_3487, i_3488, i_3489, i_3490, i_3491, i_3492, i_3493, i_3502, i_3503, i_3504, i_3505, i_3506, i_3507, i_3508, i_3509, i_3510, i_3511, i_3512, i_3513, i_3514, i_3515, i_3558, i_3559, i_3560, i_3561, i_3562, i_3563, i_3605, i_3606, i_3607, i_3608, i_3609, i_3610, i_3614, i_3615, i_3616, i_3617, i_3618, i_3619, i_3620, i_3621, i_3622, i_3623, i_3624, i_3625, i_3626, i_3627, i_3628, i_3629, i_3630, i_3631, i_3632, i_3633, i_3634, i_3635, i_3636, i_3637, i_3638, i_3639, i_3640, i_3641, i_3642, i_3643, i_3644, i_3645, i_3646, i_3647, i_3648, i_3649, i_3650, i_3651, i_3652, i_3653, i_3654, i_3655, i_3656, i_3657, i_3658, i_3659, i_3660, i_3661, i_3662, i_3663, i_3664, i_3665, i_3666, i_3667, i_3668, i_3669, i_3670, i_3671, i_3672, i_3673, i_3674, i_3675, i_3676, i_3677, i_3678, i_3679, i_3680, i_3681, i_3682, i_3683, i_3684, i_3685, i_3686, i_3687, i_3688, i_3689, i_3691, i_3700, i_3701, i_3702, i_3703, i_3704, i_3705, i_3708, i_3709, i_3710, i_3711, i_3712, i_3713, i_3715, i_3716, i_3717, i_3718, i_3719, i_3720, i_3721, i_3722, i_3723, i_3724, i_3725, i_3726, i_3727, i_3728, i_3729, i_3730, i_3731, i_3732, i_3738, i_3739, i_3740, i_3741, i_3742, i_3743, i_3744, i_3745, i_3746, i_3747, i_3748, i_3749, i_3750, i_3751, i_3752, i_3753, i_3754, i_3755, i_3756, i_3757, i_3758, i_3759, i_3760, i_3761, i_3762, i_3763, i_3764, i_3765, i_3766, i_3767, i_3768, i_3769, i_3770, i_3771, i_3775, i_3779, i_3780, i_3781, i_3782, i_3783, i_3784, i_3785, i_3786, i_3787, i_3788, i_3789, i_3793, i_3797, i_3800, i_3801, i_3802, i_3803, i_3804, i_3805, i_3806, i_3807, i_3808, i_3809, i_3810, i_3813, i_3816, i_3819, i_3822, i_3823, i_3824, i_3827, i_3828, i_3829, i_3830, i_3831, i_3834, i_3835, i_3836, i_3837, i_3838, i_3839, i_3840, i_3841, i_3842, i_3849, i_3855, i_3861, i_3867, i_3873, i_3881, i_3887, i_3893, i_3908, i_3909, i_3911, i_3914, i_3915, i_3916, i_3917, i_3918, i_3919, i_3920, i_3921, i_3927, i_3933, i_3942, i_3948, i_3956, i_3962, i_3968, i_3975, i_3976, i_3977, i_3978, i_3979, i_3980, i_3981, i_3982, i_3983, i_3984, i_3987, i_3988, i_3989, i_3990, i_3991, i_3998, i_4008, i_4011, i_4021, i_4024, i_4027, i_4031, i_4032, i_4033, i_4034, i_4035, i_4036, i_4037, i_4038, i_4039, i_4040, i_4041, i_4042, i_4067, i_4080, i_4088, i_4091, i_4094, i_4097, i_4100, i_4103, i_4106, i_4109, i_4144, i_4147, i_4150, i_4153, i_4156, i_4159, i_4183, i_4184, i_4185, i_4186, i_4188, i_4191, i_4196, i_4197, i_4198, i_4199, i_4200, i_4203, i_4206, i_4209, i_4212, i_4215, i_4219, i_4223, i_4224, i_4225, i_4228, i_4231, i_4234, i_4237, i_4240, i_4243, i_4246, i_4249, i_4252, i_4255, i_4258, i_4263, i_4264, i_4267, i_4268, i_4269, i_4270, i_4271, i_4273, i_4274, i_4276, i_4277, i_4280, i_4284, i_4290, i_4297, i_4298, i_4301, i_4305, i_4310, i_4316, i_4320, i_4325, i_4331, i_4332, i_4336, i_4342, i_4349, i_4357, i_4364, i_4375, i_4379, i_4385, i_4392, i_4396, i_4400, i_4405, i_4412, i_4418, i_4425, i_4436, i_4440, i_4445, i_4451, i_4456, i_4462, i_4469, i_4477, i_4512, i_4515, i_4516, i_4521, i_4523, i_4524, i_4532, i_4547, i_4548, i_4551, i_4554, i_4557, i_4560, i_4563, i_4566, i_4569, i_4572, i_4575, i_4578, i_4581, i_4584, i_4587, i_4590, i_4593, i_4596, i_4599, i_4602, i_4605, i_4608, i_4611, i_4614, i_4617, i_4621, i_4624, i_4627, i_4630, i_4633, i_4637, i_4640, i_4643, i_4646, i_4649, i_4652, i_4655, i_4658, i_4662, i_4665, i_4668, i_4671, i_4674, i_4677, i_4680, i_4683, i_4686, i_4689, i_4692, i_4695, i_4698, i_4701, i_4702, i_4720, i_4721, i_4724, i_4725, i_4726, i_4727, i_4728, i_4729, i_4730, i_4731, i_4732, i_4733, i_4734, i_4735, i_4736, i_4741, i_4855, i_4856, i_4908, i_4909, i_4939, i_4942, i_4947, i_4953, i_4954, i_4955, i_4956, i_4957, i_4958, i_4959, i_4960, i_4961, i_4965, i_4966, i_4967, i_4968, i_4972, i_4973, i_4974, i_4975, i_4976, i_4977, i_4978, i_4979, i_4980, i_4981, i_4982, i_4983, i_4984, i_4985, i_4986, i_4987, i_5049, i_5052, i_5053, i_5054, i_5055, i_5056, i_5057, i_5058, i_5059, i_5060, i_5061, i_5062, i_5063, i_5065, i_5066, i_5067, i_5068, i_5069, i_5070, i_5071, i_5072, i_5073, i_5074, i_5075, i_5076, i_5077, i_5078, i_5079, i_5080, i_5081, i_5082, i_5083, i_5084, i_5085, i_5086, i_5087, i_5088, i_5089, i_5090, i_5091, i_5092, i_5093, i_5094, i_5095, i_5096, i_5097, i_5098, i_5099, i_5100, i_5101, i_5102, i_5103, i_5104, i_5105, i_5106, i_5107, i_5108, i_5109, i_5110, i_5111, i_5112, i_5113, i_5114, i_5115, i_5116, i_5117, i_5118, i_5119, i_5120, i_5121, i_5122, i_5123, i_5124, i_5125, i_5126, i_5127, i_5128, i_5129, i_5130, i_5131, i_5132, i_5133, i_5135, i_5136, i_5137, i_5138, i_5139, i_5140, i_5141, i_5142, i_5143, i_5144, i_5145, i_5146, i_5147, i_5148, i_5150, i_5153, i_5154, i_5155, i_5156, i_5157, i_5160, i_5161, i_5162, i_5163, i_5164, i_5165, i_5166, i_5169, i_5172, i_5173, i_5176, i_5177, i_5180, i_5183, i_5186, i_5189, i_5192, i_5195, i_5198, i_5199, i_5202, i_5205, i_5208, i_5211, i_5214, i_5217, i_5220, i_5223, i_5224, i_5225, i_5226, i_5227, i_5228, i_5229, i_5230, i_5232, i_5233, i_5234, i_5235, i_5236, i_5239, i_5241, i_5242, i_5243, i_5244, i_5245, i_5246, i_5247, i_5248, i_5249, i_5250, i_5252, i_5253, i_5254, i_5255, i_5256, i_5257, i_5258, i_5259, i_5260, i_5261, i_5262, i_5263, i_5264, i_5274, i_5275, i_5282, i_5283, i_5284, i_5298, i_5299, i_5300, i_5303, i_5304, i_5305, i_5306, i_5307, i_5308, i_5309, i_5310, i_5311, i_5312, i_5315, i_5319, i_5324, i_5328, i_5331, i_5332, i_5346, i_5363, i_5364, i_5365, i_5366, i_5367, i_5368, i_5369, i_5370, i_5371, i_5374, i_5377, i_5382, i_5385, i_5389, i_5396, i_5407, i_5418, i_5424, i_5431, i_5441, i_5452, i_5462, i_5469, i_5470, i_5477, i_5488, i_5498, i_5506, i_5520, i_5536, i_5549, i_5555, i_5562, i_5573, i_5579, i_5595, i_5606, i_5616, i_5617, i_5618, i_5619, i_5620, i_5621, i_5622, i_5624, i_5634, i_5655, i_5671, i_5684, i_5690, i_5691, i_5692, i_5696, i_5700, i_5703, i_5707, i_5711, i_5726, i_5727, i_5728, i_5730, i_5731, i_5732, i_5733, i_5734, i_5735, i_5736, i_5739, i_5742, i_5745, i_5755, i_5756, i_5954, i_5955, i_5956, i_6005, i_6006, i_6023, i_6024, i_6025, i_6028, i_6031, i_6034, i_6037, i_6040, i_6044, i_6045, i_6048, i_6051, i_6054, i_6065, i_6066, i_6067, i_6068, i_6069, i_6071, i_6072, i_6073, i_6074, i_6075, i_6076, i_6077, i_6078, i_6079, i_6080, i_6083, i_6084, i_6085, i_6086, i_6087, i_6088, i_6089, i_6090, i_6091, i_6094, i_6095, i_6096, i_6097, i_6098, i_6099, i_6100, i_6101, i_6102, i_6103, i_6104, i_6105, i_6106, i_6107, i_6108, i_6111, i_6112, i_6113, i_6114, i_6115, i_6116, i_6117, i_6120, i_6121, i_6122, i_6123, i_6124, i_6125, i_6126, i_6127, i_6128, i_6129, i_6130, i_6131, i_6132, i_6133, i_6134, i_6135, i_6136, i_6137, i_6138, i_6139, i_6140, i_6143, i_6144, i_6145, i_6146, i_6147, i_6148, i_6149, i_6152, i_6153, i_6154, i_6155, i_6156, i_6157, i_6158, i_6159, i_6160, i_6161, i_6162, i_6163, i_6164, i_6168, i_6171, i_6172, i_6173, i_6174, i_6175, i_6178, i_6179, i_6180, i_6181, i_6182, i_6183, i_6184, i_6185, i_6186, i_6187, i_6188, i_6189, i_6190, i_6191, i_6192, i_6193, i_6194, i_6197, i_6200, i_6203, i_6206, i_6209, i_6212, i_6215, i_6218, i_6221, i_6234, i_6235, i_6238, i_6241, i_6244, i_6247, i_6250, i_6253, i_6256, i_6259, i_6262, i_6265, i_6268, i_6271, i_6274, i_6277, i_6280, i_6283, i_6286, i_6289, i_6292, i_6295, i_6298, i_6301, i_6304, i_6307, i_6310, i_6313, i_6316, i_6319, i_6322, i_6325, i_6328, i_6331, i_6335, i_6338, i_6341, i_6344, i_6347, i_6350, i_6353, i_6356, i_6359, i_6364, i_6367, i_6370, i_6373, i_6374, i_6375, i_6376, i_6377, i_6378, i_6382, i_6386, i_6388, i_6392, i_6397, i_6411, i_6415, i_6419, i_6427, i_6434, i_6437, i_6441, i_6445, i_6448, i_6449, i_6466, i_6469, i_6470, i_6471, i_6472, i_6473, i_6474, i_6475, i_6476, i_6477, i_6478, i_6482, i_6486, i_6490, i_6494, i_6500, i_6504, i_6508, i_6512, i_6516, i_6526, i_6536, i_6539, i_6553, i_6556, i_6566, i_6569, i_6572, i_6575, i_6580, i_6584, i_6587, i_6592, i_6599, i_6606, i_6609, i_6619, i_6622, i_6630, i_6631, i_6632, i_6633, i_6634, i_6637, i_6640, i_6650, i_6651, i_6653, i_6655, i_6657, i_6659, i_6660, i_6661, i_6662, i_6663, i_6664, i_6666, i_6668, i_6670, i_6672, i_6675, i_6680, i_6681, i_6682, i_6683, i_6689, i_6690, i_6691, i_6692, i_6693, i_6695, i_6698, i_6699, i_6700, i_6703, i_6708, i_6709, i_6710, i_6711, i_6712, i_6713, i_6714, i_6715, i_6718, i_6719, i_6720, i_6721, i_6722, i_6724, i_6739, i_6740, i_6741, i_6744, i_6745, i_6746, i_6751, i_6752, i_6753, i_6754, i_6755, i_6760, i_6761, i_6762, i_6772, i_6773, i_6776, i_6777, i_6782, i_6783, i_6784, i_6785, i_6790, i_6791, i_6792, i_6795, i_6801, i_6802, i_6803, i_6804, i_6805, i_6806, i_6807, i_6808, i_6809, i_6810, i_6811, i_6812, i_6813, i_6814, i_6815, i_6816, i_6817, i_6823, i_6824, i_6825, i_6826, i_6827, i_6828, i_6829, i_6830, i_6831, i_6834, i_6835, i_6836, i_6837, i_6838, i_6839, i_6840, i_6841, i_6842, i_6843, i_6844, i_6850, i_6851, i_6852, i_6853, i_6854, i_6855, i_6856, i_6857, i_6860, i_6861, i_6862, i_6863, i_6866, i_6872, i_6873, i_6874, i_6875, i_6876, i_6879, i_6880, i_6881, i_6884, i_6885, i_6888, i_6889, i_6890, i_6891, i_6894, i_6895, i_6896, i_6897, i_6900, i_6901, i_6904, i_6905, i_6908, i_6909, i_6912, i_6913, i_6914, i_6915, i_6916, i_6919, i_6922, i_6923, i_6930, i_6932, i_6935, i_6936, i_6937, i_6938, i_6939, i_6940, i_6946, i_6947, i_6948, i_6949, i_6953, i_6954, i_6955, i_6956, i_6957, i_6958, i_6964, i_6965, i_6966, i_6967, i_6973, i_6974, i_6975, i_6976, i_6977, i_6978, i_6979, i_6987, i_6990, i_6999, i_7002, i_7003, i_7006, i_7011, i_7012, i_7013, i_7016, i_7018, i_7019, i_7020, i_7021, i_7022, i_7023, i_7028, i_7031, i_7034, i_7037, i_7040, i_7041, i_7044, i_7045, i_7046, i_7047, i_7048, i_7049, i_7054, i_7057, i_7060, i_7064, i_7065, i_7072, i_7073, i_7074, i_7075, i_7076, i_7079, i_7080, i_7083, i_7084, i_7085, i_7086, i_7087, i_7088, i_7089, i_7090, i_7093, i_7094, i_7097, i_7101, i_7105, i_7110, i_7114, i_7115, i_7116, i_7125, i_7126, i_7127, i_7130, i_7131, i_7139, i_7140, i_7141, i_7146, i_7147, i_7149, i_7150, i_7151, i_7152, i_7153, i_7158, i_7159, i_7160, i_7166, i_7167, i_7168, i_7169, i_7170, i_7171, i_7172, i_7173, i_7174, i_7175, i_7176, i_7177, i_7178, i_7179, i_7180, i_7181, i_7182, i_7183, i_7184, i_7185, i_7186, i_7187, i_7188, i_7189, i_7190, i_7196, i_7197, i_7198, i_7204, i_7205, i_7206, i_7207, i_7208, i_7209, i_7212, i_7215, i_7216, i_7217, i_7218, i_7219, i_7222, i_7225, i_7228, i_7229, i_7236, i_7239, i_7242, i_7245, i_7250, i_7257, i_7260, i_7263, i_7268, i_7269, i_7270, i_7276, i_7282, i_7288, i_7294, i_7300, i_7301, i_7304, i_7310, i_7320, i_7321, i_7328, i_7338, i_7339, i_7340, i_7341, i_7342, i_7349, i_7357, i_7364, i_7394, i_7397, i_7402, i_7405, i_7406, i_7407, i_7408, i_7409, i_7412, i_7415, i_7416, i_7417, i_7418, i_7419, i_7420, i_7421, i_7424, i_7425, i_7426, i_7427, i_7428, i_7429, i_7430, i_7431, i_7433, i_7434, i_7435, i_7436, i_7437, i_7438, i_7439, i_7440, i_7441, i_7442, i_7443, i_7444, i_7445, i_7446, i_7447, i_7448, i_7450, i_7451, i_7452, i_7453, i_7454, i_7455, i_7456, i_7457, i_7458, i_7459, i_7460, i_7461, i_7462, i_7463, i_7464, i_7468, i_7479, i_7481, i_7482, i_7483, i_7484, i_7485, i_7486, i_7487, i_7488, i_7489, i_7492, i_7493, i_7498, i_7499, i_7500, i_7505, i_7507, i_7508, i_7509, i_7510, i_7512, i_7513, i_7514, i_7525, i_7526, i_7527, i_7528, i_7529, i_7530, i_7531, i_7537, i_7543, i_7549, i_7555, i_7561, i_7567, i_7573, i_7579, i_7582, i_7585, i_7586, i_7587, i_7588, i_7589, i_7592, i_7595, i_7598, i_7599, i_7624, i_7625, i_7631, i_7636, i_7657, i_7658, i_7665, i_7666, i_7667, i_7668, i_7669, i_7670, i_7671, i_7672, i_7673, i_7674, i_7675, i_7676, i_7677, i_7678, i_7679, i_7680, i_7681, i_7682, i_7683, i_7684, i_7685, i_7686, i_7687, i_7688, i_7689, i_7690, i_7691, i_7692, i_7693, i_7694, i_7695, i_7696, i_7697, i_7708, i_7709, i_7710, i_7711, i_7712, i_7715, i_7718, i_7719, i_7720, i_7721, i_7722, i_7723, i_7724, i_7727, i_7728, i_7729, i_7730, i_7731, i_7732, i_7733, i_7734, i_7743, i_7744, i_7749, i_7750, i_7751, i_7762, i_7765, i_7768, i_7769, i_7770, i_7771, i_7772, i_7775, i_7778, i_7781, i_7782, i_7787, i_7788, i_7795, i_7796, i_7797, i_7798, i_7799, i_7800, i_7803, i_7806, i_7807, i_7808, i_7809, i_7810, i_7811, i_7812, i_7815, i_7816, i_7821, i_7822, i_7823, i_7826, i_7829, i_7832, i_7833, i_7834, i_7835, i_7836, i_7839, i_7842, i_7845, i_7846, i_7851, i_7852, i_7859, i_7860, i_7861, i_7862, i_7863, i_7864, i_7867, i_7870, i_7871, i_7872, i_7873, i_7874, i_7875, i_7876, i_7879, i_7880, i_7885, i_7886, i_7887, i_7890, i_7893, i_7896, i_7897, i_7898, i_7899, i_7900, i_7903, i_7906, i_7909, i_7910, i_7917, i_7918, i_7923, i_7924, i_7925, i_7926, i_7927, i_7928, i_7929, i_7930, i_7931, i_7932, i_7935, i_7938, i_7939, i_7940, i_7943, i_7944, i_7945, i_7946, i_7951, i_7954, i_7957, i_7960, i_7963, i_7966, i_7967, i_7968, i_7969, i_7970, i_7973, i_7974, i_7984, i_7985, i_7987, i_7988, i_7989, i_7990, i_7991, i_7992, i_7993, i_7994, i_7995, i_7996, i_7997, i_7998, i_8001, i_8004, i_8009, i_8013, i_8017, i_8020, i_8021, i_8022, i_8023, i_8025, i_8026, i_8027, i_8031, i_8032, i_8033, i_8034, i_8035, i_8036, i_8037, i_8038, i_8039, i_8040, i_8041, i_8042, i_8043, i_8044, i_8045, i_8048, i_8055, i_8056, i_8057, i_8058, i_8059, i_8060, i_8061, i_8064, i_8071, i_8072, i_8073, i_8074, i_8077, i_8078, i_8079, i_8082, i_8089, i_8090, i_8091, i_8092, i_8093, i_8096, i_8099, i_8102, i_8113, i_8114, i_8115, i_8116, i_8117, i_8118, i_8119, i_8120, i_8121, i_8122, i_8125, i_8126, i_7701_in, flip_signal;

  and ginst2 (i_1042, i_135, i_631);
  not ginst3 (i_1043, i_591);
  not ginst4 (i_1066, i_592);
  not ginst5 (i_1067, i_595);
  not ginst6 (i_1080, i_596);
  not ginst7 (i_1092, i_597);
  not ginst8 (i_1104, i_598);
  not ginst9 (i_1137, i_545);
  not ginst10 (i_1138, i_348);
  not ginst11 (i_1139, i_366);
  and ginst12 (i_1140, i_552, i_562);
  not ginst13 (i_1141, i_549);
  not ginst14 (i_1142, i_545);
  not ginst15 (i_1143, i_545);
  not ginst16 (i_1144, i_338);
  not ginst17 (i_1145, i_358);
  nand ginst18 (i_1146, i_1, i_373);
  and ginst19 (i_1147, i_141, i_145);
  not ginst20 (i_1148, i_592);
  not ginst21 (i_1149, i_1042);
  and ginst22 (i_1150, i_27, i_1043);
  and ginst23 (i_1151, i_386, i_556);
  not ginst24 (i_1152, i_245);
  not ginst25 (i_1153, i_552);
  not ginst26 (i_1154, i_562);
  not ginst27 (i_1155, i_559);
  and ginst28 (i_1156, i_386, i_552, i_556, i_559);
  not ginst29 (i_1157, i_566);
  not ginst30 (i_1161, i_571);
  not ginst31 (i_1173, i_574);
  not ginst32 (i_1185, i_571);
  not ginst33 (i_1197, i_574);
  not ginst34 (i_1209, i_137);
  not ginst35 (i_1213, i_137);
  not ginst36 (i_1216, i_141);
  not ginst37 (i_1219, i_583);
  not ginst38 (i_1223, i_577);
  not ginst39 (i_1235, i_580);
  not ginst40 (i_1247, i_577);
  not ginst41 (i_1259, i_580);
  not ginst42 (i_1271, i_254);
  not ginst43 (i_1280, i_251);
  not ginst44 (i_1292, i_251);
  not ginst45 (i_1303, i_248);
  not ginst46 (i_1315, i_248);
  not ginst47 (i_1327, i_610);
  not ginst48 (i_1339, i_607);
  not ginst49 (i_1351, i_613);
  not ginst50 (i_1363, i_616);
  not ginst51 (i_1375, i_210);
  not ginst52 (i_1378, i_210);
  not ginst53 (i_1381, i_218);
  not ginst54 (i_1384, i_218);
  not ginst55 (i_1387, i_226);
  not ginst56 (i_1390, i_226);
  not ginst57 (i_1393, i_234);
  not ginst58 (i_1396, i_234);
  not ginst59 (i_1415, i_257);
  not ginst60 (i_1418, i_257);
  not ginst61 (i_1421, i_265);
  not ginst62 (i_1424, i_265);
  not ginst63 (i_1427, i_273);
  not ginst64 (i_1430, i_273);
  not ginst65 (i_1433, i_281);
  not ginst66 (i_1436, i_281);
  not ginst67 (i_1455, i_335);
  not ginst68 (i_1462, i_335);
  not ginst69 (i_1469, i_206);
  and ginst70 (i_1475, i_27, i_31);
  not ginst71 (i_1479, i_1);
  not ginst72 (i_1482, i_588);
  not ginst73 (i_1492, i_293);
  not ginst74 (i_1495, i_302);
  not ginst75 (i_1498, i_308);
  not ginst76 (i_1501, i_308);
  not ginst77 (i_1504, i_316);
  not ginst78 (i_1507, i_316);
  not ginst79 (i_1510, i_324);
  not ginst80 (i_1513, i_324);
  not ginst81 (i_1516, i_341);
  not ginst82 (i_1519, i_341);
  not ginst83 (i_1522, i_351);
  not ginst84 (i_1525, i_351);
  not ginst85 (i_1542, i_257);
  not ginst86 (i_1545, i_257);
  not ginst87 (i_1548, i_265);
  not ginst88 (i_1551, i_265);
  not ginst89 (i_1554, i_273);
  not ginst90 (i_1557, i_273);
  not ginst91 (i_1560, i_281);
  not ginst92 (i_1563, i_281);
  not ginst93 (i_1566, i_332);
  not ginst94 (i_1573, i_332);
  not ginst95 (i_1580, i_549);
  and ginst96 (i_1583, i_27, i_31);
  not ginst97 (i_1588, i_588);
  not ginst98 (i_1594, i_324);
  not ginst99 (i_1597, i_324);
  not ginst100 (i_1600, i_341);
  not ginst101 (i_1603, i_341);
  not ginst102 (i_1606, i_351);
  not ginst103 (i_1609, i_351);
  not ginst104 (i_1612, i_293);
  not ginst105 (i_1615, i_302);
  not ginst106 (i_1618, i_308);
  not ginst107 (i_1621, i_308);
  not ginst108 (i_1624, i_316);
  not ginst109 (i_1627, i_316);
  not ginst110 (i_1630, i_361);
  not ginst111 (i_1633, i_361);
  not ginst112 (i_1636, i_210);
  not ginst113 (i_1639, i_210);
  not ginst114 (i_1642, i_218);
  not ginst115 (i_1645, i_218);
  not ginst116 (i_1648, i_226);
  not ginst117 (i_1651, i_226);
  not ginst118 (i_1654, i_234);
  not ginst119 (i_1657, i_234);
  not ginst120 (i_1660, i_324);
  not ginst121 (i_1663, i_242);
  not ginst122 (i_1675, i_242);
  not ginst123 (i_1685, i_254);
  not ginst124 (i_1697, i_610);
  not ginst125 (i_1709, i_607);
  not ginst126 (i_1721, i_625);
  not ginst127 (i_1727, i_619);
  not ginst128 (i_1731, i_613);
  not ginst129 (i_1743, i_616);
  not ginst130 (i_1755, i_599);
  not ginst131 (i_1758, i_603);
  not ginst132 (i_1761, i_619);
  not ginst133 (i_1769, i_625);
  not ginst134 (i_1777, i_619);
  not ginst135 (i_1785, i_625);
  not ginst136 (i_1793, i_619);
  not ginst137 (i_1800, i_625);
  not ginst138 (i_1807, i_619);
  not ginst139 (i_1814, i_625);
  not ginst140 (i_1821, i_299);
  not ginst141 (i_1824, i_446);
  not ginst142 (i_1827, i_457);
  not ginst143 (i_1830, i_468);
  not ginst144 (i_1833, i_422);
  not ginst145 (i_1836, i_435);
  not ginst146 (i_1839, i_389);
  not ginst147 (i_1842, i_400);
  not ginst148 (i_1845, i_411);
  not ginst149 (i_1848, i_374);
  not ginst150 (i_1851, i_4);
  not ginst151 (i_1854, i_446);
  not ginst152 (i_1857, i_457);
  not ginst153 (i_1860, i_468);
  not ginst154 (i_1863, i_435);
  not ginst155 (i_1866, i_389);
  not ginst156 (i_1869, i_400);
  not ginst157 (i_1872, i_411);
  not ginst158 (i_1875, i_422);
  not ginst159 (i_1878, i_374);
  not ginst160 (i_1881, i_479);
  not ginst161 (i_1884, i_490);
  not ginst162 (i_1887, i_503);
  not ginst163 (i_1890, i_514);
  not ginst164 (i_1893, i_523);
  not ginst165 (i_1896, i_534);
  not ginst166 (i_1899, i_54);
  not ginst167 (i_1902, i_479);
  not ginst168 (i_1905, i_503);
  not ginst169 (i_1908, i_514);
  not ginst170 (i_1911, i_523);
  not ginst171 (i_1914, i_534);
  not ginst172 (i_1917, i_490);
  not ginst173 (i_1920, i_361);
  not ginst174 (i_1923, i_369);
  not ginst175 (i_1926, i_341);
  not ginst176 (i_1929, i_351);
  not ginst177 (i_1932, i_308);
  not ginst178 (i_1935, i_316);
  not ginst179 (i_1938, i_293);
  not ginst180 (i_1941, i_302);
  not ginst181 (i_1944, i_281);
  not ginst182 (i_1947, i_289);
  not ginst183 (i_1950, i_265);
  not ginst184 (i_1953, i_273);
  not ginst185 (i_1956, i_234);
  not ginst186 (i_1959, i_257);
  not ginst187 (i_1962, i_218);
  not ginst188 (i_1965, i_226);
  not ginst189 (i_1968, i_210);
  not ginst190 (i_1972, i_1146);
  and ginst191 (i_2054, i_136, i_1148);
  not ginst192 (i_2060, i_1150);
  not ginst193 (i_2061, i_1151);
  not ginst194 (i_2139, i_1209);
  not ginst195 (i_2142, i_1216);
  not ginst196 (i_2309, i_1479);
  and ginst197 (i_2349, i_514, i_1104);
  or ginst198 (i_2350, i_514, i_1067);
  not ginst199 (i_2387, i_1580);
  not ginst200 (i_2527, i_1821);
  not ginst201 (i_2584, i_1580);
  and ginst202 (i_2585, i_170, i_1161, i_1173);
  and ginst203 (i_2586, i_173, i_1161, i_1173);
  and ginst204 (i_2587, i_167, i_1161, i_1173);
  and ginst205 (i_2588, i_164, i_1161, i_1173);
  and ginst206 (i_2589, i_161, i_1161, i_1173);
  nand ginst207 (i_2590, i_140, i_1475);
  and ginst208 (i_2591, i_185, i_1185, i_1197);
  and ginst209 (i_2592, i_158, i_1185, i_1197);
  and ginst210 (i_2593, i_152, i_1185, i_1197);
  and ginst211 (i_2594, i_146, i_1185, i_1197);
  and ginst212 (i_2595, i_170, i_1223, i_1235);
  and ginst213 (i_2596, i_173, i_1223, i_1235);
  and ginst214 (i_2597, i_167, i_1223, i_1235);
  and ginst215 (i_2598, i_164, i_1223, i_1235);
  and ginst216 (i_2599, i_161, i_1223, i_1235);
  and ginst217 (i_2600, i_185, i_1247, i_1259);
  and ginst218 (i_2601, i_158, i_1247, i_1259);
  and ginst219 (i_2602, i_152, i_1247, i_1259);
  and ginst220 (i_2603, i_146, i_1247, i_1259);
  and ginst221 (i_2604, i_106, i_1731, i_1743);
  and ginst222 (i_2605, i_61, i_1327, i_1339);
  and ginst223 (i_2606, i_106, i_1697, i_1709);
  and ginst224 (i_2607, i_49, i_1697, i_1709);
  and ginst225 (i_2608, i_103, i_1697, i_1709);
  and ginst226 (i_2609, i_40, i_1697, i_1709);
  and ginst227 (i_2610, i_37, i_1697, i_1709);
  and ginst228 (i_2611, i_20, i_1327, i_1339);
  and ginst229 (i_2612, i_17, i_1327, i_1339);
  and ginst230 (i_2613, i_70, i_1327, i_1339);
  and ginst231 (i_2614, i_64, i_1327, i_1339);
  and ginst232 (i_2615, i_49, i_1731, i_1743);
  and ginst233 (i_2616, i_103, i_1731, i_1743);
  and ginst234 (i_2617, i_40, i_1731, i_1743);
  and ginst235 (i_2618, i_37, i_1731, i_1743);
  and ginst236 (i_2619, i_20, i_1351, i_1363);
  and ginst237 (i_2620, i_17, i_1351, i_1363);
  and ginst238 (i_2621, i_70, i_1351, i_1363);
  and ginst239 (i_2622, i_64, i_1351, i_1363);
  not ginst240 (i_2623, i_1475);
  and ginst241 (i_2624, i_123, i_599, i_1758);
  and ginst242 (i_2625, i_1777, i_1785);
  and ginst243 (i_2626, i_61, i_1351, i_1363);
  and ginst244 (i_2627, i_1761, i_1769);
  not ginst245 (i_2628, i_1824);
  not ginst246 (i_2629, i_1827);
  not ginst247 (i_2630, i_1830);
  not ginst248 (i_2631, i_1833);
  not ginst249 (i_2632, i_1836);
  not ginst250 (i_2633, i_1839);
  not ginst251 (i_2634, i_1842);
  not ginst252 (i_2635, i_1845);
  not ginst253 (i_2636, i_1848);
  not ginst254 (i_2637, i_1851);
  not ginst255 (i_2638, i_1854);
  not ginst256 (i_2639, i_1857);
  not ginst257 (i_2640, i_1860);
  not ginst258 (i_2641, i_1863);
  not ginst259 (i_2642, i_1866);
  not ginst260 (i_2643, i_1869);
  not ginst261 (i_2644, i_1872);
  not ginst262 (i_2645, i_1875);
  not ginst263 (i_2646, i_1878);
  not ginst264 (i_2647, i_1209);
  not ginst265 (i_2653, i_1161);
  not ginst266 (i_2664, i_1173);
  not ginst267 (i_2675, i_1209);
  not ginst268 (i_2681, i_1185);
  not ginst269 (i_2692, i_1197);
  and ginst270 (i_2703, i_179, i_1185, i_1197);
  not ginst271 (i_2704, i_1479);
  not ginst272 (i_2709, i_1881);
  not ginst273 (i_2710, i_1884);
  not ginst274 (i_2711, i_1887);
  not ginst275 (i_2712, i_1890);
  not ginst276 (i_2713, i_1893);
  not ginst277 (i_2714, i_1896);
  not ginst278 (i_2715, i_1899);
  not ginst279 (i_2716, i_1902);
  not ginst280 (i_2717, i_1905);
  not ginst281 (i_2718, i_1908);
  not ginst282 (i_2719, i_1911);
  not ginst283 (i_2720, i_1914);
  not ginst284 (i_2721, i_1917);
  not ginst285 (i_2722, i_1213);
  not ginst286 (i_2728, i_1223);
  not ginst287 (i_2739, i_1235);
  not ginst288 (i_2750, i_1213);
  not ginst289 (i_2756, i_1247);
  not ginst290 (i_2767, i_1259);
  and ginst291 (i_2778, i_179, i_1247, i_1259);
  not ginst292 (i_2779, i_1327);
  not ginst293 (i_2790, i_1339);
  not ginst294 (i_2801, i_1351);
  not ginst295 (i_2812, i_1363);
  not ginst296 (i_2823, i_1375);
  not ginst297 (i_2824, i_1378);
  not ginst298 (i_2825, i_1381);
  not ginst299 (i_2826, i_1384);
  not ginst300 (i_2827, i_1387);
  not ginst301 (i_2828, i_1390);
  not ginst302 (i_2829, i_1393);
  not ginst303 (i_2830, i_1396);
  and ginst304 (i_2831, i_457, i_1104, i_1378);
  and ginst305 (i_2832, i_468, i_1104, i_1384);
  and ginst306 (i_2833, i_422, i_1104, i_1390);
  and ginst307 (i_2834, i_435, i_1104, i_1396);
  and ginst308 (i_2835, i_1067, i_1375);
  and ginst309 (i_2836, i_1067, i_1381);
  and ginst310 (i_2837, i_1067, i_1387);
  and ginst311 (i_2838, i_1067, i_1393);
  not ginst312 (i_2839, i_1415);
  not ginst313 (i_2840, i_1418);
  not ginst314 (i_2841, i_1421);
  not ginst315 (i_2842, i_1424);
  not ginst316 (i_2843, i_1427);
  not ginst317 (i_2844, i_1430);
  not ginst318 (i_2845, i_1433);
  not ginst319 (i_2846, i_1436);
  and ginst320 (i_2847, i_389, i_1104, i_1418);
  and ginst321 (i_2848, i_400, i_1104, i_1424);
  and ginst322 (i_2849, i_411, i_1104, i_1430);
  and ginst323 (i_2850, i_374, i_1104, i_1436);
  and ginst324 (i_2851, i_1067, i_1415);
  and ginst325 (i_2852, i_1067, i_1421);
  and ginst326 (i_2853, i_1067, i_1427);
  and ginst327 (i_2854, i_1067, i_1433);
  not ginst328 (i_2855, i_1455);
  not ginst329 (i_2861, i_1462);
  and ginst330 (i_2867, i_292, i_1455);
  and ginst331 (i_2868, i_288, i_1455);
  and ginst332 (i_2869, i_280, i_1455);
  and ginst333 (i_2870, i_272, i_1455);
  and ginst334 (i_2871, i_264, i_1455);
  and ginst335 (i_2872, i_241, i_1462);
  and ginst336 (i_2873, i_233, i_1462);
  and ginst337 (i_2874, i_225, i_1462);
  and ginst338 (i_2875, i_217, i_1462);
  and ginst339 (i_2876, i_209, i_1462);
  not ginst340 (i_2877, i_1216);
  not ginst341 (i_2882, i_1482);
  not ginst342 (i_2891, i_1475);
  not ginst343 (i_2901, i_1492);
  not ginst344 (i_2902, i_1495);
  not ginst345 (i_2903, i_1498);
  not ginst346 (i_2904, i_1501);
  not ginst347 (i_2905, i_1504);
  not ginst348 (i_2906, i_1507);
  and ginst349 (i_2907, i_1303, i_1495);
  and ginst350 (i_2908, i_479, i_1303, i_1501);
  and ginst351 (i_2909, i_490, i_1303, i_1507);
  and ginst352 (i_2910, i_1492, i_1663);
  and ginst353 (i_2911, i_1498, i_1663);
  and ginst354 (i_2912, i_1504, i_1663);
  not ginst355 (i_2913, i_1510);
  not ginst356 (i_2914, i_1513);
  not ginst357 (i_2915, i_1516);
  not ginst358 (i_2916, i_1519);
  not ginst359 (i_2917, i_1522);
  not ginst360 (i_2918, i_1525);
  and ginst361 (i_2919, i_503, i_1104, i_1513);
  not ginst362 (i_2920, i_2349);
  and ginst363 (i_2921, i_523, i_1104, i_1519);
  and ginst364 (i_2922, i_534, i_1104, i_1525);
  and ginst365 (i_2923, i_1067, i_1510);
  and ginst366 (i_2924, i_1067, i_1516);
  and ginst367 (i_2925, i_1067, i_1522);
  not ginst368 (i_2926, i_1542);
  not ginst369 (i_2927, i_1545);
  not ginst370 (i_2928, i_1548);
  not ginst371 (i_2929, i_1551);
  not ginst372 (i_2930, i_1554);
  not ginst373 (i_2931, i_1557);
  not ginst374 (i_2932, i_1560);
  not ginst375 (i_2933, i_1563);
  and ginst376 (i_2934, i_389, i_1303, i_1545);
  and ginst377 (i_2935, i_400, i_1303, i_1551);
  and ginst378 (i_2936, i_411, i_1303, i_1557);
  and ginst379 (i_2937, i_374, i_1303, i_1563);
  and ginst380 (i_2938, i_1542, i_1663);
  and ginst381 (i_2939, i_1548, i_1663);
  and ginst382 (i_2940, i_1554, i_1663);
  and ginst383 (i_2941, i_1560, i_1663);
  not ginst384 (i_2942, i_1566);
  not ginst385 (i_2948, i_1573);
  and ginst386 (i_2954, i_372, i_1566);
  and ginst387 (i_2955, i_366, i_1566);
  and ginst388 (i_2956, i_358, i_1566);
  and ginst389 (i_2957, i_348, i_1566);
  and ginst390 (i_2958, i_338, i_1566);
  and ginst391 (i_2959, i_331, i_1573);
  and ginst392 (i_2960, i_323, i_1573);
  and ginst393 (i_2961, i_315, i_1573);
  and ginst394 (i_2962, i_307, i_1573);
  and ginst395 (i_2963, i_299, i_1573);
  not ginst396 (i_2964, i_1588);
  and ginst397 (i_2969, i_83, i_1588);
  and ginst398 (i_2970, i_86, i_1588);
  and ginst399 (i_2971, i_88, i_1588);
  and ginst400 (i_2972, i_88, i_1588);
  not ginst401 (i_2973, i_1594);
  not ginst402 (i_2974, i_1597);
  not ginst403 (i_2975, i_1600);
  not ginst404 (i_2976, i_1603);
  not ginst405 (i_2977, i_1606);
  not ginst406 (i_2978, i_1609);
  and ginst407 (i_2979, i_503, i_1315, i_1597);
  and ginst408 (i_2980, i_514, i_1315);
  and ginst409 (i_2981, i_523, i_1315, i_1603);
  and ginst410 (i_2982, i_534, i_1315, i_1609);
  and ginst411 (i_2983, i_1594, i_1675);
  or ginst412 (i_2984, i_514, i_1675);
  and ginst413 (i_2985, i_1600, i_1675);
  and ginst414 (i_2986, i_1606, i_1675);
  not ginst415 (i_2987, i_1612);
  not ginst416 (i_2988, i_1615);
  not ginst417 (i_2989, i_1618);
  not ginst418 (i_2990, i_1621);
  not ginst419 (i_2991, i_1624);
  not ginst420 (i_2992, i_1627);
  and ginst421 (i_2993, i_1315, i_1615);
  and ginst422 (i_2994, i_479, i_1315, i_1621);
  and ginst423 (i_2995, i_490, i_1315, i_1627);
  and ginst424 (i_2996, i_1612, i_1675);
  and ginst425 (i_2997, i_1618, i_1675);
  and ginst426 (i_2998, i_1624, i_1675);
  not ginst427 (i_2999, i_1630);
  not ginst428 (i_3000, i_1469);
  not ginst429 (i_3003, i_1469);
  not ginst430 (i_3006, i_1633);
  not ginst431 (i_3007, i_1469);
  not ginst432 (i_3010, i_1469);
  and ginst433 (i_3013, i_1315, i_1630);
  and ginst434 (i_3014, i_1315, i_1633);
  not ginst435 (i_3015, i_1636);
  not ginst436 (i_3016, i_1639);
  not ginst437 (i_3017, i_1642);
  not ginst438 (i_3018, i_1645);
  not ginst439 (i_3019, i_1648);
  not ginst440 (i_3020, i_1651);
  not ginst441 (i_3021, i_1654);
  not ginst442 (i_3022, i_1657);
  and ginst443 (i_3023, i_457, i_1303, i_1639);
  and ginst444 (i_3024, i_468, i_1303, i_1645);
  and ginst445 (i_3025, i_422, i_1303, i_1651);
  and ginst446 (i_3026, i_435, i_1303, i_1657);
  and ginst447 (i_3027, i_1636, i_1663);
  and ginst448 (i_3028, i_1642, i_1663);
  and ginst449 (i_3029, i_1648, i_1663);
  and ginst450 (i_3030, i_1654, i_1663);
  not ginst451 (i_3031, i_1920);
  not ginst452 (i_3032, i_1923);
  not ginst453 (i_3033, i_1926);
  not ginst454 (i_3034, i_1929);
  not ginst455 (i_3035, i_1660);
  not ginst456 (i_3038, i_1660);
  not ginst457 (i_3041, i_1697);
  not ginst458 (i_3052, i_1709);
  not ginst459 (i_3063, i_1721);
  not ginst460 (i_3068, i_1727);
  and ginst461 (i_3071, i_97, i_1721);
  and ginst462 (i_3072, i_94, i_1721);
  and ginst463 (i_3073, i_97, i_1721);
  and ginst464 (i_3074, i_94, i_1721);
  not ginst465 (i_3075, i_1731);
  not ginst466 (i_3086, i_1743);
  not ginst467 (i_3097, i_1761);
  not ginst468 (i_3108, i_1769);
  not ginst469 (i_3119, i_1777);
  not ginst470 (i_3130, i_1785);
  not ginst471 (i_3141, i_1944);
  not ginst472 (i_3142, i_1947);
  not ginst473 (i_3143, i_1950);
  not ginst474 (i_3144, i_1953);
  not ginst475 (i_3145, i_1956);
  not ginst476 (i_3146, i_1959);
  not ginst477 (i_3147, i_1793);
  not ginst478 (i_3158, i_1800);
  not ginst479 (i_3169, i_1807);
  not ginst480 (i_3180, i_1814);
  not ginst481 (i_3191, i_1821);
  not ginst482 (i_3194, i_1932);
  not ginst483 (i_3195, i_1935);
  not ginst484 (i_3196, i_1938);
  not ginst485 (i_3197, i_1941);
  not ginst486 (i_3198, i_1962);
  not ginst487 (i_3199, i_1965);
  not ginst488 (i_3200, i_1469);
  not ginst489 (i_3203, i_1968);
  not ginst490 (i_3357, i_2704);
  not ginst491 (i_3358, i_2704);
  not ginst492 (i_3359, i_2704);
  not ginst493 (i_3360, i_2704);
  and ginst494 (i_3401, i_457, i_1092, i_2824);
  and ginst495 (i_3402, i_468, i_1092, i_2826);
  and ginst496 (i_3403, i_422, i_1092, i_2828);
  and ginst497 (i_3404, i_435, i_1092, i_2830);
  and ginst498 (i_3405, i_1080, i_2823);
  and ginst499 (i_3406, i_1080, i_2825);
  and ginst500 (i_3407, i_1080, i_2827);
  and ginst501 (i_3408, i_1080, i_2829);
  and ginst502 (i_3409, i_389, i_1092, i_2840);
  and ginst503 (i_3410, i_400, i_1092, i_2842);
  and ginst504 (i_3411, i_411, i_1092, i_2844);
  and ginst505 (i_3412, i_374, i_1092, i_2846);
  and ginst506 (i_3413, i_1080, i_2839);
  and ginst507 (i_3414, i_1080, i_2841);
  and ginst508 (i_3415, i_1080, i_2843);
  and ginst509 (i_3416, i_1080, i_2845);
  and ginst510 (i_3444, i_1280, i_2902);
  and ginst511 (i_3445, i_479, i_1280, i_2904);
  and ginst512 (i_3446, i_490, i_1280, i_2906);
  and ginst513 (i_3447, i_1685, i_2901);
  and ginst514 (i_3448, i_1685, i_2903);
  and ginst515 (i_3449, i_1685, i_2905);
  and ginst516 (i_3450, i_503, i_1092, i_2914);
  and ginst517 (i_3451, i_523, i_1092, i_2916);
  and ginst518 (i_3452, i_534, i_1092, i_2918);
  and ginst519 (i_3453, i_1080, i_2913);
  and ginst520 (i_3454, i_1080, i_2915);
  and ginst521 (i_3455, i_1080, i_2917);
  and ginst522 (i_3456, i_2350, i_2920);
  and ginst523 (i_3459, i_389, i_1280, i_2927);
  and ginst524 (i_3460, i_400, i_1280, i_2929);
  and ginst525 (i_3461, i_411, i_1280, i_2931);
  and ginst526 (i_3462, i_374, i_1280, i_2933);
  and ginst527 (i_3463, i_1685, i_2926);
  and ginst528 (i_3464, i_1685, i_2928);
  and ginst529 (i_3465, i_1685, i_2930);
  and ginst530 (i_3466, i_1685, i_2932);
  and ginst531 (i_3481, i_503, i_1292, i_2974);
  not ginst532 (i_3482, i_2980);
  and ginst533 (i_3483, i_523, i_1292, i_2976);
  and ginst534 (i_3484, i_534, i_1292, i_2978);
  and ginst535 (i_3485, i_1271, i_2973);
  and ginst536 (i_3486, i_1271, i_2975);
  and ginst537 (i_3487, i_1271, i_2977);
  and ginst538 (i_3488, i_1292, i_2988);
  and ginst539 (i_3489, i_479, i_1292, i_2990);
  and ginst540 (i_3490, i_490, i_1292, i_2992);
  and ginst541 (i_3491, i_1271, i_2987);
  and ginst542 (i_3492, i_1271, i_2989);
  and ginst543 (i_3493, i_1271, i_2991);
  and ginst544 (i_3502, i_1292, i_2999);
  and ginst545 (i_3503, i_1292, i_3006);
  and ginst546 (i_3504, i_457, i_1280, i_3016);
  and ginst547 (i_3505, i_468, i_1280, i_3018);
  and ginst548 (i_3506, i_422, i_1280, i_3020);
  and ginst549 (i_3507, i_435, i_1280, i_3022);
  and ginst550 (i_3508, i_1685, i_3015);
  and ginst551 (i_3509, i_1685, i_3017);
  and ginst552 (i_3510, i_1685, i_3019);
  and ginst553 (i_3511, i_1685, i_3021);
  nand ginst554 (i_3512, i_1923, i_3031);
  nand ginst555 (i_3513, i_1920, i_3032);
  nand ginst556 (i_3514, i_1929, i_3033);
  nand ginst557 (i_3515, i_1926, i_3034);
  nand ginst558 (i_3558, i_1947, i_3141);
  nand ginst559 (i_3559, i_1944, i_3142);
  nand ginst560 (i_3560, i_1953, i_3143);
  nand ginst561 (i_3561, i_1950, i_3144);
  nand ginst562 (i_3562, i_1959, i_3145);
  nand ginst563 (i_3563, i_1956, i_3146);
  not ginst564 (i_3604, i_3191);
  nand ginst565 (i_3605, i_1935, i_3194);
  nand ginst566 (i_3606, i_1932, i_3195);
  nand ginst567 (i_3607, i_1941, i_3196);
  nand ginst568 (i_3608, i_1938, i_3197);
  nand ginst569 (i_3609, i_1965, i_3198);
  nand ginst570 (i_3610, i_1962, i_3199);
  not ginst571 (i_3613, i_3191);
  and ginst572 (i_3614, i_2882, i_2891);
  and ginst573 (i_3615, i_1482, i_2891);
  and ginst574 (i_3616, i_200, i_1173, i_2653);
  and ginst575 (i_3617, i_203, i_1173, i_2653);
  and ginst576 (i_3618, i_197, i_1173, i_2653);
  and ginst577 (i_3619, i_194, i_1173, i_2653);
  and ginst578 (i_3620, i_191, i_1173, i_2653);
  and ginst579 (i_3621, i_182, i_1197, i_2681);
  and ginst580 (i_3622, i_188, i_1197, i_2681);
  and ginst581 (i_3623, i_155, i_1197, i_2681);
  and ginst582 (i_3624, i_149, i_1197, i_2681);
  and ginst583 (i_3625, i_2882, i_2891);
  and ginst584 (i_3626, i_1482, i_2891);
  and ginst585 (i_3627, i_200, i_1235, i_2728);
  and ginst586 (i_3628, i_203, i_1235, i_2728);
  and ginst587 (i_3629, i_197, i_1235, i_2728);
  and ginst588 (i_3630, i_194, i_1235, i_2728);
  and ginst589 (i_3631, i_191, i_1235, i_2728);
  and ginst590 (i_3632, i_182, i_1259, i_2756);
  and ginst591 (i_3633, i_188, i_1259, i_2756);
  and ginst592 (i_3634, i_155, i_1259, i_2756);
  and ginst593 (i_3635, i_149, i_1259, i_2756);
  and ginst594 (i_3636, i_2882, i_2891);
  and ginst595 (i_3637, i_1482, i_2891);
  and ginst596 (i_3638, i_109, i_1743, i_3075);
  and ginst597 (i_3639, i_2882, i_2891);
  and ginst598 (i_3640, i_1482, i_2891);
  and ginst599 (i_3641, i_11, i_1339, i_2779);
  and ginst600 (i_3642, i_109, i_1709, i_3041);
  and ginst601 (i_3643, i_46, i_1709, i_3041);
  and ginst602 (i_3644, i_100, i_1709, i_3041);
  and ginst603 (i_3645, i_91, i_1709, i_3041);
  and ginst604 (i_3646, i_43, i_1709, i_3041);
  and ginst605 (i_3647, i_76, i_1339, i_2779);
  and ginst606 (i_3648, i_73, i_1339, i_2779);
  and ginst607 (i_3649, i_67, i_1339, i_2779);
  and ginst608 (i_3650, i_14, i_1339, i_2779);
  and ginst609 (i_3651, i_46, i_1743, i_3075);
  and ginst610 (i_3652, i_100, i_1743, i_3075);
  and ginst611 (i_3653, i_91, i_1743, i_3075);
  and ginst612 (i_3654, i_43, i_1743, i_3075);
  and ginst613 (i_3655, i_76, i_1363, i_2801);
  and ginst614 (i_3656, i_73, i_1363, i_2801);
  and ginst615 (i_3657, i_67, i_1363, i_2801);
  and ginst616 (i_3658, i_14, i_1363, i_2801);
  and ginst617 (i_3659, i_120, i_1785, i_3119);
  and ginst618 (i_3660, i_11, i_1363, i_2801);
  and ginst619 (i_3661, i_118, i_1769, i_3097);
  and ginst620 (i_3662, i_176, i_1197, i_2681);
  and ginst621 (i_3663, i_176, i_1259, i_2756);
  or ginst622 (i_3664, i_2831, i_3401);
  or ginst623 (i_3665, i_2832, i_3402);
  or ginst624 (i_3666, i_2833, i_3403);
  or ginst625 (i_3667, i_2834, i_3404);
  or ginst626 (i_3668, i_457, i_2835, i_3405);
  or ginst627 (i_3669, i_468, i_2836, i_3406);
  or ginst628 (i_3670, i_422, i_2837, i_3407);
  or ginst629 (i_3671, i_435, i_2838, i_3408);
  or ginst630 (i_3672, i_2847, i_3409);
  or ginst631 (i_3673, i_2848, i_3410);
  or ginst632 (i_3674, i_2849, i_3411);
  or ginst633 (i_3675, i_2850, i_3412);
  or ginst634 (i_3676, i_389, i_2851, i_3413);
  or ginst635 (i_3677, i_400, i_2852, i_3414);
  or ginst636 (i_3678, i_411, i_2853, i_3415);
  or ginst637 (i_3679, i_374, i_2854, i_3416);
  and ginst638 (i_3680, i_289, i_2855);
  and ginst639 (i_3681, i_281, i_2855);
  and ginst640 (i_3682, i_273, i_2855);
  and ginst641 (i_3683, i_265, i_2855);
  and ginst642 (i_3684, i_257, i_2855);
  and ginst643 (i_3685, i_234, i_2861);
  and ginst644 (i_3686, i_226, i_2861);
  and ginst645 (i_3687, i_218, i_2861);
  and ginst646 (i_3688, i_210, i_2861);
  and ginst647 (i_3689, i_206, i_2861);
  not ginst648 (i_3691, i_2891);
  or ginst649 (i_3700, i_2907, i_3444);
  or ginst650 (i_3701, i_2908, i_3445);
  or ginst651 (i_3702, i_2909, i_3446);
  or ginst652 (i_3703, i_479, i_2911, i_3448);
  or ginst653 (i_3704, i_490, i_2912, i_3449);
  or ginst654 (i_3705, i_2910, i_3447);
  or ginst655 (i_3708, i_2919, i_3450);
  or ginst656 (i_3709, i_2921, i_3451);
  or ginst657 (i_3710, i_2922, i_3452);
  or ginst658 (i_3711, i_503, i_2923, i_3453);
  or ginst659 (i_3712, i_523, i_2924, i_3454);
  or ginst660 (i_3713, i_534, i_2925, i_3455);
  or ginst661 (i_3715, i_2934, i_3459);
  or ginst662 (i_3716, i_2935, i_3460);
  or ginst663 (i_3717, i_2936, i_3461);
  or ginst664 (i_3718, i_2937, i_3462);
  or ginst665 (i_3719, i_389, i_2938, i_3463);
  or ginst666 (i_3720, i_400, i_2939, i_3464);
  or ginst667 (i_3721, i_411, i_2940, i_3465);
  or ginst668 (i_3722, i_374, i_2941, i_3466);
  and ginst669 (i_3723, i_369, i_2942);
  and ginst670 (i_3724, i_361, i_2942);
  and ginst671 (i_3725, i_351, i_2942);
  and ginst672 (i_3726, i_341, i_2942);
  and ginst673 (i_3727, i_324, i_2948);
  and ginst674 (i_3728, i_316, i_2948);
  and ginst675 (i_3729, i_308, i_2948);
  and ginst676 (i_3730, i_302, i_2948);
  and ginst677 (i_3731, i_293, i_2948);
  or ginst678 (i_3732, i_2942, i_2958);
  and ginst679 (i_3738, i_83, i_2964);
  and ginst680 (i_3739, i_87, i_2964);
  and ginst681 (i_3740, i_34, i_2964);
  and ginst682 (i_3741, i_34, i_2964);
  or ginst683 (i_3742, i_2979, i_3481);
  or ginst684 (i_3743, i_2981, i_3483);
  or ginst685 (i_3744, i_2982, i_3484);
  or ginst686 (i_3745, i_503, i_2983, i_3485);
  or ginst687 (i_3746, i_523, i_2985, i_3486);
  or ginst688 (i_3747, i_534, i_2986, i_3487);
  or ginst689 (i_3748, i_2993, i_3488);
  or ginst690 (i_3749, i_2994, i_3489);
  or ginst691 (i_3750, i_2995, i_3490);
  or ginst692 (i_3751, i_479, i_2997, i_3492);
  or ginst693 (i_3752, i_490, i_2998, i_3493);
  not ginst694 (i_3753, i_3000);
  not ginst695 (i_3754, i_3003);
  not ginst696 (i_3755, i_3007);
  not ginst697 (i_3756, i_3010);
  or ginst698 (i_3757, i_3013, i_3502);
  and ginst699 (i_3758, i_446, i_1315, i_3003);
  or ginst700 (i_3759, i_3014, i_3503);
  and ginst701 (i_3760, i_446, i_1315, i_3010);
  and ginst702 (i_3761, i_1675, i_3000);
  and ginst703 (i_3762, i_1675, i_3007);
  or ginst704 (i_3763, i_3023, i_3504);
  or ginst705 (i_3764, i_3024, i_3505);
  or ginst706 (i_3765, i_3025, i_3506);
  or ginst707 (i_3766, i_3026, i_3507);
  or ginst708 (i_3767, i_457, i_3027, i_3508);
  or ginst709 (i_3768, i_468, i_3028, i_3509);
  or ginst710 (i_3769, i_422, i_3029, i_3510);
  or ginst711 (i_3770, i_435, i_3030, i_3511);
  nand ginst712 (i_3771, i_3512, i_3513);
  nand ginst713 (i_3775, i_3514, i_3515);
  not ginst714 (i_3779, i_3035);
  not ginst715 (i_3780, i_3038);
  and ginst716 (i_3781, i_117, i_1769, i_3097);
  and ginst717 (i_3782, i_126, i_1769, i_3097);
  and ginst718 (i_3783, i_127, i_1769, i_3097);
  and ginst719 (i_3784, i_128, i_1769, i_3097);
  and ginst720 (i_3785, i_131, i_1785, i_3119);
  and ginst721 (i_3786, i_129, i_1785, i_3119);
  and ginst722 (i_3787, i_119, i_1785, i_3119);
  and ginst723 (i_3788, i_130, i_1785, i_3119);
  nand ginst724 (i_3789, i_3558, i_3559);
  nand ginst725 (i_3793, i_3560, i_3561);
  nand ginst726 (i_3797, i_3562, i_3563);
  and ginst727 (i_3800, i_122, i_1800, i_3147);
  and ginst728 (i_3801, i_113, i_1800, i_3147);
  and ginst729 (i_3802, i_53, i_1800, i_3147);
  and ginst730 (i_3803, i_114, i_1800, i_3147);
  and ginst731 (i_3804, i_115, i_1800, i_3147);
  and ginst732 (i_3805, i_52, i_1814, i_3169);
  and ginst733 (i_3806, i_112, i_1814, i_3169);
  and ginst734 (i_3807, i_116, i_1814, i_3169);
  and ginst735 (i_3808, i_121, i_1814, i_3169);
  and ginst736 (i_3809, i_123, i_1814, i_3169);
  nand ginst737 (i_3810, i_3607, i_3608);
  nand ginst738 (i_3813, i_3605, i_3606);
  and ginst739 (i_3816, i_2984, i_3482);
  or ginst740 (i_3819, i_2996, i_3491);
  not ginst741 (i_3822, i_3200);
  nand ginst742 (i_3823, i_3200, i_3203);
  nand ginst743 (i_3824, i_3609, i_3610);
  not ginst744 (i_3827, i_3456);
  or ginst745 (i_3828, i_2970, i_3739);
  or ginst746 (i_3829, i_2971, i_3740);
  or ginst747 (i_3830, i_2972, i_3741);
  or ginst748 (i_3831, i_2969, i_3738);
  not ginst749 (i_3834, i_3664);
  not ginst750 (i_3835, i_3665);
  not ginst751 (i_3836, i_3666);
  not ginst752 (i_3837, i_3667);
  not ginst753 (i_3838, i_3672);
  not ginst754 (i_3839, i_3673);
  not ginst755 (i_3840, i_3674);
  not ginst756 (i_3841, i_3675);
  or ginst757 (i_3842, i_2868, i_3681);
  or ginst758 (i_3849, i_2869, i_3682);
  or ginst759 (i_3855, i_2870, i_3683);
  or ginst760 (i_3861, i_2871, i_3684);
  or ginst761 (i_3867, i_2872, i_3685);
  or ginst762 (i_3873, i_2873, i_3686);
  or ginst763 (i_3881, i_2874, i_3687);
  or ginst764 (i_3887, i_2875, i_3688);
  or ginst765 (i_3893, i_2876, i_3689);
  not ginst766 (i_3908, i_3701);
  not ginst767 (i_3909, i_3702);
  not ginst768 (i_3911, i_3700);
  not ginst769 (i_3914, i_3708);
  not ginst770 (i_3915, i_3709);
  not ginst771 (i_3916, i_3710);
  not ginst772 (i_3917, i_3715);
  not ginst773 (i_3918, i_3716);
  not ginst774 (i_3919, i_3717);
  not ginst775 (i_3920, i_3718);
  or ginst776 (i_3921, i_2955, i_3724);
  or ginst777 (i_3927, i_2956, i_3725);
  or ginst778 (i_3933, i_2957, i_3726);
  or ginst779 (i_3942, i_2959, i_3727);
  or ginst780 (i_3948, i_2960, i_3728);
  or ginst781 (i_3956, i_2961, i_3729);
  or ginst782 (i_3962, i_2962, i_3730);
  or ginst783 (i_3968, i_2963, i_3731);
  not ginst784 (i_3975, i_3742);
  not ginst785 (i_3976, i_3743);
  not ginst786 (i_3977, i_3744);
  not ginst787 (i_3978, i_3749);
  not ginst788 (i_3979, i_3750);
  and ginst789 (i_3980, i_446, i_1292, i_3754);
  and ginst790 (i_3981, i_446, i_1292, i_3756);
  and ginst791 (i_3982, i_1271, i_3753);
  and ginst792 (i_3983, i_1271, i_3755);
  not ginst793 (i_3984, i_3757);
  not ginst794 (i_3987, i_3759);
  not ginst795 (i_3988, i_3763);
  not ginst796 (i_3989, i_3764);
  not ginst797 (i_3990, i_3765);
  not ginst798 (i_3991, i_3766);
  and ginst799 (i_3998, i_3119, i_3130, i_3456);
  or ginst800 (i_4008, i_2954, i_3723);
  or ginst801 (i_4011, i_2867, i_3680);
  not ginst802 (i_4021, i_3748);
  nand ginst803 (i_4024, i_1968, i_3822);
  not ginst804 (i_4027, i_3705);
  and ginst805 (i_4031, i_1583, i_3828);
  and ginst806 (i_4032, i_24, i_2882, i_3691);
  and ginst807 (i_4033, i_25, i_1482, i_3691);
  and ginst808 (i_4034, i_26, i_2882, i_3691);
  and ginst809 (i_4035, i_81, i_1482, i_3691);
  and ginst810 (i_4036, i_1583, i_3829);
  and ginst811 (i_4037, i_79, i_2882, i_3691);
  and ginst812 (i_4038, i_23, i_1482, i_3691);
  and ginst813 (i_4039, i_82, i_2882, i_3691);
  and ginst814 (i_4040, i_80, i_1482, i_3691);
  and ginst815 (i_4041, i_1583, i_3830);
  and ginst816 (i_4042, i_1583, i_3831);
  and ginst817 (i_4067, i_514, i_3732);
  and ginst818 (i_4080, i_514, i_3732);
  and ginst819 (i_4088, i_3668, i_3834);
  and ginst820 (i_4091, i_3669, i_3835);
  and ginst821 (i_4094, i_3670, i_3836);
  and ginst822 (i_4097, i_3671, i_3837);
  and ginst823 (i_4100, i_3676, i_3838);
  and ginst824 (i_4103, i_3677, i_3839);
  and ginst825 (i_4106, i_3678, i_3840);
  and ginst826 (i_4109, i_3679, i_3841);
  and ginst827 (i_4144, i_3703, i_3908);
  and ginst828 (i_4147, i_3704, i_3909);
  not ginst829 (i_4150, i_3705);
  and ginst830 (i_4153, i_3711, i_3914);
  and ginst831 (i_4156, i_3712, i_3915);
  and ginst832 (i_4159, i_3713, i_3916);
  or ginst833 (i_4183, i_3758, i_3980);
  or ginst834 (i_4184, i_3760, i_3981);
  or ginst835 (i_4185, i_446, i_3761, i_3982);
  or ginst836 (i_4186, i_446, i_3762, i_3983);
  not ginst837 (i_4188, i_3771);
  not ginst838 (i_4191, i_3775);
  and ginst839 (i_4196, i_3035, i_3771, i_3775);
  and ginst840 (i_4197, i_3119, i_3130, i_3987);
  and ginst841 (i_4198, i_3722, i_3920);
  not ginst842 (i_4199, i_3816);
  not ginst843 (i_4200, i_3789);
  not ginst844 (i_4203, i_3793);
  not ginst845 (i_4206, i_3797);
  not ginst846 (i_4209, i_3797);
  not ginst847 (i_4212, i_3732);
  not ginst848 (i_4215, i_3732);
  not ginst849 (i_4219, i_3732);
  not ginst850 (i_4223, i_3810);
  not ginst851 (i_4224, i_3813);
  and ginst852 (i_4225, i_3720, i_3918);
  and ginst853 (i_4228, i_3721, i_3919);
  and ginst854 (i_4231, i_3770, i_3991);
  and ginst855 (i_4234, i_3719, i_3917);
  and ginst856 (i_4237, i_3768, i_3989);
  and ginst857 (i_4240, i_3769, i_3990);
  and ginst858 (i_4243, i_3767, i_3988);
  and ginst859 (i_4246, i_3746, i_3976);
  and ginst860 (i_4249, i_3747, i_3977);
  and ginst861 (i_4252, i_3745, i_3975);
  and ginst862 (i_4255, i_3751, i_3978);
  and ginst863 (i_4258, i_3752, i_3979);
  not ginst864 (i_4263, i_3819);
  nand ginst865 (i_4264, i_3823, i_4024);
  not ginst866 (i_4267, i_3824);
  and ginst867 (i_4268, i_446, i_3893);
  not ginst868 (i_4269, i_3911);
  not ginst869 (i_4270, i_3984);
  and ginst870 (i_4271, i_446, i_3893);
  not ginst871 (i_4272, i_4031);
  or ginst872 (i_4273, i_3614, i_3615, i_4032, i_4033);
  or ginst873 (i_4274, i_3625, i_3626, i_4034, i_4035);
  not ginst874 (i_4275, i_4036);
  or ginst875 (i_4276, i_3636, i_3637, i_4037, i_4038);
  or ginst876 (i_4277, i_3639, i_3640, i_4039, i_4040);
  not ginst877 (i_4278, i_4041);
  not ginst878 (i_4279, i_4042);
  and ginst879 (i_4280, i_457, i_3887);
  and ginst880 (i_4284, i_468, i_3881);
  and ginst881 (i_4290, i_422, i_3873);
  and ginst882 (i_4297, i_435, i_3867);
  and ginst883 (i_4298, i_389, i_3861);
  and ginst884 (i_4301, i_400, i_3855);
  and ginst885 (i_4305, i_411, i_3849);
  and ginst886 (i_4310, i_374, i_3842);
  and ginst887 (i_4316, i_457, i_3887);
  and ginst888 (i_4320, i_468, i_3881);
  and ginst889 (i_4325, i_422, i_3873);
  and ginst890 (i_4331, i_435, i_3867);
  and ginst891 (i_4332, i_389, i_3861);
  and ginst892 (i_4336, i_400, i_3855);
  and ginst893 (i_4342, i_411, i_3849);
  and ginst894 (i_4349, i_374, i_3842);
  not ginst895 (i_4357, i_3968);
  not ginst896 (i_4364, i_3962);
  not ginst897 (i_4375, i_3962);
  and ginst898 (i_4379, i_479, i_3956);
  and ginst899 (i_4385, i_490, i_3948);
  and ginst900 (i_4392, i_503, i_3942);
  and ginst901 (i_4396, i_523, i_3933);
  and ginst902 (i_4400, i_534, i_3927);
  not ginst903 (i_4405, i_3921);
  not ginst904 (i_4412, i_3921);
  not ginst905 (i_4418, i_3968);
  not ginst906 (i_4425, i_3962);
  not ginst907 (i_4436, i_3962);
  and ginst908 (i_4440, i_479, i_3956);
  and ginst909 (i_4445, i_490, i_3948);
  and ginst910 (i_4451, i_503, i_3942);
  and ginst911 (i_4456, i_523, i_3933);
  and ginst912 (i_4462, i_534, i_3927);
  not ginst913 (i_4469, i_3921);
  not ginst914 (i_4477, i_3921);
  not ginst915 (i_4512, i_3968);
  not ginst916 (i_4515, i_4183);
  not ginst917 (i_4516, i_4184);
  not ginst918 (i_4521, i_4008);
  not ginst919 (i_4523, i_4011);
  not ginst920 (i_4524, i_4198);
  not ginst921 (i_4532, i_3984);
  and ginst922 (i_4547, i_3169, i_3180, i_3911);
  not ginst923 (i_4548, i_3893);
  not ginst924 (i_4551, i_3887);
  not ginst925 (i_4554, i_3881);
  not ginst926 (i_4557, i_3873);
  not ginst927 (i_4560, i_3867);
  not ginst928 (i_4563, i_3861);
  not ginst929 (i_4566, i_3855);
  not ginst930 (i_4569, i_3849);
  not ginst931 (i_4572, i_3842);
  nor ginst932 (i_4575, i_422, i_3873);
  not ginst933 (i_4578, i_3893);
  not ginst934 (i_4581, i_3887);
  not ginst935 (i_4584, i_3881);
  not ginst936 (i_4587, i_3867);
  not ginst937 (i_4590, i_3861);
  not ginst938 (i_4593, i_3855);
  not ginst939 (i_4596, i_3849);
  not ginst940 (i_4599, i_3873);
  not ginst941 (i_4602, i_3842);
  nor ginst942 (i_4605, i_422, i_3873);
  nor ginst943 (i_4608, i_374, i_3842);
  not ginst944 (i_4611, i_3956);
  not ginst945 (i_4614, i_3948);
  not ginst946 (i_4617, i_3942);
  not ginst947 (i_4621, i_3933);
  not ginst948 (i_4624, i_3927);
  nor ginst949 (i_4627, i_490, i_3948);
  not ginst950 (i_4630, i_3956);
  not ginst951 (i_4633, i_3942);
  not ginst952 (i_4637, i_3933);
  not ginst953 (i_4640, i_3927);
  not ginst954 (i_4643, i_3948);
  nor ginst955 (i_4646, i_490, i_3948);
  not ginst956 (i_4649, i_3927);
  not ginst957 (i_4652, i_3933);
  not ginst958 (i_4655, i_3921);
  not ginst959 (i_4658, i_3942);
  not ginst960 (i_4662, i_3956);
  not ginst961 (i_4665, i_3948);
  not ginst962 (i_4668, i_3968);
  not ginst963 (i_4671, i_3962);
  not ginst964 (i_4674, i_3873);
  not ginst965 (i_4677, i_3867);
  not ginst966 (i_4680, i_3887);
  not ginst967 (i_4683, i_3881);
  not ginst968 (i_4686, i_3893);
  not ginst969 (i_4689, i_3849);
  not ginst970 (i_4692, i_3842);
  not ginst971 (i_4695, i_3861);
  not ginst972 (i_4698, i_3855);
  nand ginst973 (i_4701, i_3813, i_4223);
  nand ginst974 (i_4702, i_3810, i_4224);
  not ginst975 (i_4720, i_4021);
  nand ginst976 (i_4721, i_4021, i_4263);
  not ginst977 (i_4724, i_4147);
  not ginst978 (i_4725, i_4144);
  not ginst979 (i_4726, i_4159);
  not ginst980 (i_4727, i_4156);
  not ginst981 (i_4728, i_4153);
  not ginst982 (i_4729, i_4097);
  not ginst983 (i_4730, i_4094);
  not ginst984 (i_4731, i_4091);
  not ginst985 (i_4732, i_4088);
  not ginst986 (i_4733, i_4109);
  not ginst987 (i_4734, i_4106);
  not ginst988 (i_4735, i_4103);
  not ginst989 (i_4736, i_4100);
  and ginst990 (i_4737, i_2877, i_4273);
  and ginst991 (i_4738, i_2877, i_4274);
  and ginst992 (i_4739, i_2877, i_4276);
  and ginst993 (i_4740, i_2877, i_4277);
  and ginst994 (i_4741, i_1755, i_1758, i_4150);
  not ginst995 (i_4855, i_4212);
  nand ginst996 (i_4856, i_2712, i_4212);
  nand ginst997 (i_4908, i_2718, i_4215);
  not ginst998 (i_4909, i_4215);
  and ginst999 (i_4939, i_4185, i_4515);
  and ginst1000 (i_4942, i_4186, i_4516);
  not ginst1001 (i_4947, i_4219);
  and ginst1002 (i_4953, i_3775, i_3779, i_4188);
  and ginst1003 (i_4954, i_3771, i_3780, i_4191);
  and ginst1004 (i_4955, i_3038, i_4188, i_4191);
  and ginst1005 (i_4956, i_3097, i_3108, i_4109);
  and ginst1006 (i_4957, i_3097, i_3108, i_4106);
  and ginst1007 (i_4958, i_3097, i_3108, i_4103);
  and ginst1008 (i_4959, i_3097, i_3108, i_4100);
  and ginst1009 (i_4960, i_3119, i_3130, i_4159);
  and ginst1010 (i_4961, i_3119, i_3130, i_4156);
  not ginst1011 (i_4965, i_4225);
  not ginst1012 (i_4966, i_4228);
  not ginst1013 (i_4967, i_4231);
  not ginst1014 (i_4968, i_4234);
  not ginst1015 (i_4972, i_4246);
  not ginst1016 (i_4973, i_4249);
  not ginst1017 (i_4974, i_4252);
  nand ginst1018 (i_4975, i_4199, i_4252);
  not ginst1019 (i_4976, i_4206);
  not ginst1020 (i_4977, i_4209);
  and ginst1021 (i_4978, i_3789, i_3793, i_4206);
  and ginst1022 (i_4979, i_4200, i_4203, i_4209);
  and ginst1023 (i_4980, i_3147, i_3158, i_4097);
  and ginst1024 (i_4981, i_3147, i_3158, i_4094);
  and ginst1025 (i_4982, i_3147, i_3158, i_4091);
  and ginst1026 (i_4983, i_3147, i_3158, i_4088);
  and ginst1027 (i_4984, i_3169, i_3180, i_4153);
  and ginst1028 (i_4985, i_3169, i_3180, i_4147);
  and ginst1029 (i_4986, i_3169, i_3180, i_4144);
  and ginst1030 (i_4987, i_3169, i_3180, i_4150);
  nand ginst1031 (i_5049, i_4701, i_4702);
  not ginst1032 (i_5052, i_4237);
  not ginst1033 (i_5053, i_4240);
  not ginst1034 (i_5054, i_4243);
  not ginst1035 (i_5055, i_4255);
  not ginst1036 (i_5056, i_4258);
  nand ginst1037 (i_5057, i_3819, i_4720);
  not ginst1038 (i_5058, i_4264);
  nand ginst1039 (i_5059, i_4264, i_4267);
  and ginst1040 (i_5060, i_4027, i_4269, i_4724, i_4725);
  and ginst1041 (i_5061, i_3827, i_4726, i_4727, i_4728);
  and ginst1042 (i_5062, i_4729, i_4730, i_4731, i_4732);
  and ginst1043 (i_5063, i_4733, i_4734, i_4735, i_4736);
  and ginst1044 (i_5065, i_4357, i_4375);
  and ginst1045 (i_5066, i_4357, i_4364, i_4379);
  and ginst1046 (i_5067, i_4418, i_4436);
  and ginst1047 (i_5068, i_4418, i_4425, i_4440);
  not ginst1048 (i_5069, i_4548);
  nand ginst1049 (i_5070, i_2628, i_4548);
  not ginst1050 (i_5071, i_4551);
  nand ginst1051 (i_5072, i_2629, i_4551);
  not ginst1052 (i_5073, i_4554);
  nand ginst1053 (i_5074, i_2630, i_4554);
  not ginst1054 (i_5075, i_4557);
  nand ginst1055 (i_5076, i_2631, i_4557);
  not ginst1056 (i_5077, i_4560);
  nand ginst1057 (i_5078, i_2632, i_4560);
  not ginst1058 (i_5079, i_4563);
  nand ginst1059 (i_5080, i_2633, i_4563);
  not ginst1060 (i_5081, i_4566);
  nand ginst1061 (i_5082, i_2634, i_4566);
  not ginst1062 (i_5083, i_4569);
  nand ginst1063 (i_5084, i_2635, i_4569);
  not ginst1064 (i_5085, i_4572);
  nand ginst1065 (i_5086, i_2636, i_4572);
  not ginst1066 (i_5087, i_4575);
  nand ginst1067 (i_5088, i_2638, i_4578);
  not ginst1068 (i_5089, i_4578);
  nand ginst1069 (i_5090, i_2639, i_4581);
  not ginst1070 (i_5091, i_4581);
  nand ginst1071 (i_5092, i_2640, i_4584);
  not ginst1072 (i_5093, i_4584);
  nand ginst1073 (i_5094, i_2641, i_4587);
  not ginst1074 (i_5095, i_4587);
  nand ginst1075 (i_5096, i_2642, i_4590);
  not ginst1076 (i_5097, i_4590);
  nand ginst1077 (i_5098, i_2643, i_4593);
  not ginst1078 (i_5099, i_4593);
  nand ginst1079 (i_5100, i_2644, i_4596);
  not ginst1080 (i_5101, i_4596);
  nand ginst1081 (i_5102, i_2645, i_4599);
  not ginst1082 (i_5103, i_4599);
  nand ginst1083 (i_5104, i_2646, i_4602);
  not ginst1084 (i_5105, i_4602);
  not ginst1085 (i_5106, i_4611);
  nand ginst1086 (i_5107, i_2709, i_4611);
  not ginst1087 (i_5108, i_4614);
  nand ginst1088 (i_5109, i_2710, i_4614);
  not ginst1089 (i_5110, i_4617);
  nand ginst1090 (i_5111, i_2711, i_4617);
  nand ginst1091 (i_5112, i_1890, i_4855);
  not ginst1092 (i_5113, i_4621);
  nand ginst1093 (i_5114, i_2713, i_4621);
  not ginst1094 (i_5115, i_4624);
  nand ginst1095 (i_5116, i_2714, i_4624);
  and ginst1096 (i_5117, i_4364, i_4379);
  and ginst1097 (i_5118, i_4364, i_4379);
  and ginst1098 (i_5119, i_54, i_4405);
  not ginst1099 (i_5120, i_4627);
  nand ginst1100 (i_5121, i_2716, i_4630);
  not ginst1101 (i_5122, i_4630);
  nand ginst1102 (i_5123, i_2717, i_4633);
  not ginst1103 (i_5124, i_4633);
  nand ginst1104 (i_5125, i_1908, i_4909);
  nand ginst1105 (i_5126, i_2719, i_4637);
  not ginst1106 (i_5127, i_4637);
  nand ginst1107 (i_5128, i_2720, i_4640);
  not ginst1108 (i_5129, i_4640);
  nand ginst1109 (i_5130, i_2721, i_4643);
  not ginst1110 (i_5131, i_4643);
  and ginst1111 (i_5132, i_4425, i_4440);
  and ginst1112 (i_5133, i_4425, i_4440);
  not ginst1113 (i_5135, i_4649);
  not ginst1114 (i_5136, i_4652);
  nand ginst1115 (i_5137, i_4521, i_4655);
  not ginst1116 (i_5138, i_4655);
  not ginst1117 (i_5139, i_4658);
  nand ginst1118 (i_5140, i_4658, i_4947);
  not ginst1119 (i_5141, i_4674);
  not ginst1120 (i_5142, i_4677);
  not ginst1121 (i_5143, i_4680);
  not ginst1122 (i_5144, i_4683);
  nand ginst1123 (i_5145, i_4523, i_4686);
  not ginst1124 (i_5146, i_4686);
  nor ginst1125 (i_5147, i_4196, i_4953);
  nor ginst1126 (i_5148, i_4954, i_4955);
  not ginst1127 (i_5150, i_4524);
  nand ginst1128 (i_5153, i_4228, i_4965);
  nand ginst1129 (i_5154, i_4225, i_4966);
  nand ginst1130 (i_5155, i_4234, i_4967);
  nand ginst1131 (i_5156, i_4231, i_4968);
  not ginst1132 (i_5157, i_4532);
  nand ginst1133 (i_5160, i_4249, i_4972);
  nand ginst1134 (i_5161, i_4246, i_4973);
  nand ginst1135 (i_5162, i_3816, i_4974);
  and ginst1136 (i_5163, i_3793, i_4200, i_4976);
  and ginst1137 (i_5164, i_3789, i_4203, i_4977);
  and ginst1138 (i_5165, i_3147, i_3158, i_4942);
  not ginst1139 (i_5166, i_4512);
  not ginst1140 (i_5169, i_4290);
  not ginst1141 (i_5172, i_4605);
  not ginst1142 (i_5173, i_4325);
  not ginst1143 (i_5176, i_4608);
  not ginst1144 (i_5177, i_4349);
  not ginst1145 (i_5180, i_4405);
  not ginst1146 (i_5183, i_4357);
  not ginst1147 (i_5186, i_4357);
  not ginst1148 (i_5189, i_4364);
  not ginst1149 (i_5192, i_4364);
  not ginst1150 (i_5195, i_4385);
  not ginst1151 (i_5198, i_4646);
  not ginst1152 (i_5199, i_4418);
  not ginst1153 (i_5202, i_4425);
  not ginst1154 (i_5205, i_4445);
  not ginst1155 (i_5208, i_4418);
  not ginst1156 (i_5211, i_4425);
  not ginst1157 (i_5214, i_4477);
  not ginst1158 (i_5217, i_4469);
  not ginst1159 (i_5220, i_4477);
  not ginst1160 (i_5223, i_4662);
  not ginst1161 (i_5224, i_4665);
  not ginst1162 (i_5225, i_4668);
  not ginst1163 (i_5226, i_4671);
  not ginst1164 (i_5227, i_4689);
  not ginst1165 (i_5228, i_4692);
  not ginst1166 (i_5229, i_4695);
  not ginst1167 (i_5230, i_4698);
  nand ginst1168 (i_5232, i_4240, i_5052);
  nand ginst1169 (i_5233, i_4237, i_5053);
  nand ginst1170 (i_5234, i_4258, i_5055);
  nand ginst1171 (i_5235, i_4255, i_5056);
  nand ginst1172 (i_5236, i_4721, i_5057);
  nand ginst1173 (i_5239, i_3824, i_5058);
  and ginst1174 (i_5240, i_4270, i_5060, i_5061);
  not ginst1175 (i_5241, i_4939);
  nand ginst1176 (i_5242, i_1824, i_5069);
  nand ginst1177 (i_5243, i_1827, i_5071);
  nand ginst1178 (i_5244, i_1830, i_5073);
  nand ginst1179 (i_5245, i_1833, i_5075);
  nand ginst1180 (i_5246, i_1836, i_5077);
  nand ginst1181 (i_5247, i_1839, i_5079);
  nand ginst1182 (i_5248, i_1842, i_5081);
  nand ginst1183 (i_5249, i_1845, i_5083);
  nand ginst1184 (i_5250, i_1848, i_5085);
  nand ginst1185 (i_5252, i_1854, i_5089);
  nand ginst1186 (i_5253, i_1857, i_5091);
  nand ginst1187 (i_5254, i_1860, i_5093);
  nand ginst1188 (i_5255, i_1863, i_5095);
  nand ginst1189 (i_5256, i_1866, i_5097);
  nand ginst1190 (i_5257, i_1869, i_5099);
  nand ginst1191 (i_5258, i_1872, i_5101);
  nand ginst1192 (i_5259, i_1875, i_5103);
  nand ginst1193 (i_5260, i_1878, i_5105);
  nand ginst1194 (i_5261, i_1881, i_5106);
  nand ginst1195 (i_5262, i_1884, i_5108);
  nand ginst1196 (i_5263, i_1887, i_5110);
  nand ginst1197 (i_5264, i_4856, i_5112);
  nand ginst1198 (i_5274, i_1893, i_5113);
  nand ginst1199 (i_5275, i_1896, i_5115);
  nand ginst1200 (i_5282, i_1902, i_5122);
  nand ginst1201 (i_5283, i_1905, i_5124);
  nand ginst1202 (i_5284, i_4908, i_5125);
  nand ginst1203 (i_5298, i_1911, i_5127);
  nand ginst1204 (i_5299, i_1914, i_5129);
  nand ginst1205 (i_5300, i_1917, i_5131);
  nand ginst1206 (i_5303, i_4652, i_5135);
  nand ginst1207 (i_5304, i_4649, i_5136);
  nand ginst1208 (i_5305, i_4008, i_5138);
  nand ginst1209 (i_5306, i_4219, i_5139);
  nand ginst1210 (i_5307, i_4677, i_5141);
  nand ginst1211 (i_5308, i_4674, i_5142);
  nand ginst1212 (i_5309, i_4683, i_5143);
  nand ginst1213 (i_5310, i_4680, i_5144);
  nand ginst1214 (i_5311, i_4011, i_5146);
  not ginst1215 (i_5312, i_5049);
  nand ginst1216 (i_5315, i_5153, i_5154);
  nand ginst1217 (i_5319, i_5155, i_5156);
  nand ginst1218 (i_5324, i_5160, i_5161);
  nand ginst1219 (i_5328, i_4975, i_5162);
  nor ginst1220 (i_5331, i_4978, i_5163);
  nor ginst1221 (i_5332, i_4979, i_5164);
  or ginst1222 (i_5346, i_4412, i_5119);
  nand ginst1223 (i_5363, i_4665, i_5223);
  nand ginst1224 (i_5364, i_4662, i_5224);
  nand ginst1225 (i_5365, i_4671, i_5225);
  nand ginst1226 (i_5366, i_4668, i_5226);
  nand ginst1227 (i_5367, i_4692, i_5227);
  nand ginst1228 (i_5368, i_4689, i_5228);
  nand ginst1229 (i_5369, i_4698, i_5229);
  nand ginst1230 (i_5370, i_4695, i_5230);
  nand ginst1231 (i_5371, i_5147, i_5148);
  not ginst1232 (i_5374, i_4939);
  nand ginst1233 (i_5377, i_5232, i_5233);
  nand ginst1234 (i_5382, i_5234, i_5235);
  nand ginst1235 (i_5385, i_5059, i_5239);
  and ginst1236 (i_5388, i_5062, i_5063, i_5241);
  nand ginst1237 (i_5389, i_5070, i_5242);
  nand ginst1238 (i_5396, i_5072, i_5243);
  nand ginst1239 (i_5407, i_5074, i_5244);
  nand ginst1240 (i_5418, i_5076, i_5245);
  nand ginst1241 (i_5424, i_5078, i_5246);
  nand ginst1242 (i_5431, i_5080, i_5247);
  nand ginst1243 (i_5441, i_5082, i_5248);
  nand ginst1244 (i_5452, i_5084, i_5249);
  nand ginst1245 (i_5462, i_5086, i_5250);
  not ginst1246 (i_5469, i_5169);
  nand ginst1247 (i_5470, i_5088, i_5252);
  nand ginst1248 (i_5477, i_5090, i_5253);
  nand ginst1249 (i_5488, i_5092, i_5254);
  nand ginst1250 (i_5498, i_5094, i_5255);
  nand ginst1251 (i_5506, i_5096, i_5256);
  nand ginst1252 (i_5520, i_5098, i_5257);
  nand ginst1253 (i_5536, i_5100, i_5258);
  nand ginst1254 (i_5549, i_5102, i_5259);
  nand ginst1255 (i_5555, i_5104, i_5260);
  nand ginst1256 (i_5562, i_5107, i_5261);
  nand ginst1257 (i_5573, i_5109, i_5262);
  nand ginst1258 (i_5579, i_5111, i_5263);
  nand ginst1259 (i_5595, i_5114, i_5274);
  nand ginst1260 (i_5606, i_5116, i_5275);
  nand ginst1261 (i_5616, i_2715, i_5180);
  not ginst1262 (i_5617, i_5180);
  not ginst1263 (i_5618, i_5183);
  not ginst1264 (i_5619, i_5186);
  not ginst1265 (i_5620, i_5189);
  not ginst1266 (i_5621, i_5192);
  not ginst1267 (i_5622, i_5195);
  nand ginst1268 (i_5624, i_5121, i_5282);
  nand ginst1269 (i_5634, i_5123, i_5283);
  nand ginst1270 (i_5655, i_5126, i_5298);
  nand ginst1271 (i_5671, i_5128, i_5299);
  nand ginst1272 (i_5684, i_5130, i_5300);
  not ginst1273 (i_5690, i_5202);
  not ginst1274 (i_5691, i_5211);
  nand ginst1275 (i_5692, i_5303, i_5304);
  nand ginst1276 (i_5696, i_5137, i_5305);
  nand ginst1277 (i_5700, i_5140, i_5306);
  nand ginst1278 (i_5703, i_5307, i_5308);
  nand ginst1279 (i_5707, i_5309, i_5310);
  nand ginst1280 (i_5711, i_5145, i_5311);
  and ginst1281 (i_5726, i_4512, i_5166);
  not ginst1282 (i_5727, i_5173);
  not ginst1283 (i_5728, i_5177);
  not ginst1284 (i_5730, i_5199);
  not ginst1285 (i_5731, i_5205);
  not ginst1286 (i_5732, i_5208);
  not ginst1287 (i_5733, i_5214);
  not ginst1288 (i_5734, i_5217);
  not ginst1289 (i_5735, i_5220);
  nand ginst1290 (i_5736, i_5365, i_5366);
  nand ginst1291 (i_5739, i_5363, i_5364);
  nand ginst1292 (i_5742, i_5369, i_5370);
  nand ginst1293 (i_5745, i_5367, i_5368);
  not ginst1294 (i_5755, i_5236);
  nand ginst1295 (i_5756, i_5331, i_5332);
  and ginst1296 (i_5954, i_4396, i_5264);
  nand ginst1297 (i_5955, i_1899, i_5617);
  not ginst1298 (i_5956, i_5346);
  and ginst1299 (i_6005, i_4456, i_5284);
  and ginst1300 (i_6006, i_4456, i_5284);
  not ginst1301 (i_6023, i_5371);
  nand ginst1302 (i_6024, i_5312, i_5371);
  not ginst1303 (i_6025, i_5315);
  not ginst1304 (i_6028, i_5324);
  not ginst1305 (i_6031, i_5319);
  not ginst1306 (i_6034, i_5319);
  not ginst1307 (i_6037, i_5328);
  not ginst1308 (i_6040, i_5328);
  not ginst1309 (i_6044, i_5385);
  or ginst1310 (i_6045, i_5166, i_5726);
  not ginst1311 (i_6048, i_5264);
  not ginst1312 (i_6051, i_5284);
  not ginst1313 (i_6054, i_5284);
  not ginst1314 (i_6065, i_5374);
  nand ginst1315 (i_6066, i_5054, i_5374);
  not ginst1316 (i_6067, i_5377);
  not ginst1317 (i_6068, i_5382);
  nand ginst1318 (i_6069, i_5382, i_5755);
  and ginst1319 (i_6071, i_4316, i_5470);
  and ginst1320 (i_6072, i_4320, i_5470, i_5477);
  and ginst1321 (i_6073, i_4325, i_5470, i_5477, i_5488);
  and ginst1322 (i_6074, i_4357, i_4364, i_4385, i_5562);
  and ginst1323 (i_6075, i_4280, i_5389);
  and ginst1324 (i_6076, i_4284, i_5389, i_5396);
  and ginst1325 (i_6077, i_4290, i_5389, i_5396, i_5407);
  and ginst1326 (i_6078, i_4418, i_4425, i_4445, i_5624);
  not ginst1327 (i_6079, i_5418);
  and ginst1328 (i_6080, i_5389, i_5396, i_5407, i_5418);
  and ginst1329 (i_6083, i_4284, i_5396);
  and ginst1330 (i_6084, i_4290, i_5396, i_5407);
  and ginst1331 (i_6085, i_5396, i_5407, i_5418);
  and ginst1332 (i_6086, i_4284, i_5396);
  and ginst1333 (i_6087, i_4290, i_5396, i_5407);
  and ginst1334 (i_6088, i_4290, i_5407);
  and ginst1335 (i_6089, i_5407, i_5418);
  and ginst1336 (i_6090, i_4290, i_5407);
  and ginst1337 (i_6091, i_5424, i_5431, i_5441, i_5452, i_5462);
  and ginst1338 (i_6094, i_4298, i_5424);
  and ginst1339 (i_6095, i_4301, i_5424, i_5431);
  and ginst1340 (i_6096, i_4305, i_5424, i_5431, i_5441);
  and ginst1341 (i_6097, i_4310, i_5424, i_5431, i_5441, i_5452);
  and ginst1342 (i_6098, i_4301, i_5431);
  and ginst1343 (i_6099, i_4305, i_5431, i_5441);
  and ginst1344 (i_6100, i_4310, i_5431, i_5441, i_5452);
  and ginst1345 (i_6101, i_4, i_5431, i_5441, i_5452, i_5462);
  and ginst1346 (i_6102, i_4305, i_5441);
  and ginst1347 (i_6103, i_4310, i_5441, i_5452);
  and ginst1348 (i_6104, i_4, i_5441, i_5452, i_5462);
  and ginst1349 (i_6105, i_4310, i_5452);
  and ginst1350 (i_6106, i_4, i_5452, i_5462);
  and ginst1351 (i_6107, i_4, i_5462);
  and ginst1352 (i_6108, i_5470, i_5477, i_5488, i_5549);
  and ginst1353 (i_6111, i_4320, i_5477);
  and ginst1354 (i_6112, i_4325, i_5477, i_5488);
  and ginst1355 (i_6113, i_5477, i_5488, i_5549);
  and ginst1356 (i_6114, i_4320, i_5477);
  and ginst1357 (i_6115, i_4325, i_5477, i_5488);
  and ginst1358 (i_6116, i_4325, i_5488);
  and ginst1359 (i_6117, i_5498, i_5506, i_5520, i_5536, i_5555);
  and ginst1360 (i_6120, i_4332, i_5498);
  and ginst1361 (i_6121, i_4336, i_5498, i_5506);
  and ginst1362 (i_6122, i_4342, i_5498, i_5506, i_5520);
  and ginst1363 (i_6123, i_4349, i_5498, i_5506, i_5520, i_5536);
  and ginst1364 (i_6124, i_4336, i_5506);
  and ginst1365 (i_6125, i_4342, i_5506, i_5520);
  and ginst1366 (i_6126, i_4349, i_5506, i_5520, i_5536);
  and ginst1367 (i_6127, i_5506, i_5520, i_5536, i_5555);
  and ginst1368 (i_6128, i_4336, i_5506);
  and ginst1369 (i_6129, i_4342, i_5506, i_5520);
  and ginst1370 (i_6130, i_4349, i_5506, i_5520, i_5536);
  and ginst1371 (i_6131, i_4342, i_5520);
  and ginst1372 (i_6132, i_4349, i_5520, i_5536);
  and ginst1373 (i_6133, i_5520, i_5536, i_5555);
  and ginst1374 (i_6134, i_4342, i_5520);
  and ginst1375 (i_6135, i_4349, i_5520, i_5536);
  and ginst1376 (i_6136, i_4349, i_5536);
  and ginst1377 (i_6137, i_5488, i_5549);
  and ginst1378 (i_6138, i_5536, i_5555);
  not ginst1379 (i_6139, i_5573);
  and ginst1380 (i_6140, i_4357, i_4364, i_5562, i_5573);
  and ginst1381 (i_6143, i_4364, i_4385, i_5562);
  and ginst1382 (i_6144, i_4364, i_5562, i_5573);
  and ginst1383 (i_6145, i_4364, i_4385, i_5562);
  and ginst1384 (i_6146, i_4385, i_5562);
  and ginst1385 (i_6147, i_5562, i_5573);
  and ginst1386 (i_6148, i_4385, i_5562);
  and ginst1387 (i_6149, i_4405, i_5264, i_5579, i_5595, i_5606);
  and ginst1388 (i_6152, i_4067, i_5579);
  and ginst1389 (i_6153, i_4396, i_5264, i_5579);
  and ginst1390 (i_6154, i_4400, i_5264, i_5579, i_5595);
  and ginst1391 (i_6155, i_4412, i_5264, i_5579, i_5595, i_5606);
  and ginst1392 (i_6156, i_4400, i_5264, i_5595);
  and ginst1393 (i_6157, i_4412, i_5264, i_5595, i_5606);
  and ginst1394 (i_6158, i_54, i_4405, i_5264, i_5595, i_5606);
  and ginst1395 (i_6159, i_4400, i_5595);
  and ginst1396 (i_6160, i_4412, i_5595, i_5606);
  and ginst1397 (i_6161, i_54, i_4405, i_5595, i_5606);
  and ginst1398 (i_6162, i_4412, i_5606);
  and ginst1399 (i_6163, i_54, i_4405, i_5606);
  nand ginst1400 (i_6164, i_5616, i_5955);
  and ginst1401 (i_6168, i_4418, i_4425, i_5624, i_5684);
  and ginst1402 (i_6171, i_4425, i_4445, i_5624);
  and ginst1403 (i_6172, i_4425, i_5624, i_5684);
  and ginst1404 (i_6173, i_4425, i_4445, i_5624);
  and ginst1405 (i_6174, i_4445, i_5624);
  and ginst1406 (i_6175, i_4477, i_5284, i_5634, i_5655, i_5671);
  and ginst1407 (i_6178, i_4080, i_5634);
  and ginst1408 (i_6179, i_4456, i_5284, i_5634);
  and ginst1409 (i_6180, i_4462, i_5284, i_5634, i_5655);
  and ginst1410 (i_6181, i_4469, i_5284, i_5634, i_5655, i_5671);
  and ginst1411 (i_6182, i_4462, i_5284, i_5655);
  and ginst1412 (i_6183, i_4469, i_5284, i_5655, i_5671);
  and ginst1413 (i_6184, i_4477, i_5284, i_5655, i_5671);
  and ginst1414 (i_6185, i_4462, i_5284, i_5655);
  and ginst1415 (i_6186, i_4469, i_5284, i_5655, i_5671);
  and ginst1416 (i_6187, i_4462, i_5655);
  and ginst1417 (i_6188, i_4469, i_5655, i_5671);
  and ginst1418 (i_6189, i_4477, i_5655, i_5671);
  and ginst1419 (i_6190, i_4462, i_5655);
  and ginst1420 (i_6191, i_4469, i_5655, i_5671);
  and ginst1421 (i_6192, i_4469, i_5671);
  and ginst1422 (i_6193, i_5624, i_5684);
  and ginst1423 (i_6194, i_4477, i_5671);
  not ginst1424 (i_6197, i_5692);
  not ginst1425 (i_6200, i_5696);
  not ginst1426 (i_6203, i_5703);
  not ginst1427 (i_6206, i_5707);
  not ginst1428 (i_6209, i_5700);
  not ginst1429 (i_6212, i_5700);
  not ginst1430 (i_6215, i_5711);
  not ginst1431 (i_6218, i_5711);
  nand ginst1432 (i_6221, i_5049, i_6023);
  not ginst1433 (i_6234, i_5756);
  nand ginst1434 (i_6235, i_5756, i_6044);
  not ginst1435 (i_6238, i_5462);
  not ginst1436 (i_6241, i_5389);
  not ginst1437 (i_6244, i_5389);
  not ginst1438 (i_6247, i_5396);
  not ginst1439 (i_6250, i_5396);
  not ginst1440 (i_6253, i_5407);
  not ginst1441 (i_6256, i_5407);
  not ginst1442 (i_6259, i_5424);
  not ginst1443 (i_6262, i_5431);
  not ginst1444 (i_6265, i_5441);
  not ginst1445 (i_6268, i_5452);
  not ginst1446 (i_6271, i_5549);
  not ginst1447 (i_6274, i_5488);
  not ginst1448 (i_6277, i_5470);
  not ginst1449 (i_6280, i_5477);
  not ginst1450 (i_6283, i_5549);
  not ginst1451 (i_6286, i_5488);
  not ginst1452 (i_6289, i_5470);
  not ginst1453 (i_6292, i_5477);
  not ginst1454 (i_6295, i_5555);
  not ginst1455 (i_6298, i_5536);
  not ginst1456 (i_6301, i_5498);
  not ginst1457 (i_6304, i_5520);
  not ginst1458 (i_6307, i_5506);
  not ginst1459 (i_6310, i_5506);
  not ginst1460 (i_6313, i_5555);
  not ginst1461 (i_6316, i_5536);
  not ginst1462 (i_6319, i_5498);
  not ginst1463 (i_6322, i_5520);
  not ginst1464 (i_6325, i_5562);
  not ginst1465 (i_6328, i_5562);
  not ginst1466 (i_6331, i_5579);
  not ginst1467 (i_6335, i_5595);
  not ginst1468 (i_6338, i_5606);
  not ginst1469 (i_6341, i_5684);
  not ginst1470 (i_6344, i_5624);
  not ginst1471 (i_6347, i_5684);
  not ginst1472 (i_6350, i_5624);
  not ginst1473 (i_6353, i_5671);
  not ginst1474 (i_6356, i_5634);
  not ginst1475 (i_6359, i_5655);
  not ginst1476 (i_6364, i_5671);
  not ginst1477 (i_6367, i_5634);
  not ginst1478 (i_6370, i_5655);
  not ginst1479 (i_6373, i_5736);
  not ginst1480 (i_6374, i_5739);
  not ginst1481 (i_6375, i_5742);
  not ginst1482 (i_6376, i_5745);
  nand ginst1483 (i_6377, i_4243, i_6065);
  nand ginst1484 (i_6378, i_5236, i_6068);
  or ginst1485 (i_6382, i_4268, i_6071, i_6072, i_6073);
  or ginst1486 (i_6386, i_3968, i_5065, i_5066, i_6074);
  or ginst1487 (i_6388, i_4271, i_6075, i_6076, i_6077);
  or ginst1488 (i_6392, i_3968, i_5067, i_5068, i_6078);
  or ginst1489 (i_6397, i_4297, i_6094, i_6095, i_6096, i_6097);
  or ginst1490 (i_6411, i_4320, i_6116);
  or ginst1491 (i_6415, i_4331, i_6120, i_6121, i_6122, i_6123);
  or ginst1492 (i_6419, i_4342, i_6136);
  or ginst1493 (i_6427, i_4392, i_6152, i_6153, i_6154, i_6155);
  not ginst1494 (i_6434, i_6048);
  or ginst1495 (i_6437, i_4440, i_6174);
  or ginst1496 (i_6441, i_4451, i_6178, i_6179, i_6180, i_6181);
  or ginst1497 (i_6445, i_4462, i_6192);
  not ginst1498 (i_6448, i_6051);
  not ginst1499 (i_6449, i_6054);
  nand ginst1500 (i_6466, i_6024, i_6221);
  not ginst1501 (i_6469, i_6031);
  not ginst1502 (i_6470, i_6034);
  not ginst1503 (i_6471, i_6037);
  not ginst1504 (i_6472, i_6040);
  and ginst1505 (i_6473, i_4524, i_5315, i_6031);
  and ginst1506 (i_6474, i_5150, i_6025, i_6034);
  and ginst1507 (i_6475, i_4532, i_5324, i_6037);
  and ginst1508 (i_6476, i_5157, i_6028, i_6040);
  nand ginst1509 (i_6477, i_5385, i_6234);
  nand ginst1510 (i_6478, i_132, i_6045);
  or ginst1511 (i_6482, i_4280, i_6083, i_6084, i_6085);
  nor ginst1512 (i_6486, i_4280, i_6086, i_6087);
  or ginst1513 (i_6490, i_4284, i_6088, i_6089);
  nor ginst1514 (i_6494, i_4284, i_6090);
  or ginst1515 (i_6500, i_4298, i_6098, i_6099, i_6100, i_6101);
  or ginst1516 (i_6504, i_4301, i_6102, i_6103, i_6104);
  or ginst1517 (i_6508, i_4305, i_6105, i_6106);
  or ginst1518 (i_6512, i_4310, i_6107);
  or ginst1519 (i_6516, i_4316, i_6111, i_6112, i_6113);
  nor ginst1520 (i_6526, i_4316, i_6114, i_6115);
  or ginst1521 (i_6536, i_4336, i_6131, i_6132, i_6133);
  or ginst1522 (i_6539, i_4332, i_6124, i_6125, i_6126, i_6127);
  nor ginst1523 (i_6553, i_4336, i_6134, i_6135);
  nor ginst1524 (i_6556, i_4332, i_6128, i_6129, i_6130);
  or ginst1525 (i_6566, i_4375, i_5117, i_6143, i_6144);
  nor ginst1526 (i_6569, i_4375, i_5118, i_6145);
  or ginst1527 (i_6572, i_4379, i_6146, i_6147);
  nor ginst1528 (i_6575, i_4379, i_6148);
  or ginst1529 (i_6580, i_4067, i_5954, i_6156, i_6157, i_6158);
  or ginst1530 (i_6584, i_4396, i_6159, i_6160, i_6161);
  or ginst1531 (i_6587, i_4400, i_6162, i_6163);
  or ginst1532 (i_6592, i_4436, i_5132, i_6171, i_6172);
  nor ginst1533 (i_6599, i_4436, i_5133, i_6173);
  or ginst1534 (i_6606, i_4456, i_6187, i_6188, i_6189);
  or ginst1535 (i_6609, i_4080, i_6005, i_6182, i_6183, i_6184);
  nor ginst1536 (i_6619, i_4456, i_6190, i_6191);
  nor ginst1537 (i_6622, i_4080, i_6006, i_6185, i_6186);
  nand ginst1538 (i_6630, i_5739, i_6373);
  nand ginst1539 (i_6631, i_5736, i_6374);
  nand ginst1540 (i_6632, i_5745, i_6375);
  nand ginst1541 (i_6633, i_5742, i_6376);
  nand ginst1542 (i_6634, i_6066, i_6377);
  nand ginst1543 (i_6637, i_6069, i_6378);
  not ginst1544 (i_6640, i_6164);
  and ginst1545 (i_6641, i_6108, i_6117);
  and ginst1546 (i_6643, i_6140, i_6149);
  and ginst1547 (i_6646, i_6168, i_6175);
  and ginst1548 (i_6648, i_6080, i_6091);
  nand ginst1549 (i_6650, i_2637, i_6238);
  not ginst1550 (i_6651, i_6238);
  not ginst1551 (i_6653, i_6241);
  not ginst1552 (i_6655, i_6244);
  not ginst1553 (i_6657, i_6247);
  not ginst1554 (i_6659, i_6250);
  nand ginst1555 (i_6660, i_5087, i_6253);
  not ginst1556 (i_6661, i_6253);
  nand ginst1557 (i_6662, i_5469, i_6256);
  not ginst1558 (i_6663, i_6256);
  and ginst1559 (i_6664, i_4, i_6091);
  not ginst1560 (i_6666, i_6259);
  not ginst1561 (i_6668, i_6262);
  not ginst1562 (i_6670, i_6265);
  not ginst1563 (i_6672, i_6268);
  not ginst1564 (i_6675, i_6117);
  not ginst1565 (i_6680, i_6280);
  not ginst1566 (i_6681, i_6292);
  not ginst1567 (i_6682, i_6307);
  not ginst1568 (i_6683, i_6310);
  nand ginst1569 (i_6689, i_5120, i_6325);
  not ginst1570 (i_6690, i_6325);
  nand ginst1571 (i_6691, i_5622, i_6328);
  not ginst1572 (i_6692, i_6328);
  and ginst1573 (i_6693, i_54, i_6149);
  not ginst1574 (i_6695, i_6331);
  not ginst1575 (i_6698, i_6335);
  nand ginst1576 (i_6699, i_5956, i_6338);
  not ginst1577 (i_6700, i_6338);
  not ginst1578 (i_6703, i_6175);
  not ginst1579 (i_6708, i_6209);
  not ginst1580 (i_6709, i_6212);
  not ginst1581 (i_6710, i_6215);
  not ginst1582 (i_6711, i_6218);
  and ginst1583 (i_6712, i_5692, i_5696, i_6209);
  and ginst1584 (i_6713, i_6197, i_6200, i_6212);
  and ginst1585 (i_6714, i_5703, i_5707, i_6215);
  and ginst1586 (i_6715, i_6203, i_6206, i_6218);
  not ginst1587 (i_6716, i_6466);
  and ginst1588 (i_6718, i_1777, i_3130, i_6164);
  and ginst1589 (i_6719, i_5150, i_5315, i_6469);
  and ginst1590 (i_6720, i_4524, i_6025, i_6470);
  and ginst1591 (i_6721, i_5157, i_5324, i_6471);
  and ginst1592 (i_6722, i_4532, i_6028, i_6472);
  nand ginst1593 (i_6724, i_6235, i_6477);
  not ginst1594 (i_6739, i_6271);
  not ginst1595 (i_6740, i_6274);
  not ginst1596 (i_6741, i_6277);
  not ginst1597 (i_6744, i_6283);
  not ginst1598 (i_6745, i_6286);
  not ginst1599 (i_6746, i_6289);
  not ginst1600 (i_6751, i_6295);
  not ginst1601 (i_6752, i_6298);
  not ginst1602 (i_6753, i_6301);
  not ginst1603 (i_6754, i_6304);
  not ginst1604 (i_6755, i_6322);
  not ginst1605 (i_6760, i_6313);
  not ginst1606 (i_6761, i_6316);
  not ginst1607 (i_6762, i_6319);
  not ginst1608 (i_6772, i_6341);
  not ginst1609 (i_6773, i_6344);
  not ginst1610 (i_6776, i_6347);
  not ginst1611 (i_6777, i_6350);
  not ginst1612 (i_6782, i_6353);
  not ginst1613 (i_6783, i_6356);
  not ginst1614 (i_6784, i_6359);
  not ginst1615 (i_6785, i_6370);
  not ginst1616 (i_6790, i_6364);
  not ginst1617 (i_6791, i_6367);
  nand ginst1618 (i_6792, i_6630, i_6631);
  nand ginst1619 (i_6795, i_6632, i_6633);
  and ginst1620 (i_6801, i_6108, i_6415);
  and ginst1621 (i_6802, i_6140, i_6427);
  and ginst1622 (i_6803, i_6080, i_6397);
  and ginst1623 (i_6804, i_6168, i_6441);
  not ginst1624 (i_6805, i_6466);
  nand ginst1625 (i_6806, i_1851, i_6651);
  not ginst1626 (i_6807, i_6482);
  nand ginst1627 (i_6808, i_6482, i_6653);
  not ginst1628 (i_6809, i_6486);
  nand ginst1629 (i_6810, i_6486, i_6655);
  not ginst1630 (i_6811, i_6490);
  nand ginst1631 (i_6812, i_6490, i_6657);
  not ginst1632 (i_6813, i_6494);
  nand ginst1633 (i_6814, i_6494, i_6659);
  nand ginst1634 (i_6815, i_4575, i_6661);
  nand ginst1635 (i_6816, i_5169, i_6663);
  or ginst1636 (i_6817, i_6397, i_6664);
  not ginst1637 (i_6823, i_6500);
  nand ginst1638 (i_6824, i_6500, i_6666);
  not ginst1639 (i_6825, i_6504);
  nand ginst1640 (i_6826, i_6504, i_6668);
  not ginst1641 (i_6827, i_6508);
  nand ginst1642 (i_6828, i_6508, i_6670);
  not ginst1643 (i_6829, i_6512);
  nand ginst1644 (i_6830, i_6512, i_6672);
  not ginst1645 (i_6831, i_6415);
  not ginst1646 (i_6834, i_6566);
  nand ginst1647 (i_6835, i_5618, i_6566);
  not ginst1648 (i_6836, i_6569);
  nand ginst1649 (i_6837, i_5619, i_6569);
  not ginst1650 (i_6838, i_6572);
  nand ginst1651 (i_6839, i_5620, i_6572);
  not ginst1652 (i_6840, i_6575);
  nand ginst1653 (i_6841, i_5621, i_6575);
  nand ginst1654 (i_6842, i_4627, i_6690);
  nand ginst1655 (i_6843, i_5195, i_6692);
  or ginst1656 (i_6844, i_6427, i_6693);
  not ginst1657 (i_6850, i_6580);
  nand ginst1658 (i_6851, i_6580, i_6695);
  not ginst1659 (i_6852, i_6584);
  nand ginst1660 (i_6853, i_6434, i_6584);
  not ginst1661 (i_6854, i_6587);
  nand ginst1662 (i_6855, i_6587, i_6698);
  nand ginst1663 (i_6856, i_5346, i_6700);
  not ginst1664 (i_6857, i_6441);
  and ginst1665 (i_6860, i_5696, i_6197, i_6708);
  and ginst1666 (i_6861, i_5692, i_6200, i_6709);
  and ginst1667 (i_6862, i_5707, i_6203, i_6710);
  and ginst1668 (i_6863, i_5703, i_6206, i_6711);
  or ginst1669 (i_6866, i_3785, i_4197, i_6718);
  nor ginst1670 (i_6872, i_6473, i_6719);
  nor ginst1671 (i_6873, i_6474, i_6720);
  nor ginst1672 (i_6874, i_6475, i_6721);
  nor ginst1673 (i_6875, i_6476, i_6722);
  not ginst1674 (i_6876, i_6637);
  not ginst1675 (i_6877, i_6724);
  and ginst1676 (i_6879, i_6045, i_6478);
  and ginst1677 (i_6880, i_132, i_6478);
  or ginst1678 (i_6881, i_6137, i_6411);
  not ginst1679 (i_6884, i_6516);
  not ginst1680 (i_6885, i_6411);
  not ginst1681 (i_6888, i_6526);
  not ginst1682 (i_6889, i_6536);
  nand ginst1683 (i_6890, i_5176, i_6536);
  or ginst1684 (i_6891, i_6138, i_6419);
  not ginst1685 (i_6894, i_6539);
  not ginst1686 (i_6895, i_6553);
  nand ginst1687 (i_6896, i_5728, i_6553);
  not ginst1688 (i_6897, i_6419);
  not ginst1689 (i_6900, i_6556);
  or ginst1690 (i_6901, i_6193, i_6437);
  not ginst1691 (i_6904, i_6592);
  not ginst1692 (i_6905, i_6437);
  not ginst1693 (i_6908, i_6599);
  or ginst1694 (i_6909, i_6194, i_6445);
  not ginst1695 (i_6912, i_6606);
  not ginst1696 (i_6913, i_6609);
  not ginst1697 (i_6914, i_6619);
  nand ginst1698 (i_6915, i_5734, i_6619);
  not ginst1699 (i_6916, i_6445);
  not ginst1700 (i_6919, i_6622);
  not ginst1701 (i_6922, i_6634);
  nand ginst1702 (i_6923, i_6067, i_6634);
  or ginst1703 (i_6924, i_6382, i_6801);
  or ginst1704 (i_6925, i_6386, i_6802);
  or ginst1705 (i_6926, i_6388, i_6803);
  or ginst1706 (i_6927, i_6392, i_6804);
  not ginst1707 (i_6930, i_6724);
  nand ginst1708 (i_6932, i_6650, i_6806);
  nand ginst1709 (i_6935, i_6241, i_6807);
  nand ginst1710 (i_6936, i_6244, i_6809);
  nand ginst1711 (i_6937, i_6247, i_6811);
  nand ginst1712 (i_6938, i_6250, i_6813);
  nand ginst1713 (i_6939, i_6660, i_6815);
  nand ginst1714 (i_6940, i_6662, i_6816);
  nand ginst1715 (i_6946, i_6259, i_6823);
  nand ginst1716 (i_6947, i_6262, i_6825);
  nand ginst1717 (i_6948, i_6265, i_6827);
  nand ginst1718 (i_6949, i_6268, i_6829);
  nand ginst1719 (i_6953, i_5183, i_6834);
  nand ginst1720 (i_6954, i_5186, i_6836);
  nand ginst1721 (i_6955, i_5189, i_6838);
  nand ginst1722 (i_6956, i_5192, i_6840);
  nand ginst1723 (i_6957, i_6689, i_6842);
  nand ginst1724 (i_6958, i_6691, i_6843);
  nand ginst1725 (i_6964, i_6331, i_6850);
  nand ginst1726 (i_6965, i_6048, i_6852);
  nand ginst1727 (i_6966, i_6335, i_6854);
  nand ginst1728 (i_6967, i_6699, i_6856);
  nor ginst1729 (i_6973, i_6712, i_6860);
  nor ginst1730 (i_6974, i_6713, i_6861);
  nor ginst1731 (i_6975, i_6714, i_6862);
  nor ginst1732 (i_6976, i_6715, i_6863);
  not ginst1733 (i_6977, i_6792);
  not ginst1734 (i_6978, i_6795);
  or ginst1735 (i_6979, i_6879, i_6880);
  nand ginst1736 (i_6987, i_4608, i_6889);
  nand ginst1737 (i_6990, i_5177, i_6895);
  nand ginst1738 (i_6999, i_5217, i_6914);
  nand ginst1739 (i_7002, i_5377, i_6922);
  nand ginst1740 (i_7003, i_6872, i_6873);
  nand ginst1741 (i_7006, i_6874, i_6875);
  and ginst1742 (i_7011, i_2681, i_2692, i_6866);
  and ginst1743 (i_7012, i_2756, i_2767, i_6866);
  and ginst1744 (i_7013, i_2779, i_2790, i_6866);
  not ginst1745 (i_7015, i_6866);
  and ginst1746 (i_7016, i_2801, i_2812, i_6866);
  nand ginst1747 (i_7018, i_6808, i_6935);
  nand ginst1748 (i_7019, i_6810, i_6936);
  nand ginst1749 (i_7020, i_6812, i_6937);
  nand ginst1750 (i_7021, i_6814, i_6938);
  not ginst1751 (i_7022, i_6939);
  not ginst1752 (i_7023, i_6817);
  nand ginst1753 (i_7028, i_6824, i_6946);
  nand ginst1754 (i_7031, i_6826, i_6947);
  nand ginst1755 (i_7034, i_6828, i_6948);
  nand ginst1756 (i_7037, i_6830, i_6949);
  and ginst1757 (i_7040, i_6079, i_6817);
  and ginst1758 (i_7041, i_6675, i_6831);
  nand ginst1759 (i_7044, i_6835, i_6953);
  nand ginst1760 (i_7045, i_6837, i_6954);
  nand ginst1761 (i_7046, i_6839, i_6955);
  nand ginst1762 (i_7047, i_6841, i_6956);
  not ginst1763 (i_7048, i_6957);
  not ginst1764 (i_7049, i_6844);
  nand ginst1765 (i_7054, i_6851, i_6964);
  nand ginst1766 (i_7057, i_6853, i_6965);
  nand ginst1767 (i_7060, i_6855, i_6966);
  and ginst1768 (i_7064, i_6139, i_6844);
  and ginst1769 (i_7065, i_6703, i_6857);
  not ginst1770 (i_7072, i_6881);
  nand ginst1771 (i_7073, i_5172, i_6881);
  not ginst1772 (i_7074, i_6885);
  nand ginst1773 (i_7075, i_5727, i_6885);
  nand ginst1774 (i_7076, i_6890, i_6987);
  not ginst1775 (i_7079, i_6891);
  nand ginst1776 (i_7080, i_6896, i_6990);
  not ginst1777 (i_7083, i_6897);
  not ginst1778 (i_7084, i_6901);
  nand ginst1779 (i_7085, i_5198, i_6901);
  not ginst1780 (i_7086, i_6905);
  nand ginst1781 (i_7087, i_5731, i_6905);
  not ginst1782 (i_7088, i_6909);
  nand ginst1783 (i_7089, i_6909, i_6912);
  not ginst1784 (i_709, i_141);
  nand ginst1785 (i_7090, i_6915, i_6999);
  not ginst1786 (i_7093, i_6916);
  nand ginst1787 (i_7094, i_6973, i_6974);
  nand ginst1788 (i_7097, i_6975, i_6976);
  nand ginst1789 (i_7101, i_6923, i_7002);
  not ginst1790 (i_7105, i_6932);
  not ginst1791 (i_7110, i_6967);
  and ginst1792 (i_7114, i_603, i_1755, i_6979);
  not ginst1793 (i_7115, i_7019);
  not ginst1794 (i_7116, i_7021);
  and ginst1795 (i_7125, i_6817, i_7018);
  and ginst1796 (i_7126, i_6817, i_7020);
  and ginst1797 (i_7127, i_6817, i_7022);
  not ginst1798 (i_7130, i_7045);
  not ginst1799 (i_7131, i_7047);
  and ginst1800 (i_7139, i_6844, i_7044);
  and ginst1801 (i_7140, i_6844, i_7046);
  and ginst1802 (i_7141, i_6844, i_7048);
  and ginst1803 (i_7146, i_1761, i_3108, i_6932);
  and ginst1804 (i_7147, i_1777, i_3130, i_6967);
  not ginst1805 (i_7149, i_7003);
  not ginst1806 (i_7150, i_7006);
  nand ginst1807 (i_7151, i_6876, i_7006);
  nand ginst1808 (i_7152, i_4605, i_7072);
  nand ginst1809 (i_7153, i_5173, i_7074);
  nand ginst1810 (i_7158, i_4646, i_7084);
  nand ginst1811 (i_7159, i_5205, i_7086);
  nand ginst1812 (i_7160, i_6606, i_7088);
  not ginst1813 (i_7166, i_7037);
  not ginst1814 (i_7167, i_7034);
  not ginst1815 (i_7168, i_7031);
  not ginst1816 (i_7169, i_7028);
  not ginst1817 (i_7170, i_7060);
  not ginst1818 (i_7171, i_7057);
  not ginst1819 (i_7172, i_7054);
  and ginst1820 (i_7173, i_7023, i_7115);
  and ginst1821 (i_7174, i_7023, i_7116);
  and ginst1822 (i_7175, i_6940, i_7023);
  and ginst1823 (i_7176, i_5418, i_7023);
  not ginst1824 (i_7177, i_7041);
  and ginst1825 (i_7178, i_7049, i_7130);
  and ginst1826 (i_7179, i_7049, i_7131);
  and ginst1827 (i_7180, i_6958, i_7049);
  and ginst1828 (i_7181, i_5573, i_7049);
  not ginst1829 (i_7182, i_7065);
  not ginst1830 (i_7183, i_7094);
  nand ginst1831 (i_7184, i_6977, i_7094);
  not ginst1832 (i_7185, i_7097);
  nand ginst1833 (i_7186, i_6978, i_7097);
  and ginst1834 (i_7187, i_1761, i_3108, i_7037);
  and ginst1835 (i_7188, i_1761, i_3108, i_7034);
  and ginst1836 (i_7189, i_1761, i_3108, i_7031);
  or ginst1837 (i_7190, i_3781, i_4956, i_7146);
  and ginst1838 (i_7196, i_1777, i_3130, i_7060);
  and ginst1839 (i_7197, i_1777, i_3130, i_7057);
  or ginst1840 (i_7198, i_3786, i_4960, i_7147);
  nand ginst1841 (i_7204, i_7101, i_7149);
  not ginst1842 (i_7205, i_7101);
  nand ginst1843 (i_7206, i_6637, i_7150);
  and ginst1844 (i_7207, i_1793, i_3158, i_7028);
  and ginst1845 (i_7208, i_1807, i_3180, i_7054);
  nand ginst1846 (i_7209, i_7073, i_7152);
  nand ginst1847 (i_7212, i_7075, i_7153);
  not ginst1848 (i_7215, i_7076);
  nand ginst1849 (i_7216, i_7076, i_7079);
  not ginst1850 (i_7217, i_7080);
  nand ginst1851 (i_7218, i_7080, i_7083);
  nand ginst1852 (i_7219, i_7085, i_7158);
  nand ginst1853 (i_7222, i_7087, i_7159);
  nand ginst1854 (i_7225, i_7089, i_7160);
  not ginst1855 (i_7228, i_7090);
  nand ginst1856 (i_7229, i_7090, i_7093);
  or ginst1857 (i_7236, i_7125, i_7173);
  or ginst1858 (i_7239, i_7126, i_7174);
  or ginst1859 (i_7242, i_7127, i_7175);
  or ginst1860 (i_7245, i_7040, i_7176);
  or ginst1861 (i_7250, i_7139, i_7178);
  or ginst1862 (i_7257, i_7140, i_7179);
  or ginst1863 (i_7260, i_7141, i_7180);
  or ginst1864 (i_7263, i_7064, i_7181);
  nand ginst1865 (i_7268, i_6792, i_7183);
  nand ginst1866 (i_7269, i_6795, i_7185);
  or ginst1867 (i_7270, i_3782, i_4957, i_7187);
  or ginst1868 (i_7276, i_3783, i_4958, i_7188);
  or ginst1869 (i_7282, i_3784, i_4959, i_7189);
  or ginst1870 (i_7288, i_3787, i_4961, i_7196);
  or ginst1871 (i_7294, i_3788, i_3998, i_7197);
  nand ginst1872 (i_7300, i_7003, i_7205);
  nand ginst1873 (i_7301, i_7151, i_7206);
  or ginst1874 (i_7304, i_3800, i_4980, i_7207);
  or ginst1875 (i_7310, i_3805, i_4984, i_7208);
  nand ginst1876 (i_7320, i_6891, i_7215);
  nand ginst1877 (i_7321, i_6897, i_7217);
  nand ginst1878 (i_7328, i_6916, i_7228);
  and ginst1879 (i_7338, i_1185, i_2692, i_7190);
  and ginst1880 (i_7339, i_2681, i_2692, i_7198);
  and ginst1881 (i_7340, i_1247, i_2767, i_7190);
  and ginst1882 (i_7341, i_2756, i_2767, i_7198);
  and ginst1883 (i_7342, i_1327, i_2790, i_7190);
  and ginst1884 (i_7349, i_2779, i_2790, i_7198);
  and ginst1885 (i_7357, i_2801, i_2812, i_7198);
  not ginst1886 (i_7363, i_7198);
  and ginst1887 (i_7364, i_1351, i_2812, i_7190);
  not ginst1888 (i_7365, i_7190);
  nand ginst1889 (i_7394, i_7184, i_7268);
  nand ginst1890 (i_7397, i_7186, i_7269);
  nand ginst1891 (i_7402, i_7204, i_7300);
  not ginst1892 (i_7405, i_7209);
  nand ginst1893 (i_7406, i_6884, i_7209);
  not ginst1894 (i_7407, i_7212);
  nand ginst1895 (i_7408, i_6888, i_7212);
  nand ginst1896 (i_7409, i_7216, i_7320);
  nand ginst1897 (i_7412, i_7218, i_7321);
  not ginst1898 (i_7415, i_7219);
  nand ginst1899 (i_7416, i_6904, i_7219);
  not ginst1900 (i_7417, i_7222);
  nand ginst1901 (i_7418, i_6908, i_7222);
  not ginst1902 (i_7419, i_7225);
  nand ginst1903 (i_7420, i_6913, i_7225);
  nand ginst1904 (i_7421, i_7229, i_7328);
  not ginst1905 (i_7424, i_7245);
  not ginst1906 (i_7425, i_7242);
  not ginst1907 (i_7426, i_7239);
  not ginst1908 (i_7427, i_7236);
  not ginst1909 (i_7428, i_7263);
  not ginst1910 (i_7429, i_7260);
  not ginst1911 (i_7430, i_7257);
  not ginst1912 (i_7431, i_7250);
  not ginst1913 (i_7432, i_7250);
  and ginst1914 (i_7433, i_2653, i_2664, i_7310);
  and ginst1915 (i_7434, i_1161, i_2664, i_7304);
  or ginst1916 (i_7435, i_2591, i_3621, i_7011, i_7338);
  and ginst1917 (i_7436, i_1185, i_2692, i_7270);
  and ginst1918 (i_7437, i_2681, i_2692, i_7288);
  and ginst1919 (i_7438, i_1185, i_2692, i_7276);
  and ginst1920 (i_7439, i_2681, i_2692, i_7294);
  and ginst1921 (i_7440, i_1185, i_2692, i_7282);
  and ginst1922 (i_7441, i_2728, i_2739, i_7310);
  and ginst1923 (i_7442, i_1223, i_2739, i_7304);
  or ginst1924 (i_7443, i_2600, i_3632, i_7012, i_7340);
  and ginst1925 (i_7444, i_1247, i_2767, i_7270);
  and ginst1926 (i_7445, i_2756, i_2767, i_7288);
  and ginst1927 (i_7446, i_1247, i_2767, i_7276);
  and ginst1928 (i_7447, i_2756, i_2767, i_7294);
  and ginst1929 (i_7448, i_1247, i_2767, i_7282);
  or ginst1930 (i_7449, i_2605, i_3641, i_7013, i_7342);
  and ginst1931 (i_7450, i_3041, i_3052, i_7310);
  and ginst1932 (i_7451, i_1697, i_3052, i_7304);
  and ginst1933 (i_7452, i_2779, i_2790, i_7294);
  and ginst1934 (i_7453, i_1327, i_2790, i_7282);
  and ginst1935 (i_7454, i_2779, i_2790, i_7288);
  and ginst1936 (i_7455, i_1327, i_2790, i_7276);
  and ginst1937 (i_7456, i_1327, i_2790, i_7270);
  and ginst1938 (i_7457, i_3075, i_3086, i_7310);
  and ginst1939 (i_7458, i_1731, i_3086, i_7304);
  and ginst1940 (i_7459, i_2801, i_2812, i_7294);
  and ginst1941 (i_7460, i_1351, i_2812, i_7282);
  and ginst1942 (i_7461, i_2801, i_2812, i_7288);
  and ginst1943 (i_7462, i_1351, i_2812, i_7276);
  and ginst1944 (i_7463, i_1351, i_2812, i_7270);
  and ginst1945 (i_7464, i_599, i_603, i_7250);
  not ginst1946 (i_7465, i_7310);
  not ginst1947 (i_7466, i_7294);
  not ginst1948 (i_7467, i_7288);
  not ginst1949 (i_7468, i_7301);
  or ginst1950 (i_7469, i_2626, i_3660, i_7016, i_7364);
  not ginst1951 (i_7470, i_7304);
  not ginst1952 (i_7471, i_7282);
  not ginst1953 (i_7472, i_7276);
  not ginst1954 (i_7473, i_7270);
  not ginst1955 (i_7474, i_7394);
  not ginst1956 (i_7476, i_7397);
  and ginst1957 (i_7479, i_3068, i_7301);
  and ginst1958 (i_7481, i_1793, i_3158, i_7245);
  and ginst1959 (i_7482, i_1793, i_3158, i_7242);
  and ginst1960 (i_7483, i_1793, i_3158, i_7239);
  and ginst1961 (i_7484, i_1793, i_3158, i_7236);
  and ginst1962 (i_7485, i_1807, i_3180, i_7263);
  and ginst1963 (i_7486, i_1807, i_3180, i_7260);
  and ginst1964 (i_7487, i_1807, i_3180, i_7257);
  and ginst1965 (i_7488, i_1807, i_3180, i_7250);
  nand ginst1966 (i_7489, i_6979, i_7250);
  nand ginst1967 (i_7492, i_6516, i_7405);
  nand ginst1968 (i_7493, i_6526, i_7407);
  nand ginst1969 (i_7498, i_6592, i_7415);
  nand ginst1970 (i_7499, i_6599, i_7417);
  nand ginst1971 (i_7500, i_6609, i_7419);
  and ginst1972 (i_7503, i_7105, i_7166, i_7167, i_7168, i_7169, i_7424, i_7425, i_7426, i_7427);
  and ginst1973 (i_7504, i_6640, i_7110, i_7170, i_7171, i_7172, i_7428, i_7429, i_7430, i_7431);
  or ginst1974 (i_7505, i_2585, i_3616, i_7433, i_7434);
  and ginst1975 (i_7506, i_2675, i_7435);
  or ginst1976 (i_7507, i_2592, i_3622, i_7339, i_7436);
  or ginst1977 (i_7508, i_2593, i_3623, i_7437, i_7438);
  or ginst1978 (i_7509, i_2594, i_3624, i_7439, i_7440);
  or ginst1979 (i_7510, i_2595, i_3627, i_7441, i_7442);
  and ginst1980 (i_7511, i_2750, i_7443);
  or ginst1981 (i_7512, i_2601, i_3633, i_7341, i_7444);
  or ginst1982 (i_7513, i_2602, i_3634, i_7445, i_7446);
  or ginst1983 (i_7514, i_2603, i_3635, i_7447, i_7448);
  or ginst1984 (i_7515, i_2610, i_3646, i_7450, i_7451);
  or ginst1985 (i_7516, i_2611, i_3647, i_7452, i_7453);
  or ginst1986 (i_7517, i_2612, i_3648, i_7454, i_7455);
  or ginst1987 (i_7518, i_2613, i_3649, i_7349, i_7456);
  or ginst1988 (i_7519, i_2618, i_3654, i_7457, i_7458);
  or ginst1989 (i_7520, i_2619, i_3655, i_7459, i_7460);
  or ginst1990 (i_7521, i_2620, i_3656, i_7461, i_7462);
  or ginst1991 (i_7522, i_2621, i_3657, i_7357, i_7463);
  or ginst1992 (i_7525, i_2624, i_4741, i_7114, i_7464);
  and ginst1993 (i_7526, i_3119, i_3130, i_7468);
  not ginst1994 (i_7527, i_7394);
  not ginst1995 (i_7528, i_7397);
  not ginst1996 (i_7529, i_7402);
  and ginst1997 (i_7530, i_3068, i_7402);
  or ginst1998 (i_7531, i_3801, i_4981, i_7481);
  or ginst1999 (i_7537, i_3802, i_4982, i_7482);
  or ginst2000 (i_7543, i_3803, i_4983, i_7483);
  or ginst2001 (i_7549, i_3804, i_5165, i_7484);
  or ginst2002 (i_7555, i_3806, i_4985, i_7485);
  or ginst2003 (i_7561, i_3807, i_4986, i_7486);
  or ginst2004 (i_7567, i_3808, i_4547, i_7487);
  or ginst2005 (i_7573, i_3809, i_4987, i_7488);
  nand ginst2006 (i_7579, i_7406, i_7492);
  nand ginst2007 (i_7582, i_7408, i_7493);
  not ginst2008 (i_7585, i_7409);
  nand ginst2009 (i_7586, i_6894, i_7409);
  not ginst2010 (i_7587, i_7412);
  nand ginst2011 (i_7588, i_6900, i_7412);
  nand ginst2012 (i_7589, i_7416, i_7498);
  nand ginst2013 (i_7592, i_7418, i_7499);
  nand ginst2014 (i_7595, i_7420, i_7500);
  not ginst2015 (i_7598, i_7421);
  nand ginst2016 (i_7599, i_6919, i_7421);
  and ginst2017 (i_7600, i_2647, i_7505);
  and ginst2018 (i_7601, i_2675, i_7507);
  and ginst2019 (i_7602, i_2675, i_7508);
  and ginst2020 (i_7603, i_2675, i_7509);
  and ginst2021 (i_7604, i_2722, i_7510);
  and ginst2022 (i_7605, i_2750, i_7512);
  and ginst2023 (i_7606, i_2750, i_7513);
  and ginst2024 (i_7607, i_2750, i_7514);
  and ginst2025 (i_7624, i_6979, i_7489);
  and ginst2026 (i_7625, i_7250, i_7489);
  and ginst2027 (i_7626, i_1149, i_7525);
  and ginst2028 (i_7631, i_562, i_6805, i_6930, i_7527, i_7528);
  and ginst2029 (i_7636, i_3097, i_3108, i_7529);
  nand ginst2030 (i_7657, i_6539, i_7585);
  nand ginst2031 (i_7658, i_6556, i_7587);
  nand ginst2032 (i_7665, i_6622, i_7598);
  and ginst2033 (i_7666, i_2653, i_2664, i_7555);
  and ginst2034 (i_7667, i_1161, i_2664, i_7531);
  and ginst2035 (i_7668, i_2653, i_2664, i_7561);
  and ginst2036 (i_7669, i_1161, i_2664, i_7537);
  and ginst2037 (i_7670, i_2653, i_2664, i_7567);
  and ginst2038 (i_7671, i_1161, i_2664, i_7543);
  and ginst2039 (i_7672, i_2653, i_2664, i_7573);
  and ginst2040 (i_7673, i_1161, i_2664, i_7549);
  and ginst2041 (i_7674, i_2728, i_2739, i_7555);
  and ginst2042 (i_7675, i_1223, i_2739, i_7531);
  and ginst2043 (i_7676, i_2728, i_2739, i_7561);
  and ginst2044 (i_7677, i_1223, i_2739, i_7537);
  and ginst2045 (i_7678, i_2728, i_2739, i_7567);
  and ginst2046 (i_7679, i_1223, i_2739, i_7543);
  and ginst2047 (i_7680, i_2728, i_2739, i_7573);
  and ginst2048 (i_7681, i_1223, i_2739, i_7549);
  and ginst2049 (i_7682, i_3075, i_3086, i_7573);
  and ginst2050 (i_7683, i_1731, i_3086, i_7549);
  and ginst2051 (i_7684, i_3041, i_3052, i_7573);
  and ginst2052 (i_7685, i_1697, i_3052, i_7549);
  and ginst2053 (i_7686, i_3041, i_3052, i_7567);
  and ginst2054 (i_7687, i_1697, i_3052, i_7543);
  and ginst2055 (i_7688, i_3041, i_3052, i_7561);
  and ginst2056 (i_7689, i_1697, i_3052, i_7537);
  and ginst2057 (i_7690, i_3041, i_3052, i_7555);
  and ginst2058 (i_7691, i_1697, i_3052, i_7531);
  and ginst2059 (i_7692, i_3075, i_3086, i_7567);
  and ginst2060 (i_7693, i_1731, i_3086, i_7543);
  and ginst2061 (i_7694, i_3075, i_3086, i_7561);
  and ginst2062 (i_7695, i_1731, i_3086, i_7537);
  and ginst2063 (i_7696, i_3075, i_3086, i_7555);
  and ginst2064 (i_7697, i_1731, i_3086, i_7531);
  or ginst2065 (i_7698, i_7624, i_7625);
  not ginst2066 (i_7699, i_7573);
  not ginst2067 (i_7700, i_7567);
  xor ginst2068 (i_7701, i_7701_in, flip_signal);
  not ginst2069 (i_7701_in, i_7561);
  not ginst2070 (i_7702, i_7555);
  and ginst2071 (i_7703, i_245, i_1156, i_7631);
  not ginst2072 (i_7704, i_7549);
  not ginst2073 (i_7705, i_7543);
  not ginst2074 (i_7706, i_7537);
  not ginst2075 (i_7707, i_7531);
  not ginst2076 (i_7708, i_7579);
  nand ginst2077 (i_7709, i_6739, i_7579);
  not ginst2078 (i_7710, i_7582);
  nand ginst2079 (i_7711, i_6744, i_7582);
  nand ginst2080 (i_7712, i_7586, i_7657);
  nand ginst2081 (i_7715, i_7588, i_7658);
  not ginst2082 (i_7718, i_7589);
  nand ginst2083 (i_7719, i_6772, i_7589);
  not ginst2084 (i_7720, i_7592);
  nand ginst2085 (i_7721, i_6776, i_7592);
  not ginst2086 (i_7722, i_7595);
  nand ginst2087 (i_7723, i_5733, i_7595);
  nand ginst2088 (i_7724, i_7599, i_7665);
  or ginst2089 (i_7727, i_2586, i_3617, i_7666, i_7667);
  or ginst2090 (i_7728, i_2587, i_3618, i_7668, i_7669);
  or ginst2091 (i_7729, i_2588, i_3619, i_7670, i_7671);
  or ginst2092 (i_7730, i_2589, i_3620, i_7672, i_7673);
  or ginst2093 (i_7731, i_2596, i_3628, i_7674, i_7675);
  or ginst2094 (i_7732, i_2597, i_3629, i_7676, i_7677);
  or ginst2095 (i_7733, i_2598, i_3630, i_7678, i_7679);
  or ginst2096 (i_7734, i_2599, i_3631, i_7680, i_7681);
  or ginst2097 (i_7735, i_2604, i_3638, i_7682, i_7683);
  or ginst2098 (i_7736, i_2606, i_3642, i_7684, i_7685);
  or ginst2099 (i_7737, i_2607, i_3643, i_7686, i_7687);
  or ginst2100 (i_7738, i_2608, i_3644, i_7688, i_7689);
  or ginst2101 (i_7739, i_2609, i_3645, i_7690, i_7691);
  or ginst2102 (i_7740, i_2615, i_3651, i_7692, i_7693);
  or ginst2103 (i_7741, i_2616, i_3652, i_7694, i_7695);
  or ginst2104 (i_7742, i_2617, i_3653, i_7696, i_7697);
  nand ginst2105 (i_7743, i_6271, i_7708);
  nand ginst2106 (i_7744, i_6283, i_7710);
  nand ginst2107 (i_7749, i_6341, i_7718);
  nand ginst2108 (i_7750, i_6347, i_7720);
  nand ginst2109 (i_7751, i_5214, i_7722);
  and ginst2110 (i_7754, i_2647, i_7727);
  and ginst2111 (i_7755, i_2647, i_7728);
  and ginst2112 (i_7756, i_2647, i_7729);
  and ginst2113 (i_7757, i_2647, i_7730);
  and ginst2114 (i_7758, i_2722, i_7731);
  and ginst2115 (i_7759, i_2722, i_7732);
  and ginst2116 (i_7760, i_2722, i_7733);
  and ginst2117 (i_7761, i_2722, i_7734);
  nand ginst2118 (i_7762, i_7709, i_7743);
  nand ginst2119 (i_7765, i_7711, i_7744);
  not ginst2120 (i_7768, i_7712);
  nand ginst2121 (i_7769, i_6751, i_7712);
  not ginst2122 (i_7770, i_7715);
  nand ginst2123 (i_7771, i_6760, i_7715);
  nand ginst2124 (i_7772, i_7719, i_7749);
  nand ginst2125 (i_7775, i_7721, i_7750);
  nand ginst2126 (i_7778, i_7723, i_7751);
  not ginst2127 (i_7781, i_7724);
  nand ginst2128 (i_7782, i_5735, i_7724);
  nand ginst2129 (i_7787, i_6295, i_7768);
  nand ginst2130 (i_7788, i_6313, i_7770);
  nand ginst2131 (i_7795, i_5220, i_7781);
  not ginst2132 (i_7796, i_7762);
  nand ginst2133 (i_7797, i_6740, i_7762);
  not ginst2134 (i_7798, i_7765);
  nand ginst2135 (i_7799, i_6745, i_7765);
  nand ginst2136 (i_7800, i_7769, i_7787);
  nand ginst2137 (i_7803, i_7771, i_7788);
  not ginst2138 (i_7806, i_7772);
  nand ginst2139 (i_7807, i_6773, i_7772);
  not ginst2140 (i_7808, i_7775);
  nand ginst2141 (i_7809, i_6777, i_7775);
  not ginst2142 (i_7810, i_7778);
  nand ginst2143 (i_7811, i_6782, i_7778);
  nand ginst2144 (i_7812, i_7782, i_7795);
  nand ginst2145 (i_7815, i_6274, i_7796);
  nand ginst2146 (i_7816, i_6286, i_7798);
  nand ginst2147 (i_7821, i_6344, i_7806);
  nand ginst2148 (i_7822, i_6350, i_7808);
  nand ginst2149 (i_7823, i_6353, i_7810);
  nand ginst2150 (i_7826, i_7797, i_7815);
  nand ginst2151 (i_7829, i_7799, i_7816);
  not ginst2152 (i_7832, i_7800);
  nand ginst2153 (i_7833, i_6752, i_7800);
  not ginst2154 (i_7834, i_7803);
  nand ginst2155 (i_7835, i_6761, i_7803);
  nand ginst2156 (i_7836, i_7807, i_7821);
  nand ginst2157 (i_7839, i_7809, i_7822);
  nand ginst2158 (i_7842, i_7811, i_7823);
  not ginst2159 (i_7845, i_7812);
  nand ginst2160 (i_7846, i_6790, i_7812);
  nand ginst2161 (i_7851, i_6298, i_7832);
  nand ginst2162 (i_7852, i_6316, i_7834);
  nand ginst2163 (i_7859, i_6364, i_7845);
  not ginst2164 (i_7860, i_7826);
  nand ginst2165 (i_7861, i_6741, i_7826);
  not ginst2166 (i_7862, i_7829);
  nand ginst2167 (i_7863, i_6746, i_7829);
  nand ginst2168 (i_7864, i_7833, i_7851);
  nand ginst2169 (i_7867, i_7835, i_7852);
  not ginst2170 (i_7870, i_7836);
  nand ginst2171 (i_7871, i_5730, i_7836);
  not ginst2172 (i_7872, i_7839);
  nand ginst2173 (i_7873, i_5732, i_7839);
  not ginst2174 (i_7874, i_7842);
  nand ginst2175 (i_7875, i_6783, i_7842);
  nand ginst2176 (i_7876, i_7846, i_7859);
  nand ginst2177 (i_7879, i_6277, i_7860);
  nand ginst2178 (i_7880, i_6289, i_7862);
  nand ginst2179 (i_7885, i_5199, i_7870);
  nand ginst2180 (i_7886, i_5208, i_7872);
  nand ginst2181 (i_7887, i_6356, i_7874);
  nand ginst2182 (i_7890, i_7861, i_7879);
  nand ginst2183 (i_7893, i_7863, i_7880);
  not ginst2184 (i_7896, i_7864);
  nand ginst2185 (i_7897, i_6753, i_7864);
  not ginst2186 (i_7898, i_7867);
  nand ginst2187 (i_7899, i_6762, i_7867);
  nand ginst2188 (i_7900, i_7871, i_7885);
  nand ginst2189 (i_7903, i_7873, i_7886);
  nand ginst2190 (i_7906, i_7875, i_7887);
  not ginst2191 (i_7909, i_7876);
  nand ginst2192 (i_7910, i_6791, i_7876);
  nand ginst2193 (i_7917, i_6301, i_7896);
  nand ginst2194 (i_7918, i_6319, i_7898);
  nand ginst2195 (i_7923, i_6367, i_7909);
  not ginst2196 (i_7924, i_7890);
  nand ginst2197 (i_7925, i_6680, i_7890);
  not ginst2198 (i_7926, i_7893);
  nand ginst2199 (i_7927, i_6681, i_7893);
  not ginst2200 (i_7928, i_7900);
  nand ginst2201 (i_7929, i_5690, i_7900);
  not ginst2202 (i_7930, i_7903);
  nand ginst2203 (i_7931, i_5691, i_7903);
  nand ginst2204 (i_7932, i_7897, i_7917);
  nand ginst2205 (i_7935, i_7899, i_7918);
  not ginst2206 (i_7938, i_7906);
  nand ginst2207 (i_7939, i_6784, i_7906);
  nand ginst2208 (i_7940, i_7910, i_7923);
  nand ginst2209 (i_7943, i_6280, i_7924);
  nand ginst2210 (i_7944, i_6292, i_7926);
  nand ginst2211 (i_7945, i_5202, i_7928);
  nand ginst2212 (i_7946, i_5211, i_7930);
  nand ginst2213 (i_7951, i_6359, i_7938);
  nand ginst2214 (i_7954, i_7925, i_7943);
  nand ginst2215 (i_7957, i_7927, i_7944);
  nand ginst2216 (i_7960, i_7929, i_7945);
  nand ginst2217 (i_7963, i_7931, i_7946);
  not ginst2218 (i_7966, i_7932);
  nand ginst2219 (i_7967, i_6754, i_7932);
  not ginst2220 (i_7968, i_7935);
  nand ginst2221 (i_7969, i_6755, i_7935);
  nand ginst2222 (i_7970, i_7939, i_7951);
  not ginst2223 (i_7973, i_7940);
  nand ginst2224 (i_7974, i_6785, i_7940);
  nand ginst2225 (i_7984, i_6304, i_7966);
  nand ginst2226 (i_7985, i_6322, i_7968);
  nand ginst2227 (i_7987, i_6370, i_7973);
  and ginst2228 (i_7988, i_1157, i_6831, i_7957);
  and ginst2229 (i_7989, i_1157, i_6415, i_7954);
  and ginst2230 (i_7990, i_566, i_7041, i_7957);
  and ginst2231 (i_7991, i_566, i_7177, i_7954);
  not ginst2232 (i_7992, i_7970);
  nand ginst2233 (i_7993, i_6448, i_7970);
  and ginst2234 (i_7994, i_1219, i_6857, i_7963);
  and ginst2235 (i_7995, i_1219, i_6441, i_7960);
  and ginst2236 (i_7996, i_583, i_7065, i_7963);
  and ginst2237 (i_7997, i_583, i_7182, i_7960);
  nand ginst2238 (i_7998, i_7967, i_7984);
  nand ginst2239 (i_8001, i_7969, i_7985);
  nand ginst2240 (i_8004, i_7974, i_7987);
  nand ginst2241 (i_8009, i_6051, i_7992);
  or ginst2242 (i_8013, i_7988, i_7989, i_7990, i_7991);
  or ginst2243 (i_8017, i_7994, i_7995, i_7996, i_7997);
  not ginst2244 (i_8020, i_7998);
  nand ginst2245 (i_8021, i_6682, i_7998);
  not ginst2246 (i_8022, i_8001);
  nand ginst2247 (i_8023, i_6683, i_8001);
  nand ginst2248 (i_8025, i_7993, i_8009);
  not ginst2249 (i_8026, i_8004);
  nand ginst2250 (i_8027, i_6449, i_8004);
  nand ginst2251 (i_8031, i_6307, i_8020);
  nand ginst2252 (i_8032, i_6310, i_8022);
  not ginst2253 (i_8033, i_8013);
  nand ginst2254 (i_8034, i_6054, i_8026);
  and ginst2255 (i_8035, i_583, i_8025);
  not ginst2256 (i_8036, i_8017);
  nand ginst2257 (i_8037, i_8021, i_8031);
  nand ginst2258 (i_8038, i_8023, i_8032);
  nand ginst2259 (i_8039, i_8027, i_8034);
  not ginst2260 (i_8040, i_8038);
  and ginst2261 (i_8041, i_566, i_8037);
  not ginst2262 (i_8042, i_8039);
  and ginst2263 (i_8043, i_1157, i_8040);
  and ginst2264 (i_8044, i_1219, i_8042);
  or ginst2265 (i_8045, i_8041, i_8043);
  or ginst2266 (i_8048, i_8035, i_8044);
  nand ginst2267 (i_8055, i_8033, i_8045);
  not ginst2268 (i_8056, i_8045);
  nand ginst2269 (i_8057, i_8036, i_8048);
  not ginst2270 (i_8058, i_8048);
  nand ginst2271 (i_8059, i_8013, i_8056);
  nand ginst2272 (i_8060, i_8017, i_8058);
  nand ginst2273 (i_8061, i_8055, i_8059);
  nand ginst2274 (i_8064, i_8057, i_8060);
  and ginst2275 (i_8071, i_1777, i_3130, i_8064);
  and ginst2276 (i_8072, i_1761, i_3108, i_8061);
  not ginst2277 (i_8073, i_8061);
  not ginst2278 (i_8074, i_8064);
  or ginst2279 (i_8075, i_2625, i_3659, i_7526, i_8071);
  or ginst2280 (i_8076, i_2627, i_3661, i_7636, i_8072);
  and ginst2281 (i_8077, i_1727, i_8073);
  and ginst2282 (i_8078, i_1727, i_8074);
  or ginst2283 (i_8079, i_7530, i_8077);
  or ginst2284 (i_8082, i_7479, i_8078);
  and ginst2285 (i_8089, i_3063, i_8079);
  and ginst2286 (i_8090, i_3063, i_8082);
  and ginst2287 (i_8091, i_3063, i_8079);
  and ginst2288 (i_8092, i_3063, i_8082);
  or ginst2289 (i_8093, i_3071, i_8089);
  or ginst2290 (i_8096, i_3072, i_8090);
  or ginst2291 (i_8099, i_3073, i_8091);
  or ginst2292 (i_8102, i_3074, i_8092);
  and ginst2293 (i_8113, i_2779, i_2790, i_8102);
  and ginst2294 (i_8114, i_1327, i_2790, i_8099);
  and ginst2295 (i_8115, i_2801, i_2812, i_8102);
  and ginst2296 (i_8116, i_1351, i_2812, i_8099);
  and ginst2297 (i_8117, i_2681, i_2692, i_8096);
  and ginst2298 (i_8118, i_1185, i_2692, i_8093);
  and ginst2299 (i_8119, i_2756, i_2767, i_8096);
  and ginst2300 (i_8120, i_1247, i_2767, i_8093);
  or ginst2301 (i_8121, i_2703, i_3662, i_8117, i_8118);
  or ginst2302 (i_8122, i_2778, i_3663, i_8119, i_8120);
  or ginst2303 (i_8123, i_2614, i_3650, i_8113, i_8114);
  or ginst2304 (i_8124, i_2622, i_3658, i_8115, i_8116);
  and ginst2305 (i_8125, i_2675, i_8121);
  and ginst2306 (i_8126, i_2750, i_8122);
  not ginst2307 (i_8127, i_8125);
  not ginst2308 (i_8128, i_8126);
  not ginst2309 (i_816, i_293);

SatHard block1 (flip_signal, i_242, i_5261, i_5606, i_1887, i_2714, i_7048, i_248, i_5120, keyinput0, keyinput1, keyinput2, keyinput3, keyinput4, keyinput5, keyinput6, keyinput7, keyinput8, keyinput9, keyinput10, keyinput11, keyinput12, keyinput13, keyinput14, keyinput15);

endmodule
/*************** SatHard block ***************/
module SatHard (flip_signal, i_242, i_5261, i_5606, i_1887, i_2714, i_7048, i_248, i_5120, keyinput0, keyinput1, keyinput2, keyinput3, keyinput4, keyinput5, keyinput6, keyinput7, keyinput8, keyinput9, keyinput10, keyinput11, keyinput12, keyinput13, keyinput14, keyinput15);

  input i_242, i_5261, i_5606, i_1887, i_2714, i_7048, i_248, i_5120, keyinput0, keyinput1, keyinput2, keyinput3, keyinput4, keyinput5, keyinput6, keyinput7, keyinput8, keyinput9, keyinput10, keyinput11, keyinput12, keyinput13, keyinput14, keyinput15;
  output flip_signal;
  //SatHard key=0110110100101000
  wire [7:0] sat_res_inputs;
  assign sat_res_inputs[7:0] = {i_242, i_5261, i_5606, i_1887, i_2714, i_7048, i_248, i_5120};
  wire [15:0] keyinputs, keyvalue;
  assign keyinputs[15:0] = {keyinput0, keyinput1, keyinput2, keyinput3, keyinput4, keyinput5, keyinput6, keyinput7, keyinput8, keyinput9, keyinput10, keyinput11, keyinput12, keyinput13, keyinput14, keyinput15};
  assign keyvalue[15:0] = 16'b0110110100101000;

  wire g, g_bar;
  assign g = &(keyinputs[7:0] ^ sat_res_inputs ^ keyvalue[7:0]);
  assign g_bar = ~&(keyinputs[15:8] ^ sat_res_inputs ^ keyvalue[15:8]);
  assign flip_signal = g & g_bar;

endmodule
/*************** SatHard block ***************/
