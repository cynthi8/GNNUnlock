//key=01000001
// Main module
module c7552_AntiSAT_8_1(i_1, i_5, i_9, i_12, i_15, i_18, i_23, i_26, i_29, i_32, i_35, i_38, i_41, i_44, i_47, i_50, i_53, i_54, i_55, i_56, i_57, i_58, i_59, i_60, i_61, i_62, i_63, i_64, i_65, i_66, i_69, i_70, i_73, i_74, i_75, i_76, i_77, i_78, i_79, i_80, i_81, i_82, i_83, i_84, i_85, i_86, i_87, i_88, i_89, i_94, i_97, i_100, i_103, i_106, i_109, i_110, i_111, i_112, i_113, i_114, i_115, i_118, i_121, i_124, i_127, i_130, i_133, i_134, i_135, i_138, i_141, i_144, i_147, i_150, i_151, i_152, i_153, i_154, i_155, i_156, i_157, i_158, i_159, i_160, i_161, i_162, i_163, i_164, i_165, i_166, i_167, i_168, i_169, i_170, i_171, i_172, i_173, i_174, i_175, i_176, i_177, i_178, i_179, i_180, i_181, i_182, i_183, i_184, i_185, i_186, i_187, i_188, i_189, i_190, i_191, i_192, i_193, i_194, i_195, i_196, i_197, i_198, i_199, i_200, i_201, i_202, i_203, i_204, i_205, i_206, i_207, i_208, i_209, i_210, i_211, i_212, i_213, i_214, i_215, i_216, i_217, i_218, i_219, i_220, i_221, i_222, i_223, i_224, i_225, i_226, i_227, i_228, i_229, i_230, i_231, i_232, i_233, i_234, i_235, i_236, i_237, i_238, i_239, i_240, i_241, i_242, i_245, i_248, i_251, i_254, i_257, i_260, i_263, i_267, i_271, i_274, i_277, i_280, i_283, i_286, i_289, i_293, i_296, i_299, i_303, i_307, i_310, i_313, i_316, i_319, i_322, i_325, i_328, i_331, i_334, i_337, i_340, i_343, i_346, i_349, i_352, i_355, i_358, i_361, i_364, i_367, i_382, keyinput0, keyinput1, keyinput2, keyinput3, keyinput4, keyinput5, keyinput6, keyinput7, i_241, i_387, i_388, i_478, i_482, i_484, i_486, i_489, i_492, i_501, i_505, i_507, i_509, i_511, i_513, i_515, i_517, i_519, i_535, i_537, i_539, i_541, i_543, i_545, i_547, i_549, i_551, i_553, i_556, i_559, i_561, i_563, i_565, i_567, i_569, i_571, i_573, i_582, i_643, i_707, i_813, i_881, i_882, i_883, i_884, i_885, i_889, i_945, i_1110, i_1111, i_1112, i_1113, i_1114, i_1489, i_1490, i_1781, i_10025, i_10101, i_10102, i_10103, i_10104, i_10109, i_10110, i_10111, i_10112, i_10350, i_10351, i_10352, i_10353, i_10574, i_10575, i_10576, i_10628, i_10632, i_10641, i_10704, i_10706, i_10711, i_10712, i_10713, i_10714, i_10715, i_10716, i_10717, i_10718, i_10729, i_10759, i_10760, i_10761, i_10762, i_10763, i_10827, i_10837, i_10838, i_10839, i_10840, i_10868, i_10869, i_10870, i_10871, i_10905, i_10906, i_10907, i_10908, i_11333, i_11334, i_11340, i_11342);

  input i_1, i_5, i_9, i_12, i_15, i_18, i_23, i_26, i_29, i_32, i_35, i_38, i_41, i_44, i_47, i_50, i_53, i_54, i_55, i_56, i_57, i_58, i_59, i_60, i_61, i_62, i_63, i_64, i_65, i_66, i_69, i_70, i_73, i_74, i_75, i_76, i_77, i_78, i_79, i_80, i_81, i_82, i_83, i_84, i_85, i_86, i_87, i_88, i_89, i_94, i_97, i_100, i_103, i_106, i_109, i_110, i_111, i_112, i_113, i_114, i_115, i_118, i_121, i_124, i_127, i_130, i_133, i_134, i_135, i_138, i_141, i_144, i_147, i_150, i_151, i_152, i_153, i_154, i_155, i_156, i_157, i_158, i_159, i_160, i_161, i_162, i_163, i_164, i_165, i_166, i_167, i_168, i_169, i_170, i_171, i_172, i_173, i_174, i_175, i_176, i_177, i_178, i_179, i_180, i_181, i_182, i_183, i_184, i_185, i_186, i_187, i_188, i_189, i_190, i_191, i_192, i_193, i_194, i_195, i_196, i_197, i_198, i_199, i_200, i_201, i_202, i_203, i_204, i_205, i_206, i_207, i_208, i_209, i_210, i_211, i_212, i_213, i_214, i_215, i_216, i_217, i_218, i_219, i_220, i_221, i_222, i_223, i_224, i_225, i_226, i_227, i_228, i_229, i_230, i_231, i_232, i_233, i_234, i_235, i_236, i_237, i_238, i_239, i_240, i_241, i_242, i_245, i_248, i_251, i_254, i_257, i_260, i_263, i_267, i_271, i_274, i_277, i_280, i_283, i_286, i_289, i_293, i_296, i_299, i_303, i_307, i_310, i_313, i_316, i_319, i_322, i_325, i_328, i_331, i_334, i_337, i_340, i_343, i_346, i_349, i_352, i_355, i_358, i_361, i_364, i_367, i_382, keyinput0, keyinput1, keyinput2, keyinput3, keyinput4, keyinput5, keyinput6, keyinput7;
  output i_241, i_387, i_388, i_478, i_482, i_484, i_486, i_489, i_492, i_501, i_505, i_507, i_509, i_511, i_513, i_515, i_517, i_519, i_535, i_537, i_539, i_541, i_543, i_545, i_547, i_549, i_551, i_553, i_556, i_559, i_561, i_563, i_565, i_567, i_569, i_571, i_573, i_582, i_643, i_707, i_813, i_881, i_882, i_883, i_884, i_885, i_889, i_945, i_1110, i_1111, i_1112, i_1113, i_1114, i_1489, i_1490, i_1781, i_10025, i_10101, i_10102, i_10103, i_10104, i_10109, i_10110, i_10111, i_10112, i_10350, i_10351, i_10352, i_10353, i_10574, i_10575, i_10576, i_10628, i_10632, i_10641, i_10704, i_10706, i_10711, i_10712, i_10713, i_10714, i_10715, i_10716, i_10717, i_10718, i_10729, i_10759, i_10760, i_10761, i_10762, i_10763, i_10827, i_10837, i_10838, i_10839, i_10840, i_10868, i_10869, i_10870, i_10871, i_10905, i_10906, i_10907, i_10908, i_11333, i_11334, i_11340, i_11342;
  wire i_10002, i_10003, i_10006, i_10007, i_10010, i_10013, i_10014, i_10015, i_10016, i_10017, i_10018, i_10019, i_10020, i_10021, i_10022, i_10023, i_10024, i_10026, i_10028, i_10032, i_10033, i_10034, i_10035, i_10036, i_10037, i_10038, i_10039, i_10040, i_10041, i_10042, i_10043, i_10050, i_10053, i_10054, i_10055, i_10056, i_10057, i_10058, i_10059, i_10060, i_10061, i_10062, i_10067, i_10070, i_10073, i_10076, i_10077, i_10082, i_10083, i_10084, i_10085, i_10086, i_10093, i_10094, i_10105, i_10106, i_10107, i_10108, i_10113, i_10114, i_10115, i_10116, i_10119, i_10124, i_10130, i_10131, i_10132, i_10133, i_10134, i_10135, i_10136, i_10137, i_10138, i_10139, i_10140, i_10141, i_10148, i_10155, i_10156, i_10157, i_10158, i_10159, i_10160, i_10161, i_10162, i_10163, i_10164, i_10165, i_10170, i_10173, i_10176, i_10177, i_10178, i_10179, i_10180, i_10183, i_10186, i_10189, i_10192, i_10195, i_10196, i_10197, i_10200, i_10203, i_10204, i_10205, i_10206, i_10212, i_10213, i_10230, i_10231, i_10232, i_10233, i_10234, i_10237, i_10238, i_10239, i_10240, i_10241, i_10242, i_10247, i_10248, i_10259, i_10264, i_10265, i_10266, i_10267, i_10268, i_10269, i_10270, i_10271, i_10272, i_10273, i_10278, i_10279, i_1028, i_10280, i_10281, i_10282, i_10283, i_10287, i_10288, i_10289, i_1029, i_10290, i_10291, i_10292, i_10293, i_10294, i_10295, i_10296, i_10299, i_10300, i_10301, i_10306, i_10307, i_10308, i_10311, i_10314, i_10315, i_10316, i_10317, i_10318, i_10321, i_10324, i_10325, i_10326, i_10327, i_10328, i_10329, i_10330, i_10331, i_10332, i_10333, i_10334, i_10337, i_10338, i_10339, i_10340, i_10341, i_10344, i_10354, i_10357, i_10360, i_10367, i_10375, i_10381, i_10388, i_10391, i_10399, i_10402, i_10406, i_10409, i_10412, i_10415, i_10419, i_10422, i_10425, i_10428, i_10431, i_10432, i_10437, i_10438, i_10439, i_10440, i_10441, i_10444, i_10445, i_10450, i_10451, i_10455, i_10456, i_10465, i_10466, i_10479, i_10497, i_10509, i_10512, i_10515, i_10516, i_10517, i_10518, i_10519, i_10522, i_10525, i_10528, i_10531, i_10534, i_10535, i_10536, i_10539, i_10542, i_10543, i_10544, i_10545, i_10546, i_10547, i_10548, i_10549, i_10550, i_10551, i_10552, i_10553, i_10554, i_10555, i_10556, i_10557, i_10558, i_10559, i_10560, i_10561, i_10562, i_10563, i_10564, i_10565, i_10566, i_10567, i_10568, i_10569, i_10570, i_10571, i_10572, i_10573, i_10577, i_10581, i_10582, i_10583, i_10587, i_10588, i_10589, i_10594, i_10595, i_10596, i_10597, i_10598, i_10602, i_10609, i_10610, i_10621, i_10626, i_10627, i_10629, i_10631, i_10637, i_10638, i_10639, i_10640, i_10642, i_10643, i_10644, i_10645, i_10647, i_10648, i_10649, i_10652, i_10659, i_10662, i_10665, i_10668, i_10671, i_10672, i_10673, i_10674, i_10675, i_10678, i_10681, i_10682, i_10683, i_10684, i_10685, i_10686, i_10687, i_10688, i_10689, i_10690, i_10691, i_10694, i_10695, i_10696, i_10697, i_10698, i_10701, i_10705, i_10707, i_10708, i_10709, i_10710, i_10719, i_10720, i_10730, i_10731, i_10737, i_10738, i_10739, i_10746, i_10747, i_10748, i_10749, i_10750, i_10753, i_10754, i_10764, i_10765, i_10766, i_10767, i_10768, i_10769, i_10770, i_10771, i_10772, i_10773, i_10774, i_10775, i_10776, i_10778, i_10781, i_10784, i_10789, i_10792, i_10796, i_10797, i_10798, i_10799, i_10800, i_10803, i_10806, i_10809, i_10812, i_10815, i_10816, i_10817, i_10820, i_10823, i_10824, i_10825, i_10826, i_10832, i_10833, i_10834, i_10835, i_10836, i_10845, i_10846, i_10857, i_10862, i_10863, i_10864, i_10865, i_10866, i_10867, i_10872, i_10873, i_10874, i_10875, i_10876, i_10879, i_10882, i_10883, i_10884, i_10885, i_10886, i_10887, i_10888, i_10889, i_10890, i_10891, i_10892, i_10895, i_10896, i_10897, i_10898, i_10899, i_10902, i_10909, i_10910, i_10915, i_10916, i_10917, i_10918, i_10919, i_10922, i_10923, i_10928, i_10931, i_10934, i_10935, i_10936, i_10937, i_10938, i_10941, i_10944, i_10947, i_10950, i_10953, i_10954, i_10955, i_10958, i_10961, i_10962, i_10963, i_10964, i_10969, i_10970, i_10981, i_10986, i_10987, i_10988, i_10989, i_10990, i_10991, i_10992, i_10995, i_10998, i_10999, i_11000, i_11001, i_11002, i_11003, i_11004, i_11005, i_11006, i_11007, i_11008, i_11011, i_11012, i_11013, i_11014, i_11015, i_11018, i_11023, i_11024, i_11027, i_11028, i_11029, i_11030, i_11031, i_11034, i_11035, i_11040, i_11041, i_11042, i_11043, i_11044, i_11047, i_11050, i_11053, i_11056, i_11059, i_11062, i_11065, i_11066, i_11067, i_11070, i_11073, i_11074, i_11075, i_11076, i_11077, i_11078, i_1109, i_11095, i_11098, i_11099, i_11100, i_11103, i_11106, i_11107, i_11108, i_11109, i_11110, i_11111, i_11112, i_11113, i_11114, i_11115, i_11116, i_11117, i_11118, i_11119, i_11120, i_11121, i_11122, i_11123, i_11124, i_11127, i_11130, i_11137, i_11138, i_11139, i_11140, i_11141, i_11142, i_11143, i_11144, i_11145, i_1115, i_11152, i_11153, i_11154, i_11155, i_11156, i_11159, i_1116, i_11162, i_11165, i_11168, i_11171, i_11174, i_11177, i_11180, i_11183, i_11184, i_11185, i_11186, i_11187, i_11188, i_1119, i_11205, i_11210, i_11211, i_11212, i_11213, i_11214, i_11215, i_11216, i_11217, i_11218, i_11219, i_11220, i_11222, i_11223, i_11224, i_11225, i_11226, i_11227, i_11228, i_11229, i_11231, i_11232, i_11233, i_11236, i_11239, i_11242, i_11243, i_11244, i_11245, i_11246, i_1125, i_11250, i_11252, i_11257, i_11260, i_11261, i_11262, i_11263, i_11264, i_11265, i_11267, i_11268, i_11269, i_11270, i_11272, i_11277, i_11278, i_11279, i_11280, i_11282, i_11283, i_11284, i_11285, i_11286, i_11288, i_11289, i_11290, i_11291, i_11292, i_11293, i_11294, i_11295, i_11296, i_11297, i_11298, i_11299, i_11302, i_11307, i_11308, i_11309, i_11312, i_11313, i_11314, i_11315, i_11316, i_11317, i_1132, i_11320, i_11321, i_11323, i_11327, i_11328, i_11329, i_11331, i_11335, i_11336, i_11337, i_11338, i_11339, i_11341, i_1136, i_1141, i_1147, i_1154, i_1160, i_1167, i_1174, i_1175, i_1182, i_1189, i_1194, i_1199, i_1206, i_1211, i_1218, i_1222, i_1227, i_1233, i_1240, i_1244, i_1249, i_1256, i_1263, i_1270, i_1277, i_1284, i_1287, i_1290, i_1293, i_1296, i_1299, i_1302, i_1305, i_1308, i_1311, i_1314, i_1317, i_1320, i_1323, i_1326, i_1329, i_1332, i_1335, i_1338, i_1341, i_1344, i_1347, i_1350, i_1353, i_1356, i_1359, i_1362, i_1365, i_1368, i_1371, i_1374, i_1377, i_1380, i_1383, i_1386, i_1389, i_1392, i_1395, i_1398, i_1401, i_1404, i_1407, i_1410, i_1413, i_1416, i_1419, i_1422, i_1425, i_1428, i_1431, i_1434, i_1437, i_1440, i_1443, i_1446, i_1449, i_1452, i_1455, i_1458, i_1461, i_1464, i_1467, i_1470, i_1473, i_1476, i_1479, i_1482, i_1485, i_1537, i_1551, i_1649, i_1703, i_1708, i_1713, i_1721, i_1758, i_1782, i_1783, i_1789, i_1793, i_1794, i_1795, i_1796, i_1797, i_1798, i_1799, i_1805, i_1811, i_1812, i_1813, i_1814, i_1815, i_1816, i_1817, i_1818, i_1819, i_1820, i_1821, i_1822, i_1828, i_1829, i_1830, i_1832, i_1833, i_1834, i_1835, i_1839, i_1840, i_1841, i_1842, i_1843, i_1845, i_1851, i_1857, i_1858, i_1859, i_1860, i_1861, i_1862, i_1863, i_1864, i_1865, i_1866, i_1867, i_1868, i_1869, i_1870, i_1871, i_1872, i_1873, i_1874, i_1875, i_1876, i_1877, i_1878, i_1879, i_1880, i_1881, i_1882, i_1883, i_1884, i_1885, i_1892, i_1899, i_1906, i_1913, i_1919, i_1926, i_1927, i_1928, i_1929, i_1930, i_1931, i_1932, i_1933, i_1934, i_1935, i_1936, i_1937, i_1938, i_1939, i_1940, i_1941, i_1942, i_1943, i_1944, i_1945, i_1946, i_1947, i_1953, i_1957, i_1958, i_1959, i_1960, i_1961, i_1962, i_1963, i_1965, i_1966, i_1967, i_1968, i_1969, i_1970, i_1971, i_1972, i_1973, i_1974, i_1975, i_1976, i_1977, i_1983, i_1989, i_1990, i_1991, i_1992, i_1993, i_1994, i_1995, i_1996, i_1997, i_2003, i_2010, i_2011, i_2012, i_2013, i_2014, i_2015, i_2016, i_2017, i_2018, i_2019, i_2020, i_2021, i_2022, i_2023, i_2024, i_2031, i_2038, i_2045, i_2052, i_2058, i_2064, i_2065, i_2066, i_2067, i_2068, i_2069, i_2070, i_2071, i_2072, i_2073, i_2074, i_2081, i_2086, i_2107, i_2108, i_2110, i_2111, i_2112, i_2113, i_2114, i_2115, i_2117, i_2171, i_2172, i_2230, i_2231, i_2235, i_2239, i_2240, i_2241, i_2242, i_2243, i_2244, i_2245, i_2246, i_2247, i_2248, i_2249, i_2250, i_2251, i_2252, i_2253, i_2254, i_2255, i_2256, i_2257, i_2267, i_2268, i_2269, i_2274, i_2275, i_2277, i_2278, i_2279, i_2280, i_2281, i_2282, i_2283, i_2284, i_2285, i_2286, i_2287, i_2293, i_2299, i_2300, i_2301, i_2302, i_2303, i_2304, i_2305, i_2306, i_2307, i_2308, i_2309, i_2315, i_2321, i_2322, i_2323, i_2324, i_2325, i_2326, i_2327, i_2328, i_2329, i_2330, i_2331, i_2337, i_2338, i_2339, i_2340, i_2341, i_2342, i_2343, i_2344, i_2345, i_2346, i_2347, i_2348, i_2349, i_2350, i_2351, i_2352, i_2353, i_2354, i_2355, i_2356, i_2357, i_2358, i_2359, i_2360, i_2361, i_2362, i_2363, i_2364, i_2365, i_2366, i_2367, i_2368, i_2374, i_2375, i_2376, i_2377, i_2378, i_2379, i_2380, i_2381, i_2382, i_2383, i_2384, i_2390, i_2396, i_2397, i_2398, i_2399, i_2400, i_2401, i_2402, i_2403, i_2404, i_2405, i_2406, i_2412, i_2418, i_2419, i_2420, i_2421, i_2422, i_2423, i_2424, i_2425, i_2426, i_2427, i_2428, i_2429, i_2430, i_2431, i_2432, i_2433, i_2434, i_2435, i_2436, i_2437, i_2441, i_2442, i_2446, i_2450, i_2454, i_2458, i_2462, i_2466, i_2470, i_2474, i_2478, i_2482, i_2488, i_2496, i_2502, i_2508, i_2523, i_2533, i_2537, i_2538, i_2542, i_2546, i_2550, i_2554, i_2561, i_2567, i_2573, i_2604, i_2607, i_2611, i_2615, i_2619, i_2626, i_2632, i_2638, i_2644, i_2650, i_2653, i_2654, i_2658, i_2662, i_2666, i_2670, i_2674, i_2680, i_2688, i_2692, i_2696, i_2700, i_2704, i_2728, i_2729, i_2733, i_2737, i_2741, i_2745, i_2749, i_2753, i_2757, i_2761, i_2765, i_2766, i_2769, i_2772, i_2775, i_2778, i_2781, i_2784, i_2787, i_2790, i_2793, i_2796, i_2866, i_2867, i_2868, i_2869, i_2878, i_2913, i_2914, i_2915, i_2916, i_2917, i_2918, i_2919, i_2920, i_2921, i_2922, i_2923, i_2924, i_2925, i_2926, i_2927, i_2928, i_2929, i_2930, i_2931, i_2932, i_2933, i_2934, i_2935, i_2936, i_2937, i_2988, i_3005, i_3006, i_3007, i_3008, i_3009, i_3020, i_3021, i_3022, i_3023, i_3024, i_3025, i_3026, i_3027, i_3028, i_3029, i_3032, i_3033, i_3034, i_3035, i_3036, i_3037, i_3038, i_3039, i_3040, i_3041, i_3061, i_3064, i_3067, i_3070, i_3073, i_3080, i_3096, i_3097, i_3101, i_3107, i_3114, i_3122, i_3126, i_3130, i_3131, i_3134, i_3135, i_3136, i_3137, i_3140, i_3144, i_3149, i_3155, i_3159, i_3167, i_3168, i_3169, i_3173, i_3178, i_3184, i_3185, i_3189, i_3195, i_3202, i_3210, i_3211, i_3215, i_3221, i_3228, i_3229, i_3232, i_3236, i_3241, i_3247, i_3251, i_3255, i_3259, i_3263, i_3267, i_3273, i_3281, i_3287, i_3293, i_3299, i_3303, i_3307, i_3311, i_3315, i_3322, i_3328, i_3334, i_3340, i_3343, i_3349, i_3355, i_3361, i_3362, i_3363, i_3364, i_3365, i_3366, i_3367, i_3368, i_3369, i_3370, i_3371, i_3372, i_3373, i_3374, i_3375, i_3379, i_3380, i_3381, i_3384, i_3390, i_3398, i_3404, i_3410, i_3416, i_3420, i_3424, i_3428, i_3432, i_3436, i_3440, i_3444, i_3448, i_3452, i_3453, i_3454, i_3458, i_3462, i_3466, i_3470, i_3474, i_3478, i_3482, i_3486, i_3487, i_3490, i_3493, i_3496, i_3499, i_3502, i_3507, i_3510, i_3515, i_3518, i_3521, i_3524, i_3527, i_3530, i_3535, i_3539, i_3542, i_3545, i_3548, i_3551, i_3552, i_3553, i_3557, i_3560, i_3563, i_3566, i_3569, i_3570, i_3571, i_3574, i_3577, i_3580, i_3583, i_3586, i_3589, i_3592, i_3595, i_3598, i_3601, i_3604, i_3607, i_3610, i_3613, i_3616, i_3619, i_3622, i_3625, i_3628, i_3631, i_3634, i_3637, i_3640, i_3643, i_3646, i_3649, i_3652, i_3655, i_3658, i_3661, i_3664, i_3667, i_3670, i_3673, i_3676, i_3679, i_3682, i_3685, i_3688, i_3691, i_3694, i_3697, i_3700, i_3703, i_3706, i_3709, i_3712, i_3715, i_3718, i_3721, i_3724, i_3727, i_3730, i_3733, i_3736, i_3739, i_3742, i_3745, i_3748, i_3751, i_3754, i_3757, i_3760, i_3763, i_3766, i_3769, i_3772, i_3775, i_3778, i_3781, i_3782, i_3783, i_3786, i_3789, i_3792, i_3795, i_3798, i_3801, i_3804, i_3807, i_3810, i_3813, i_3816, i_3819, i_3822, i_3825, i_3828, i_3831, i_3834, i_3837, i_3840, i_3843, i_3846, i_3849, i_3852, i_3855, i_3858, i_3861, i_3864, i_3867, i_3870, i_3873, i_3876, i_3879, i_3882, i_3885, i_3888, i_3891, i_3953, i_3954, i_3955, i_3956, i_3958, i_3964, i_4193, i_4303, i_4308, i_4313, i_4326, i_4327, i_4333, i_4334, i_4411, i_4412, i_4463, i_4464, i_4465, i_4466, i_4467, i_4468, i_4469, i_4470, i_4471, i_4472, i_4473, i_4474, i_4475, i_4476, i_4477, i_4478, i_4479, i_4480, i_4481, i_4482, i_4483, i_4484, i_4485, i_4486, i_4487, i_4488, i_4489, i_4490, i_4491, i_4492, i_4493, i_4494, i_4495, i_4496, i_4497, i_4498, i_4499, i_4500, i_4501, i_4502, i_4503, i_4504, i_4505, i_4506, i_4507, i_4508, i_4509, i_4510, i_4511, i_4512, i_4513, i_4514, i_4515, i_4516, i_4517, i_4518, i_4519, i_4520, i_4521, i_4522, i_4523, i_4524, i_4525, i_4526, i_4527, i_4528, i_4529, i_4530, i_4531, i_4532, i_4533, i_4534, i_4535, i_4536, i_4537, i_4538, i_4539, i_4540, i_4541, i_4542, i_4543, i_4544, i_4545, i_4549, i_4555, i_4562, i_4563, i_4566, i_4570, i_4575, i_4576, i_4577, i_4581, i_4586, i_4592, i_4593, i_4597, i_4603, i_4610, i_4611, i_4612, i_4613, i_4614, i_4615, i_4616, i_4617, i_4618, i_4619, i_4620, i_4621, i_4622, i_4623, i_4624, i_4625, i_4626, i_4627, i_4628, i_4629, i_4630, i_4631, i_4632, i_4633, i_4634, i_4635, i_4636, i_4637, i_4638, i_4639, i_4640, i_4641, i_4642, i_4643, i_4644, i_4645, i_4646, i_4647, i_4648, i_4649, i_4650, i_4651, i_4652, i_4653, i_4656, i_4657, i_4661, i_4667, i_467, i_4674, i_4675, i_4678, i_4682, i_4687, i_469, i_4693, i_4694, i_4695, i_4696, i_4697, i_4698, i_4699, i_4700, i_4701, i_4702, i_4706, i_4711, i_4717, i_4718, i_4722, i_4728, i_4735, i_4743, i_4744, i_4745, i_4746, i_4747, i_4748, i_4749, i_4750, i_4751, i_4752, i_4753, i_4754, i_4755, i_4756, i_4757, i_4758, i_4759, i_4760, i_4761, i_4762, i_4763, i_4764, i_4765, i_4766, i_4767, i_4768, i_4769, i_4775, i_4776, i_4777, i_4778, i_4779, i_4780, i_4781, i_4782, i_4783, i_4784, i_4789, i_4790, i_4793, i_4794, i_4795, i_4796, i_4799, i_4800, i_4801, i_4802, i_4803, i_4806, i_4809, i_4810, i_4813, i_4814, i_4817, i_4820, i_4823, i_4826, i_4829, i_4832, i_4835, i_4838, i_4841, i_4844, i_4847, i_4850, i_4853, i_4856, i_4859, i_4862, i_4865, i_4868, i_4871, i_4874, i_4877, i_4880, i_4883, i_4886, i_4889, i_4892, i_4895, i_4898, i_4901, i_4904, i_4907, i_4910, i_4913, i_4916, i_4919, i_4922, i_4925, i_4928, i_4931, i_4934, i_4937, i_494, i_4940, i_4943, i_4946, i_4949, i_4952, i_4955, i_4958, i_4961, i_4964, i_4967, i_4970, i_4973, i_4976, i_4979, i_4982, i_4985, i_4988, i_4991, i_4994, i_4997, i_5000, i_5003, i_5006, i_5009, i_5012, i_5015, i_5018, i_5021, i_5024, i_5027, i_5030, i_5033, i_5036, i_5039, i_5042, i_5045, i_5046, i_5047, i_5048, i_5049, i_5052, i_5055, i_5058, i_5061, i_5064, i_5065, i_5066, i_5067, i_5068, i_5071, i_5074, i_5077, i_5080, i_5083, i_5086, i_5089, i_5092, i_5095, i_5098, i_5101, i_5104, i_5107, i_5110, i_5111, i_5112, i_5113, i_5114, i_5117, i_5120, i_5123, i_5126, i_5129, i_5132, i_5135, i_5138, i_5141, i_5144, i_5147, i_5150, i_5153, i_5156, i_5159, i_5162, i_5165, i_5166, i_5167, i_5168, i_5169, i_5170, i_5171, i_5172, i_5173, i_5174, i_5175, i_5176, i_5177, i_5178, i_5179, i_5180, i_5181, i_5182, i_5183, i_5184, i_5185, i_5186, i_5187, i_5188, i_5189, i_5190, i_5191, i_5192, i_5193, i_5196, i_5197, i_5198, i_5199, i_5200, i_5201, i_5202, i_5203, i_5204, i_5205, i_5206, i_5207, i_5208, i_5209, i_5210, i_5211, i_5212, i_5213, i_528, i_5283, i_5284, i_5285, i_5286, i_5287, i_5288, i_5289, i_5290, i_5291, i_5292, i_5293, i_5294, i_5295, i_5296, i_5297, i_5298, i_5299, i_5300, i_5314, i_5315, i_5316, i_5317, i_5318, i_5319, i_5320, i_5321, i_5322, i_5323, i_5324, i_5363, i_5364, i_5365, i_5366, i_5367, i_5425, i_5426, i_5427, i_5429, i_5430, i_5431, i_5432, i_5433, i_5451, i_5452, i_5453, i_5454, i_5455, i_5456, i_5457, i_5469, i_5474, i_5475, i_5476, i_5477, i_5571, i_5572, i_5573, i_5574, i_5584, i_5585, i_5586, i_5587, i_5602, i_5603, i_5604, i_5605, i_5631, i_5632, i_5640, i_5654, i_5670, i_5683, i_5690, i_5697, i_5707, i_5718, i_5728, i_5735, i_5736, i_5740, i_5744, i_5747, i_575, i_5751, i_5755, i_5758, i_5762, i_5766, i_5769, i_5770, i_5771, i_5778, i_578, i_5789, i_5799, i_5807, i_5821, i_5837, i_585, i_5850, i_5856, i_5863, i_5870, i_5881, i_5892, i_5898, i_590, i_5905, i_5915, i_5926, i_593, i_5936, i_5943, i_5944, i_5945, i_5946, i_5947, i_5948, i_5949, i_5950, i_5951, i_5952, i_5953, i_5954, i_5955, i_5956, i_5957, i_5958, i_5959, i_596, i_5960, i_5966, i_5967, i_5968, i_5969, i_5970, i_5971, i_5972, i_5973, i_5974, i_5975, i_5976, i_5977, i_5978, i_5979, i_5980, i_5981, i_5989, i_599, i_5990, i_5991, i_5996, i_6000, i_6003, i_6009, i_6014, i_6018, i_6021, i_6022, i_6023, i_6024, i_6025, i_6026, i_6027, i_6028, i_6029, i_6030, i_6031, i_6032, i_6033, i_6034, i_6035, i_6036, i_6037, i_6038, i_6039, i_604, i_6040, i_6041, i_6047, i_6052, i_6056, i_6059, i_6060, i_6061, i_6062, i_6063, i_6064, i_6065, i_6066, i_6067, i_6068, i_6069, i_6070, i_6071, i_6072, i_6073, i_6074, i_6075, i_6076, i_6077, i_6078, i_6079, i_6083, i_6087, i_609, i_6090, i_6091, i_6092, i_6093, i_6094, i_6095, i_6096, i_6097, i_6098, i_6099, i_6100, i_6101, i_6102, i_6103, i_6104, i_6105, i_6106, i_6107, i_6108, i_6109, i_6110, i_6111, i_6112, i_6113, i_6114, i_6115, i_6116, i_6117, i_6118, i_6119, i_6120, i_6121, i_6122, i_6123, i_6124, i_6125, i_6126, i_6127, i_6131, i_6135, i_6136, i_6137, i_614, i_6141, i_6145, i_6148, i_6149, i_6150, i_6151, i_6152, i_6153, i_6154, i_6155, i_6156, i_6157, i_6158, i_6159, i_6160, i_6161, i_6162, i_6163, i_6164, i_6165, i_6166, i_6170, i_6174, i_6177, i_6181, i_6182, i_6183, i_6184, i_6185, i_6186, i_6187, i_6188, i_6189, i_6190, i_6191, i_6192, i_6193, i_6194, i_6195, i_6196, i_6199, i_6202, i_6203, i_6204, i_6207, i_6210, i_6213, i_6214, i_6217, i_6220, i_6223, i_6224, i_6225, i_6226, i_6227, i_6228, i_6229, i_6230, i_6231, i_6232, i_6235, i_6236, i_6239, i_6240, i_6241, i_6242, i_6243, i_6246, i_6249, i_625, i_6252, i_6255, i_6256, i_6257, i_6258, i_6259, i_6260, i_6261, i_6262, i_6263, i_6266, i_628, i_632, i_636, i_641, i_642, i_644, i_651, i_6540, i_6541, i_6542, i_6543, i_6544, i_6545, i_6546, i_6547, i_6555, i_6556, i_6557, i_6558, i_6559, i_6560, i_6561, i_6569, i_657, i_6594, i_6595, i_6596, i_6597, i_6598, i_6599, i_660, i_6600, i_6601, i_6602, i_6603, i_6604, i_6605, i_6606, i_6621, i_6622, i_6623, i_6624, i_6625, i_6626, i_6627, i_6628, i_6629, i_6639, i_6640, i_6641, i_6642, i_6643, i_6644, i_6645, i_6646, i_6647, i_6648, i_6649, i_6650, i_6651, i_6652, i_6653, i_6654, i_6655, i_6656, i_6657, i_6658, i_6659, i_666, i_6660, i_6661, i_6668, i_6677, i_6678, i_6679, i_6680, i_6681, i_6682, i_6683, i_6684, i_6685, i_6686, i_6687, i_6688, i_6689, i_6690, i_6702, i_6703, i_6704, i_6705, i_6706, i_6707, i_6708, i_6709, i_6710, i_6711, i_6712, i_672, i_6729, i_673, i_6730, i_6731, i_6732, i_6733, i_6734, i_6735, i_6736, i_674, i_6741, i_6742, i_6743, i_6744, i_6751, i_6752, i_6753, i_6754, i_6755, i_6756, i_6757, i_6758, i_676, i_6761, i_6762, i_6766, i_6767, i_6768, i_6769, i_6770, i_6771, i_6772, i_6773, i_6774, i_6775, i_6776, i_6777, i_6778, i_6779, i_6780, i_6781, i_6782, i_6783, i_6784, i_6787, i_6788, i_6789, i_6790, i_6791, i_6792, i_6793, i_6794, i_6795, i_6796, i_6797, i_6800, i_6803, i_6806, i_6809, i_6812, i_6815, i_6818, i_682, i_6821, i_6824, i_6827, i_6830, i_6833, i_6836, i_6837, i_6838, i_6839, i_6840, i_6841, i_6842, i_6843, i_6844, i_6845, i_6848, i_6849, i_6850, i_6851, i_6852, i_6853, i_6854, i_6855, i_6856, i_6857, i_6858, i_6859, i_6860, i_6861, i_6862, i_6863, i_6864, i_6865, i_6866, i_6867, i_6870, i_6871, i_6872, i_6873, i_6874, i_6875, i_6876, i_6877, i_6878, i_6879, i_688, i_6880, i_6881, i_6884, i_6885, i_6886, i_6887, i_6888, i_6889, i_689, i_6890, i_6891, i_6892, i_6893, i_6894, i_6901, i_6912, i_6923, i_6929, i_6936, i_6946, i_695, i_6957, i_6967, i_6968, i_6969, i_6970, i_6977, i_6988, i_6998, i_700, i_7006, i_7020, i_7036, i_7049, i_705, i_7055, i_7056, i_7057, i_706, i_7060, i_7061, i_7062, i_7063, i_7064, i_7065, i_7066, i_7067, i_7068, i_7073, i_7077, i_708, i_7080, i_7086, i_7091, i_7095, i_7098, i_7099, i_7100, i_7103, i_7104, i_7105, i_7106, i_7107, i_7114, i_7125, i_7136, i_7142, i_7149, i_715, i_7159, i_7170, i_7180, i_7187, i_7188, i_7191, i_7194, i_7198, i_7202, i_7205, i_7209, i_721, i_7213, i_7216, i_7219, i_7222, i_7229, i_7240, i_7250, i_7258, i_727, i_7272, i_7288, i_7301, i_7307, i_7314, i_7318, i_7322, i_7325, i_7328, i_733, i_7331, i_7334, i_7337, i_734, i_7340, i_7343, i_7346, i_7351, i_7355, i_7358, i_7364, i_7369, i_7373, i_7376, i_7377, i_7378, i_7381, i_7384, i_7387, i_7391, i_7394, i_7398, i_7402, i_7405, i_7408, i_7411, i_7414, i_7417, i_742, i_7420, i_7423, i_7426, i_7429, i_7432, i_7435, i_7438, i_7441, i_7444, i_7447, i_7450, i_7453, i_7456, i_7459, i_7462, i_7465, i_7468, i_7471, i_7474, i_7477, i_7478, i_7479, i_748, i_7482, i_7485, i_7488, i_749, i_7491, i_7494, i_7497, i_750, i_7500, i_7503, i_7506, i_7509, i_7512, i_7515, i_7518, i_7521, i_7524, i_7527, i_7530, i_7533, i_7536, i_7539, i_7542, i_7545, i_7548, i_7551, i_7552, i_7553, i_7556, i_7557, i_7558, i_7559, i_7560, i_7563, i_7566, i_7569, i_7572, i_7573, i_7574, i_7577, i_758, i_7580, i_7581, i_7582, i_7585, i_7588, i_759, i_7591, i_7609, i_7613, i_762, i_7620, i_7649, i_7650, i_7655, i_7659, i_7668, i_7671, i_768, i_774, i_7744, i_780, i_7822, i_7825, i_7826, i_7852, i_786, i_794, i_800, i_806, i_8114, i_8117, i_812, i_8131, i_8134, i_814, i_8144, i_8145, i_8146, i_8156, i_8166, i_8169, i_8183, i_8186, i_8196, i_8200, i_8204, i_8208, i_821, i_8216, i_8217, i_8218, i_8219, i_8232, i_8233, i_8242, i_8243, i_8244, i_8245, i_8246, i_8247, i_8248, i_8249, i_8250, i_8251, i_8252, i_8253, i_8254, i_8260, i_8261, i_8262, i_8269, i_827, i_8274, i_8275, i_8276, i_8277, i_8278, i_8279, i_8280, i_8281, i_8282, i_8283, i_8284, i_8285, i_8288, i_8294, i_8295, i_8296, i_8297, i_8298, i_8307, i_8315, i_8317, i_8319, i_8321, i_8322, i_8323, i_8324, i_8325, i_8326, i_833, i_8333, i_8337, i_8338, i_8339, i_8340, i_8341, i_8342, i_8343, i_8344, i_8345, i_8346, i_8347, i_8348, i_8349, i_8350, i_8351, i_8352, i_8353, i_8354, i_8355, i_8356, i_8357, i_8358, i_8365, i_8369, i_8370, i_8371, i_8372, i_8373, i_8374, i_8375, i_8376, i_8377, i_8378, i_8379, i_8380, i_8381, i_8382, i_8383, i_8384, i_8385, i_8386, i_8387, i_8388, i_8389, i_839, i_8390, i_8391, i_8392, i_8393, i_8394, i_8404, i_8405, i_8409, i_8410, i_8411, i_8412, i_8415, i_8416, i_8417, i_8418, i_8421, i_8430, i_8433, i_8434, i_8435, i_8436, i_8437, i_8438, i_8439, i_8440, i_8441, i_8442, i_8443, i_8444, i_8447, i_8448, i_8449, i_845, i_8450, i_8451, i_8452, i_8453, i_8454, i_8455, i_8456, i_8457, i_8460, i_8463, i_8466, i_8469, i_8470, i_8471, i_8474, i_8477, i_8480, i_8483, i_8484, i_8485, i_8488, i_8489, i_8490, i_8491, i_8492, i_8493, i_8494, i_8495, i_8496, i_8497, i_8500, i_8501, i_8502, i_8503, i_8504, i_8505, i_8506, i_8507, i_8508, i_8509, i_8510, i_8511, i_8512, i_8513, i_8514, i_8515, i_8516, i_8517, i_8518, i_8519, i_8522, i_8525, i_8528, i_853, i_8531, i_8534, i_8537, i_8538, i_8539, i_8540, i_8541, i_8545, i_8546, i_8547, i_8548, i_8551, i_8552, i_8553, i_8554, i_8555, i_8558, i_8561, i_8564, i_8565, i_8566, i_8569, i_8572, i_8575, i_8578, i_8579, i_8580, i_8583, i_8586, i_8589, i_859, i_8592, i_8595, i_8598, i_8601, i_8604, i_8607, i_8608, i_8609, i_8610, i_8615, i_8616, i_8617, i_8618, i_8619, i_8624, i_8625, i_8626, i_8627, i_8632, i_8633, i_8634, i_8637, i_8638, i_8639, i_8644, i_8645, i_8646, i_8647, i_8648, i_865, i_8653, i_8654, i_8655, i_8660, i_8663, i_8666, i_8669, i_8672, i_8675, i_8678, i_8681, i_8684, i_8687, i_8690, i_8693, i_8696, i_8699, i_8702, i_8705, i_8708, i_871, i_8711, i_8714, i_8717, i_8718, i_8721, i_8724, i_8727, i_8730, i_8733, i_8734, i_8735, i_8738, i_8741, i_8744, i_8747, i_8750, i_8753, i_8754, i_8755, i_8756, i_8757, i_8760, i_8763, i_8766, i_8769, i_8772, i_8775, i_8778, i_8781, i_8784, i_8787, i_8790, i_8793, i_8796, i_8799, i_8802, i_8805, i_8808, i_8811, i_8814, i_8815, i_8816, i_8817, i_8818, i_8840, i_8857, i_886, i_8861, i_8862, i_8863, i_8864, i_8865, i_8866, i_887, i_8871, i_8874, i_8878, i_8879, i_8880, i_8881, i_8882, i_8883, i_8884, i_8885, i_8886, i_8887, i_8888, i_8898, i_8902, i_8920, i_8924, i_8927, i_8931, i_8943, i_8950, i_8956, i_8959, i_8960, i_8963, i_8966, i_8991, i_8992, i_8995, i_8996, i_9001, i_9005, i_9024, i_9025, i_9029, i_9035, i_9053, i_9054, i_9064, i_9065, i_9066, i_9067, i_9068, i_9071, i_9072, i_9073, i_9074, i_9077, i_9079, i_9082, i_9083, i_9086, i_9087, i_9088, i_9089, i_9092, i_9093, i_9094, i_9095, i_9098, i_9099, i_9103, i_9107, i_9111, i_9117, i_9127, i_9146, i_9149, i_9159, i_9160, i_9161, i_9165, i_9169, i_9173, i_9179, i_9180, i_9181, i_9182, i_9183, i_9193, i_9203, i_9206, i_9220, i_9223, i_9234, i_9235, i_9236, i_9237, i_9238, i_9242, i_9243, i_9244, i_9245, i_9246, i_9247, i_9248, i_9249, i_9250, i_9251, i_9252, i_9256, i_9257, i_9258, i_9259, i_9260, i_9261, i_9262, i_9265, i_9268, i_9271, i_9272, i_9273, i_9274, i_9275, i_9276, i_9280, i_9285, i_9286, i_9287, i_9288, i_9290, i_9292, i_9294, i_9296, i_9297, i_9298, i_9299, i_9300, i_9301, i_9307, i_9314, i_9315, i_9318, i_9319, i_9320, i_9321, i_9322, i_9323, i_9324, i_9326, i_9332, i_9339, i_9344, i_9352, i_9354, i_9356, i_9358, i_9359, i_9360, i_9361, i_9362, i_9363, i_9364, i_9365, i_9366, i_9367, i_9368, i_9369, i_9370, i_9371, i_9372, i_9375, i_9381, i_9382, i_9383, i_9384, i_9385, i_9392, i_9393, i_9394, i_9395, i_9396, i_9397, i_9398, i_9399, i_9400, i_9401, i_9402, i_9407, i_9408, i_9412, i_9413, i_9414, i_9415, i_9416, i_9417, i_9418, i_9419, i_9420, i_9421, i_9422, i_9423, i_9426, i_9429, i_9432, i_9435, i_9442, i_9445, i_9454, i_9455, i_9456, i_9459, i_9460, i_9461, i_9462, i_9465, i_9466, i_9467, i_9468, i_9473, i_9476, i_9477, i_9478, i_9485, i_9488, i_9493, i_9494, i_9495, i_9498, i_9499, i_9500, i_9505, i_9506, i_9507, i_9508, i_9509, i_9514, i_9515, i_9516, i_9517, i_9520, i_9526, i_9531, i_9539, i_9540, i_9541, i_9543, i_9551, i_9555, i_9556, i_9557, i_9560, i_9561, i_9562, i_9563, i_9564, i_9565, i_9566, i_9567, i_9568, i_9569, i_957, i_9570, i_9571, i_9575, i_9579, i_9581, i_9582, i_9585, i_9591, i_9592, i_9593, i_9594, i_9595, i_9596, i_9597, i_9598, i_9599, i_9600, i_9601, i_9602, i_9603, i_9604, i_9605, i_9608, i_9611, i_9612, i_9613, i_9614, i_9615, i_9616, i_9617, i_9618, i_9621, i_9622, i_9623, i_9624, i_9626, i_9629, i_9632, i_9635, i_9642, i_9645, i_9646, i_9649, i_9650, i_9653, i_9656, i_9659, i_9660, i_9661, i_9662, i_9663, i_9666, i_9667, i_9670, i_9671, i_9674, i_9675, i_9678, i_9679, i_9682, i_9685, i_9690, i_9691, i_9692, i_9695, i_9698, i_9702, i_9707, i_9710, i_9711, i_9714, i_9715, i_9716, i_9717, i_9720, i_9721, i_9722, i_9723, i_9726, i_9727, i_9732, i_9733, i_9734, i_9735, i_9736, i_9737, i_9738, i_9739, i_9740, i_9741, i_9742, i_9754, i_9758, i_9762, i_9763, i_9764, i_9765, i_9766, i_9767, i_9768, i_9769, i_9773, i_9774, i_9775, i_9779, i_9784, i_9785, i_9786, i_9790, i_9791, i_9795, i_9796, i_9797, i_9798, i_9799, i_9800, i_9801, i_9802, i_9803, i_9805, i_9806, i_9809, i_9813, i_9814, i_9815, i_9816, i_9817, i_9820, i_9825, i_9826, i_9827, i_9828, i_9829, i_9830, i_9835, i_9836, i_9837, i_9838, i_9846, i_9847, i_9862, i_9863, i_9866, i_9873, i_9876, i_9890, i_9891, i_9892, i_9893, i_9894, i_9895, i_9896, i_9897, i_9898, i_9899, i_9900, i_9901, i_9902, i_9903, i_9904, i_9905, i_9906, i_9907, i_9908, i_9909, i_9910, i_9911, i_9917, i_9923, i_9924, i_9925, i_9932, i_9935, i_9938, i_9939, i_9945, i_9946, i_9947, i_9948, i_9949, i_9953, i_9954, i_9955, i_9956, i_9957, i_9958, i_9959, i_9960, i_9961, i_9964, i_9967, i_9968, i_9969, i_9970, i_9971, i_9972, i_9973, i_9974, i_9975, i_9976, i_9977, i_9978, i_9979, i_9982, i_9983, i_9986, i_9989, i_9992, i_9995, i_9996, i_9997, i_9998, i_9999, i_10111_in, flip_signal;

  not ginst2 (i_10002, i_9717);
  nand ginst3 (i_10003, i_9722, i_9876);
  not ginst4 (i_10006, i_9723);
  nand ginst5 (i_10007, i_9829, i_9830);
  nand ginst6 (i_10010, i_9827, i_9828);
  and ginst7 (i_10013, i_8269, i_8307, i_9791);
  and ginst8 (i_10014, i_8269, i_8307, i_9344, i_9758);
  and ginst9 (i_10015, i_367, i_8269, i_8307, i_9344, i_9754);
  and ginst10 (i_10016, i_8394, i_8421, i_9786);
  and ginst11 (i_10017, i_8394, i_8421, i_9332, i_9820);
  and ginst12 (i_10018, i_8394, i_8421, i_9786);
  and ginst13 (i_10019, i_8394, i_8421, i_9332, i_9820);
  and ginst14 (i_10020, i_8262, i_8298, i_9809);
  and ginst15 (i_10021, i_8262, i_8298, i_9385, i_9779);
  and ginst16 (i_10022, i_367, i_8262, i_8298, i_9385, i_9775);
  not ginst17 (i_10023, i_9945);
  not ginst18 (i_10024, i_9946);
  nand ginst19 (i_10025, i_9740, i_9893);
  not ginst20 (i_10026, i_9923);
  not ginst21 (i_10028, i_9924);
  nand ginst22 (i_10032, i_8595, i_9897);
  nand ginst23 (i_10033, i_8598, i_9899);
  nand ginst24 (i_10034, i_8601, i_9901);
  nand ginst25 (i_10035, i_8604, i_9903);
  nand ginst26 (i_10036, i_4803, i_9906);
  nand ginst27 (i_10037, i_4806, i_9908);
  nand ginst28 (i_10038, i_8627, i_9910);
  and ginst29 (i_10039, i_8298, i_9809);
  and ginst30 (i_10040, i_8298, i_9385, i_9779);
  and ginst31 (i_10041, i_367, i_8298, i_9385, i_9775);
  and ginst32 (i_10042, i_9385, i_9779);
  and ginst33 (i_10043, i_367, i_9385, i_9775);
  nand ginst34 (i_10050, i_8727, i_9938);
  not ginst35 (i_10053, i_9817);
  and ginst36 (i_10054, i_9029, i_9817);
  and ginst37 (i_10055, i_8394, i_9786);
  and ginst38 (i_10056, i_8394, i_9332, i_9820);
  and ginst39 (i_10057, i_8307, i_9791);
  and ginst40 (i_10058, i_8307, i_9344, i_9758);
  and ginst41 (i_10059, i_367, i_8307, i_9344, i_9754);
  and ginst42 (i_10060, i_9344, i_9758);
  and ginst43 (i_10061, i_367, i_9344, i_9754);
  nand ginst44 (i_10062, i_4997, i_9947);
  nand ginst45 (i_10067, i_8811, i_9953);
  nand ginst46 (i_10070, i_9836, i_9955);
  nand ginst47 (i_10073, i_9838, i_9956);
  nand ginst48 (i_10076, i_9068, i_9957);
  nand ginst49 (i_10077, i_9074, i_9959);
  nand ginst50 (i_10082, i_9089, i_9967);
  nand ginst51 (i_10083, i_9095, i_9969);
  nand ginst52 (i_10084, i_4871, i_9971);
  nand ginst53 (i_10085, i_6214, i_9973);
  nand ginst54 (i_10086, i_6217, i_9975);
  nand ginst55 (i_10093, i_5027, i_9995);
  nand ginst56 (i_10094, i_6232, i_9997);
  or ginst57 (i_10101, i_10013, i_10014, i_10015, i_9238, i_9732);
  or ginst58 (i_10102, i_10016, i_10017, i_9339, i_9526, i_9734);
  or ginst59 (i_10103, i_10018, i_10019, i_9339, i_9531, i_9735);
  or ginst60 (i_10104, i_10020, i_10021, i_10022, i_9242, i_9736);
  and ginst61 (i_10105, i_9894, i_9925);
  and ginst62 (i_10106, i_9895, i_9925);
  and ginst63 (i_10107, i_9896, i_9925);
  and ginst64 (i_10108, i_8253, i_9925);
  nand ginst65 (i_10109, i_10032, i_9898);
  nand ginst66 (i_10110, i_10033, i_9900);
  xor ginst67 (i_10111, i_10111_in, flip_signal);
  nand ginst68 (i_10111_in, i_10034, i_9902);
  nand ginst69 (i_10112, i_10035, i_9904);
  nand ginst70 (i_10113, i_10036, i_9907);
  nand ginst71 (i_10114, i_10037, i_9909);
  nand ginst72 (i_10115, i_10038, i_9911);
  or ginst73 (i_10116, i_10039, i_10040, i_10041, i_9265);
  or ginst74 (i_10119, i_10042, i_10043, i_9809);
  not ginst75 (i_10124, i_9925);
  and ginst76 (i_10130, i_9768, i_9925);
  not ginst77 (i_10131, i_9932);
  not ginst78 (i_10132, i_9935);
  and ginst79 (i_10133, i_8920, i_9932);
  nand ginst80 (i_10134, i_10050, i_9939);
  not ginst81 (i_10135, i_9983);
  nand ginst82 (i_10136, i_9324, i_9983);
  not ginst83 (i_10137, i_9986);
  nand ginst84 (i_10138, i_9784, i_9986);
  and ginst85 (i_10139, i_10053, i_9785);
  or ginst86 (i_10140, i_10055, i_10056, i_8943, i_9790);
  or ginst87 (i_10141, i_10057, i_10058, i_10059, i_9268);
  or ginst88 (i_10148, i_10060, i_10061, i_9791);
  nand ginst89 (i_10155, i_10062, i_9948);
  not ginst90 (i_10156, i_9989);
  nand ginst91 (i_10157, i_9805, i_9989);
  not ginst92 (i_10158, i_9992);
  nand ginst93 (i_10159, i_9806, i_9992);
  not ginst94 (i_10160, i_9949);
  nand ginst95 (i_10161, i_10067, i_9954);
  not ginst96 (i_10162, i_10007);
  nand ginst97 (i_10163, i_10007, i_9825);
  not ginst98 (i_10164, i_10010);
  nand ginst99 (i_10165, i_10010, i_9826);
  nand ginst100 (i_10170, i_10076, i_9958);
  nand ginst101 (i_10173, i_10077, i_9960);
  not ginst102 (i_10176, i_9961);
  nand ginst103 (i_10177, i_9082, i_9961);
  not ginst104 (i_10178, i_9964);
  nand ginst105 (i_10179, i_9086, i_9964);
  nand ginst106 (i_10180, i_10082, i_9968);
  nand ginst107 (i_10183, i_10083, i_9970);
  nand ginst108 (i_10186, i_10084, i_9972);
  nand ginst109 (i_10189, i_10085, i_9974);
  nand ginst110 (i_10192, i_10086, i_9976);
  not ginst111 (i_10195, i_9979);
  nand ginst112 (i_10196, i_9979, i_9982);
  nand ginst113 (i_10197, i_10093, i_9996);
  nand ginst114 (i_10200, i_10094, i_9998);
  not ginst115 (i_10203, i_9999);
  nand ginst116 (i_10204, i_10002, i_9999);
  not ginst117 (i_10205, i_10003);
  nand ginst118 (i_10206, i_10003, i_10006);
  nand ginst119 (i_10212, i_10070, i_4308);
  nand ginst120 (i_10213, i_10073, i_4313);
  and ginst121 (i_10230, i_10131, i_9774);
  nand ginst122 (i_10231, i_10135, i_8730);
  nand ginst123 (i_10232, i_10137, i_9478);
  or ginst124 (i_10233, i_10054, i_10139);
  nand ginst125 (i_10234, i_10140, i_7100);
  nand ginst126 (i_10237, i_10156, i_9485);
  nand ginst127 (i_10238, i_10158, i_9488);
  nand ginst128 (i_10239, i_10162, i_9517);
  nand ginst129 (i_10240, i_10164, i_9520);
  not ginst130 (i_10241, i_10070);
  not ginst131 (i_10242, i_10073);
  nand ginst132 (i_10247, i_10176, i_8146);
  nand ginst133 (i_10248, i_10178, i_8156);
  nand ginst134 (i_10259, i_10195, i_9692);
  nand ginst135 (i_10264, i_10203, i_9717);
  nand ginst136 (i_10265, i_10205, i_9723);
  and ginst137 (i_10266, i_10026, i_10124);
  and ginst138 (i_10267, i_10028, i_10124);
  and ginst139 (i_10268, i_10124, i_9742);
  and ginst140 (i_10269, i_10124, i_6923);
  nand ginst141 (i_10270, i_10116, i_6762);
  nand ginst142 (i_10271, i_10241, i_3061);
  nand ginst143 (i_10272, i_10242, i_3064);
  not ginst144 (i_10273, i_10116);
  and ginst145 (i_10278, i_10141, i_5697, i_5707, i_5718, i_5728);
  and ginst146 (i_10279, i_10141, i_5707, i_5718, i_5728);
  and ginst147 (i_1028, i_382, i_641);
  and ginst148 (i_10280, i_10141, i_5718, i_5728);
  and ginst149 (i_10281, i_10141, i_5728);
  and ginst150 (i_10282, i_10141, i_6784);
  not ginst151 (i_10283, i_10119);
  and ginst152 (i_10287, i_10148, i_5905, i_5915, i_5926, i_5936);
  and ginst153 (i_10288, i_10148, i_5915, i_5926, i_5936);
  and ginst154 (i_10289, i_10148, i_5926, i_5936);
  nand ginst155 (i_1029, i_382, i_705);
  and ginst156 (i_10290, i_10148, i_5936);
  and ginst157 (i_10291, i_10148, i_6881);
  and ginst158 (i_10292, i_10124, i_8898);
  nand ginst159 (i_10293, i_10136, i_10231);
  nand ginst160 (i_10294, i_10138, i_10232);
  nand ginst161 (i_10295, i_10233, i_8412);
  and ginst162 (i_10296, i_10234, i_8959);
  nand ginst163 (i_10299, i_10157, i_10237);
  nand ginst164 (i_10300, i_10159, i_10238);
  or ginst165 (i_10301, i_10133, i_10230);
  nand ginst166 (i_10306, i_10163, i_10239);
  nand ginst167 (i_10307, i_10165, i_10240);
  not ginst168 (i_10308, i_10148);
  not ginst169 (i_10311, i_10141);
  not ginst170 (i_10314, i_10170);
  nand ginst171 (i_10315, i_10170, i_9071);
  not ginst172 (i_10316, i_10173);
  nand ginst173 (i_10317, i_10173, i_9077);
  nand ginst174 (i_10318, i_10177, i_10247);
  nand ginst175 (i_10321, i_10179, i_10248);
  not ginst176 (i_10324, i_10180);
  nand ginst177 (i_10325, i_10180, i_9092);
  not ginst178 (i_10326, i_10183);
  nand ginst179 (i_10327, i_10183, i_9098);
  not ginst180 (i_10328, i_10186);
  nand ginst181 (i_10329, i_10186, i_9674);
  not ginst182 (i_10330, i_10189);
  nand ginst183 (i_10331, i_10189, i_9678);
  not ginst184 (i_10332, i_10192);
  nand ginst185 (i_10333, i_10192, i_9977);
  nand ginst186 (i_10334, i_10196, i_10259);
  not ginst187 (i_10337, i_10197);
  nand ginst188 (i_10338, i_10197, i_9710);
  not ginst189 (i_10339, i_10200);
  nand ginst190 (i_10340, i_10200, i_9714);
  nand ginst191 (i_10341, i_10204, i_10264);
  nand ginst192 (i_10344, i_10206, i_10265);
  or ginst193 (i_10350, i_10105, i_10266);
  or ginst194 (i_10351, i_10106, i_10267);
  or ginst195 (i_10352, i_10107, i_10268);
  or ginst196 (i_10353, i_10108, i_10269);
  and ginst197 (i_10354, i_10270, i_8857);
  nand ginst198 (i_10357, i_10212, i_10271);
  nand ginst199 (i_10360, i_10213, i_10272);
  or ginst200 (i_10367, i_10282, i_7620);
  or ginst201 (i_10375, i_10291, i_7671);
  or ginst202 (i_10381, i_10130, i_10292);
  and ginst203 (i_10388, i_10114, i_10134, i_10293, i_10294);
  and ginst204 (i_10391, i_10295, i_9582);
  and ginst205 (i_10399, i_10113, i_10115, i_10299, i_10300);
  and ginst206 (i_10402, i_10155, i_10161, i_10306, i_10307);
  or ginst207 (i_10406, i_10287, i_3229, i_6888, i_6889, i_6890);
  or ginst208 (i_10409, i_10288, i_3232, i_6891, i_6892);
  or ginst209 (i_10412, i_10289, i_3236, i_6893);
  or ginst210 (i_10415, i_10290, i_3241);
  or ginst211 (i_10419, i_10278, i_3137, i_6791, i_6792, i_6793);
  or ginst212 (i_10422, i_10279, i_3140, i_6794, i_6795);
  or ginst213 (i_10425, i_10280, i_3144, i_6796);
  or ginst214 (i_10428, i_10281, i_3149);
  nand ginst215 (i_10431, i_10314, i_8117);
  nand ginst216 (i_10432, i_10316, i_8134);
  nand ginst217 (i_10437, i_10324, i_8169);
  nand ginst218 (i_10438, i_10326, i_8186);
  nand ginst219 (i_10439, i_10328, i_9117);
  nand ginst220 (i_10440, i_10330, i_9127);
  nand ginst221 (i_10441, i_10332, i_9682);
  nand ginst222 (i_10444, i_10337, i_9183);
  nand ginst223 (i_10445, i_10339, i_9193);
  not ginst224 (i_10450, i_10296);
  and ginst225 (i_10451, i_10296, i_4193);
  not ginst226 (i_10455, i_10308);
  nand ginst227 (i_10456, i_10308, i_8242);
  not ginst228 (i_10465, i_10311);
  nand ginst229 (i_10466, i_10311, i_8247);
  not ginst230 (i_10479, i_10273);
  not ginst231 (i_10497, i_10301);
  nand ginst232 (i_10509, i_10315, i_10431);
  nand ginst233 (i_10512, i_10317, i_10432);
  not ginst234 (i_10515, i_10318);
  nand ginst235 (i_10516, i_10318, i_8632);
  not ginst236 (i_10517, i_10321);
  nand ginst237 (i_10518, i_10321, i_8637);
  nand ginst238 (i_10519, i_10325, i_10437);
  nand ginst239 (i_10522, i_10327, i_10438);
  nand ginst240 (i_10525, i_10329, i_10439);
  nand ginst241 (i_10528, i_10331, i_10440);
  nand ginst242 (i_10531, i_10333, i_10441);
  not ginst243 (i_10534, i_10334);
  nand ginst244 (i_10535, i_10334, i_9695);
  nand ginst245 (i_10536, i_10338, i_10444);
  nand ginst246 (i_10539, i_10340, i_10445);
  not ginst247 (i_10542, i_10341);
  nand ginst248 (i_10543, i_10341, i_9720);
  not ginst249 (i_10544, i_10344);
  nand ginst250 (i_10545, i_10344, i_9726);
  and ginst251 (i_10546, i_10450, i_5631);
  not ginst252 (i_10547, i_10391);
  and ginst253 (i_10548, i_10391, i_8950);
  and ginst254 (i_10549, i_10367, i_5165);
  not ginst255 (i_10550, i_10354);
  and ginst256 (i_10551, i_10354, i_3126);
  nand ginst257 (i_10552, i_10455, i_7411);
  and ginst258 (i_10553, i_10375, i_9539);
  and ginst259 (i_10554, i_10375, i_9540);
  and ginst260 (i_10555, i_10375, i_9541);
  and ginst261 (i_10556, i_10375, i_6761);
  not ginst262 (i_10557, i_10406);
  nand ginst263 (i_10558, i_10406, i_8243);
  not ginst264 (i_10559, i_10409);
  nand ginst265 (i_10560, i_10409, i_8244);
  not ginst266 (i_10561, i_10412);
  nand ginst267 (i_10562, i_10412, i_8245);
  not ginst268 (i_10563, i_10415);
  nand ginst269 (i_10564, i_10415, i_8246);
  nand ginst270 (i_10565, i_10465, i_7426);
  not ginst271 (i_10566, i_10419);
  nand ginst272 (i_10567, i_10419, i_8248);
  not ginst273 (i_10568, i_10422);
  nand ginst274 (i_10569, i_10422, i_8249);
  not ginst275 (i_10570, i_10425);
  nand ginst276 (i_10571, i_10425, i_8250);
  not ginst277 (i_10572, i_10428);
  nand ginst278 (i_10573, i_10428, i_8251);
  not ginst279 (i_10574, i_10399);
  not ginst280 (i_10575, i_10402);
  not ginst281 (i_10576, i_10388);
  and ginst282 (i_10577, i_10388, i_10399, i_10402);
  and ginst283 (i_10581, i_10273, i_10360, i_9543);
  and ginst284 (i_10582, i_10273, i_10357, i_9905);
  not ginst285 (i_10583, i_10367);
  and ginst286 (i_10587, i_10367, i_5735);
  and ginst287 (i_10588, i_10367, i_3135);
  not ginst288 (i_10589, i_10375);
  and ginst289 (i_10594, i_10381, i_7149, i_7159, i_7170, i_7180);
  and ginst290 (i_10595, i_10381, i_7159, i_7170, i_7180);
  and ginst291 (i_10596, i_10381, i_7170, i_7180);
  and ginst292 (i_10597, i_10381, i_7180);
  and ginst293 (i_10598, i_10381, i_8444);
  not ginst294 (i_10602, i_10381);
  nand ginst295 (i_10609, i_10515, i_7479);
  nand ginst296 (i_10610, i_10517, i_7491);
  nand ginst297 (i_10621, i_10534, i_9149);
  nand ginst298 (i_10626, i_10542, i_9206);
  nand ginst299 (i_10627, i_10544, i_9223);
  or ginst300 (i_10628, i_10451, i_10546);
  and ginst301 (i_10629, i_10547, i_9733);
  and ginst302 (i_10631, i_10550, i_5166);
  nand ginst303 (i_10632, i_10456, i_10552);
  nand ginst304 (i_10637, i_10557, i_7414);
  nand ginst305 (i_10638, i_10559, i_7417);
  nand ginst306 (i_10639, i_10561, i_7420);
  nand ginst307 (i_10640, i_10563, i_7423);
  nand ginst308 (i_10641, i_10466, i_10565);
  nand ginst309 (i_10642, i_10566, i_7429);
  nand ginst310 (i_10643, i_10568, i_7432);
  nand ginst311 (i_10644, i_10570, i_7435);
  nand ginst312 (i_10645, i_10572, i_7438);
  and ginst313 (i_10647, i_10577, i_886, i_887);
  and ginst314 (i_10648, i_10360, i_10479, i_8857);
  and ginst315 (i_10649, i_10357, i_10479, i_7609);
  or ginst316 (i_10652, i_10598, i_8966);
  or ginst317 (i_10659, i_10594, i_4675, i_8451, i_8452, i_8453);
  or ginst318 (i_10662, i_10595, i_4678, i_8454, i_8455);
  or ginst319 (i_10665, i_10596, i_4682, i_8456);
  or ginst320 (i_10668, i_10597, i_4687);
  not ginst321 (i_10671, i_10509);
  nand ginst322 (i_10672, i_10509, i_8615);
  not ginst323 (i_10673, i_10512);
  nand ginst324 (i_10674, i_10512, i_8624);
  nand ginst325 (i_10675, i_10516, i_10609);
  nand ginst326 (i_10678, i_10518, i_10610);
  not ginst327 (i_10681, i_10519);
  nand ginst328 (i_10682, i_10519, i_8644);
  not ginst329 (i_10683, i_10522);
  nand ginst330 (i_10684, i_10522, i_8653);
  not ginst331 (i_10685, i_10525);
  nand ginst332 (i_10686, i_10525, i_9454);
  not ginst333 (i_10687, i_10528);
  nand ginst334 (i_10688, i_10528, i_9459);
  not ginst335 (i_10689, i_10531);
  nand ginst336 (i_10690, i_10531, i_9978);
  nand ginst337 (i_10691, i_10535, i_10621);
  not ginst338 (i_10694, i_10536);
  nand ginst339 (i_10695, i_10536, i_9493);
  not ginst340 (i_10696, i_10539);
  nand ginst341 (i_10697, i_10539, i_9498);
  nand ginst342 (i_10698, i_10543, i_10626);
  nand ginst343 (i_10701, i_10545, i_10627);
  or ginst344 (i_10704, i_10548, i_10629);
  and ginst345 (i_10705, i_10583, i_3159);
  or ginst346 (i_10706, i_10551, i_10631);
  and ginst347 (i_10707, i_10589, i_9737);
  and ginst348 (i_10708, i_10589, i_9738);
  and ginst349 (i_10709, i_10589, i_9243);
  and ginst350 (i_10710, i_10589, i_5892);
  nand ginst351 (i_10711, i_10558, i_10637);
  nand ginst352 (i_10712, i_10560, i_10638);
  nand ginst353 (i_10713, i_10562, i_10639);
  nand ginst354 (i_10714, i_10564, i_10640);
  nand ginst355 (i_10715, i_10567, i_10642);
  nand ginst356 (i_10716, i_10569, i_10643);
  nand ginst357 (i_10717, i_10571, i_10644);
  nand ginst358 (i_10718, i_10573, i_10645);
  not ginst359 (i_10719, i_10602);
  nand ginst360 (i_10720, i_10602, i_9244);
  not ginst361 (i_10729, i_10647);
  and ginst362 (i_10730, i_10583, i_5178);
  and ginst363 (i_10731, i_10583, i_2533);
  nand ginst364 (i_10737, i_10671, i_7447);
  nand ginst365 (i_10738, i_10673, i_7465);
  or ginst366 (i_10739, i_10581, i_10582, i_10648, i_10649);
  nand ginst367 (i_10746, i_10681, i_7503);
  nand ginst368 (i_10747, i_10683, i_7521);
  nand ginst369 (i_10748, i_10685, i_8678);
  nand ginst370 (i_10749, i_10687, i_8690);
  nand ginst371 (i_10750, i_10689, i_9685);
  nand ginst372 (i_10753, i_10694, i_8757);
  nand ginst373 (i_10754, i_10696, i_8769);
  or ginst374 (i_10759, i_10549, i_10705);
  or ginst375 (i_10760, i_10553, i_10707);
  or ginst376 (i_10761, i_10554, i_10708);
  or ginst377 (i_10762, i_10555, i_10709);
  or ginst378 (i_10763, i_10556, i_10710);
  nand ginst379 (i_10764, i_10719, i_8580);
  and ginst380 (i_10765, i_10652, i_9890);
  and ginst381 (i_10766, i_10652, i_9891);
  and ginst382 (i_10767, i_10652, i_9892);
  and ginst383 (i_10768, i_10652, i_8252);
  not ginst384 (i_10769, i_10659);
  nand ginst385 (i_10770, i_10659, i_9245);
  not ginst386 (i_10771, i_10662);
  nand ginst387 (i_10772, i_10662, i_9246);
  not ginst388 (i_10773, i_10665);
  nand ginst389 (i_10774, i_10665, i_9247);
  not ginst390 (i_10775, i_10668);
  nand ginst391 (i_10776, i_10668, i_9248);
  or ginst392 (i_10778, i_10587, i_10730);
  or ginst393 (i_10781, i_10588, i_10731);
  not ginst394 (i_10784, i_10652);
  nand ginst395 (i_10789, i_10672, i_10737);
  nand ginst396 (i_10792, i_10674, i_10738);
  not ginst397 (i_10796, i_10675);
  nand ginst398 (i_10797, i_10675, i_8633);
  not ginst399 (i_10798, i_10678);
  nand ginst400 (i_10799, i_10678, i_8638);
  nand ginst401 (i_10800, i_10682, i_10746);
  nand ginst402 (i_10803, i_10684, i_10747);
  nand ginst403 (i_10806, i_10686, i_10748);
  nand ginst404 (i_10809, i_10688, i_10749);
  nand ginst405 (i_10812, i_10690, i_10750);
  not ginst406 (i_10815, i_10691);
  nand ginst407 (i_10816, i_10691, i_9866);
  nand ginst408 (i_10817, i_10695, i_10753);
  nand ginst409 (i_10820, i_10697, i_10754);
  not ginst410 (i_10823, i_10698);
  nand ginst411 (i_10824, i_10698, i_9505);
  not ginst412 (i_10825, i_10701);
  nand ginst413 (i_10826, i_10701, i_9514);
  nand ginst414 (i_10827, i_10720, i_10764);
  nand ginst415 (i_10832, i_10769, i_8583);
  nand ginst416 (i_10833, i_10771, i_8586);
  nand ginst417 (i_10834, i_10773, i_8589);
  nand ginst418 (i_10835, i_10775, i_8592);
  not ginst419 (i_10836, i_10739);
  not ginst420 (i_10837, i_10778);
  not ginst421 (i_10838, i_10778);
  not ginst422 (i_10839, i_10781);
  not ginst423 (i_10840, i_10781);
  nand ginst424 (i_10845, i_10796, i_7482);
  nand ginst425 (i_10846, i_10798, i_7494);
  nand ginst426 (i_10857, i_10815, i_9473);
  nand ginst427 (i_10862, i_10823, i_8781);
  nand ginst428 (i_10863, i_10825, i_8799);
  and ginst429 (i_10864, i_10023, i_10784);
  and ginst430 (i_10865, i_10024, i_10784);
  and ginst431 (i_10866, i_10784, i_9739);
  and ginst432 (i_10867, i_10784, i_7136);
  nand ginst433 (i_10868, i_10770, i_10832);
  nand ginst434 (i_10869, i_10772, i_10833);
  nand ginst435 (i_10870, i_10774, i_10834);
  nand ginst436 (i_10871, i_10776, i_10835);
  not ginst437 (i_10872, i_10789);
  nand ginst438 (i_10873, i_10789, i_8616);
  not ginst439 (i_10874, i_10792);
  nand ginst440 (i_10875, i_10792, i_8625);
  nand ginst441 (i_10876, i_10797, i_10845);
  nand ginst442 (i_10879, i_10799, i_10846);
  not ginst443 (i_10882, i_10800);
  nand ginst444 (i_10883, i_10800, i_8645);
  not ginst445 (i_10884, i_10803);
  nand ginst446 (i_10885, i_10803, i_8654);
  not ginst447 (i_10886, i_10806);
  nand ginst448 (i_10887, i_10806, i_9455);
  not ginst449 (i_10888, i_10809);
  nand ginst450 (i_10889, i_10809, i_9460);
  not ginst451 (i_10890, i_10812);
  nand ginst452 (i_10891, i_10812, i_9862);
  nand ginst453 (i_10892, i_10816, i_10857);
  not ginst454 (i_10895, i_10817);
  nand ginst455 (i_10896, i_10817, i_9494);
  not ginst456 (i_10897, i_10820);
  nand ginst457 (i_10898, i_10820, i_9499);
  nand ginst458 (i_10899, i_10824, i_10862);
  nand ginst459 (i_10902, i_10826, i_10863);
  or ginst460 (i_10905, i_10765, i_10864);
  or ginst461 (i_10906, i_10766, i_10865);
  or ginst462 (i_10907, i_10767, i_10866);
  or ginst463 (i_10908, i_10768, i_10867);
  nand ginst464 (i_10909, i_10872, i_7450);
  nand ginst465 (i_10910, i_10874, i_7468);
  nand ginst466 (i_10915, i_10882, i_7506);
  nand ginst467 (i_10916, i_10884, i_7524);
  nand ginst468 (i_10917, i_10886, i_8681);
  nand ginst469 (i_10918, i_10888, i_8693);
  nand ginst470 (i_10919, i_10890, i_9462);
  nand ginst471 (i_10922, i_10895, i_8760);
  nand ginst472 (i_10923, i_10897, i_8772);
  nand ginst473 (i_10928, i_10873, i_10909);
  nand ginst474 (i_10931, i_10875, i_10910);
  not ginst475 (i_10934, i_10876);
  nand ginst476 (i_10935, i_10876, i_8634);
  not ginst477 (i_10936, i_10879);
  nand ginst478 (i_10937, i_10879, i_8639);
  nand ginst479 (i_10938, i_10883, i_10915);
  nand ginst480 (i_10941, i_10885, i_10916);
  nand ginst481 (i_10944, i_10887, i_10917);
  nand ginst482 (i_10947, i_10889, i_10918);
  nand ginst483 (i_10950, i_10891, i_10919);
  not ginst484 (i_10953, i_10892);
  nand ginst485 (i_10954, i_10892, i_9476);
  nand ginst486 (i_10955, i_10896, i_10922);
  nand ginst487 (i_10958, i_10898, i_10923);
  not ginst488 (i_10961, i_10899);
  nand ginst489 (i_10962, i_10899, i_9506);
  not ginst490 (i_10963, i_10902);
  nand ginst491 (i_10964, i_10902, i_9515);
  nand ginst492 (i_10969, i_10934, i_7485);
  nand ginst493 (i_10970, i_10936, i_7497);
  nand ginst494 (i_10981, i_10953, i_8718);
  nand ginst495 (i_10986, i_10961, i_8784);
  nand ginst496 (i_10987, i_10963, i_8802);
  not ginst497 (i_10988, i_10928);
  nand ginst498 (i_10989, i_10928, i_8617);
  not ginst499 (i_10990, i_10931);
  nand ginst500 (i_10991, i_10931, i_8626);
  nand ginst501 (i_10992, i_10935, i_10969);
  nand ginst502 (i_10995, i_10937, i_10970);
  not ginst503 (i_10998, i_10938);
  nand ginst504 (i_10999, i_10938, i_8646);
  not ginst505 (i_11000, i_10941);
  nand ginst506 (i_11001, i_10941, i_8655);
  not ginst507 (i_11002, i_10944);
  nand ginst508 (i_11003, i_10944, i_9456);
  not ginst509 (i_11004, i_10947);
  nand ginst510 (i_11005, i_10947, i_9461);
  not ginst511 (i_11006, i_10950);
  nand ginst512 (i_11007, i_10950, i_9465);
  nand ginst513 (i_11008, i_10954, i_10981);
  not ginst514 (i_11011, i_10955);
  nand ginst515 (i_11012, i_10955, i_9495);
  not ginst516 (i_11013, i_10958);
  nand ginst517 (i_11014, i_10958, i_9500);
  nand ginst518 (i_11015, i_10962, i_10986);
  nand ginst519 (i_11018, i_10964, i_10987);
  nand ginst520 (i_11023, i_10988, i_7453);
  nand ginst521 (i_11024, i_10990, i_7471);
  nand ginst522 (i_11027, i_10998, i_7509);
  nand ginst523 (i_11028, i_11000, i_7527);
  nand ginst524 (i_11029, i_11002, i_8684);
  nand ginst525 (i_11030, i_11004, i_8696);
  nand ginst526 (i_11031, i_11006, i_8702);
  nand ginst527 (i_11034, i_11011, i_8763);
  nand ginst528 (i_11035, i_11013, i_8775);
  not ginst529 (i_11040, i_10992);
  nand ginst530 (i_11041, i_10992, i_8294);
  not ginst531 (i_11042, i_10995);
  nand ginst532 (i_11043, i_10995, i_8295);
  nand ginst533 (i_11044, i_10989, i_11023);
  nand ginst534 (i_11047, i_10991, i_11024);
  nand ginst535 (i_11050, i_10999, i_11027);
  nand ginst536 (i_11053, i_11001, i_11028);
  nand ginst537 (i_11056, i_11003, i_11029);
  nand ginst538 (i_11059, i_11005, i_11030);
  nand ginst539 (i_11062, i_11007, i_11031);
  not ginst540 (i_11065, i_11008);
  nand ginst541 (i_11066, i_11008, i_9477);
  nand ginst542 (i_11067, i_11012, i_11034);
  nand ginst543 (i_11070, i_11014, i_11035);
  not ginst544 (i_11073, i_11015);
  nand ginst545 (i_11074, i_11015, i_9507);
  not ginst546 (i_11075, i_11018);
  nand ginst547 (i_11076, i_11018, i_9516);
  nand ginst548 (i_11077, i_11040, i_7488);
  nand ginst549 (i_11078, i_11042, i_7500);
  and ginst550 (i_1109, i_469, i_596);
  nand ginst551 (i_11095, i_11065, i_8721);
  nand ginst552 (i_11098, i_11073, i_8787);
  nand ginst553 (i_11099, i_11075, i_8805);
  nand ginst554 (i_1110, i_242, i_593);
  nand ginst555 (i_11100, i_11041, i_11077);
  nand ginst556 (i_11103, i_11043, i_11078);
  not ginst557 (i_11106, i_11056);
  nand ginst558 (i_11107, i_11056, i_9319);
  not ginst559 (i_11108, i_11059);
  nand ginst560 (i_11109, i_11059, i_9320);
  not ginst561 (i_1111, i_625);
  not ginst562 (i_11110, i_11067);
  nand ginst563 (i_11111, i_11067, i_9381);
  not ginst564 (i_11112, i_11070);
  nand ginst565 (i_11113, i_11070, i_9382);
  not ginst566 (i_11114, i_11044);
  nand ginst567 (i_11115, i_11044, i_8618);
  not ginst568 (i_11116, i_11047);
  nand ginst569 (i_11117, i_11047, i_8619);
  not ginst570 (i_11118, i_11050);
  nand ginst571 (i_11119, i_11050, i_8647);
  nand ginst572 (i_1112, i_242, i_593);
  not ginst573 (i_11120, i_11053);
  nand ginst574 (i_11121, i_11053, i_8648);
  not ginst575 (i_11122, i_11062);
  nand ginst576 (i_11123, i_11062, i_9466);
  nand ginst577 (i_11124, i_11066, i_11095);
  nand ginst578 (i_11127, i_11074, i_11098);
  nand ginst579 (i_1113, i_469, i_596);
  nand ginst580 (i_11130, i_11076, i_11099);
  nand ginst581 (i_11137, i_11106, i_8687);
  nand ginst582 (i_11138, i_11108, i_8699);
  nand ginst583 (i_11139, i_11110, i_8766);
  not ginst584 (i_1114, i_625);
  nand ginst585 (i_11140, i_11112, i_8778);
  nand ginst586 (i_11141, i_11114, i_7456);
  nand ginst587 (i_11142, i_11116, i_7474);
  nand ginst588 (i_11143, i_11118, i_7512);
  nand ginst589 (i_11144, i_11120, i_7530);
  nand ginst590 (i_11145, i_11122, i_8705);
  not ginst591 (i_1115, i_871);
  and ginst592 (i_11152, i_10283, i_11103, i_8871);
  and ginst593 (i_11153, i_10283, i_11100, i_7655);
  and ginst594 (i_11154, i_10119, i_11103, i_9551);
  and ginst595 (i_11155, i_10119, i_11100, i_9917);
  nand ginst596 (i_11156, i_11107, i_11137);
  nand ginst597 (i_11159, i_11109, i_11138);
  not ginst598 (i_1116, i_590);
  nand ginst599 (i_11162, i_11111, i_11139);
  nand ginst600 (i_11165, i_11113, i_11140);
  nand ginst601 (i_11168, i_11115, i_11141);
  nand ginst602 (i_11171, i_11117, i_11142);
  nand ginst603 (i_11174, i_11119, i_11143);
  nand ginst604 (i_11177, i_11121, i_11144);
  nand ginst605 (i_11180, i_11123, i_11145);
  not ginst606 (i_11183, i_11124);
  nand ginst607 (i_11184, i_11124, i_9468);
  not ginst608 (i_11185, i_11127);
  nand ginst609 (i_11186, i_11127, i_9508);
  not ginst610 (i_11187, i_11130);
  nand ginst611 (i_11188, i_11130, i_9509);
  not ginst612 (i_1119, i_628);
  or ginst613 (i_11205, i_11152, i_11153, i_11154, i_11155);
  nand ginst614 (i_11210, i_11183, i_8724);
  nand ginst615 (i_11211, i_11185, i_8790);
  nand ginst616 (i_11212, i_11187, i_8808);
  not ginst617 (i_11213, i_11168);
  nand ginst618 (i_11214, i_11168, i_8260);
  not ginst619 (i_11215, i_11171);
  nand ginst620 (i_11216, i_11171, i_8261);
  not ginst621 (i_11217, i_11174);
  nand ginst622 (i_11218, i_11174, i_8296);
  not ginst623 (i_11219, i_11177);
  nand ginst624 (i_11220, i_11177, i_8297);
  and ginst625 (i_11222, i_11159, i_1218, i_9575);
  and ginst626 (i_11223, i_11156, i_1218, i_8927);
  and ginst627 (i_11224, i_11159, i_750, i_9935);
  and ginst628 (i_11225, i_10132, i_11156, i_750);
  and ginst629 (i_11226, i_10497, i_11165, i_9608);
  and ginst630 (i_11227, i_10497, i_11162, i_9001);
  and ginst631 (i_11228, i_10301, i_11165, i_9949);
  and ginst632 (i_11229, i_10160, i_10301, i_11162);
  not ginst633 (i_11231, i_11180);
  nand ginst634 (i_11232, i_11180, i_9467);
  nand ginst635 (i_11233, i_11184, i_11210);
  nand ginst636 (i_11236, i_11186, i_11211);
  nand ginst637 (i_11239, i_11188, i_11212);
  nand ginst638 (i_11242, i_11213, i_7459);
  nand ginst639 (i_11243, i_11215, i_7462);
  nand ginst640 (i_11244, i_11217, i_7515);
  nand ginst641 (i_11245, i_11219, i_7518);
  not ginst642 (i_11246, i_11205);
  not ginst643 (i_1125, i_682);
  nand ginst644 (i_11250, i_11231, i_8708);
  or ginst645 (i_11252, i_11222, i_11223, i_11224, i_11225);
  or ginst646 (i_11257, i_11226, i_11227, i_11228, i_11229);
  nand ginst647 (i_11260, i_11214, i_11242);
  nand ginst648 (i_11261, i_11216, i_11243);
  nand ginst649 (i_11262, i_11218, i_11244);
  nand ginst650 (i_11263, i_11220, i_11245);
  not ginst651 (i_11264, i_11233);
  nand ginst652 (i_11265, i_11233, i_9322);
  not ginst653 (i_11267, i_11236);
  nand ginst654 (i_11268, i_11236, i_9383);
  not ginst655 (i_11269, i_11239);
  nand ginst656 (i_11270, i_11239, i_9384);
  nand ginst657 (i_11272, i_11232, i_11250);
  not ginst658 (i_11277, i_11261);
  and ginst659 (i_11278, i_10273, i_11260);
  not ginst660 (i_11279, i_11263);
  and ginst661 (i_11280, i_10119, i_11262);
  nand ginst662 (i_11282, i_11264, i_8714);
  not ginst663 (i_11283, i_11252);
  nand ginst664 (i_11284, i_11267, i_8793);
  nand ginst665 (i_11285, i_11269, i_8796);
  not ginst666 (i_11286, i_11257);
  and ginst667 (i_11288, i_10479, i_11277);
  and ginst668 (i_11289, i_10283, i_11279);
  not ginst669 (i_11290, i_11272);
  nand ginst670 (i_11291, i_11272, i_9321);
  nand ginst671 (i_11292, i_11265, i_11282);
  nand ginst672 (i_11293, i_11268, i_11284);
  nand ginst673 (i_11294, i_11270, i_11285);
  nand ginst674 (i_11295, i_11290, i_8711);
  not ginst675 (i_11296, i_11292);
  not ginst676 (i_11297, i_11294);
  and ginst677 (i_11298, i_10301, i_11293);
  or ginst678 (i_11299, i_11278, i_11288);
  or ginst679 (i_11302, i_11280, i_11289);
  nand ginst680 (i_11307, i_11291, i_11295);
  and ginst681 (i_11308, i_11296, i_1218);
  and ginst682 (i_11309, i_10497, i_11297);
  nand ginst683 (i_11312, i_11246, i_11302);
  nand ginst684 (i_11313, i_10836, i_11299);
  not ginst685 (i_11314, i_11299);
  not ginst686 (i_11315, i_11302);
  and ginst687 (i_11316, i_11307, i_750);
  or ginst688 (i_11317, i_11298, i_11309);
  not ginst689 (i_1132, i_628);
  nand ginst690 (i_11320, i_11205, i_11315);
  nand ginst691 (i_11321, i_10739, i_11314);
  or ginst692 (i_11323, i_11308, i_11316);
  nand ginst693 (i_11327, i_11312, i_11320);
  nand ginst694 (i_11328, i_11313, i_11321);
  nand ginst695 (i_11329, i_11286, i_11317);
  not ginst696 (i_11331, i_11317);
  not ginst697 (i_11333, i_11327);
  not ginst698 (i_11334, i_11328);
  nand ginst699 (i_11335, i_11257, i_11331);
  nand ginst700 (i_11336, i_11283, i_11323);
  not ginst701 (i_11337, i_11323);
  nand ginst702 (i_11338, i_11329, i_11335);
  nand ginst703 (i_11339, i_11252, i_11337);
  not ginst704 (i_11340, i_11338);
  nand ginst705 (i_11341, i_11336, i_11339);
  not ginst706 (i_11342, i_11341);
  not ginst707 (i_1136, i_682);
  not ginst708 (i_1141, i_628);
  not ginst709 (i_1147, i_682);
  not ginst710 (i_1154, i_632);
  not ginst711 (i_1160, i_676);
  and ginst712 (i_1167, i_614, i_700);
  and ginst713 (i_1174, i_614, i_700);
  not ginst714 (i_1175, i_682);
  not ginst715 (i_1182, i_676);
  not ginst716 (i_1189, i_657);
  not ginst717 (i_1194, i_676);
  not ginst718 (i_1199, i_682);
  not ginst719 (i_1206, i_689);
  not ginst720 (i_1211, i_695);
  not ginst721 (i_1218, i_750);
  not ginst722 (i_1222, i_1028);
  not ginst723 (i_1227, i_632);
  not ginst724 (i_1233, i_676);
  not ginst725 (i_1240, i_632);
  not ginst726 (i_1244, i_676);
  not ginst727 (i_1249, i_689);
  not ginst728 (i_1256, i_689);
  not ginst729 (i_1263, i_695);
  not ginst730 (i_1270, i_689);
  not ginst731 (i_1277, i_689);
  not ginst732 (i_1284, i_700);
  not ginst733 (i_1287, i_614);
  not ginst734 (i_1290, i_666);
  not ginst735 (i_1293, i_660);
  not ginst736 (i_1296, i_651);
  not ginst737 (i_1299, i_614);
  not ginst738 (i_1302, i_644);
  not ginst739 (i_1305, i_700);
  not ginst740 (i_1308, i_614);
  not ginst741 (i_1311, i_614);
  not ginst742 (i_1314, i_666);
  not ginst743 (i_1317, i_660);
  not ginst744 (i_1320, i_651);
  not ginst745 (i_1323, i_644);
  not ginst746 (i_1326, i_609);
  not ginst747 (i_1329, i_604);
  not ginst748 (i_1332, i_742);
  not ginst749 (i_1335, i_599);
  not ginst750 (i_1338, i_727);
  not ginst751 (i_1341, i_721);
  not ginst752 (i_1344, i_715);
  not ginst753 (i_1347, i_734);
  not ginst754 (i_1350, i_708);
  not ginst755 (i_1353, i_609);
  not ginst756 (i_1356, i_604);
  not ginst757 (i_1359, i_742);
  not ginst758 (i_1362, i_734);
  not ginst759 (i_1365, i_599);
  not ginst760 (i_1368, i_727);
  not ginst761 (i_1371, i_721);
  not ginst762 (i_1374, i_715);
  not ginst763 (i_1377, i_708);
  not ginst764 (i_1380, i_806);
  not ginst765 (i_1383, i_800);
  not ginst766 (i_1386, i_794);
  not ginst767 (i_1389, i_786);
  not ginst768 (i_1392, i_780);
  not ginst769 (i_1395, i_774);
  not ginst770 (i_1398, i_768);
  not ginst771 (i_1401, i_762);
  not ginst772 (i_1404, i_806);
  not ginst773 (i_1407, i_800);
  not ginst774 (i_1410, i_794);
  not ginst775 (i_1413, i_780);
  not ginst776 (i_1416, i_774);
  not ginst777 (i_1419, i_768);
  not ginst778 (i_1422, i_762);
  not ginst779 (i_1425, i_786);
  not ginst780 (i_1428, i_636);
  not ginst781 (i_1431, i_636);
  not ginst782 (i_1434, i_865);
  not ginst783 (i_1437, i_859);
  not ginst784 (i_1440, i_853);
  not ginst785 (i_1443, i_845);
  not ginst786 (i_1446, i_839);
  not ginst787 (i_1449, i_833);
  not ginst788 (i_1452, i_827);
  not ginst789 (i_1455, i_821);
  not ginst790 (i_1458, i_814);
  not ginst791 (i_1461, i_865);
  not ginst792 (i_1464, i_859);
  not ginst793 (i_1467, i_853);
  not ginst794 (i_1470, i_839);
  not ginst795 (i_1473, i_833);
  not ginst796 (i_1476, i_827);
  not ginst797 (i_1479, i_821);
  not ginst798 (i_1482, i_845);
  not ginst799 (i_1485, i_814);
  not ginst800 (i_1489, i_1109);
  not ginst801 (i_1490, i_1116);
  and ginst802 (i_1537, i_614, i_957);
  and ginst803 (i_1551, i_614, i_957);
  and ginst804 (i_1649, i_1029, i_636);
  not ginst805 (i_1703, i_957);
  nor ginst806 (i_1708, i_614, i_957);
  not ginst807 (i_1713, i_957);
  nor ginst808 (i_1721, i_614, i_957);
  not ginst809 (i_1758, i_1029);
  and ginst810 (i_1781, i_163, i_1116);
  and ginst811 (i_1782, i_170, i_1125);
  not ginst812 (i_1783, i_1125);
  not ginst813 (i_1789, i_1136);
  and ginst814 (i_1793, i_169, i_1125);
  and ginst815 (i_1794, i_168, i_1125);
  and ginst816 (i_1795, i_167, i_1125);
  and ginst817 (i_1796, i_166, i_1136);
  and ginst818 (i_1797, i_165, i_1136);
  and ginst819 (i_1798, i_164, i_1136);
  not ginst820 (i_1799, i_1147);
  not ginst821 (i_1805, i_1160);
  and ginst822 (i_1811, i_177, i_1147);
  and ginst823 (i_1812, i_176, i_1147);
  and ginst824 (i_1813, i_175, i_1147);
  and ginst825 (i_1814, i_174, i_1147);
  and ginst826 (i_1815, i_173, i_1147);
  and ginst827 (i_1816, i_157, i_1160);
  and ginst828 (i_1817, i_156, i_1160);
  and ginst829 (i_1818, i_155, i_1160);
  and ginst830 (i_1819, i_154, i_1160);
  and ginst831 (i_1820, i_153, i_1160);
  not ginst832 (i_1821, i_1284);
  not ginst833 (i_1822, i_1287);
  not ginst834 (i_1828, i_1290);
  not ginst835 (i_1829, i_1293);
  not ginst836 (i_1830, i_1296);
  not ginst837 (i_1832, i_1299);
  not ginst838 (i_1833, i_1302);
  not ginst839 (i_1834, i_1305);
  not ginst840 (i_1835, i_1308);
  not ginst841 (i_1839, i_1311);
  not ginst842 (i_1840, i_1314);
  not ginst843 (i_1841, i_1317);
  not ginst844 (i_1842, i_1320);
  not ginst845 (i_1843, i_1323);
  not ginst846 (i_1845, i_1175);
  not ginst847 (i_1851, i_1182);
  and ginst848 (i_1857, i_181, i_1175);
  and ginst849 (i_1858, i_171, i_1175);
  and ginst850 (i_1859, i_180, i_1175);
  and ginst851 (i_1860, i_179, i_1175);
  and ginst852 (i_1861, i_178, i_1175);
  and ginst853 (i_1862, i_161, i_1182);
  and ginst854 (i_1863, i_151, i_1182);
  and ginst855 (i_1864, i_160, i_1182);
  and ginst856 (i_1865, i_159, i_1182);
  and ginst857 (i_1866, i_158, i_1182);
  not ginst858 (i_1867, i_1326);
  not ginst859 (i_1868, i_1329);
  not ginst860 (i_1869, i_1332);
  not ginst861 (i_1870, i_1335);
  not ginst862 (i_1871, i_1338);
  not ginst863 (i_1872, i_1341);
  not ginst864 (i_1873, i_1344);
  not ginst865 (i_1874, i_1347);
  not ginst866 (i_1875, i_1350);
  not ginst867 (i_1876, i_1353);
  not ginst868 (i_1877, i_1356);
  not ginst869 (i_1878, i_1359);
  not ginst870 (i_1879, i_1362);
  not ginst871 (i_1880, i_1365);
  not ginst872 (i_1881, i_1368);
  not ginst873 (i_1882, i_1371);
  not ginst874 (i_1883, i_1374);
  not ginst875 (i_1884, i_1377);
  not ginst876 (i_1885, i_1199);
  not ginst877 (i_1892, i_1194);
  not ginst878 (i_1899, i_1199);
  not ginst879 (i_1906, i_1194);
  not ginst880 (i_1913, i_1211);
  not ginst881 (i_1919, i_1194);
  and ginst882 (i_1926, i_44, i_1211);
  and ginst883 (i_1927, i_41, i_1211);
  and ginst884 (i_1928, i_29, i_1211);
  and ginst885 (i_1929, i_26, i_1211);
  and ginst886 (i_1930, i_23, i_1211);
  not ginst887 (i_1931, i_1380);
  not ginst888 (i_1932, i_1383);
  not ginst889 (i_1933, i_1386);
  not ginst890 (i_1934, i_1389);
  not ginst891 (i_1935, i_1392);
  not ginst892 (i_1936, i_1395);
  not ginst893 (i_1937, i_1398);
  not ginst894 (i_1938, i_1401);
  not ginst895 (i_1939, i_1404);
  not ginst896 (i_1940, i_1407);
  not ginst897 (i_1941, i_1410);
  not ginst898 (i_1942, i_1413);
  not ginst899 (i_1943, i_1416);
  not ginst900 (i_1944, i_1419);
  not ginst901 (i_1945, i_1422);
  not ginst902 (i_1946, i_1425);
  not ginst903 (i_1947, i_1233);
  not ginst904 (i_1953, i_1244);
  and ginst905 (i_1957, i_209, i_1233);
  and ginst906 (i_1958, i_216, i_1233);
  and ginst907 (i_1959, i_215, i_1233);
  and ginst908 (i_1960, i_214, i_1233);
  and ginst909 (i_1961, i_213, i_1244);
  and ginst910 (i_1962, i_212, i_1244);
  and ginst911 (i_1963, i_211, i_1244);
  not ginst912 (i_1965, i_1428);
  and ginst913 (i_1966, i_1222, i_636);
  not ginst914 (i_1967, i_1431);
  not ginst915 (i_1968, i_1434);
  not ginst916 (i_1969, i_1437);
  not ginst917 (i_1970, i_1440);
  not ginst918 (i_1971, i_1443);
  not ginst919 (i_1972, i_1446);
  not ginst920 (i_1973, i_1449);
  not ginst921 (i_1974, i_1452);
  not ginst922 (i_1975, i_1455);
  not ginst923 (i_1976, i_1458);
  not ginst924 (i_1977, i_1249);
  not ginst925 (i_1983, i_1256);
  and ginst926 (i_1989, i_1249, i_642);
  and ginst927 (i_1990, i_1249, i_644);
  and ginst928 (i_1991, i_1249, i_651);
  and ginst929 (i_1992, i_1249, i_674);
  and ginst930 (i_1993, i_1249, i_660);
  and ginst931 (i_1994, i_1256, i_666);
  and ginst932 (i_1995, i_1256, i_672);
  and ginst933 (i_1996, i_1256, i_673);
  not ginst934 (i_1997, i_1263);
  not ginst935 (i_2003, i_1194);
  and ginst936 (i_2010, i_47, i_1263);
  and ginst937 (i_2011, i_35, i_1263);
  and ginst938 (i_2012, i_32, i_1263);
  and ginst939 (i_2013, i_50, i_1263);
  and ginst940 (i_2014, i_66, i_1263);
  not ginst941 (i_2015, i_1461);
  not ginst942 (i_2016, i_1464);
  not ginst943 (i_2017, i_1467);
  not ginst944 (i_2018, i_1470);
  not ginst945 (i_2019, i_1473);
  not ginst946 (i_2020, i_1476);
  not ginst947 (i_2021, i_1479);
  not ginst948 (i_2022, i_1482);
  not ginst949 (i_2023, i_1485);
  not ginst950 (i_2024, i_1206);
  not ginst951 (i_2031, i_1206);
  not ginst952 (i_2038, i_1206);
  not ginst953 (i_2045, i_1206);
  not ginst954 (i_2052, i_1270);
  not ginst955 (i_2058, i_1277);
  and ginst956 (i_2064, i_1270, i_706);
  and ginst957 (i_2065, i_1270, i_708);
  and ginst958 (i_2066, i_1270, i_715);
  and ginst959 (i_2067, i_1270, i_721);
  and ginst960 (i_2068, i_1270, i_727);
  and ginst961 (i_2069, i_1277, i_733);
  and ginst962 (i_2070, i_1277, i_734);
  and ginst963 (i_2071, i_1277, i_742);
  and ginst964 (i_2072, i_1277, i_748);
  and ginst965 (i_2073, i_1277, i_749);
  not ginst966 (i_2074, i_1189);
  not ginst967 (i_2081, i_1189);
  not ginst968 (i_2086, i_1222);
  nand ginst969 (i_2107, i_1287, i_1821);
  nand ginst970 (i_2108, i_1284, i_1822);
  not ginst971 (i_2110, i_1703);
  nand ginst972 (i_2111, i_1703, i_1832);
  nand ginst973 (i_2112, i_1308, i_1834);
  nand ginst974 (i_2113, i_1305, i_1835);
  not ginst975 (i_2114, i_1713);
  nand ginst976 (i_2115, i_1713, i_1839);
  not ginst977 (i_2117, i_1721);
  not ginst978 (i_2171, i_1758);
  nand ginst979 (i_2172, i_1758, i_1965);
  not ginst980 (i_2230, i_1708);
  not ginst981 (i_2231, i_1537);
  not ginst982 (i_2235, i_1551);
  or ginst983 (i_2239, i_1782, i_1783);
  or ginst984 (i_2240, i_1125, i_1783);
  or ginst985 (i_2241, i_1783, i_1793);
  or ginst986 (i_2242, i_1783, i_1794);
  or ginst987 (i_2243, i_1783, i_1795);
  or ginst988 (i_2244, i_1789, i_1796);
  or ginst989 (i_2245, i_1789, i_1797);
  or ginst990 (i_2246, i_1789, i_1798);
  or ginst991 (i_2247, i_1799, i_1811);
  or ginst992 (i_2248, i_1799, i_1812);
  or ginst993 (i_2249, i_1799, i_1813);
  or ginst994 (i_2250, i_1799, i_1814);
  or ginst995 (i_2251, i_1799, i_1815);
  or ginst996 (i_2252, i_1805, i_1816);
  or ginst997 (i_2253, i_1805, i_1817);
  or ginst998 (i_2254, i_1805, i_1818);
  or ginst999 (i_2255, i_1805, i_1819);
  or ginst1000 (i_2256, i_1805, i_1820);
  nand ginst1001 (i_2257, i_2107, i_2108);
  not ginst1002 (i_2267, i_2074);
  nand ginst1003 (i_2268, i_1299, i_2110);
  nand ginst1004 (i_2269, i_2112, i_2113);
  nand ginst1005 (i_2274, i_1311, i_2114);
  not ginst1006 (i_2275, i_2081);
  and ginst1007 (i_2277, i_141, i_1845);
  and ginst1008 (i_2278, i_147, i_1845);
  and ginst1009 (i_2279, i_138, i_1845);
  and ginst1010 (i_2280, i_144, i_1845);
  and ginst1011 (i_2281, i_135, i_1845);
  and ginst1012 (i_2282, i_141, i_1851);
  and ginst1013 (i_2283, i_147, i_1851);
  and ginst1014 (i_2284, i_138, i_1851);
  and ginst1015 (i_2285, i_144, i_1851);
  and ginst1016 (i_2286, i_135, i_1851);
  not ginst1017 (i_2287, i_1885);
  not ginst1018 (i_2293, i_1892);
  and ginst1019 (i_2299, i_103, i_1885);
  and ginst1020 (i_2300, i_130, i_1885);
  and ginst1021 (i_2301, i_127, i_1885);
  and ginst1022 (i_2302, i_124, i_1885);
  and ginst1023 (i_2303, i_100, i_1885);
  and ginst1024 (i_2304, i_103, i_1892);
  and ginst1025 (i_2305, i_130, i_1892);
  and ginst1026 (i_2306, i_127, i_1892);
  and ginst1027 (i_2307, i_124, i_1892);
  and ginst1028 (i_2308, i_100, i_1892);
  not ginst1029 (i_2309, i_1899);
  not ginst1030 (i_2315, i_1906);
  and ginst1031 (i_2321, i_115, i_1899);
  and ginst1032 (i_2322, i_118, i_1899);
  and ginst1033 (i_2323, i_97, i_1899);
  and ginst1034 (i_2324, i_94, i_1899);
  and ginst1035 (i_2325, i_121, i_1899);
  and ginst1036 (i_2326, i_115, i_1906);
  and ginst1037 (i_2327, i_118, i_1906);
  and ginst1038 (i_2328, i_97, i_1906);
  and ginst1039 (i_2329, i_94, i_1906);
  and ginst1040 (i_2330, i_121, i_1906);
  not ginst1041 (i_2331, i_1919);
  and ginst1042 (i_2337, i_208, i_1913);
  and ginst1043 (i_2338, i_198, i_1913);
  and ginst1044 (i_2339, i_207, i_1913);
  and ginst1045 (i_2340, i_206, i_1913);
  and ginst1046 (i_2341, i_205, i_1913);
  and ginst1047 (i_2342, i_44, i_1919);
  and ginst1048 (i_2343, i_41, i_1919);
  and ginst1049 (i_2344, i_29, i_1919);
  and ginst1050 (i_2345, i_26, i_1919);
  and ginst1051 (i_2346, i_23, i_1919);
  or ginst1052 (i_2347, i_1233, i_1947);
  or ginst1053 (i_2348, i_1947, i_1957);
  or ginst1054 (i_2349, i_1947, i_1958);
  or ginst1055 (i_2350, i_1947, i_1959);
  or ginst1056 (i_2351, i_1947, i_1960);
  or ginst1057 (i_2352, i_1953, i_1961);
  or ginst1058 (i_2353, i_1953, i_1962);
  or ginst1059 (i_2354, i_1953, i_1963);
  nand ginst1060 (i_2355, i_1428, i_2171);
  not ginst1061 (i_2356, i_2086);
  nand ginst1062 (i_2357, i_1967, i_2086);
  and ginst1063 (i_2358, i_114, i_1977);
  and ginst1064 (i_2359, i_113, i_1977);
  and ginst1065 (i_2360, i_111, i_1977);
  and ginst1066 (i_2361, i_87, i_1977);
  and ginst1067 (i_2362, i_112, i_1977);
  and ginst1068 (i_2363, i_88, i_1983);
  and ginst1069 (i_2364, i_245, i_1983);
  and ginst1070 (i_2365, i_271, i_1983);
  and ginst1071 (i_2366, i_1983, i_759);
  and ginst1072 (i_2367, i_70, i_1983);
  not ginst1073 (i_2368, i_2003);
  and ginst1074 (i_2374, i_193, i_1997);
  and ginst1075 (i_2375, i_192, i_1997);
  and ginst1076 (i_2376, i_191, i_1997);
  and ginst1077 (i_2377, i_190, i_1997);
  and ginst1078 (i_2378, i_189, i_1997);
  and ginst1079 (i_2379, i_47, i_2003);
  and ginst1080 (i_2380, i_35, i_2003);
  and ginst1081 (i_2381, i_32, i_2003);
  and ginst1082 (i_2382, i_50, i_2003);
  and ginst1083 (i_2383, i_66, i_2003);
  not ginst1084 (i_2384, i_2024);
  not ginst1085 (i_2390, i_2031);
  and ginst1086 (i_2396, i_58, i_2024);
  and ginst1087 (i_2397, i_77, i_2024);
  and ginst1088 (i_2398, i_78, i_2024);
  and ginst1089 (i_2399, i_59, i_2024);
  and ginst1090 (i_2400, i_81, i_2024);
  and ginst1091 (i_2401, i_80, i_2031);
  and ginst1092 (i_2402, i_79, i_2031);
  and ginst1093 (i_2403, i_60, i_2031);
  and ginst1094 (i_2404, i_61, i_2031);
  and ginst1095 (i_2405, i_62, i_2031);
  not ginst1096 (i_2406, i_2038);
  not ginst1097 (i_2412, i_2045);
  and ginst1098 (i_2418, i_69, i_2038);
  and ginst1099 (i_2419, i_70, i_2038);
  and ginst1100 (i_2420, i_74, i_2038);
  and ginst1101 (i_2421, i_76, i_2038);
  and ginst1102 (i_2422, i_75, i_2038);
  and ginst1103 (i_2423, i_73, i_2045);
  and ginst1104 (i_2424, i_53, i_2045);
  and ginst1105 (i_2425, i_54, i_2045);
  and ginst1106 (i_2426, i_55, i_2045);
  and ginst1107 (i_2427, i_56, i_2045);
  and ginst1108 (i_2428, i_82, i_2052);
  and ginst1109 (i_2429, i_65, i_2052);
  and ginst1110 (i_2430, i_83, i_2052);
  and ginst1111 (i_2431, i_84, i_2052);
  and ginst1112 (i_2432, i_85, i_2052);
  and ginst1113 (i_2433, i_64, i_2058);
  and ginst1114 (i_2434, i_63, i_2058);
  and ginst1115 (i_2435, i_86, i_2058);
  and ginst1116 (i_2436, i_109, i_2058);
  and ginst1117 (i_2437, i_110, i_2058);
  and ginst1118 (i_2441, i_1119, i_2239);
  and ginst1119 (i_2442, i_1119, i_2240);
  and ginst1120 (i_2446, i_1119, i_2241);
  and ginst1121 (i_2450, i_1119, i_2242);
  and ginst1122 (i_2454, i_1119, i_2243);
  and ginst1123 (i_2458, i_1132, i_2244);
  and ginst1124 (i_2462, i_1141, i_2247);
  and ginst1125 (i_2466, i_1141, i_2248);
  and ginst1126 (i_2470, i_1141, i_2249);
  and ginst1127 (i_2474, i_1141, i_2250);
  and ginst1128 (i_2478, i_1141, i_2251);
  and ginst1129 (i_2482, i_1154, i_2252);
  and ginst1130 (i_2488, i_1154, i_2253);
  and ginst1131 (i_2496, i_1154, i_2254);
  and ginst1132 (i_2502, i_1154, i_2255);
  and ginst1133 (i_2508, i_1154, i_2256);
  nand ginst1134 (i_2523, i_2111, i_2268);
  nand ginst1135 (i_2533, i_2115, i_2274);
  not ginst1136 (i_2537, i_2235);
  or ginst1137 (i_2538, i_1858, i_2278);
  or ginst1138 (i_2542, i_1859, i_2279);
  or ginst1139 (i_2546, i_1860, i_2280);
  or ginst1140 (i_2550, i_1861, i_2281);
  or ginst1141 (i_2554, i_1863, i_2283);
  or ginst1142 (i_2561, i_1864, i_2284);
  or ginst1143 (i_2567, i_1865, i_2285);
  or ginst1144 (i_2573, i_1866, i_2286);
  or ginst1145 (i_2604, i_1927, i_2338);
  or ginst1146 (i_2607, i_1928, i_2339);
  or ginst1147 (i_2611, i_1929, i_2340);
  or ginst1148 (i_2615, i_1930, i_2341);
  and ginst1149 (i_2619, i_1227, i_2348);
  and ginst1150 (i_2626, i_1227, i_2349);
  and ginst1151 (i_2632, i_1227, i_2350);
  and ginst1152 (i_2638, i_1227, i_2351);
  and ginst1153 (i_2644, i_1240, i_2352);
  nand ginst1154 (i_2650, i_2172, i_2355);
  nand ginst1155 (i_2653, i_1431, i_2356);
  or ginst1156 (i_2654, i_1990, i_2359);
  or ginst1157 (i_2658, i_1991, i_2360);
  or ginst1158 (i_2662, i_1992, i_2361);
  or ginst1159 (i_2666, i_1993, i_2362);
  or ginst1160 (i_2670, i_1994, i_2363);
  or ginst1161 (i_2674, i_1256, i_2366);
  or ginst1162 (i_2680, i_1256, i_2367);
  or ginst1163 (i_2688, i_2010, i_2374);
  or ginst1164 (i_2692, i_2011, i_2375);
  or ginst1165 (i_2696, i_2012, i_2376);
  or ginst1166 (i_2700, i_2013, i_2377);
  or ginst1167 (i_2704, i_2014, i_2378);
  and ginst1168 (i_2728, i_1227, i_2347);
  or ginst1169 (i_2729, i_2065, i_2429);
  or ginst1170 (i_2733, i_2066, i_2430);
  or ginst1171 (i_2737, i_2067, i_2431);
  or ginst1172 (i_2741, i_2068, i_2432);
  or ginst1173 (i_2745, i_2069, i_2433);
  or ginst1174 (i_2749, i_2070, i_2434);
  or ginst1175 (i_2753, i_2071, i_2435);
  or ginst1176 (i_2757, i_2072, i_2436);
  or ginst1177 (i_2761, i_2073, i_2437);
  not ginst1178 (i_2765, i_2231);
  and ginst1179 (i_2766, i_1240, i_2354);
  and ginst1180 (i_2769, i_1240, i_2353);
  and ginst1181 (i_2772, i_1132, i_2246);
  and ginst1182 (i_2775, i_1132, i_2245);
  or ginst1183 (i_2778, i_1862, i_2282);
  or ginst1184 (i_2781, i_1989, i_2358);
  or ginst1185 (i_2784, i_1996, i_2365);
  or ginst1186 (i_2787, i_1995, i_2364);
  or ginst1187 (i_2790, i_1926, i_2337);
  or ginst1188 (i_2793, i_1857, i_2277);
  or ginst1189 (i_2796, i_2064, i_2428);
  and ginst1190 (i_2866, i_1537, i_2257);
  and ginst1191 (i_2867, i_1537, i_2257);
  and ginst1192 (i_2868, i_1537, i_2257);
  and ginst1193 (i_2869, i_1537, i_2257);
  and ginst1194 (i_2878, i_1551, i_2269);
  and ginst1195 (i_2913, i_204, i_2287);
  and ginst1196 (i_2914, i_203, i_2287);
  and ginst1197 (i_2915, i_202, i_2287);
  and ginst1198 (i_2916, i_201, i_2287);
  and ginst1199 (i_2917, i_200, i_2287);
  and ginst1200 (i_2918, i_235, i_2293);
  and ginst1201 (i_2919, i_234, i_2293);
  and ginst1202 (i_2920, i_233, i_2293);
  and ginst1203 (i_2921, i_232, i_2293);
  and ginst1204 (i_2922, i_231, i_2293);
  and ginst1205 (i_2923, i_197, i_2309);
  and ginst1206 (i_2924, i_187, i_2309);
  and ginst1207 (i_2925, i_196, i_2309);
  and ginst1208 (i_2926, i_195, i_2309);
  and ginst1209 (i_2927, i_194, i_2309);
  and ginst1210 (i_2928, i_227, i_2315);
  and ginst1211 (i_2929, i_217, i_2315);
  and ginst1212 (i_2930, i_226, i_2315);
  and ginst1213 (i_2931, i_225, i_2315);
  and ginst1214 (i_2932, i_224, i_2315);
  and ginst1215 (i_2933, i_239, i_2331);
  and ginst1216 (i_2934, i_229, i_2331);
  and ginst1217 (i_2935, i_238, i_2331);
  and ginst1218 (i_2936, i_237, i_2331);
  and ginst1219 (i_2937, i_236, i_2331);
  nand ginst1220 (i_2988, i_2357, i_2653);
  and ginst1221 (i_3005, i_223, i_2368);
  and ginst1222 (i_3006, i_222, i_2368);
  and ginst1223 (i_3007, i_221, i_2368);
  and ginst1224 (i_3008, i_220, i_2368);
  and ginst1225 (i_3009, i_219, i_2368);
  and ginst1226 (i_3020, i_2384, i_812);
  and ginst1227 (i_3021, i_2384, i_814);
  and ginst1228 (i_3022, i_2384, i_821);
  and ginst1229 (i_3023, i_2384, i_827);
  and ginst1230 (i_3024, i_2384, i_833);
  and ginst1231 (i_3025, i_2390, i_839);
  and ginst1232 (i_3026, i_2390, i_845);
  and ginst1233 (i_3027, i_2390, i_853);
  and ginst1234 (i_3028, i_2390, i_859);
  and ginst1235 (i_3029, i_2390, i_865);
  and ginst1236 (i_3032, i_2406, i_758);
  and ginst1237 (i_3033, i_2406, i_759);
  and ginst1238 (i_3034, i_2406, i_762);
  and ginst1239 (i_3035, i_2406, i_768);
  and ginst1240 (i_3036, i_2406, i_774);
  and ginst1241 (i_3037, i_2412, i_780);
  and ginst1242 (i_3038, i_2412, i_786);
  and ginst1243 (i_3039, i_2412, i_794);
  and ginst1244 (i_3040, i_2412, i_800);
  and ginst1245 (i_3041, i_2412, i_806);
  not ginst1246 (i_3061, i_2257);
  not ginst1247 (i_3064, i_2257);
  not ginst1248 (i_3067, i_2269);
  not ginst1249 (i_3070, i_2269);
  not ginst1250 (i_3073, i_2728);
  not ginst1251 (i_3080, i_2441);
  and ginst1252 (i_3096, i_2644, i_666);
  and ginst1253 (i_3097, i_2638, i_660);
  and ginst1254 (i_3101, i_1189, i_2632);
  and ginst1255 (i_3107, i_2626, i_651);
  and ginst1256 (i_3114, i_2619, i_644);
  and ginst1257 (i_3122, i_2257, i_2523);
  or ginst1258 (i_3126, i_1167, i_2866);
  and ginst1259 (i_3130, i_2257, i_2523);
  or ginst1260 (i_3131, i_1167, i_2869);
  and ginst1261 (i_3134, i_2257, i_2523);
  not ginst1262 (i_3135, i_2533);
  and ginst1263 (i_3136, i_2644, i_666);
  and ginst1264 (i_3137, i_2638, i_660);
  and ginst1265 (i_3140, i_1189, i_2632);
  and ginst1266 (i_3144, i_2626, i_651);
  and ginst1267 (i_3149, i_2619, i_644);
  and ginst1268 (i_3155, i_2269, i_2533);
  or ginst1269 (i_3159, i_1174, i_2878);
  not ginst1270 (i_3167, i_2778);
  and ginst1271 (i_3168, i_2508, i_609);
  and ginst1272 (i_3169, i_2502, i_604);
  and ginst1273 (i_3173, i_2496, i_742);
  and ginst1274 (i_3178, i_2488, i_734);
  and ginst1275 (i_3184, i_2482, i_599);
  and ginst1276 (i_3185, i_2573, i_727);
  and ginst1277 (i_3189, i_2567, i_721);
  and ginst1278 (i_3195, i_2561, i_715);
  and ginst1279 (i_3202, i_2554, i_708);
  and ginst1280 (i_3210, i_2508, i_609);
  and ginst1281 (i_3211, i_2502, i_604);
  and ginst1282 (i_3215, i_2496, i_742);
  and ginst1283 (i_3221, i_2488, i_734);
  and ginst1284 (i_3228, i_2482, i_599);
  and ginst1285 (i_3229, i_2573, i_727);
  and ginst1286 (i_3232, i_2567, i_721);
  and ginst1287 (i_3236, i_2561, i_715);
  and ginst1288 (i_3241, i_2554, i_708);
  or ginst1289 (i_3247, i_2299, i_2913);
  or ginst1290 (i_3251, i_2300, i_2914);
  or ginst1291 (i_3255, i_2301, i_2915);
  or ginst1292 (i_3259, i_2302, i_2916);
  or ginst1293 (i_3263, i_2303, i_2917);
  or ginst1294 (i_3267, i_2304, i_2918);
  or ginst1295 (i_3273, i_2305, i_2919);
  or ginst1296 (i_3281, i_2306, i_2920);
  or ginst1297 (i_3287, i_2307, i_2921);
  or ginst1298 (i_3293, i_2308, i_2922);
  or ginst1299 (i_3299, i_2322, i_2924);
  or ginst1300 (i_3303, i_2323, i_2925);
  or ginst1301 (i_3307, i_2324, i_2926);
  or ginst1302 (i_3311, i_2325, i_2927);
  or ginst1303 (i_3315, i_2327, i_2929);
  or ginst1304 (i_3322, i_2328, i_2930);
  or ginst1305 (i_3328, i_2329, i_2931);
  or ginst1306 (i_3334, i_2330, i_2932);
  or ginst1307 (i_3340, i_2343, i_2934);
  or ginst1308 (i_3343, i_2344, i_2935);
  or ginst1309 (i_3349, i_2345, i_2936);
  or ginst1310 (i_3355, i_2346, i_2937);
  and ginst1311 (i_3361, i_2478, i_2761);
  and ginst1312 (i_3362, i_2474, i_2757);
  and ginst1313 (i_3363, i_2470, i_2753);
  and ginst1314 (i_3364, i_2466, i_2749);
  and ginst1315 (i_3365, i_2462, i_2745);
  and ginst1316 (i_3366, i_2550, i_2741);
  and ginst1317 (i_3367, i_2546, i_2737);
  and ginst1318 (i_3368, i_2542, i_2733);
  and ginst1319 (i_3369, i_2538, i_2729);
  and ginst1320 (i_3370, i_2458, i_2670);
  and ginst1321 (i_3371, i_2454, i_2666);
  and ginst1322 (i_3372, i_2450, i_2662);
  and ginst1323 (i_3373, i_2446, i_2658);
  and ginst1324 (i_3374, i_2442, i_2654);
  and ginst1325 (i_3375, i_2650, i_2988);
  and ginst1326 (i_3379, i_1966, i_2650);
  not ginst1327 (i_3380, i_2781);
  and ginst1328 (i_3381, i_2604, i_695);
  or ginst1329 (i_3384, i_2379, i_3005);
  or ginst1330 (i_3390, i_2380, i_3006);
  or ginst1331 (i_3398, i_2381, i_3007);
  or ginst1332 (i_3404, i_2382, i_3008);
  or ginst1333 (i_3410, i_2383, i_3009);
  or ginst1334 (i_3416, i_2397, i_3021);
  or ginst1335 (i_3420, i_2398, i_3022);
  or ginst1336 (i_3424, i_2399, i_3023);
  or ginst1337 (i_3428, i_2400, i_3024);
  or ginst1338 (i_3432, i_2401, i_3025);
  or ginst1339 (i_3436, i_2402, i_3026);
  or ginst1340 (i_3440, i_2403, i_3027);
  or ginst1341 (i_3444, i_2404, i_3028);
  or ginst1342 (i_3448, i_2405, i_3029);
  not ginst1343 (i_3452, i_2790);
  not ginst1344 (i_3453, i_2793);
  or ginst1345 (i_3454, i_2420, i_3034);
  or ginst1346 (i_3458, i_2421, i_3035);
  or ginst1347 (i_3462, i_2422, i_3036);
  or ginst1348 (i_3466, i_2423, i_3037);
  or ginst1349 (i_3470, i_2424, i_3038);
  or ginst1350 (i_3474, i_2425, i_3039);
  or ginst1351 (i_3478, i_2426, i_3040);
  or ginst1352 (i_3482, i_2427, i_3041);
  not ginst1353 (i_3486, i_2796);
  not ginst1354 (i_3487, i_2644);
  not ginst1355 (i_3490, i_2638);
  not ginst1356 (i_3493, i_2632);
  not ginst1357 (i_3496, i_2626);
  not ginst1358 (i_3499, i_2619);
  not ginst1359 (i_3502, i_2523);
  nor ginst1360 (i_3507, i_1167, i_2868);
  not ginst1361 (i_3510, i_2523);
  nor ginst1362 (i_3515, i_2619, i_644);
  not ginst1363 (i_3518, i_2644);
  not ginst1364 (i_3521, i_2638);
  not ginst1365 (i_3524, i_2632);
  not ginst1366 (i_3527, i_2626);
  not ginst1367 (i_3530, i_2619);
  not ginst1368 (i_3535, i_2619);
  not ginst1369 (i_3539, i_2632);
  not ginst1370 (i_3542, i_2626);
  not ginst1371 (i_3545, i_2644);
  not ginst1372 (i_3548, i_2638);
  not ginst1373 (i_3551, i_2766);
  not ginst1374 (i_3552, i_2769);
  not ginst1375 (i_3553, i_2442);
  not ginst1376 (i_3557, i_2450);
  not ginst1377 (i_3560, i_2446);
  not ginst1378 (i_3563, i_2458);
  not ginst1379 (i_3566, i_2454);
  not ginst1380 (i_3569, i_2772);
  not ginst1381 (i_3570, i_2775);
  not ginst1382 (i_3571, i_2554);
  not ginst1383 (i_3574, i_2567);
  not ginst1384 (i_3577, i_2561);
  not ginst1385 (i_3580, i_2482);
  not ginst1386 (i_3583, i_2573);
  not ginst1387 (i_3586, i_2496);
  not ginst1388 (i_3589, i_2488);
  not ginst1389 (i_3592, i_2508);
  not ginst1390 (i_3595, i_2502);
  not ginst1391 (i_3598, i_2508);
  not ginst1392 (i_3601, i_2502);
  not ginst1393 (i_3604, i_2496);
  not ginst1394 (i_3607, i_2482);
  not ginst1395 (i_3610, i_2573);
  not ginst1396 (i_3613, i_2567);
  not ginst1397 (i_3616, i_2561);
  not ginst1398 (i_3619, i_2488);
  not ginst1399 (i_3622, i_2554);
  nor ginst1400 (i_3625, i_2488, i_734);
  nor ginst1401 (i_3628, i_2554, i_708);
  not ginst1402 (i_3631, i_2508);
  not ginst1403 (i_3634, i_2502);
  not ginst1404 (i_3637, i_2496);
  not ginst1405 (i_3640, i_2488);
  not ginst1406 (i_3643, i_2482);
  not ginst1407 (i_3646, i_2573);
  not ginst1408 (i_3649, i_2567);
  not ginst1409 (i_3652, i_2561);
  not ginst1410 (i_3655, i_2554);
  nor ginst1411 (i_3658, i_2488, i_734);
  not ginst1412 (i_3661, i_2674);
  not ginst1413 (i_3664, i_2674);
  not ginst1414 (i_3667, i_2761);
  not ginst1415 (i_3670, i_2478);
  not ginst1416 (i_3673, i_2757);
  not ginst1417 (i_3676, i_2474);
  not ginst1418 (i_3679, i_2753);
  not ginst1419 (i_3682, i_2470);
  not ginst1420 (i_3685, i_2745);
  not ginst1421 (i_3688, i_2462);
  not ginst1422 (i_3691, i_2741);
  not ginst1423 (i_3694, i_2550);
  not ginst1424 (i_3697, i_2737);
  not ginst1425 (i_3700, i_2546);
  not ginst1426 (i_3703, i_2733);
  not ginst1427 (i_3706, i_2542);
  not ginst1428 (i_3709, i_2749);
  not ginst1429 (i_3712, i_2466);
  not ginst1430 (i_3715, i_2729);
  not ginst1431 (i_3718, i_2538);
  not ginst1432 (i_3721, i_2704);
  not ginst1433 (i_3724, i_2700);
  not ginst1434 (i_3727, i_2696);
  not ginst1435 (i_3730, i_2688);
  not ginst1436 (i_3733, i_2692);
  not ginst1437 (i_3736, i_2670);
  not ginst1438 (i_3739, i_2458);
  not ginst1439 (i_3742, i_2666);
  not ginst1440 (i_3745, i_2454);
  not ginst1441 (i_3748, i_2662);
  not ginst1442 (i_3751, i_2450);
  not ginst1443 (i_3754, i_2658);
  not ginst1444 (i_3757, i_2446);
  not ginst1445 (i_3760, i_2654);
  not ginst1446 (i_3763, i_2442);
  not ginst1447 (i_3766, i_2654);
  not ginst1448 (i_3769, i_2662);
  not ginst1449 (i_3772, i_2658);
  not ginst1450 (i_3775, i_2670);
  not ginst1451 (i_3778, i_2666);
  not ginst1452 (i_3781, i_2784);
  not ginst1453 (i_3782, i_2787);
  or ginst1454 (i_3783, i_2326, i_2928);
  or ginst1455 (i_3786, i_2342, i_2933);
  or ginst1456 (i_3789, i_2321, i_2923);
  not ginst1457 (i_3792, i_2688);
  not ginst1458 (i_3795, i_2696);
  not ginst1459 (i_3798, i_2692);
  not ginst1460 (i_3801, i_2704);
  not ginst1461 (i_3804, i_2700);
  not ginst1462 (i_3807, i_2604);
  not ginst1463 (i_3810, i_2611);
  not ginst1464 (i_3813, i_2607);
  not ginst1465 (i_3816, i_2615);
  not ginst1466 (i_3819, i_2538);
  not ginst1467 (i_3822, i_2546);
  not ginst1468 (i_3825, i_2542);
  not ginst1469 (i_3828, i_2462);
  not ginst1470 (i_3831, i_2550);
  not ginst1471 (i_3834, i_2470);
  not ginst1472 (i_3837, i_2466);
  not ginst1473 (i_3840, i_2478);
  not ginst1474 (i_3843, i_2474);
  not ginst1475 (i_3846, i_2615);
  not ginst1476 (i_3849, i_2611);
  not ginst1477 (i_3852, i_2607);
  not ginst1478 (i_3855, i_2680);
  not ginst1479 (i_3858, i_2729);
  not ginst1480 (i_3861, i_2737);
  not ginst1481 (i_3864, i_2733);
  not ginst1482 (i_3867, i_2745);
  not ginst1483 (i_387, i_1);
  not ginst1484 (i_3870, i_2741);
  not ginst1485 (i_3873, i_2753);
  not ginst1486 (i_3876, i_2749);
  not ginst1487 (i_3879, i_2761);
  not ginst1488 (i_388, i_1);
  not ginst1489 (i_3882, i_2757);
  or ginst1490 (i_3885, i_2419, i_3033);
  or ginst1491 (i_3888, i_2418, i_3032);
  or ginst1492 (i_3891, i_2396, i_3020);
  nand ginst1493 (i_3953, i_2117, i_3067);
  not ginst1494 (i_3954, i_3067);
  nand ginst1495 (i_3955, i_2537, i_3070);
  not ginst1496 (i_3956, i_3070);
  not ginst1497 (i_3958, i_3073);
  not ginst1498 (i_3964, i_3080);
  or ginst1499 (i_4193, i_1649, i_3379);
  or ginst1500 (i_4303, i_1167, i_2867, i_3130);
  not ginst1501 (i_4308, i_3061);
  not ginst1502 (i_4313, i_3064);
  nand ginst1503 (i_4326, i_2769, i_3551);
  nand ginst1504 (i_4327, i_2766, i_3552);
  nand ginst1505 (i_4333, i_2775, i_3569);
  nand ginst1506 (i_4334, i_2772, i_3570);
  nand ginst1507 (i_4411, i_2787, i_3781);
  nand ginst1508 (i_4412, i_2784, i_3782);
  nand ginst1509 (i_4463, i_1828, i_3487);
  not ginst1510 (i_4464, i_3487);
  nand ginst1511 (i_4465, i_1829, i_3490);
  not ginst1512 (i_4466, i_3490);
  nand ginst1513 (i_4467, i_2267, i_3493);
  not ginst1514 (i_4468, i_3493);
  nand ginst1515 (i_4469, i_1830, i_3496);
  not ginst1516 (i_4470, i_3496);
  nand ginst1517 (i_4471, i_1833, i_3499);
  not ginst1518 (i_4472, i_3499);
  not ginst1519 (i_4473, i_3122);
  not ginst1520 (i_4474, i_3126);
  nand ginst1521 (i_4475, i_1840, i_3518);
  not ginst1522 (i_4476, i_3518);
  nand ginst1523 (i_4477, i_1841, i_3521);
  not ginst1524 (i_4478, i_3521);
  nand ginst1525 (i_4479, i_2275, i_3524);
  not ginst1526 (i_4480, i_3524);
  nand ginst1527 (i_4481, i_1842, i_3527);
  not ginst1528 (i_4482, i_3527);
  nand ginst1529 (i_4483, i_1843, i_3530);
  not ginst1530 (i_4484, i_3530);
  not ginst1531 (i_4485, i_3155);
  not ginst1532 (i_4486, i_3159);
  nand ginst1533 (i_4487, i_1721, i_3954);
  nand ginst1534 (i_4488, i_2235, i_3956);
  not ginst1535 (i_4489, i_3535);
  nand ginst1536 (i_4490, i_3535, i_3958);
  not ginst1537 (i_4491, i_3539);
  not ginst1538 (i_4492, i_3542);
  not ginst1539 (i_4493, i_3545);
  not ginst1540 (i_4494, i_3548);
  not ginst1541 (i_4495, i_3553);
  nand ginst1542 (i_4496, i_3553, i_3964);
  not ginst1543 (i_4497, i_3557);
  not ginst1544 (i_4498, i_3560);
  not ginst1545 (i_4499, i_3563);
  not ginst1546 (i_4500, i_3566);
  not ginst1547 (i_4501, i_3571);
  nand ginst1548 (i_4502, i_3167, i_3571);
  not ginst1549 (i_4503, i_3574);
  not ginst1550 (i_4504, i_3577);
  not ginst1551 (i_4505, i_3580);
  not ginst1552 (i_4506, i_3583);
  nand ginst1553 (i_4507, i_1867, i_3598);
  not ginst1554 (i_4508, i_3598);
  nand ginst1555 (i_4509, i_1868, i_3601);
  not ginst1556 (i_4510, i_3601);
  nand ginst1557 (i_4511, i_1869, i_3604);
  not ginst1558 (i_4512, i_3604);
  nand ginst1559 (i_4513, i_1870, i_3607);
  not ginst1560 (i_4514, i_3607);
  nand ginst1561 (i_4515, i_1871, i_3610);
  not ginst1562 (i_4516, i_3610);
  nand ginst1563 (i_4517, i_1872, i_3613);
  not ginst1564 (i_4518, i_3613);
  nand ginst1565 (i_4519, i_1873, i_3616);
  not ginst1566 (i_4520, i_3616);
  nand ginst1567 (i_4521, i_1874, i_3619);
  not ginst1568 (i_4522, i_3619);
  nand ginst1569 (i_4523, i_1875, i_3622);
  not ginst1570 (i_4524, i_3622);
  nand ginst1571 (i_4525, i_1876, i_3631);
  not ginst1572 (i_4526, i_3631);
  nand ginst1573 (i_4527, i_1877, i_3634);
  not ginst1574 (i_4528, i_3634);
  nand ginst1575 (i_4529, i_1878, i_3637);
  not ginst1576 (i_4530, i_3637);
  nand ginst1577 (i_4531, i_1879, i_3640);
  not ginst1578 (i_4532, i_3640);
  nand ginst1579 (i_4533, i_1880, i_3643);
  not ginst1580 (i_4534, i_3643);
  nand ginst1581 (i_4535, i_1881, i_3646);
  not ginst1582 (i_4536, i_3646);
  nand ginst1583 (i_4537, i_1882, i_3649);
  not ginst1584 (i_4538, i_3649);
  nand ginst1585 (i_4539, i_1883, i_3652);
  not ginst1586 (i_4540, i_3652);
  nand ginst1587 (i_4541, i_1884, i_3655);
  not ginst1588 (i_4542, i_3655);
  not ginst1589 (i_4543, i_3658);
  and ginst1590 (i_4544, i_3293, i_806);
  and ginst1591 (i_4545, i_3287, i_800);
  and ginst1592 (i_4549, i_3281, i_794);
  and ginst1593 (i_4555, i_3273, i_786);
  and ginst1594 (i_4562, i_3267, i_780);
  and ginst1595 (i_4563, i_3355, i_774);
  and ginst1596 (i_4566, i_3349, i_768);
  and ginst1597 (i_4570, i_3343, i_762);
  not ginst1598 (i_4575, i_3661);
  and ginst1599 (i_4576, i_3293, i_806);
  and ginst1600 (i_4577, i_3287, i_800);
  and ginst1601 (i_4581, i_3281, i_794);
  and ginst1602 (i_4586, i_3273, i_786);
  and ginst1603 (i_4592, i_3267, i_780);
  and ginst1604 (i_4593, i_3355, i_774);
  and ginst1605 (i_4597, i_3349, i_768);
  and ginst1606 (i_4603, i_3343, i_762);
  not ginst1607 (i_4610, i_3664);
  not ginst1608 (i_4611, i_3667);
  not ginst1609 (i_4612, i_3670);
  not ginst1610 (i_4613, i_3673);
  not ginst1611 (i_4614, i_3676);
  not ginst1612 (i_4615, i_3679);
  not ginst1613 (i_4616, i_3682);
  not ginst1614 (i_4617, i_3685);
  not ginst1615 (i_4618, i_3688);
  not ginst1616 (i_4619, i_3691);
  not ginst1617 (i_4620, i_3694);
  not ginst1618 (i_4621, i_3697);
  not ginst1619 (i_4622, i_3700);
  not ginst1620 (i_4623, i_3703);
  not ginst1621 (i_4624, i_3706);
  not ginst1622 (i_4625, i_3709);
  not ginst1623 (i_4626, i_3712);
  not ginst1624 (i_4627, i_3715);
  not ginst1625 (i_4628, i_3718);
  not ginst1626 (i_4629, i_3721);
  and ginst1627 (i_4630, i_2704, i_3448);
  not ginst1628 (i_4631, i_3724);
  and ginst1629 (i_4632, i_2700, i_3444);
  not ginst1630 (i_4633, i_3727);
  and ginst1631 (i_4634, i_2696, i_3440);
  and ginst1632 (i_4635, i_2692, i_3436);
  not ginst1633 (i_4636, i_3730);
  and ginst1634 (i_4637, i_2688, i_3432);
  and ginst1635 (i_4638, i_3311, i_3428);
  and ginst1636 (i_4639, i_3307, i_3424);
  and ginst1637 (i_4640, i_3303, i_3420);
  and ginst1638 (i_4641, i_3299, i_3416);
  not ginst1639 (i_4642, i_3733);
  not ginst1640 (i_4643, i_3736);
  not ginst1641 (i_4644, i_3739);
  not ginst1642 (i_4645, i_3742);
  not ginst1643 (i_4646, i_3745);
  not ginst1644 (i_4647, i_3748);
  not ginst1645 (i_4648, i_3751);
  not ginst1646 (i_4649, i_3754);
  not ginst1647 (i_4650, i_3757);
  not ginst1648 (i_4651, i_3760);
  not ginst1649 (i_4652, i_3763);
  not ginst1650 (i_4653, i_3375);
  and ginst1651 (i_4656, i_3410, i_865);
  and ginst1652 (i_4657, i_3404, i_859);
  and ginst1653 (i_4661, i_3398, i_853);
  and ginst1654 (i_4667, i_3390, i_845);
  not ginst1655 (i_467, i_57);
  and ginst1656 (i_4674, i_3384, i_839);
  and ginst1657 (i_4675, i_3334, i_833);
  and ginst1658 (i_4678, i_3328, i_827);
  and ginst1659 (i_4682, i_3322, i_821);
  and ginst1660 (i_4687, i_3315, i_814);
  and ginst1661 (i_469, i_133, i_134);
  not ginst1662 (i_4693, i_3766);
  nand ginst1663 (i_4694, i_3380, i_3766);
  not ginst1664 (i_4695, i_3769);
  not ginst1665 (i_4696, i_3772);
  not ginst1666 (i_4697, i_3775);
  not ginst1667 (i_4698, i_3778);
  not ginst1668 (i_4699, i_3783);
  not ginst1669 (i_4700, i_3786);
  and ginst1670 (i_4701, i_3410, i_865);
  and ginst1671 (i_4702, i_3404, i_859);
  and ginst1672 (i_4706, i_3398, i_853);
  and ginst1673 (i_4711, i_3390, i_845);
  and ginst1674 (i_4717, i_3384, i_839);
  and ginst1675 (i_4718, i_3334, i_833);
  and ginst1676 (i_4722, i_3328, i_827);
  and ginst1677 (i_4728, i_3322, i_821);
  and ginst1678 (i_4735, i_3315, i_814);
  not ginst1679 (i_4743, i_3789);
  not ginst1680 (i_4744, i_3792);
  not ginst1681 (i_4745, i_3807);
  nand ginst1682 (i_4746, i_3452, i_3807);
  not ginst1683 (i_4747, i_3810);
  not ginst1684 (i_4748, i_3813);
  not ginst1685 (i_4749, i_3816);
  not ginst1686 (i_4750, i_3819);
  nand ginst1687 (i_4751, i_3453, i_3819);
  not ginst1688 (i_4752, i_3822);
  not ginst1689 (i_4753, i_3825);
  not ginst1690 (i_4754, i_3828);
  not ginst1691 (i_4755, i_3831);
  and ginst1692 (i_4756, i_3263, i_3482);
  and ginst1693 (i_4757, i_3259, i_3478);
  and ginst1694 (i_4758, i_3255, i_3474);
  and ginst1695 (i_4759, i_3251, i_3470);
  and ginst1696 (i_4760, i_3247, i_3466);
  not ginst1697 (i_4761, i_3846);
  and ginst1698 (i_4762, i_2615, i_3462);
  not ginst1699 (i_4763, i_3849);
  and ginst1700 (i_4764, i_2611, i_3458);
  not ginst1701 (i_4765, i_3852);
  and ginst1702 (i_4766, i_2607, i_3454);
  and ginst1703 (i_4767, i_2680, i_3381);
  not ginst1704 (i_4768, i_3855);
  and ginst1705 (i_4769, i_3340, i_695);
  not ginst1706 (i_4775, i_3858);
  nand ginst1707 (i_4776, i_3486, i_3858);
  not ginst1708 (i_4777, i_3861);
  not ginst1709 (i_4778, i_3864);
  not ginst1710 (i_4779, i_3867);
  not ginst1711 (i_478, i_248);
  not ginst1712 (i_4780, i_3870);
  not ginst1713 (i_4781, i_3885);
  not ginst1714 (i_4782, i_3888);
  not ginst1715 (i_4783, i_3891);
  or ginst1716 (i_4784, i_3131, i_3134);
  not ginst1717 (i_4789, i_3502);
  not ginst1718 (i_4790, i_3131);
  not ginst1719 (i_4793, i_3507);
  not ginst1720 (i_4794, i_3510);
  not ginst1721 (i_4795, i_3515);
  not ginst1722 (i_4796, i_3114);
  not ginst1723 (i_4799, i_3586);
  not ginst1724 (i_4800, i_3589);
  not ginst1725 (i_4801, i_3592);
  not ginst1726 (i_4802, i_3595);
  nand ginst1727 (i_4803, i_4326, i_4327);
  nand ginst1728 (i_4806, i_4333, i_4334);
  not ginst1729 (i_4809, i_3625);
  not ginst1730 (i_4810, i_3178);
  not ginst1731 (i_4813, i_3628);
  not ginst1732 (i_4814, i_3202);
  not ginst1733 (i_4817, i_3221);
  not ginst1734 (i_482, i_254);
  not ginst1735 (i_4820, i_3293);
  not ginst1736 (i_4823, i_3287);
  not ginst1737 (i_4826, i_3281);
  not ginst1738 (i_4829, i_3273);
  not ginst1739 (i_4832, i_3267);
  not ginst1740 (i_4835, i_3355);
  not ginst1741 (i_4838, i_3349);
  not ginst1742 (i_484, i_257);
  not ginst1743 (i_4841, i_3343);
  nor ginst1744 (i_4844, i_3273, i_786);
  not ginst1745 (i_4847, i_3293);
  not ginst1746 (i_4850, i_3287);
  not ginst1747 (i_4853, i_3281);
  not ginst1748 (i_4856, i_3267);
  not ginst1749 (i_4859, i_3355);
  not ginst1750 (i_486, i_260);
  not ginst1751 (i_4862, i_3349);
  not ginst1752 (i_4865, i_3343);
  not ginst1753 (i_4868, i_3273);
  nor ginst1754 (i_4871, i_3273, i_786);
  not ginst1755 (i_4874, i_3448);
  not ginst1756 (i_4877, i_3444);
  not ginst1757 (i_4880, i_3440);
  not ginst1758 (i_4883, i_3432);
  not ginst1759 (i_4886, i_3428);
  not ginst1760 (i_4889, i_3311);
  not ginst1761 (i_489, i_263);
  not ginst1762 (i_4892, i_3424);
  not ginst1763 (i_4895, i_3307);
  not ginst1764 (i_4898, i_3420);
  not ginst1765 (i_4901, i_3303);
  not ginst1766 (i_4904, i_3436);
  not ginst1767 (i_4907, i_3416);
  not ginst1768 (i_4910, i_3299);
  not ginst1769 (i_4913, i_3410);
  not ginst1770 (i_4916, i_3404);
  not ginst1771 (i_4919, i_3398);
  not ginst1772 (i_492, i_267);
  not ginst1773 (i_4922, i_3390);
  not ginst1774 (i_4925, i_3384);
  not ginst1775 (i_4928, i_3334);
  not ginst1776 (i_4931, i_3328);
  not ginst1777 (i_4934, i_3322);
  not ginst1778 (i_4937, i_3315);
  and ginst1779 (i_494, i_162, i_172, i_188, i_199);
  nor ginst1780 (i_4940, i_3390, i_845);
  not ginst1781 (i_4943, i_3315);
  not ginst1782 (i_4946, i_3328);
  not ginst1783 (i_4949, i_3322);
  not ginst1784 (i_4952, i_3384);
  not ginst1785 (i_4955, i_3334);
  not ginst1786 (i_4958, i_3398);
  not ginst1787 (i_4961, i_3390);
  not ginst1788 (i_4964, i_3410);
  not ginst1789 (i_4967, i_3404);
  not ginst1790 (i_4970, i_3340);
  not ginst1791 (i_4973, i_3349);
  not ginst1792 (i_4976, i_3343);
  not ginst1793 (i_4979, i_3267);
  not ginst1794 (i_4982, i_3355);
  not ginst1795 (i_4985, i_3281);
  not ginst1796 (i_4988, i_3273);
  not ginst1797 (i_4991, i_3293);
  not ginst1798 (i_4994, i_3287);
  nand ginst1799 (i_4997, i_4411, i_4412);
  not ginst1800 (i_5000, i_3410);
  not ginst1801 (i_5003, i_3404);
  not ginst1802 (i_5006, i_3398);
  not ginst1803 (i_5009, i_3384);
  not ginst1804 (i_501, i_274);
  not ginst1805 (i_5012, i_3334);
  not ginst1806 (i_5015, i_3328);
  not ginst1807 (i_5018, i_3322);
  not ginst1808 (i_5021, i_3390);
  not ginst1809 (i_5024, i_3315);
  nor ginst1810 (i_5027, i_3390, i_845);
  nor ginst1811 (i_5030, i_3315, i_814);
  not ginst1812 (i_5033, i_3299);
  not ginst1813 (i_5036, i_3307);
  not ginst1814 (i_5039, i_3303);
  not ginst1815 (i_5042, i_3311);
  not ginst1816 (i_5045, i_3795);
  not ginst1817 (i_5046, i_3798);
  not ginst1818 (i_5047, i_3801);
  not ginst1819 (i_5048, i_3804);
  not ginst1820 (i_5049, i_3247);
  not ginst1821 (i_505, i_280);
  not ginst1822 (i_5052, i_3255);
  not ginst1823 (i_5055, i_3251);
  not ginst1824 (i_5058, i_3263);
  not ginst1825 (i_5061, i_3259);
  not ginst1826 (i_5064, i_3834);
  not ginst1827 (i_5065, i_3837);
  not ginst1828 (i_5066, i_3840);
  not ginst1829 (i_5067, i_3843);
  not ginst1830 (i_5068, i_3482);
  not ginst1831 (i_507, i_283);
  not ginst1832 (i_5071, i_3263);
  not ginst1833 (i_5074, i_3478);
  not ginst1834 (i_5077, i_3259);
  not ginst1835 (i_5080, i_3474);
  not ginst1836 (i_5083, i_3255);
  not ginst1837 (i_5086, i_3466);
  not ginst1838 (i_5089, i_3247);
  not ginst1839 (i_509, i_286);
  not ginst1840 (i_5092, i_3462);
  not ginst1841 (i_5095, i_3458);
  not ginst1842 (i_5098, i_3454);
  not ginst1843 (i_5101, i_3470);
  not ginst1844 (i_5104, i_3251);
  not ginst1845 (i_5107, i_3381);
  not ginst1846 (i_511, i_289);
  not ginst1847 (i_5110, i_3873);
  not ginst1848 (i_5111, i_3876);
  not ginst1849 (i_5112, i_3879);
  not ginst1850 (i_5113, i_3882);
  not ginst1851 (i_5114, i_3458);
  not ginst1852 (i_5117, i_3454);
  not ginst1853 (i_5120, i_3466);
  not ginst1854 (i_5123, i_3462);
  not ginst1855 (i_5126, i_3474);
  not ginst1856 (i_5129, i_3470);
  not ginst1857 (i_513, i_293);
  not ginst1858 (i_5132, i_3482);
  not ginst1859 (i_5135, i_3478);
  not ginst1860 (i_5138, i_3416);
  not ginst1861 (i_5141, i_3424);
  not ginst1862 (i_5144, i_3420);
  not ginst1863 (i_5147, i_3432);
  not ginst1864 (i_515, i_296);
  not ginst1865 (i_5150, i_3428);
  not ginst1866 (i_5153, i_3440);
  not ginst1867 (i_5156, i_3436);
  not ginst1868 (i_5159, i_3448);
  not ginst1869 (i_5162, i_3444);
  nand ginst1870 (i_5165, i_4485, i_4486);
  nand ginst1871 (i_5166, i_4473, i_4474);
  nand ginst1872 (i_5167, i_1290, i_4464);
  nand ginst1873 (i_5168, i_1293, i_4466);
  nand ginst1874 (i_5169, i_2074, i_4468);
  not ginst1875 (i_517, i_299);
  nand ginst1876 (i_5170, i_1296, i_4470);
  nand ginst1877 (i_5171, i_1302, i_4472);
  nand ginst1878 (i_5172, i_1314, i_4476);
  nand ginst1879 (i_5173, i_1317, i_4478);
  nand ginst1880 (i_5174, i_2081, i_4480);
  nand ginst1881 (i_5175, i_1320, i_4482);
  nand ginst1882 (i_5176, i_1323, i_4484);
  nand ginst1883 (i_5177, i_3953, i_4487);
  nand ginst1884 (i_5178, i_3955, i_4488);
  nand ginst1885 (i_5179, i_3073, i_4489);
  nand ginst1886 (i_5180, i_3542, i_4491);
  nand ginst1887 (i_5181, i_3539, i_4492);
  nand ginst1888 (i_5182, i_3548, i_4493);
  nand ginst1889 (i_5183, i_3545, i_4494);
  nand ginst1890 (i_5184, i_3080, i_4495);
  nand ginst1891 (i_5185, i_3560, i_4497);
  nand ginst1892 (i_5186, i_3557, i_4498);
  nand ginst1893 (i_5187, i_3566, i_4499);
  nand ginst1894 (i_5188, i_3563, i_4500);
  nand ginst1895 (i_5189, i_2778, i_4501);
  not ginst1896 (i_519, i_303);
  nand ginst1897 (i_5190, i_3577, i_4503);
  nand ginst1898 (i_5191, i_3574, i_4504);
  nand ginst1899 (i_5192, i_3583, i_4505);
  nand ginst1900 (i_5193, i_3580, i_4506);
  nand ginst1901 (i_5196, i_1326, i_4508);
  nand ginst1902 (i_5197, i_1329, i_4510);
  nand ginst1903 (i_5198, i_1332, i_4512);
  nand ginst1904 (i_5199, i_1335, i_4514);
  nand ginst1905 (i_5200, i_1338, i_4516);
  nand ginst1906 (i_5201, i_1341, i_4518);
  nand ginst1907 (i_5202, i_1344, i_4520);
  nand ginst1908 (i_5203, i_1347, i_4522);
  nand ginst1909 (i_5204, i_1350, i_4524);
  nand ginst1910 (i_5205, i_1353, i_4526);
  nand ginst1911 (i_5206, i_1356, i_4528);
  nand ginst1912 (i_5207, i_1359, i_4530);
  nand ginst1913 (i_5208, i_1362, i_4532);
  nand ginst1914 (i_5209, i_1365, i_4534);
  nand ginst1915 (i_5210, i_1368, i_4536);
  nand ginst1916 (i_5211, i_1371, i_4538);
  nand ginst1917 (i_5212, i_1374, i_4540);
  nand ginst1918 (i_5213, i_1377, i_4542);
  and ginst1919 (i_528, i_150, i_184, i_228, i_240);
  nand ginst1920 (i_5283, i_3670, i_4611);
  nand ginst1921 (i_5284, i_3667, i_4612);
  nand ginst1922 (i_5285, i_3676, i_4613);
  nand ginst1923 (i_5286, i_3673, i_4614);
  nand ginst1924 (i_5287, i_3682, i_4615);
  nand ginst1925 (i_5288, i_3679, i_4616);
  nand ginst1926 (i_5289, i_3688, i_4617);
  nand ginst1927 (i_5290, i_3685, i_4618);
  nand ginst1928 (i_5291, i_3694, i_4619);
  nand ginst1929 (i_5292, i_3691, i_4620);
  nand ginst1930 (i_5293, i_3700, i_4621);
  nand ginst1931 (i_5294, i_3697, i_4622);
  nand ginst1932 (i_5295, i_3706, i_4623);
  nand ginst1933 (i_5296, i_3703, i_4624);
  nand ginst1934 (i_5297, i_3712, i_4625);
  nand ginst1935 (i_5298, i_3709, i_4626);
  nand ginst1936 (i_5299, i_3718, i_4627);
  nand ginst1937 (i_5300, i_3715, i_4628);
  nand ginst1938 (i_5314, i_3739, i_4643);
  nand ginst1939 (i_5315, i_3736, i_4644);
  nand ginst1940 (i_5316, i_3745, i_4645);
  nand ginst1941 (i_5317, i_3742, i_4646);
  nand ginst1942 (i_5318, i_3751, i_4647);
  nand ginst1943 (i_5319, i_3748, i_4648);
  nand ginst1944 (i_5320, i_3757, i_4649);
  nand ginst1945 (i_5321, i_3754, i_4650);
  nand ginst1946 (i_5322, i_3763, i_4651);
  nand ginst1947 (i_5323, i_3760, i_4652);
  not ginst1948 (i_5324, i_4193);
  not ginst1949 (i_535, i_307);
  nand ginst1950 (i_5363, i_2781, i_4693);
  nand ginst1951 (i_5364, i_3772, i_4695);
  nand ginst1952 (i_5365, i_3769, i_4696);
  nand ginst1953 (i_5366, i_3778, i_4697);
  nand ginst1954 (i_5367, i_3775, i_4698);
  not ginst1955 (i_537, i_310);
  not ginst1956 (i_539, i_313);
  not ginst1957 (i_541, i_316);
  nand ginst1958 (i_5425, i_2790, i_4745);
  nand ginst1959 (i_5426, i_3813, i_4747);
  nand ginst1960 (i_5427, i_3810, i_4748);
  nand ginst1961 (i_5429, i_2793, i_4750);
  not ginst1962 (i_543, i_319);
  nand ginst1963 (i_5430, i_3825, i_4752);
  nand ginst1964 (i_5431, i_3822, i_4753);
  nand ginst1965 (i_5432, i_3831, i_4754);
  nand ginst1966 (i_5433, i_3828, i_4755);
  not ginst1967 (i_545, i_322);
  nand ginst1968 (i_5451, i_2796, i_4775);
  nand ginst1969 (i_5452, i_3864, i_4777);
  nand ginst1970 (i_5453, i_3861, i_4778);
  nand ginst1971 (i_5454, i_3870, i_4779);
  nand ginst1972 (i_5455, i_3867, i_4780);
  nand ginst1973 (i_5456, i_3888, i_4781);
  nand ginst1974 (i_5457, i_3885, i_4782);
  not ginst1975 (i_5469, i_4303);
  not ginst1976 (i_547, i_325);
  nand ginst1977 (i_5474, i_3589, i_4799);
  nand ginst1978 (i_5475, i_3586, i_4800);
  nand ginst1979 (i_5476, i_3595, i_4801);
  nand ginst1980 (i_5477, i_3592, i_4802);
  not ginst1981 (i_549, i_328);
  not ginst1982 (i_551, i_331);
  not ginst1983 (i_553, i_334);
  not ginst1984 (i_556, i_337);
  nand ginst1985 (i_5571, i_3798, i_5045);
  nand ginst1986 (i_5572, i_3795, i_5046);
  nand ginst1987 (i_5573, i_3804, i_5047);
  nand ginst1988 (i_5574, i_3801, i_5048);
  nand ginst1989 (i_5584, i_3837, i_5064);
  nand ginst1990 (i_5585, i_3834, i_5065);
  nand ginst1991 (i_5586, i_3843, i_5066);
  nand ginst1992 (i_5587, i_3840, i_5067);
  not ginst1993 (i_559, i_343);
  nand ginst1994 (i_5602, i_3876, i_5110);
  nand ginst1995 (i_5603, i_3873, i_5111);
  nand ginst1996 (i_5604, i_3882, i_5112);
  nand ginst1997 (i_5605, i_3879, i_5113);
  not ginst1998 (i_561, i_346);
  not ginst1999 (i_563, i_349);
  nand ginst2000 (i_5631, i_4653, i_5324);
  nand ginst2001 (i_5632, i_4463, i_5167);
  nand ginst2002 (i_5640, i_4465, i_5168);
  not ginst2003 (i_565, i_352);
  nand ginst2004 (i_5654, i_4467, i_5169);
  not ginst2005 (i_567, i_355);
  nand ginst2006 (i_5670, i_4469, i_5170);
  nand ginst2007 (i_5683, i_4471, i_5171);
  not ginst2008 (i_569, i_358);
  nand ginst2009 (i_5690, i_4475, i_5172);
  nand ginst2010 (i_5697, i_4477, i_5173);
  nand ginst2011 (i_5707, i_4479, i_5174);
  not ginst2012 (i_571, i_361);
  nand ginst2013 (i_5718, i_4481, i_5175);
  nand ginst2014 (i_5728, i_4483, i_5176);
  not ginst2015 (i_573, i_364);
  not ginst2016 (i_5735, i_5177);
  nand ginst2017 (i_5736, i_4490, i_5179);
  nand ginst2018 (i_5740, i_5180, i_5181);
  nand ginst2019 (i_5744, i_5182, i_5183);
  nand ginst2020 (i_5747, i_4496, i_5184);
  and ginst2021 (i_575, i_182, i_183, i_185, i_186);
  nand ginst2022 (i_5751, i_5185, i_5186);
  nand ginst2023 (i_5755, i_5187, i_5188);
  nand ginst2024 (i_5758, i_4502, i_5189);
  nand ginst2025 (i_5762, i_5190, i_5191);
  nand ginst2026 (i_5766, i_5192, i_5193);
  not ginst2027 (i_5769, i_4803);
  not ginst2028 (i_5770, i_4806);
  nand ginst2029 (i_5771, i_4507, i_5196);
  nand ginst2030 (i_5778, i_4509, i_5197);
  and ginst2031 (i_578, i_152, i_210, i_218, i_230);
  nand ginst2032 (i_5789, i_4511, i_5198);
  nand ginst2033 (i_5799, i_4513, i_5199);
  nand ginst2034 (i_5807, i_4515, i_5200);
  not ginst2035 (i_582, i_15);
  nand ginst2036 (i_5821, i_4517, i_5201);
  nand ginst2037 (i_5837, i_4519, i_5202);
  not ginst2038 (i_585, i_5);
  nand ginst2039 (i_5850, i_4521, i_5203);
  nand ginst2040 (i_5856, i_4523, i_5204);
  nand ginst2041 (i_5863, i_4525, i_5205);
  nand ginst2042 (i_5870, i_4527, i_5206);
  nand ginst2043 (i_5881, i_4529, i_5207);
  nand ginst2044 (i_5892, i_4531, i_5208);
  nand ginst2045 (i_5898, i_4533, i_5209);
  not ginst2046 (i_590, i_1);
  nand ginst2047 (i_5905, i_4535, i_5210);
  nand ginst2048 (i_5915, i_4537, i_5211);
  nand ginst2049 (i_5926, i_4539, i_5212);
  not ginst2050 (i_593, i_5);
  nand ginst2051 (i_5936, i_4541, i_5213);
  not ginst2052 (i_5943, i_4817);
  nand ginst2053 (i_5944, i_1931, i_4820);
  not ginst2054 (i_5945, i_4820);
  nand ginst2055 (i_5946, i_1932, i_4823);
  not ginst2056 (i_5947, i_4823);
  nand ginst2057 (i_5948, i_1933, i_4826);
  not ginst2058 (i_5949, i_4826);
  nand ginst2059 (i_5950, i_1934, i_4829);
  not ginst2060 (i_5951, i_4829);
  nand ginst2061 (i_5952, i_1935, i_4832);
  not ginst2062 (i_5953, i_4832);
  nand ginst2063 (i_5954, i_1936, i_4835);
  not ginst2064 (i_5955, i_4835);
  nand ginst2065 (i_5956, i_1937, i_4838);
  not ginst2066 (i_5957, i_4838);
  nand ginst2067 (i_5958, i_1938, i_4841);
  not ginst2068 (i_5959, i_4841);
  not ginst2069 (i_596, i_5);
  and ginst2070 (i_5960, i_2674, i_4769);
  not ginst2071 (i_5966, i_4844);
  nand ginst2072 (i_5967, i_1939, i_4847);
  not ginst2073 (i_5968, i_4847);
  nand ginst2074 (i_5969, i_1940, i_4850);
  not ginst2075 (i_5970, i_4850);
  nand ginst2076 (i_5971, i_1941, i_4853);
  not ginst2077 (i_5972, i_4853);
  nand ginst2078 (i_5973, i_1942, i_4856);
  not ginst2079 (i_5974, i_4856);
  nand ginst2080 (i_5975, i_1943, i_4859);
  not ginst2081 (i_5976, i_4859);
  nand ginst2082 (i_5977, i_1944, i_4862);
  not ginst2083 (i_5978, i_4862);
  nand ginst2084 (i_5979, i_1945, i_4865);
  not ginst2085 (i_5980, i_4865);
  and ginst2086 (i_5981, i_2674, i_4769);
  nand ginst2087 (i_5989, i_1946, i_4868);
  not ginst2088 (i_599, i_289);
  not ginst2089 (i_5990, i_4868);
  nand ginst2090 (i_5991, i_5283, i_5284);
  nand ginst2091 (i_5996, i_5285, i_5286);
  nand ginst2092 (i_6000, i_5287, i_5288);
  nand ginst2093 (i_6003, i_5289, i_5290);
  nand ginst2094 (i_6009, i_5291, i_5292);
  nand ginst2095 (i_6014, i_5293, i_5294);
  nand ginst2096 (i_6018, i_5295, i_5296);
  nand ginst2097 (i_6021, i_5297, i_5298);
  nand ginst2098 (i_6022, i_5299, i_5300);
  not ginst2099 (i_6023, i_4874);
  nand ginst2100 (i_6024, i_4629, i_4874);
  not ginst2101 (i_6025, i_4877);
  nand ginst2102 (i_6026, i_4631, i_4877);
  not ginst2103 (i_6027, i_4880);
  nand ginst2104 (i_6028, i_4633, i_4880);
  not ginst2105 (i_6029, i_4883);
  nand ginst2106 (i_6030, i_4636, i_4883);
  not ginst2107 (i_6031, i_4886);
  not ginst2108 (i_6032, i_4889);
  not ginst2109 (i_6033, i_4892);
  not ginst2110 (i_6034, i_4895);
  not ginst2111 (i_6035, i_4898);
  not ginst2112 (i_6036, i_4901);
  not ginst2113 (i_6037, i_4904);
  nand ginst2114 (i_6038, i_4642, i_4904);
  not ginst2115 (i_6039, i_4907);
  not ginst2116 (i_604, i_299);
  not ginst2117 (i_6040, i_4910);
  nand ginst2118 (i_6041, i_5314, i_5315);
  nand ginst2119 (i_6047, i_5316, i_5317);
  nand ginst2120 (i_6052, i_5318, i_5319);
  nand ginst2121 (i_6056, i_5320, i_5321);
  nand ginst2122 (i_6059, i_5322, i_5323);
  nand ginst2123 (i_6060, i_1968, i_4913);
  not ginst2124 (i_6061, i_4913);
  nand ginst2125 (i_6062, i_1969, i_4916);
  not ginst2126 (i_6063, i_4916);
  nand ginst2127 (i_6064, i_1970, i_4919);
  not ginst2128 (i_6065, i_4919);
  nand ginst2129 (i_6066, i_1971, i_4922);
  not ginst2130 (i_6067, i_4922);
  nand ginst2131 (i_6068, i_1972, i_4925);
  not ginst2132 (i_6069, i_4925);
  nand ginst2133 (i_6070, i_1973, i_4928);
  not ginst2134 (i_6071, i_4928);
  nand ginst2135 (i_6072, i_1974, i_4931);
  not ginst2136 (i_6073, i_4931);
  nand ginst2137 (i_6074, i_1975, i_4934);
  not ginst2138 (i_6075, i_4934);
  nand ginst2139 (i_6076, i_1976, i_4937);
  not ginst2140 (i_6077, i_4937);
  not ginst2141 (i_6078, i_4940);
  nand ginst2142 (i_6079, i_4694, i_5363);
  nand ginst2143 (i_6083, i_5364, i_5365);
  nand ginst2144 (i_6087, i_5366, i_5367);
  not ginst2145 (i_609, i_303);
  not ginst2146 (i_6090, i_4943);
  nand ginst2147 (i_6091, i_4699, i_4943);
  not ginst2148 (i_6092, i_4946);
  not ginst2149 (i_6093, i_4949);
  not ginst2150 (i_6094, i_4952);
  not ginst2151 (i_6095, i_4955);
  not ginst2152 (i_6096, i_4970);
  nand ginst2153 (i_6097, i_4700, i_4970);
  not ginst2154 (i_6098, i_4973);
  not ginst2155 (i_6099, i_4976);
  not ginst2156 (i_6100, i_4979);
  not ginst2157 (i_6101, i_4982);
  not ginst2158 (i_6102, i_4997);
  nand ginst2159 (i_6103, i_2015, i_5000);
  not ginst2160 (i_6104, i_5000);
  nand ginst2161 (i_6105, i_2016, i_5003);
  not ginst2162 (i_6106, i_5003);
  nand ginst2163 (i_6107, i_2017, i_5006);
  not ginst2164 (i_6108, i_5006);
  nand ginst2165 (i_6109, i_2018, i_5009);
  not ginst2166 (i_6110, i_5009);
  nand ginst2167 (i_6111, i_2019, i_5012);
  not ginst2168 (i_6112, i_5012);
  nand ginst2169 (i_6113, i_2020, i_5015);
  not ginst2170 (i_6114, i_5015);
  nand ginst2171 (i_6115, i_2021, i_5018);
  not ginst2172 (i_6116, i_5018);
  nand ginst2173 (i_6117, i_2022, i_5021);
  not ginst2174 (i_6118, i_5021);
  nand ginst2175 (i_6119, i_2023, i_5024);
  not ginst2176 (i_6120, i_5024);
  not ginst2177 (i_6121, i_5033);
  nand ginst2178 (i_6122, i_4743, i_5033);
  not ginst2179 (i_6123, i_5036);
  not ginst2180 (i_6124, i_5039);
  nand ginst2181 (i_6125, i_4744, i_5042);
  not ginst2182 (i_6126, i_5042);
  nand ginst2183 (i_6127, i_4746, i_5425);
  nand ginst2184 (i_6131, i_5426, i_5427);
  not ginst2185 (i_6135, i_5049);
  nand ginst2186 (i_6136, i_4749, i_5049);
  nand ginst2187 (i_6137, i_4751, i_5429);
  not ginst2188 (i_614, i_38);
  nand ginst2189 (i_6141, i_5430, i_5431);
  nand ginst2190 (i_6145, i_5432, i_5433);
  not ginst2191 (i_6148, i_5068);
  not ginst2192 (i_6149, i_5071);
  not ginst2193 (i_6150, i_5074);
  not ginst2194 (i_6151, i_5077);
  not ginst2195 (i_6152, i_5080);
  not ginst2196 (i_6153, i_5083);
  not ginst2197 (i_6154, i_5086);
  not ginst2198 (i_6155, i_5089);
  not ginst2199 (i_6156, i_5092);
  nand ginst2200 (i_6157, i_4761, i_5092);
  not ginst2201 (i_6158, i_5095);
  nand ginst2202 (i_6159, i_4763, i_5095);
  not ginst2203 (i_6160, i_5098);
  nand ginst2204 (i_6161, i_4765, i_5098);
  not ginst2205 (i_6162, i_5101);
  not ginst2206 (i_6163, i_5104);
  nand ginst2207 (i_6164, i_4768, i_5107);
  not ginst2208 (i_6165, i_5107);
  nand ginst2209 (i_6166, i_4776, i_5451);
  nand ginst2210 (i_6170, i_5452, i_5453);
  nand ginst2211 (i_6174, i_5454, i_5455);
  nand ginst2212 (i_6177, i_5456, i_5457);
  not ginst2213 (i_6181, i_5114);
  not ginst2214 (i_6182, i_5117);
  not ginst2215 (i_6183, i_5120);
  not ginst2216 (i_6184, i_5123);
  not ginst2217 (i_6185, i_5138);
  nand ginst2218 (i_6186, i_4783, i_5138);
  not ginst2219 (i_6187, i_5141);
  not ginst2220 (i_6188, i_5144);
  not ginst2221 (i_6189, i_5147);
  not ginst2222 (i_6190, i_5150);
  not ginst2223 (i_6191, i_4784);
  nand ginst2224 (i_6192, i_2230, i_4784);
  not ginst2225 (i_6193, i_4790);
  nand ginst2226 (i_6194, i_2765, i_4790);
  not ginst2227 (i_6195, i_4796);
  nand ginst2228 (i_6196, i_5476, i_5477);
  nand ginst2229 (i_6199, i_5474, i_5475);
  not ginst2230 (i_6202, i_4810);
  not ginst2231 (i_6203, i_4814);
  not ginst2232 (i_6204, i_4769);
  not ginst2233 (i_6207, i_4555);
  not ginst2234 (i_6210, i_4769);
  not ginst2235 (i_6213, i_4871);
  not ginst2236 (i_6214, i_4586);
  nor ginst2237 (i_6217, i_2674, i_4769);
  not ginst2238 (i_6220, i_4667);
  not ginst2239 (i_6223, i_4958);
  not ginst2240 (i_6224, i_4961);
  not ginst2241 (i_6225, i_4964);
  not ginst2242 (i_6226, i_4967);
  not ginst2243 (i_6227, i_4985);
  not ginst2244 (i_6228, i_4988);
  not ginst2245 (i_6229, i_4991);
  not ginst2246 (i_6230, i_4994);
  not ginst2247 (i_6231, i_5027);
  not ginst2248 (i_6232, i_4711);
  not ginst2249 (i_6235, i_5030);
  not ginst2250 (i_6236, i_4735);
  not ginst2251 (i_6239, i_5052);
  not ginst2252 (i_6240, i_5055);
  not ginst2253 (i_6241, i_5058);
  not ginst2254 (i_6242, i_5061);
  nand ginst2255 (i_6243, i_5573, i_5574);
  nand ginst2256 (i_6246, i_5571, i_5572);
  nand ginst2257 (i_6249, i_5586, i_5587);
  not ginst2258 (i_625, i_15);
  nand ginst2259 (i_6252, i_5584, i_5585);
  not ginst2260 (i_6255, i_5126);
  not ginst2261 (i_6256, i_5129);
  not ginst2262 (i_6257, i_5132);
  not ginst2263 (i_6258, i_5135);
  not ginst2264 (i_6259, i_5153);
  not ginst2265 (i_6260, i_5156);
  not ginst2266 (i_6261, i_5159);
  not ginst2267 (i_6262, i_5162);
  nand ginst2268 (i_6263, i_5604, i_5605);
  nand ginst2269 (i_6266, i_5602, i_5603);
  nand ginst2270 (i_628, i_9, i_12);
  nand ginst2271 (i_632, i_9, i_12);
  not ginst2272 (i_636, i_38);
  not ginst2273 (i_641, i_245);
  not ginst2274 (i_642, i_248);
  not ginst2275 (i_643, i_251);
  not ginst2276 (i_644, i_251);
  not ginst2277 (i_651, i_254);
  nand ginst2278 (i_6540, i_1380, i_5945);
  nand ginst2279 (i_6541, i_1383, i_5947);
  nand ginst2280 (i_6542, i_1386, i_5949);
  nand ginst2281 (i_6543, i_1389, i_5951);
  nand ginst2282 (i_6544, i_1392, i_5953);
  nand ginst2283 (i_6545, i_1395, i_5955);
  nand ginst2284 (i_6546, i_1398, i_5957);
  nand ginst2285 (i_6547, i_1401, i_5959);
  nand ginst2286 (i_6555, i_1404, i_5968);
  nand ginst2287 (i_6556, i_1407, i_5970);
  nand ginst2288 (i_6557, i_1410, i_5972);
  nand ginst2289 (i_6558, i_1413, i_5974);
  nand ginst2290 (i_6559, i_1416, i_5976);
  nand ginst2291 (i_6560, i_1419, i_5978);
  nand ginst2292 (i_6561, i_1422, i_5980);
  nand ginst2293 (i_6569, i_1425, i_5990);
  not ginst2294 (i_657, i_106);
  nand ginst2295 (i_6594, i_3721, i_6023);
  nand ginst2296 (i_6595, i_3724, i_6025);
  nand ginst2297 (i_6596, i_3727, i_6027);
  nand ginst2298 (i_6597, i_3730, i_6029);
  nand ginst2299 (i_6598, i_4889, i_6031);
  nand ginst2300 (i_6599, i_4886, i_6032);
  not ginst2301 (i_660, i_257);
  nand ginst2302 (i_6600, i_4895, i_6033);
  nand ginst2303 (i_6601, i_4892, i_6034);
  nand ginst2304 (i_6602, i_4901, i_6035);
  nand ginst2305 (i_6603, i_4898, i_6036);
  nand ginst2306 (i_6604, i_3733, i_6037);
  nand ginst2307 (i_6605, i_4910, i_6039);
  nand ginst2308 (i_6606, i_4907, i_6040);
  nand ginst2309 (i_6621, i_1434, i_6061);
  nand ginst2310 (i_6622, i_1437, i_6063);
  nand ginst2311 (i_6623, i_1440, i_6065);
  nand ginst2312 (i_6624, i_1443, i_6067);
  nand ginst2313 (i_6625, i_1446, i_6069);
  nand ginst2314 (i_6626, i_1449, i_6071);
  nand ginst2315 (i_6627, i_1452, i_6073);
  nand ginst2316 (i_6628, i_1455, i_6075);
  nand ginst2317 (i_6629, i_1458, i_6077);
  nand ginst2318 (i_6639, i_3783, i_6090);
  nand ginst2319 (i_6640, i_4949, i_6092);
  nand ginst2320 (i_6641, i_4946, i_6093);
  nand ginst2321 (i_6642, i_4955, i_6094);
  nand ginst2322 (i_6643, i_4952, i_6095);
  nand ginst2323 (i_6644, i_3786, i_6096);
  nand ginst2324 (i_6645, i_4976, i_6098);
  nand ginst2325 (i_6646, i_4973, i_6099);
  nand ginst2326 (i_6647, i_4982, i_6100);
  nand ginst2327 (i_6648, i_4979, i_6101);
  nand ginst2328 (i_6649, i_1461, i_6104);
  nand ginst2329 (i_6650, i_1464, i_6106);
  nand ginst2330 (i_6651, i_1467, i_6108);
  nand ginst2331 (i_6652, i_1470, i_6110);
  nand ginst2332 (i_6653, i_1473, i_6112);
  nand ginst2333 (i_6654, i_1476, i_6114);
  nand ginst2334 (i_6655, i_1479, i_6116);
  nand ginst2335 (i_6656, i_1482, i_6118);
  nand ginst2336 (i_6657, i_1485, i_6120);
  nand ginst2337 (i_6658, i_3789, i_6121);
  nand ginst2338 (i_6659, i_5039, i_6123);
  not ginst2339 (i_666, i_260);
  nand ginst2340 (i_6660, i_5036, i_6124);
  nand ginst2341 (i_6661, i_3792, i_6126);
  nand ginst2342 (i_6668, i_3816, i_6135);
  nand ginst2343 (i_6677, i_5071, i_6148);
  nand ginst2344 (i_6678, i_5068, i_6149);
  nand ginst2345 (i_6679, i_5077, i_6150);
  nand ginst2346 (i_6680, i_5074, i_6151);
  nand ginst2347 (i_6681, i_5083, i_6152);
  nand ginst2348 (i_6682, i_5080, i_6153);
  nand ginst2349 (i_6683, i_5089, i_6154);
  nand ginst2350 (i_6684, i_5086, i_6155);
  nand ginst2351 (i_6685, i_3846, i_6156);
  nand ginst2352 (i_6686, i_3849, i_6158);
  nand ginst2353 (i_6687, i_3852, i_6160);
  nand ginst2354 (i_6688, i_5104, i_6162);
  nand ginst2355 (i_6689, i_5101, i_6163);
  nand ginst2356 (i_6690, i_3855, i_6165);
  nand ginst2357 (i_6702, i_5117, i_6181);
  nand ginst2358 (i_6703, i_5114, i_6182);
  nand ginst2359 (i_6704, i_5123, i_6183);
  nand ginst2360 (i_6705, i_5120, i_6184);
  nand ginst2361 (i_6706, i_3891, i_6185);
  nand ginst2362 (i_6707, i_5144, i_6187);
  nand ginst2363 (i_6708, i_5141, i_6188);
  nand ginst2364 (i_6709, i_5150, i_6189);
  nand ginst2365 (i_6710, i_5147, i_6190);
  nand ginst2366 (i_6711, i_1708, i_6191);
  nand ginst2367 (i_6712, i_2231, i_6193);
  not ginst2368 (i_672, i_263);
  nand ginst2369 (i_6729, i_4961, i_6223);
  not ginst2370 (i_673, i_267);
  nand ginst2371 (i_6730, i_4958, i_6224);
  nand ginst2372 (i_6731, i_4967, i_6225);
  nand ginst2373 (i_6732, i_4964, i_6226);
  nand ginst2374 (i_6733, i_4988, i_6227);
  nand ginst2375 (i_6734, i_4985, i_6228);
  nand ginst2376 (i_6735, i_4994, i_6229);
  nand ginst2377 (i_6736, i_4991, i_6230);
  not ginst2378 (i_674, i_106);
  nand ginst2379 (i_6741, i_5055, i_6239);
  nand ginst2380 (i_6742, i_5052, i_6240);
  nand ginst2381 (i_6743, i_5061, i_6241);
  nand ginst2382 (i_6744, i_5058, i_6242);
  nand ginst2383 (i_6751, i_5129, i_6255);
  nand ginst2384 (i_6752, i_5126, i_6256);
  nand ginst2385 (i_6753, i_5135, i_6257);
  nand ginst2386 (i_6754, i_5132, i_6258);
  nand ginst2387 (i_6755, i_5156, i_6259);
  nand ginst2388 (i_6756, i_5153, i_6260);
  nand ginst2389 (i_6757, i_5162, i_6261);
  nand ginst2390 (i_6758, i_5159, i_6262);
  not ginst2391 (i_676, i_18);
  not ginst2392 (i_6761, i_5892);
  and ginst2393 (i_6762, i_5632, i_5640, i_5654, i_5670, i_5683);
  and ginst2394 (i_6766, i_3097, i_5632);
  and ginst2395 (i_6767, i_3101, i_5632, i_5640);
  and ginst2396 (i_6768, i_3107, i_5632, i_5640, i_5654);
  and ginst2397 (i_6769, i_3114, i_5632, i_5640, i_5654, i_5670);
  and ginst2398 (i_6770, i_3101, i_5640);
  and ginst2399 (i_6771, i_3107, i_5640, i_5654);
  and ginst2400 (i_6772, i_3114, i_5640, i_5654, i_5670);
  and ginst2401 (i_6773, i_5640, i_5654, i_5670, i_5683);
  and ginst2402 (i_6774, i_3101, i_5640);
  and ginst2403 (i_6775, i_3107, i_5640, i_5654);
  and ginst2404 (i_6776, i_3114, i_5640, i_5654, i_5670);
  and ginst2405 (i_6777, i_3107, i_5654);
  and ginst2406 (i_6778, i_3114, i_5654, i_5670);
  and ginst2407 (i_6779, i_5654, i_5670, i_5683);
  and ginst2408 (i_6780, i_3107, i_5654);
  and ginst2409 (i_6781, i_3114, i_5654, i_5670);
  and ginst2410 (i_6782, i_3114, i_5670);
  and ginst2411 (i_6783, i_5670, i_5683);
  and ginst2412 (i_6784, i_5690, i_5697, i_5707, i_5718, i_5728);
  and ginst2413 (i_6787, i_3137, i_5690);
  and ginst2414 (i_6788, i_3140, i_5690, i_5697);
  and ginst2415 (i_6789, i_3144, i_5690, i_5697, i_5707);
  and ginst2416 (i_6790, i_3149, i_5690, i_5697, i_5707, i_5718);
  and ginst2417 (i_6791, i_3140, i_5697);
  and ginst2418 (i_6792, i_3144, i_5697, i_5707);
  and ginst2419 (i_6793, i_3149, i_5697, i_5707, i_5718);
  and ginst2420 (i_6794, i_3144, i_5707);
  and ginst2421 (i_6795, i_3149, i_5707, i_5718);
  and ginst2422 (i_6796, i_3149, i_5718);
  not ginst2423 (i_6797, i_5736);
  not ginst2424 (i_6800, i_5740);
  not ginst2425 (i_6803, i_5747);
  not ginst2426 (i_6806, i_5751);
  not ginst2427 (i_6809, i_5758);
  not ginst2428 (i_6812, i_5762);
  not ginst2429 (i_6815, i_5744);
  not ginst2430 (i_6818, i_5744);
  not ginst2431 (i_682, i_18);
  not ginst2432 (i_6821, i_5755);
  not ginst2433 (i_6824, i_5755);
  not ginst2434 (i_6827, i_5766);
  not ginst2435 (i_6830, i_5766);
  and ginst2436 (i_6833, i_5771, i_5778, i_5789, i_5850);
  and ginst2437 (i_6836, i_3169, i_5771);
  and ginst2438 (i_6837, i_3173, i_5771, i_5778);
  and ginst2439 (i_6838, i_3178, i_5771, i_5778, i_5789);
  and ginst2440 (i_6839, i_3173, i_5778);
  and ginst2441 (i_6840, i_3178, i_5778, i_5789);
  and ginst2442 (i_6841, i_5778, i_5789, i_5850);
  and ginst2443 (i_6842, i_3173, i_5778);
  and ginst2444 (i_6843, i_3178, i_5778, i_5789);
  and ginst2445 (i_6844, i_3178, i_5789);
  and ginst2446 (i_6845, i_5799, i_5807, i_5821, i_5837, i_5856);
  and ginst2447 (i_6848, i_3185, i_5799);
  and ginst2448 (i_6849, i_3189, i_5799, i_5807);
  and ginst2449 (i_6850, i_3195, i_5799, i_5807, i_5821);
  and ginst2450 (i_6851, i_3202, i_5799, i_5807, i_5821, i_5837);
  and ginst2451 (i_6852, i_3189, i_5807);
  and ginst2452 (i_6853, i_3195, i_5807, i_5821);
  and ginst2453 (i_6854, i_3202, i_5807, i_5821, i_5837);
  and ginst2454 (i_6855, i_5807, i_5821, i_5837, i_5856);
  and ginst2455 (i_6856, i_3189, i_5807);
  and ginst2456 (i_6857, i_3195, i_5807, i_5821);
  and ginst2457 (i_6858, i_3202, i_5807, i_5821, i_5837);
  and ginst2458 (i_6859, i_3195, i_5821);
  and ginst2459 (i_6860, i_3202, i_5821, i_5837);
  and ginst2460 (i_6861, i_5821, i_5837, i_5856);
  and ginst2461 (i_6862, i_3195, i_5821);
  and ginst2462 (i_6863, i_3202, i_5821, i_5837);
  and ginst2463 (i_6864, i_3202, i_5837);
  and ginst2464 (i_6865, i_5789, i_5850);
  and ginst2465 (i_6866, i_5837, i_5856);
  and ginst2466 (i_6867, i_5863, i_5870, i_5881, i_5892);
  and ginst2467 (i_6870, i_3211, i_5863);
  and ginst2468 (i_6871, i_3215, i_5863, i_5870);
  and ginst2469 (i_6872, i_3221, i_5863, i_5870, i_5881);
  and ginst2470 (i_6873, i_3215, i_5870);
  and ginst2471 (i_6874, i_3221, i_5870, i_5881);
  and ginst2472 (i_6875, i_5870, i_5881, i_5892);
  and ginst2473 (i_6876, i_3215, i_5870);
  and ginst2474 (i_6877, i_3221, i_5870, i_5881);
  and ginst2475 (i_6878, i_3221, i_5881);
  and ginst2476 (i_6879, i_5881, i_5892);
  and ginst2477 (i_688, i_263, i_382);
  and ginst2478 (i_6880, i_3221, i_5881);
  and ginst2479 (i_6881, i_5898, i_5905, i_5915, i_5926, i_5936);
  and ginst2480 (i_6884, i_3229, i_5898);
  and ginst2481 (i_6885, i_3232, i_5898, i_5905);
  and ginst2482 (i_6886, i_3236, i_5898, i_5905, i_5915);
  and ginst2483 (i_6887, i_3241, i_5898, i_5905, i_5915, i_5926);
  and ginst2484 (i_6888, i_3232, i_5905);
  and ginst2485 (i_6889, i_3236, i_5905, i_5915);
  not ginst2486 (i_689, i_18);
  and ginst2487 (i_6890, i_3241, i_5905, i_5915, i_5926);
  and ginst2488 (i_6891, i_3236, i_5915);
  and ginst2489 (i_6892, i_3241, i_5915, i_5926);
  and ginst2490 (i_6893, i_3241, i_5926);
  nand ginst2491 (i_6894, i_5944, i_6540);
  nand ginst2492 (i_6901, i_5946, i_6541);
  nand ginst2493 (i_6912, i_5948, i_6542);
  nand ginst2494 (i_6923, i_5950, i_6543);
  nand ginst2495 (i_6929, i_5952, i_6544);
  nand ginst2496 (i_6936, i_5954, i_6545);
  nand ginst2497 (i_6946, i_5956, i_6546);
  not ginst2498 (i_695, i_18);
  nand ginst2499 (i_6957, i_5958, i_6547);
  nand ginst2500 (i_6967, i_4575, i_6204);
  not ginst2501 (i_6968, i_6204);
  not ginst2502 (i_6969, i_6207);
  nand ginst2503 (i_6970, i_5967, i_6555);
  nand ginst2504 (i_6977, i_5969, i_6556);
  nand ginst2505 (i_6988, i_5971, i_6557);
  nand ginst2506 (i_6998, i_5973, i_6558);
  nand ginst2507 (i_700, i_267, i_382);
  nand ginst2508 (i_7006, i_5975, i_6559);
  nand ginst2509 (i_7020, i_5977, i_6560);
  nand ginst2510 (i_7036, i_5979, i_6561);
  nand ginst2511 (i_7049, i_5989, i_6569);
  not ginst2512 (i_705, i_271);
  nand ginst2513 (i_7055, i_4610, i_6210);
  not ginst2514 (i_7056, i_6210);
  and ginst2515 (i_7057, i_5991, i_5996, i_6000, i_6021);
  not ginst2516 (i_706, i_274);
  and ginst2517 (i_7060, i_3362, i_5991);
  and ginst2518 (i_7061, i_3363, i_5991, i_5996);
  and ginst2519 (i_7062, i_3364, i_5991, i_5996, i_6000);
  and ginst2520 (i_7063, i_6003, i_6009, i_6014, i_6018, i_6022);
  and ginst2521 (i_7064, i_3366, i_6003);
  and ginst2522 (i_7065, i_3367, i_6003, i_6009);
  and ginst2523 (i_7066, i_3368, i_6003, i_6009, i_6014);
  and ginst2524 (i_7067, i_3369, i_6003, i_6009, i_6014, i_6018);
  nand ginst2525 (i_7068, i_6024, i_6594);
  not ginst2526 (i_707, i_277);
  nand ginst2527 (i_7073, i_6026, i_6595);
  nand ginst2528 (i_7077, i_6028, i_6596);
  not ginst2529 (i_708, i_277);
  nand ginst2530 (i_7080, i_6030, i_6597);
  nand ginst2531 (i_7086, i_6598, i_6599);
  nand ginst2532 (i_7091, i_6600, i_6601);
  nand ginst2533 (i_7095, i_6602, i_6603);
  nand ginst2534 (i_7098, i_6038, i_6604);
  nand ginst2535 (i_7099, i_6605, i_6606);
  and ginst2536 (i_7100, i_6041, i_6047, i_6052, i_6056, i_6059);
  and ginst2537 (i_7103, i_3371, i_6041);
  and ginst2538 (i_7104, i_3372, i_6041, i_6047);
  and ginst2539 (i_7105, i_3373, i_6041, i_6047, i_6052);
  and ginst2540 (i_7106, i_3374, i_6041, i_6047, i_6052, i_6056);
  nand ginst2541 (i_7107, i_6060, i_6621);
  nand ginst2542 (i_7114, i_6062, i_6622);
  nand ginst2543 (i_7125, i_6064, i_6623);
  nand ginst2544 (i_7136, i_6066, i_6624);
  nand ginst2545 (i_7142, i_6068, i_6625);
  nand ginst2546 (i_7149, i_6070, i_6626);
  not ginst2547 (i_715, i_280);
  nand ginst2548 (i_7159, i_6072, i_6627);
  nand ginst2549 (i_7170, i_6074, i_6628);
  nand ginst2550 (i_7180, i_6076, i_6629);
  not ginst2551 (i_7187, i_6220);
  not ginst2552 (i_7188, i_6079);
  not ginst2553 (i_7191, i_6083);
  nand ginst2554 (i_7194, i_6091, i_6639);
  nand ginst2555 (i_7198, i_6640, i_6641);
  nand ginst2556 (i_7202, i_6642, i_6643);
  nand ginst2557 (i_7205, i_6097, i_6644);
  nand ginst2558 (i_7209, i_6645, i_6646);
  not ginst2559 (i_721, i_283);
  nand ginst2560 (i_7213, i_6647, i_6648);
  not ginst2561 (i_7216, i_6087);
  not ginst2562 (i_7219, i_6087);
  nand ginst2563 (i_7222, i_6103, i_6649);
  nand ginst2564 (i_7229, i_6105, i_6650);
  nand ginst2565 (i_7240, i_6107, i_6651);
  nand ginst2566 (i_7250, i_6109, i_6652);
  nand ginst2567 (i_7258, i_6111, i_6653);
  not ginst2568 (i_727, i_286);
  nand ginst2569 (i_7272, i_6113, i_6654);
  nand ginst2570 (i_7288, i_6115, i_6655);
  nand ginst2571 (i_7301, i_6117, i_6656);
  nand ginst2572 (i_7307, i_6119, i_6657);
  nand ginst2573 (i_7314, i_6122, i_6658);
  nand ginst2574 (i_7318, i_6659, i_6660);
  nand ginst2575 (i_7322, i_6125, i_6661);
  not ginst2576 (i_7325, i_6127);
  not ginst2577 (i_7328, i_6131);
  not ginst2578 (i_733, i_289);
  nand ginst2579 (i_7331, i_6136, i_6668);
  not ginst2580 (i_7334, i_6137);
  not ginst2581 (i_7337, i_6141);
  not ginst2582 (i_734, i_293);
  not ginst2583 (i_7340, i_6145);
  not ginst2584 (i_7343, i_6145);
  nand ginst2585 (i_7346, i_6677, i_6678);
  nand ginst2586 (i_7351, i_6679, i_6680);
  nand ginst2587 (i_7355, i_6681, i_6682);
  nand ginst2588 (i_7358, i_6683, i_6684);
  nand ginst2589 (i_7364, i_6157, i_6685);
  nand ginst2590 (i_7369, i_6159, i_6686);
  nand ginst2591 (i_7373, i_6161, i_6687);
  nand ginst2592 (i_7376, i_6688, i_6689);
  nand ginst2593 (i_7377, i_6164, i_6690);
  not ginst2594 (i_7378, i_6166);
  not ginst2595 (i_7381, i_6170);
  not ginst2596 (i_7384, i_6177);
  nand ginst2597 (i_7387, i_6702, i_6703);
  nand ginst2598 (i_7391, i_6704, i_6705);
  nand ginst2599 (i_7394, i_6186, i_6706);
  nand ginst2600 (i_7398, i_6707, i_6708);
  nand ginst2601 (i_7402, i_6709, i_6710);
  not ginst2602 (i_7405, i_6174);
  not ginst2603 (i_7408, i_6174);
  not ginst2604 (i_7411, i_5936);
  not ginst2605 (i_7414, i_5898);
  not ginst2606 (i_7417, i_5905);
  not ginst2607 (i_742, i_296);
  not ginst2608 (i_7420, i_5915);
  not ginst2609 (i_7423, i_5926);
  not ginst2610 (i_7426, i_5728);
  not ginst2611 (i_7429, i_5690);
  not ginst2612 (i_7432, i_5697);
  not ginst2613 (i_7435, i_5707);
  not ginst2614 (i_7438, i_5718);
  nand ginst2615 (i_7441, i_6192, i_6711);
  nand ginst2616 (i_7444, i_6194, i_6712);
  not ginst2617 (i_7447, i_5683);
  not ginst2618 (i_7450, i_5670);
  not ginst2619 (i_7453, i_5632);
  not ginst2620 (i_7456, i_5654);
  not ginst2621 (i_7459, i_5640);
  not ginst2622 (i_7462, i_5640);
  not ginst2623 (i_7465, i_5683);
  not ginst2624 (i_7468, i_5670);
  not ginst2625 (i_7471, i_5632);
  not ginst2626 (i_7474, i_5654);
  not ginst2627 (i_7477, i_6196);
  not ginst2628 (i_7478, i_6199);
  not ginst2629 (i_7479, i_5850);
  not ginst2630 (i_748, i_299);
  not ginst2631 (i_7482, i_5789);
  not ginst2632 (i_7485, i_5771);
  not ginst2633 (i_7488, i_5778);
  not ginst2634 (i_749, i_303);
  not ginst2635 (i_7491, i_5850);
  not ginst2636 (i_7494, i_5789);
  not ginst2637 (i_7497, i_5771);
  not ginst2638 (i_750, i_367);
  not ginst2639 (i_7500, i_5778);
  not ginst2640 (i_7503, i_5856);
  not ginst2641 (i_7506, i_5837);
  not ginst2642 (i_7509, i_5799);
  not ginst2643 (i_7512, i_5821);
  not ginst2644 (i_7515, i_5807);
  not ginst2645 (i_7518, i_5807);
  not ginst2646 (i_7521, i_5856);
  not ginst2647 (i_7524, i_5837);
  not ginst2648 (i_7527, i_5799);
  not ginst2649 (i_7530, i_5821);
  not ginst2650 (i_7533, i_5863);
  not ginst2651 (i_7536, i_5863);
  not ginst2652 (i_7539, i_5870);
  not ginst2653 (i_7542, i_5870);
  not ginst2654 (i_7545, i_5881);
  not ginst2655 (i_7548, i_5881);
  not ginst2656 (i_7551, i_6214);
  not ginst2657 (i_7552, i_6217);
  not ginst2658 (i_7553, i_5981);
  not ginst2659 (i_7556, i_6249);
  not ginst2660 (i_7557, i_6252);
  not ginst2661 (i_7558, i_6243);
  not ginst2662 (i_7559, i_6246);
  nand ginst2663 (i_7560, i_6731, i_6732);
  nand ginst2664 (i_7563, i_6729, i_6730);
  nand ginst2665 (i_7566, i_6735, i_6736);
  nand ginst2666 (i_7569, i_6733, i_6734);
  not ginst2667 (i_7572, i_6232);
  not ginst2668 (i_7573, i_6236);
  nand ginst2669 (i_7574, i_6743, i_6744);
  nand ginst2670 (i_7577, i_6741, i_6742);
  not ginst2671 (i_758, i_307);
  not ginst2672 (i_7580, i_6263);
  not ginst2673 (i_7581, i_6266);
  nand ginst2674 (i_7582, i_6753, i_6754);
  nand ginst2675 (i_7585, i_6751, i_6752);
  nand ginst2676 (i_7588, i_6757, i_6758);
  not ginst2677 (i_759, i_310);
  nand ginst2678 (i_7591, i_6755, i_6756);
  or ginst2679 (i_7609, i_3096, i_6766, i_6767, i_6768, i_6769);
  or ginst2680 (i_7613, i_3107, i_6782);
  not ginst2681 (i_762, i_313);
  or ginst2682 (i_7620, i_3136, i_6787, i_6788, i_6789, i_6790);
  or ginst2683 (i_7649, i_3168, i_6836, i_6837, i_6838);
  or ginst2684 (i_7650, i_3173, i_6844);
  or ginst2685 (i_7655, i_3184, i_6848, i_6849, i_6850, i_6851);
  or ginst2686 (i_7659, i_3195, i_6864);
  or ginst2687 (i_7668, i_3210, i_6870, i_6871, i_6872);
  or ginst2688 (i_7671, i_3228, i_6884, i_6885, i_6886, i_6887);
  not ginst2689 (i_768, i_316);
  not ginst2690 (i_774, i_319);
  nand ginst2691 (i_7744, i_3661, i_6968);
  not ginst2692 (i_780, i_322);
  nand ginst2693 (i_7822, i_3664, i_7056);
  or ginst2694 (i_7825, i_3361, i_7060, i_7061, i_7062);
  or ginst2695 (i_7826, i_3365, i_7064, i_7065, i_7066, i_7067);
  or ginst2696 (i_7852, i_3370, i_7103, i_7104, i_7105, i_7106);
  not ginst2697 (i_786, i_325);
  not ginst2698 (i_794, i_328);
  not ginst2699 (i_800, i_331);
  not ginst2700 (i_806, i_334);
  or ginst2701 (i_8114, i_3101, i_6777, i_6778, i_6779);
  or ginst2702 (i_8117, i_3097, i_6770, i_6771, i_6772, i_6773);
  not ginst2703 (i_812, i_337);
  not ginst2704 (i_813, i_340);
  nor ginst2705 (i_8131, i_3101, i_6780, i_6781);
  nor ginst2706 (i_8134, i_3097, i_6774, i_6775, i_6776);
  not ginst2707 (i_814, i_340);
  nand ginst2708 (i_8144, i_6199, i_7477);
  nand ginst2709 (i_8145, i_6196, i_7478);
  or ginst2710 (i_8146, i_3169, i_6839, i_6840, i_6841);
  nor ginst2711 (i_8156, i_3169, i_6842, i_6843);
  or ginst2712 (i_8166, i_3189, i_6859, i_6860, i_6861);
  or ginst2713 (i_8169, i_3185, i_6852, i_6853, i_6854, i_6855);
  nor ginst2714 (i_8183, i_3189, i_6862, i_6863);
  nor ginst2715 (i_8186, i_3185, i_6856, i_6857, i_6858);
  or ginst2716 (i_8196, i_3211, i_6873, i_6874, i_6875);
  nor ginst2717 (i_8200, i_3211, i_6876, i_6877);
  or ginst2718 (i_8204, i_3215, i_6878, i_6879);
  nor ginst2719 (i_8208, i_3215, i_6880);
  not ginst2720 (i_821, i_343);
  nand ginst2721 (i_8216, i_6252, i_7556);
  nand ginst2722 (i_8217, i_6249, i_7557);
  nand ginst2723 (i_8218, i_6246, i_7558);
  nand ginst2724 (i_8219, i_6243, i_7559);
  nand ginst2725 (i_8232, i_6266, i_7580);
  nand ginst2726 (i_8233, i_6263, i_7581);
  not ginst2727 (i_8242, i_7411);
  not ginst2728 (i_8243, i_7414);
  not ginst2729 (i_8244, i_7417);
  not ginst2730 (i_8245, i_7420);
  not ginst2731 (i_8246, i_7423);
  not ginst2732 (i_8247, i_7426);
  not ginst2733 (i_8248, i_7429);
  not ginst2734 (i_8249, i_7432);
  not ginst2735 (i_8250, i_7435);
  not ginst2736 (i_8251, i_7438);
  not ginst2737 (i_8252, i_7136);
  not ginst2738 (i_8253, i_6923);
  not ginst2739 (i_8254, i_6762);
  not ginst2740 (i_8260, i_7459);
  not ginst2741 (i_8261, i_7462);
  and ginst2742 (i_8262, i_3122, i_6762);
  and ginst2743 (i_8269, i_3155, i_6784);
  not ginst2744 (i_827, i_346);
  not ginst2745 (i_8274, i_6815);
  not ginst2746 (i_8275, i_6818);
  not ginst2747 (i_8276, i_6821);
  not ginst2748 (i_8277, i_6824);
  not ginst2749 (i_8278, i_6827);
  not ginst2750 (i_8279, i_6830);
  and ginst2751 (i_8280, i_5736, i_5740, i_6815);
  and ginst2752 (i_8281, i_6797, i_6800, i_6818);
  and ginst2753 (i_8282, i_5747, i_5751, i_6821);
  and ginst2754 (i_8283, i_6803, i_6806, i_6824);
  and ginst2755 (i_8284, i_5758, i_5762, i_6827);
  and ginst2756 (i_8285, i_6809, i_6812, i_6830);
  not ginst2757 (i_8288, i_6845);
  not ginst2758 (i_8294, i_7488);
  not ginst2759 (i_8295, i_7500);
  not ginst2760 (i_8296, i_7515);
  not ginst2761 (i_8297, i_7518);
  and ginst2762 (i_8298, i_6833, i_6845);
  and ginst2763 (i_8307, i_6867, i_6881);
  not ginst2764 (i_8315, i_7533);
  not ginst2765 (i_8317, i_7536);
  not ginst2766 (i_8319, i_7539);
  not ginst2767 (i_8321, i_7542);
  nand ginst2768 (i_8322, i_4543, i_7545);
  not ginst2769 (i_8323, i_7545);
  nand ginst2770 (i_8324, i_5943, i_7548);
  not ginst2771 (i_8325, i_7548);
  nand ginst2772 (i_8326, i_6967, i_7744);
  not ginst2773 (i_833, i_349);
  and ginst2774 (i_8333, i_6894, i_6901, i_6912, i_6923);
  and ginst2775 (i_8337, i_4545, i_6894);
  and ginst2776 (i_8338, i_4549, i_6894, i_6901);
  and ginst2777 (i_8339, i_4555, i_6894, i_6901, i_6912);
  and ginst2778 (i_8340, i_4549, i_6901);
  and ginst2779 (i_8341, i_4555, i_6901, i_6912);
  and ginst2780 (i_8342, i_6901, i_6912, i_6923);
  and ginst2781 (i_8343, i_4549, i_6901);
  and ginst2782 (i_8344, i_4555, i_6901, i_6912);
  and ginst2783 (i_8345, i_4555, i_6912);
  and ginst2784 (i_8346, i_6912, i_6923);
  and ginst2785 (i_8347, i_4555, i_6912);
  and ginst2786 (i_8348, i_4563, i_6929);
  and ginst2787 (i_8349, i_4566, i_6929, i_6936);
  and ginst2788 (i_8350, i_4570, i_6929, i_6936, i_6946);
  and ginst2789 (i_8351, i_5960, i_6929, i_6936, i_6946, i_6957);
  and ginst2790 (i_8352, i_4566, i_6936);
  and ginst2791 (i_8353, i_4570, i_6936, i_6946);
  and ginst2792 (i_8354, i_5960, i_6936, i_6946, i_6957);
  and ginst2793 (i_8355, i_4570, i_6946);
  and ginst2794 (i_8356, i_5960, i_6946, i_6957);
  and ginst2795 (i_8357, i_5960, i_6957);
  nand ginst2796 (i_8358, i_7055, i_7822);
  and ginst2797 (i_8365, i_6970, i_6977, i_6988, i_7049);
  and ginst2798 (i_8369, i_4577, i_6970);
  and ginst2799 (i_8370, i_4581, i_6970, i_6977);
  and ginst2800 (i_8371, i_4586, i_6970, i_6977, i_6988);
  and ginst2801 (i_8372, i_4581, i_6977);
  and ginst2802 (i_8373, i_4586, i_6977, i_6988);
  and ginst2803 (i_8374, i_6977, i_6988, i_7049);
  and ginst2804 (i_8375, i_4581, i_6977);
  and ginst2805 (i_8376, i_4586, i_6977, i_6988);
  and ginst2806 (i_8377, i_4586, i_6988);
  and ginst2807 (i_8378, i_4593, i_6998);
  and ginst2808 (i_8379, i_4597, i_6998, i_7006);
  and ginst2809 (i_8380, i_4603, i_6998, i_7006, i_7020);
  and ginst2810 (i_8381, i_5981, i_6998, i_7006, i_7020, i_7036);
  and ginst2811 (i_8382, i_4597, i_7006);
  and ginst2812 (i_8383, i_4603, i_7006, i_7020);
  and ginst2813 (i_8384, i_5981, i_7006, i_7020, i_7036);
  and ginst2814 (i_8385, i_4597, i_7006);
  and ginst2815 (i_8386, i_4603, i_7006, i_7020);
  and ginst2816 (i_8387, i_5981, i_7006, i_7020, i_7036);
  and ginst2817 (i_8388, i_4603, i_7020);
  and ginst2818 (i_8389, i_5981, i_7020, i_7036);
  not ginst2819 (i_839, i_352);
  and ginst2820 (i_8390, i_4603, i_7020);
  and ginst2821 (i_8391, i_5981, i_7020, i_7036);
  and ginst2822 (i_8392, i_5981, i_7036);
  and ginst2823 (i_8393, i_6988, i_7049);
  and ginst2824 (i_8394, i_7057, i_7063);
  and ginst2825 (i_8404, i_7057, i_7826);
  and ginst2826 (i_8405, i_7068, i_7073, i_7077, i_7098);
  and ginst2827 (i_8409, i_4632, i_7068);
  and ginst2828 (i_8410, i_4634, i_7068, i_7073);
  and ginst2829 (i_8411, i_4635, i_7068, i_7073, i_7077);
  and ginst2830 (i_8412, i_7080, i_7086, i_7091, i_7095, i_7099);
  and ginst2831 (i_8415, i_4638, i_7080);
  and ginst2832 (i_8416, i_4639, i_7080, i_7086);
  and ginst2833 (i_8417, i_4640, i_7080, i_7086, i_7091);
  and ginst2834 (i_8418, i_4641, i_7080, i_7086, i_7091, i_7095);
  and ginst2835 (i_8421, i_3375, i_7100);
  and ginst2836 (i_8430, i_7107, i_7114, i_7125, i_7136);
  and ginst2837 (i_8433, i_4657, i_7107);
  and ginst2838 (i_8434, i_4661, i_7107, i_7114);
  and ginst2839 (i_8435, i_4667, i_7107, i_7114, i_7125);
  and ginst2840 (i_8436, i_4661, i_7114);
  and ginst2841 (i_8437, i_4667, i_7114, i_7125);
  and ginst2842 (i_8438, i_7114, i_7125, i_7136);
  and ginst2843 (i_8439, i_4661, i_7114);
  and ginst2844 (i_8440, i_4667, i_7114, i_7125);
  and ginst2845 (i_8441, i_4667, i_7125);
  and ginst2846 (i_8442, i_7125, i_7136);
  and ginst2847 (i_8443, i_4667, i_7125);
  and ginst2848 (i_8444, i_7142, i_7149, i_7159, i_7170, i_7180);
  and ginst2849 (i_8447, i_4675, i_7142);
  and ginst2850 (i_8448, i_4678, i_7142, i_7149);
  and ginst2851 (i_8449, i_4682, i_7142, i_7149, i_7159);
  not ginst2852 (i_845, i_355);
  and ginst2853 (i_8450, i_4687, i_7142, i_7149, i_7159, i_7170);
  and ginst2854 (i_8451, i_4678, i_7149);
  and ginst2855 (i_8452, i_4682, i_7149, i_7159);
  and ginst2856 (i_8453, i_4687, i_7149, i_7159, i_7170);
  and ginst2857 (i_8454, i_4682, i_7159);
  and ginst2858 (i_8455, i_4687, i_7159, i_7170);
  and ginst2859 (i_8456, i_4687, i_7170);
  not ginst2860 (i_8457, i_7194);
  not ginst2861 (i_8460, i_7198);
  not ginst2862 (i_8463, i_7205);
  not ginst2863 (i_8466, i_7209);
  not ginst2864 (i_8469, i_7216);
  not ginst2865 (i_8470, i_7219);
  not ginst2866 (i_8471, i_7202);
  not ginst2867 (i_8474, i_7202);
  not ginst2868 (i_8477, i_7213);
  not ginst2869 (i_8480, i_7213);
  and ginst2870 (i_8483, i_6079, i_6083, i_7216);
  and ginst2871 (i_8484, i_7188, i_7191, i_7219);
  and ginst2872 (i_8485, i_7222, i_7229, i_7240, i_7301);
  and ginst2873 (i_8488, i_4702, i_7222);
  and ginst2874 (i_8489, i_4706, i_7222, i_7229);
  and ginst2875 (i_8490, i_4711, i_7222, i_7229, i_7240);
  and ginst2876 (i_8491, i_4706, i_7229);
  and ginst2877 (i_8492, i_4711, i_7229, i_7240);
  and ginst2878 (i_8493, i_7229, i_7240, i_7301);
  and ginst2879 (i_8494, i_4706, i_7229);
  and ginst2880 (i_8495, i_4711, i_7229, i_7240);
  and ginst2881 (i_8496, i_4711, i_7240);
  and ginst2882 (i_8497, i_7250, i_7258, i_7272, i_7288, i_7307);
  and ginst2883 (i_8500, i_4718, i_7250);
  and ginst2884 (i_8501, i_4722, i_7250, i_7258);
  and ginst2885 (i_8502, i_4728, i_7250, i_7258, i_7272);
  and ginst2886 (i_8503, i_4735, i_7250, i_7258, i_7272, i_7288);
  and ginst2887 (i_8504, i_4722, i_7258);
  and ginst2888 (i_8505, i_4728, i_7258, i_7272);
  and ginst2889 (i_8506, i_4735, i_7258, i_7272, i_7288);
  and ginst2890 (i_8507, i_7258, i_7272, i_7288, i_7307);
  and ginst2891 (i_8508, i_4722, i_7258);
  and ginst2892 (i_8509, i_4728, i_7258, i_7272);
  and ginst2893 (i_8510, i_4735, i_7258, i_7272, i_7288);
  and ginst2894 (i_8511, i_4728, i_7272);
  and ginst2895 (i_8512, i_4735, i_7272, i_7288);
  and ginst2896 (i_8513, i_7272, i_7288, i_7307);
  and ginst2897 (i_8514, i_4728, i_7272);
  and ginst2898 (i_8515, i_4735, i_7272, i_7288);
  and ginst2899 (i_8516, i_4735, i_7288);
  and ginst2900 (i_8517, i_7240, i_7301);
  and ginst2901 (i_8518, i_7288, i_7307);
  not ginst2902 (i_8519, i_7314);
  not ginst2903 (i_8522, i_7318);
  not ginst2904 (i_8525, i_7322);
  not ginst2905 (i_8528, i_7322);
  not ginst2906 (i_853, i_358);
  not ginst2907 (i_8531, i_7331);
  not ginst2908 (i_8534, i_7331);
  not ginst2909 (i_8537, i_7340);
  not ginst2910 (i_8538, i_7343);
  and ginst2911 (i_8539, i_6137, i_6141, i_7340);
  and ginst2912 (i_8540, i_7334, i_7337, i_7343);
  and ginst2913 (i_8541, i_7346, i_7351, i_7355, i_7376);
  and ginst2914 (i_8545, i_4757, i_7346);
  and ginst2915 (i_8546, i_4758, i_7346, i_7351);
  and ginst2916 (i_8547, i_4759, i_7346, i_7351, i_7355);
  and ginst2917 (i_8548, i_7358, i_7364, i_7369, i_7373, i_7377);
  and ginst2918 (i_8551, i_4762, i_7358);
  and ginst2919 (i_8552, i_4764, i_7358, i_7364);
  and ginst2920 (i_8553, i_4766, i_7358, i_7364, i_7369);
  and ginst2921 (i_8554, i_4767, i_7358, i_7364, i_7369, i_7373);
  not ginst2922 (i_8555, i_7387);
  not ginst2923 (i_8558, i_7394);
  not ginst2924 (i_8561, i_7398);
  not ginst2925 (i_8564, i_7405);
  not ginst2926 (i_8565, i_7408);
  not ginst2927 (i_8566, i_7391);
  not ginst2928 (i_8569, i_7391);
  not ginst2929 (i_8572, i_7402);
  not ginst2930 (i_8575, i_7402);
  and ginst2931 (i_8578, i_6166, i_6170, i_7405);
  and ginst2932 (i_8579, i_7378, i_7381, i_7408);
  not ginst2933 (i_8580, i_7180);
  not ginst2934 (i_8583, i_7142);
  not ginst2935 (i_8586, i_7149);
  not ginst2936 (i_8589, i_7159);
  not ginst2937 (i_859, i_361);
  not ginst2938 (i_8592, i_7170);
  not ginst2939 (i_8595, i_6929);
  not ginst2940 (i_8598, i_6936);
  not ginst2941 (i_8601, i_6946);
  not ginst2942 (i_8604, i_6957);
  not ginst2943 (i_8607, i_7441);
  nand ginst2944 (i_8608, i_5469, i_7441);
  not ginst2945 (i_8609, i_7444);
  nand ginst2946 (i_8610, i_4793, i_7444);
  not ginst2947 (i_8615, i_7447);
  not ginst2948 (i_8616, i_7450);
  not ginst2949 (i_8617, i_7453);
  not ginst2950 (i_8618, i_7456);
  not ginst2951 (i_8619, i_7474);
  not ginst2952 (i_8624, i_7465);
  not ginst2953 (i_8625, i_7468);
  not ginst2954 (i_8626, i_7471);
  nand ginst2955 (i_8627, i_8144, i_8145);
  not ginst2956 (i_8632, i_7479);
  not ginst2957 (i_8633, i_7482);
  not ginst2958 (i_8634, i_7485);
  not ginst2959 (i_8637, i_7491);
  not ginst2960 (i_8638, i_7494);
  not ginst2961 (i_8639, i_7497);
  not ginst2962 (i_8644, i_7503);
  not ginst2963 (i_8645, i_7506);
  not ginst2964 (i_8646, i_7509);
  not ginst2965 (i_8647, i_7512);
  not ginst2966 (i_8648, i_7530);
  not ginst2967 (i_865, i_364);
  not ginst2968 (i_8653, i_7521);
  not ginst2969 (i_8654, i_7524);
  not ginst2970 (i_8655, i_7527);
  not ginst2971 (i_8660, i_6894);
  not ginst2972 (i_8663, i_6894);
  not ginst2973 (i_8666, i_6901);
  not ginst2974 (i_8669, i_6901);
  not ginst2975 (i_8672, i_6912);
  not ginst2976 (i_8675, i_6912);
  not ginst2977 (i_8678, i_7049);
  not ginst2978 (i_8681, i_6988);
  not ginst2979 (i_8684, i_6970);
  not ginst2980 (i_8687, i_6977);
  not ginst2981 (i_8690, i_7049);
  not ginst2982 (i_8693, i_6988);
  not ginst2983 (i_8696, i_6970);
  not ginst2984 (i_8699, i_6977);
  not ginst2985 (i_8702, i_7036);
  not ginst2986 (i_8705, i_6998);
  not ginst2987 (i_8708, i_7020);
  not ginst2988 (i_871, i_367);
  not ginst2989 (i_8711, i_7006);
  not ginst2990 (i_8714, i_7006);
  not ginst2991 (i_8717, i_7553);
  not ginst2992 (i_8718, i_7036);
  not ginst2993 (i_8721, i_6998);
  not ginst2994 (i_8724, i_7020);
  nand ginst2995 (i_8727, i_8216, i_8217);
  nand ginst2996 (i_8730, i_8218, i_8219);
  not ginst2997 (i_8733, i_7574);
  not ginst2998 (i_8734, i_7577);
  not ginst2999 (i_8735, i_7107);
  not ginst3000 (i_8738, i_7107);
  not ginst3001 (i_8741, i_7114);
  not ginst3002 (i_8744, i_7114);
  not ginst3003 (i_8747, i_7125);
  not ginst3004 (i_8750, i_7125);
  not ginst3005 (i_8753, i_7560);
  not ginst3006 (i_8754, i_7563);
  not ginst3007 (i_8755, i_7566);
  not ginst3008 (i_8756, i_7569);
  not ginst3009 (i_8757, i_7301);
  not ginst3010 (i_8760, i_7240);
  not ginst3011 (i_8763, i_7222);
  not ginst3012 (i_8766, i_7229);
  not ginst3013 (i_8769, i_7301);
  not ginst3014 (i_8772, i_7240);
  not ginst3015 (i_8775, i_7222);
  not ginst3016 (i_8778, i_7229);
  not ginst3017 (i_8781, i_7307);
  not ginst3018 (i_8784, i_7288);
  not ginst3019 (i_8787, i_7250);
  not ginst3020 (i_8790, i_7272);
  not ginst3021 (i_8793, i_7258);
  not ginst3022 (i_8796, i_7258);
  not ginst3023 (i_8799, i_7307);
  not ginst3024 (i_8802, i_7288);
  not ginst3025 (i_8805, i_7250);
  not ginst3026 (i_8808, i_7272);
  nand ginst3027 (i_881, i_467, i_585);
  nand ginst3028 (i_8811, i_8232, i_8233);
  not ginst3029 (i_8814, i_7588);
  not ginst3030 (i_8815, i_7591);
  not ginst3031 (i_8816, i_7582);
  not ginst3032 (i_8817, i_7585);
  and ginst3033 (i_8818, i_3155, i_7620);
  not ginst3034 (i_882, i_528);
  not ginst3035 (i_883, i_578);
  not ginst3036 (i_884, i_575);
  and ginst3037 (i_8840, i_3122, i_7609);
  not ginst3038 (i_885, i_494);
  not ginst3039 (i_8857, i_7609);
  and ginst3040 (i_886, i_528, i_578);
  and ginst3041 (i_8861, i_5740, i_6797, i_8274);
  and ginst3042 (i_8862, i_5736, i_6800, i_8275);
  and ginst3043 (i_8863, i_5751, i_6803, i_8276);
  and ginst3044 (i_8864, i_5747, i_6806, i_8277);
  and ginst3045 (i_8865, i_5762, i_6809, i_8278);
  and ginst3046 (i_8866, i_5758, i_6812, i_8279);
  and ginst3047 (i_887, i_494, i_575);
  not ginst3048 (i_8871, i_7655);
  and ginst3049 (i_8874, i_6833, i_7655);
  and ginst3050 (i_8878, i_6867, i_7671);
  not ginst3051 (i_8879, i_8196);
  nand ginst3052 (i_8880, i_8196, i_8315);
  not ginst3053 (i_8881, i_8200);
  nand ginst3054 (i_8882, i_8200, i_8317);
  not ginst3055 (i_8883, i_8204);
  nand ginst3056 (i_8884, i_8204, i_8319);
  not ginst3057 (i_8885, i_8208);
  nand ginst3058 (i_8886, i_8208, i_8321);
  nand ginst3059 (i_8887, i_3658, i_8323);
  nand ginst3060 (i_8888, i_4817, i_8325);
  not ginst3061 (i_889, i_590);
  or ginst3062 (i_8898, i_4544, i_8337, i_8338, i_8339);
  or ginst3063 (i_8902, i_4562, i_8348, i_8349, i_8350, i_8351);
  or ginst3064 (i_8920, i_4576, i_8369, i_8370, i_8371);
  or ginst3065 (i_8924, i_4581, i_8377);
  or ginst3066 (i_8927, i_4592, i_8378, i_8379, i_8380, i_8381);
  or ginst3067 (i_8931, i_4603, i_8392);
  or ginst3068 (i_8943, i_7825, i_8404);
  or ginst3069 (i_8950, i_4630, i_8409, i_8410, i_8411);
  or ginst3070 (i_8956, i_4637, i_8415, i_8416, i_8417, i_8418);
  not ginst3071 (i_8959, i_7852);
  and ginst3072 (i_8960, i_3375, i_7852);
  or ginst3073 (i_8963, i_4656, i_8433, i_8434, i_8435);
  or ginst3074 (i_8966, i_4674, i_8447, i_8448, i_8449, i_8450);
  and ginst3075 (i_8991, i_6083, i_7188, i_8469);
  and ginst3076 (i_8992, i_6079, i_7191, i_8470);
  or ginst3077 (i_8995, i_4701, i_8488, i_8489, i_8490);
  or ginst3078 (i_8996, i_4706, i_8496);
  or ginst3079 (i_9001, i_4717, i_8500, i_8501, i_8502, i_8503);
  or ginst3080 (i_9005, i_4728, i_8516);
  and ginst3081 (i_9024, i_6141, i_7334, i_8537);
  and ginst3082 (i_9025, i_6137, i_7337, i_8538);
  or ginst3083 (i_9029, i_4756, i_8545, i_8546, i_8547);
  or ginst3084 (i_9035, i_4760, i_8551, i_8552, i_8553, i_8554);
  and ginst3085 (i_9053, i_6170, i_7378, i_8564);
  and ginst3086 (i_9054, i_6166, i_7381, i_8565);
  nand ginst3087 (i_9064, i_4303, i_8607);
  nand ginst3088 (i_9065, i_3507, i_8609);
  not ginst3089 (i_9066, i_8114);
  nand ginst3090 (i_9067, i_4795, i_8114);
  or ginst3091 (i_9068, i_6783, i_7613);
  not ginst3092 (i_9071, i_8117);
  not ginst3093 (i_9072, i_8131);
  nand ginst3094 (i_9073, i_6195, i_8131);
  not ginst3095 (i_9074, i_7613);
  not ginst3096 (i_9077, i_8134);
  or ginst3097 (i_9079, i_6865, i_7650);
  not ginst3098 (i_9082, i_8146);
  not ginst3099 (i_9083, i_7650);
  not ginst3100 (i_9086, i_8156);
  not ginst3101 (i_9087, i_8166);
  nand ginst3102 (i_9088, i_4813, i_8166);
  or ginst3103 (i_9089, i_6866, i_7659);
  not ginst3104 (i_9092, i_8169);
  not ginst3105 (i_9093, i_8183);
  nand ginst3106 (i_9094, i_6203, i_8183);
  not ginst3107 (i_9095, i_7659);
  not ginst3108 (i_9098, i_8186);
  or ginst3109 (i_9099, i_4545, i_8340, i_8341, i_8342);
  nor ginst3110 (i_9103, i_4545, i_8343, i_8344);
  or ginst3111 (i_9107, i_4549, i_8345, i_8346);
  nor ginst3112 (i_9111, i_4549, i_8347);
  or ginst3113 (i_9117, i_4577, i_8372, i_8373, i_8374);
  nor ginst3114 (i_9127, i_4577, i_8375, i_8376);
  nor ginst3115 (i_9146, i_4597, i_8390, i_8391);
  nor ginst3116 (i_9149, i_4593, i_8385, i_8386, i_8387);
  nand ginst3117 (i_9159, i_7577, i_8733);
  nand ginst3118 (i_9160, i_7574, i_8734);
  or ginst3119 (i_9161, i_4657, i_8436, i_8437, i_8438);
  nor ginst3120 (i_9165, i_4657, i_8439, i_8440);
  or ginst3121 (i_9169, i_4661, i_8441, i_8442);
  nor ginst3122 (i_9173, i_4661, i_8443);
  nand ginst3123 (i_9179, i_7563, i_8753);
  nand ginst3124 (i_9180, i_7560, i_8754);
  nand ginst3125 (i_9181, i_7569, i_8755);
  nand ginst3126 (i_9182, i_7566, i_8756);
  or ginst3127 (i_9183, i_4702, i_8491, i_8492, i_8493);
  nor ginst3128 (i_9193, i_4702, i_8494, i_8495);
  or ginst3129 (i_9203, i_4722, i_8511, i_8512, i_8513);
  or ginst3130 (i_9206, i_4718, i_8504, i_8505, i_8506, i_8507);
  nor ginst3131 (i_9220, i_4722, i_8514, i_8515);
  nor ginst3132 (i_9223, i_4718, i_8508, i_8509, i_8510);
  nand ginst3133 (i_9234, i_7591, i_8814);
  nand ginst3134 (i_9235, i_7588, i_8815);
  nand ginst3135 (i_9236, i_7585, i_8816);
  nand ginst3136 (i_9237, i_7582, i_8817);
  or ginst3137 (i_9238, i_3159, i_8818);
  or ginst3138 (i_9242, i_3126, i_8840);
  nand ginst3139 (i_9243, i_8324, i_8888);
  not ginst3140 (i_9244, i_8580);
  not ginst3141 (i_9245, i_8583);
  not ginst3142 (i_9246, i_8586);
  not ginst3143 (i_9247, i_8589);
  not ginst3144 (i_9248, i_8592);
  not ginst3145 (i_9249, i_8595);
  not ginst3146 (i_9250, i_8598);
  not ginst3147 (i_9251, i_8601);
  not ginst3148 (i_9252, i_8604);
  nor ginst3149 (i_9256, i_8280, i_8861);
  nor ginst3150 (i_9257, i_8281, i_8862);
  nor ginst3151 (i_9258, i_8282, i_8863);
  nor ginst3152 (i_9259, i_8283, i_8864);
  nor ginst3153 (i_9260, i_8284, i_8865);
  nor ginst3154 (i_9261, i_8285, i_8866);
  not ginst3155 (i_9262, i_8627);
  or ginst3156 (i_9265, i_7649, i_8874);
  or ginst3157 (i_9268, i_7668, i_8878);
  nand ginst3158 (i_9271, i_7533, i_8879);
  nand ginst3159 (i_9272, i_7536, i_8881);
  nand ginst3160 (i_9273, i_7539, i_8883);
  nand ginst3161 (i_9274, i_7542, i_8885);
  nand ginst3162 (i_9275, i_8322, i_8887);
  not ginst3163 (i_9276, i_8333);
  and ginst3164 (i_9280, i_6929, i_6936, i_6946, i_6957, i_8326);
  and ginst3165 (i_9285, i_367, i_6936, i_6946, i_6957, i_8326);
  and ginst3166 (i_9286, i_367, i_6946, i_6957, i_8326);
  and ginst3167 (i_9287, i_367, i_6957, i_8326);
  and ginst3168 (i_9288, i_367, i_8326);
  not ginst3169 (i_9290, i_8660);
  not ginst3170 (i_9292, i_8663);
  not ginst3171 (i_9294, i_8666);
  not ginst3172 (i_9296, i_8669);
  nand ginst3173 (i_9297, i_5966, i_8672);
  not ginst3174 (i_9298, i_8672);
  nand ginst3175 (i_9299, i_6969, i_8675);
  not ginst3176 (i_9300, i_8675);
  not ginst3177 (i_9301, i_8365);
  and ginst3178 (i_9307, i_6998, i_7006, i_7020, i_7036, i_8358);
  and ginst3179 (i_9314, i_7006, i_7020, i_7036, i_8358);
  and ginst3180 (i_9315, i_7020, i_7036, i_8358);
  and ginst3181 (i_9318, i_7036, i_8358);
  not ginst3182 (i_9319, i_8687);
  not ginst3183 (i_9320, i_8699);
  not ginst3184 (i_9321, i_8711);
  not ginst3185 (i_9322, i_8714);
  not ginst3186 (i_9323, i_8727);
  not ginst3187 (i_9324, i_8730);
  not ginst3188 (i_9326, i_8405);
  and ginst3189 (i_9332, i_8405, i_8412);
  or ginst3190 (i_9339, i_4193, i_8960);
  and ginst3191 (i_9344, i_8430, i_8444);
  not ginst3192 (i_9352, i_8735);
  not ginst3193 (i_9354, i_8738);
  not ginst3194 (i_9356, i_8741);
  not ginst3195 (i_9358, i_8744);
  nand ginst3196 (i_9359, i_6078, i_8747);
  not ginst3197 (i_9360, i_8747);
  nand ginst3198 (i_9361, i_7187, i_8750);
  not ginst3199 (i_9362, i_8750);
  not ginst3200 (i_9363, i_8471);
  not ginst3201 (i_9364, i_8474);
  not ginst3202 (i_9365, i_8477);
  not ginst3203 (i_9366, i_8480);
  nor ginst3204 (i_9367, i_8483, i_8991);
  nor ginst3205 (i_9368, i_8484, i_8992);
  and ginst3206 (i_9369, i_7194, i_7198, i_8471);
  and ginst3207 (i_9370, i_8457, i_8460, i_8474);
  and ginst3208 (i_9371, i_7205, i_7209, i_8477);
  and ginst3209 (i_9372, i_8463, i_8466, i_8480);
  not ginst3210 (i_9375, i_8497);
  not ginst3211 (i_9381, i_8766);
  not ginst3212 (i_9382, i_8778);
  not ginst3213 (i_9383, i_8793);
  not ginst3214 (i_9384, i_8796);
  and ginst3215 (i_9385, i_8485, i_8497);
  not ginst3216 (i_9392, i_8525);
  not ginst3217 (i_9393, i_8528);
  not ginst3218 (i_9394, i_8531);
  not ginst3219 (i_9395, i_8534);
  and ginst3220 (i_9396, i_7314, i_7318, i_8525);
  and ginst3221 (i_9397, i_8519, i_8522, i_8528);
  and ginst3222 (i_9398, i_6127, i_6131, i_8531);
  and ginst3223 (i_9399, i_7325, i_7328, i_8534);
  nor ginst3224 (i_9400, i_8539, i_9024);
  nor ginst3225 (i_9401, i_8540, i_9025);
  not ginst3226 (i_9402, i_8541);
  nand ginst3227 (i_9407, i_89, i_8548);
  and ginst3228 (i_9408, i_8541, i_8548);
  not ginst3229 (i_9412, i_8811);
  not ginst3230 (i_9413, i_8566);
  not ginst3231 (i_9414, i_8569);
  not ginst3232 (i_9415, i_8572);
  not ginst3233 (i_9416, i_8575);
  nor ginst3234 (i_9417, i_8578, i_9053);
  nor ginst3235 (i_9418, i_8579, i_9054);
  and ginst3236 (i_9419, i_6177, i_7387, i_8566);
  and ginst3237 (i_9420, i_7384, i_8555, i_8569);
  and ginst3238 (i_9421, i_7394, i_7398, i_8572);
  and ginst3239 (i_9422, i_8558, i_8561, i_8575);
  not ginst3240 (i_9423, i_8326);
  nand ginst3241 (i_9426, i_8608, i_9064);
  nand ginst3242 (i_9429, i_8610, i_9065);
  nand ginst3243 (i_9432, i_3515, i_9066);
  nand ginst3244 (i_9435, i_4796, i_9072);
  nand ginst3245 (i_9442, i_3628, i_9087);
  nand ginst3246 (i_9445, i_4814, i_9093);
  not ginst3247 (i_945, i_657);
  not ginst3248 (i_9454, i_8678);
  not ginst3249 (i_9455, i_8681);
  not ginst3250 (i_9456, i_8684);
  not ginst3251 (i_9459, i_8690);
  not ginst3252 (i_9460, i_8693);
  not ginst3253 (i_9461, i_8696);
  not ginst3254 (i_9462, i_8358);
  not ginst3255 (i_9465, i_8702);
  not ginst3256 (i_9466, i_8705);
  not ginst3257 (i_9467, i_8708);
  not ginst3258 (i_9468, i_8724);
  not ginst3259 (i_9473, i_8358);
  not ginst3260 (i_9476, i_8718);
  not ginst3261 (i_9477, i_8721);
  nand ginst3262 (i_9478, i_9159, i_9160);
  nand ginst3263 (i_9485, i_9179, i_9180);
  nand ginst3264 (i_9488, i_9181, i_9182);
  not ginst3265 (i_9493, i_8757);
  not ginst3266 (i_9494, i_8760);
  not ginst3267 (i_9495, i_8763);
  not ginst3268 (i_9498, i_8769);
  not ginst3269 (i_9499, i_8772);
  not ginst3270 (i_9500, i_8775);
  not ginst3271 (i_9505, i_8781);
  not ginst3272 (i_9506, i_8784);
  not ginst3273 (i_9507, i_8787);
  not ginst3274 (i_9508, i_8790);
  not ginst3275 (i_9509, i_8808);
  not ginst3276 (i_9514, i_8799);
  not ginst3277 (i_9515, i_8802);
  not ginst3278 (i_9516, i_8805);
  nand ginst3279 (i_9517, i_9234, i_9235);
  nand ginst3280 (i_9520, i_9236, i_9237);
  and ginst3281 (i_9526, i_8421, i_8943);
  and ginst3282 (i_9531, i_8421, i_8943);
  nand ginst3283 (i_9539, i_8880, i_9271);
  nand ginst3284 (i_9540, i_8884, i_9273);
  not ginst3285 (i_9541, i_9275);
  and ginst3286 (i_9543, i_8254, i_8857);
  and ginst3287 (i_9551, i_8288, i_8871);
  nand ginst3288 (i_9555, i_8882, i_9272);
  nand ginst3289 (i_9556, i_8886, i_9274);
  not ginst3290 (i_9557, i_8898);
  and ginst3291 (i_9560, i_8333, i_8902);
  not ginst3292 (i_9561, i_9099);
  nand ginst3293 (i_9562, i_9099, i_9290);
  not ginst3294 (i_9563, i_9103);
  nand ginst3295 (i_9564, i_9103, i_9292);
  not ginst3296 (i_9565, i_9107);
  nand ginst3297 (i_9566, i_9107, i_9294);
  not ginst3298 (i_9567, i_9111);
  nand ginst3299 (i_9568, i_9111, i_9296);
  nand ginst3300 (i_9569, i_4844, i_9298);
  not ginst3301 (i_957, i_688);
  nand ginst3302 (i_9570, i_6207, i_9300);
  not ginst3303 (i_9571, i_8920);
  not ginst3304 (i_9575, i_8927);
  and ginst3305 (i_9579, i_8365, i_8927);
  not ginst3306 (i_9581, i_8950);
  not ginst3307 (i_9582, i_8956);
  and ginst3308 (i_9585, i_8405, i_8956);
  and ginst3309 (i_9591, i_8430, i_8966);
  not ginst3310 (i_9592, i_9161);
  nand ginst3311 (i_9593, i_9161, i_9352);
  not ginst3312 (i_9594, i_9165);
  nand ginst3313 (i_9595, i_9165, i_9354);
  not ginst3314 (i_9596, i_9169);
  nand ginst3315 (i_9597, i_9169, i_9356);
  not ginst3316 (i_9598, i_9173);
  nand ginst3317 (i_9599, i_9173, i_9358);
  nand ginst3318 (i_9600, i_4940, i_9360);
  nand ginst3319 (i_9601, i_6220, i_9362);
  and ginst3320 (i_9602, i_7198, i_8457, i_9363);
  and ginst3321 (i_9603, i_7194, i_8460, i_9364);
  and ginst3322 (i_9604, i_7209, i_8463, i_9365);
  and ginst3323 (i_9605, i_7205, i_8466, i_9366);
  not ginst3324 (i_9608, i_9001);
  and ginst3325 (i_9611, i_8485, i_9001);
  and ginst3326 (i_9612, i_7318, i_8519, i_9392);
  and ginst3327 (i_9613, i_7314, i_8522, i_9393);
  and ginst3328 (i_9614, i_6131, i_7325, i_9394);
  and ginst3329 (i_9615, i_6127, i_7328, i_9395);
  not ginst3330 (i_9616, i_9029);
  not ginst3331 (i_9617, i_9035);
  and ginst3332 (i_9618, i_8541, i_9035);
  and ginst3333 (i_9621, i_7384, i_7387, i_9413);
  and ginst3334 (i_9622, i_6177, i_8555, i_9414);
  and ginst3335 (i_9623, i_7398, i_8558, i_9415);
  and ginst3336 (i_9624, i_7394, i_8561, i_9416);
  or ginst3337 (i_9626, i_4563, i_8352, i_8353, i_8354, i_9285);
  or ginst3338 (i_9629, i_4566, i_8355, i_8356, i_9286);
  or ginst3339 (i_9632, i_4570, i_8357, i_9287);
  or ginst3340 (i_9635, i_5960, i_9288);
  nand ginst3341 (i_9642, i_9067, i_9432);
  not ginst3342 (i_9645, i_9068);
  nand ginst3343 (i_9646, i_9073, i_9435);
  not ginst3344 (i_9649, i_9074);
  nand ginst3345 (i_9650, i_9256, i_9257);
  nand ginst3346 (i_9653, i_9258, i_9259);
  nand ginst3347 (i_9656, i_9260, i_9261);
  not ginst3348 (i_9659, i_9079);
  nand ginst3349 (i_9660, i_4809, i_9079);
  not ginst3350 (i_9661, i_9083);
  nand ginst3351 (i_9662, i_6202, i_9083);
  nand ginst3352 (i_9663, i_9088, i_9442);
  not ginst3353 (i_9666, i_9089);
  nand ginst3354 (i_9667, i_9094, i_9445);
  not ginst3355 (i_9670, i_9095);
  or ginst3356 (i_9671, i_8393, i_8924);
  not ginst3357 (i_9674, i_9117);
  not ginst3358 (i_9675, i_8924);
  not ginst3359 (i_9678, i_9127);
  or ginst3360 (i_9679, i_4597, i_8388, i_8389, i_9315);
  or ginst3361 (i_9682, i_8931, i_9318);
  or ginst3362 (i_9685, i_4593, i_8382, i_8383, i_8384, i_9314);
  not ginst3363 (i_9690, i_9146);
  nand ginst3364 (i_9691, i_8717, i_9146);
  not ginst3365 (i_9692, i_8931);
  not ginst3366 (i_9695, i_9149);
  nand ginst3367 (i_9698, i_9400, i_9401);
  nand ginst3368 (i_9702, i_9367, i_9368);
  or ginst3369 (i_9707, i_8517, i_8996);
  not ginst3370 (i_9710, i_9183);
  not ginst3371 (i_9711, i_8996);
  not ginst3372 (i_9714, i_9193);
  not ginst3373 (i_9715, i_9203);
  nand ginst3374 (i_9716, i_6235, i_9203);
  or ginst3375 (i_9717, i_8518, i_9005);
  not ginst3376 (i_9720, i_9206);
  not ginst3377 (i_9721, i_9220);
  nand ginst3378 (i_9722, i_7573, i_9220);
  not ginst3379 (i_9723, i_9005);
  not ginst3380 (i_9726, i_9223);
  nand ginst3381 (i_9727, i_9417, i_9418);
  and ginst3382 (i_9732, i_8269, i_9268);
  nand ginst3383 (i_9733, i_9326, i_9581);
  and ginst3384 (i_9734, i_89, i_8394, i_8421, i_9332, i_9408);
  and ginst3385 (i_9735, i_89, i_8394, i_8421, i_9332, i_9408);
  and ginst3386 (i_9736, i_8262, i_9265);
  not ginst3387 (i_9737, i_9555);
  not ginst3388 (i_9738, i_9556);
  nand ginst3389 (i_9739, i_9361, i_9601);
  nand ginst3390 (i_9740, i_1115, i_9423);
  not ginst3391 (i_9741, i_9423);
  nand ginst3392 (i_9742, i_9299, i_9570);
  and ginst3393 (i_9754, i_8333, i_9280);
  or ginst3394 (i_9758, i_8898, i_9560);
  nand ginst3395 (i_9762, i_8660, i_9561);
  nand ginst3396 (i_9763, i_8663, i_9563);
  nand ginst3397 (i_9764, i_8666, i_9565);
  nand ginst3398 (i_9765, i_8669, i_9567);
  nand ginst3399 (i_9766, i_9297, i_9569);
  and ginst3400 (i_9767, i_367, i_9280);
  nand ginst3401 (i_9768, i_9276, i_9557);
  not ginst3402 (i_9769, i_9307);
  nand ginst3403 (i_9773, i_367, i_9307);
  nand ginst3404 (i_9774, i_9301, i_9571);
  and ginst3405 (i_9775, i_8365, i_9307);
  or ginst3406 (i_9779, i_8920, i_9579);
  not ginst3407 (i_9784, i_9478);
  nand ginst3408 (i_9785, i_9402, i_9616);
  or ginst3409 (i_9786, i_8950, i_9585);
  and ginst3410 (i_9790, i_89, i_8394, i_9332, i_9408);
  or ginst3411 (i_9791, i_8963, i_9591);
  nand ginst3412 (i_9795, i_8735, i_9592);
  nand ginst3413 (i_9796, i_8738, i_9594);
  nand ginst3414 (i_9797, i_8741, i_9596);
  nand ginst3415 (i_9798, i_8744, i_9598);
  nand ginst3416 (i_9799, i_9359, i_9600);
  nor ginst3417 (i_9800, i_9369, i_9602);
  nor ginst3418 (i_9801, i_9370, i_9603);
  nor ginst3419 (i_9802, i_9371, i_9604);
  nor ginst3420 (i_9803, i_9372, i_9605);
  not ginst3421 (i_9805, i_9485);
  not ginst3422 (i_9806, i_9488);
  or ginst3423 (i_9809, i_8995, i_9611);
  nor ginst3424 (i_9813, i_9396, i_9612);
  nor ginst3425 (i_9814, i_9397, i_9613);
  nor ginst3426 (i_9815, i_9398, i_9614);
  nor ginst3427 (i_9816, i_9399, i_9615);
  and ginst3428 (i_9817, i_9407, i_9617);
  or ginst3429 (i_9820, i_9029, i_9618);
  not ginst3430 (i_9825, i_9517);
  not ginst3431 (i_9826, i_9520);
  nor ginst3432 (i_9827, i_9419, i_9621);
  nor ginst3433 (i_9828, i_9420, i_9622);
  nor ginst3434 (i_9829, i_9421, i_9623);
  nor ginst3435 (i_9830, i_9422, i_9624);
  not ginst3436 (i_9835, i_9426);
  nand ginst3437 (i_9836, i_4789, i_9426);
  not ginst3438 (i_9837, i_9429);
  nand ginst3439 (i_9838, i_4794, i_9429);
  nand ginst3440 (i_9846, i_3625, i_9659);
  nand ginst3441 (i_9847, i_4810, i_9661);
  not ginst3442 (i_9862, i_9462);
  nand ginst3443 (i_9863, i_7553, i_9690);
  not ginst3444 (i_9866, i_9473);
  nand ginst3445 (i_9873, i_5030, i_9715);
  nand ginst3446 (i_9876, i_6236, i_9721);
  nand ginst3447 (i_9890, i_9593, i_9795);
  nand ginst3448 (i_9891, i_9597, i_9797);
  not ginst3449 (i_9892, i_9799);
  nand ginst3450 (i_9893, i_871, i_9741);
  nand ginst3451 (i_9894, i_9562, i_9762);
  nand ginst3452 (i_9895, i_9566, i_9764);
  not ginst3453 (i_9896, i_9766);
  not ginst3454 (i_9897, i_9626);
  nand ginst3455 (i_9898, i_9249, i_9626);
  not ginst3456 (i_9899, i_9629);
  nand ginst3457 (i_9900, i_9250, i_9629);
  not ginst3458 (i_9901, i_9632);
  nand ginst3459 (i_9902, i_9251, i_9632);
  not ginst3460 (i_9903, i_9635);
  nand ginst3461 (i_9904, i_9252, i_9635);
  not ginst3462 (i_9905, i_9543);
  not ginst3463 (i_9906, i_9650);
  nand ginst3464 (i_9907, i_5769, i_9650);
  not ginst3465 (i_9908, i_9653);
  nand ginst3466 (i_9909, i_5770, i_9653);
  not ginst3467 (i_9910, i_9656);
  nand ginst3468 (i_9911, i_9262, i_9656);
  not ginst3469 (i_9917, i_9551);
  nand ginst3470 (i_9923, i_9564, i_9763);
  nand ginst3471 (i_9924, i_9568, i_9765);
  or ginst3472 (i_9925, i_8902, i_9767);
  and ginst3473 (i_9932, i_9575, i_9773);
  and ginst3474 (i_9935, i_9575, i_9769);
  not ginst3475 (i_9938, i_9698);
  nand ginst3476 (i_9939, i_9323, i_9698);
  nand ginst3477 (i_9945, i_9595, i_9796);
  nand ginst3478 (i_9946, i_9599, i_9798);
  not ginst3479 (i_9947, i_9702);
  nand ginst3480 (i_9948, i_6102, i_9702);
  and ginst3481 (i_9949, i_9375, i_9608);
  not ginst3482 (i_9953, i_9727);
  nand ginst3483 (i_9954, i_9412, i_9727);
  nand ginst3484 (i_9955, i_3502, i_9835);
  nand ginst3485 (i_9956, i_3510, i_9837);
  not ginst3486 (i_9957, i_9642);
  nand ginst3487 (i_9958, i_9642, i_9645);
  not ginst3488 (i_9959, i_9646);
  nand ginst3489 (i_9960, i_9646, i_9649);
  nand ginst3490 (i_9961, i_9660, i_9846);
  nand ginst3491 (i_9964, i_9662, i_9847);
  not ginst3492 (i_9967, i_9663);
  nand ginst3493 (i_9968, i_9663, i_9666);
  not ginst3494 (i_9969, i_9667);
  nand ginst3495 (i_9970, i_9667, i_9670);
  not ginst3496 (i_9971, i_9671);
  nand ginst3497 (i_9972, i_6213, i_9671);
  not ginst3498 (i_9973, i_9675);
  nand ginst3499 (i_9974, i_7551, i_9675);
  not ginst3500 (i_9975, i_9679);
  nand ginst3501 (i_9976, i_7552, i_9679);
  not ginst3502 (i_9977, i_9682);
  not ginst3503 (i_9978, i_9685);
  nand ginst3504 (i_9979, i_9691, i_9863);
  not ginst3505 (i_9982, i_9692);
  nand ginst3506 (i_9983, i_9813, i_9814);
  nand ginst3507 (i_9986, i_9815, i_9816);
  nand ginst3508 (i_9989, i_9800, i_9801);
  nand ginst3509 (i_9992, i_9802, i_9803);
  not ginst3510 (i_9995, i_9707);
  nand ginst3511 (i_9996, i_6231, i_9707);
  not ginst3512 (i_9997, i_9711);
  nand ginst3513 (i_9998, i_7572, i_9711);
  nand ginst3514 (i_9999, i_9716, i_9873);

SatHard block1 (flip_signal, i_2344, i_6547, i_3343, i_4570, keyinput0, keyinput1, keyinput2, keyinput3, keyinput4, keyinput5, keyinput6, keyinput7);

endmodule
/*************** SatHard block ***************/
module SatHard (flip_signal, i_2344, i_6547, i_3343, i_4570, keyinput0, keyinput1, keyinput2, keyinput3, keyinput4, keyinput5, keyinput6, keyinput7);

  input i_2344, i_6547, i_3343, i_4570, keyinput0, keyinput1, keyinput2, keyinput3, keyinput4, keyinput5, keyinput6, keyinput7;
  output flip_signal;
  //SatHard key=01000001
  wire [3:0] sat_res_inputs;
  assign sat_res_inputs[3:0] = {i_2344, i_6547, i_3343, i_4570};
  wire [7:0] keyinputs, keyvalue;
  assign keyinputs[7:0] = {keyinput0, keyinput1, keyinput2, keyinput3, keyinput4, keyinput5, keyinput6, keyinput7};
  assign keyvalue[7:0] = 8'b01000001;

  wire g, g_bar;
  assign g = &(keyinputs[3:0] ^ sat_res_inputs ^ keyvalue[3:0]);
  assign g_bar = ~&(keyinputs[7:4] ^ sat_res_inputs ^ keyvalue[7:4]);
  assign flip_signal = g & g_bar;

endmodule
/*************** SatHard block ***************/
