//key=10011010110001101101000011100100
// Main module
module b20_C_SFLL-HD(0)_32_0(P2_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, SI_28_, SI_27_, SI_26_, SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, SI_19_, SI_18_, SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, SI_10_, SI_9_, SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, SI_0_, P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN, P2_REG3_REG_7__SCAN_IN, P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_14__SCAN_IN, P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_10__SCAN_IN, P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_19__SCAN_IN, P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_8__SCAN_IN, P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_21__SCAN_IN, P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_25__SCAN_IN, P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_5__SCAN_IN, P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_24__SCAN_IN, P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_9__SCAN_IN, P2_REG3_REG_0__SCAN_IN, P2_REG3_REG_20__SCAN_IN, P2_REG3_REG_13__SCAN_IN, P2_REG3_REG_22__SCAN_IN, P2_REG3_REG_11__SCAN_IN, P2_REG3_REG_2__SCAN_IN, P2_REG3_REG_18__SCAN_IN, P2_REG3_REG_6__SCAN_IN, P2_REG3_REG_26__SCAN_IN, P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN, P2_DATAO_REG_31__SCAN_IN, P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_29__SCAN_IN, P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_27__SCAN_IN, P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_25__SCAN_IN, P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_23__SCAN_IN, P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_21__SCAN_IN, P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_19__SCAN_IN, P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_17__SCAN_IN, P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_15__SCAN_IN, P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_13__SCAN_IN, P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_11__SCAN_IN, P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_9__SCAN_IN, P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_7__SCAN_IN, P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN, P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN, P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN, P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN, P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN, P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN, P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN, P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN, P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN, P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN, P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN, P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN, P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN, P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN, P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN, P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN, P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN, P1_REG1_REG_3__SCAN_IN, P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN, P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN, P1_REG1_REG_9__SCAN_IN, P1_REG1_REG_10__SCAN_IN, P1_REG1_REG_11__SCAN_IN, P1_REG1_REG_12__SCAN_IN, P1_REG1_REG_13__SCAN_IN, P1_REG1_REG_14__SCAN_IN, P1_REG1_REG_15__SCAN_IN, P1_REG1_REG_16__SCAN_IN, P1_REG1_REG_17__SCAN_IN, P1_REG1_REG_18__SCAN_IN, P1_REG1_REG_19__SCAN_IN, P1_REG1_REG_20__SCAN_IN, P1_REG1_REG_21__SCAN_IN, P1_REG1_REG_22__SCAN_IN, P1_REG1_REG_23__SCAN_IN, P1_REG1_REG_24__SCAN_IN, P1_REG1_REG_25__SCAN_IN, P1_REG1_REG_26__SCAN_IN, P1_REG1_REG_27__SCAN_IN, P1_REG1_REG_28__SCAN_IN, P1_REG1_REG_29__SCAN_IN, P1_REG1_REG_30__SCAN_IN, P1_REG1_REG_31__SCAN_IN, P1_REG2_REG_0__SCAN_IN, P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN, P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN, P1_REG2_REG_6__SCAN_IN, P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN, P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN, P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN, P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN, P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN, P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN, P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN, P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN, P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN, P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN, P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN, P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN, P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN, P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN, P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN, P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN, P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN, P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN, P1_ADDR_REG_6__SCAN_IN, P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN, P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN, P1_ADDR_REG_0__SCAN_IN, P1_DATAO_REG_0__SCAN_IN, P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, P1_REG3_REG_15__SCAN_IN, P1_REG3_REG_26__SCAN_IN, P1_REG3_REG_6__SCAN_IN, P1_REG3_REG_18__SCAN_IN, P1_REG3_REG_2__SCAN_IN, P1_REG3_REG_11__SCAN_IN, P1_REG3_REG_22__SCAN_IN, P1_REG3_REG_13__SCAN_IN, P1_REG3_REG_20__SCAN_IN, P1_REG3_REG_0__SCAN_IN, P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN, P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN, P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN, P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN, P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN, P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN, P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN, P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN, P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN, P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN, P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN, P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN, P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN, P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN, P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN, P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN, P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN, P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN, P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN, P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN, P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN, P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN, P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN, P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN, P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN, P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN, P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN, P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN, P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN, P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN, P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN, P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN, P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN, P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN, P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN, P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN, P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN, P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN, P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN, P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN, P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN, P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN, P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN, P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN, P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN, P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN, P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN, P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN, P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN, P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN, P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN, P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN, P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN, P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN, P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN, P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN, P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN, P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN, P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN, P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN, P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN, P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN, P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN, P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN, P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN, P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN, P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN, P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN, P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN, P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN, P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN, P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN, P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN, P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN, P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN, P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN, P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN, P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN, P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN, P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN, P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN, P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN, P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN, P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN, P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN, P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN, P2_DATAO_REG_5__SCAN_IN, P2_DATAO_REG_6__SCAN_IN, keyinput0, keyinput1, keyinput2, keyinput3, keyinput4, keyinput5, keyinput6, keyinput7, keyinput8, keyinput9, keyinput10, keyinput11, keyinput12, keyinput13, keyinput14, keyinput15, keyinput16, keyinput17, keyinput18, keyinput19, keyinput20, keyinput21, keyinput22, keyinput23, keyinput24, keyinput25, keyinput26, keyinput27, keyinput28, keyinput29, keyinput30, keyinput31, ADD_1068_U4, ADD_1068_U55, ADD_1068_U56, ADD_1068_U57, ADD_1068_U58, ADD_1068_U59, ADD_1068_U60, ADD_1068_U61, ADD_1068_U62, ADD_1068_U63, ADD_1068_U47, ADD_1068_U48, ADD_1068_U49, ADD_1068_U50, ADD_1068_U51, ADD_1068_U52, ADD_1068_U53, ADD_1068_U54, ADD_1068_U5, ADD_1068_U46, U126, U123, P1_U3355, P1_U3354, P1_U3353, P1_U3352, P1_U3351, P1_U3350, P1_U3349, P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, P1_U3343, P1_U3342, P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, P1_U3336, P1_U3335, P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, P1_U3329, P1_U3328, P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3439, P1_U3440, P1_U3323, P1_U3322, P1_U3321, P1_U3320, P1_U3319, P1_U3318, P1_U3317, P1_U3316, P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, P1_U3310, P1_U3309, P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, P1_U3303, P1_U3302, P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, P1_U3296, P1_U3295, P1_U3294, P1_U3453, P1_U3456, P1_U3459, P1_U3462, P1_U3465, P1_U3468, P1_U3471, P1_U3474, P1_U3477, P1_U3480, P1_U3483, P1_U3486, P1_U3489, P1_U3492, P1_U3495, P1_U3498, P1_U3501, P1_U3504, P1_U3507, P1_U3509, P1_U3510, P1_U3511, P1_U3512, P1_U3513, P1_U3514, P1_U3515, P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521, P1_U3522, P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528, P1_U3529, P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535, P1_U3536, P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542, P1_U3543, P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549, P1_U3550, P1_U3551, P1_U3552, P1_U3553, P1_U3293, P1_U3292, P1_U3291, P1_U3290, P1_U3289, P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, P1_U3283, P1_U3282, P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, P1_U3276, P1_U3275, P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, P1_U3269, P1_U3268, P1_U3267, P1_U3266, P1_U3265, P1_U3356, P1_U3264, P1_U3263, P1_U3262, P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, P1_U3256, P1_U3255, P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, P1_U3249, P1_U3248, P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, P1_U3554, P1_U3555, P1_U3556, P1_U3557, P1_U3558, P1_U3559, P1_U3560, P1_U3561, P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567, P1_U3568, P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574, P1_U3575, P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581, P1_U3582, P1_U3583, P1_U3584, P1_U3585, P1_U3242, P1_U3241, P1_U3240, P1_U3239, P1_U3238, P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, P1_U3232, P1_U3231, P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, P1_U3225, P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218, P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3086, P1_U3085, P1_U3973, P2_U3295, P2_U3294, P2_U3293, P2_U3292, P2_U3291, P2_U3290, P2_U3289, P2_U3288, P2_U3287, P2_U3286, P2_U3285, P2_U3284, P2_U3283, P2_U3282, P2_U3281, P2_U3280, P2_U3279, P2_U3278, P2_U3277, P2_U3276, P2_U3275, P2_U3274, P2_U3273, P2_U3272, P2_U3271, P2_U3270, P2_U3269, P2_U3268, P2_U3267, P2_U3266, P2_U3265, P2_U3264, P2_U3376, P2_U3377, P2_U3263, P2_U3262, P2_U3261, P2_U3260, P2_U3259, P2_U3258, P2_U3257, P2_U3256, P2_U3255, P2_U3254, P2_U3253, P2_U3252, P2_U3251, P2_U3250, P2_U3249, P2_U3248, P2_U3247, P2_U3246, P2_U3245, P2_U3244, P2_U3243, P2_U3242, P2_U3241, P2_U3240, P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234, P2_U3390, P2_U3393, P2_U3396, P2_U3399, P2_U3402, P2_U3405, P2_U3408, P2_U3411, P2_U3414, P2_U3417, P2_U3420, P2_U3423, P2_U3426, P2_U3429, P2_U3432, P2_U3435, P2_U3438, P2_U3441, P2_U3444, P2_U3446, P2_U3447, P2_U3448, P2_U3449, P2_U3450, P2_U3451, P2_U3452, P2_U3453, P2_U3454, P2_U3455, P2_U3456, P2_U3457, P2_U3458, P2_U3459, P2_U3460, P2_U3461, P2_U3462, P2_U3463, P2_U3464, P2_U3465, P2_U3466, P2_U3467, P2_U3468, P2_U3469, P2_U3470, P2_U3471, P2_U3472, P2_U3473, P2_U3474, P2_U3475, P2_U3476, P2_U3477, P2_U3478, P2_U3479, P2_U3480, P2_U3481, P2_U3482, P2_U3483, P2_U3484, P2_U3485, P2_U3486, P2_U3487, P2_U3488, P2_U3489, P2_U3490, P2_U3233, P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227, P2_U3226, P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220, P2_U3219, P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3214, P2_U3213, P2_U3212, P2_U3211, P2_U3210, P2_U3209, P2_U3208, P2_U3207, P2_U3206, P2_U3205, P2_U3204, P2_U3203, P2_U3202, P2_U3201, P2_U3200, P2_U3199, P2_U3198, P2_U3197, P2_U3196, P2_U3195, P2_U3194, P2_U3193, P2_U3192, P2_U3191, P2_U3190, P2_U3189, P2_U3188, P2_U3187, P2_U3186, P2_U3185, P2_U3184, P2_U3183, P2_U3182, P2_U3491, P2_U3492, P2_U3493, P2_U3494, P2_U3495, P2_U3496, P2_U3497, P2_U3498, P2_U3499, P2_U3500, P2_U3501, P2_U3502, P2_U3503, P2_U3504, P2_U3505, P2_U3506, P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511, P2_U3512, P2_U3513, P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518, P2_U3519, P2_U3520, P2_U3521, P2_U3522, P2_U3296, P2_U3181, P2_U3180, P2_U3179, P2_U3178, P2_U3177, P2_U3176, P2_U3175, P2_U3174, P2_U3173, P2_U3172, P2_U3171, P2_U3170, P2_U3169, P2_U3168, P2_U3167, P2_U3166, P2_U3165, P2_U3164, P2_U3163, P2_U3162, P2_U3161, P2_U3160, P2_U3159, P2_U3158, P2_U3157, P2_U3156, P2_U3155, P2_U3154, P2_U3153, P2_U3151, P2_U3150, P2_U3893);

  input P2_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, SI_28_, SI_27_, SI_26_, SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, SI_19_, SI_18_, SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, SI_10_, SI_9_, SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, SI_0_, P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN, P2_REG3_REG_7__SCAN_IN, P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_14__SCAN_IN, P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_10__SCAN_IN, P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_19__SCAN_IN, P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_8__SCAN_IN, P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_21__SCAN_IN, P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_25__SCAN_IN, P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_5__SCAN_IN, P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_24__SCAN_IN, P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_9__SCAN_IN, P2_REG3_REG_0__SCAN_IN, P2_REG3_REG_20__SCAN_IN, P2_REG3_REG_13__SCAN_IN, P2_REG3_REG_22__SCAN_IN, P2_REG3_REG_11__SCAN_IN, P2_REG3_REG_2__SCAN_IN, P2_REG3_REG_18__SCAN_IN, P2_REG3_REG_6__SCAN_IN, P2_REG3_REG_26__SCAN_IN, P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN, P2_DATAO_REG_31__SCAN_IN, P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_29__SCAN_IN, P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_27__SCAN_IN, P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_25__SCAN_IN, P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_23__SCAN_IN, P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_21__SCAN_IN, P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_19__SCAN_IN, P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_17__SCAN_IN, P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_15__SCAN_IN, P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_13__SCAN_IN, P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_11__SCAN_IN, P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_9__SCAN_IN, P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_7__SCAN_IN, P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN, P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN, P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN, P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN, P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN, P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN, P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN, P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN, P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN, P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN, P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN, P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN, P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN, P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN, P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN, P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN, P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN, P1_REG1_REG_3__SCAN_IN, P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN, P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN, P1_REG1_REG_9__SCAN_IN, P1_REG1_REG_10__SCAN_IN, P1_REG1_REG_11__SCAN_IN, P1_REG1_REG_12__SCAN_IN, P1_REG1_REG_13__SCAN_IN, P1_REG1_REG_14__SCAN_IN, P1_REG1_REG_15__SCAN_IN, P1_REG1_REG_16__SCAN_IN, P1_REG1_REG_17__SCAN_IN, P1_REG1_REG_18__SCAN_IN, P1_REG1_REG_19__SCAN_IN, P1_REG1_REG_20__SCAN_IN, P1_REG1_REG_21__SCAN_IN, P1_REG1_REG_22__SCAN_IN, P1_REG1_REG_23__SCAN_IN, P1_REG1_REG_24__SCAN_IN, P1_REG1_REG_25__SCAN_IN, P1_REG1_REG_26__SCAN_IN, P1_REG1_REG_27__SCAN_IN, P1_REG1_REG_28__SCAN_IN, P1_REG1_REG_29__SCAN_IN, P1_REG1_REG_30__SCAN_IN, P1_REG1_REG_31__SCAN_IN, P1_REG2_REG_0__SCAN_IN, P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN, P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN, P1_REG2_REG_6__SCAN_IN, P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN, P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN, P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN, P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN, P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN, P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN, P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN, P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN, P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN, P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN, P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN, P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN, P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN, P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN, P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN, P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN, P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN, P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN, P1_ADDR_REG_6__SCAN_IN, P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN, P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN, P1_ADDR_REG_0__SCAN_IN, P1_DATAO_REG_0__SCAN_IN, P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, P1_REG3_REG_15__SCAN_IN, P1_REG3_REG_26__SCAN_IN, P1_REG3_REG_6__SCAN_IN, P1_REG3_REG_18__SCAN_IN, P1_REG3_REG_2__SCAN_IN, P1_REG3_REG_11__SCAN_IN, P1_REG3_REG_22__SCAN_IN, P1_REG3_REG_13__SCAN_IN, P1_REG3_REG_20__SCAN_IN, P1_REG3_REG_0__SCAN_IN, P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN, P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN, P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN, P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN, P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN, P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN, P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN, P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN, P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN, P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN, P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN, P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN, P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN, P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN, P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN, P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN, P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN, P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN, P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN, P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN, P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN, P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN, P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN, P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN, P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN, P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN, P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN, P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN, P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN, P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN, P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN, P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN, P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN, P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN, P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN, P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN, P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN, P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN, P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN, P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN, P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN, P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN, P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN, P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN, P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN, P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN, P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN, P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN, P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN, P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN, P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN, P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN, P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN, P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN, P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN, P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN, P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN, P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN, P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN, P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN, P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN, P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN, P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN, P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN, P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN, P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN, P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN, P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN, P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN, P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN, P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN, P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN, P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN, P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN, P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN, P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN, P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN, P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN, P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN, P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN, P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN, P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN, P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN, P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN, P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN, P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN, P2_DATAO_REG_5__SCAN_IN, P2_DATAO_REG_6__SCAN_IN, keyinput0, keyinput1, keyinput2, keyinput3, keyinput4, keyinput5, keyinput6, keyinput7, keyinput8, keyinput9, keyinput10, keyinput11, keyinput12, keyinput13, keyinput14, keyinput15, keyinput16, keyinput17, keyinput18, keyinput19, keyinput20, keyinput21, keyinput22, keyinput23, keyinput24, keyinput25, keyinput26, keyinput27, keyinput28, keyinput29, keyinput30, keyinput31;
  output ADD_1068_U4, ADD_1068_U55, ADD_1068_U56, ADD_1068_U57, ADD_1068_U58, ADD_1068_U59, ADD_1068_U60, ADD_1068_U61, ADD_1068_U62, ADD_1068_U63, ADD_1068_U47, ADD_1068_U48, ADD_1068_U49, ADD_1068_U50, ADD_1068_U51, ADD_1068_U52, ADD_1068_U53, ADD_1068_U54, ADD_1068_U5, ADD_1068_U46, U126, U123, P1_U3355, P1_U3354, P1_U3353, P1_U3352, P1_U3351, P1_U3350, P1_U3349, P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, P1_U3343, P1_U3342, P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, P1_U3336, P1_U3335, P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, P1_U3329, P1_U3328, P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3439, P1_U3440, P1_U3323, P1_U3322, P1_U3321, P1_U3320, P1_U3319, P1_U3318, P1_U3317, P1_U3316, P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, P1_U3310, P1_U3309, P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, P1_U3303, P1_U3302, P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, P1_U3296, P1_U3295, P1_U3294, P1_U3453, P1_U3456, P1_U3459, P1_U3462, P1_U3465, P1_U3468, P1_U3471, P1_U3474, P1_U3477, P1_U3480, P1_U3483, P1_U3486, P1_U3489, P1_U3492, P1_U3495, P1_U3498, P1_U3501, P1_U3504, P1_U3507, P1_U3509, P1_U3510, P1_U3511, P1_U3512, P1_U3513, P1_U3514, P1_U3515, P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521, P1_U3522, P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528, P1_U3529, P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535, P1_U3536, P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542, P1_U3543, P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549, P1_U3550, P1_U3551, P1_U3552, P1_U3553, P1_U3293, P1_U3292, P1_U3291, P1_U3290, P1_U3289, P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, P1_U3283, P1_U3282, P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, P1_U3276, P1_U3275, P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, P1_U3269, P1_U3268, P1_U3267, P1_U3266, P1_U3265, P1_U3356, P1_U3264, P1_U3263, P1_U3262, P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, P1_U3256, P1_U3255, P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, P1_U3249, P1_U3248, P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, P1_U3554, P1_U3555, P1_U3556, P1_U3557, P1_U3558, P1_U3559, P1_U3560, P1_U3561, P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567, P1_U3568, P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574, P1_U3575, P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581, P1_U3582, P1_U3583, P1_U3584, P1_U3585, P1_U3242, P1_U3241, P1_U3240, P1_U3239, P1_U3238, P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, P1_U3232, P1_U3231, P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, P1_U3225, P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218, P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3086, P1_U3085, P1_U3973, P2_U3295, P2_U3294, P2_U3293, P2_U3292, P2_U3291, P2_U3290, P2_U3289, P2_U3288, P2_U3287, P2_U3286, P2_U3285, P2_U3284, P2_U3283, P2_U3282, P2_U3281, P2_U3280, P2_U3279, P2_U3278, P2_U3277, P2_U3276, P2_U3275, P2_U3274, P2_U3273, P2_U3272, P2_U3271, P2_U3270, P2_U3269, P2_U3268, P2_U3267, P2_U3266, P2_U3265, P2_U3264, P2_U3376, P2_U3377, P2_U3263, P2_U3262, P2_U3261, P2_U3260, P2_U3259, P2_U3258, P2_U3257, P2_U3256, P2_U3255, P2_U3254, P2_U3253, P2_U3252, P2_U3251, P2_U3250, P2_U3249, P2_U3248, P2_U3247, P2_U3246, P2_U3245, P2_U3244, P2_U3243, P2_U3242, P2_U3241, P2_U3240, P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234, P2_U3390, P2_U3393, P2_U3396, P2_U3399, P2_U3402, P2_U3405, P2_U3408, P2_U3411, P2_U3414, P2_U3417, P2_U3420, P2_U3423, P2_U3426, P2_U3429, P2_U3432, P2_U3435, P2_U3438, P2_U3441, P2_U3444, P2_U3446, P2_U3447, P2_U3448, P2_U3449, P2_U3450, P2_U3451, P2_U3452, P2_U3453, P2_U3454, P2_U3455, P2_U3456, P2_U3457, P2_U3458, P2_U3459, P2_U3460, P2_U3461, P2_U3462, P2_U3463, P2_U3464, P2_U3465, P2_U3466, P2_U3467, P2_U3468, P2_U3469, P2_U3470, P2_U3471, P2_U3472, P2_U3473, P2_U3474, P2_U3475, P2_U3476, P2_U3477, P2_U3478, P2_U3479, P2_U3480, P2_U3481, P2_U3482, P2_U3483, P2_U3484, P2_U3485, P2_U3486, P2_U3487, P2_U3488, P2_U3489, P2_U3490, P2_U3233, P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227, P2_U3226, P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220, P2_U3219, P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3214, P2_U3213, P2_U3212, P2_U3211, P2_U3210, P2_U3209, P2_U3208, P2_U3207, P2_U3206, P2_U3205, P2_U3204, P2_U3203, P2_U3202, P2_U3201, P2_U3200, P2_U3199, P2_U3198, P2_U3197, P2_U3196, P2_U3195, P2_U3194, P2_U3193, P2_U3192, P2_U3191, P2_U3190, P2_U3189, P2_U3188, P2_U3187, P2_U3186, P2_U3185, P2_U3184, P2_U3183, P2_U3182, P2_U3491, P2_U3492, P2_U3493, P2_U3494, P2_U3495, P2_U3496, P2_U3497, P2_U3498, P2_U3499, P2_U3500, P2_U3501, P2_U3502, P2_U3503, P2_U3504, P2_U3505, P2_U3506, P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511, P2_U3512, P2_U3513, P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518, P2_U3519, P2_U3520, P2_U3521, P2_U3522, P2_U3296, P2_U3181, P2_U3180, P2_U3179, P2_U3178, P2_U3177, P2_U3176, P2_U3175, P2_U3174, P2_U3173, P2_U3172, P2_U3171, P2_U3170, P2_U3169, P2_U3168, P2_U3167, P2_U3166, P2_U3165, P2_U3164, P2_U3163, P2_U3162, P2_U3161, P2_U3160, P2_U3159, P2_U3158, P2_U3157, P2_U3156, P2_U3155, P2_U3154, P2_U3153, P2_U3151, P2_U3150, P2_U3893;
  wire ADD_1068_U10, ADD_1068_U100, ADD_1068_U101, ADD_1068_U102, ADD_1068_U103, ADD_1068_U104, ADD_1068_U105, ADD_1068_U106, ADD_1068_U107, ADD_1068_U108, ADD_1068_U109, ADD_1068_U11, ADD_1068_U110, ADD_1068_U111, ADD_1068_U112, ADD_1068_U113, ADD_1068_U114, ADD_1068_U115, ADD_1068_U116, ADD_1068_U117, ADD_1068_U118, ADD_1068_U119, ADD_1068_U12, ADD_1068_U120, ADD_1068_U121, ADD_1068_U122, ADD_1068_U123, ADD_1068_U124, ADD_1068_U125, ADD_1068_U126, ADD_1068_U127, ADD_1068_U128, ADD_1068_U129, ADD_1068_U13, ADD_1068_U130, ADD_1068_U131, ADD_1068_U132, ADD_1068_U133, ADD_1068_U134, ADD_1068_U135, ADD_1068_U136, ADD_1068_U137, ADD_1068_U138, ADD_1068_U139, ADD_1068_U14, ADD_1068_U140, ADD_1068_U141, ADD_1068_U142, ADD_1068_U143, ADD_1068_U144, ADD_1068_U145, ADD_1068_U146, ADD_1068_U147, ADD_1068_U148, ADD_1068_U149, ADD_1068_U15, ADD_1068_U150, ADD_1068_U151, ADD_1068_U152, ADD_1068_U153, ADD_1068_U154, ADD_1068_U155, ADD_1068_U156, ADD_1068_U157, ADD_1068_U158, ADD_1068_U159, ADD_1068_U16, ADD_1068_U160, ADD_1068_U161, ADD_1068_U162, ADD_1068_U163, ADD_1068_U164, ADD_1068_U165, ADD_1068_U166, ADD_1068_U167, ADD_1068_U168, ADD_1068_U169, ADD_1068_U17, ADD_1068_U170, ADD_1068_U171, ADD_1068_U172, ADD_1068_U173, ADD_1068_U174, ADD_1068_U175, ADD_1068_U176, ADD_1068_U177, ADD_1068_U178, ADD_1068_U179, ADD_1068_U18, ADD_1068_U180, ADD_1068_U181, ADD_1068_U182, ADD_1068_U183, ADD_1068_U184, ADD_1068_U185, ADD_1068_U186, ADD_1068_U187, ADD_1068_U188, ADD_1068_U189, ADD_1068_U19, ADD_1068_U190, ADD_1068_U191, ADD_1068_U192, ADD_1068_U193, ADD_1068_U194, ADD_1068_U195, ADD_1068_U196, ADD_1068_U197, ADD_1068_U198, ADD_1068_U199, ADD_1068_U20, ADD_1068_U200, ADD_1068_U201, ADD_1068_U202, ADD_1068_U203, ADD_1068_U204, ADD_1068_U205, ADD_1068_U206, ADD_1068_U207, ADD_1068_U208, ADD_1068_U209, ADD_1068_U21, ADD_1068_U210, ADD_1068_U211, ADD_1068_U212, ADD_1068_U213, ADD_1068_U214, ADD_1068_U215, ADD_1068_U216, ADD_1068_U217, ADD_1068_U218, ADD_1068_U219, ADD_1068_U22, ADD_1068_U220, ADD_1068_U221, ADD_1068_U222, ADD_1068_U223, ADD_1068_U224, ADD_1068_U225, ADD_1068_U226, ADD_1068_U227, ADD_1068_U228, ADD_1068_U229, ADD_1068_U23, ADD_1068_U230, ADD_1068_U231, ADD_1068_U232, ADD_1068_U233, ADD_1068_U234, ADD_1068_U235, ADD_1068_U236, ADD_1068_U237, ADD_1068_U238, ADD_1068_U239, ADD_1068_U24, ADD_1068_U240, ADD_1068_U241, ADD_1068_U242, ADD_1068_U243, ADD_1068_U244, ADD_1068_U245, ADD_1068_U246, ADD_1068_U247, ADD_1068_U248, ADD_1068_U249, ADD_1068_U25, ADD_1068_U250, ADD_1068_U251, ADD_1068_U252, ADD_1068_U253, ADD_1068_U254, ADD_1068_U255, ADD_1068_U256, ADD_1068_U257, ADD_1068_U258, ADD_1068_U259, ADD_1068_U26, ADD_1068_U260, ADD_1068_U261, ADD_1068_U262, ADD_1068_U263, ADD_1068_U264, ADD_1068_U265, ADD_1068_U266, ADD_1068_U267, ADD_1068_U268, ADD_1068_U269, ADD_1068_U27, ADD_1068_U270, ADD_1068_U271, ADD_1068_U272, ADD_1068_U273, ADD_1068_U274, ADD_1068_U275, ADD_1068_U276, ADD_1068_U277, ADD_1068_U278, ADD_1068_U279, ADD_1068_U28, ADD_1068_U280, ADD_1068_U281, ADD_1068_U282, ADD_1068_U283, ADD_1068_U284, ADD_1068_U285, ADD_1068_U286, ADD_1068_U287, ADD_1068_U288, ADD_1068_U289, ADD_1068_U29, ADD_1068_U290, ADD_1068_U291, ADD_1068_U30, ADD_1068_U31, ADD_1068_U32, ADD_1068_U33, ADD_1068_U34, ADD_1068_U35, ADD_1068_U36, ADD_1068_U37, ADD_1068_U38, ADD_1068_U39, ADD_1068_U40, ADD_1068_U41, ADD_1068_U42, ADD_1068_U43, ADD_1068_U44, ADD_1068_U45, ADD_1068_U6, ADD_1068_U64, ADD_1068_U65, ADD_1068_U66, ADD_1068_U67, ADD_1068_U68, ADD_1068_U69, ADD_1068_U7, ADD_1068_U70, ADD_1068_U71, ADD_1068_U72, ADD_1068_U73, ADD_1068_U74, ADD_1068_U75, ADD_1068_U76, ADD_1068_U77, ADD_1068_U78, ADD_1068_U79, ADD_1068_U8, ADD_1068_U80, ADD_1068_U81, ADD_1068_U82, ADD_1068_U83, ADD_1068_U84, ADD_1068_U85, ADD_1068_U86, ADD_1068_U87, ADD_1068_U88, ADD_1068_U89, ADD_1068_U9, ADD_1068_U90, ADD_1068_U91, ADD_1068_U92, ADD_1068_U93, ADD_1068_U94, ADD_1068_U95, ADD_1068_U96, ADD_1068_U97, ADD_1068_U98, ADD_1068_U99, LT_1075_19_U6, LT_1075_U6, P1_ADD_95_U10, P1_ADD_95_U100, P1_ADD_95_U101, P1_ADD_95_U102, P1_ADD_95_U103, P1_ADD_95_U104, P1_ADD_95_U105, P1_ADD_95_U106, P1_ADD_95_U107, P1_ADD_95_U108, P1_ADD_95_U109, P1_ADD_95_U11, P1_ADD_95_U110, P1_ADD_95_U111, P1_ADD_95_U112, P1_ADD_95_U113, P1_ADD_95_U114, P1_ADD_95_U115, P1_ADD_95_U116, P1_ADD_95_U117, P1_ADD_95_U118, P1_ADD_95_U119, P1_ADD_95_U12, P1_ADD_95_U120, P1_ADD_95_U121, P1_ADD_95_U122, P1_ADD_95_U123, P1_ADD_95_U124, P1_ADD_95_U125, P1_ADD_95_U126, P1_ADD_95_U127, P1_ADD_95_U128, P1_ADD_95_U129, P1_ADD_95_U13, P1_ADD_95_U130, P1_ADD_95_U131, P1_ADD_95_U132, P1_ADD_95_U133, P1_ADD_95_U134, P1_ADD_95_U135, P1_ADD_95_U136, P1_ADD_95_U137, P1_ADD_95_U138, P1_ADD_95_U139, P1_ADD_95_U14, P1_ADD_95_U140, P1_ADD_95_U141, P1_ADD_95_U142, P1_ADD_95_U143, P1_ADD_95_U144, P1_ADD_95_U145, P1_ADD_95_U146, P1_ADD_95_U147, P1_ADD_95_U148, P1_ADD_95_U149, P1_ADD_95_U15, P1_ADD_95_U150, P1_ADD_95_U151, P1_ADD_95_U152, P1_ADD_95_U153, P1_ADD_95_U16, P1_ADD_95_U17, P1_ADD_95_U18, P1_ADD_95_U19, P1_ADD_95_U20, P1_ADD_95_U21, P1_ADD_95_U22, P1_ADD_95_U23, P1_ADD_95_U24, P1_ADD_95_U25, P1_ADD_95_U26, P1_ADD_95_U27, P1_ADD_95_U28, P1_ADD_95_U29, P1_ADD_95_U30, P1_ADD_95_U31, P1_ADD_95_U32, P1_ADD_95_U33, P1_ADD_95_U34, P1_ADD_95_U35, P1_ADD_95_U36, P1_ADD_95_U37, P1_ADD_95_U38, P1_ADD_95_U39, P1_ADD_95_U4, P1_ADD_95_U40, P1_ADD_95_U41, P1_ADD_95_U42, P1_ADD_95_U43, P1_ADD_95_U44, P1_ADD_95_U45, P1_ADD_95_U46, P1_ADD_95_U47, P1_ADD_95_U48, P1_ADD_95_U49, P1_ADD_95_U5, P1_ADD_95_U50, P1_ADD_95_U51, P1_ADD_95_U52, P1_ADD_95_U53, P1_ADD_95_U54, P1_ADD_95_U55, P1_ADD_95_U56, P1_ADD_95_U57, P1_ADD_95_U58, P1_ADD_95_U59, P1_ADD_95_U6, P1_ADD_95_U60, P1_ADD_95_U61, P1_ADD_95_U62, P1_ADD_95_U63, P1_ADD_95_U64, P1_ADD_95_U65, P1_ADD_95_U66, P1_ADD_95_U67, P1_ADD_95_U68, P1_ADD_95_U69, P1_ADD_95_U7, P1_ADD_95_U70, P1_ADD_95_U71, P1_ADD_95_U72, P1_ADD_95_U73, P1_ADD_95_U74, P1_ADD_95_U75, P1_ADD_95_U76, P1_ADD_95_U77, P1_ADD_95_U78, P1_ADD_95_U79, P1_ADD_95_U8, P1_ADD_95_U80, P1_ADD_95_U81, P1_ADD_95_U82, P1_ADD_95_U83, P1_ADD_95_U84, P1_ADD_95_U85, P1_ADD_95_U86, P1_ADD_95_U87, P1_ADD_95_U88, P1_ADD_95_U89, P1_ADD_95_U9, P1_ADD_95_U90, P1_ADD_95_U91, P1_ADD_95_U92, P1_ADD_95_U93, P1_ADD_95_U94, P1_ADD_95_U95, P1_ADD_95_U96, P1_ADD_95_U97, P1_ADD_95_U98, P1_ADD_95_U99, P1_LT_197_U10, P1_LT_197_U100, P1_LT_197_U101, P1_LT_197_U102, P1_LT_197_U103, P1_LT_197_U104, P1_LT_197_U105, P1_LT_197_U106, P1_LT_197_U107, P1_LT_197_U108, P1_LT_197_U109, P1_LT_197_U11, P1_LT_197_U110, P1_LT_197_U111, P1_LT_197_U112, P1_LT_197_U113, P1_LT_197_U114, P1_LT_197_U115, P1_LT_197_U116, P1_LT_197_U117, P1_LT_197_U118, P1_LT_197_U119, P1_LT_197_U12, P1_LT_197_U120, P1_LT_197_U121, P1_LT_197_U122, P1_LT_197_U123, P1_LT_197_U124, P1_LT_197_U125, P1_LT_197_U126, P1_LT_197_U127, P1_LT_197_U128, P1_LT_197_U129, P1_LT_197_U13, P1_LT_197_U130, P1_LT_197_U131, P1_LT_197_U132, P1_LT_197_U133, P1_LT_197_U134, P1_LT_197_U135, P1_LT_197_U136, P1_LT_197_U137, P1_LT_197_U138, P1_LT_197_U139, P1_LT_197_U14, P1_LT_197_U140, P1_LT_197_U141, P1_LT_197_U142, P1_LT_197_U143, P1_LT_197_U144, P1_LT_197_U145, P1_LT_197_U146, P1_LT_197_U147, P1_LT_197_U148, P1_LT_197_U149, P1_LT_197_U15, P1_LT_197_U150, P1_LT_197_U151, P1_LT_197_U152, P1_LT_197_U153, P1_LT_197_U154, P1_LT_197_U155, P1_LT_197_U156, P1_LT_197_U157, P1_LT_197_U158, P1_LT_197_U159, P1_LT_197_U16, P1_LT_197_U160, P1_LT_197_U161, P1_LT_197_U162, P1_LT_197_U163, P1_LT_197_U164, P1_LT_197_U165, P1_LT_197_U166, P1_LT_197_U167, P1_LT_197_U168, P1_LT_197_U169, P1_LT_197_U17, P1_LT_197_U170, P1_LT_197_U171, P1_LT_197_U172, P1_LT_197_U173, P1_LT_197_U174, P1_LT_197_U175, P1_LT_197_U176, P1_LT_197_U177, P1_LT_197_U178, P1_LT_197_U179, P1_LT_197_U18, P1_LT_197_U180, P1_LT_197_U181, P1_LT_197_U182, P1_LT_197_U183, P1_LT_197_U184, P1_LT_197_U185, P1_LT_197_U186, P1_LT_197_U187, P1_LT_197_U188, P1_LT_197_U189, P1_LT_197_U19, P1_LT_197_U190, P1_LT_197_U191, P1_LT_197_U192, P1_LT_197_U193, P1_LT_197_U194, P1_LT_197_U195, P1_LT_197_U196, P1_LT_197_U197, P1_LT_197_U198, P1_LT_197_U199, P1_LT_197_U20, P1_LT_197_U200, P1_LT_197_U21, P1_LT_197_U22, P1_LT_197_U23, P1_LT_197_U24, P1_LT_197_U25, P1_LT_197_U26, P1_LT_197_U27, P1_LT_197_U28, P1_LT_197_U29, P1_LT_197_U30, P1_LT_197_U31, P1_LT_197_U32, P1_LT_197_U33, P1_LT_197_U34, P1_LT_197_U35, P1_LT_197_U36, P1_LT_197_U37, P1_LT_197_U38, P1_LT_197_U39, P1_LT_197_U40, P1_LT_197_U41, P1_LT_197_U42, P1_LT_197_U43, P1_LT_197_U44, P1_LT_197_U45, P1_LT_197_U46, P1_LT_197_U47, P1_LT_197_U48, P1_LT_197_U49, P1_LT_197_U50, P1_LT_197_U51, P1_LT_197_U52, P1_LT_197_U53, P1_LT_197_U54, P1_LT_197_U55, P1_LT_197_U56, P1_LT_197_U57, P1_LT_197_U58, P1_LT_197_U59, P1_LT_197_U6, P1_LT_197_U60, P1_LT_197_U61, P1_LT_197_U62, P1_LT_197_U63, P1_LT_197_U64, P1_LT_197_U65, P1_LT_197_U66, P1_LT_197_U67, P1_LT_197_U68, P1_LT_197_U69, P1_LT_197_U7, P1_LT_197_U70, P1_LT_197_U71, P1_LT_197_U72, P1_LT_197_U73, P1_LT_197_U74, P1_LT_197_U75, P1_LT_197_U76, P1_LT_197_U77, P1_LT_197_U78, P1_LT_197_U79, P1_LT_197_U8, P1_LT_197_U80, P1_LT_197_U81, P1_LT_197_U82, P1_LT_197_U83, P1_LT_197_U84, P1_LT_197_U85, P1_LT_197_U86, P1_LT_197_U87, P1_LT_197_U88, P1_LT_197_U89, P1_LT_197_U9, P1_LT_197_U90, P1_LT_197_U91, P1_LT_197_U92, P1_LT_197_U93, P1_LT_197_U94, P1_LT_197_U95, P1_LT_197_U96, P1_LT_197_U97, P1_LT_197_U98, P1_LT_197_U99, P1_R1105_U10, P1_R1105_U100, P1_R1105_U101, P1_R1105_U102, P1_R1105_U103, P1_R1105_U104, P1_R1105_U105, P1_R1105_U106, P1_R1105_U107, P1_R1105_U108, P1_R1105_U109, P1_R1105_U11, P1_R1105_U110, P1_R1105_U111, P1_R1105_U112, P1_R1105_U113, P1_R1105_U114, P1_R1105_U115, P1_R1105_U116, P1_R1105_U117, P1_R1105_U118, P1_R1105_U119, P1_R1105_U12, P1_R1105_U120, P1_R1105_U121, P1_R1105_U122, P1_R1105_U123, P1_R1105_U124, P1_R1105_U125, P1_R1105_U126, P1_R1105_U127, P1_R1105_U128, P1_R1105_U129, P1_R1105_U13, P1_R1105_U130, P1_R1105_U131, P1_R1105_U132, P1_R1105_U133, P1_R1105_U134, P1_R1105_U135, P1_R1105_U136, P1_R1105_U137, P1_R1105_U138, P1_R1105_U139, P1_R1105_U14, P1_R1105_U140, P1_R1105_U141, P1_R1105_U142, P1_R1105_U143, P1_R1105_U144, P1_R1105_U145, P1_R1105_U146, P1_R1105_U147, P1_R1105_U148, P1_R1105_U149, P1_R1105_U15, P1_R1105_U150, P1_R1105_U151, P1_R1105_U152, P1_R1105_U153, P1_R1105_U154, P1_R1105_U155, P1_R1105_U156, P1_R1105_U157, P1_R1105_U158, P1_R1105_U159, P1_R1105_U16, P1_R1105_U160, P1_R1105_U161, P1_R1105_U162, P1_R1105_U163, P1_R1105_U164, P1_R1105_U165, P1_R1105_U166, P1_R1105_U167, P1_R1105_U168, P1_R1105_U169, P1_R1105_U17, P1_R1105_U170, P1_R1105_U171, P1_R1105_U172, P1_R1105_U173, P1_R1105_U174, P1_R1105_U175, P1_R1105_U176, P1_R1105_U177, P1_R1105_U178, P1_R1105_U179, P1_R1105_U18, P1_R1105_U180, P1_R1105_U181, P1_R1105_U182, P1_R1105_U183, P1_R1105_U184, P1_R1105_U185, P1_R1105_U186, P1_R1105_U187, P1_R1105_U188, P1_R1105_U189, P1_R1105_U19, P1_R1105_U190, P1_R1105_U191, P1_R1105_U192, P1_R1105_U193, P1_R1105_U194, P1_R1105_U195, P1_R1105_U196, P1_R1105_U197, P1_R1105_U198, P1_R1105_U199, P1_R1105_U20, P1_R1105_U200, P1_R1105_U201, P1_R1105_U202, P1_R1105_U203, P1_R1105_U204, P1_R1105_U205, P1_R1105_U206, P1_R1105_U207, P1_R1105_U208, P1_R1105_U209, P1_R1105_U21, P1_R1105_U210, P1_R1105_U211, P1_R1105_U212, P1_R1105_U213, P1_R1105_U214, P1_R1105_U215, P1_R1105_U216, P1_R1105_U217, P1_R1105_U218, P1_R1105_U219, P1_R1105_U22, P1_R1105_U220, P1_R1105_U221, P1_R1105_U222, P1_R1105_U223, P1_R1105_U224, P1_R1105_U225, P1_R1105_U226, P1_R1105_U227, P1_R1105_U228, P1_R1105_U229, P1_R1105_U23, P1_R1105_U230, P1_R1105_U231, P1_R1105_U232, P1_R1105_U233, P1_R1105_U234, P1_R1105_U235, P1_R1105_U236, P1_R1105_U237, P1_R1105_U238, P1_R1105_U239, P1_R1105_U24, P1_R1105_U240, P1_R1105_U241, P1_R1105_U242, P1_R1105_U243, P1_R1105_U244, P1_R1105_U245, P1_R1105_U246, P1_R1105_U247, P1_R1105_U248, P1_R1105_U249, P1_R1105_U25, P1_R1105_U250, P1_R1105_U251, P1_R1105_U252, P1_R1105_U253, P1_R1105_U254, P1_R1105_U255, P1_R1105_U256, P1_R1105_U257, P1_R1105_U258, P1_R1105_U259, P1_R1105_U26, P1_R1105_U260, P1_R1105_U261, P1_R1105_U262, P1_R1105_U263, P1_R1105_U264, P1_R1105_U265, P1_R1105_U266, P1_R1105_U267, P1_R1105_U268, P1_R1105_U269, P1_R1105_U27, P1_R1105_U270, P1_R1105_U271, P1_R1105_U272, P1_R1105_U273, P1_R1105_U274, P1_R1105_U275, P1_R1105_U276, P1_R1105_U277, P1_R1105_U278, P1_R1105_U279, P1_R1105_U28, P1_R1105_U280, P1_R1105_U281, P1_R1105_U282, P1_R1105_U283, P1_R1105_U284, P1_R1105_U285, P1_R1105_U286, P1_R1105_U287, P1_R1105_U288, P1_R1105_U289, P1_R1105_U29, P1_R1105_U290, P1_R1105_U291, P1_R1105_U292, P1_R1105_U293, P1_R1105_U294, P1_R1105_U295, P1_R1105_U296, P1_R1105_U297, P1_R1105_U298, P1_R1105_U299, P1_R1105_U30, P1_R1105_U300, P1_R1105_U301, P1_R1105_U302, P1_R1105_U303, P1_R1105_U304, P1_R1105_U305, P1_R1105_U306, P1_R1105_U307, P1_R1105_U308, P1_R1105_U31, P1_R1105_U32, P1_R1105_U33, P1_R1105_U34, P1_R1105_U35, P1_R1105_U36, P1_R1105_U37, P1_R1105_U38, P1_R1105_U39, P1_R1105_U4, P1_R1105_U40, P1_R1105_U41, P1_R1105_U42, P1_R1105_U43, P1_R1105_U44, P1_R1105_U45, P1_R1105_U46, P1_R1105_U47, P1_R1105_U48, P1_R1105_U49, P1_R1105_U5, P1_R1105_U50, P1_R1105_U51, P1_R1105_U52, P1_R1105_U53, P1_R1105_U54, P1_R1105_U55, P1_R1105_U56, P1_R1105_U57, P1_R1105_U58, P1_R1105_U59, P1_R1105_U6, P1_R1105_U60, P1_R1105_U61, P1_R1105_U62, P1_R1105_U63, P1_R1105_U64, P1_R1105_U65, P1_R1105_U66, P1_R1105_U67, P1_R1105_U68, P1_R1105_U69, P1_R1105_U7, P1_R1105_U70, P1_R1105_U71, P1_R1105_U72, P1_R1105_U73, P1_R1105_U74, P1_R1105_U75, P1_R1105_U76, P1_R1105_U77, P1_R1105_U78, P1_R1105_U79, P1_R1105_U8, P1_R1105_U80, P1_R1105_U81, P1_R1105_U82, P1_R1105_U83, P1_R1105_U84, P1_R1105_U85, P1_R1105_U86, P1_R1105_U87, P1_R1105_U88, P1_R1105_U89, P1_R1105_U9, P1_R1105_U90, P1_R1105_U91, P1_R1105_U92, P1_R1105_U93, P1_R1105_U94, P1_R1105_U95, P1_R1105_U96, P1_R1105_U97, P1_R1105_U98, P1_R1105_U99, P1_R1117_U10, P1_R1117_U100, P1_R1117_U101, P1_R1117_U102, P1_R1117_U103, P1_R1117_U104, P1_R1117_U105, P1_R1117_U106, P1_R1117_U107, P1_R1117_U108, P1_R1117_U109, P1_R1117_U11, P1_R1117_U110, P1_R1117_U111, P1_R1117_U112, P1_R1117_U113, P1_R1117_U114, P1_R1117_U115, P1_R1117_U116, P1_R1117_U117, P1_R1117_U118, P1_R1117_U119, P1_R1117_U12, P1_R1117_U120, P1_R1117_U121, P1_R1117_U122, P1_R1117_U123, P1_R1117_U124, P1_R1117_U125, P1_R1117_U126, P1_R1117_U127, P1_R1117_U128, P1_R1117_U129, P1_R1117_U13, P1_R1117_U130, P1_R1117_U131, P1_R1117_U132, P1_R1117_U133, P1_R1117_U134, P1_R1117_U135, P1_R1117_U136, P1_R1117_U137, P1_R1117_U138, P1_R1117_U139, P1_R1117_U14, P1_R1117_U140, P1_R1117_U141, P1_R1117_U142, P1_R1117_U143, P1_R1117_U144, P1_R1117_U145, P1_R1117_U146, P1_R1117_U147, P1_R1117_U148, P1_R1117_U149, P1_R1117_U15, P1_R1117_U150, P1_R1117_U151, P1_R1117_U152, P1_R1117_U153, P1_R1117_U154, P1_R1117_U155, P1_R1117_U156, P1_R1117_U157, P1_R1117_U158, P1_R1117_U159, P1_R1117_U16, P1_R1117_U160, P1_R1117_U161, P1_R1117_U162, P1_R1117_U163, P1_R1117_U164, P1_R1117_U165, P1_R1117_U166, P1_R1117_U167, P1_R1117_U168, P1_R1117_U169, P1_R1117_U17, P1_R1117_U170, P1_R1117_U171, P1_R1117_U172, P1_R1117_U173, P1_R1117_U174, P1_R1117_U175, P1_R1117_U176, P1_R1117_U177, P1_R1117_U178, P1_R1117_U179, P1_R1117_U18, P1_R1117_U180, P1_R1117_U181, P1_R1117_U182, P1_R1117_U183, P1_R1117_U184, P1_R1117_U185, P1_R1117_U186, P1_R1117_U187, P1_R1117_U188, P1_R1117_U189, P1_R1117_U19, P1_R1117_U190, P1_R1117_U191, P1_R1117_U192, P1_R1117_U193, P1_R1117_U194, P1_R1117_U195, P1_R1117_U196, P1_R1117_U197, P1_R1117_U198, P1_R1117_U199, P1_R1117_U20, P1_R1117_U200, P1_R1117_U201, P1_R1117_U202, P1_R1117_U203, P1_R1117_U204, P1_R1117_U205, P1_R1117_U206, P1_R1117_U207, P1_R1117_U208, P1_R1117_U209, P1_R1117_U21, P1_R1117_U210, P1_R1117_U211, P1_R1117_U212, P1_R1117_U213, P1_R1117_U214, P1_R1117_U215, P1_R1117_U216, P1_R1117_U217, P1_R1117_U218, P1_R1117_U219, P1_R1117_U22, P1_R1117_U220, P1_R1117_U221, P1_R1117_U222, P1_R1117_U223, P1_R1117_U224, P1_R1117_U225, P1_R1117_U226, P1_R1117_U227, P1_R1117_U228, P1_R1117_U229, P1_R1117_U23, P1_R1117_U230, P1_R1117_U231, P1_R1117_U232, P1_R1117_U233, P1_R1117_U234, P1_R1117_U235, P1_R1117_U236, P1_R1117_U237, P1_R1117_U238, P1_R1117_U239, P1_R1117_U24, P1_R1117_U240, P1_R1117_U241, P1_R1117_U242, P1_R1117_U243, P1_R1117_U244, P1_R1117_U245, P1_R1117_U246, P1_R1117_U247, P1_R1117_U248, P1_R1117_U249, P1_R1117_U25, P1_R1117_U250, P1_R1117_U251, P1_R1117_U252, P1_R1117_U253, P1_R1117_U254, P1_R1117_U255, P1_R1117_U256, P1_R1117_U257, P1_R1117_U258, P1_R1117_U259, P1_R1117_U26, P1_R1117_U260, P1_R1117_U261, P1_R1117_U262, P1_R1117_U263, P1_R1117_U264, P1_R1117_U265, P1_R1117_U266, P1_R1117_U267, P1_R1117_U268, P1_R1117_U269, P1_R1117_U27, P1_R1117_U270, P1_R1117_U271, P1_R1117_U272, P1_R1117_U273, P1_R1117_U274, P1_R1117_U275, P1_R1117_U276, P1_R1117_U277, P1_R1117_U278, P1_R1117_U279, P1_R1117_U28, P1_R1117_U280, P1_R1117_U281, P1_R1117_U282, P1_R1117_U283, P1_R1117_U284, P1_R1117_U285, P1_R1117_U286, P1_R1117_U287, P1_R1117_U288, P1_R1117_U289, P1_R1117_U29, P1_R1117_U290, P1_R1117_U291, P1_R1117_U292, P1_R1117_U293, P1_R1117_U294, P1_R1117_U295, P1_R1117_U296, P1_R1117_U297, P1_R1117_U298, P1_R1117_U299, P1_R1117_U30, P1_R1117_U300, P1_R1117_U301, P1_R1117_U302, P1_R1117_U303, P1_R1117_U304, P1_R1117_U305, P1_R1117_U306, P1_R1117_U307, P1_R1117_U308, P1_R1117_U309, P1_R1117_U31, P1_R1117_U310, P1_R1117_U311, P1_R1117_U312, P1_R1117_U313, P1_R1117_U314, P1_R1117_U315, P1_R1117_U316, P1_R1117_U317, P1_R1117_U318, P1_R1117_U319, P1_R1117_U32, P1_R1117_U320, P1_R1117_U321, P1_R1117_U322, P1_R1117_U323, P1_R1117_U324, P1_R1117_U325, P1_R1117_U326, P1_R1117_U327, P1_R1117_U328, P1_R1117_U329, P1_R1117_U33, P1_R1117_U330, P1_R1117_U331, P1_R1117_U332, P1_R1117_U333, P1_R1117_U334, P1_R1117_U335, P1_R1117_U336, P1_R1117_U337, P1_R1117_U338, P1_R1117_U339, P1_R1117_U34, P1_R1117_U340, P1_R1117_U341, P1_R1117_U342, P1_R1117_U343, P1_R1117_U344, P1_R1117_U345, P1_R1117_U346, P1_R1117_U347, P1_R1117_U348, P1_R1117_U349, P1_R1117_U35, P1_R1117_U350, P1_R1117_U351, P1_R1117_U352, P1_R1117_U353, P1_R1117_U354, P1_R1117_U355, P1_R1117_U356, P1_R1117_U357, P1_R1117_U358, P1_R1117_U359, P1_R1117_U36, P1_R1117_U360, P1_R1117_U361, P1_R1117_U362, P1_R1117_U363, P1_R1117_U364, P1_R1117_U365, P1_R1117_U366, P1_R1117_U367, P1_R1117_U368, P1_R1117_U369, P1_R1117_U37, P1_R1117_U370, P1_R1117_U371, P1_R1117_U372, P1_R1117_U373, P1_R1117_U374, P1_R1117_U375, P1_R1117_U376, P1_R1117_U377, P1_R1117_U378, P1_R1117_U379, P1_R1117_U38, P1_R1117_U380, P1_R1117_U381, P1_R1117_U382, P1_R1117_U383, P1_R1117_U384, P1_R1117_U385, P1_R1117_U386, P1_R1117_U387, P1_R1117_U388, P1_R1117_U389, P1_R1117_U39, P1_R1117_U390, P1_R1117_U391, P1_R1117_U392, P1_R1117_U393, P1_R1117_U394, P1_R1117_U395, P1_R1117_U396, P1_R1117_U397, P1_R1117_U398, P1_R1117_U399, P1_R1117_U40, P1_R1117_U400, P1_R1117_U401, P1_R1117_U402, P1_R1117_U403, P1_R1117_U404, P1_R1117_U405, P1_R1117_U406, P1_R1117_U407, P1_R1117_U408, P1_R1117_U409, P1_R1117_U41, P1_R1117_U410, P1_R1117_U411, P1_R1117_U412, P1_R1117_U413, P1_R1117_U414, P1_R1117_U415, P1_R1117_U416, P1_R1117_U417, P1_R1117_U418, P1_R1117_U419, P1_R1117_U42, P1_R1117_U420, P1_R1117_U421, P1_R1117_U422, P1_R1117_U423, P1_R1117_U424, P1_R1117_U425, P1_R1117_U426, P1_R1117_U427, P1_R1117_U428, P1_R1117_U429, P1_R1117_U43, P1_R1117_U430, P1_R1117_U431, P1_R1117_U432, P1_R1117_U433, P1_R1117_U434, P1_R1117_U435, P1_R1117_U436, P1_R1117_U437, P1_R1117_U438, P1_R1117_U439, P1_R1117_U44, P1_R1117_U440, P1_R1117_U441, P1_R1117_U442, P1_R1117_U443, P1_R1117_U444, P1_R1117_U445, P1_R1117_U446, P1_R1117_U447, P1_R1117_U448, P1_R1117_U449, P1_R1117_U45, P1_R1117_U450, P1_R1117_U451, P1_R1117_U452, P1_R1117_U453, P1_R1117_U454, P1_R1117_U455, P1_R1117_U456, P1_R1117_U457, P1_R1117_U458, P1_R1117_U459, P1_R1117_U46, P1_R1117_U460, P1_R1117_U461, P1_R1117_U462, P1_R1117_U463, P1_R1117_U464, P1_R1117_U465, P1_R1117_U466, P1_R1117_U467, P1_R1117_U468, P1_R1117_U469, P1_R1117_U47, P1_R1117_U470, P1_R1117_U471, P1_R1117_U472, P1_R1117_U473, P1_R1117_U48, P1_R1117_U49, P1_R1117_U50, P1_R1117_U51, P1_R1117_U52, P1_R1117_U53, P1_R1117_U54, P1_R1117_U55, P1_R1117_U56, P1_R1117_U57, P1_R1117_U58, P1_R1117_U59, P1_R1117_U6, P1_R1117_U60, P1_R1117_U61, P1_R1117_U62, P1_R1117_U63, P1_R1117_U64, P1_R1117_U65, P1_R1117_U66, P1_R1117_U67, P1_R1117_U68, P1_R1117_U69, P1_R1117_U7, P1_R1117_U70, P1_R1117_U71, P1_R1117_U72, P1_R1117_U73, P1_R1117_U74, P1_R1117_U75, P1_R1117_U76, P1_R1117_U77, P1_R1117_U78, P1_R1117_U79, P1_R1117_U8, P1_R1117_U80, P1_R1117_U81, P1_R1117_U82, P1_R1117_U83, P1_R1117_U84, P1_R1117_U85, P1_R1117_U86, P1_R1117_U87, P1_R1117_U88, P1_R1117_U89, P1_R1117_U9, P1_R1117_U90, P1_R1117_U91, P1_R1117_U92, P1_R1117_U93, P1_R1117_U94, P1_R1117_U95, P1_R1117_U96, P1_R1117_U97, P1_R1117_U98, P1_R1117_U99, P1_R1138_U10, P1_R1138_U100, P1_R1138_U101, P1_R1138_U102, P1_R1138_U103, P1_R1138_U104, P1_R1138_U105, P1_R1138_U106, P1_R1138_U107, P1_R1138_U108, P1_R1138_U109, P1_R1138_U11, P1_R1138_U110, P1_R1138_U111, P1_R1138_U112, P1_R1138_U113, P1_R1138_U114, P1_R1138_U115, P1_R1138_U116, P1_R1138_U117, P1_R1138_U118, P1_R1138_U119, P1_R1138_U12, P1_R1138_U120, P1_R1138_U121, P1_R1138_U122, P1_R1138_U123, P1_R1138_U124, P1_R1138_U125, P1_R1138_U126, P1_R1138_U127, P1_R1138_U128, P1_R1138_U129, P1_R1138_U13, P1_R1138_U130, P1_R1138_U131, P1_R1138_U132, P1_R1138_U133, P1_R1138_U134, P1_R1138_U135, P1_R1138_U136, P1_R1138_U137, P1_R1138_U138, P1_R1138_U139, P1_R1138_U14, P1_R1138_U140, P1_R1138_U141, P1_R1138_U142, P1_R1138_U143, P1_R1138_U144, P1_R1138_U145, P1_R1138_U146, P1_R1138_U147, P1_R1138_U148, P1_R1138_U149, P1_R1138_U15, P1_R1138_U150, P1_R1138_U151, P1_R1138_U152, P1_R1138_U153, P1_R1138_U154, P1_R1138_U155, P1_R1138_U156, P1_R1138_U157, P1_R1138_U158, P1_R1138_U159, P1_R1138_U16, P1_R1138_U160, P1_R1138_U161, P1_R1138_U162, P1_R1138_U163, P1_R1138_U164, P1_R1138_U165, P1_R1138_U166, P1_R1138_U167, P1_R1138_U168, P1_R1138_U169, P1_R1138_U17, P1_R1138_U170, P1_R1138_U171, P1_R1138_U172, P1_R1138_U173, P1_R1138_U174, P1_R1138_U175, P1_R1138_U176, P1_R1138_U177, P1_R1138_U178, P1_R1138_U179, P1_R1138_U18, P1_R1138_U180, P1_R1138_U181, P1_R1138_U182, P1_R1138_U183, P1_R1138_U184, P1_R1138_U185, P1_R1138_U186, P1_R1138_U187, P1_R1138_U188, P1_R1138_U189, P1_R1138_U19, P1_R1138_U190, P1_R1138_U191, P1_R1138_U192, P1_R1138_U193, P1_R1138_U194, P1_R1138_U195, P1_R1138_U196, P1_R1138_U197, P1_R1138_U198, P1_R1138_U199, P1_R1138_U20, P1_R1138_U200, P1_R1138_U201, P1_R1138_U202, P1_R1138_U203, P1_R1138_U204, P1_R1138_U205, P1_R1138_U206, P1_R1138_U207, P1_R1138_U208, P1_R1138_U209, P1_R1138_U21, P1_R1138_U210, P1_R1138_U211, P1_R1138_U212, P1_R1138_U213, P1_R1138_U214, P1_R1138_U215, P1_R1138_U216, P1_R1138_U217, P1_R1138_U218, P1_R1138_U219, P1_R1138_U22, P1_R1138_U220, P1_R1138_U221, P1_R1138_U222, P1_R1138_U223, P1_R1138_U224, P1_R1138_U225, P1_R1138_U226, P1_R1138_U227, P1_R1138_U228, P1_R1138_U229, P1_R1138_U23, P1_R1138_U230, P1_R1138_U231, P1_R1138_U232, P1_R1138_U233, P1_R1138_U234, P1_R1138_U235, P1_R1138_U236, P1_R1138_U237, P1_R1138_U238, P1_R1138_U239, P1_R1138_U24, P1_R1138_U240, P1_R1138_U241, P1_R1138_U242, P1_R1138_U243, P1_R1138_U244, P1_R1138_U245, P1_R1138_U246, P1_R1138_U247, P1_R1138_U248, P1_R1138_U249, P1_R1138_U25, P1_R1138_U250, P1_R1138_U251, P1_R1138_U252, P1_R1138_U253, P1_R1138_U254, P1_R1138_U255, P1_R1138_U256, P1_R1138_U257, P1_R1138_U258, P1_R1138_U259, P1_R1138_U26, P1_R1138_U260, P1_R1138_U261, P1_R1138_U262, P1_R1138_U263, P1_R1138_U264, P1_R1138_U265, P1_R1138_U266, P1_R1138_U267, P1_R1138_U268, P1_R1138_U269, P1_R1138_U27, P1_R1138_U270, P1_R1138_U271, P1_R1138_U272, P1_R1138_U273, P1_R1138_U274, P1_R1138_U275, P1_R1138_U276, P1_R1138_U277, P1_R1138_U278, P1_R1138_U279, P1_R1138_U28, P1_R1138_U280, P1_R1138_U281, P1_R1138_U282, P1_R1138_U283, P1_R1138_U284, P1_R1138_U285, P1_R1138_U286, P1_R1138_U287, P1_R1138_U288, P1_R1138_U289, P1_R1138_U29, P1_R1138_U290, P1_R1138_U291, P1_R1138_U292, P1_R1138_U293, P1_R1138_U294, P1_R1138_U295, P1_R1138_U296, P1_R1138_U297, P1_R1138_U298, P1_R1138_U299, P1_R1138_U30, P1_R1138_U300, P1_R1138_U301, P1_R1138_U302, P1_R1138_U303, P1_R1138_U304, P1_R1138_U305, P1_R1138_U306, P1_R1138_U307, P1_R1138_U308, P1_R1138_U309, P1_R1138_U31, P1_R1138_U310, P1_R1138_U311, P1_R1138_U312, P1_R1138_U313, P1_R1138_U314, P1_R1138_U315, P1_R1138_U316, P1_R1138_U317, P1_R1138_U318, P1_R1138_U319, P1_R1138_U32, P1_R1138_U320, P1_R1138_U321, P1_R1138_U322, P1_R1138_U323, P1_R1138_U324, P1_R1138_U325, P1_R1138_U326, P1_R1138_U327, P1_R1138_U328, P1_R1138_U329, P1_R1138_U33, P1_R1138_U330, P1_R1138_U331, P1_R1138_U332, P1_R1138_U333, P1_R1138_U334, P1_R1138_U335, P1_R1138_U336, P1_R1138_U337, P1_R1138_U338, P1_R1138_U339, P1_R1138_U34, P1_R1138_U340, P1_R1138_U341, P1_R1138_U342, P1_R1138_U343, P1_R1138_U344, P1_R1138_U345, P1_R1138_U346, P1_R1138_U347, P1_R1138_U348, P1_R1138_U349, P1_R1138_U35, P1_R1138_U350, P1_R1138_U351, P1_R1138_U352, P1_R1138_U353, P1_R1138_U354, P1_R1138_U355, P1_R1138_U356, P1_R1138_U357, P1_R1138_U358, P1_R1138_U359, P1_R1138_U36, P1_R1138_U360, P1_R1138_U361, P1_R1138_U362, P1_R1138_U363, P1_R1138_U364, P1_R1138_U365, P1_R1138_U366, P1_R1138_U367, P1_R1138_U368, P1_R1138_U369, P1_R1138_U37, P1_R1138_U370, P1_R1138_U371, P1_R1138_U372, P1_R1138_U373, P1_R1138_U374, P1_R1138_U375, P1_R1138_U376, P1_R1138_U377, P1_R1138_U378, P1_R1138_U379, P1_R1138_U38, P1_R1138_U380, P1_R1138_U381, P1_R1138_U382, P1_R1138_U383, P1_R1138_U384, P1_R1138_U385, P1_R1138_U386, P1_R1138_U387, P1_R1138_U388, P1_R1138_U389, P1_R1138_U39, P1_R1138_U390, P1_R1138_U391, P1_R1138_U392, P1_R1138_U393, P1_R1138_U394, P1_R1138_U395, P1_R1138_U396, P1_R1138_U397, P1_R1138_U398, P1_R1138_U399, P1_R1138_U4, P1_R1138_U40, P1_R1138_U400, P1_R1138_U401, P1_R1138_U402, P1_R1138_U403, P1_R1138_U404, P1_R1138_U405, P1_R1138_U406, P1_R1138_U407, P1_R1138_U408, P1_R1138_U409, P1_R1138_U41, P1_R1138_U410, P1_R1138_U411, P1_R1138_U412, P1_R1138_U413, P1_R1138_U414, P1_R1138_U415, P1_R1138_U416, P1_R1138_U417, P1_R1138_U418, P1_R1138_U419, P1_R1138_U42, P1_R1138_U420, P1_R1138_U421, P1_R1138_U422, P1_R1138_U423, P1_R1138_U424, P1_R1138_U425, P1_R1138_U426, P1_R1138_U427, P1_R1138_U428, P1_R1138_U429, P1_R1138_U43, P1_R1138_U430, P1_R1138_U431, P1_R1138_U432, P1_R1138_U433, P1_R1138_U434, P1_R1138_U435, P1_R1138_U436, P1_R1138_U437, P1_R1138_U438, P1_R1138_U439, P1_R1138_U44, P1_R1138_U440, P1_R1138_U441, P1_R1138_U442, P1_R1138_U443, P1_R1138_U444, P1_R1138_U445, P1_R1138_U446, P1_R1138_U447, P1_R1138_U448, P1_R1138_U449, P1_R1138_U45, P1_R1138_U450, P1_R1138_U451, P1_R1138_U452, P1_R1138_U453, P1_R1138_U454, P1_R1138_U455, P1_R1138_U456, P1_R1138_U457, P1_R1138_U458, P1_R1138_U459, P1_R1138_U46, P1_R1138_U460, P1_R1138_U461, P1_R1138_U462, P1_R1138_U463, P1_R1138_U464, P1_R1138_U465, P1_R1138_U466, P1_R1138_U467, P1_R1138_U468, P1_R1138_U469, P1_R1138_U47, P1_R1138_U470, P1_R1138_U471, P1_R1138_U472, P1_R1138_U473, P1_R1138_U474, P1_R1138_U475, P1_R1138_U476, P1_R1138_U477, P1_R1138_U478, P1_R1138_U479, P1_R1138_U48, P1_R1138_U480, P1_R1138_U481, P1_R1138_U482, P1_R1138_U483, P1_R1138_U484, P1_R1138_U485, P1_R1138_U486, P1_R1138_U487, P1_R1138_U488, P1_R1138_U489, P1_R1138_U49, P1_R1138_U490, P1_R1138_U491, P1_R1138_U492, P1_R1138_U493, P1_R1138_U494, P1_R1138_U495, P1_R1138_U496, P1_R1138_U497, P1_R1138_U498, P1_R1138_U499, P1_R1138_U5, P1_R1138_U50, P1_R1138_U500, P1_R1138_U501, P1_R1138_U502, P1_R1138_U503, P1_R1138_U51, P1_R1138_U52, P1_R1138_U53, P1_R1138_U54, P1_R1138_U55, P1_R1138_U56, P1_R1138_U57, P1_R1138_U58, P1_R1138_U59, P1_R1138_U6, P1_R1138_U60, P1_R1138_U61, P1_R1138_U62, P1_R1138_U63, P1_R1138_U64, P1_R1138_U65, P1_R1138_U66, P1_R1138_U67, P1_R1138_U68, P1_R1138_U69, P1_R1138_U7, P1_R1138_U70, P1_R1138_U71, P1_R1138_U72, P1_R1138_U73, P1_R1138_U74, P1_R1138_U75, P1_R1138_U76, P1_R1138_U77, P1_R1138_U78, P1_R1138_U79, P1_R1138_U8, P1_R1138_U80, P1_R1138_U81, P1_R1138_U82, P1_R1138_U83, P1_R1138_U84, P1_R1138_U85, P1_R1138_U86, P1_R1138_U87, P1_R1138_U88, P1_R1138_U89, P1_R1138_U9, P1_R1138_U90, P1_R1138_U91, P1_R1138_U92, P1_R1138_U93, P1_R1138_U94, P1_R1138_U95, P1_R1138_U96, P1_R1138_U97, P1_R1138_U98, P1_R1138_U99, P1_R1150_U10, P1_R1150_U100, P1_R1150_U101, P1_R1150_U102, P1_R1150_U103, P1_R1150_U104, P1_R1150_U105, P1_R1150_U106, P1_R1150_U107, P1_R1150_U108, P1_R1150_U109, P1_R1150_U11, P1_R1150_U110, P1_R1150_U111, P1_R1150_U112, P1_R1150_U113, P1_R1150_U114, P1_R1150_U115, P1_R1150_U116, P1_R1150_U117, P1_R1150_U118, P1_R1150_U119, P1_R1150_U12, P1_R1150_U120, P1_R1150_U121, P1_R1150_U122, P1_R1150_U123, P1_R1150_U124, P1_R1150_U125, P1_R1150_U126, P1_R1150_U127, P1_R1150_U128, P1_R1150_U129, P1_R1150_U13, P1_R1150_U130, P1_R1150_U131, P1_R1150_U132, P1_R1150_U133, P1_R1150_U134, P1_R1150_U135, P1_R1150_U136, P1_R1150_U137, P1_R1150_U138, P1_R1150_U139, P1_R1150_U14, P1_R1150_U140, P1_R1150_U141, P1_R1150_U142, P1_R1150_U143, P1_R1150_U144, P1_R1150_U145, P1_R1150_U146, P1_R1150_U147, P1_R1150_U148, P1_R1150_U149, P1_R1150_U15, P1_R1150_U150, P1_R1150_U151, P1_R1150_U152, P1_R1150_U153, P1_R1150_U154, P1_R1150_U155, P1_R1150_U156, P1_R1150_U157, P1_R1150_U158, P1_R1150_U159, P1_R1150_U16, P1_R1150_U160, P1_R1150_U161, P1_R1150_U162, P1_R1150_U163, P1_R1150_U164, P1_R1150_U165, P1_R1150_U166, P1_R1150_U167, P1_R1150_U168, P1_R1150_U169, P1_R1150_U17, P1_R1150_U170, P1_R1150_U171, P1_R1150_U172, P1_R1150_U173, P1_R1150_U174, P1_R1150_U175, P1_R1150_U176, P1_R1150_U177, P1_R1150_U178, P1_R1150_U179, P1_R1150_U18, P1_R1150_U180, P1_R1150_U181, P1_R1150_U182, P1_R1150_U183, P1_R1150_U184, P1_R1150_U185, P1_R1150_U186, P1_R1150_U187, P1_R1150_U188, P1_R1150_U189, P1_R1150_U19, P1_R1150_U190, P1_R1150_U191, P1_R1150_U192, P1_R1150_U193, P1_R1150_U194, P1_R1150_U195, P1_R1150_U196, P1_R1150_U197, P1_R1150_U198, P1_R1150_U199, P1_R1150_U20, P1_R1150_U200, P1_R1150_U201, P1_R1150_U202, P1_R1150_U203, P1_R1150_U204, P1_R1150_U205, P1_R1150_U206, P1_R1150_U207, P1_R1150_U208, P1_R1150_U209, P1_R1150_U21, P1_R1150_U210, P1_R1150_U211, P1_R1150_U212, P1_R1150_U213, P1_R1150_U214, P1_R1150_U215, P1_R1150_U216, P1_R1150_U217, P1_R1150_U218, P1_R1150_U219, P1_R1150_U22, P1_R1150_U220, P1_R1150_U221, P1_R1150_U222, P1_R1150_U223, P1_R1150_U224, P1_R1150_U225, P1_R1150_U226, P1_R1150_U227, P1_R1150_U228, P1_R1150_U229, P1_R1150_U23, P1_R1150_U230, P1_R1150_U231, P1_R1150_U232, P1_R1150_U233, P1_R1150_U234, P1_R1150_U235, P1_R1150_U236, P1_R1150_U237, P1_R1150_U238, P1_R1150_U239, P1_R1150_U24, P1_R1150_U240, P1_R1150_U241, P1_R1150_U242, P1_R1150_U243, P1_R1150_U244, P1_R1150_U245, P1_R1150_U246, P1_R1150_U247, P1_R1150_U248, P1_R1150_U249, P1_R1150_U25, P1_R1150_U250, P1_R1150_U251, P1_R1150_U252, P1_R1150_U253, P1_R1150_U254, P1_R1150_U255, P1_R1150_U256, P1_R1150_U257, P1_R1150_U258, P1_R1150_U259, P1_R1150_U26, P1_R1150_U260, P1_R1150_U261, P1_R1150_U262, P1_R1150_U263, P1_R1150_U264, P1_R1150_U265, P1_R1150_U266, P1_R1150_U267, P1_R1150_U268, P1_R1150_U269, P1_R1150_U27, P1_R1150_U270, P1_R1150_U271, P1_R1150_U272, P1_R1150_U273, P1_R1150_U274, P1_R1150_U275, P1_R1150_U276, P1_R1150_U277, P1_R1150_U278, P1_R1150_U279, P1_R1150_U28, P1_R1150_U280, P1_R1150_U281, P1_R1150_U282, P1_R1150_U283, P1_R1150_U284, P1_R1150_U285, P1_R1150_U286, P1_R1150_U287, P1_R1150_U288, P1_R1150_U289, P1_R1150_U29, P1_R1150_U290, P1_R1150_U291, P1_R1150_U292, P1_R1150_U293, P1_R1150_U294, P1_R1150_U295, P1_R1150_U296, P1_R1150_U297, P1_R1150_U298, P1_R1150_U299, P1_R1150_U30, P1_R1150_U300, P1_R1150_U301, P1_R1150_U302, P1_R1150_U303, P1_R1150_U304, P1_R1150_U305, P1_R1150_U306, P1_R1150_U307, P1_R1150_U308, P1_R1150_U309, P1_R1150_U31, P1_R1150_U310, P1_R1150_U311, P1_R1150_U312, P1_R1150_U313, P1_R1150_U314, P1_R1150_U315, P1_R1150_U316, P1_R1150_U317, P1_R1150_U318, P1_R1150_U319, P1_R1150_U32, P1_R1150_U320, P1_R1150_U321, P1_R1150_U322, P1_R1150_U323, P1_R1150_U324, P1_R1150_U325, P1_R1150_U326, P1_R1150_U327, P1_R1150_U328, P1_R1150_U329, P1_R1150_U33, P1_R1150_U330, P1_R1150_U331, P1_R1150_U332, P1_R1150_U333, P1_R1150_U334, P1_R1150_U335, P1_R1150_U336, P1_R1150_U337, P1_R1150_U338, P1_R1150_U339, P1_R1150_U34, P1_R1150_U340, P1_R1150_U341, P1_R1150_U342, P1_R1150_U343, P1_R1150_U344, P1_R1150_U345, P1_R1150_U346, P1_R1150_U347, P1_R1150_U348, P1_R1150_U349, P1_R1150_U35, P1_R1150_U350, P1_R1150_U351, P1_R1150_U352, P1_R1150_U353, P1_R1150_U354, P1_R1150_U355, P1_R1150_U356, P1_R1150_U357, P1_R1150_U358, P1_R1150_U359, P1_R1150_U36, P1_R1150_U360, P1_R1150_U361, P1_R1150_U362, P1_R1150_U363, P1_R1150_U364, P1_R1150_U365, P1_R1150_U366, P1_R1150_U367, P1_R1150_U368, P1_R1150_U369, P1_R1150_U37, P1_R1150_U370, P1_R1150_U371, P1_R1150_U372, P1_R1150_U373, P1_R1150_U374, P1_R1150_U375, P1_R1150_U376, P1_R1150_U377, P1_R1150_U378, P1_R1150_U379, P1_R1150_U38, P1_R1150_U380, P1_R1150_U381, P1_R1150_U382, P1_R1150_U383, P1_R1150_U384, P1_R1150_U385, P1_R1150_U386, P1_R1150_U387, P1_R1150_U388, P1_R1150_U389, P1_R1150_U39, P1_R1150_U390, P1_R1150_U391, P1_R1150_U392, P1_R1150_U393, P1_R1150_U394, P1_R1150_U395, P1_R1150_U396, P1_R1150_U397, P1_R1150_U398, P1_R1150_U399, P1_R1150_U40, P1_R1150_U400, P1_R1150_U401, P1_R1150_U402, P1_R1150_U403, P1_R1150_U404, P1_R1150_U405, P1_R1150_U406, P1_R1150_U407, P1_R1150_U408, P1_R1150_U409, P1_R1150_U41, P1_R1150_U410, P1_R1150_U411, P1_R1150_U412, P1_R1150_U413, P1_R1150_U414, P1_R1150_U415, P1_R1150_U416, P1_R1150_U417, P1_R1150_U418, P1_R1150_U419, P1_R1150_U42, P1_R1150_U420, P1_R1150_U421, P1_R1150_U422, P1_R1150_U423, P1_R1150_U424, P1_R1150_U425, P1_R1150_U426, P1_R1150_U427, P1_R1150_U428, P1_R1150_U429, P1_R1150_U43, P1_R1150_U430, P1_R1150_U431, P1_R1150_U432, P1_R1150_U433, P1_R1150_U434, P1_R1150_U435, P1_R1150_U436, P1_R1150_U437, P1_R1150_U438, P1_R1150_U439, P1_R1150_U44, P1_R1150_U440, P1_R1150_U441, P1_R1150_U442, P1_R1150_U443, P1_R1150_U444, P1_R1150_U445, P1_R1150_U446, P1_R1150_U447, P1_R1150_U448, P1_R1150_U449, P1_R1150_U45, P1_R1150_U450, P1_R1150_U451, P1_R1150_U452, P1_R1150_U453, P1_R1150_U454, P1_R1150_U455, P1_R1150_U456, P1_R1150_U457, P1_R1150_U458, P1_R1150_U459, P1_R1150_U46, P1_R1150_U460, P1_R1150_U461, P1_R1150_U462, P1_R1150_U463, P1_R1150_U464, P1_R1150_U465, P1_R1150_U466, P1_R1150_U467, P1_R1150_U468, P1_R1150_U469, P1_R1150_U47, P1_R1150_U470, P1_R1150_U471, P1_R1150_U472, P1_R1150_U473, P1_R1150_U48, P1_R1150_U49, P1_R1150_U50, P1_R1150_U51, P1_R1150_U52, P1_R1150_U53, P1_R1150_U54, P1_R1150_U55, P1_R1150_U56, P1_R1150_U57, P1_R1150_U58, P1_R1150_U59, P1_R1150_U6, P1_R1150_U60, P1_R1150_U61, P1_R1150_U62, P1_R1150_U63, P1_R1150_U64, P1_R1150_U65, P1_R1150_U66, P1_R1150_U67, P1_R1150_U68, P1_R1150_U69, P1_R1150_U7, P1_R1150_U70, P1_R1150_U71, P1_R1150_U72, P1_R1150_U73, P1_R1150_U74, P1_R1150_U75, P1_R1150_U76, P1_R1150_U77, P1_R1150_U78, P1_R1150_U79, P1_R1150_U8, P1_R1150_U80, P1_R1150_U81, P1_R1150_U82, P1_R1150_U83, P1_R1150_U84, P1_R1150_U85, P1_R1150_U86, P1_R1150_U87, P1_R1150_U88, P1_R1150_U89, P1_R1150_U9, P1_R1150_U90, P1_R1150_U91, P1_R1150_U92, P1_R1150_U93, P1_R1150_U94, P1_R1150_U95, P1_R1150_U96, P1_R1150_U97, P1_R1150_U98, P1_R1150_U99, P1_R1162_U10, P1_R1162_U100, P1_R1162_U101, P1_R1162_U102, P1_R1162_U103, P1_R1162_U104, P1_R1162_U105, P1_R1162_U106, P1_R1162_U107, P1_R1162_U108, P1_R1162_U109, P1_R1162_U11, P1_R1162_U110, P1_R1162_U111, P1_R1162_U112, P1_R1162_U113, P1_R1162_U114, P1_R1162_U115, P1_R1162_U116, P1_R1162_U117, P1_R1162_U118, P1_R1162_U119, P1_R1162_U12, P1_R1162_U120, P1_R1162_U121, P1_R1162_U122, P1_R1162_U123, P1_R1162_U124, P1_R1162_U125, P1_R1162_U126, P1_R1162_U127, P1_R1162_U128, P1_R1162_U129, P1_R1162_U13, P1_R1162_U130, P1_R1162_U131, P1_R1162_U132, P1_R1162_U133, P1_R1162_U134, P1_R1162_U135, P1_R1162_U136, P1_R1162_U137, P1_R1162_U138, P1_R1162_U139, P1_R1162_U14, P1_R1162_U140, P1_R1162_U141, P1_R1162_U142, P1_R1162_U143, P1_R1162_U144, P1_R1162_U145, P1_R1162_U146, P1_R1162_U147, P1_R1162_U148, P1_R1162_U149, P1_R1162_U15, P1_R1162_U150, P1_R1162_U151, P1_R1162_U152, P1_R1162_U153, P1_R1162_U154, P1_R1162_U155, P1_R1162_U156, P1_R1162_U157, P1_R1162_U158, P1_R1162_U159, P1_R1162_U16, P1_R1162_U160, P1_R1162_U161, P1_R1162_U162, P1_R1162_U163, P1_R1162_U164, P1_R1162_U165, P1_R1162_U166, P1_R1162_U167, P1_R1162_U168, P1_R1162_U169, P1_R1162_U17, P1_R1162_U170, P1_R1162_U171, P1_R1162_U172, P1_R1162_U173, P1_R1162_U174, P1_R1162_U175, P1_R1162_U176, P1_R1162_U177, P1_R1162_U178, P1_R1162_U179, P1_R1162_U18, P1_R1162_U180, P1_R1162_U181, P1_R1162_U182, P1_R1162_U183, P1_R1162_U184, P1_R1162_U185, P1_R1162_U186, P1_R1162_U187, P1_R1162_U188, P1_R1162_U189, P1_R1162_U19, P1_R1162_U190, P1_R1162_U191, P1_R1162_U192, P1_R1162_U193, P1_R1162_U194, P1_R1162_U195, P1_R1162_U196, P1_R1162_U197, P1_R1162_U198, P1_R1162_U199, P1_R1162_U20, P1_R1162_U200, P1_R1162_U201, P1_R1162_U202, P1_R1162_U203, P1_R1162_U204, P1_R1162_U205, P1_R1162_U206, P1_R1162_U207, P1_R1162_U208, P1_R1162_U209, P1_R1162_U21, P1_R1162_U210, P1_R1162_U211, P1_R1162_U212, P1_R1162_U213, P1_R1162_U214, P1_R1162_U215, P1_R1162_U216, P1_R1162_U217, P1_R1162_U218, P1_R1162_U219, P1_R1162_U22, P1_R1162_U220, P1_R1162_U221, P1_R1162_U222, P1_R1162_U223, P1_R1162_U224, P1_R1162_U225, P1_R1162_U226, P1_R1162_U227, P1_R1162_U228, P1_R1162_U229, P1_R1162_U23, P1_R1162_U230, P1_R1162_U231, P1_R1162_U232, P1_R1162_U233, P1_R1162_U234, P1_R1162_U235, P1_R1162_U236, P1_R1162_U237, P1_R1162_U238, P1_R1162_U239, P1_R1162_U24, P1_R1162_U240, P1_R1162_U241, P1_R1162_U242, P1_R1162_U243, P1_R1162_U244, P1_R1162_U245, P1_R1162_U246, P1_R1162_U247, P1_R1162_U248, P1_R1162_U249, P1_R1162_U25, P1_R1162_U250, P1_R1162_U251, P1_R1162_U252, P1_R1162_U253, P1_R1162_U254, P1_R1162_U255, P1_R1162_U256, P1_R1162_U257, P1_R1162_U258, P1_R1162_U259, P1_R1162_U26, P1_R1162_U260, P1_R1162_U261, P1_R1162_U262, P1_R1162_U263, P1_R1162_U264, P1_R1162_U265, P1_R1162_U266, P1_R1162_U267, P1_R1162_U268, P1_R1162_U269, P1_R1162_U27, P1_R1162_U270, P1_R1162_U271, P1_R1162_U272, P1_R1162_U273, P1_R1162_U274, P1_R1162_U275, P1_R1162_U276, P1_R1162_U277, P1_R1162_U278, P1_R1162_U279, P1_R1162_U28, P1_R1162_U280, P1_R1162_U281, P1_R1162_U282, P1_R1162_U283, P1_R1162_U284, P1_R1162_U285, P1_R1162_U286, P1_R1162_U287, P1_R1162_U288, P1_R1162_U289, P1_R1162_U29, P1_R1162_U290, P1_R1162_U291, P1_R1162_U292, P1_R1162_U293, P1_R1162_U294, P1_R1162_U295, P1_R1162_U296, P1_R1162_U297, P1_R1162_U298, P1_R1162_U299, P1_R1162_U30, P1_R1162_U300, P1_R1162_U301, P1_R1162_U302, P1_R1162_U303, P1_R1162_U304, P1_R1162_U305, P1_R1162_U306, P1_R1162_U307, P1_R1162_U308, P1_R1162_U31, P1_R1162_U32, P1_R1162_U33, P1_R1162_U34, P1_R1162_U35, P1_R1162_U36, P1_R1162_U37, P1_R1162_U38, P1_R1162_U39, P1_R1162_U4, P1_R1162_U40, P1_R1162_U41, P1_R1162_U42, P1_R1162_U43, P1_R1162_U44, P1_R1162_U45, P1_R1162_U46, P1_R1162_U47, P1_R1162_U48, P1_R1162_U49, P1_R1162_U5, P1_R1162_U50, P1_R1162_U51, P1_R1162_U52, P1_R1162_U53, P1_R1162_U54, P1_R1162_U55, P1_R1162_U56, P1_R1162_U57, P1_R1162_U58, P1_R1162_U59, P1_R1162_U6, P1_R1162_U60, P1_R1162_U61, P1_R1162_U62, P1_R1162_U63, P1_R1162_U64, P1_R1162_U65, P1_R1162_U66, P1_R1162_U67, P1_R1162_U68, P1_R1162_U69, P1_R1162_U7, P1_R1162_U70, P1_R1162_U71, P1_R1162_U72, P1_R1162_U73, P1_R1162_U74, P1_R1162_U75, P1_R1162_U76, P1_R1162_U77, P1_R1162_U78, P1_R1162_U79, P1_R1162_U8, P1_R1162_U80, P1_R1162_U81, P1_R1162_U82, P1_R1162_U83, P1_R1162_U84, P1_R1162_U85, P1_R1162_U86, P1_R1162_U87, P1_R1162_U88, P1_R1162_U89, P1_R1162_U9, P1_R1162_U90, P1_R1162_U91, P1_R1162_U92, P1_R1162_U93, P1_R1162_U94, P1_R1162_U95, P1_R1162_U96, P1_R1162_U97, P1_R1162_U98, P1_R1162_U99, P1_R1165_U10, P1_R1165_U100, P1_R1165_U101, P1_R1165_U102, P1_R1165_U103, P1_R1165_U104, P1_R1165_U105, P1_R1165_U106, P1_R1165_U107, P1_R1165_U108, P1_R1165_U109, P1_R1165_U11, P1_R1165_U110, P1_R1165_U111, P1_R1165_U112, P1_R1165_U113, P1_R1165_U114, P1_R1165_U115, P1_R1165_U116, P1_R1165_U117, P1_R1165_U118, P1_R1165_U119, P1_R1165_U12, P1_R1165_U120, P1_R1165_U121, P1_R1165_U122, P1_R1165_U123, P1_R1165_U124, P1_R1165_U125, P1_R1165_U126, P1_R1165_U127, P1_R1165_U128, P1_R1165_U129, P1_R1165_U13, P1_R1165_U130, P1_R1165_U131, P1_R1165_U132, P1_R1165_U133, P1_R1165_U134, P1_R1165_U135, P1_R1165_U136, P1_R1165_U137, P1_R1165_U138, P1_R1165_U139, P1_R1165_U14, P1_R1165_U140, P1_R1165_U141, P1_R1165_U142, P1_R1165_U143, P1_R1165_U144, P1_R1165_U145, P1_R1165_U146, P1_R1165_U147, P1_R1165_U148, P1_R1165_U149, P1_R1165_U15, P1_R1165_U150, P1_R1165_U151, P1_R1165_U152, P1_R1165_U153, P1_R1165_U154, P1_R1165_U155, P1_R1165_U156, P1_R1165_U157, P1_R1165_U158, P1_R1165_U159, P1_R1165_U16, P1_R1165_U160, P1_R1165_U161, P1_R1165_U162, P1_R1165_U163, P1_R1165_U164, P1_R1165_U165, P1_R1165_U166, P1_R1165_U167, P1_R1165_U168, P1_R1165_U169, P1_R1165_U17, P1_R1165_U170, P1_R1165_U171, P1_R1165_U172, P1_R1165_U173, P1_R1165_U174, P1_R1165_U175, P1_R1165_U176, P1_R1165_U177, P1_R1165_U178, P1_R1165_U179, P1_R1165_U18, P1_R1165_U180, P1_R1165_U181, P1_R1165_U182, P1_R1165_U183, P1_R1165_U184, P1_R1165_U185, P1_R1165_U186, P1_R1165_U187, P1_R1165_U188, P1_R1165_U189, P1_R1165_U19, P1_R1165_U190, P1_R1165_U191, P1_R1165_U192, P1_R1165_U193, P1_R1165_U194, P1_R1165_U195, P1_R1165_U196, P1_R1165_U197, P1_R1165_U198, P1_R1165_U199, P1_R1165_U20, P1_R1165_U200, P1_R1165_U201, P1_R1165_U202, P1_R1165_U203, P1_R1165_U204, P1_R1165_U205, P1_R1165_U206, P1_R1165_U207, P1_R1165_U208, P1_R1165_U209, P1_R1165_U21, P1_R1165_U210, P1_R1165_U211, P1_R1165_U212, P1_R1165_U213, P1_R1165_U214, P1_R1165_U215, P1_R1165_U216, P1_R1165_U217, P1_R1165_U218, P1_R1165_U219, P1_R1165_U22, P1_R1165_U220, P1_R1165_U221, P1_R1165_U222, P1_R1165_U223, P1_R1165_U224, P1_R1165_U225, P1_R1165_U226, P1_R1165_U227, P1_R1165_U228, P1_R1165_U229, P1_R1165_U23, P1_R1165_U230, P1_R1165_U231, P1_R1165_U232, P1_R1165_U233, P1_R1165_U234, P1_R1165_U235, P1_R1165_U236, P1_R1165_U237, P1_R1165_U238, P1_R1165_U239, P1_R1165_U24, P1_R1165_U240, P1_R1165_U241, P1_R1165_U242, P1_R1165_U243, P1_R1165_U244, P1_R1165_U245, P1_R1165_U246, P1_R1165_U247, P1_R1165_U248, P1_R1165_U249, P1_R1165_U25, P1_R1165_U250, P1_R1165_U251, P1_R1165_U252, P1_R1165_U253, P1_R1165_U254, P1_R1165_U255, P1_R1165_U256, P1_R1165_U257, P1_R1165_U258, P1_R1165_U259, P1_R1165_U26, P1_R1165_U260, P1_R1165_U261, P1_R1165_U262, P1_R1165_U263, P1_R1165_U264, P1_R1165_U265, P1_R1165_U266, P1_R1165_U267, P1_R1165_U268, P1_R1165_U269, P1_R1165_U27, P1_R1165_U270, P1_R1165_U271, P1_R1165_U272, P1_R1165_U273, P1_R1165_U274, P1_R1165_U275, P1_R1165_U276, P1_R1165_U277, P1_R1165_U278, P1_R1165_U279, P1_R1165_U28, P1_R1165_U280, P1_R1165_U281, P1_R1165_U282, P1_R1165_U283, P1_R1165_U284, P1_R1165_U285, P1_R1165_U286, P1_R1165_U287, P1_R1165_U288, P1_R1165_U289, P1_R1165_U29, P1_R1165_U290, P1_R1165_U291, P1_R1165_U292, P1_R1165_U293, P1_R1165_U294, P1_R1165_U295, P1_R1165_U296, P1_R1165_U297, P1_R1165_U298, P1_R1165_U299, P1_R1165_U30, P1_R1165_U300, P1_R1165_U301, P1_R1165_U302, P1_R1165_U303, P1_R1165_U304, P1_R1165_U305, P1_R1165_U306, P1_R1165_U307, P1_R1165_U308, P1_R1165_U309, P1_R1165_U31, P1_R1165_U310, P1_R1165_U311, P1_R1165_U312, P1_R1165_U313, P1_R1165_U314, P1_R1165_U315, P1_R1165_U316, P1_R1165_U317, P1_R1165_U318, P1_R1165_U319, P1_R1165_U32, P1_R1165_U320, P1_R1165_U321, P1_R1165_U322, P1_R1165_U323, P1_R1165_U324, P1_R1165_U325, P1_R1165_U326, P1_R1165_U327, P1_R1165_U328, P1_R1165_U329, P1_R1165_U33, P1_R1165_U330, P1_R1165_U331, P1_R1165_U332, P1_R1165_U333, P1_R1165_U334, P1_R1165_U335, P1_R1165_U336, P1_R1165_U337, P1_R1165_U338, P1_R1165_U339, P1_R1165_U34, P1_R1165_U340, P1_R1165_U341, P1_R1165_U342, P1_R1165_U343, P1_R1165_U344, P1_R1165_U345, P1_R1165_U346, P1_R1165_U347, P1_R1165_U348, P1_R1165_U349, P1_R1165_U35, P1_R1165_U350, P1_R1165_U351, P1_R1165_U352, P1_R1165_U353, P1_R1165_U354, P1_R1165_U355, P1_R1165_U356, P1_R1165_U357, P1_R1165_U358, P1_R1165_U359, P1_R1165_U36, P1_R1165_U360, P1_R1165_U361, P1_R1165_U362, P1_R1165_U363, P1_R1165_U364, P1_R1165_U365, P1_R1165_U366, P1_R1165_U367, P1_R1165_U368, P1_R1165_U369, P1_R1165_U37, P1_R1165_U370, P1_R1165_U371, P1_R1165_U372, P1_R1165_U373, P1_R1165_U374, P1_R1165_U375, P1_R1165_U376, P1_R1165_U377, P1_R1165_U378, P1_R1165_U379, P1_R1165_U38, P1_R1165_U380, P1_R1165_U381, P1_R1165_U382, P1_R1165_U383, P1_R1165_U384, P1_R1165_U385, P1_R1165_U386, P1_R1165_U387, P1_R1165_U388, P1_R1165_U389, P1_R1165_U39, P1_R1165_U390, P1_R1165_U391, P1_R1165_U392, P1_R1165_U393, P1_R1165_U394, P1_R1165_U395, P1_R1165_U396, P1_R1165_U397, P1_R1165_U398, P1_R1165_U399, P1_R1165_U4, P1_R1165_U40, P1_R1165_U400, P1_R1165_U401, P1_R1165_U402, P1_R1165_U403, P1_R1165_U404, P1_R1165_U405, P1_R1165_U406, P1_R1165_U407, P1_R1165_U408, P1_R1165_U409, P1_R1165_U41, P1_R1165_U410, P1_R1165_U411, P1_R1165_U412, P1_R1165_U413, P1_R1165_U414, P1_R1165_U415, P1_R1165_U416, P1_R1165_U417, P1_R1165_U418, P1_R1165_U419, P1_R1165_U42, P1_R1165_U420, P1_R1165_U421, P1_R1165_U422, P1_R1165_U423, P1_R1165_U424, P1_R1165_U425, P1_R1165_U426, P1_R1165_U427, P1_R1165_U428, P1_R1165_U429, P1_R1165_U43, P1_R1165_U430, P1_R1165_U431, P1_R1165_U432, P1_R1165_U433, P1_R1165_U434, P1_R1165_U435, P1_R1165_U436, P1_R1165_U437, P1_R1165_U438, P1_R1165_U439, P1_R1165_U44, P1_R1165_U440, P1_R1165_U441, P1_R1165_U442, P1_R1165_U443, P1_R1165_U444, P1_R1165_U445, P1_R1165_U446, P1_R1165_U447, P1_R1165_U448, P1_R1165_U449, P1_R1165_U45, P1_R1165_U450, P1_R1165_U451, P1_R1165_U452, P1_R1165_U453, P1_R1165_U454, P1_R1165_U455, P1_R1165_U456, P1_R1165_U457, P1_R1165_U458, P1_R1165_U459, P1_R1165_U46, P1_R1165_U460, P1_R1165_U461, P1_R1165_U462, P1_R1165_U463, P1_R1165_U464, P1_R1165_U465, P1_R1165_U466, P1_R1165_U467, P1_R1165_U468, P1_R1165_U469, P1_R1165_U47, P1_R1165_U470, P1_R1165_U471, P1_R1165_U472, P1_R1165_U473, P1_R1165_U474, P1_R1165_U475, P1_R1165_U476, P1_R1165_U477, P1_R1165_U478, P1_R1165_U479, P1_R1165_U48, P1_R1165_U480, P1_R1165_U481, P1_R1165_U482, P1_R1165_U483, P1_R1165_U484, P1_R1165_U485, P1_R1165_U486, P1_R1165_U487, P1_R1165_U488, P1_R1165_U489, P1_R1165_U49, P1_R1165_U490, P1_R1165_U491, P1_R1165_U492, P1_R1165_U493, P1_R1165_U494, P1_R1165_U495, P1_R1165_U496, P1_R1165_U497, P1_R1165_U498, P1_R1165_U499, P1_R1165_U5, P1_R1165_U50, P1_R1165_U500, P1_R1165_U501, P1_R1165_U502, P1_R1165_U503, P1_R1165_U504, P1_R1165_U505, P1_R1165_U506, P1_R1165_U507, P1_R1165_U508, P1_R1165_U509, P1_R1165_U51, P1_R1165_U510, P1_R1165_U511, P1_R1165_U512, P1_R1165_U513, P1_R1165_U514, P1_R1165_U515, P1_R1165_U516, P1_R1165_U517, P1_R1165_U518, P1_R1165_U519, P1_R1165_U52, P1_R1165_U520, P1_R1165_U521, P1_R1165_U522, P1_R1165_U523, P1_R1165_U524, P1_R1165_U525, P1_R1165_U526, P1_R1165_U527, P1_R1165_U528, P1_R1165_U529, P1_R1165_U53, P1_R1165_U530, P1_R1165_U531, P1_R1165_U532, P1_R1165_U533, P1_R1165_U534, P1_R1165_U535, P1_R1165_U536, P1_R1165_U537, P1_R1165_U538, P1_R1165_U539, P1_R1165_U54, P1_R1165_U540, P1_R1165_U541, P1_R1165_U542, P1_R1165_U543, P1_R1165_U544, P1_R1165_U545, P1_R1165_U546, P1_R1165_U547, P1_R1165_U548, P1_R1165_U549, P1_R1165_U55, P1_R1165_U550, P1_R1165_U551, P1_R1165_U552, P1_R1165_U553, P1_R1165_U554, P1_R1165_U555, P1_R1165_U556, P1_R1165_U557, P1_R1165_U558, P1_R1165_U559, P1_R1165_U56, P1_R1165_U560, P1_R1165_U561, P1_R1165_U562, P1_R1165_U563, P1_R1165_U564, P1_R1165_U565, P1_R1165_U566, P1_R1165_U567, P1_R1165_U568, P1_R1165_U569, P1_R1165_U57, P1_R1165_U570, P1_R1165_U571, P1_R1165_U572, P1_R1165_U573, P1_R1165_U574, P1_R1165_U575, P1_R1165_U576, P1_R1165_U577, P1_R1165_U578, P1_R1165_U579, P1_R1165_U58, P1_R1165_U580, P1_R1165_U581, P1_R1165_U582, P1_R1165_U583, P1_R1165_U584, P1_R1165_U585, P1_R1165_U586, P1_R1165_U587, P1_R1165_U588, P1_R1165_U589, P1_R1165_U59, P1_R1165_U590, P1_R1165_U591, P1_R1165_U592, P1_R1165_U593, P1_R1165_U594, P1_R1165_U595, P1_R1165_U596, P1_R1165_U597, P1_R1165_U598, P1_R1165_U599, P1_R1165_U6, P1_R1165_U60, P1_R1165_U600, P1_R1165_U601, P1_R1165_U602, P1_R1165_U61, P1_R1165_U62, P1_R1165_U63, P1_R1165_U64, P1_R1165_U65, P1_R1165_U66, P1_R1165_U67, P1_R1165_U68, P1_R1165_U69, P1_R1165_U7, P1_R1165_U70, P1_R1165_U71, P1_R1165_U72, P1_R1165_U73, P1_R1165_U74, P1_R1165_U75, P1_R1165_U76, P1_R1165_U77, P1_R1165_U78, P1_R1165_U79, P1_R1165_U8, P1_R1165_U80, P1_R1165_U81, P1_R1165_U82, P1_R1165_U83, P1_R1165_U84, P1_R1165_U85, P1_R1165_U86, P1_R1165_U87, P1_R1165_U88, P1_R1165_U89, P1_R1165_U9, P1_R1165_U90, P1_R1165_U91, P1_R1165_U92, P1_R1165_U93, P1_R1165_U94, P1_R1165_U95, P1_R1165_U96, P1_R1165_U97, P1_R1165_U98, P1_R1165_U99, P1_R1171_U10, P1_R1171_U100, P1_R1171_U101, P1_R1171_U102, P1_R1171_U103, P1_R1171_U104, P1_R1171_U105, P1_R1171_U106, P1_R1171_U107, P1_R1171_U108, P1_R1171_U109, P1_R1171_U11, P1_R1171_U110, P1_R1171_U111, P1_R1171_U112, P1_R1171_U113, P1_R1171_U114, P1_R1171_U115, P1_R1171_U116, P1_R1171_U117, P1_R1171_U118, P1_R1171_U119, P1_R1171_U12, P1_R1171_U120, P1_R1171_U121, P1_R1171_U122, P1_R1171_U123, P1_R1171_U124, P1_R1171_U125, P1_R1171_U126, P1_R1171_U127, P1_R1171_U128, P1_R1171_U129, P1_R1171_U13, P1_R1171_U130, P1_R1171_U131, P1_R1171_U132, P1_R1171_U133, P1_R1171_U134, P1_R1171_U135, P1_R1171_U136, P1_R1171_U137, P1_R1171_U138, P1_R1171_U139, P1_R1171_U14, P1_R1171_U140, P1_R1171_U141, P1_R1171_U142, P1_R1171_U143, P1_R1171_U144, P1_R1171_U145, P1_R1171_U146, P1_R1171_U147, P1_R1171_U148, P1_R1171_U149, P1_R1171_U15, P1_R1171_U150, P1_R1171_U151, P1_R1171_U152, P1_R1171_U153, P1_R1171_U154, P1_R1171_U155, P1_R1171_U156, P1_R1171_U157, P1_R1171_U158, P1_R1171_U159, P1_R1171_U16, P1_R1171_U160, P1_R1171_U161, P1_R1171_U162, P1_R1171_U163, P1_R1171_U164, P1_R1171_U165, P1_R1171_U166, P1_R1171_U167, P1_R1171_U168, P1_R1171_U169, P1_R1171_U17, P1_R1171_U170, P1_R1171_U171, P1_R1171_U172, P1_R1171_U173, P1_R1171_U174, P1_R1171_U175, P1_R1171_U176, P1_R1171_U177, P1_R1171_U178, P1_R1171_U179, P1_R1171_U18, P1_R1171_U180, P1_R1171_U181, P1_R1171_U182, P1_R1171_U183, P1_R1171_U184, P1_R1171_U185, P1_R1171_U186, P1_R1171_U187, P1_R1171_U188, P1_R1171_U189, P1_R1171_U19, P1_R1171_U190, P1_R1171_U191, P1_R1171_U192, P1_R1171_U193, P1_R1171_U194, P1_R1171_U195, P1_R1171_U196, P1_R1171_U197, P1_R1171_U198, P1_R1171_U199, P1_R1171_U20, P1_R1171_U200, P1_R1171_U201, P1_R1171_U202, P1_R1171_U203, P1_R1171_U204, P1_R1171_U205, P1_R1171_U206, P1_R1171_U207, P1_R1171_U208, P1_R1171_U209, P1_R1171_U21, P1_R1171_U210, P1_R1171_U211, P1_R1171_U212, P1_R1171_U213, P1_R1171_U214, P1_R1171_U215, P1_R1171_U216, P1_R1171_U217, P1_R1171_U218, P1_R1171_U219, P1_R1171_U22, P1_R1171_U220, P1_R1171_U221, P1_R1171_U222, P1_R1171_U223, P1_R1171_U224, P1_R1171_U225, P1_R1171_U226, P1_R1171_U227, P1_R1171_U228, P1_R1171_U229, P1_R1171_U23, P1_R1171_U230, P1_R1171_U231, P1_R1171_U232, P1_R1171_U233, P1_R1171_U234, P1_R1171_U235, P1_R1171_U236, P1_R1171_U237, P1_R1171_U238, P1_R1171_U239, P1_R1171_U24, P1_R1171_U240, P1_R1171_U241, P1_R1171_U242, P1_R1171_U243, P1_R1171_U244, P1_R1171_U245, P1_R1171_U246, P1_R1171_U247, P1_R1171_U248, P1_R1171_U249, P1_R1171_U25, P1_R1171_U250, P1_R1171_U251, P1_R1171_U252, P1_R1171_U253, P1_R1171_U254, P1_R1171_U255, P1_R1171_U256, P1_R1171_U257, P1_R1171_U258, P1_R1171_U259, P1_R1171_U26, P1_R1171_U260, P1_R1171_U261, P1_R1171_U262, P1_R1171_U263, P1_R1171_U264, P1_R1171_U265, P1_R1171_U266, P1_R1171_U267, P1_R1171_U268, P1_R1171_U269, P1_R1171_U27, P1_R1171_U270, P1_R1171_U271, P1_R1171_U272, P1_R1171_U273, P1_R1171_U274, P1_R1171_U275, P1_R1171_U276, P1_R1171_U277, P1_R1171_U278, P1_R1171_U279, P1_R1171_U28, P1_R1171_U280, P1_R1171_U281, P1_R1171_U282, P1_R1171_U283, P1_R1171_U284, P1_R1171_U285, P1_R1171_U286, P1_R1171_U287, P1_R1171_U288, P1_R1171_U289, P1_R1171_U29, P1_R1171_U290, P1_R1171_U291, P1_R1171_U292, P1_R1171_U293, P1_R1171_U294, P1_R1171_U295, P1_R1171_U296, P1_R1171_U297, P1_R1171_U298, P1_R1171_U299, P1_R1171_U30, P1_R1171_U300, P1_R1171_U301, P1_R1171_U302, P1_R1171_U303, P1_R1171_U304, P1_R1171_U305, P1_R1171_U306, P1_R1171_U307, P1_R1171_U308, P1_R1171_U309, P1_R1171_U31, P1_R1171_U310, P1_R1171_U311, P1_R1171_U312, P1_R1171_U313, P1_R1171_U314, P1_R1171_U315, P1_R1171_U316, P1_R1171_U317, P1_R1171_U318, P1_R1171_U319, P1_R1171_U32, P1_R1171_U320, P1_R1171_U321, P1_R1171_U322, P1_R1171_U323, P1_R1171_U324, P1_R1171_U325, P1_R1171_U326, P1_R1171_U327, P1_R1171_U328, P1_R1171_U329, P1_R1171_U33, P1_R1171_U330, P1_R1171_U331, P1_R1171_U332, P1_R1171_U333, P1_R1171_U334, P1_R1171_U335, P1_R1171_U336, P1_R1171_U337, P1_R1171_U338, P1_R1171_U339, P1_R1171_U34, P1_R1171_U340, P1_R1171_U341, P1_R1171_U342, P1_R1171_U343, P1_R1171_U344, P1_R1171_U345, P1_R1171_U346, P1_R1171_U347, P1_R1171_U348, P1_R1171_U349, P1_R1171_U35, P1_R1171_U350, P1_R1171_U351, P1_R1171_U352, P1_R1171_U353, P1_R1171_U354, P1_R1171_U355, P1_R1171_U356, P1_R1171_U357, P1_R1171_U358, P1_R1171_U359, P1_R1171_U36, P1_R1171_U360, P1_R1171_U361, P1_R1171_U362, P1_R1171_U363, P1_R1171_U364, P1_R1171_U365, P1_R1171_U366, P1_R1171_U367, P1_R1171_U368, P1_R1171_U369, P1_R1171_U37, P1_R1171_U370, P1_R1171_U371, P1_R1171_U372, P1_R1171_U373, P1_R1171_U374, P1_R1171_U375, P1_R1171_U376, P1_R1171_U377, P1_R1171_U378, P1_R1171_U379, P1_R1171_U38, P1_R1171_U380, P1_R1171_U381, P1_R1171_U382, P1_R1171_U383, P1_R1171_U384, P1_R1171_U385, P1_R1171_U386, P1_R1171_U387, P1_R1171_U388, P1_R1171_U389, P1_R1171_U39, P1_R1171_U390, P1_R1171_U391, P1_R1171_U392, P1_R1171_U393, P1_R1171_U394, P1_R1171_U395, P1_R1171_U396, P1_R1171_U397, P1_R1171_U398, P1_R1171_U399, P1_R1171_U4, P1_R1171_U40, P1_R1171_U400, P1_R1171_U401, P1_R1171_U402, P1_R1171_U403, P1_R1171_U404, P1_R1171_U405, P1_R1171_U406, P1_R1171_U407, P1_R1171_U408, P1_R1171_U409, P1_R1171_U41, P1_R1171_U410, P1_R1171_U411, P1_R1171_U412, P1_R1171_U413, P1_R1171_U414, P1_R1171_U415, P1_R1171_U416, P1_R1171_U417, P1_R1171_U418, P1_R1171_U419, P1_R1171_U42, P1_R1171_U420, P1_R1171_U421, P1_R1171_U422, P1_R1171_U423, P1_R1171_U424, P1_R1171_U425, P1_R1171_U426, P1_R1171_U427, P1_R1171_U428, P1_R1171_U429, P1_R1171_U43, P1_R1171_U430, P1_R1171_U431, P1_R1171_U432, P1_R1171_U433, P1_R1171_U434, P1_R1171_U435, P1_R1171_U436, P1_R1171_U437, P1_R1171_U438, P1_R1171_U439, P1_R1171_U44, P1_R1171_U440, P1_R1171_U441, P1_R1171_U442, P1_R1171_U443, P1_R1171_U444, P1_R1171_U445, P1_R1171_U446, P1_R1171_U447, P1_R1171_U448, P1_R1171_U449, P1_R1171_U45, P1_R1171_U450, P1_R1171_U451, P1_R1171_U452, P1_R1171_U453, P1_R1171_U454, P1_R1171_U455, P1_R1171_U456, P1_R1171_U457, P1_R1171_U458, P1_R1171_U459, P1_R1171_U46, P1_R1171_U460, P1_R1171_U461, P1_R1171_U462, P1_R1171_U463, P1_R1171_U464, P1_R1171_U465, P1_R1171_U466, P1_R1171_U467, P1_R1171_U468, P1_R1171_U469, P1_R1171_U47, P1_R1171_U470, P1_R1171_U471, P1_R1171_U472, P1_R1171_U473, P1_R1171_U474, P1_R1171_U475, P1_R1171_U476, P1_R1171_U477, P1_R1171_U478, P1_R1171_U479, P1_R1171_U48, P1_R1171_U480, P1_R1171_U481, P1_R1171_U482, P1_R1171_U483, P1_R1171_U484, P1_R1171_U485, P1_R1171_U486, P1_R1171_U487, P1_R1171_U488, P1_R1171_U489, P1_R1171_U49, P1_R1171_U490, P1_R1171_U491, P1_R1171_U492, P1_R1171_U493, P1_R1171_U494, P1_R1171_U495, P1_R1171_U496, P1_R1171_U497, P1_R1171_U498, P1_R1171_U499, P1_R1171_U5, P1_R1171_U50, P1_R1171_U500, P1_R1171_U501, P1_R1171_U502, P1_R1171_U503, P1_R1171_U51, P1_R1171_U52, P1_R1171_U53, P1_R1171_U54, P1_R1171_U55, P1_R1171_U56, P1_R1171_U57, P1_R1171_U58, P1_R1171_U59, P1_R1171_U6, P1_R1171_U60, P1_R1171_U61, P1_R1171_U62, P1_R1171_U63, P1_R1171_U64, P1_R1171_U65, P1_R1171_U66, P1_R1171_U67, P1_R1171_U68, P1_R1171_U69, P1_R1171_U7, P1_R1171_U70, P1_R1171_U71, P1_R1171_U72, P1_R1171_U73, P1_R1171_U74, P1_R1171_U75, P1_R1171_U76, P1_R1171_U77, P1_R1171_U78, P1_R1171_U79, P1_R1171_U8, P1_R1171_U80, P1_R1171_U81, P1_R1171_U82, P1_R1171_U83, P1_R1171_U84, P1_R1171_U85, P1_R1171_U86, P1_R1171_U87, P1_R1171_U88, P1_R1171_U89, P1_R1171_U9, P1_R1171_U90, P1_R1171_U91, P1_R1171_U92, P1_R1171_U93, P1_R1171_U94, P1_R1171_U95, P1_R1171_U96, P1_R1171_U97, P1_R1171_U98, P1_R1171_U99, P1_R1192_U10, P1_R1192_U100, P1_R1192_U101, P1_R1192_U102, P1_R1192_U103, P1_R1192_U104, P1_R1192_U105, P1_R1192_U106, P1_R1192_U107, P1_R1192_U108, P1_R1192_U109, P1_R1192_U11, P1_R1192_U110, P1_R1192_U111, P1_R1192_U112, P1_R1192_U113, P1_R1192_U114, P1_R1192_U115, P1_R1192_U116, P1_R1192_U117, P1_R1192_U118, P1_R1192_U119, P1_R1192_U12, P1_R1192_U120, P1_R1192_U121, P1_R1192_U122, P1_R1192_U123, P1_R1192_U124, P1_R1192_U125, P1_R1192_U126, P1_R1192_U127, P1_R1192_U128, P1_R1192_U129, P1_R1192_U13, P1_R1192_U130, P1_R1192_U131, P1_R1192_U132, P1_R1192_U133, P1_R1192_U134, P1_R1192_U135, P1_R1192_U136, P1_R1192_U137, P1_R1192_U138, P1_R1192_U139, P1_R1192_U14, P1_R1192_U140, P1_R1192_U141, P1_R1192_U142, P1_R1192_U143, P1_R1192_U144, P1_R1192_U145, P1_R1192_U146, P1_R1192_U147, P1_R1192_U148, P1_R1192_U149, P1_R1192_U15, P1_R1192_U150, P1_R1192_U151, P1_R1192_U152, P1_R1192_U153, P1_R1192_U154, P1_R1192_U155, P1_R1192_U156, P1_R1192_U157, P1_R1192_U158, P1_R1192_U159, P1_R1192_U16, P1_R1192_U160, P1_R1192_U161, P1_R1192_U162, P1_R1192_U163, P1_R1192_U164, P1_R1192_U165, P1_R1192_U166, P1_R1192_U167, P1_R1192_U168, P1_R1192_U169, P1_R1192_U17, P1_R1192_U170, P1_R1192_U171, P1_R1192_U172, P1_R1192_U173, P1_R1192_U174, P1_R1192_U175, P1_R1192_U176, P1_R1192_U177, P1_R1192_U178, P1_R1192_U179, P1_R1192_U18, P1_R1192_U180, P1_R1192_U181, P1_R1192_U182, P1_R1192_U183, P1_R1192_U184, P1_R1192_U185, P1_R1192_U186, P1_R1192_U187, P1_R1192_U188, P1_R1192_U189, P1_R1192_U19, P1_R1192_U190, P1_R1192_U191, P1_R1192_U192, P1_R1192_U193, P1_R1192_U194, P1_R1192_U195, P1_R1192_U196, P1_R1192_U197, P1_R1192_U198, P1_R1192_U199, P1_R1192_U20, P1_R1192_U200, P1_R1192_U201, P1_R1192_U202, P1_R1192_U203, P1_R1192_U204, P1_R1192_U205, P1_R1192_U206, P1_R1192_U207, P1_R1192_U208, P1_R1192_U209, P1_R1192_U21, P1_R1192_U210, P1_R1192_U211, P1_R1192_U212, P1_R1192_U213, P1_R1192_U214, P1_R1192_U215, P1_R1192_U216, P1_R1192_U217, P1_R1192_U218, P1_R1192_U219, P1_R1192_U22, P1_R1192_U220, P1_R1192_U221, P1_R1192_U222, P1_R1192_U223, P1_R1192_U224, P1_R1192_U225, P1_R1192_U226, P1_R1192_U227, P1_R1192_U228, P1_R1192_U229, P1_R1192_U23, P1_R1192_U230, P1_R1192_U231, P1_R1192_U232, P1_R1192_U233, P1_R1192_U234, P1_R1192_U235, P1_R1192_U236, P1_R1192_U237, P1_R1192_U238, P1_R1192_U239, P1_R1192_U24, P1_R1192_U240, P1_R1192_U241, P1_R1192_U242, P1_R1192_U243, P1_R1192_U244, P1_R1192_U245, P1_R1192_U246, P1_R1192_U247, P1_R1192_U248, P1_R1192_U249, P1_R1192_U25, P1_R1192_U250, P1_R1192_U251, P1_R1192_U252, P1_R1192_U253, P1_R1192_U254, P1_R1192_U255, P1_R1192_U256, P1_R1192_U257, P1_R1192_U258, P1_R1192_U259, P1_R1192_U26, P1_R1192_U260, P1_R1192_U261, P1_R1192_U262, P1_R1192_U263, P1_R1192_U264, P1_R1192_U265, P1_R1192_U266, P1_R1192_U267, P1_R1192_U268, P1_R1192_U269, P1_R1192_U27, P1_R1192_U270, P1_R1192_U271, P1_R1192_U272, P1_R1192_U273, P1_R1192_U274, P1_R1192_U275, P1_R1192_U276, P1_R1192_U277, P1_R1192_U278, P1_R1192_U279, P1_R1192_U28, P1_R1192_U280, P1_R1192_U281, P1_R1192_U282, P1_R1192_U283, P1_R1192_U284, P1_R1192_U285, P1_R1192_U286, P1_R1192_U287, P1_R1192_U288, P1_R1192_U289, P1_R1192_U29, P1_R1192_U290, P1_R1192_U291, P1_R1192_U292, P1_R1192_U293, P1_R1192_U294, P1_R1192_U295, P1_R1192_U296, P1_R1192_U297, P1_R1192_U298, P1_R1192_U299, P1_R1192_U30, P1_R1192_U300, P1_R1192_U301, P1_R1192_U302, P1_R1192_U303, P1_R1192_U304, P1_R1192_U305, P1_R1192_U306, P1_R1192_U307, P1_R1192_U308, P1_R1192_U309, P1_R1192_U31, P1_R1192_U310, P1_R1192_U311, P1_R1192_U312, P1_R1192_U313, P1_R1192_U314, P1_R1192_U315, P1_R1192_U316, P1_R1192_U317, P1_R1192_U318, P1_R1192_U319, P1_R1192_U32, P1_R1192_U320, P1_R1192_U321, P1_R1192_U322, P1_R1192_U323, P1_R1192_U324, P1_R1192_U325, P1_R1192_U326, P1_R1192_U327, P1_R1192_U328, P1_R1192_U329, P1_R1192_U33, P1_R1192_U330, P1_R1192_U331, P1_R1192_U332, P1_R1192_U333, P1_R1192_U334, P1_R1192_U335, P1_R1192_U336, P1_R1192_U337, P1_R1192_U338, P1_R1192_U339, P1_R1192_U34, P1_R1192_U340, P1_R1192_U341, P1_R1192_U342, P1_R1192_U343, P1_R1192_U344, P1_R1192_U345, P1_R1192_U346, P1_R1192_U347, P1_R1192_U348, P1_R1192_U349, P1_R1192_U35, P1_R1192_U350, P1_R1192_U351, P1_R1192_U352, P1_R1192_U353, P1_R1192_U354, P1_R1192_U355, P1_R1192_U356, P1_R1192_U357, P1_R1192_U358, P1_R1192_U359, P1_R1192_U36, P1_R1192_U360, P1_R1192_U361, P1_R1192_U362, P1_R1192_U363, P1_R1192_U364, P1_R1192_U365, P1_R1192_U366, P1_R1192_U367, P1_R1192_U368, P1_R1192_U369, P1_R1192_U37, P1_R1192_U370, P1_R1192_U371, P1_R1192_U372, P1_R1192_U373, P1_R1192_U374, P1_R1192_U375, P1_R1192_U376, P1_R1192_U377, P1_R1192_U378, P1_R1192_U379, P1_R1192_U38, P1_R1192_U380, P1_R1192_U381, P1_R1192_U382, P1_R1192_U383, P1_R1192_U384, P1_R1192_U385, P1_R1192_U386, P1_R1192_U387, P1_R1192_U388, P1_R1192_U389, P1_R1192_U39, P1_R1192_U390, P1_R1192_U391, P1_R1192_U392, P1_R1192_U393, P1_R1192_U394, P1_R1192_U395, P1_R1192_U396, P1_R1192_U397, P1_R1192_U398, P1_R1192_U399, P1_R1192_U40, P1_R1192_U400, P1_R1192_U401, P1_R1192_U402, P1_R1192_U403, P1_R1192_U404, P1_R1192_U405, P1_R1192_U406, P1_R1192_U407, P1_R1192_U408, P1_R1192_U409, P1_R1192_U41, P1_R1192_U410, P1_R1192_U411, P1_R1192_U412, P1_R1192_U413, P1_R1192_U414, P1_R1192_U415, P1_R1192_U416, P1_R1192_U417, P1_R1192_U418, P1_R1192_U419, P1_R1192_U42, P1_R1192_U420, P1_R1192_U421, P1_R1192_U422, P1_R1192_U423, P1_R1192_U424, P1_R1192_U425, P1_R1192_U426, P1_R1192_U427, P1_R1192_U428, P1_R1192_U429, P1_R1192_U43, P1_R1192_U430, P1_R1192_U431, P1_R1192_U432, P1_R1192_U433, P1_R1192_U434, P1_R1192_U435, P1_R1192_U436, P1_R1192_U437, P1_R1192_U438, P1_R1192_U439, P1_R1192_U44, P1_R1192_U440, P1_R1192_U441, P1_R1192_U442, P1_R1192_U443, P1_R1192_U444, P1_R1192_U445, P1_R1192_U446, P1_R1192_U447, P1_R1192_U448, P1_R1192_U449, P1_R1192_U45, P1_R1192_U450, P1_R1192_U451, P1_R1192_U452, P1_R1192_U453, P1_R1192_U454, P1_R1192_U455, P1_R1192_U456, P1_R1192_U457, P1_R1192_U458, P1_R1192_U459, P1_R1192_U46, P1_R1192_U460, P1_R1192_U461, P1_R1192_U462, P1_R1192_U463, P1_R1192_U464, P1_R1192_U465, P1_R1192_U466, P1_R1192_U467, P1_R1192_U468, P1_R1192_U469, P1_R1192_U47, P1_R1192_U470, P1_R1192_U471, P1_R1192_U472, P1_R1192_U473, P1_R1192_U48, P1_R1192_U49, P1_R1192_U50, P1_R1192_U51, P1_R1192_U52, P1_R1192_U53, P1_R1192_U54, P1_R1192_U55, P1_R1192_U56, P1_R1192_U57, P1_R1192_U58, P1_R1192_U59, P1_R1192_U6, P1_R1192_U60, P1_R1192_U61, P1_R1192_U62, P1_R1192_U63, P1_R1192_U64, P1_R1192_U65, P1_R1192_U66, P1_R1192_U67, P1_R1192_U68, P1_R1192_U69, P1_R1192_U7, P1_R1192_U70, P1_R1192_U71, P1_R1192_U72, P1_R1192_U73, P1_R1192_U74, P1_R1192_U75, P1_R1192_U76, P1_R1192_U77, P1_R1192_U78, P1_R1192_U79, P1_R1192_U8, P1_R1192_U80, P1_R1192_U81, P1_R1192_U82, P1_R1192_U83, P1_R1192_U84, P1_R1192_U85, P1_R1192_U86, P1_R1192_U87, P1_R1192_U88, P1_R1192_U89, P1_R1192_U9, P1_R1192_U90, P1_R1192_U91, P1_R1192_U92, P1_R1192_U93, P1_R1192_U94, P1_R1192_U95, P1_R1192_U96, P1_R1192_U97, P1_R1192_U98, P1_R1192_U99, P1_R1207_U10, P1_R1207_U100, P1_R1207_U101, P1_R1207_U102, P1_R1207_U103, P1_R1207_U104, P1_R1207_U105, P1_R1207_U106, P1_R1207_U107, P1_R1207_U108, P1_R1207_U109, P1_R1207_U11, P1_R1207_U110, P1_R1207_U111, P1_R1207_U112, P1_R1207_U113, P1_R1207_U114, P1_R1207_U115, P1_R1207_U116, P1_R1207_U117, P1_R1207_U118, P1_R1207_U119, P1_R1207_U12, P1_R1207_U120, P1_R1207_U121, P1_R1207_U122, P1_R1207_U123, P1_R1207_U124, P1_R1207_U125, P1_R1207_U126, P1_R1207_U127, P1_R1207_U128, P1_R1207_U129, P1_R1207_U13, P1_R1207_U130, P1_R1207_U131, P1_R1207_U132, P1_R1207_U133, P1_R1207_U134, P1_R1207_U135, P1_R1207_U136, P1_R1207_U137, P1_R1207_U138, P1_R1207_U139, P1_R1207_U14, P1_R1207_U140, P1_R1207_U141, P1_R1207_U142, P1_R1207_U143, P1_R1207_U144, P1_R1207_U145, P1_R1207_U146, P1_R1207_U147, P1_R1207_U148, P1_R1207_U149, P1_R1207_U15, P1_R1207_U150, P1_R1207_U151, P1_R1207_U152, P1_R1207_U153, P1_R1207_U154, P1_R1207_U155, P1_R1207_U156, P1_R1207_U157, P1_R1207_U158, P1_R1207_U159, P1_R1207_U16, P1_R1207_U160, P1_R1207_U161, P1_R1207_U162, P1_R1207_U163, P1_R1207_U164, P1_R1207_U165, P1_R1207_U166, P1_R1207_U167, P1_R1207_U168, P1_R1207_U169, P1_R1207_U17, P1_R1207_U170, P1_R1207_U171, P1_R1207_U172, P1_R1207_U173, P1_R1207_U174, P1_R1207_U175, P1_R1207_U176, P1_R1207_U177, P1_R1207_U178, P1_R1207_U179, P1_R1207_U18, P1_R1207_U180, P1_R1207_U181, P1_R1207_U182, P1_R1207_U183, P1_R1207_U184, P1_R1207_U185, P1_R1207_U186, P1_R1207_U187, P1_R1207_U188, P1_R1207_U189, P1_R1207_U19, P1_R1207_U190, P1_R1207_U191, P1_R1207_U192, P1_R1207_U193, P1_R1207_U194, P1_R1207_U195, P1_R1207_U196, P1_R1207_U197, P1_R1207_U198, P1_R1207_U199, P1_R1207_U20, P1_R1207_U200, P1_R1207_U201, P1_R1207_U202, P1_R1207_U203, P1_R1207_U204, P1_R1207_U205, P1_R1207_U206, P1_R1207_U207, P1_R1207_U208, P1_R1207_U209, P1_R1207_U21, P1_R1207_U210, P1_R1207_U211, P1_R1207_U212, P1_R1207_U213, P1_R1207_U214, P1_R1207_U215, P1_R1207_U216, P1_R1207_U217, P1_R1207_U218, P1_R1207_U219, P1_R1207_U22, P1_R1207_U220, P1_R1207_U221, P1_R1207_U222, P1_R1207_U223, P1_R1207_U224, P1_R1207_U225, P1_R1207_U226, P1_R1207_U227, P1_R1207_U228, P1_R1207_U229, P1_R1207_U23, P1_R1207_U230, P1_R1207_U231, P1_R1207_U232, P1_R1207_U233, P1_R1207_U234, P1_R1207_U235, P1_R1207_U236, P1_R1207_U237, P1_R1207_U238, P1_R1207_U239, P1_R1207_U24, P1_R1207_U240, P1_R1207_U241, P1_R1207_U242, P1_R1207_U243, P1_R1207_U244, P1_R1207_U245, P1_R1207_U246, P1_R1207_U247, P1_R1207_U248, P1_R1207_U249, P1_R1207_U25, P1_R1207_U250, P1_R1207_U251, P1_R1207_U252, P1_R1207_U253, P1_R1207_U254, P1_R1207_U255, P1_R1207_U256, P1_R1207_U257, P1_R1207_U258, P1_R1207_U259, P1_R1207_U26, P1_R1207_U260, P1_R1207_U261, P1_R1207_U262, P1_R1207_U263, P1_R1207_U264, P1_R1207_U265, P1_R1207_U266, P1_R1207_U267, P1_R1207_U268, P1_R1207_U269, P1_R1207_U27, P1_R1207_U270, P1_R1207_U271, P1_R1207_U272, P1_R1207_U273, P1_R1207_U274, P1_R1207_U275, P1_R1207_U276, P1_R1207_U277, P1_R1207_U278, P1_R1207_U279, P1_R1207_U28, P1_R1207_U280, P1_R1207_U281, P1_R1207_U282, P1_R1207_U283, P1_R1207_U284, P1_R1207_U285, P1_R1207_U286, P1_R1207_U287, P1_R1207_U288, P1_R1207_U289, P1_R1207_U29, P1_R1207_U290, P1_R1207_U291, P1_R1207_U292, P1_R1207_U293, P1_R1207_U294, P1_R1207_U295, P1_R1207_U296, P1_R1207_U297, P1_R1207_U298, P1_R1207_U299, P1_R1207_U30, P1_R1207_U300, P1_R1207_U301, P1_R1207_U302, P1_R1207_U303, P1_R1207_U304, P1_R1207_U305, P1_R1207_U306, P1_R1207_U307, P1_R1207_U308, P1_R1207_U309, P1_R1207_U31, P1_R1207_U310, P1_R1207_U311, P1_R1207_U312, P1_R1207_U313, P1_R1207_U314, P1_R1207_U315, P1_R1207_U316, P1_R1207_U317, P1_R1207_U318, P1_R1207_U319, P1_R1207_U32, P1_R1207_U320, P1_R1207_U321, P1_R1207_U322, P1_R1207_U323, P1_R1207_U324, P1_R1207_U325, P1_R1207_U326, P1_R1207_U327, P1_R1207_U328, P1_R1207_U329, P1_R1207_U33, P1_R1207_U330, P1_R1207_U331, P1_R1207_U332, P1_R1207_U333, P1_R1207_U334, P1_R1207_U335, P1_R1207_U336, P1_R1207_U337, P1_R1207_U338, P1_R1207_U339, P1_R1207_U34, P1_R1207_U340, P1_R1207_U341, P1_R1207_U342, P1_R1207_U343, P1_R1207_U344, P1_R1207_U345, P1_R1207_U346, P1_R1207_U347, P1_R1207_U348, P1_R1207_U349, P1_R1207_U35, P1_R1207_U350, P1_R1207_U351, P1_R1207_U352, P1_R1207_U353, P1_R1207_U354, P1_R1207_U355, P1_R1207_U356, P1_R1207_U357, P1_R1207_U358, P1_R1207_U359, P1_R1207_U36, P1_R1207_U360, P1_R1207_U361, P1_R1207_U362, P1_R1207_U363, P1_R1207_U364, P1_R1207_U365, P1_R1207_U366, P1_R1207_U367, P1_R1207_U368, P1_R1207_U369, P1_R1207_U37, P1_R1207_U370, P1_R1207_U371, P1_R1207_U372, P1_R1207_U373, P1_R1207_U374, P1_R1207_U375, P1_R1207_U376, P1_R1207_U377, P1_R1207_U378, P1_R1207_U379, P1_R1207_U38, P1_R1207_U380, P1_R1207_U381, P1_R1207_U382, P1_R1207_U383, P1_R1207_U384, P1_R1207_U385, P1_R1207_U386, P1_R1207_U387, P1_R1207_U388, P1_R1207_U389, P1_R1207_U39, P1_R1207_U390, P1_R1207_U391, P1_R1207_U392, P1_R1207_U393, P1_R1207_U394, P1_R1207_U395, P1_R1207_U396, P1_R1207_U397, P1_R1207_U398, P1_R1207_U399, P1_R1207_U40, P1_R1207_U400, P1_R1207_U401, P1_R1207_U402, P1_R1207_U403, P1_R1207_U404, P1_R1207_U405, P1_R1207_U406, P1_R1207_U407, P1_R1207_U408, P1_R1207_U409, P1_R1207_U41, P1_R1207_U410, P1_R1207_U411, P1_R1207_U412, P1_R1207_U413, P1_R1207_U414, P1_R1207_U415, P1_R1207_U416, P1_R1207_U417, P1_R1207_U418, P1_R1207_U419, P1_R1207_U42, P1_R1207_U420, P1_R1207_U421, P1_R1207_U422, P1_R1207_U423, P1_R1207_U424, P1_R1207_U425, P1_R1207_U426, P1_R1207_U427, P1_R1207_U428, P1_R1207_U429, P1_R1207_U43, P1_R1207_U430, P1_R1207_U431, P1_R1207_U432, P1_R1207_U433, P1_R1207_U434, P1_R1207_U435, P1_R1207_U436, P1_R1207_U437, P1_R1207_U438, P1_R1207_U439, P1_R1207_U44, P1_R1207_U440, P1_R1207_U441, P1_R1207_U442, P1_R1207_U443, P1_R1207_U444, P1_R1207_U445, P1_R1207_U446, P1_R1207_U447, P1_R1207_U448, P1_R1207_U449, P1_R1207_U45, P1_R1207_U450, P1_R1207_U451, P1_R1207_U452, P1_R1207_U453, P1_R1207_U454, P1_R1207_U455, P1_R1207_U456, P1_R1207_U457, P1_R1207_U458, P1_R1207_U459, P1_R1207_U46, P1_R1207_U460, P1_R1207_U461, P1_R1207_U462, P1_R1207_U463, P1_R1207_U464, P1_R1207_U465, P1_R1207_U466, P1_R1207_U467, P1_R1207_U468, P1_R1207_U469, P1_R1207_U47, P1_R1207_U470, P1_R1207_U471, P1_R1207_U472, P1_R1207_U473, P1_R1207_U48, P1_R1207_U49, P1_R1207_U50, P1_R1207_U51, P1_R1207_U52, P1_R1207_U53, P1_R1207_U54, P1_R1207_U55, P1_R1207_U56, P1_R1207_U57, P1_R1207_U58, P1_R1207_U59, P1_R1207_U6, P1_R1207_U60, P1_R1207_U61, P1_R1207_U62, P1_R1207_U63, P1_R1207_U64, P1_R1207_U65, P1_R1207_U66, P1_R1207_U67, P1_R1207_U68, P1_R1207_U69, P1_R1207_U7, P1_R1207_U70, P1_R1207_U71, P1_R1207_U72, P1_R1207_U73, P1_R1207_U74, P1_R1207_U75, P1_R1207_U76, P1_R1207_U77, P1_R1207_U78, P1_R1207_U79, P1_R1207_U8, P1_R1207_U80, P1_R1207_U81, P1_R1207_U82, P1_R1207_U83, P1_R1207_U84, P1_R1207_U85, P1_R1207_U86, P1_R1207_U87, P1_R1207_U88, P1_R1207_U89, P1_R1207_U9, P1_R1207_U90, P1_R1207_U91, P1_R1207_U92, P1_R1207_U93, P1_R1207_U94, P1_R1207_U95, P1_R1207_U96, P1_R1207_U97, P1_R1207_U98, P1_R1207_U99, P1_R1222_U10, P1_R1222_U100, P1_R1222_U101, P1_R1222_U102, P1_R1222_U103, P1_R1222_U104, P1_R1222_U105, P1_R1222_U106, P1_R1222_U107, P1_R1222_U108, P1_R1222_U109, P1_R1222_U11, P1_R1222_U110, P1_R1222_U111, P1_R1222_U112, P1_R1222_U113, P1_R1222_U114, P1_R1222_U115, P1_R1222_U116, P1_R1222_U117, P1_R1222_U118, P1_R1222_U119, P1_R1222_U12, P1_R1222_U120, P1_R1222_U121, P1_R1222_U122, P1_R1222_U123, P1_R1222_U124, P1_R1222_U125, P1_R1222_U126, P1_R1222_U127, P1_R1222_U128, P1_R1222_U129, P1_R1222_U13, P1_R1222_U130, P1_R1222_U131, P1_R1222_U132, P1_R1222_U133, P1_R1222_U134, P1_R1222_U135, P1_R1222_U136, P1_R1222_U137, P1_R1222_U138, P1_R1222_U139, P1_R1222_U14, P1_R1222_U140, P1_R1222_U141, P1_R1222_U142, P1_R1222_U143, P1_R1222_U144, P1_R1222_U145, P1_R1222_U146, P1_R1222_U147, P1_R1222_U148, P1_R1222_U149, P1_R1222_U15, P1_R1222_U150, P1_R1222_U151, P1_R1222_U152, P1_R1222_U153, P1_R1222_U154, P1_R1222_U155, P1_R1222_U156, P1_R1222_U157, P1_R1222_U158, P1_R1222_U159, P1_R1222_U16, P1_R1222_U160, P1_R1222_U161, P1_R1222_U162, P1_R1222_U163, P1_R1222_U164, P1_R1222_U165, P1_R1222_U166, P1_R1222_U167, P1_R1222_U168, P1_R1222_U169, P1_R1222_U17, P1_R1222_U170, P1_R1222_U171, P1_R1222_U172, P1_R1222_U173, P1_R1222_U174, P1_R1222_U175, P1_R1222_U176, P1_R1222_U177, P1_R1222_U178, P1_R1222_U179, P1_R1222_U18, P1_R1222_U180, P1_R1222_U181, P1_R1222_U182, P1_R1222_U183, P1_R1222_U184, P1_R1222_U185, P1_R1222_U186, P1_R1222_U187, P1_R1222_U188, P1_R1222_U189, P1_R1222_U19, P1_R1222_U190, P1_R1222_U191, P1_R1222_U192, P1_R1222_U193, P1_R1222_U194, P1_R1222_U195, P1_R1222_U196, P1_R1222_U197, P1_R1222_U198, P1_R1222_U199, P1_R1222_U20, P1_R1222_U200, P1_R1222_U201, P1_R1222_U202, P1_R1222_U203, P1_R1222_U204, P1_R1222_U205, P1_R1222_U206, P1_R1222_U207, P1_R1222_U208, P1_R1222_U209, P1_R1222_U21, P1_R1222_U210, P1_R1222_U211, P1_R1222_U212, P1_R1222_U213, P1_R1222_U214, P1_R1222_U215, P1_R1222_U216, P1_R1222_U217, P1_R1222_U218, P1_R1222_U219, P1_R1222_U22, P1_R1222_U220, P1_R1222_U221, P1_R1222_U222, P1_R1222_U223, P1_R1222_U224, P1_R1222_U225, P1_R1222_U226, P1_R1222_U227, P1_R1222_U228, P1_R1222_U229, P1_R1222_U23, P1_R1222_U230, P1_R1222_U231, P1_R1222_U232, P1_R1222_U233, P1_R1222_U234, P1_R1222_U235, P1_R1222_U236, P1_R1222_U237, P1_R1222_U238, P1_R1222_U239, P1_R1222_U24, P1_R1222_U240, P1_R1222_U241, P1_R1222_U242, P1_R1222_U243, P1_R1222_U244, P1_R1222_U245, P1_R1222_U246, P1_R1222_U247, P1_R1222_U248, P1_R1222_U249, P1_R1222_U25, P1_R1222_U250, P1_R1222_U251, P1_R1222_U252, P1_R1222_U253, P1_R1222_U254, P1_R1222_U255, P1_R1222_U256, P1_R1222_U257, P1_R1222_U258, P1_R1222_U259, P1_R1222_U26, P1_R1222_U260, P1_R1222_U261, P1_R1222_U262, P1_R1222_U263, P1_R1222_U264, P1_R1222_U265, P1_R1222_U266, P1_R1222_U267, P1_R1222_U268, P1_R1222_U269, P1_R1222_U27, P1_R1222_U270, P1_R1222_U271, P1_R1222_U272, P1_R1222_U273, P1_R1222_U274, P1_R1222_U275, P1_R1222_U276, P1_R1222_U277, P1_R1222_U278, P1_R1222_U279, P1_R1222_U28, P1_R1222_U280, P1_R1222_U281, P1_R1222_U282, P1_R1222_U283, P1_R1222_U284, P1_R1222_U285, P1_R1222_U286, P1_R1222_U287, P1_R1222_U288, P1_R1222_U289, P1_R1222_U29, P1_R1222_U290, P1_R1222_U291, P1_R1222_U292, P1_R1222_U293, P1_R1222_U294, P1_R1222_U295, P1_R1222_U296, P1_R1222_U297, P1_R1222_U298, P1_R1222_U299, P1_R1222_U30, P1_R1222_U300, P1_R1222_U301, P1_R1222_U302, P1_R1222_U303, P1_R1222_U304, P1_R1222_U305, P1_R1222_U306, P1_R1222_U307, P1_R1222_U308, P1_R1222_U309, P1_R1222_U31, P1_R1222_U310, P1_R1222_U311, P1_R1222_U312, P1_R1222_U313, P1_R1222_U314, P1_R1222_U315, P1_R1222_U316, P1_R1222_U317, P1_R1222_U318, P1_R1222_U319, P1_R1222_U32, P1_R1222_U320, P1_R1222_U321, P1_R1222_U322, P1_R1222_U323, P1_R1222_U324, P1_R1222_U325, P1_R1222_U326, P1_R1222_U327, P1_R1222_U328, P1_R1222_U329, P1_R1222_U33, P1_R1222_U330, P1_R1222_U331, P1_R1222_U332, P1_R1222_U333, P1_R1222_U334, P1_R1222_U335, P1_R1222_U336, P1_R1222_U337, P1_R1222_U338, P1_R1222_U339, P1_R1222_U34, P1_R1222_U340, P1_R1222_U341, P1_R1222_U342, P1_R1222_U343, P1_R1222_U344, P1_R1222_U345, P1_R1222_U346, P1_R1222_U347, P1_R1222_U348, P1_R1222_U349, P1_R1222_U35, P1_R1222_U350, P1_R1222_U351, P1_R1222_U352, P1_R1222_U353, P1_R1222_U354, P1_R1222_U355, P1_R1222_U356, P1_R1222_U357, P1_R1222_U358, P1_R1222_U359, P1_R1222_U36, P1_R1222_U360, P1_R1222_U361, P1_R1222_U362, P1_R1222_U363, P1_R1222_U364, P1_R1222_U365, P1_R1222_U366, P1_R1222_U367, P1_R1222_U368, P1_R1222_U369, P1_R1222_U37, P1_R1222_U370, P1_R1222_U371, P1_R1222_U372, P1_R1222_U373, P1_R1222_U374, P1_R1222_U375, P1_R1222_U376, P1_R1222_U377, P1_R1222_U378, P1_R1222_U379, P1_R1222_U38, P1_R1222_U380, P1_R1222_U381, P1_R1222_U382, P1_R1222_U383, P1_R1222_U384, P1_R1222_U385, P1_R1222_U386, P1_R1222_U387, P1_R1222_U388, P1_R1222_U389, P1_R1222_U39, P1_R1222_U390, P1_R1222_U391, P1_R1222_U392, P1_R1222_U393, P1_R1222_U394, P1_R1222_U395, P1_R1222_U396, P1_R1222_U397, P1_R1222_U398, P1_R1222_U399, P1_R1222_U4, P1_R1222_U40, P1_R1222_U400, P1_R1222_U401, P1_R1222_U402, P1_R1222_U403, P1_R1222_U404, P1_R1222_U405, P1_R1222_U406, P1_R1222_U407, P1_R1222_U408, P1_R1222_U409, P1_R1222_U41, P1_R1222_U410, P1_R1222_U411, P1_R1222_U412, P1_R1222_U413, P1_R1222_U414, P1_R1222_U415, P1_R1222_U416, P1_R1222_U417, P1_R1222_U418, P1_R1222_U419, P1_R1222_U42, P1_R1222_U420, P1_R1222_U421, P1_R1222_U422, P1_R1222_U423, P1_R1222_U424, P1_R1222_U425, P1_R1222_U426, P1_R1222_U427, P1_R1222_U428, P1_R1222_U429, P1_R1222_U43, P1_R1222_U430, P1_R1222_U431, P1_R1222_U432, P1_R1222_U433, P1_R1222_U434, P1_R1222_U435, P1_R1222_U436, P1_R1222_U437, P1_R1222_U438, P1_R1222_U439, P1_R1222_U44, P1_R1222_U440, P1_R1222_U441, P1_R1222_U442, P1_R1222_U443, P1_R1222_U444, P1_R1222_U445, P1_R1222_U446, P1_R1222_U447, P1_R1222_U448, P1_R1222_U449, P1_R1222_U45, P1_R1222_U450, P1_R1222_U451, P1_R1222_U452, P1_R1222_U453, P1_R1222_U454, P1_R1222_U455, P1_R1222_U456, P1_R1222_U457, P1_R1222_U458, P1_R1222_U459, P1_R1222_U46, P1_R1222_U460, P1_R1222_U461, P1_R1222_U462, P1_R1222_U463, P1_R1222_U464, P1_R1222_U465, P1_R1222_U466, P1_R1222_U467, P1_R1222_U468, P1_R1222_U469, P1_R1222_U47, P1_R1222_U470, P1_R1222_U471, P1_R1222_U472, P1_R1222_U473, P1_R1222_U474, P1_R1222_U475, P1_R1222_U476, P1_R1222_U477, P1_R1222_U478, P1_R1222_U479, P1_R1222_U48, P1_R1222_U480, P1_R1222_U481, P1_R1222_U482, P1_R1222_U483, P1_R1222_U484, P1_R1222_U485, P1_R1222_U486, P1_R1222_U487, P1_R1222_U488, P1_R1222_U489, P1_R1222_U49, P1_R1222_U490, P1_R1222_U491, P1_R1222_U492, P1_R1222_U493, P1_R1222_U494, P1_R1222_U495, P1_R1222_U496, P1_R1222_U497, P1_R1222_U498, P1_R1222_U499, P1_R1222_U5, P1_R1222_U50, P1_R1222_U500, P1_R1222_U501, P1_R1222_U502, P1_R1222_U503, P1_R1222_U51, P1_R1222_U52, P1_R1222_U53, P1_R1222_U54, P1_R1222_U55, P1_R1222_U56, P1_R1222_U57, P1_R1222_U58, P1_R1222_U59, P1_R1222_U6, P1_R1222_U60, P1_R1222_U61, P1_R1222_U62, P1_R1222_U63, P1_R1222_U64, P1_R1222_U65, P1_R1222_U66, P1_R1222_U67, P1_R1222_U68, P1_R1222_U69, P1_R1222_U7, P1_R1222_U70, P1_R1222_U71, P1_R1222_U72, P1_R1222_U73, P1_R1222_U74, P1_R1222_U75, P1_R1222_U76, P1_R1222_U77, P1_R1222_U78, P1_R1222_U79, P1_R1222_U8, P1_R1222_U80, P1_R1222_U81, P1_R1222_U82, P1_R1222_U83, P1_R1222_U84, P1_R1222_U85, P1_R1222_U86, P1_R1222_U87, P1_R1222_U88, P1_R1222_U89, P1_R1222_U9, P1_R1222_U90, P1_R1222_U91, P1_R1222_U92, P1_R1222_U93, P1_R1222_U94, P1_R1222_U95, P1_R1222_U96, P1_R1222_U97, P1_R1222_U98, P1_R1222_U99, P1_R1240_U10, P1_R1240_U100, P1_R1240_U101, P1_R1240_U102, P1_R1240_U103, P1_R1240_U104, P1_R1240_U105, P1_R1240_U106, P1_R1240_U107, P1_R1240_U108, P1_R1240_U109, P1_R1240_U11, P1_R1240_U110, P1_R1240_U111, P1_R1240_U112, P1_R1240_U113, P1_R1240_U114, P1_R1240_U115, P1_R1240_U116, P1_R1240_U117, P1_R1240_U118, P1_R1240_U119, P1_R1240_U12, P1_R1240_U120, P1_R1240_U121, P1_R1240_U122, P1_R1240_U123, P1_R1240_U124, P1_R1240_U125, P1_R1240_U126, P1_R1240_U127, P1_R1240_U128, P1_R1240_U129, P1_R1240_U13, P1_R1240_U130, P1_R1240_U131, P1_R1240_U132, P1_R1240_U133, P1_R1240_U134, P1_R1240_U135, P1_R1240_U136, P1_R1240_U137, P1_R1240_U138, P1_R1240_U139, P1_R1240_U14, P1_R1240_U140, P1_R1240_U141, P1_R1240_U142, P1_R1240_U143, P1_R1240_U144, P1_R1240_U145, P1_R1240_U146, P1_R1240_U147, P1_R1240_U148, P1_R1240_U149, P1_R1240_U15, P1_R1240_U150, P1_R1240_U151, P1_R1240_U152, P1_R1240_U153, P1_R1240_U154, P1_R1240_U155, P1_R1240_U156, P1_R1240_U157, P1_R1240_U158, P1_R1240_U159, P1_R1240_U16, P1_R1240_U160, P1_R1240_U161, P1_R1240_U162, P1_R1240_U163, P1_R1240_U164, P1_R1240_U165, P1_R1240_U166, P1_R1240_U167, P1_R1240_U168, P1_R1240_U169, P1_R1240_U17, P1_R1240_U170, P1_R1240_U171, P1_R1240_U172, P1_R1240_U173, P1_R1240_U174, P1_R1240_U175, P1_R1240_U176, P1_R1240_U177, P1_R1240_U178, P1_R1240_U179, P1_R1240_U18, P1_R1240_U180, P1_R1240_U181, P1_R1240_U182, P1_R1240_U183, P1_R1240_U184, P1_R1240_U185, P1_R1240_U186, P1_R1240_U187, P1_R1240_U188, P1_R1240_U189, P1_R1240_U19, P1_R1240_U190, P1_R1240_U191, P1_R1240_U192, P1_R1240_U193, P1_R1240_U194, P1_R1240_U195, P1_R1240_U196, P1_R1240_U197, P1_R1240_U198, P1_R1240_U199, P1_R1240_U20, P1_R1240_U200, P1_R1240_U201, P1_R1240_U202, P1_R1240_U203, P1_R1240_U204, P1_R1240_U205, P1_R1240_U206, P1_R1240_U207, P1_R1240_U208, P1_R1240_U209, P1_R1240_U21, P1_R1240_U210, P1_R1240_U211, P1_R1240_U212, P1_R1240_U213, P1_R1240_U214, P1_R1240_U215, P1_R1240_U216, P1_R1240_U217, P1_R1240_U218, P1_R1240_U219, P1_R1240_U22, P1_R1240_U220, P1_R1240_U221, P1_R1240_U222, P1_R1240_U223, P1_R1240_U224, P1_R1240_U225, P1_R1240_U226, P1_R1240_U227, P1_R1240_U228, P1_R1240_U229, P1_R1240_U23, P1_R1240_U230, P1_R1240_U231, P1_R1240_U232, P1_R1240_U233, P1_R1240_U234, P1_R1240_U235, P1_R1240_U236, P1_R1240_U237, P1_R1240_U238, P1_R1240_U239, P1_R1240_U24, P1_R1240_U240, P1_R1240_U241, P1_R1240_U242, P1_R1240_U243, P1_R1240_U244, P1_R1240_U245, P1_R1240_U246, P1_R1240_U247, P1_R1240_U248, P1_R1240_U249, P1_R1240_U25, P1_R1240_U250, P1_R1240_U251, P1_R1240_U252, P1_R1240_U253, P1_R1240_U254, P1_R1240_U255, P1_R1240_U256, P1_R1240_U257, P1_R1240_U258, P1_R1240_U259, P1_R1240_U26, P1_R1240_U260, P1_R1240_U261, P1_R1240_U262, P1_R1240_U263, P1_R1240_U264, P1_R1240_U265, P1_R1240_U266, P1_R1240_U267, P1_R1240_U268, P1_R1240_U269, P1_R1240_U27, P1_R1240_U270, P1_R1240_U271, P1_R1240_U272, P1_R1240_U273, P1_R1240_U274, P1_R1240_U275, P1_R1240_U276, P1_R1240_U277, P1_R1240_U278, P1_R1240_U279, P1_R1240_U28, P1_R1240_U280, P1_R1240_U281, P1_R1240_U282, P1_R1240_U283, P1_R1240_U284, P1_R1240_U285, P1_R1240_U286, P1_R1240_U287, P1_R1240_U288, P1_R1240_U289, P1_R1240_U29, P1_R1240_U290, P1_R1240_U291, P1_R1240_U292, P1_R1240_U293, P1_R1240_U294, P1_R1240_U295, P1_R1240_U296, P1_R1240_U297, P1_R1240_U298, P1_R1240_U299, P1_R1240_U30, P1_R1240_U300, P1_R1240_U301, P1_R1240_U302, P1_R1240_U303, P1_R1240_U304, P1_R1240_U305, P1_R1240_U306, P1_R1240_U307, P1_R1240_U308, P1_R1240_U309, P1_R1240_U31, P1_R1240_U310, P1_R1240_U311, P1_R1240_U312, P1_R1240_U313, P1_R1240_U314, P1_R1240_U315, P1_R1240_U316, P1_R1240_U317, P1_R1240_U318, P1_R1240_U319, P1_R1240_U32, P1_R1240_U320, P1_R1240_U321, P1_R1240_U322, P1_R1240_U323, P1_R1240_U324, P1_R1240_U325, P1_R1240_U326, P1_R1240_U327, P1_R1240_U328, P1_R1240_U329, P1_R1240_U33, P1_R1240_U330, P1_R1240_U331, P1_R1240_U332, P1_R1240_U333, P1_R1240_U334, P1_R1240_U335, P1_R1240_U336, P1_R1240_U337, P1_R1240_U338, P1_R1240_U339, P1_R1240_U34, P1_R1240_U340, P1_R1240_U341, P1_R1240_U342, P1_R1240_U343, P1_R1240_U344, P1_R1240_U345, P1_R1240_U346, P1_R1240_U347, P1_R1240_U348, P1_R1240_U349, P1_R1240_U35, P1_R1240_U350, P1_R1240_U351, P1_R1240_U352, P1_R1240_U353, P1_R1240_U354, P1_R1240_U355, P1_R1240_U356, P1_R1240_U357, P1_R1240_U358, P1_R1240_U359, P1_R1240_U36, P1_R1240_U360, P1_R1240_U361, P1_R1240_U362, P1_R1240_U363, P1_R1240_U364, P1_R1240_U365, P1_R1240_U366, P1_R1240_U367, P1_R1240_U368, P1_R1240_U369, P1_R1240_U37, P1_R1240_U370, P1_R1240_U371, P1_R1240_U372, P1_R1240_U373, P1_R1240_U374, P1_R1240_U375, P1_R1240_U376, P1_R1240_U377, P1_R1240_U378, P1_R1240_U379, P1_R1240_U38, P1_R1240_U380, P1_R1240_U381, P1_R1240_U382, P1_R1240_U383, P1_R1240_U384, P1_R1240_U385, P1_R1240_U386, P1_R1240_U387, P1_R1240_U388, P1_R1240_U389, P1_R1240_U39, P1_R1240_U390, P1_R1240_U391, P1_R1240_U392, P1_R1240_U393, P1_R1240_U394, P1_R1240_U395, P1_R1240_U396, P1_R1240_U397, P1_R1240_U398, P1_R1240_U399, P1_R1240_U4, P1_R1240_U40, P1_R1240_U400, P1_R1240_U401, P1_R1240_U402, P1_R1240_U403, P1_R1240_U404, P1_R1240_U405, P1_R1240_U406, P1_R1240_U407, P1_R1240_U408, P1_R1240_U409, P1_R1240_U41, P1_R1240_U410, P1_R1240_U411, P1_R1240_U412, P1_R1240_U413, P1_R1240_U414, P1_R1240_U415, P1_R1240_U416, P1_R1240_U417, P1_R1240_U418, P1_R1240_U419, P1_R1240_U42, P1_R1240_U420, P1_R1240_U421, P1_R1240_U422, P1_R1240_U423, P1_R1240_U424, P1_R1240_U425, P1_R1240_U426, P1_R1240_U427, P1_R1240_U428, P1_R1240_U429, P1_R1240_U43, P1_R1240_U430, P1_R1240_U431, P1_R1240_U432, P1_R1240_U433, P1_R1240_U434, P1_R1240_U435, P1_R1240_U436, P1_R1240_U437, P1_R1240_U438, P1_R1240_U439, P1_R1240_U44, P1_R1240_U440, P1_R1240_U441, P1_R1240_U442, P1_R1240_U443, P1_R1240_U444, P1_R1240_U445, P1_R1240_U446, P1_R1240_U447, P1_R1240_U448, P1_R1240_U449, P1_R1240_U45, P1_R1240_U450, P1_R1240_U451, P1_R1240_U452, P1_R1240_U453, P1_R1240_U454, P1_R1240_U455, P1_R1240_U456, P1_R1240_U457, P1_R1240_U458, P1_R1240_U459, P1_R1240_U46, P1_R1240_U460, P1_R1240_U461, P1_R1240_U462, P1_R1240_U463, P1_R1240_U464, P1_R1240_U465, P1_R1240_U466, P1_R1240_U467, P1_R1240_U468, P1_R1240_U469, P1_R1240_U47, P1_R1240_U470, P1_R1240_U471, P1_R1240_U472, P1_R1240_U473, P1_R1240_U474, P1_R1240_U475, P1_R1240_U476, P1_R1240_U477, P1_R1240_U478, P1_R1240_U479, P1_R1240_U48, P1_R1240_U480, P1_R1240_U481, P1_R1240_U482, P1_R1240_U483, P1_R1240_U484, P1_R1240_U485, P1_R1240_U486, P1_R1240_U487, P1_R1240_U488, P1_R1240_U489, P1_R1240_U49, P1_R1240_U490, P1_R1240_U491, P1_R1240_U492, P1_R1240_U493, P1_R1240_U494, P1_R1240_U495, P1_R1240_U496, P1_R1240_U497, P1_R1240_U498, P1_R1240_U499, P1_R1240_U5, P1_R1240_U50, P1_R1240_U500, P1_R1240_U501, P1_R1240_U502, P1_R1240_U503, P1_R1240_U51, P1_R1240_U52, P1_R1240_U53, P1_R1240_U54, P1_R1240_U55, P1_R1240_U56, P1_R1240_U57, P1_R1240_U58, P1_R1240_U59, P1_R1240_U6, P1_R1240_U60, P1_R1240_U61, P1_R1240_U62, P1_R1240_U63, P1_R1240_U64, P1_R1240_U65, P1_R1240_U66, P1_R1240_U67, P1_R1240_U68, P1_R1240_U69, P1_R1240_U7, P1_R1240_U70, P1_R1240_U71, P1_R1240_U72, P1_R1240_U73, P1_R1240_U74, P1_R1240_U75, P1_R1240_U76, P1_R1240_U77, P1_R1240_U78, P1_R1240_U79, P1_R1240_U8, P1_R1240_U80, P1_R1240_U81, P1_R1240_U82, P1_R1240_U83, P1_R1240_U84, P1_R1240_U85, P1_R1240_U86, P1_R1240_U87, P1_R1240_U88, P1_R1240_U89, P1_R1240_U9, P1_R1240_U90, P1_R1240_U91, P1_R1240_U92, P1_R1240_U93, P1_R1240_U94, P1_R1240_U95, P1_R1240_U96, P1_R1240_U97, P1_R1240_U98, P1_R1240_U99, P1_R1282_U10, P1_R1282_U100, P1_R1282_U101, P1_R1282_U102, P1_R1282_U103, P1_R1282_U104, P1_R1282_U105, P1_R1282_U106, P1_R1282_U107, P1_R1282_U108, P1_R1282_U109, P1_R1282_U11, P1_R1282_U110, P1_R1282_U111, P1_R1282_U112, P1_R1282_U113, P1_R1282_U114, P1_R1282_U115, P1_R1282_U116, P1_R1282_U117, P1_R1282_U118, P1_R1282_U119, P1_R1282_U12, P1_R1282_U120, P1_R1282_U121, P1_R1282_U122, P1_R1282_U123, P1_R1282_U124, P1_R1282_U125, P1_R1282_U126, P1_R1282_U127, P1_R1282_U128, P1_R1282_U129, P1_R1282_U13, P1_R1282_U130, P1_R1282_U131, P1_R1282_U132, P1_R1282_U133, P1_R1282_U134, P1_R1282_U135, P1_R1282_U136, P1_R1282_U137, P1_R1282_U138, P1_R1282_U139, P1_R1282_U14, P1_R1282_U140, P1_R1282_U141, P1_R1282_U142, P1_R1282_U143, P1_R1282_U144, P1_R1282_U145, P1_R1282_U146, P1_R1282_U147, P1_R1282_U148, P1_R1282_U149, P1_R1282_U15, P1_R1282_U150, P1_R1282_U151, P1_R1282_U152, P1_R1282_U153, P1_R1282_U154, P1_R1282_U155, P1_R1282_U156, P1_R1282_U157, P1_R1282_U158, P1_R1282_U159, P1_R1282_U16, P1_R1282_U17, P1_R1282_U18, P1_R1282_U19, P1_R1282_U20, P1_R1282_U21, P1_R1282_U22, P1_R1282_U23, P1_R1282_U24, P1_R1282_U25, P1_R1282_U26, P1_R1282_U27, P1_R1282_U28, P1_R1282_U29, P1_R1282_U30, P1_R1282_U31, P1_R1282_U32, P1_R1282_U33, P1_R1282_U34, P1_R1282_U35, P1_R1282_U36, P1_R1282_U37, P1_R1282_U38, P1_R1282_U39, P1_R1282_U40, P1_R1282_U41, P1_R1282_U42, P1_R1282_U43, P1_R1282_U44, P1_R1282_U45, P1_R1282_U46, P1_R1282_U47, P1_R1282_U48, P1_R1282_U49, P1_R1282_U50, P1_R1282_U51, P1_R1282_U52, P1_R1282_U53, P1_R1282_U54, P1_R1282_U55, P1_R1282_U56, P1_R1282_U57, P1_R1282_U58, P1_R1282_U59, P1_R1282_U6, P1_R1282_U60, P1_R1282_U61, P1_R1282_U62, P1_R1282_U63, P1_R1282_U64, P1_R1282_U65, P1_R1282_U66, P1_R1282_U67, P1_R1282_U68, P1_R1282_U69, P1_R1282_U7, P1_R1282_U70, P1_R1282_U71, P1_R1282_U72, P1_R1282_U73, P1_R1282_U74, P1_R1282_U75, P1_R1282_U76, P1_R1282_U77, P1_R1282_U78, P1_R1282_U79, P1_R1282_U8, P1_R1282_U80, P1_R1282_U81, P1_R1282_U82, P1_R1282_U83, P1_R1282_U84, P1_R1282_U85, P1_R1282_U86, P1_R1282_U87, P1_R1282_U88, P1_R1282_U89, P1_R1282_U9, P1_R1282_U90, P1_R1282_U91, P1_R1282_U92, P1_R1282_U93, P1_R1282_U94, P1_R1282_U95, P1_R1282_U96, P1_R1282_U97, P1_R1282_U98, P1_R1282_U99, P1_R1309_U10, P1_R1309_U6, P1_R1309_U7, P1_R1309_U8, P1_R1309_U9, P1_R1352_U6, P1_R1352_U7, P1_R1360_U10, P1_R1360_U100, P1_R1360_U101, P1_R1360_U102, P1_R1360_U103, P1_R1360_U104, P1_R1360_U105, P1_R1360_U106, P1_R1360_U107, P1_R1360_U108, P1_R1360_U109, P1_R1360_U11, P1_R1360_U110, P1_R1360_U111, P1_R1360_U112, P1_R1360_U113, P1_R1360_U114, P1_R1360_U115, P1_R1360_U116, P1_R1360_U117, P1_R1360_U118, P1_R1360_U119, P1_R1360_U12, P1_R1360_U120, P1_R1360_U121, P1_R1360_U122, P1_R1360_U123, P1_R1360_U124, P1_R1360_U125, P1_R1360_U126, P1_R1360_U127, P1_R1360_U128, P1_R1360_U129, P1_R1360_U13, P1_R1360_U130, P1_R1360_U131, P1_R1360_U132, P1_R1360_U133, P1_R1360_U134, P1_R1360_U135, P1_R1360_U136, P1_R1360_U137, P1_R1360_U138, P1_R1360_U139, P1_R1360_U14, P1_R1360_U140, P1_R1360_U141, P1_R1360_U142, P1_R1360_U143, P1_R1360_U144, P1_R1360_U145, P1_R1360_U146, P1_R1360_U147, P1_R1360_U148, P1_R1360_U149, P1_R1360_U15, P1_R1360_U150, P1_R1360_U151, P1_R1360_U152, P1_R1360_U153, P1_R1360_U154, P1_R1360_U155, P1_R1360_U156, P1_R1360_U157, P1_R1360_U158, P1_R1360_U159, P1_R1360_U16, P1_R1360_U160, P1_R1360_U161, P1_R1360_U162, P1_R1360_U163, P1_R1360_U164, P1_R1360_U165, P1_R1360_U166, P1_R1360_U167, P1_R1360_U168, P1_R1360_U169, P1_R1360_U17, P1_R1360_U170, P1_R1360_U171, P1_R1360_U172, P1_R1360_U173, P1_R1360_U174, P1_R1360_U175, P1_R1360_U176, P1_R1360_U177, P1_R1360_U178, P1_R1360_U179, P1_R1360_U18, P1_R1360_U180, P1_R1360_U181, P1_R1360_U182, P1_R1360_U183, P1_R1360_U184, P1_R1360_U185, P1_R1360_U186, P1_R1360_U187, P1_R1360_U188, P1_R1360_U189, P1_R1360_U19, P1_R1360_U190, P1_R1360_U191, P1_R1360_U192, P1_R1360_U193, P1_R1360_U194, P1_R1360_U195, P1_R1360_U196, P1_R1360_U197, P1_R1360_U198, P1_R1360_U199, P1_R1360_U20, P1_R1360_U200, P1_R1360_U201, P1_R1360_U202, P1_R1360_U203, P1_R1360_U204, P1_R1360_U205, P1_R1360_U21, P1_R1360_U22, P1_R1360_U23, P1_R1360_U24, P1_R1360_U25, P1_R1360_U26, P1_R1360_U27, P1_R1360_U28, P1_R1360_U29, P1_R1360_U30, P1_R1360_U31, P1_R1360_U32, P1_R1360_U33, P1_R1360_U34, P1_R1360_U35, P1_R1360_U36, P1_R1360_U37, P1_R1360_U38, P1_R1360_U39, P1_R1360_U40, P1_R1360_U41, P1_R1360_U42, P1_R1360_U43, P1_R1360_U44, P1_R1360_U45, P1_R1360_U46, P1_R1360_U47, P1_R1360_U48, P1_R1360_U49, P1_R1360_U50, P1_R1360_U51, P1_R1360_U52, P1_R1360_U53, P1_R1360_U54, P1_R1360_U55, P1_R1360_U56, P1_R1360_U57, P1_R1360_U58, P1_R1360_U59, P1_R1360_U6, P1_R1360_U60, P1_R1360_U61, P1_R1360_U62, P1_R1360_U63, P1_R1360_U64, P1_R1360_U65, P1_R1360_U66, P1_R1360_U67, P1_R1360_U68, P1_R1360_U69, P1_R1360_U7, P1_R1360_U70, P1_R1360_U71, P1_R1360_U72, P1_R1360_U73, P1_R1360_U74, P1_R1360_U75, P1_R1360_U76, P1_R1360_U77, P1_R1360_U78, P1_R1360_U79, P1_R1360_U8, P1_R1360_U80, P1_R1360_U81, P1_R1360_U82, P1_R1360_U83, P1_R1360_U84, P1_R1360_U85, P1_R1360_U86, P1_R1360_U87, P1_R1360_U88, P1_R1360_U89, P1_R1360_U9, P1_R1360_U90, P1_R1360_U91, P1_R1360_U92, P1_R1360_U93, P1_R1360_U94, P1_R1360_U95, P1_R1360_U96, P1_R1360_U97, P1_R1360_U98, P1_R1360_U99, P1_R1375_U10, P1_R1375_U100, P1_R1375_U101, P1_R1375_U102, P1_R1375_U103, P1_R1375_U104, P1_R1375_U105, P1_R1375_U106, P1_R1375_U107, P1_R1375_U108, P1_R1375_U109, P1_R1375_U11, P1_R1375_U110, P1_R1375_U111, P1_R1375_U112, P1_R1375_U113, P1_R1375_U114, P1_R1375_U115, P1_R1375_U116, P1_R1375_U117, P1_R1375_U118, P1_R1375_U119, P1_R1375_U12, P1_R1375_U120, P1_R1375_U121, P1_R1375_U122, P1_R1375_U123, P1_R1375_U124, P1_R1375_U125, P1_R1375_U126, P1_R1375_U127, P1_R1375_U128, P1_R1375_U129, P1_R1375_U13, P1_R1375_U130, P1_R1375_U131, P1_R1375_U132, P1_R1375_U133, P1_R1375_U134, P1_R1375_U135, P1_R1375_U136, P1_R1375_U137, P1_R1375_U138, P1_R1375_U139, P1_R1375_U14, P1_R1375_U140, P1_R1375_U141, P1_R1375_U142, P1_R1375_U143, P1_R1375_U144, P1_R1375_U145, P1_R1375_U146, P1_R1375_U147, P1_R1375_U148, P1_R1375_U149, P1_R1375_U15, P1_R1375_U150, P1_R1375_U151, P1_R1375_U152, P1_R1375_U153, P1_R1375_U154, P1_R1375_U155, P1_R1375_U156, P1_R1375_U157, P1_R1375_U158, P1_R1375_U159, P1_R1375_U16, P1_R1375_U160, P1_R1375_U161, P1_R1375_U162, P1_R1375_U163, P1_R1375_U164, P1_R1375_U165, P1_R1375_U166, P1_R1375_U167, P1_R1375_U168, P1_R1375_U169, P1_R1375_U17, P1_R1375_U170, P1_R1375_U171, P1_R1375_U172, P1_R1375_U173, P1_R1375_U174, P1_R1375_U175, P1_R1375_U176, P1_R1375_U177, P1_R1375_U178, P1_R1375_U179, P1_R1375_U18, P1_R1375_U180, P1_R1375_U181, P1_R1375_U182, P1_R1375_U183, P1_R1375_U184, P1_R1375_U185, P1_R1375_U186, P1_R1375_U187, P1_R1375_U188, P1_R1375_U189, P1_R1375_U19, P1_R1375_U190, P1_R1375_U191, P1_R1375_U192, P1_R1375_U193, P1_R1375_U194, P1_R1375_U195, P1_R1375_U196, P1_R1375_U197, P1_R1375_U198, P1_R1375_U199, P1_R1375_U20, P1_R1375_U200, P1_R1375_U201, P1_R1375_U202, P1_R1375_U203, P1_R1375_U204, P1_R1375_U205, P1_R1375_U206, P1_R1375_U207, P1_R1375_U21, P1_R1375_U22, P1_R1375_U23, P1_R1375_U24, P1_R1375_U25, P1_R1375_U26, P1_R1375_U27, P1_R1375_U28, P1_R1375_U29, P1_R1375_U30, P1_R1375_U31, P1_R1375_U32, P1_R1375_U33, P1_R1375_U34, P1_R1375_U35, P1_R1375_U36, P1_R1375_U37, P1_R1375_U38, P1_R1375_U39, P1_R1375_U40, P1_R1375_U41, P1_R1375_U42, P1_R1375_U43, P1_R1375_U44, P1_R1375_U45, P1_R1375_U46, P1_R1375_U47, P1_R1375_U48, P1_R1375_U49, P1_R1375_U50, P1_R1375_U51, P1_R1375_U52, P1_R1375_U53, P1_R1375_U54, P1_R1375_U55, P1_R1375_U56, P1_R1375_U57, P1_R1375_U58, P1_R1375_U59, P1_R1375_U6, P1_R1375_U60, P1_R1375_U61, P1_R1375_U62, P1_R1375_U63, P1_R1375_U64, P1_R1375_U65, P1_R1375_U66, P1_R1375_U67, P1_R1375_U68, P1_R1375_U69, P1_R1375_U7, P1_R1375_U70, P1_R1375_U71, P1_R1375_U72, P1_R1375_U73, P1_R1375_U74, P1_R1375_U75, P1_R1375_U76, P1_R1375_U77, P1_R1375_U78, P1_R1375_U79, P1_R1375_U8, P1_R1375_U80, P1_R1375_U81, P1_R1375_U82, P1_R1375_U83, P1_R1375_U84, P1_R1375_U85, P1_R1375_U86, P1_R1375_U87, P1_R1375_U88, P1_R1375_U89, P1_R1375_U9, P1_R1375_U90, P1_R1375_U91, P1_R1375_U92, P1_R1375_U93, P1_R1375_U94, P1_R1375_U95, P1_R1375_U96, P1_R1375_U97, P1_R1375_U98, P1_R1375_U99, P1_SUB_84_U10, P1_SUB_84_U100, P1_SUB_84_U101, P1_SUB_84_U102, P1_SUB_84_U103, P1_SUB_84_U104, P1_SUB_84_U105, P1_SUB_84_U106, P1_SUB_84_U107, P1_SUB_84_U108, P1_SUB_84_U109, P1_SUB_84_U11, P1_SUB_84_U110, P1_SUB_84_U111, P1_SUB_84_U112, P1_SUB_84_U113, P1_SUB_84_U114, P1_SUB_84_U115, P1_SUB_84_U116, P1_SUB_84_U117, P1_SUB_84_U118, P1_SUB_84_U119, P1_SUB_84_U12, P1_SUB_84_U120, P1_SUB_84_U121, P1_SUB_84_U122, P1_SUB_84_U123, P1_SUB_84_U124, P1_SUB_84_U125, P1_SUB_84_U126, P1_SUB_84_U127, P1_SUB_84_U128, P1_SUB_84_U129, P1_SUB_84_U13, P1_SUB_84_U130, P1_SUB_84_U131, P1_SUB_84_U132, P1_SUB_84_U133, P1_SUB_84_U134, P1_SUB_84_U135, P1_SUB_84_U136, P1_SUB_84_U137, P1_SUB_84_U138, P1_SUB_84_U139, P1_SUB_84_U14, P1_SUB_84_U140, P1_SUB_84_U141, P1_SUB_84_U142, P1_SUB_84_U143, P1_SUB_84_U144, P1_SUB_84_U145, P1_SUB_84_U146, P1_SUB_84_U147, P1_SUB_84_U148, P1_SUB_84_U149, P1_SUB_84_U15, P1_SUB_84_U150, P1_SUB_84_U151, P1_SUB_84_U152, P1_SUB_84_U153, P1_SUB_84_U154, P1_SUB_84_U155, P1_SUB_84_U156, P1_SUB_84_U157, P1_SUB_84_U158, P1_SUB_84_U159, P1_SUB_84_U16, P1_SUB_84_U160, P1_SUB_84_U161, P1_SUB_84_U162, P1_SUB_84_U163, P1_SUB_84_U164, P1_SUB_84_U165, P1_SUB_84_U166, P1_SUB_84_U167, P1_SUB_84_U168, P1_SUB_84_U169, P1_SUB_84_U17, P1_SUB_84_U170, P1_SUB_84_U171, P1_SUB_84_U172, P1_SUB_84_U173, P1_SUB_84_U174, P1_SUB_84_U175, P1_SUB_84_U176, P1_SUB_84_U177, P1_SUB_84_U178, P1_SUB_84_U179, P1_SUB_84_U18, P1_SUB_84_U180, P1_SUB_84_U181, P1_SUB_84_U182, P1_SUB_84_U183, P1_SUB_84_U184, P1_SUB_84_U185, P1_SUB_84_U186, P1_SUB_84_U187, P1_SUB_84_U188, P1_SUB_84_U189, P1_SUB_84_U19, P1_SUB_84_U190, P1_SUB_84_U191, P1_SUB_84_U192, P1_SUB_84_U193, P1_SUB_84_U194, P1_SUB_84_U195, P1_SUB_84_U196, P1_SUB_84_U197, P1_SUB_84_U198, P1_SUB_84_U199, P1_SUB_84_U20, P1_SUB_84_U200, P1_SUB_84_U201, P1_SUB_84_U202, P1_SUB_84_U203, P1_SUB_84_U204, P1_SUB_84_U205, P1_SUB_84_U206, P1_SUB_84_U207, P1_SUB_84_U208, P1_SUB_84_U209, P1_SUB_84_U21, P1_SUB_84_U210, P1_SUB_84_U211, P1_SUB_84_U212, P1_SUB_84_U213, P1_SUB_84_U214, P1_SUB_84_U215, P1_SUB_84_U216, P1_SUB_84_U217, P1_SUB_84_U218, P1_SUB_84_U219, P1_SUB_84_U22, P1_SUB_84_U220, P1_SUB_84_U221, P1_SUB_84_U222, P1_SUB_84_U223, P1_SUB_84_U224, P1_SUB_84_U225, P1_SUB_84_U226, P1_SUB_84_U227, P1_SUB_84_U228, P1_SUB_84_U229, P1_SUB_84_U23, P1_SUB_84_U230, P1_SUB_84_U231, P1_SUB_84_U232, P1_SUB_84_U233, P1_SUB_84_U234, P1_SUB_84_U235, P1_SUB_84_U236, P1_SUB_84_U237, P1_SUB_84_U238, P1_SUB_84_U239, P1_SUB_84_U24, P1_SUB_84_U240, P1_SUB_84_U241, P1_SUB_84_U242, P1_SUB_84_U243, P1_SUB_84_U244, P1_SUB_84_U245, P1_SUB_84_U246, P1_SUB_84_U247, P1_SUB_84_U248, P1_SUB_84_U249, P1_SUB_84_U25, P1_SUB_84_U250, P1_SUB_84_U251, P1_SUB_84_U26, P1_SUB_84_U27, P1_SUB_84_U28, P1_SUB_84_U29, P1_SUB_84_U30, P1_SUB_84_U31, P1_SUB_84_U32, P1_SUB_84_U33, P1_SUB_84_U34, P1_SUB_84_U35, P1_SUB_84_U36, P1_SUB_84_U37, P1_SUB_84_U38, P1_SUB_84_U39, P1_SUB_84_U40, P1_SUB_84_U41, P1_SUB_84_U42, P1_SUB_84_U43, P1_SUB_84_U44, P1_SUB_84_U45, P1_SUB_84_U46, P1_SUB_84_U47, P1_SUB_84_U48, P1_SUB_84_U49, P1_SUB_84_U50, P1_SUB_84_U51, P1_SUB_84_U52, P1_SUB_84_U53, P1_SUB_84_U54, P1_SUB_84_U55, P1_SUB_84_U56, P1_SUB_84_U57, P1_SUB_84_U58, P1_SUB_84_U59, P1_SUB_84_U6, P1_SUB_84_U60, P1_SUB_84_U61, P1_SUB_84_U62, P1_SUB_84_U63, P1_SUB_84_U64, P1_SUB_84_U65, P1_SUB_84_U66, P1_SUB_84_U67, P1_SUB_84_U68, P1_SUB_84_U69, P1_SUB_84_U7, P1_SUB_84_U70, P1_SUB_84_U71, P1_SUB_84_U72, P1_SUB_84_U73, P1_SUB_84_U74, P1_SUB_84_U75, P1_SUB_84_U76, P1_SUB_84_U77, P1_SUB_84_U78, P1_SUB_84_U79, P1_SUB_84_U8, P1_SUB_84_U80, P1_SUB_84_U81, P1_SUB_84_U82, P1_SUB_84_U83, P1_SUB_84_U84, P1_SUB_84_U85, P1_SUB_84_U86, P1_SUB_84_U87, P1_SUB_84_U88, P1_SUB_84_U89, P1_SUB_84_U9, P1_SUB_84_U90, P1_SUB_84_U91, P1_SUB_84_U92, P1_SUB_84_U93, P1_SUB_84_U94, P1_SUB_84_U95, P1_SUB_84_U96, P1_SUB_84_U97, P1_SUB_84_U98, P1_SUB_84_U99, P1_U3014, P1_U3015, P1_U3016, P1_U3017, P1_U3018, P1_U3019, P1_U3020, P1_U3021, P1_U3022, P1_U3023, P1_U3024, P1_U3025, P1_U3026, P1_U3027, P1_U3028, P1_U3029, P1_U3030, P1_U3031, P1_U3032, P1_U3033, P1_U3034, P1_U3035, P1_U3036, P1_U3037, P1_U3038, P1_U3039, P1_U3040, P1_U3041, P1_U3042, P1_U3043, P1_U3044, P1_U3045, P1_U3046, P1_U3047, P1_U3048, P1_U3049, P1_U3050, P1_U3051, P1_U3052, P1_U3053, P1_U3054, P1_U3055, P1_U3056, P1_U3057, P1_U3058, P1_U3059, P1_U3060, P1_U3061, P1_U3062, P1_U3063, P1_U3064, P1_U3065, P1_U3066, P1_U3067, P1_U3068, P1_U3069, P1_U3070, P1_U3071, P1_U3072, P1_U3073, P1_U3074, P1_U3075, P1_U3076, P1_U3077, P1_U3078, P1_U3079, P1_U3080, P1_U3081, P1_U3082, P1_U3083, P1_U3084, P1_U3087, P1_U3088, P1_U3089, P1_U3090, P1_U3091, P1_U3092, P1_U3093, P1_U3094, P1_U3095, P1_U3096, P1_U3097, P1_U3098, P1_U3099, P1_U3100, P1_U3101, P1_U3102, P1_U3103, P1_U3104, P1_U3105, P1_U3106, P1_U3107, P1_U3108, P1_U3109, P1_U3110, P1_U3111, P1_U3112, P1_U3113, P1_U3114, P1_U3115, P1_U3116, P1_U3117, P1_U3118, P1_U3119, P1_U3120, P1_U3121, P1_U3122, P1_U3123, P1_U3124, P1_U3125, P1_U3126, P1_U3127, P1_U3128, P1_U3129, P1_U3130, P1_U3131, P1_U3132, P1_U3133, P1_U3134, P1_U3135, P1_U3136, P1_U3137, P1_U3138, P1_U3139, P1_U3140, P1_U3141, P1_U3142, P1_U3143, P1_U3144, P1_U3145, P1_U3146, P1_U3147, P1_U3148, P1_U3149, P1_U3150, P1_U3151, P1_U3152, P1_U3153, P1_U3154, P1_U3155, P1_U3156, P1_U3157, P1_U3158, P1_U3159, P1_U3160, P1_U3161, P1_U3162, P1_U3163, P1_U3164, P1_U3165, P1_U3166, P1_U3167, P1_U3168, P1_U3169, P1_U3170, P1_U3171, P1_U3172, P1_U3173, P1_U3174, P1_U3175, P1_U3176, P1_U3177, P1_U3178, P1_U3179, P1_U3180, P1_U3181, P1_U3182, P1_U3183, P1_U3184, P1_U3185, P1_U3186, P1_U3187, P1_U3188, P1_U3189, P1_U3190, P1_U3191, P1_U3192, P1_U3193, P1_U3194, P1_U3195, P1_U3196, P1_U3197, P1_U3198, P1_U3199, P1_U3200, P1_U3201, P1_U3202, P1_U3203, P1_U3204, P1_U3205, P1_U3206, P1_U3207, P1_U3208, P1_U3209, P1_U3210, P1_U3211, P1_U3212, P1_U3357, P1_U3358, P1_U3359, P1_U3360, P1_U3361, P1_U3362, P1_U3363, P1_U3364, P1_U3365, P1_U3366, P1_U3367, P1_U3368, P1_U3369, P1_U3370, P1_U3371, P1_U3372, P1_U3373, P1_U3374, P1_U3375, P1_U3376, P1_U3377, P1_U3378, P1_U3379, P1_U3380, P1_U3381, P1_U3382, P1_U3383, P1_U3384, P1_U3385, P1_U3386, P1_U3387, P1_U3388, P1_U3389, P1_U3390, P1_U3391, P1_U3392, P1_U3393, P1_U3394, P1_U3395, P1_U3396, P1_U3397, P1_U3398, P1_U3399, P1_U3400, P1_U3401, P1_U3402, P1_U3403, P1_U3404, P1_U3405, P1_U3406, P1_U3407, P1_U3408, P1_U3409, P1_U3410, P1_U3411, P1_U3412, P1_U3413, P1_U3414, P1_U3415, P1_U3416, P1_U3417, P1_U3418, P1_U3419, P1_U3420, P1_U3421, P1_U3422, P1_U3423, P1_U3424, P1_U3425, P1_U3426, P1_U3427, P1_U3428, P1_U3429, P1_U3430, P1_U3431, P1_U3432, P1_U3433, P1_U3434, P1_U3435, P1_U3436, P1_U3437, P1_U3438, P1_U3441, P1_U3442, P1_U3443, P1_U3444, P1_U3445, P1_U3446, P1_U3447, P1_U3448, P1_U3449, P1_U3450, P1_U3451, P1_U3452, P1_U3454, P1_U3455, P1_U3457, P1_U3458, P1_U3460, P1_U3461, P1_U3463, P1_U3464, P1_U3466, P1_U3467, P1_U3469, P1_U3470, P1_U3472, P1_U3473, P1_U3475, P1_U3476, P1_U3478, P1_U3479, P1_U3481, P1_U3482, P1_U3484, P1_U3485, P1_U3487, P1_U3488, P1_U3490, P1_U3491, P1_U3493, P1_U3494, P1_U3496, P1_U3497, P1_U3499, P1_U3500, P1_U3502, P1_U3503, P1_U3505, P1_U3506, P1_U3508, P1_U3586, P1_U3587, P1_U3588, P1_U3589, P1_U3590, P1_U3591, P1_U3592, P1_U3593, P1_U3594, P1_U3595, P1_U3596, P1_U3597, P1_U3598, P1_U3599, P1_U3600, P1_U3601, P1_U3602, P1_U3603, P1_U3604, P1_U3605, P1_U3606, P1_U3607, P1_U3608, P1_U3609, P1_U3610, P1_U3611, P1_U3612, P1_U3613, P1_U3614, P1_U3615, P1_U3616, P1_U3617, P1_U3618, P1_U3619, P1_U3620, P1_U3621, P1_U3622, P1_U3623, P1_U3624, P1_U3625, P1_U3626, P1_U3627, P1_U3628, P1_U3629, P1_U3630, P1_U3631, P1_U3632, P1_U3633, P1_U3634, P1_U3635, P1_U3636, P1_U3637, P1_U3638, P1_U3639, P1_U3640, P1_U3641, P1_U3642, P1_U3643, P1_U3644, P1_U3645, P1_U3646, P1_U3647, P1_U3648, P1_U3649, P1_U3650, P1_U3651, P1_U3652, P1_U3653, P1_U3654, P1_U3655, P1_U3656, P1_U3657, P1_U3658, P1_U3659, P1_U3660, P1_U3661, P1_U3662, P1_U3663, P1_U3664, P1_U3665, P1_U3666, P1_U3667, P1_U3668, P1_U3669, P1_U3670, P1_U3671, P1_U3672, P1_U3673, P1_U3674, P1_U3675, P1_U3676, P1_U3677, P1_U3678, P1_U3679, P1_U3680, P1_U3681, P1_U3682, P1_U3683, P1_U3684, P1_U3685, P1_U3686, P1_U3687, P1_U3688, P1_U3689, P1_U3690, P1_U3691, P1_U3692, P1_U3693, P1_U3694, P1_U3695, P1_U3696, P1_U3697, P1_U3698, P1_U3699, P1_U3700, P1_U3701, P1_U3702, P1_U3703, P1_U3704, P1_U3705, P1_U3706, P1_U3707, P1_U3708, P1_U3709, P1_U3710, P1_U3711, P1_U3712, P1_U3713, P1_U3714, P1_U3715, P1_U3716, P1_U3717, P1_U3718, P1_U3719, P1_U3720, P1_U3721, P1_U3722, P1_U3723, P1_U3724, P1_U3725, P1_U3726, P1_U3727, P1_U3728, P1_U3729, P1_U3730, P1_U3731, P1_U3732, P1_U3733, P1_U3734, P1_U3735, P1_U3736, P1_U3737, P1_U3738, P1_U3739, P1_U3740, P1_U3741, P1_U3742, P1_U3743, P1_U3744, P1_U3745, P1_U3746, P1_U3747, P1_U3748, P1_U3749, P1_U3750, P1_U3751, P1_U3752, P1_U3753, P1_U3754, P1_U3755, P1_U3756, P1_U3757, P1_U3758, P1_U3759, P1_U3760, P1_U3761, P1_U3762, P1_U3763, P1_U3764, P1_U3765, P1_U3766, P1_U3767, P1_U3768, P1_U3769, P1_U3770, P1_U3771, P1_U3772, P1_U3773, P1_U3774, P1_U3775, P1_U3776, P1_U3777, P1_U3778, P1_U3779, P1_U3780, P1_U3781, P1_U3782, P1_U3783, P1_U3784, P1_U3785, P1_U3786, P1_U3787, P1_U3788, P1_U3789, P1_U3790, P1_U3791, P1_U3792, P1_U3793, P1_U3794, P1_U3795, P1_U3796, P1_U3797, P1_U3798, P1_U3799, P1_U3800, P1_U3801, P1_U3802, P1_U3803, P1_U3804, P1_U3805, P1_U3806, P1_U3807, P1_U3808, P1_U3809, P1_U3810, P1_U3811, P1_U3812, P1_U3813, P1_U3814, P1_U3815, P1_U3816, P1_U3817, P1_U3818, P1_U3819, P1_U3820, P1_U3821, P1_U3822, P1_U3823, P1_U3824, P1_U3825, P1_U3826, P1_U3827, P1_U3828, P1_U3829, P1_U3830, P1_U3831, P1_U3832, P1_U3833, P1_U3834, P1_U3835, P1_U3836, P1_U3837, P1_U3838, P1_U3839, P1_U3840, P1_U3841, P1_U3842, P1_U3843, P1_U3844, P1_U3845, P1_U3846, P1_U3847, P1_U3848, P1_U3849, P1_U3850, P1_U3851, P1_U3852, P1_U3853, P1_U3854, P1_U3855, P1_U3856, P1_U3857, P1_U3858, P1_U3859, P1_U3860, P1_U3861, P1_U3862, P1_U3863, P1_U3864, P1_U3865, P1_U3866, P1_U3867, P1_U3868, P1_U3869, P1_U3870, P1_U3871, P1_U3872, P1_U3873, P1_U3874, P1_U3875, P1_U3876, P1_U3877, P1_U3878, P1_U3879, P1_U3880, P1_U3881, P1_U3882, P1_U3883, P1_U3884, P1_U3885, P1_U3886, P1_U3887, P1_U3888, P1_U3889, P1_U3890, P1_U3891, P1_U3892, P1_U3893, P1_U3894, P1_U3895, P1_U3896, P1_U3897, P1_U3898, P1_U3899, P1_U3900, P1_U3901, P1_U3902, P1_U3903, P1_U3904, P1_U3905, P1_U3906, P1_U3907, P1_U3908, P1_U3909, P1_U3910, P1_U3911, P1_U3912, P1_U3913, P1_U3914, P1_U3915, P1_U3916, P1_U3917, P1_U3918, P1_U3919, P1_U3920, P1_U3921, P1_U3922, P1_U3923, P1_U3924, P1_U3925, P1_U3926, P1_U3927, P1_U3928, P1_U3929, P1_U3930, P1_U3931, P1_U3932, P1_U3933, P1_U3934, P1_U3935, P1_U3936, P1_U3937, P1_U3938, P1_U3939, P1_U3940, P1_U3941, P1_U3942, P1_U3943, P1_U3944, P1_U3945, P1_U3946, P1_U3947, P1_U3948, P1_U3949, P1_U3950, P1_U3951, P1_U3952, P1_U3953, P1_U3954, P1_U3955, P1_U3956, P1_U3957, P1_U3958, P1_U3959, P1_U3960, P1_U3961, P1_U3962, P1_U3963, P1_U3964, P1_U3965, P1_U3966, P1_U3967, P1_U3968, P1_U3969, P1_U3970, P1_U3971, P1_U3972, P1_U3974, P1_U3975, P1_U3976, P1_U3977, P1_U3978, P1_U3979, P1_U3980, P1_U3981, P1_U3982, P1_U3983, P1_U3984, P1_U3985, P1_U3986, P1_U3987, P1_U3988, P1_U3989, P1_U3990, P1_U3991, P1_U3992, P1_U3993, P1_U3994, P1_U3995, P1_U3996, P1_U3997, P1_U3998, P1_U3999, P1_U4000, P1_U4001, P1_U4002, P1_U4003, P1_U4004, P1_U4005, P1_U4006, P1_U4007, P1_U4008, P1_U4009, P1_U4010, P1_U4011, P1_U4012, P1_U4013, P1_U4014, P1_U4015, P1_U4016, P1_U4017, P1_U4018, P1_U4019, P1_U4020, P1_U4021, P1_U4022, P1_U4023, P1_U4024, P1_U4025, P1_U4026, P1_U4027, P1_U4028, P1_U4029, P1_U4030, P1_U4031, P1_U4032, P1_U4033, P1_U4034, P1_U4035, P1_U4036, P1_U4037, P1_U4038, P1_U4039, P1_U4040, P1_U4041, P1_U4042, P1_U4043, P1_U4044, P1_U4045, P1_U4046, P1_U4047, P1_U4048, P1_U4049, P1_U4050, P1_U4051, P1_U4052, P1_U4053, P1_U4054, P1_U4055, P1_U4056, P1_U4057, P1_U4058, P1_U4059, P1_U4060, P1_U4061, P1_U4062, P1_U4063, P1_U4064, P1_U4065, P1_U4066, P1_U4067, P1_U4068, P1_U4069, P1_U4070, P1_U4071, P1_U4072, P1_U4073, P1_U4074, P1_U4075, P1_U4076, P1_U4077, P1_U4078, P1_U4079, P1_U4080, P1_U4081, P1_U4082, P1_U4083, P1_U4084, P1_U4085, P1_U4086, P1_U4087, P1_U4088, P1_U4089, P1_U4090, P1_U4091, P1_U4092, P1_U4093, P1_U4094, P1_U4095, P1_U4096, P1_U4097, P1_U4098, P1_U4099, P1_U4100, P1_U4101, P1_U4102, P1_U4103, P1_U4104, P1_U4105, P1_U4106, P1_U4107, P1_U4108, P1_U4109, P1_U4110, P1_U4111, P1_U4112, P1_U4113, P1_U4114, P1_U4115, P1_U4116, P1_U4117, P1_U4118, P1_U4119, P1_U4120, P1_U4121, P1_U4122, P1_U4123, P1_U4124, P1_U4125, P1_U4126, P1_U4127, P1_U4128, P1_U4129, P1_U4130, P1_U4131, P1_U4132, P1_U4133, P1_U4134, P1_U4135, P1_U4136, P1_U4137, P1_U4138, P1_U4139, P1_U4140, P1_U4141, P1_U4142, P1_U4143, P1_U4144, P1_U4145, P1_U4146, P1_U4147, P1_U4148, P1_U4149, P1_U4150, P1_U4151, P1_U4152, P1_U4153, P1_U4154, P1_U4155, P1_U4156, P1_U4157, P1_U4158, P1_U4159, P1_U4160, P1_U4161, P1_U4162, P1_U4163, P1_U4164, P1_U4165, P1_U4166, P1_U4167, P1_U4168, P1_U4169, P1_U4170, P1_U4171, P1_U4172, P1_U4173, P1_U4174, P1_U4175, P1_U4176, P1_U4177, P1_U4178, P1_U4179, P1_U4180, P1_U4181, P1_U4182, P1_U4183, P1_U4184, P1_U4185, P1_U4186, P1_U4187, P1_U4188, P1_U4189, P1_U4190, P1_U4191, P1_U4192, P1_U4193, P1_U4194, P1_U4195, P1_U4196, P1_U4197, P1_U4198, P1_U4199, P1_U4200, P1_U4201, P1_U4202, P1_U4203, P1_U4204, P1_U4205, P1_U4206, P1_U4207, P1_U4208, P1_U4209, P1_U4210, P1_U4211, P1_U4212, P1_U4213, P1_U4214, P1_U4215, P1_U4216, P1_U4217, P1_U4218, P1_U4219, P1_U4220, P1_U4221, P1_U4222, P1_U4223, P1_U4224, P1_U4225, P1_U4226, P1_U4227, P1_U4228, P1_U4229, P1_U4230, P1_U4231, P1_U4232, P1_U4233, P1_U4234, P1_U4235, P1_U4236, P1_U4237, P1_U4238, P1_U4239, P1_U4240, P1_U4241, P1_U4242, P1_U4243, P1_U4244, P1_U4245, P1_U4246, P1_U4247, P1_U4248, P1_U4249, P1_U4250, P1_U4251, P1_U4252, P1_U4253, P1_U4254, P1_U4255, P1_U4256, P1_U4257, P1_U4258, P1_U4259, P1_U4260, P1_U4261, P1_U4262, P1_U4263, P1_U4264, P1_U4265, P1_U4266, P1_U4267, P1_U4268, P1_U4269, P1_U4270, P1_U4271, P1_U4272, P1_U4273, P1_U4274, P1_U4275, P1_U4276, P1_U4277, P1_U4278, P1_U4279, P1_U4280, P1_U4281, P1_U4282, P1_U4283, P1_U4284, P1_U4285, P1_U4286, P1_U4287, P1_U4288, P1_U4289, P1_U4290, P1_U4291, P1_U4292, P1_U4293, P1_U4294, P1_U4295, P1_U4296, P1_U4297, P1_U4298, P1_U4299, P1_U4300, P1_U4301, P1_U4302, P1_U4303, P1_U4304, P1_U4305, P1_U4306, P1_U4307, P1_U4308, P1_U4309, P1_U4310, P1_U4311, P1_U4312, P1_U4313, P1_U4314, P1_U4315, P1_U4316, P1_U4317, P1_U4318, P1_U4319, P1_U4320, P1_U4321, P1_U4322, P1_U4323, P1_U4324, P1_U4325, P1_U4326, P1_U4327, P1_U4328, P1_U4329, P1_U4330, P1_U4331, P1_U4332, P1_U4333, P1_U4334, P1_U4335, P1_U4336, P1_U4337, P1_U4338, P1_U4339, P1_U4340, P1_U4341, P1_U4342, P1_U4343, P1_U4344, P1_U4345, P1_U4346, P1_U4347, P1_U4348, P1_U4349, P1_U4350, P1_U4351, P1_U4352, P1_U4353, P1_U4354, P1_U4355, P1_U4356, P1_U4357, P1_U4358, P1_U4359, P1_U4360, P1_U4361, P1_U4362, P1_U4363, P1_U4364, P1_U4365, P1_U4366, P1_U4367, P1_U4368, P1_U4369, P1_U4370, P1_U4371, P1_U4372, P1_U4373, P1_U4374, P1_U4375, P1_U4376, P1_U4377, P1_U4378, P1_U4379, P1_U4380, P1_U4381, P1_U4382, P1_U4383, P1_U4384, P1_U4385, P1_U4386, P1_U4387, P1_U4388, P1_U4389, P1_U4390, P1_U4391, P1_U4392, P1_U4393, P1_U4394, P1_U4395, P1_U4396, P1_U4397, P1_U4398, P1_U4399, P1_U4400, P1_U4401, P1_U4402, P1_U4403, P1_U4404, P1_U4405, P1_U4406, P1_U4407, P1_U4408, P1_U4409, P1_U4410, P1_U4411, P1_U4412, P1_U4413, P1_U4414, P1_U4415, P1_U4416, P1_U4417, P1_U4418, P1_U4419, P1_U4420, P1_U4421, P1_U4422, P1_U4423, P1_U4424, P1_U4425, P1_U4426, P1_U4427, P1_U4428, P1_U4429, P1_U4430, P1_U4431, P1_U4432, P1_U4433, P1_U4434, P1_U4435, P1_U4436, P1_U4437, P1_U4438, P1_U4439, P1_U4440, P1_U4441, P1_U4442, P1_U4443, P1_U4444, P1_U4445, P1_U4446, P1_U4447, P1_U4448, P1_U4449, P1_U4450, P1_U4451, P1_U4452, P1_U4453, P1_U4454, P1_U4455, P1_U4456, P1_U4457, P1_U4458, P1_U4459, P1_U4460, P1_U4461, P1_U4462, P1_U4463, P1_U4464, P1_U4465, P1_U4466, P1_U4467, P1_U4468, P1_U4469, P1_U4470, P1_U4471, P1_U4472, P1_U4473, P1_U4474, P1_U4475, P1_U4476, P1_U4477, P1_U4478, P1_U4479, P1_U4480, P1_U4481, P1_U4482, P1_U4483, P1_U4484, P1_U4485, P1_U4486, P1_U4487, P1_U4488, P1_U4489, P1_U4490, P1_U4491, P1_U4492, P1_U4493, P1_U4494, P1_U4495, P1_U4496, P1_U4497, P1_U4498, P1_U4499, P1_U4500, P1_U4501, P1_U4502, P1_U4503, P1_U4504, P1_U4505, P1_U4506, P1_U4507, P1_U4508, P1_U4509, P1_U4510, P1_U4511, P1_U4512, P1_U4513, P1_U4514, P1_U4515, P1_U4516, P1_U4517, P1_U4518, P1_U4519, P1_U4520, P1_U4521, P1_U4522, P1_U4523, P1_U4524, P1_U4525, P1_U4526, P1_U4527, P1_U4528, P1_U4529, P1_U4530, P1_U4531, P1_U4532, P1_U4533, P1_U4534, P1_U4535, P1_U4536, P1_U4537, P1_U4538, P1_U4539, P1_U4540, P1_U4541, P1_U4542, P1_U4543, P1_U4544, P1_U4545, P1_U4546, P1_U4547, P1_U4548, P1_U4549, P1_U4550, P1_U4551, P1_U4552, P1_U4553, P1_U4554, P1_U4555, P1_U4556, P1_U4557, P1_U4558, P1_U4559, P1_U4560, P1_U4561, P1_U4562, P1_U4563, P1_U4564, P1_U4565, P1_U4566, P1_U4567, P1_U4568, P1_U4569, P1_U4570, P1_U4571, P1_U4572, P1_U4573, P1_U4574, P1_U4575, P1_U4576, P1_U4577, P1_U4578, P1_U4579, P1_U4580, P1_U4581, P1_U4582, P1_U4583, P1_U4584, P1_U4585, P1_U4586, P1_U4587, P1_U4588, P1_U4589, P1_U4590, P1_U4591, P1_U4592, P1_U4593, P1_U4594, P1_U4595, P1_U4596, P1_U4597, P1_U4598, P1_U4599, P1_U4600, P1_U4601, P1_U4602, P1_U4603, P1_U4604, P1_U4605, P1_U4606, P1_U4607, P1_U4608, P1_U4609, P1_U4610, P1_U4611, P1_U4612, P1_U4613, P1_U4614, P1_U4615, P1_U4616, P1_U4617, P1_U4618, P1_U4619, P1_U4620, P1_U4621, P1_U4622, P1_U4623, P1_U4624, P1_U4625, P1_U4626, P1_U4627, P1_U4628, P1_U4629, P1_U4630, P1_U4631, P1_U4632, P1_U4633, P1_U4634, P1_U4635, P1_U4636, P1_U4637, P1_U4638, P1_U4639, P1_U4640, P1_U4641, P1_U4642, P1_U4643, P1_U4644, P1_U4645, P1_U4646, P1_U4647, P1_U4648, P1_U4649, P1_U4650, P1_U4651, P1_U4652, P1_U4653, P1_U4654, P1_U4655, P1_U4656, P1_U4657, P1_U4658, P1_U4659, P1_U4660, P1_U4661, P1_U4662, P1_U4663, P1_U4664, P1_U4665, P1_U4666, P1_U4667, P1_U4668, P1_U4669, P1_U4670, P1_U4671, P1_U4672, P1_U4673, P1_U4674, P1_U4675, P1_U4676, P1_U4677, P1_U4678, P1_U4679, P1_U4680, P1_U4681, P1_U4682, P1_U4683, P1_U4684, P1_U4685, P1_U4686, P1_U4687, P1_U4688, P1_U4689, P1_U4690, P1_U4691, P1_U4692, P1_U4693, P1_U4694, P1_U4695, P1_U4696, P1_U4697, P1_U4698, P1_U4699, P1_U4700, P1_U4701, P1_U4702, P1_U4703, P1_U4704, P1_U4705, P1_U4706, P1_U4707, P1_U4708, P1_U4709, P1_U4710, P1_U4711, P1_U4712, P1_U4713, P1_U4714, P1_U4715, P1_U4716, P1_U4717, P1_U4718, P1_U4719, P1_U4720, P1_U4721, P1_U4722, P1_U4723, P1_U4724, P1_U4725, P1_U4726, P1_U4727, P1_U4728, P1_U4729, P1_U4730, P1_U4731, P1_U4732, P1_U4733, P1_U4734, P1_U4735, P1_U4736, P1_U4737, P1_U4738, P1_U4739, P1_U4740, P1_U4741, P1_U4742, P1_U4743, P1_U4744, P1_U4745, P1_U4746, P1_U4747, P1_U4748, P1_U4749, P1_U4750, P1_U4751, P1_U4752, P1_U4753, P1_U4754, P1_U4755, P1_U4756, P1_U4757, P1_U4758, P1_U4759, P1_U4760, P1_U4761, P1_U4762, P1_U4763, P1_U4764, P1_U4765, P1_U4766, P1_U4767, P1_U4768, P1_U4769, P1_U4770, P1_U4771, P1_U4772, P1_U4773, P1_U4774, P1_U4775, P1_U4776, P1_U4777, P1_U4778, P1_U4779, P1_U4780, P1_U4781, P1_U4782, P1_U4783, P1_U4784, P1_U4785, P1_U4786, P1_U4787, P1_U4788, P1_U4789, P1_U4790, P1_U4791, P1_U4792, P1_U4793, P1_U4794, P1_U4795, P1_U4796, P1_U4797, P1_U4798, P1_U4799, P1_U4800, P1_U4801, P1_U4802, P1_U4803, P1_U4804, P1_U4805, P1_U4806, P1_U4807, P1_U4808, P1_U4809, P1_U4810, P1_U4811, P1_U4812, P1_U4813, P1_U4814, P1_U4815, P1_U4816, P1_U4817, P1_U4818, P1_U4819, P1_U4820, P1_U4821, P1_U4822, P1_U4823, P1_U4824, P1_U4825, P1_U4826, P1_U4827, P1_U4828, P1_U4829, P1_U4830, P1_U4831, P1_U4832, P1_U4833, P1_U4834, P1_U4835, P1_U4836, P1_U4837, P1_U4838, P1_U4839, P1_U4840, P1_U4841, P1_U4842, P1_U4843, P1_U4844, P1_U4845, P1_U4846, P1_U4847, P1_U4848, P1_U4849, P1_U4850, P1_U4851, P1_U4852, P1_U4853, P1_U4854, P1_U4855, P1_U4856, P1_U4857, P1_U4858, P1_U4859, P1_U4860, P1_U4861, P1_U4862, P1_U4863, P1_U4864, P1_U4865, P1_U4866, P1_U4867, P1_U4868, P1_U4869, P1_U4870, P1_U4871, P1_U4872, P1_U4873, P1_U4874, P1_U4875, P1_U4876, P1_U4877, P1_U4878, P1_U4879, P1_U4880, P1_U4881, P1_U4882, P1_U4883, P1_U4884, P1_U4885, P1_U4886, P1_U4887, P1_U4888, P1_U4889, P1_U4890, P1_U4891, P1_U4892, P1_U4893, P1_U4894, P1_U4895, P1_U4896, P1_U4897, P1_U4898, P1_U4899, P1_U4900, P1_U4901, P1_U4902, P1_U4903, P1_U4904, P1_U4905, P1_U4906, P1_U4907, P1_U4908, P1_U4909, P1_U4910, P1_U4911, P1_U4912, P1_U4913, P1_U4914, P1_U4915, P1_U4916, P1_U4917, P1_U4918, P1_U4919, P1_U4920, P1_U4921, P1_U4922, P1_U4923, P1_U4924, P1_U4925, P1_U4926, P1_U4927, P1_U4928, P1_U4929, P1_U4930, P1_U4931, P1_U4932, P1_U4933, P1_U4934, P1_U4935, P1_U4936, P1_U4937, P1_U4938, P1_U4939, P1_U4940, P1_U4941, P1_U4942, P1_U4943, P1_U4944, P1_U4945, P1_U4946, P1_U4947, P1_U4948, P1_U4949, P1_U4950, P1_U4951, P1_U4952, P1_U4953, P1_U4954, P1_U4955, P1_U4956, P1_U4957, P1_U4958, P1_U4959, P1_U4960, P1_U4961, P1_U4962, P1_U4963, P1_U4964, P1_U4965, P1_U4966, P1_U4967, P1_U4968, P1_U4969, P1_U4970, P1_U4971, P1_U4972, P1_U4973, P1_U4974, P1_U4975, P1_U4976, P1_U4977, P1_U4978, P1_U4979, P1_U4980, P1_U4981, P1_U4982, P1_U4983, P1_U4984, P1_U4985, P1_U4986, P1_U4987, P1_U4988, P1_U4989, P1_U4990, P1_U4991, P1_U4992, P1_U4993, P1_U4994, P1_U4995, P1_U4996, P1_U4997, P1_U4998, P1_U4999, P1_U5000, P1_U5001, P1_U5002, P1_U5003, P1_U5004, P1_U5005, P1_U5006, P1_U5007, P1_U5008, P1_U5009, P1_U5010, P1_U5011, P1_U5012, P1_U5013, P1_U5014, P1_U5015, P1_U5016, P1_U5017, P1_U5018, P1_U5019, P1_U5020, P1_U5021, P1_U5022, P1_U5023, P1_U5024, P1_U5025, P1_U5026, P1_U5027, P1_U5028, P1_U5029, P1_U5030, P1_U5031, P1_U5032, P1_U5033, P1_U5034, P1_U5035, P1_U5036, P1_U5037, P1_U5038, P1_U5039, P1_U5040, P1_U5041, P1_U5042, P1_U5043, P1_U5044, P1_U5045, P1_U5046, P1_U5047, P1_U5048, P1_U5049, P1_U5050, P1_U5051, P1_U5052, P1_U5053, P1_U5054, P1_U5055, P1_U5056, P1_U5057, P1_U5058, P1_U5059, P1_U5060, P1_U5061, P1_U5062, P1_U5063, P1_U5064, P1_U5065, P1_U5066, P1_U5067, P1_U5068, P1_U5069, P1_U5070, P1_U5071, P1_U5072, P1_U5073, P1_U5074, P1_U5075, P1_U5076, P1_U5077, P1_U5078, P1_U5079, P1_U5080, P1_U5081, P1_U5082, P1_U5083, P1_U5084, P1_U5085, P1_U5086, P1_U5087, P1_U5088, P1_U5089, P1_U5090, P1_U5091, P1_U5092, P1_U5093, P1_U5094, P1_U5095, P1_U5096, P1_U5097, P1_U5098, P1_U5099, P1_U5100, P1_U5101, P1_U5102, P1_U5103, P1_U5104, P1_U5105, P1_U5106, P1_U5107, P1_U5108, P1_U5109, P1_U5110, P1_U5111, P1_U5112, P1_U5113, P1_U5114, P1_U5115, P1_U5116, P1_U5117, P1_U5118, P1_U5119, P1_U5120, P1_U5121, P1_U5122, P1_U5123, P1_U5124, P1_U5125, P1_U5126, P1_U5127, P1_U5128, P1_U5129, P1_U5130, P1_U5131, P1_U5132, P1_U5133, P1_U5134, P1_U5135, P1_U5136, P1_U5137, P1_U5138, P1_U5139, P1_U5140, P1_U5141, P1_U5142, P1_U5143, P1_U5144, P1_U5145, P1_U5146, P1_U5147, P1_U5148, P1_U5149, P1_U5150, P1_U5151, P1_U5152, P1_U5153, P1_U5154, P1_U5155, P1_U5156, P1_U5157, P1_U5158, P1_U5159, P1_U5160, P1_U5161, P1_U5162, P1_U5163, P1_U5164, P1_U5165, P1_U5166, P1_U5167, P1_U5168, P1_U5169, P1_U5170, P1_U5171, P1_U5172, P1_U5173, P1_U5174, P1_U5175, P1_U5176, P1_U5177, P1_U5178, P1_U5179, P1_U5180, P1_U5181, P1_U5182, P1_U5183, P1_U5184, P1_U5185, P1_U5186, P1_U5187, P1_U5188, P1_U5189, P1_U5190, P1_U5191, P1_U5192, P1_U5193, P1_U5194, P1_U5195, P1_U5196, P1_U5197, P1_U5198, P1_U5199, P1_U5200, P1_U5201, P1_U5202, P1_U5203, P1_U5204, P1_U5205, P1_U5206, P1_U5207, P1_U5208, P1_U5209, P1_U5210, P1_U5211, P1_U5212, P1_U5213, P1_U5214, P1_U5215, P1_U5216, P1_U5217, P1_U5218, P1_U5219, P1_U5220, P1_U5221, P1_U5222, P1_U5223, P1_U5224, P1_U5225, P1_U5226, P1_U5227, P1_U5228, P1_U5229, P1_U5230, P1_U5231, P1_U5232, P1_U5233, P1_U5234, P1_U5235, P1_U5236, P1_U5237, P1_U5238, P1_U5239, P1_U5240, P1_U5241, P1_U5242, P1_U5243, P1_U5244, P1_U5245, P1_U5246, P1_U5247, P1_U5248, P1_U5249, P1_U5250, P1_U5251, P1_U5252, P1_U5253, P1_U5254, P1_U5255, P1_U5256, P1_U5257, P1_U5258, P1_U5259, P1_U5260, P1_U5261, P1_U5262, P1_U5263, P1_U5264, P1_U5265, P1_U5266, P1_U5267, P1_U5268, P1_U5269, P1_U5270, P1_U5271, P1_U5272, P1_U5273, P1_U5274, P1_U5275, P1_U5276, P1_U5277, P1_U5278, P1_U5279, P1_U5280, P1_U5281, P1_U5282, P1_U5283, P1_U5284, P1_U5285, P1_U5286, P1_U5287, P1_U5288, P1_U5289, P1_U5290, P1_U5291, P1_U5292, P1_U5293, P1_U5294, P1_U5295, P1_U5296, P1_U5297, P1_U5298, P1_U5299, P1_U5300, P1_U5301, P1_U5302, P1_U5303, P1_U5304, P1_U5305, P1_U5306, P1_U5307, P1_U5308, P1_U5309, P1_U5310, P1_U5311, P1_U5312, P1_U5313, P1_U5314, P1_U5315, P1_U5316, P1_U5317, P1_U5318, P1_U5319, P1_U5320, P1_U5321, P1_U5322, P1_U5323, P1_U5324, P1_U5325, P1_U5326, P1_U5327, P1_U5328, P1_U5329, P1_U5330, P1_U5331, P1_U5332, P1_U5333, P1_U5334, P1_U5335, P1_U5336, P1_U5337, P1_U5338, P1_U5339, P1_U5340, P1_U5341, P1_U5342, P1_U5343, P1_U5344, P1_U5345, P1_U5346, P1_U5347, P1_U5348, P1_U5349, P1_U5350, P1_U5351, P1_U5352, P1_U5353, P1_U5354, P1_U5355, P1_U5356, P1_U5357, P1_U5358, P1_U5359, P1_U5360, P1_U5361, P1_U5362, P1_U5363, P1_U5364, P1_U5365, P1_U5366, P1_U5367, P1_U5368, P1_U5369, P1_U5370, P1_U5371, P1_U5372, P1_U5373, P1_U5374, P1_U5375, P1_U5376, P1_U5377, P1_U5378, P1_U5379, P1_U5380, P1_U5381, P1_U5382, P1_U5383, P1_U5384, P1_U5385, P1_U5386, P1_U5387, P1_U5388, P1_U5389, P1_U5390, P1_U5391, P1_U5392, P1_U5393, P1_U5394, P1_U5395, P1_U5396, P1_U5397, P1_U5398, P1_U5399, P1_U5400, P1_U5401, P1_U5402, P1_U5403, P1_U5404, P1_U5405, P1_U5406, P1_U5407, P1_U5408, P1_U5409, P1_U5410, P1_U5411, P1_U5412, P1_U5413, P1_U5414, P1_U5415, P1_U5416, P1_U5417, P1_U5418, P1_U5419, P1_U5420, P1_U5421, P1_U5422, P1_U5423, P1_U5424, P1_U5425, P1_U5426, P1_U5427, P1_U5428, P1_U5429, P1_U5430, P1_U5431, P1_U5432, P1_U5433, P1_U5434, P1_U5435, P1_U5436, P1_U5437, P1_U5438, P1_U5439, P1_U5440, P1_U5441, P1_U5442, P1_U5443, P1_U5444, P1_U5445, P1_U5446, P1_U5447, P1_U5448, P1_U5449, P1_U5450, P1_U5451, P1_U5452, P1_U5453, P1_U5454, P1_U5455, P1_U5456, P1_U5457, P1_U5458, P1_U5459, P1_U5460, P1_U5461, P1_U5462, P1_U5463, P1_U5464, P1_U5465, P1_U5466, P1_U5467, P1_U5468, P1_U5469, P1_U5470, P1_U5471, P1_U5472, P1_U5473, P1_U5474, P1_U5475, P1_U5476, P1_U5477, P1_U5478, P1_U5479, P1_U5480, P1_U5481, P1_U5482, P1_U5483, P1_U5484, P1_U5485, P1_U5486, P1_U5487, P1_U5488, P1_U5489, P1_U5490, P1_U5491, P1_U5492, P1_U5493, P1_U5494, P1_U5495, P1_U5496, P1_U5497, P1_U5498, P1_U5499, P1_U5500, P1_U5501, P1_U5502, P1_U5503, P1_U5504, P1_U5505, P1_U5506, P1_U5507, P1_U5508, P1_U5509, P1_U5510, P1_U5511, P1_U5512, P1_U5513, P1_U5514, P1_U5515, P1_U5516, P1_U5517, P1_U5518, P1_U5519, P1_U5520, P1_U5521, P1_U5522, P1_U5523, P1_U5524, P1_U5525, P1_U5526, P1_U5527, P1_U5528, P1_U5529, P1_U5530, P1_U5531, P1_U5532, P1_U5533, P1_U5534, P1_U5535, P1_U5536, P1_U5537, P1_U5538, P1_U5539, P1_U5540, P1_U5541, P1_U5542, P1_U5543, P1_U5544, P1_U5545, P1_U5546, P1_U5547, P1_U5548, P1_U5549, P1_U5550, P1_U5551, P1_U5552, P1_U5553, P1_U5554, P1_U5555, P1_U5556, P1_U5557, P1_U5558, P1_U5559, P1_U5560, P1_U5561, P1_U5562, P1_U5563, P1_U5564, P1_U5565, P1_U5566, P1_U5567, P1_U5568, P1_U5569, P1_U5570, P1_U5571, P1_U5572, P1_U5573, P1_U5574, P1_U5575, P1_U5576, P1_U5577, P1_U5578, P1_U5579, P1_U5580, P1_U5581, P1_U5582, P1_U5583, P1_U5584, P1_U5585, P1_U5586, P1_U5587, P1_U5588, P1_U5589, P1_U5590, P1_U5591, P1_U5592, P1_U5593, P1_U5594, P1_U5595, P1_U5596, P1_U5597, P1_U5598, P1_U5599, P1_U5600, P1_U5601, P1_U5602, P1_U5603, P1_U5604, P1_U5605, P1_U5606, P1_U5607, P1_U5608, P1_U5609, P1_U5610, P1_U5611, P1_U5612, P1_U5613, P1_U5614, P1_U5615, P1_U5616, P1_U5617, P1_U5618, P1_U5619, P1_U5620, P1_U5621, P1_U5622, P1_U5623, P1_U5624, P1_U5625, P1_U5626, P1_U5627, P1_U5628, P1_U5629, P1_U5630, P1_U5631, P1_U5632, P1_U5633, P1_U5634, P1_U5635, P1_U5636, P1_U5637, P1_U5638, P1_U5639, P1_U5640, P1_U5641, P1_U5642, P1_U5643, P1_U5644, P1_U5645, P1_U5646, P1_U5647, P1_U5648, P1_U5649, P1_U5650, P1_U5651, P1_U5652, P1_U5653, P1_U5654, P1_U5655, P1_U5656, P1_U5657, P1_U5658, P1_U5659, P1_U5660, P1_U5661, P1_U5662, P1_U5663, P1_U5664, P1_U5665, P1_U5666, P1_U5667, P1_U5668, P1_U5669, P1_U5670, P1_U5671, P1_U5672, P1_U5673, P1_U5674, P1_U5675, P1_U5676, P1_U5677, P1_U5678, P1_U5679, P1_U5680, P1_U5681, P1_U5682, P1_U5683, P1_U5684, P1_U5685, P1_U5686, P1_U5687, P1_U5688, P1_U5689, P1_U5690, P1_U5691, P1_U5692, P1_U5693, P1_U5694, P1_U5695, P1_U5696, P1_U5697, P1_U5698, P1_U5699, P1_U5700, P1_U5701, P1_U5702, P1_U5703, P1_U5704, P1_U5705, P1_U5706, P1_U5707, P1_U5708, P1_U5709, P1_U5710, P1_U5711, P1_U5712, P1_U5713, P1_U5714, P1_U5715, P1_U5716, P1_U5717, P1_U5718, P1_U5719, P1_U5720, P1_U5721, P1_U5722, P1_U5723, P1_U5724, P1_U5725, P1_U5726, P1_U5727, P1_U5728, P1_U5729, P1_U5730, P1_U5731, P1_U5732, P1_U5733, P1_U5734, P1_U5735, P1_U5736, P1_U5737, P1_U5738, P1_U5739, P1_U5740, P1_U5741, P1_U5742, P1_U5743, P1_U5744, P1_U5745, P1_U5746, P1_U5747, P1_U5748, P1_U5749, P1_U5750, P1_U5751, P1_U5752, P1_U5753, P1_U5754, P1_U5755, P1_U5756, P1_U5757, P1_U5758, P1_U5759, P1_U5760, P1_U5761, P1_U5762, P1_U5763, P1_U5764, P1_U5765, P1_U5766, P1_U5767, P1_U5768, P1_U5769, P1_U5770, P1_U5771, P1_U5772, P1_U5773, P1_U5774, P1_U5775, P1_U5776, P1_U5777, P1_U5778, P1_U5779, P1_U5780, P1_U5781, P1_U5782, P1_U5783, P1_U5784, P1_U5785, P1_U5786, P1_U5787, P1_U5788, P1_U5789, P1_U5790, P1_U5791, P1_U5792, P1_U5793, P1_U5794, P1_U5795, P1_U5796, P1_U5797, P1_U5798, P1_U5799, P1_U5800, P1_U5801, P1_U5802, P1_U5803, P1_U5804, P1_U5805, P1_U5806, P1_U5807, P1_U5808, P1_U5809, P1_U5810, P1_U5811, P1_U5812, P1_U5813, P1_U5814, P1_U5815, P1_U5816, P1_U5817, P1_U5818, P1_U5819, P1_U5820, P1_U5821, P1_U5822, P1_U5823, P1_U5824, P1_U5825, P1_U5826, P1_U5827, P1_U5828, P1_U5829, P1_U5830, P1_U5831, P1_U5832, P1_U5833, P1_U5834, P1_U5835, P1_U5836, P1_U5837, P1_U5838, P1_U5839, P1_U5840, P1_U5841, P1_U5842, P1_U5843, P1_U5844, P1_U5845, P1_U5846, P1_U5847, P1_U5848, P1_U5849, P1_U5850, P1_U5851, P1_U5852, P1_U5853, P1_U5854, P1_U5855, P1_U5856, P1_U5857, P1_U5858, P1_U5859, P1_U5860, P1_U5861, P1_U5862, P1_U5863, P1_U5864, P1_U5865, P1_U5866, P1_U5867, P1_U5868, P1_U5869, P1_U5870, P1_U5871, P1_U5872, P1_U5873, P1_U5874, P1_U5875, P1_U5876, P1_U5877, P1_U5878, P1_U5879, P1_U5880, P1_U5881, P1_U5882, P1_U5883, P1_U5884, P1_U5885, P1_U5886, P1_U5887, P1_U5888, P1_U5889, P1_U5890, P1_U5891, P1_U5892, P1_U5893, P1_U5894, P1_U5895, P1_U5896, P1_U5897, P1_U5898, P1_U5899, P1_U5900, P1_U5901, P1_U5902, P1_U5903, P1_U5904, P1_U5905, P1_U5906, P1_U5907, P1_U5908, P1_U5909, P1_U5910, P1_U5911, P1_U5912, P1_U5913, P1_U5914, P1_U5915, P1_U5916, P1_U5917, P1_U5918, P1_U5919, P1_U5920, P1_U5921, P1_U5922, P1_U5923, P1_U5924, P1_U5925, P1_U5926, P1_U5927, P1_U5928, P1_U5929, P1_U5930, P1_U5931, P1_U5932, P1_U5933, P1_U5934, P1_U5935, P1_U5936, P1_U5937, P1_U5938, P1_U5939, P1_U5940, P1_U5941, P1_U5942, P1_U5943, P1_U5944, P1_U5945, P1_U5946, P1_U5947, P1_U5948, P1_U5949, P1_U5950, P1_U5951, P1_U5952, P1_U5953, P1_U5954, P1_U5955, P1_U5956, P1_U5957, P1_U5958, P1_U5959, P1_U5960, P1_U5961, P1_U5962, P1_U5963, P1_U5964, P1_U5965, P1_U5966, P1_U5967, P1_U5968, P1_U5969, P1_U5970, P1_U5971, P1_U5972, P1_U5973, P1_U5974, P1_U5975, P1_U5976, P1_U5977, P1_U5978, P1_U5979, P1_U5980, P1_U5981, P1_U5982, P1_U5983, P1_U5984, P1_U5985, P1_U5986, P1_U5987, P1_U5988, P1_U5989, P1_U5990, P1_U5991, P1_U5992, P1_U5993, P1_U5994, P1_U5995, P1_U5996, P1_U5997, P1_U5998, P1_U5999, P1_U6000, P1_U6001, P1_U6002, P1_U6003, P1_U6004, P1_U6005, P1_U6006, P1_U6007, P1_U6008, P1_U6009, P1_U6010, P1_U6011, P1_U6012, P1_U6013, P1_U6014, P1_U6015, P1_U6016, P1_U6017, P1_U6018, P1_U6019, P1_U6020, P1_U6021, P1_U6022, P1_U6023, P1_U6024, P1_U6025, P1_U6026, P1_U6027, P1_U6028, P1_U6029, P1_U6030, P1_U6031, P1_U6032, P1_U6033, P1_U6034, P1_U6035, P1_U6036, P1_U6037, P1_U6038, P1_U6039, P1_U6040, P1_U6041, P1_U6042, P1_U6043, P1_U6044, P1_U6045, P1_U6046, P1_U6047, P1_U6048, P1_U6049, P1_U6050, P1_U6051, P1_U6052, P1_U6053, P1_U6054, P1_U6055, P1_U6056, P1_U6057, P1_U6058, P1_U6059, P1_U6060, P1_U6061, P1_U6062, P1_U6063, P1_U6064, P1_U6065, P1_U6066, P1_U6067, P1_U6068, P1_U6069, P1_U6070, P1_U6071, P1_U6072, P1_U6073, P1_U6074, P1_U6075, P1_U6076, P1_U6077, P1_U6078, P1_U6079, P1_U6080, P1_U6081, P1_U6082, P1_U6083, P1_U6084, P1_U6085, P1_U6086, P1_U6087, P1_U6088, P1_U6089, P1_U6090, P1_U6091, P1_U6092, P1_U6093, P1_U6094, P1_U6095, P1_U6096, P1_U6097, P1_U6098, P1_U6099, P1_U6100, P1_U6101, P1_U6102, P1_U6103, P1_U6104, P1_U6105, P1_U6106, P1_U6107, P1_U6108, P1_U6109, P1_U6110, P1_U6111, P1_U6112, P1_U6113, P1_U6114, P1_U6115, P1_U6116, P1_U6117, P1_U6118, P1_U6119, P1_U6120, P1_U6121, P1_U6122, P1_U6123, P1_U6124, P1_U6125, P1_U6126, P1_U6127, P1_U6128, P1_U6129, P1_U6130, P1_U6131, P1_U6132, P1_U6133, P1_U6134, P1_U6135, P1_U6136, P1_U6137, P1_U6138, P1_U6139, P1_U6140, P1_U6141, P1_U6142, P1_U6143, P1_U6144, P1_U6145, P1_U6146, P1_U6147, P1_U6148, P1_U6149, P1_U6150, P1_U6151, P1_U6152, P1_U6153, P1_U6154, P1_U6155, P1_U6156, P1_U6157, P1_U6158, P1_U6159, P1_U6160, P1_U6161, P1_U6162, P1_U6163, P1_U6164, P1_U6165, P1_U6166, P1_U6167, P1_U6168, P1_U6169, P1_U6170, P1_U6171, P1_U6172, P1_U6173, P1_U6174, P1_U6175, P1_U6176, P1_U6177, P1_U6178, P1_U6179, P1_U6180, P1_U6181, P1_U6182, P1_U6183, P1_U6184, P1_U6185, P1_U6186, P1_U6187, P1_U6188, P1_U6189, P1_U6190, P1_U6191, P1_U6192, P1_U6193, P1_U6194, P1_U6195, P1_U6196, P1_U6197, P1_U6198, P1_U6199, P1_U6200, P1_U6201, P1_U6202, P1_U6203, P1_U6204, P1_U6205, P1_U6206, P1_U6207, P1_U6208, P1_U6209, P1_U6210, P1_U6211, P1_U6212, P1_U6213, P1_U6214, P1_U6215, P1_U6216, P1_U6217, P1_U6218, P1_U6219, P1_U6220, P1_U6221, P1_U6222, P1_U6223, P1_U6224, P1_U6225, P1_U6226, P1_U6227, P1_U6228, P1_U6229, P1_U6230, P1_U6231, P1_U6232, P1_U6233, P1_U6234, P1_U6235, P1_U6236, P2_R1054_U10, P2_R1054_U100, P2_R1054_U101, P2_R1054_U102, P2_R1054_U103, P2_R1054_U104, P2_R1054_U105, P2_R1054_U106, P2_R1054_U107, P2_R1054_U108, P2_R1054_U109, P2_R1054_U11, P2_R1054_U110, P2_R1054_U111, P2_R1054_U112, P2_R1054_U113, P2_R1054_U114, P2_R1054_U115, P2_R1054_U116, P2_R1054_U117, P2_R1054_U118, P2_R1054_U119, P2_R1054_U12, P2_R1054_U120, P2_R1054_U121, P2_R1054_U122, P2_R1054_U123, P2_R1054_U124, P2_R1054_U125, P2_R1054_U126, P2_R1054_U127, P2_R1054_U128, P2_R1054_U129, P2_R1054_U13, P2_R1054_U130, P2_R1054_U131, P2_R1054_U132, P2_R1054_U133, P2_R1054_U134, P2_R1054_U135, P2_R1054_U136, P2_R1054_U137, P2_R1054_U138, P2_R1054_U139, P2_R1054_U14, P2_R1054_U140, P2_R1054_U141, P2_R1054_U142, P2_R1054_U143, P2_R1054_U144, P2_R1054_U145, P2_R1054_U146, P2_R1054_U147, P2_R1054_U148, P2_R1054_U149, P2_R1054_U15, P2_R1054_U150, P2_R1054_U151, P2_R1054_U152, P2_R1054_U153, P2_R1054_U154, P2_R1054_U155, P2_R1054_U156, P2_R1054_U157, P2_R1054_U158, P2_R1054_U159, P2_R1054_U16, P2_R1054_U160, P2_R1054_U161, P2_R1054_U162, P2_R1054_U163, P2_R1054_U164, P2_R1054_U165, P2_R1054_U166, P2_R1054_U167, P2_R1054_U168, P2_R1054_U169, P2_R1054_U17, P2_R1054_U170, P2_R1054_U171, P2_R1054_U172, P2_R1054_U173, P2_R1054_U174, P2_R1054_U175, P2_R1054_U176, P2_R1054_U177, P2_R1054_U178, P2_R1054_U179, P2_R1054_U18, P2_R1054_U180, P2_R1054_U181, P2_R1054_U182, P2_R1054_U183, P2_R1054_U184, P2_R1054_U185, P2_R1054_U186, P2_R1054_U187, P2_R1054_U188, P2_R1054_U189, P2_R1054_U19, P2_R1054_U190, P2_R1054_U191, P2_R1054_U192, P2_R1054_U193, P2_R1054_U194, P2_R1054_U195, P2_R1054_U196, P2_R1054_U197, P2_R1054_U198, P2_R1054_U199, P2_R1054_U20, P2_R1054_U200, P2_R1054_U201, P2_R1054_U202, P2_R1054_U203, P2_R1054_U204, P2_R1054_U205, P2_R1054_U206, P2_R1054_U207, P2_R1054_U208, P2_R1054_U209, P2_R1054_U21, P2_R1054_U210, P2_R1054_U211, P2_R1054_U212, P2_R1054_U213, P2_R1054_U214, P2_R1054_U215, P2_R1054_U216, P2_R1054_U217, P2_R1054_U218, P2_R1054_U219, P2_R1054_U22, P2_R1054_U220, P2_R1054_U221, P2_R1054_U222, P2_R1054_U223, P2_R1054_U224, P2_R1054_U225, P2_R1054_U226, P2_R1054_U227, P2_R1054_U228, P2_R1054_U229, P2_R1054_U23, P2_R1054_U230, P2_R1054_U231, P2_R1054_U232, P2_R1054_U233, P2_R1054_U234, P2_R1054_U235, P2_R1054_U236, P2_R1054_U237, P2_R1054_U238, P2_R1054_U239, P2_R1054_U24, P2_R1054_U240, P2_R1054_U241, P2_R1054_U242, P2_R1054_U243, P2_R1054_U244, P2_R1054_U245, P2_R1054_U246, P2_R1054_U247, P2_R1054_U248, P2_R1054_U249, P2_R1054_U25, P2_R1054_U250, P2_R1054_U251, P2_R1054_U252, P2_R1054_U253, P2_R1054_U254, P2_R1054_U255, P2_R1054_U256, P2_R1054_U257, P2_R1054_U258, P2_R1054_U259, P2_R1054_U26, P2_R1054_U260, P2_R1054_U261, P2_R1054_U262, P2_R1054_U263, P2_R1054_U264, P2_R1054_U265, P2_R1054_U266, P2_R1054_U267, P2_R1054_U268, P2_R1054_U269, P2_R1054_U27, P2_R1054_U270, P2_R1054_U271, P2_R1054_U272, P2_R1054_U273, P2_R1054_U274, P2_R1054_U275, P2_R1054_U276, P2_R1054_U277, P2_R1054_U278, P2_R1054_U279, P2_R1054_U28, P2_R1054_U280, P2_R1054_U281, P2_R1054_U282, P2_R1054_U283, P2_R1054_U284, P2_R1054_U285, P2_R1054_U286, P2_R1054_U287, P2_R1054_U288, P2_R1054_U289, P2_R1054_U29, P2_R1054_U290, P2_R1054_U291, P2_R1054_U292, P2_R1054_U293, P2_R1054_U294, P2_R1054_U30, P2_R1054_U31, P2_R1054_U32, P2_R1054_U33, P2_R1054_U34, P2_R1054_U35, P2_R1054_U36, P2_R1054_U37, P2_R1054_U38, P2_R1054_U39, P2_R1054_U40, P2_R1054_U41, P2_R1054_U42, P2_R1054_U43, P2_R1054_U44, P2_R1054_U45, P2_R1054_U46, P2_R1054_U47, P2_R1054_U48, P2_R1054_U49, P2_R1054_U50, P2_R1054_U51, P2_R1054_U52, P2_R1054_U53, P2_R1054_U54, P2_R1054_U55, P2_R1054_U56, P2_R1054_U57, P2_R1054_U58, P2_R1054_U59, P2_R1054_U6, P2_R1054_U60, P2_R1054_U61, P2_R1054_U62, P2_R1054_U63, P2_R1054_U64, P2_R1054_U65, P2_R1054_U66, P2_R1054_U67, P2_R1054_U68, P2_R1054_U69, P2_R1054_U7, P2_R1054_U70, P2_R1054_U71, P2_R1054_U72, P2_R1054_U73, P2_R1054_U74, P2_R1054_U75, P2_R1054_U76, P2_R1054_U77, P2_R1054_U78, P2_R1054_U79, P2_R1054_U8, P2_R1054_U80, P2_R1054_U81, P2_R1054_U82, P2_R1054_U83, P2_R1054_U84, P2_R1054_U85, P2_R1054_U86, P2_R1054_U87, P2_R1054_U88, P2_R1054_U89, P2_R1054_U9, P2_R1054_U90, P2_R1054_U91, P2_R1054_U92, P2_R1054_U93, P2_R1054_U94, P2_R1054_U95, P2_R1054_U96, P2_R1054_U97, P2_R1054_U98, P2_R1054_U99, P2_R1077_U10, P2_R1077_U100, P2_R1077_U101, P2_R1077_U102, P2_R1077_U103, P2_R1077_U104, P2_R1077_U105, P2_R1077_U106, P2_R1077_U107, P2_R1077_U108, P2_R1077_U109, P2_R1077_U11, P2_R1077_U110, P2_R1077_U111, P2_R1077_U112, P2_R1077_U113, P2_R1077_U114, P2_R1077_U115, P2_R1077_U116, P2_R1077_U117, P2_R1077_U118, P2_R1077_U119, P2_R1077_U12, P2_R1077_U120, P2_R1077_U121, P2_R1077_U122, P2_R1077_U123, P2_R1077_U124, P2_R1077_U125, P2_R1077_U126, P2_R1077_U127, P2_R1077_U128, P2_R1077_U129, P2_R1077_U13, P2_R1077_U130, P2_R1077_U131, P2_R1077_U132, P2_R1077_U133, P2_R1077_U134, P2_R1077_U135, P2_R1077_U136, P2_R1077_U137, P2_R1077_U138, P2_R1077_U139, P2_R1077_U14, P2_R1077_U140, P2_R1077_U141, P2_R1077_U142, P2_R1077_U143, P2_R1077_U144, P2_R1077_U145, P2_R1077_U146, P2_R1077_U147, P2_R1077_U148, P2_R1077_U149, P2_R1077_U15, P2_R1077_U150, P2_R1077_U151, P2_R1077_U152, P2_R1077_U153, P2_R1077_U154, P2_R1077_U155, P2_R1077_U156, P2_R1077_U157, P2_R1077_U158, P2_R1077_U159, P2_R1077_U16, P2_R1077_U160, P2_R1077_U161, P2_R1077_U162, P2_R1077_U163, P2_R1077_U164, P2_R1077_U165, P2_R1077_U166, P2_R1077_U167, P2_R1077_U168, P2_R1077_U169, P2_R1077_U17, P2_R1077_U170, P2_R1077_U171, P2_R1077_U172, P2_R1077_U173, P2_R1077_U174, P2_R1077_U175, P2_R1077_U176, P2_R1077_U177, P2_R1077_U178, P2_R1077_U179, P2_R1077_U18, P2_R1077_U180, P2_R1077_U181, P2_R1077_U182, P2_R1077_U183, P2_R1077_U184, P2_R1077_U185, P2_R1077_U186, P2_R1077_U187, P2_R1077_U188, P2_R1077_U189, P2_R1077_U19, P2_R1077_U190, P2_R1077_U191, P2_R1077_U192, P2_R1077_U193, P2_R1077_U194, P2_R1077_U195, P2_R1077_U196, P2_R1077_U197, P2_R1077_U198, P2_R1077_U199, P2_R1077_U20, P2_R1077_U200, P2_R1077_U201, P2_R1077_U202, P2_R1077_U203, P2_R1077_U204, P2_R1077_U205, P2_R1077_U206, P2_R1077_U207, P2_R1077_U208, P2_R1077_U209, P2_R1077_U21, P2_R1077_U210, P2_R1077_U211, P2_R1077_U212, P2_R1077_U213, P2_R1077_U214, P2_R1077_U215, P2_R1077_U216, P2_R1077_U217, P2_R1077_U218, P2_R1077_U219, P2_R1077_U22, P2_R1077_U220, P2_R1077_U221, P2_R1077_U222, P2_R1077_U223, P2_R1077_U224, P2_R1077_U225, P2_R1077_U226, P2_R1077_U227, P2_R1077_U228, P2_R1077_U229, P2_R1077_U23, P2_R1077_U230, P2_R1077_U231, P2_R1077_U232, P2_R1077_U233, P2_R1077_U234, P2_R1077_U235, P2_R1077_U236, P2_R1077_U237, P2_R1077_U238, P2_R1077_U239, P2_R1077_U24, P2_R1077_U240, P2_R1077_U241, P2_R1077_U242, P2_R1077_U243, P2_R1077_U244, P2_R1077_U245, P2_R1077_U246, P2_R1077_U247, P2_R1077_U248, P2_R1077_U249, P2_R1077_U25, P2_R1077_U250, P2_R1077_U251, P2_R1077_U252, P2_R1077_U253, P2_R1077_U254, P2_R1077_U255, P2_R1077_U256, P2_R1077_U257, P2_R1077_U258, P2_R1077_U259, P2_R1077_U26, P2_R1077_U260, P2_R1077_U261, P2_R1077_U262, P2_R1077_U263, P2_R1077_U264, P2_R1077_U265, P2_R1077_U266, P2_R1077_U267, P2_R1077_U268, P2_R1077_U269, P2_R1077_U27, P2_R1077_U270, P2_R1077_U271, P2_R1077_U272, P2_R1077_U273, P2_R1077_U274, P2_R1077_U275, P2_R1077_U276, P2_R1077_U277, P2_R1077_U278, P2_R1077_U279, P2_R1077_U28, P2_R1077_U280, P2_R1077_U281, P2_R1077_U282, P2_R1077_U283, P2_R1077_U284, P2_R1077_U285, P2_R1077_U286, P2_R1077_U287, P2_R1077_U288, P2_R1077_U289, P2_R1077_U29, P2_R1077_U290, P2_R1077_U291, P2_R1077_U292, P2_R1077_U293, P2_R1077_U294, P2_R1077_U295, P2_R1077_U296, P2_R1077_U297, P2_R1077_U298, P2_R1077_U299, P2_R1077_U30, P2_R1077_U300, P2_R1077_U301, P2_R1077_U302, P2_R1077_U303, P2_R1077_U304, P2_R1077_U305, P2_R1077_U306, P2_R1077_U307, P2_R1077_U308, P2_R1077_U309, P2_R1077_U31, P2_R1077_U310, P2_R1077_U311, P2_R1077_U312, P2_R1077_U313, P2_R1077_U314, P2_R1077_U315, P2_R1077_U316, P2_R1077_U317, P2_R1077_U318, P2_R1077_U319, P2_R1077_U32, P2_R1077_U320, P2_R1077_U321, P2_R1077_U322, P2_R1077_U323, P2_R1077_U324, P2_R1077_U325, P2_R1077_U326, P2_R1077_U327, P2_R1077_U328, P2_R1077_U329, P2_R1077_U33, P2_R1077_U330, P2_R1077_U331, P2_R1077_U332, P2_R1077_U333, P2_R1077_U334, P2_R1077_U335, P2_R1077_U336, P2_R1077_U337, P2_R1077_U338, P2_R1077_U339, P2_R1077_U34, P2_R1077_U340, P2_R1077_U341, P2_R1077_U342, P2_R1077_U343, P2_R1077_U344, P2_R1077_U345, P2_R1077_U346, P2_R1077_U347, P2_R1077_U348, P2_R1077_U349, P2_R1077_U35, P2_R1077_U350, P2_R1077_U351, P2_R1077_U352, P2_R1077_U353, P2_R1077_U354, P2_R1077_U355, P2_R1077_U356, P2_R1077_U357, P2_R1077_U358, P2_R1077_U359, P2_R1077_U36, P2_R1077_U360, P2_R1077_U361, P2_R1077_U362, P2_R1077_U363, P2_R1077_U364, P2_R1077_U365, P2_R1077_U366, P2_R1077_U367, P2_R1077_U368, P2_R1077_U369, P2_R1077_U37, P2_R1077_U370, P2_R1077_U371, P2_R1077_U372, P2_R1077_U373, P2_R1077_U374, P2_R1077_U375, P2_R1077_U376, P2_R1077_U377, P2_R1077_U378, P2_R1077_U379, P2_R1077_U38, P2_R1077_U380, P2_R1077_U381, P2_R1077_U382, P2_R1077_U383, P2_R1077_U384, P2_R1077_U385, P2_R1077_U386, P2_R1077_U387, P2_R1077_U388, P2_R1077_U389, P2_R1077_U39, P2_R1077_U390, P2_R1077_U391, P2_R1077_U392, P2_R1077_U393, P2_R1077_U394, P2_R1077_U395, P2_R1077_U396, P2_R1077_U397, P2_R1077_U398, P2_R1077_U399, P2_R1077_U4, P2_R1077_U40, P2_R1077_U400, P2_R1077_U401, P2_R1077_U402, P2_R1077_U403, P2_R1077_U404, P2_R1077_U405, P2_R1077_U406, P2_R1077_U407, P2_R1077_U408, P2_R1077_U409, P2_R1077_U41, P2_R1077_U410, P2_R1077_U411, P2_R1077_U412, P2_R1077_U413, P2_R1077_U414, P2_R1077_U415, P2_R1077_U416, P2_R1077_U417, P2_R1077_U418, P2_R1077_U419, P2_R1077_U42, P2_R1077_U420, P2_R1077_U421, P2_R1077_U422, P2_R1077_U423, P2_R1077_U424, P2_R1077_U425, P2_R1077_U426, P2_R1077_U427, P2_R1077_U428, P2_R1077_U429, P2_R1077_U43, P2_R1077_U430, P2_R1077_U431, P2_R1077_U432, P2_R1077_U433, P2_R1077_U434, P2_R1077_U435, P2_R1077_U436, P2_R1077_U437, P2_R1077_U438, P2_R1077_U439, P2_R1077_U44, P2_R1077_U440, P2_R1077_U441, P2_R1077_U442, P2_R1077_U443, P2_R1077_U444, P2_R1077_U445, P2_R1077_U446, P2_R1077_U447, P2_R1077_U448, P2_R1077_U449, P2_R1077_U45, P2_R1077_U450, P2_R1077_U451, P2_R1077_U452, P2_R1077_U453, P2_R1077_U454, P2_R1077_U455, P2_R1077_U456, P2_R1077_U457, P2_R1077_U458, P2_R1077_U459, P2_R1077_U46, P2_R1077_U460, P2_R1077_U461, P2_R1077_U462, P2_R1077_U463, P2_R1077_U464, P2_R1077_U465, P2_R1077_U466, P2_R1077_U467, P2_R1077_U468, P2_R1077_U469, P2_R1077_U47, P2_R1077_U470, P2_R1077_U471, P2_R1077_U472, P2_R1077_U473, P2_R1077_U474, P2_R1077_U475, P2_R1077_U476, P2_R1077_U477, P2_R1077_U478, P2_R1077_U479, P2_R1077_U48, P2_R1077_U480, P2_R1077_U481, P2_R1077_U482, P2_R1077_U483, P2_R1077_U484, P2_R1077_U485, P2_R1077_U486, P2_R1077_U487, P2_R1077_U488, P2_R1077_U489, P2_R1077_U49, P2_R1077_U490, P2_R1077_U491, P2_R1077_U492, P2_R1077_U493, P2_R1077_U494, P2_R1077_U495, P2_R1077_U496, P2_R1077_U497, P2_R1077_U498, P2_R1077_U499, P2_R1077_U5, P2_R1077_U50, P2_R1077_U500, P2_R1077_U501, P2_R1077_U502, P2_R1077_U503, P2_R1077_U504, P2_R1077_U51, P2_R1077_U52, P2_R1077_U53, P2_R1077_U54, P2_R1077_U55, P2_R1077_U56, P2_R1077_U57, P2_R1077_U58, P2_R1077_U59, P2_R1077_U6, P2_R1077_U60, P2_R1077_U61, P2_R1077_U62, P2_R1077_U63, P2_R1077_U64, P2_R1077_U65, P2_R1077_U66, P2_R1077_U67, P2_R1077_U68, P2_R1077_U69, P2_R1077_U7, P2_R1077_U70, P2_R1077_U71, P2_R1077_U72, P2_R1077_U73, P2_R1077_U74, P2_R1077_U75, P2_R1077_U76, P2_R1077_U77, P2_R1077_U78, P2_R1077_U79, P2_R1077_U8, P2_R1077_U80, P2_R1077_U81, P2_R1077_U82, P2_R1077_U83, P2_R1077_U84, P2_R1077_U85, P2_R1077_U86, P2_R1077_U87, P2_R1077_U88, P2_R1077_U89, P2_R1077_U9, P2_R1077_U90, P2_R1077_U91, P2_R1077_U92, P2_R1077_U93, P2_R1077_U94, P2_R1077_U95, P2_R1077_U96, P2_R1077_U97, P2_R1077_U98, P2_R1077_U99, P2_R1095_U10, P2_R1095_U100, P2_R1095_U101, P2_R1095_U102, P2_R1095_U103, P2_R1095_U104, P2_R1095_U105, P2_R1095_U106, P2_R1095_U107, P2_R1095_U108, P2_R1095_U109, P2_R1095_U11, P2_R1095_U110, P2_R1095_U111, P2_R1095_U112, P2_R1095_U113, P2_R1095_U114, P2_R1095_U115, P2_R1095_U116, P2_R1095_U117, P2_R1095_U118, P2_R1095_U119, P2_R1095_U12, P2_R1095_U120, P2_R1095_U121, P2_R1095_U122, P2_R1095_U123, P2_R1095_U124, P2_R1095_U125, P2_R1095_U126, P2_R1095_U127, P2_R1095_U128, P2_R1095_U129, P2_R1095_U13, P2_R1095_U130, P2_R1095_U131, P2_R1095_U132, P2_R1095_U133, P2_R1095_U134, P2_R1095_U135, P2_R1095_U136, P2_R1095_U137, P2_R1095_U138, P2_R1095_U139, P2_R1095_U14, P2_R1095_U140, P2_R1095_U141, P2_R1095_U142, P2_R1095_U143, P2_R1095_U144, P2_R1095_U145, P2_R1095_U146, P2_R1095_U147, P2_R1095_U148, P2_R1095_U149, P2_R1095_U15, P2_R1095_U150, P2_R1095_U151, P2_R1095_U152, P2_R1095_U153, P2_R1095_U154, P2_R1095_U155, P2_R1095_U156, P2_R1095_U157, P2_R1095_U158, P2_R1095_U159, P2_R1095_U16, P2_R1095_U160, P2_R1095_U161, P2_R1095_U162, P2_R1095_U163, P2_R1095_U164, P2_R1095_U165, P2_R1095_U166, P2_R1095_U167, P2_R1095_U168, P2_R1095_U169, P2_R1095_U17, P2_R1095_U170, P2_R1095_U171, P2_R1095_U172, P2_R1095_U173, P2_R1095_U174, P2_R1095_U175, P2_R1095_U176, P2_R1095_U177, P2_R1095_U178, P2_R1095_U179, P2_R1095_U18, P2_R1095_U180, P2_R1095_U181, P2_R1095_U182, P2_R1095_U183, P2_R1095_U184, P2_R1095_U185, P2_R1095_U186, P2_R1095_U187, P2_R1095_U188, P2_R1095_U189, P2_R1095_U19, P2_R1095_U190, P2_R1095_U191, P2_R1095_U192, P2_R1095_U193, P2_R1095_U194, P2_R1095_U195, P2_R1095_U196, P2_R1095_U197, P2_R1095_U198, P2_R1095_U199, P2_R1095_U20, P2_R1095_U200, P2_R1095_U201, P2_R1095_U202, P2_R1095_U203, P2_R1095_U204, P2_R1095_U205, P2_R1095_U206, P2_R1095_U207, P2_R1095_U208, P2_R1095_U209, P2_R1095_U21, P2_R1095_U210, P2_R1095_U211, P2_R1095_U212, P2_R1095_U213, P2_R1095_U214, P2_R1095_U215, P2_R1095_U216, P2_R1095_U217, P2_R1095_U218, P2_R1095_U219, P2_R1095_U22, P2_R1095_U220, P2_R1095_U221, P2_R1095_U222, P2_R1095_U223, P2_R1095_U224, P2_R1095_U225, P2_R1095_U226, P2_R1095_U227, P2_R1095_U228, P2_R1095_U229, P2_R1095_U23, P2_R1095_U230, P2_R1095_U231, P2_R1095_U232, P2_R1095_U233, P2_R1095_U234, P2_R1095_U235, P2_R1095_U236, P2_R1095_U237, P2_R1095_U238, P2_R1095_U239, P2_R1095_U24, P2_R1095_U240, P2_R1095_U241, P2_R1095_U242, P2_R1095_U243, P2_R1095_U244, P2_R1095_U245, P2_R1095_U246, P2_R1095_U247, P2_R1095_U248, P2_R1095_U249, P2_R1095_U25, P2_R1095_U250, P2_R1095_U251, P2_R1095_U252, P2_R1095_U253, P2_R1095_U254, P2_R1095_U255, P2_R1095_U256, P2_R1095_U257, P2_R1095_U258, P2_R1095_U259, P2_R1095_U26, P2_R1095_U260, P2_R1095_U261, P2_R1095_U262, P2_R1095_U263, P2_R1095_U264, P2_R1095_U265, P2_R1095_U266, P2_R1095_U267, P2_R1095_U268, P2_R1095_U269, P2_R1095_U27, P2_R1095_U270, P2_R1095_U271, P2_R1095_U272, P2_R1095_U273, P2_R1095_U274, P2_R1095_U275, P2_R1095_U276, P2_R1095_U277, P2_R1095_U278, P2_R1095_U279, P2_R1095_U28, P2_R1095_U280, P2_R1095_U281, P2_R1095_U282, P2_R1095_U283, P2_R1095_U284, P2_R1095_U285, P2_R1095_U286, P2_R1095_U287, P2_R1095_U288, P2_R1095_U289, P2_R1095_U29, P2_R1095_U290, P2_R1095_U291, P2_R1095_U292, P2_R1095_U293, P2_R1095_U294, P2_R1095_U295, P2_R1095_U296, P2_R1095_U297, P2_R1095_U298, P2_R1095_U299, P2_R1095_U30, P2_R1095_U300, P2_R1095_U301, P2_R1095_U302, P2_R1095_U303, P2_R1095_U304, P2_R1095_U305, P2_R1095_U306, P2_R1095_U307, P2_R1095_U308, P2_R1095_U309, P2_R1095_U31, P2_R1095_U310, P2_R1095_U311, P2_R1095_U312, P2_R1095_U313, P2_R1095_U314, P2_R1095_U315, P2_R1095_U316, P2_R1095_U317, P2_R1095_U318, P2_R1095_U319, P2_R1095_U32, P2_R1095_U320, P2_R1095_U321, P2_R1095_U322, P2_R1095_U323, P2_R1095_U324, P2_R1095_U325, P2_R1095_U326, P2_R1095_U327, P2_R1095_U328, P2_R1095_U329, P2_R1095_U33, P2_R1095_U330, P2_R1095_U331, P2_R1095_U332, P2_R1095_U333, P2_R1095_U334, P2_R1095_U335, P2_R1095_U336, P2_R1095_U337, P2_R1095_U338, P2_R1095_U339, P2_R1095_U34, P2_R1095_U340, P2_R1095_U341, P2_R1095_U342, P2_R1095_U343, P2_R1095_U344, P2_R1095_U345, P2_R1095_U346, P2_R1095_U347, P2_R1095_U348, P2_R1095_U349, P2_R1095_U35, P2_R1095_U350, P2_R1095_U351, P2_R1095_U352, P2_R1095_U353, P2_R1095_U354, P2_R1095_U355, P2_R1095_U356, P2_R1095_U357, P2_R1095_U358, P2_R1095_U359, P2_R1095_U36, P2_R1095_U360, P2_R1095_U361, P2_R1095_U362, P2_R1095_U363, P2_R1095_U364, P2_R1095_U365, P2_R1095_U366, P2_R1095_U367, P2_R1095_U368, P2_R1095_U369, P2_R1095_U37, P2_R1095_U370, P2_R1095_U371, P2_R1095_U372, P2_R1095_U373, P2_R1095_U374, P2_R1095_U375, P2_R1095_U376, P2_R1095_U377, P2_R1095_U378, P2_R1095_U379, P2_R1095_U38, P2_R1095_U380, P2_R1095_U381, P2_R1095_U382, P2_R1095_U383, P2_R1095_U384, P2_R1095_U385, P2_R1095_U386, P2_R1095_U387, P2_R1095_U388, P2_R1095_U389, P2_R1095_U39, P2_R1095_U390, P2_R1095_U391, P2_R1095_U392, P2_R1095_U393, P2_R1095_U394, P2_R1095_U395, P2_R1095_U396, P2_R1095_U397, P2_R1095_U398, P2_R1095_U399, P2_R1095_U40, P2_R1095_U400, P2_R1095_U401, P2_R1095_U402, P2_R1095_U403, P2_R1095_U404, P2_R1095_U405, P2_R1095_U406, P2_R1095_U407, P2_R1095_U408, P2_R1095_U409, P2_R1095_U41, P2_R1095_U410, P2_R1095_U411, P2_R1095_U412, P2_R1095_U413, P2_R1095_U414, P2_R1095_U415, P2_R1095_U416, P2_R1095_U417, P2_R1095_U418, P2_R1095_U419, P2_R1095_U42, P2_R1095_U420, P2_R1095_U421, P2_R1095_U422, P2_R1095_U423, P2_R1095_U424, P2_R1095_U425, P2_R1095_U426, P2_R1095_U427, P2_R1095_U428, P2_R1095_U429, P2_R1095_U43, P2_R1095_U430, P2_R1095_U431, P2_R1095_U432, P2_R1095_U433, P2_R1095_U434, P2_R1095_U435, P2_R1095_U436, P2_R1095_U437, P2_R1095_U438, P2_R1095_U439, P2_R1095_U44, P2_R1095_U440, P2_R1095_U441, P2_R1095_U442, P2_R1095_U443, P2_R1095_U444, P2_R1095_U445, P2_R1095_U446, P2_R1095_U447, P2_R1095_U448, P2_R1095_U449, P2_R1095_U45, P2_R1095_U450, P2_R1095_U451, P2_R1095_U452, P2_R1095_U453, P2_R1095_U454, P2_R1095_U455, P2_R1095_U456, P2_R1095_U457, P2_R1095_U458, P2_R1095_U459, P2_R1095_U46, P2_R1095_U460, P2_R1095_U461, P2_R1095_U462, P2_R1095_U463, P2_R1095_U464, P2_R1095_U465, P2_R1095_U466, P2_R1095_U467, P2_R1095_U468, P2_R1095_U469, P2_R1095_U47, P2_R1095_U470, P2_R1095_U471, P2_R1095_U472, P2_R1095_U473, P2_R1095_U474, P2_R1095_U475, P2_R1095_U476, P2_R1095_U477, P2_R1095_U478, P2_R1095_U479, P2_R1095_U48, P2_R1095_U480, P2_R1095_U481, P2_R1095_U482, P2_R1095_U483, P2_R1095_U484, P2_R1095_U485, P2_R1095_U486, P2_R1095_U487, P2_R1095_U488, P2_R1095_U489, P2_R1095_U49, P2_R1095_U50, P2_R1095_U51, P2_R1095_U52, P2_R1095_U53, P2_R1095_U54, P2_R1095_U55, P2_R1095_U56, P2_R1095_U57, P2_R1095_U58, P2_R1095_U59, P2_R1095_U6, P2_R1095_U60, P2_R1095_U61, P2_R1095_U62, P2_R1095_U63, P2_R1095_U64, P2_R1095_U65, P2_R1095_U66, P2_R1095_U67, P2_R1095_U68, P2_R1095_U69, P2_R1095_U7, P2_R1095_U70, P2_R1095_U71, P2_R1095_U72, P2_R1095_U73, P2_R1095_U74, P2_R1095_U75, P2_R1095_U76, P2_R1095_U77, P2_R1095_U78, P2_R1095_U79, P2_R1095_U8, P2_R1095_U80, P2_R1095_U81, P2_R1095_U82, P2_R1095_U83, P2_R1095_U84, P2_R1095_U85, P2_R1095_U86, P2_R1095_U87, P2_R1095_U88, P2_R1095_U89, P2_R1095_U9, P2_R1095_U90, P2_R1095_U91, P2_R1095_U92, P2_R1095_U93, P2_R1095_U94, P2_R1095_U95, P2_R1095_U96, P2_R1095_U97, P2_R1095_U98, P2_R1095_U99, P2_R1110_U10, P2_R1110_U100, P2_R1110_U101, P2_R1110_U102, P2_R1110_U103, P2_R1110_U104, P2_R1110_U105, P2_R1110_U106, P2_R1110_U107, P2_R1110_U108, P2_R1110_U109, P2_R1110_U11, P2_R1110_U110, P2_R1110_U111, P2_R1110_U112, P2_R1110_U113, P2_R1110_U114, P2_R1110_U115, P2_R1110_U116, P2_R1110_U117, P2_R1110_U118, P2_R1110_U119, P2_R1110_U12, P2_R1110_U120, P2_R1110_U121, P2_R1110_U122, P2_R1110_U123, P2_R1110_U124, P2_R1110_U125, P2_R1110_U126, P2_R1110_U127, P2_R1110_U128, P2_R1110_U129, P2_R1110_U13, P2_R1110_U130, P2_R1110_U131, P2_R1110_U132, P2_R1110_U133, P2_R1110_U134, P2_R1110_U135, P2_R1110_U136, P2_R1110_U137, P2_R1110_U138, P2_R1110_U139, P2_R1110_U14, P2_R1110_U140, P2_R1110_U141, P2_R1110_U142, P2_R1110_U143, P2_R1110_U144, P2_R1110_U145, P2_R1110_U146, P2_R1110_U147, P2_R1110_U148, P2_R1110_U149, P2_R1110_U15, P2_R1110_U150, P2_R1110_U151, P2_R1110_U152, P2_R1110_U153, P2_R1110_U154, P2_R1110_U155, P2_R1110_U156, P2_R1110_U157, P2_R1110_U158, P2_R1110_U159, P2_R1110_U16, P2_R1110_U160, P2_R1110_U161, P2_R1110_U162, P2_R1110_U163, P2_R1110_U164, P2_R1110_U165, P2_R1110_U166, P2_R1110_U167, P2_R1110_U168, P2_R1110_U169, P2_R1110_U17, P2_R1110_U170, P2_R1110_U171, P2_R1110_U172, P2_R1110_U173, P2_R1110_U174, P2_R1110_U175, P2_R1110_U176, P2_R1110_U177, P2_R1110_U178, P2_R1110_U179, P2_R1110_U18, P2_R1110_U180, P2_R1110_U181, P2_R1110_U182, P2_R1110_U183, P2_R1110_U184, P2_R1110_U185, P2_R1110_U186, P2_R1110_U187, P2_R1110_U188, P2_R1110_U189, P2_R1110_U19, P2_R1110_U190, P2_R1110_U191, P2_R1110_U192, P2_R1110_U193, P2_R1110_U194, P2_R1110_U195, P2_R1110_U196, P2_R1110_U197, P2_R1110_U198, P2_R1110_U199, P2_R1110_U20, P2_R1110_U200, P2_R1110_U201, P2_R1110_U202, P2_R1110_U203, P2_R1110_U204, P2_R1110_U205, P2_R1110_U206, P2_R1110_U207, P2_R1110_U208, P2_R1110_U209, P2_R1110_U21, P2_R1110_U210, P2_R1110_U211, P2_R1110_U212, P2_R1110_U213, P2_R1110_U214, P2_R1110_U215, P2_R1110_U216, P2_R1110_U217, P2_R1110_U218, P2_R1110_U219, P2_R1110_U22, P2_R1110_U220, P2_R1110_U221, P2_R1110_U222, P2_R1110_U223, P2_R1110_U224, P2_R1110_U225, P2_R1110_U226, P2_R1110_U227, P2_R1110_U228, P2_R1110_U229, P2_R1110_U23, P2_R1110_U230, P2_R1110_U231, P2_R1110_U232, P2_R1110_U233, P2_R1110_U234, P2_R1110_U235, P2_R1110_U236, P2_R1110_U237, P2_R1110_U238, P2_R1110_U239, P2_R1110_U24, P2_R1110_U240, P2_R1110_U241, P2_R1110_U242, P2_R1110_U243, P2_R1110_U244, P2_R1110_U245, P2_R1110_U246, P2_R1110_U247, P2_R1110_U248, P2_R1110_U249, P2_R1110_U25, P2_R1110_U250, P2_R1110_U251, P2_R1110_U252, P2_R1110_U253, P2_R1110_U254, P2_R1110_U255, P2_R1110_U256, P2_R1110_U257, P2_R1110_U258, P2_R1110_U259, P2_R1110_U26, P2_R1110_U260, P2_R1110_U261, P2_R1110_U262, P2_R1110_U263, P2_R1110_U264, P2_R1110_U265, P2_R1110_U266, P2_R1110_U267, P2_R1110_U268, P2_R1110_U269, P2_R1110_U27, P2_R1110_U270, P2_R1110_U271, P2_R1110_U272, P2_R1110_U273, P2_R1110_U274, P2_R1110_U275, P2_R1110_U276, P2_R1110_U277, P2_R1110_U278, P2_R1110_U279, P2_R1110_U28, P2_R1110_U280, P2_R1110_U281, P2_R1110_U282, P2_R1110_U283, P2_R1110_U284, P2_R1110_U285, P2_R1110_U286, P2_R1110_U287, P2_R1110_U288, P2_R1110_U289, P2_R1110_U29, P2_R1110_U290, P2_R1110_U291, P2_R1110_U292, P2_R1110_U293, P2_R1110_U294, P2_R1110_U295, P2_R1110_U296, P2_R1110_U297, P2_R1110_U298, P2_R1110_U299, P2_R1110_U30, P2_R1110_U300, P2_R1110_U301, P2_R1110_U302, P2_R1110_U303, P2_R1110_U304, P2_R1110_U305, P2_R1110_U306, P2_R1110_U307, P2_R1110_U308, P2_R1110_U309, P2_R1110_U31, P2_R1110_U310, P2_R1110_U311, P2_R1110_U312, P2_R1110_U313, P2_R1110_U314, P2_R1110_U315, P2_R1110_U316, P2_R1110_U317, P2_R1110_U318, P2_R1110_U319, P2_R1110_U32, P2_R1110_U320, P2_R1110_U321, P2_R1110_U322, P2_R1110_U323, P2_R1110_U324, P2_R1110_U325, P2_R1110_U326, P2_R1110_U327, P2_R1110_U328, P2_R1110_U329, P2_R1110_U33, P2_R1110_U330, P2_R1110_U331, P2_R1110_U332, P2_R1110_U333, P2_R1110_U334, P2_R1110_U335, P2_R1110_U336, P2_R1110_U337, P2_R1110_U338, P2_R1110_U339, P2_R1110_U34, P2_R1110_U340, P2_R1110_U341, P2_R1110_U342, P2_R1110_U343, P2_R1110_U344, P2_R1110_U345, P2_R1110_U346, P2_R1110_U347, P2_R1110_U348, P2_R1110_U349, P2_R1110_U35, P2_R1110_U350, P2_R1110_U351, P2_R1110_U352, P2_R1110_U353, P2_R1110_U354, P2_R1110_U355, P2_R1110_U356, P2_R1110_U357, P2_R1110_U358, P2_R1110_U359, P2_R1110_U36, P2_R1110_U360, P2_R1110_U361, P2_R1110_U362, P2_R1110_U363, P2_R1110_U364, P2_R1110_U365, P2_R1110_U366, P2_R1110_U367, P2_R1110_U368, P2_R1110_U369, P2_R1110_U37, P2_R1110_U370, P2_R1110_U371, P2_R1110_U372, P2_R1110_U373, P2_R1110_U374, P2_R1110_U375, P2_R1110_U376, P2_R1110_U377, P2_R1110_U378, P2_R1110_U379, P2_R1110_U38, P2_R1110_U380, P2_R1110_U381, P2_R1110_U382, P2_R1110_U383, P2_R1110_U384, P2_R1110_U385, P2_R1110_U386, P2_R1110_U387, P2_R1110_U388, P2_R1110_U389, P2_R1110_U39, P2_R1110_U390, P2_R1110_U391, P2_R1110_U392, P2_R1110_U393, P2_R1110_U394, P2_R1110_U395, P2_R1110_U396, P2_R1110_U397, P2_R1110_U398, P2_R1110_U399, P2_R1110_U4, P2_R1110_U40, P2_R1110_U400, P2_R1110_U401, P2_R1110_U402, P2_R1110_U403, P2_R1110_U404, P2_R1110_U405, P2_R1110_U406, P2_R1110_U407, P2_R1110_U408, P2_R1110_U409, P2_R1110_U41, P2_R1110_U410, P2_R1110_U411, P2_R1110_U412, P2_R1110_U413, P2_R1110_U414, P2_R1110_U415, P2_R1110_U416, P2_R1110_U417, P2_R1110_U418, P2_R1110_U419, P2_R1110_U42, P2_R1110_U420, P2_R1110_U421, P2_R1110_U422, P2_R1110_U423, P2_R1110_U424, P2_R1110_U425, P2_R1110_U426, P2_R1110_U427, P2_R1110_U428, P2_R1110_U429, P2_R1110_U43, P2_R1110_U430, P2_R1110_U431, P2_R1110_U432, P2_R1110_U433, P2_R1110_U434, P2_R1110_U435, P2_R1110_U436, P2_R1110_U437, P2_R1110_U438, P2_R1110_U439, P2_R1110_U44, P2_R1110_U440, P2_R1110_U441, P2_R1110_U442, P2_R1110_U443, P2_R1110_U444, P2_R1110_U445, P2_R1110_U446, P2_R1110_U447, P2_R1110_U448, P2_R1110_U449, P2_R1110_U45, P2_R1110_U450, P2_R1110_U451, P2_R1110_U452, P2_R1110_U453, P2_R1110_U454, P2_R1110_U455, P2_R1110_U456, P2_R1110_U457, P2_R1110_U458, P2_R1110_U459, P2_R1110_U46, P2_R1110_U460, P2_R1110_U461, P2_R1110_U462, P2_R1110_U463, P2_R1110_U464, P2_R1110_U465, P2_R1110_U466, P2_R1110_U467, P2_R1110_U468, P2_R1110_U469, P2_R1110_U47, P2_R1110_U470, P2_R1110_U471, P2_R1110_U472, P2_R1110_U473, P2_R1110_U474, P2_R1110_U475, P2_R1110_U476, P2_R1110_U477, P2_R1110_U478, P2_R1110_U479, P2_R1110_U48, P2_R1110_U480, P2_R1110_U481, P2_R1110_U482, P2_R1110_U483, P2_R1110_U484, P2_R1110_U485, P2_R1110_U486, P2_R1110_U487, P2_R1110_U488, P2_R1110_U489, P2_R1110_U49, P2_R1110_U490, P2_R1110_U491, P2_R1110_U492, P2_R1110_U493, P2_R1110_U494, P2_R1110_U495, P2_R1110_U496, P2_R1110_U497, P2_R1110_U498, P2_R1110_U499, P2_R1110_U5, P2_R1110_U50, P2_R1110_U500, P2_R1110_U501, P2_R1110_U502, P2_R1110_U503, P2_R1110_U504, P2_R1110_U51, P2_R1110_U52, P2_R1110_U53, P2_R1110_U54, P2_R1110_U55, P2_R1110_U56, P2_R1110_U57, P2_R1110_U58, P2_R1110_U59, P2_R1110_U6, P2_R1110_U60, P2_R1110_U61, P2_R1110_U62, P2_R1110_U63, P2_R1110_U64, P2_R1110_U65, P2_R1110_U66, P2_R1110_U67, P2_R1110_U68, P2_R1110_U69, P2_R1110_U7, P2_R1110_U70, P2_R1110_U71, P2_R1110_U72, P2_R1110_U73, P2_R1110_U74, P2_R1110_U75, P2_R1110_U76, P2_R1110_U77, P2_R1110_U78, P2_R1110_U79, P2_R1110_U8, P2_R1110_U80, P2_R1110_U81, P2_R1110_U82, P2_R1110_U83, P2_R1110_U84, P2_R1110_U85, P2_R1110_U86, P2_R1110_U87, P2_R1110_U88, P2_R1110_U89, P2_R1110_U9, P2_R1110_U90, P2_R1110_U91, P2_R1110_U92, P2_R1110_U93, P2_R1110_U94, P2_R1110_U95, P2_R1110_U96, P2_R1110_U97, P2_R1110_U98, P2_R1110_U99, P2_R1131_U10, P2_R1131_U100, P2_R1131_U101, P2_R1131_U102, P2_R1131_U103, P2_R1131_U104, P2_R1131_U105, P2_R1131_U106, P2_R1131_U107, P2_R1131_U108, P2_R1131_U109, P2_R1131_U11, P2_R1131_U110, P2_R1131_U111, P2_R1131_U112, P2_R1131_U113, P2_R1131_U114, P2_R1131_U115, P2_R1131_U116, P2_R1131_U117, P2_R1131_U118, P2_R1131_U119, P2_R1131_U12, P2_R1131_U120, P2_R1131_U121, P2_R1131_U122, P2_R1131_U123, P2_R1131_U124, P2_R1131_U125, P2_R1131_U126, P2_R1131_U127, P2_R1131_U128, P2_R1131_U129, P2_R1131_U13, P2_R1131_U130, P2_R1131_U131, P2_R1131_U132, P2_R1131_U133, P2_R1131_U134, P2_R1131_U135, P2_R1131_U136, P2_R1131_U137, P2_R1131_U138, P2_R1131_U139, P2_R1131_U14, P2_R1131_U140, P2_R1131_U141, P2_R1131_U142, P2_R1131_U143, P2_R1131_U144, P2_R1131_U145, P2_R1131_U146, P2_R1131_U147, P2_R1131_U148, P2_R1131_U149, P2_R1131_U15, P2_R1131_U150, P2_R1131_U151, P2_R1131_U152, P2_R1131_U153, P2_R1131_U154, P2_R1131_U155, P2_R1131_U156, P2_R1131_U157, P2_R1131_U158, P2_R1131_U159, P2_R1131_U16, P2_R1131_U160, P2_R1131_U161, P2_R1131_U162, P2_R1131_U163, P2_R1131_U164, P2_R1131_U165, P2_R1131_U166, P2_R1131_U167, P2_R1131_U168, P2_R1131_U169, P2_R1131_U17, P2_R1131_U170, P2_R1131_U171, P2_R1131_U172, P2_R1131_U173, P2_R1131_U174, P2_R1131_U175, P2_R1131_U176, P2_R1131_U177, P2_R1131_U178, P2_R1131_U179, P2_R1131_U18, P2_R1131_U180, P2_R1131_U181, P2_R1131_U182, P2_R1131_U183, P2_R1131_U184, P2_R1131_U185, P2_R1131_U186, P2_R1131_U187, P2_R1131_U188, P2_R1131_U189, P2_R1131_U19, P2_R1131_U190, P2_R1131_U191, P2_R1131_U192, P2_R1131_U193, P2_R1131_U194, P2_R1131_U195, P2_R1131_U196, P2_R1131_U197, P2_R1131_U198, P2_R1131_U199, P2_R1131_U20, P2_R1131_U200, P2_R1131_U201, P2_R1131_U202, P2_R1131_U203, P2_R1131_U204, P2_R1131_U205, P2_R1131_U206, P2_R1131_U207, P2_R1131_U208, P2_R1131_U209, P2_R1131_U21, P2_R1131_U210, P2_R1131_U211, P2_R1131_U212, P2_R1131_U213, P2_R1131_U214, P2_R1131_U215, P2_R1131_U216, P2_R1131_U217, P2_R1131_U218, P2_R1131_U219, P2_R1131_U22, P2_R1131_U220, P2_R1131_U221, P2_R1131_U222, P2_R1131_U223, P2_R1131_U224, P2_R1131_U225, P2_R1131_U226, P2_R1131_U227, P2_R1131_U228, P2_R1131_U229, P2_R1131_U23, P2_R1131_U230, P2_R1131_U231, P2_R1131_U232, P2_R1131_U233, P2_R1131_U234, P2_R1131_U235, P2_R1131_U236, P2_R1131_U237, P2_R1131_U238, P2_R1131_U239, P2_R1131_U24, P2_R1131_U240, P2_R1131_U241, P2_R1131_U242, P2_R1131_U243, P2_R1131_U244, P2_R1131_U245, P2_R1131_U246, P2_R1131_U247, P2_R1131_U248, P2_R1131_U249, P2_R1131_U25, P2_R1131_U250, P2_R1131_U251, P2_R1131_U252, P2_R1131_U253, P2_R1131_U254, P2_R1131_U255, P2_R1131_U256, P2_R1131_U257, P2_R1131_U258, P2_R1131_U259, P2_R1131_U26, P2_R1131_U260, P2_R1131_U261, P2_R1131_U262, P2_R1131_U263, P2_R1131_U264, P2_R1131_U265, P2_R1131_U266, P2_R1131_U267, P2_R1131_U268, P2_R1131_U269, P2_R1131_U27, P2_R1131_U270, P2_R1131_U271, P2_R1131_U272, P2_R1131_U273, P2_R1131_U274, P2_R1131_U275, P2_R1131_U276, P2_R1131_U277, P2_R1131_U278, P2_R1131_U279, P2_R1131_U28, P2_R1131_U280, P2_R1131_U281, P2_R1131_U282, P2_R1131_U283, P2_R1131_U284, P2_R1131_U285, P2_R1131_U286, P2_R1131_U287, P2_R1131_U288, P2_R1131_U289, P2_R1131_U29, P2_R1131_U290, P2_R1131_U291, P2_R1131_U292, P2_R1131_U293, P2_R1131_U294, P2_R1131_U295, P2_R1131_U296, P2_R1131_U297, P2_R1131_U298, P2_R1131_U299, P2_R1131_U30, P2_R1131_U300, P2_R1131_U301, P2_R1131_U302, P2_R1131_U303, P2_R1131_U304, P2_R1131_U305, P2_R1131_U306, P2_R1131_U307, P2_R1131_U308, P2_R1131_U309, P2_R1131_U31, P2_R1131_U310, P2_R1131_U311, P2_R1131_U312, P2_R1131_U313, P2_R1131_U314, P2_R1131_U315, P2_R1131_U316, P2_R1131_U317, P2_R1131_U318, P2_R1131_U319, P2_R1131_U32, P2_R1131_U320, P2_R1131_U321, P2_R1131_U322, P2_R1131_U323, P2_R1131_U324, P2_R1131_U325, P2_R1131_U326, P2_R1131_U327, P2_R1131_U328, P2_R1131_U329, P2_R1131_U33, P2_R1131_U330, P2_R1131_U331, P2_R1131_U332, P2_R1131_U333, P2_R1131_U334, P2_R1131_U335, P2_R1131_U336, P2_R1131_U337, P2_R1131_U338, P2_R1131_U339, P2_R1131_U34, P2_R1131_U340, P2_R1131_U341, P2_R1131_U342, P2_R1131_U343, P2_R1131_U344, P2_R1131_U345, P2_R1131_U346, P2_R1131_U347, P2_R1131_U348, P2_R1131_U349, P2_R1131_U35, P2_R1131_U350, P2_R1131_U351, P2_R1131_U352, P2_R1131_U353, P2_R1131_U354, P2_R1131_U355, P2_R1131_U356, P2_R1131_U357, P2_R1131_U358, P2_R1131_U359, P2_R1131_U36, P2_R1131_U360, P2_R1131_U361, P2_R1131_U362, P2_R1131_U363, P2_R1131_U364, P2_R1131_U365, P2_R1131_U366, P2_R1131_U367, P2_R1131_U368, P2_R1131_U369, P2_R1131_U37, P2_R1131_U370, P2_R1131_U371, P2_R1131_U372, P2_R1131_U373, P2_R1131_U374, P2_R1131_U375, P2_R1131_U376, P2_R1131_U377, P2_R1131_U378, P2_R1131_U379, P2_R1131_U38, P2_R1131_U380, P2_R1131_U381, P2_R1131_U382, P2_R1131_U383, P2_R1131_U384, P2_R1131_U385, P2_R1131_U386, P2_R1131_U387, P2_R1131_U388, P2_R1131_U389, P2_R1131_U39, P2_R1131_U390, P2_R1131_U391, P2_R1131_U392, P2_R1131_U393, P2_R1131_U394, P2_R1131_U395, P2_R1131_U396, P2_R1131_U397, P2_R1131_U398, P2_R1131_U399, P2_R1131_U40, P2_R1131_U400, P2_R1131_U401, P2_R1131_U402, P2_R1131_U403, P2_R1131_U404, P2_R1131_U405, P2_R1131_U406, P2_R1131_U407, P2_R1131_U408, P2_R1131_U409, P2_R1131_U41, P2_R1131_U410, P2_R1131_U411, P2_R1131_U412, P2_R1131_U413, P2_R1131_U414, P2_R1131_U415, P2_R1131_U416, P2_R1131_U417, P2_R1131_U418, P2_R1131_U419, P2_R1131_U42, P2_R1131_U420, P2_R1131_U421, P2_R1131_U422, P2_R1131_U423, P2_R1131_U424, P2_R1131_U425, P2_R1131_U426, P2_R1131_U427, P2_R1131_U428, P2_R1131_U429, P2_R1131_U43, P2_R1131_U430, P2_R1131_U431, P2_R1131_U432, P2_R1131_U433, P2_R1131_U434, P2_R1131_U435, P2_R1131_U436, P2_R1131_U437, P2_R1131_U438, P2_R1131_U439, P2_R1131_U44, P2_R1131_U440, P2_R1131_U441, P2_R1131_U442, P2_R1131_U443, P2_R1131_U444, P2_R1131_U445, P2_R1131_U446, P2_R1131_U447, P2_R1131_U448, P2_R1131_U449, P2_R1131_U45, P2_R1131_U450, P2_R1131_U451, P2_R1131_U452, P2_R1131_U453, P2_R1131_U454, P2_R1131_U455, P2_R1131_U456, P2_R1131_U457, P2_R1131_U458, P2_R1131_U459, P2_R1131_U46, P2_R1131_U460, P2_R1131_U461, P2_R1131_U462, P2_R1131_U463, P2_R1131_U464, P2_R1131_U465, P2_R1131_U466, P2_R1131_U467, P2_R1131_U468, P2_R1131_U469, P2_R1131_U47, P2_R1131_U470, P2_R1131_U471, P2_R1131_U472, P2_R1131_U473, P2_R1131_U474, P2_R1131_U475, P2_R1131_U476, P2_R1131_U477, P2_R1131_U478, P2_R1131_U479, P2_R1131_U48, P2_R1131_U480, P2_R1131_U481, P2_R1131_U482, P2_R1131_U483, P2_R1131_U484, P2_R1131_U485, P2_R1131_U486, P2_R1131_U487, P2_R1131_U488, P2_R1131_U489, P2_R1131_U49, P2_R1131_U50, P2_R1131_U51, P2_R1131_U52, P2_R1131_U53, P2_R1131_U54, P2_R1131_U55, P2_R1131_U56, P2_R1131_U57, P2_R1131_U58, P2_R1131_U59, P2_R1131_U6, P2_R1131_U60, P2_R1131_U61, P2_R1131_U62, P2_R1131_U63, P2_R1131_U64, P2_R1131_U65, P2_R1131_U66, P2_R1131_U67, P2_R1131_U68, P2_R1131_U69, P2_R1131_U7, P2_R1131_U70, P2_R1131_U71, P2_R1131_U72, P2_R1131_U73, P2_R1131_U74, P2_R1131_U75, P2_R1131_U76, P2_R1131_U77, P2_R1131_U78, P2_R1131_U79, P2_R1131_U8, P2_R1131_U80, P2_R1131_U81, P2_R1131_U82, P2_R1131_U83, P2_R1131_U84, P2_R1131_U85, P2_R1131_U86, P2_R1131_U87, P2_R1131_U88, P2_R1131_U89, P2_R1131_U9, P2_R1131_U90, P2_R1131_U91, P2_R1131_U92, P2_R1131_U93, P2_R1131_U94, P2_R1131_U95, P2_R1131_U96, P2_R1131_U97, P2_R1131_U98, P2_R1131_U99, P2_R1143_U10, P2_R1143_U100, P2_R1143_U101, P2_R1143_U102, P2_R1143_U103, P2_R1143_U104, P2_R1143_U105, P2_R1143_U106, P2_R1143_U107, P2_R1143_U108, P2_R1143_U109, P2_R1143_U11, P2_R1143_U110, P2_R1143_U111, P2_R1143_U112, P2_R1143_U113, P2_R1143_U114, P2_R1143_U115, P2_R1143_U116, P2_R1143_U117, P2_R1143_U118, P2_R1143_U119, P2_R1143_U12, P2_R1143_U120, P2_R1143_U121, P2_R1143_U122, P2_R1143_U123, P2_R1143_U124, P2_R1143_U125, P2_R1143_U126, P2_R1143_U127, P2_R1143_U128, P2_R1143_U129, P2_R1143_U13, P2_R1143_U130, P2_R1143_U131, P2_R1143_U132, P2_R1143_U133, P2_R1143_U134, P2_R1143_U135, P2_R1143_U136, P2_R1143_U137, P2_R1143_U138, P2_R1143_U139, P2_R1143_U14, P2_R1143_U140, P2_R1143_U141, P2_R1143_U142, P2_R1143_U143, P2_R1143_U144, P2_R1143_U145, P2_R1143_U146, P2_R1143_U147, P2_R1143_U148, P2_R1143_U149, P2_R1143_U15, P2_R1143_U150, P2_R1143_U151, P2_R1143_U152, P2_R1143_U153, P2_R1143_U154, P2_R1143_U155, P2_R1143_U156, P2_R1143_U157, P2_R1143_U158, P2_R1143_U159, P2_R1143_U16, P2_R1143_U160, P2_R1143_U161, P2_R1143_U162, P2_R1143_U163, P2_R1143_U164, P2_R1143_U165, P2_R1143_U166, P2_R1143_U167, P2_R1143_U168, P2_R1143_U169, P2_R1143_U17, P2_R1143_U170, P2_R1143_U171, P2_R1143_U172, P2_R1143_U173, P2_R1143_U174, P2_R1143_U175, P2_R1143_U176, P2_R1143_U177, P2_R1143_U178, P2_R1143_U179, P2_R1143_U18, P2_R1143_U180, P2_R1143_U181, P2_R1143_U182, P2_R1143_U183, P2_R1143_U184, P2_R1143_U185, P2_R1143_U186, P2_R1143_U187, P2_R1143_U188, P2_R1143_U189, P2_R1143_U19, P2_R1143_U190, P2_R1143_U191, P2_R1143_U192, P2_R1143_U193, P2_R1143_U194, P2_R1143_U195, P2_R1143_U196, P2_R1143_U197, P2_R1143_U198, P2_R1143_U199, P2_R1143_U20, P2_R1143_U200, P2_R1143_U201, P2_R1143_U202, P2_R1143_U203, P2_R1143_U204, P2_R1143_U205, P2_R1143_U206, P2_R1143_U207, P2_R1143_U208, P2_R1143_U209, P2_R1143_U21, P2_R1143_U210, P2_R1143_U211, P2_R1143_U212, P2_R1143_U213, P2_R1143_U214, P2_R1143_U215, P2_R1143_U216, P2_R1143_U217, P2_R1143_U218, P2_R1143_U219, P2_R1143_U22, P2_R1143_U220, P2_R1143_U221, P2_R1143_U222, P2_R1143_U223, P2_R1143_U224, P2_R1143_U225, P2_R1143_U226, P2_R1143_U227, P2_R1143_U228, P2_R1143_U229, P2_R1143_U23, P2_R1143_U230, P2_R1143_U231, P2_R1143_U232, P2_R1143_U233, P2_R1143_U234, P2_R1143_U235, P2_R1143_U236, P2_R1143_U237, P2_R1143_U238, P2_R1143_U239, P2_R1143_U24, P2_R1143_U240, P2_R1143_U241, P2_R1143_U242, P2_R1143_U243, P2_R1143_U244, P2_R1143_U245, P2_R1143_U246, P2_R1143_U247, P2_R1143_U248, P2_R1143_U249, P2_R1143_U25, P2_R1143_U250, P2_R1143_U251, P2_R1143_U252, P2_R1143_U253, P2_R1143_U254, P2_R1143_U255, P2_R1143_U256, P2_R1143_U257, P2_R1143_U258, P2_R1143_U259, P2_R1143_U26, P2_R1143_U260, P2_R1143_U261, P2_R1143_U262, P2_R1143_U263, P2_R1143_U264, P2_R1143_U265, P2_R1143_U266, P2_R1143_U267, P2_R1143_U268, P2_R1143_U269, P2_R1143_U27, P2_R1143_U270, P2_R1143_U271, P2_R1143_U272, P2_R1143_U273, P2_R1143_U274, P2_R1143_U275, P2_R1143_U276, P2_R1143_U277, P2_R1143_U278, P2_R1143_U279, P2_R1143_U28, P2_R1143_U280, P2_R1143_U281, P2_R1143_U282, P2_R1143_U283, P2_R1143_U284, P2_R1143_U285, P2_R1143_U286, P2_R1143_U287, P2_R1143_U288, P2_R1143_U289, P2_R1143_U29, P2_R1143_U290, P2_R1143_U291, P2_R1143_U292, P2_R1143_U293, P2_R1143_U294, P2_R1143_U295, P2_R1143_U296, P2_R1143_U297, P2_R1143_U298, P2_R1143_U299, P2_R1143_U30, P2_R1143_U300, P2_R1143_U301, P2_R1143_U302, P2_R1143_U303, P2_R1143_U304, P2_R1143_U305, P2_R1143_U306, P2_R1143_U307, P2_R1143_U308, P2_R1143_U309, P2_R1143_U31, P2_R1143_U310, P2_R1143_U311, P2_R1143_U312, P2_R1143_U313, P2_R1143_U314, P2_R1143_U315, P2_R1143_U316, P2_R1143_U317, P2_R1143_U318, P2_R1143_U319, P2_R1143_U32, P2_R1143_U320, P2_R1143_U321, P2_R1143_U322, P2_R1143_U323, P2_R1143_U324, P2_R1143_U325, P2_R1143_U326, P2_R1143_U327, P2_R1143_U328, P2_R1143_U329, P2_R1143_U33, P2_R1143_U330, P2_R1143_U331, P2_R1143_U332, P2_R1143_U333, P2_R1143_U334, P2_R1143_U335, P2_R1143_U336, P2_R1143_U337, P2_R1143_U338, P2_R1143_U339, P2_R1143_U34, P2_R1143_U340, P2_R1143_U341, P2_R1143_U342, P2_R1143_U343, P2_R1143_U344, P2_R1143_U345, P2_R1143_U346, P2_R1143_U347, P2_R1143_U348, P2_R1143_U349, P2_R1143_U35, P2_R1143_U350, P2_R1143_U351, P2_R1143_U352, P2_R1143_U353, P2_R1143_U354, P2_R1143_U355, P2_R1143_U356, P2_R1143_U357, P2_R1143_U358, P2_R1143_U359, P2_R1143_U36, P2_R1143_U360, P2_R1143_U361, P2_R1143_U362, P2_R1143_U363, P2_R1143_U364, P2_R1143_U365, P2_R1143_U366, P2_R1143_U367, P2_R1143_U368, P2_R1143_U369, P2_R1143_U37, P2_R1143_U370, P2_R1143_U371, P2_R1143_U372, P2_R1143_U373, P2_R1143_U374, P2_R1143_U375, P2_R1143_U376, P2_R1143_U377, P2_R1143_U378, P2_R1143_U379, P2_R1143_U38, P2_R1143_U380, P2_R1143_U381, P2_R1143_U382, P2_R1143_U383, P2_R1143_U384, P2_R1143_U385, P2_R1143_U386, P2_R1143_U387, P2_R1143_U388, P2_R1143_U389, P2_R1143_U39, P2_R1143_U390, P2_R1143_U391, P2_R1143_U392, P2_R1143_U393, P2_R1143_U394, P2_R1143_U395, P2_R1143_U396, P2_R1143_U397, P2_R1143_U398, P2_R1143_U399, P2_R1143_U4, P2_R1143_U40, P2_R1143_U400, P2_R1143_U401, P2_R1143_U402, P2_R1143_U403, P2_R1143_U404, P2_R1143_U405, P2_R1143_U406, P2_R1143_U407, P2_R1143_U408, P2_R1143_U409, P2_R1143_U41, P2_R1143_U410, P2_R1143_U411, P2_R1143_U412, P2_R1143_U413, P2_R1143_U414, P2_R1143_U415, P2_R1143_U416, P2_R1143_U417, P2_R1143_U418, P2_R1143_U419, P2_R1143_U42, P2_R1143_U420, P2_R1143_U421, P2_R1143_U422, P2_R1143_U423, P2_R1143_U424, P2_R1143_U425, P2_R1143_U426, P2_R1143_U427, P2_R1143_U428, P2_R1143_U429, P2_R1143_U43, P2_R1143_U430, P2_R1143_U431, P2_R1143_U432, P2_R1143_U433, P2_R1143_U434, P2_R1143_U435, P2_R1143_U436, P2_R1143_U437, P2_R1143_U438, P2_R1143_U439, P2_R1143_U44, P2_R1143_U440, P2_R1143_U441, P2_R1143_U442, P2_R1143_U443, P2_R1143_U444, P2_R1143_U445, P2_R1143_U446, P2_R1143_U447, P2_R1143_U448, P2_R1143_U449, P2_R1143_U45, P2_R1143_U450, P2_R1143_U451, P2_R1143_U452, P2_R1143_U453, P2_R1143_U454, P2_R1143_U455, P2_R1143_U456, P2_R1143_U457, P2_R1143_U458, P2_R1143_U459, P2_R1143_U46, P2_R1143_U460, P2_R1143_U461, P2_R1143_U462, P2_R1143_U463, P2_R1143_U464, P2_R1143_U465, P2_R1143_U466, P2_R1143_U467, P2_R1143_U468, P2_R1143_U469, P2_R1143_U47, P2_R1143_U470, P2_R1143_U471, P2_R1143_U472, P2_R1143_U473, P2_R1143_U474, P2_R1143_U475, P2_R1143_U476, P2_R1143_U477, P2_R1143_U478, P2_R1143_U479, P2_R1143_U48, P2_R1143_U480, P2_R1143_U481, P2_R1143_U482, P2_R1143_U483, P2_R1143_U484, P2_R1143_U485, P2_R1143_U486, P2_R1143_U487, P2_R1143_U488, P2_R1143_U489, P2_R1143_U49, P2_R1143_U490, P2_R1143_U491, P2_R1143_U492, P2_R1143_U493, P2_R1143_U494, P2_R1143_U495, P2_R1143_U496, P2_R1143_U497, P2_R1143_U498, P2_R1143_U499, P2_R1143_U5, P2_R1143_U50, P2_R1143_U500, P2_R1143_U501, P2_R1143_U502, P2_R1143_U503, P2_R1143_U504, P2_R1143_U51, P2_R1143_U52, P2_R1143_U53, P2_R1143_U54, P2_R1143_U55, P2_R1143_U56, P2_R1143_U57, P2_R1143_U58, P2_R1143_U59, P2_R1143_U6, P2_R1143_U60, P2_R1143_U61, P2_R1143_U62, P2_R1143_U63, P2_R1143_U64, P2_R1143_U65, P2_R1143_U66, P2_R1143_U67, P2_R1143_U68, P2_R1143_U69, P2_R1143_U7, P2_R1143_U70, P2_R1143_U71, P2_R1143_U72, P2_R1143_U73, P2_R1143_U74, P2_R1143_U75, P2_R1143_U76, P2_R1143_U77, P2_R1143_U78, P2_R1143_U79, P2_R1143_U8, P2_R1143_U80, P2_R1143_U81, P2_R1143_U82, P2_R1143_U83, P2_R1143_U84, P2_R1143_U85, P2_R1143_U86, P2_R1143_U87, P2_R1143_U88, P2_R1143_U89, P2_R1143_U9, P2_R1143_U90, P2_R1143_U91, P2_R1143_U92, P2_R1143_U93, P2_R1143_U94, P2_R1143_U95, P2_R1143_U96, P2_R1143_U97, P2_R1143_U98, P2_R1143_U99, P2_R1158_U10, P2_R1158_U100, P2_R1158_U101, P2_R1158_U102, P2_R1158_U103, P2_R1158_U104, P2_R1158_U105, P2_R1158_U106, P2_R1158_U107, P2_R1158_U108, P2_R1158_U109, P2_R1158_U11, P2_R1158_U110, P2_R1158_U111, P2_R1158_U112, P2_R1158_U113, P2_R1158_U114, P2_R1158_U115, P2_R1158_U116, P2_R1158_U117, P2_R1158_U118, P2_R1158_U119, P2_R1158_U12, P2_R1158_U120, P2_R1158_U121, P2_R1158_U122, P2_R1158_U123, P2_R1158_U124, P2_R1158_U125, P2_R1158_U126, P2_R1158_U127, P2_R1158_U128, P2_R1158_U129, P2_R1158_U13, P2_R1158_U130, P2_R1158_U131, P2_R1158_U132, P2_R1158_U133, P2_R1158_U134, P2_R1158_U135, P2_R1158_U136, P2_R1158_U137, P2_R1158_U138, P2_R1158_U139, P2_R1158_U14, P2_R1158_U140, P2_R1158_U141, P2_R1158_U142, P2_R1158_U143, P2_R1158_U144, P2_R1158_U145, P2_R1158_U146, P2_R1158_U147, P2_R1158_U148, P2_R1158_U149, P2_R1158_U15, P2_R1158_U150, P2_R1158_U151, P2_R1158_U152, P2_R1158_U153, P2_R1158_U154, P2_R1158_U155, P2_R1158_U156, P2_R1158_U157, P2_R1158_U158, P2_R1158_U159, P2_R1158_U16, P2_R1158_U160, P2_R1158_U161, P2_R1158_U162, P2_R1158_U163, P2_R1158_U164, P2_R1158_U165, P2_R1158_U166, P2_R1158_U167, P2_R1158_U168, P2_R1158_U169, P2_R1158_U17, P2_R1158_U170, P2_R1158_U171, P2_R1158_U172, P2_R1158_U173, P2_R1158_U174, P2_R1158_U175, P2_R1158_U176, P2_R1158_U177, P2_R1158_U178, P2_R1158_U179, P2_R1158_U18, P2_R1158_U180, P2_R1158_U181, P2_R1158_U182, P2_R1158_U183, P2_R1158_U184, P2_R1158_U185, P2_R1158_U186, P2_R1158_U187, P2_R1158_U188, P2_R1158_U189, P2_R1158_U19, P2_R1158_U190, P2_R1158_U191, P2_R1158_U192, P2_R1158_U193, P2_R1158_U194, P2_R1158_U195, P2_R1158_U196, P2_R1158_U197, P2_R1158_U198, P2_R1158_U199, P2_R1158_U20, P2_R1158_U200, P2_R1158_U201, P2_R1158_U202, P2_R1158_U203, P2_R1158_U204, P2_R1158_U205, P2_R1158_U206, P2_R1158_U207, P2_R1158_U208, P2_R1158_U209, P2_R1158_U21, P2_R1158_U210, P2_R1158_U211, P2_R1158_U212, P2_R1158_U213, P2_R1158_U214, P2_R1158_U215, P2_R1158_U216, P2_R1158_U217, P2_R1158_U218, P2_R1158_U219, P2_R1158_U22, P2_R1158_U220, P2_R1158_U221, P2_R1158_U222, P2_R1158_U223, P2_R1158_U224, P2_R1158_U225, P2_R1158_U226, P2_R1158_U227, P2_R1158_U228, P2_R1158_U229, P2_R1158_U23, P2_R1158_U230, P2_R1158_U231, P2_R1158_U232, P2_R1158_U233, P2_R1158_U234, P2_R1158_U235, P2_R1158_U236, P2_R1158_U237, P2_R1158_U238, P2_R1158_U239, P2_R1158_U24, P2_R1158_U240, P2_R1158_U241, P2_R1158_U242, P2_R1158_U243, P2_R1158_U244, P2_R1158_U245, P2_R1158_U246, P2_R1158_U247, P2_R1158_U248, P2_R1158_U249, P2_R1158_U25, P2_R1158_U250, P2_R1158_U251, P2_R1158_U252, P2_R1158_U253, P2_R1158_U254, P2_R1158_U255, P2_R1158_U256, P2_R1158_U257, P2_R1158_U258, P2_R1158_U259, P2_R1158_U26, P2_R1158_U260, P2_R1158_U261, P2_R1158_U262, P2_R1158_U263, P2_R1158_U264, P2_R1158_U265, P2_R1158_U266, P2_R1158_U267, P2_R1158_U268, P2_R1158_U269, P2_R1158_U27, P2_R1158_U270, P2_R1158_U271, P2_R1158_U272, P2_R1158_U273, P2_R1158_U274, P2_R1158_U275, P2_R1158_U276, P2_R1158_U277, P2_R1158_U278, P2_R1158_U279, P2_R1158_U28, P2_R1158_U280, P2_R1158_U281, P2_R1158_U282, P2_R1158_U283, P2_R1158_U284, P2_R1158_U285, P2_R1158_U286, P2_R1158_U287, P2_R1158_U288, P2_R1158_U289, P2_R1158_U29, P2_R1158_U290, P2_R1158_U291, P2_R1158_U292, P2_R1158_U293, P2_R1158_U294, P2_R1158_U295, P2_R1158_U296, P2_R1158_U297, P2_R1158_U298, P2_R1158_U299, P2_R1158_U30, P2_R1158_U300, P2_R1158_U301, P2_R1158_U302, P2_R1158_U303, P2_R1158_U304, P2_R1158_U305, P2_R1158_U306, P2_R1158_U307, P2_R1158_U308, P2_R1158_U309, P2_R1158_U31, P2_R1158_U310, P2_R1158_U311, P2_R1158_U312, P2_R1158_U313, P2_R1158_U314, P2_R1158_U315, P2_R1158_U316, P2_R1158_U317, P2_R1158_U318, P2_R1158_U319, P2_R1158_U32, P2_R1158_U320, P2_R1158_U321, P2_R1158_U322, P2_R1158_U323, P2_R1158_U324, P2_R1158_U325, P2_R1158_U326, P2_R1158_U327, P2_R1158_U328, P2_R1158_U329, P2_R1158_U33, P2_R1158_U330, P2_R1158_U331, P2_R1158_U332, P2_R1158_U333, P2_R1158_U334, P2_R1158_U335, P2_R1158_U336, P2_R1158_U337, P2_R1158_U338, P2_R1158_U339, P2_R1158_U34, P2_R1158_U340, P2_R1158_U341, P2_R1158_U342, P2_R1158_U343, P2_R1158_U344, P2_R1158_U345, P2_R1158_U346, P2_R1158_U347, P2_R1158_U348, P2_R1158_U349, P2_R1158_U35, P2_R1158_U350, P2_R1158_U351, P2_R1158_U352, P2_R1158_U353, P2_R1158_U354, P2_R1158_U355, P2_R1158_U356, P2_R1158_U357, P2_R1158_U358, P2_R1158_U359, P2_R1158_U36, P2_R1158_U360, P2_R1158_U361, P2_R1158_U362, P2_R1158_U363, P2_R1158_U364, P2_R1158_U365, P2_R1158_U366, P2_R1158_U367, P2_R1158_U368, P2_R1158_U369, P2_R1158_U37, P2_R1158_U370, P2_R1158_U371, P2_R1158_U372, P2_R1158_U373, P2_R1158_U374, P2_R1158_U375, P2_R1158_U376, P2_R1158_U377, P2_R1158_U378, P2_R1158_U379, P2_R1158_U38, P2_R1158_U380, P2_R1158_U381, P2_R1158_U382, P2_R1158_U383, P2_R1158_U384, P2_R1158_U385, P2_R1158_U386, P2_R1158_U387, P2_R1158_U388, P2_R1158_U389, P2_R1158_U39, P2_R1158_U390, P2_R1158_U391, P2_R1158_U392, P2_R1158_U393, P2_R1158_U394, P2_R1158_U395, P2_R1158_U396, P2_R1158_U397, P2_R1158_U398, P2_R1158_U399, P2_R1158_U4, P2_R1158_U40, P2_R1158_U400, P2_R1158_U401, P2_R1158_U402, P2_R1158_U403, P2_R1158_U404, P2_R1158_U405, P2_R1158_U406, P2_R1158_U407, P2_R1158_U408, P2_R1158_U409, P2_R1158_U41, P2_R1158_U410, P2_R1158_U411, P2_R1158_U412, P2_R1158_U413, P2_R1158_U414, P2_R1158_U415, P2_R1158_U416, P2_R1158_U417, P2_R1158_U418, P2_R1158_U419, P2_R1158_U42, P2_R1158_U420, P2_R1158_U421, P2_R1158_U422, P2_R1158_U423, P2_R1158_U424, P2_R1158_U425, P2_R1158_U426, P2_R1158_U427, P2_R1158_U428, P2_R1158_U429, P2_R1158_U43, P2_R1158_U430, P2_R1158_U431, P2_R1158_U432, P2_R1158_U433, P2_R1158_U434, P2_R1158_U435, P2_R1158_U436, P2_R1158_U437, P2_R1158_U438, P2_R1158_U439, P2_R1158_U44, P2_R1158_U440, P2_R1158_U441, P2_R1158_U442, P2_R1158_U443, P2_R1158_U444, P2_R1158_U445, P2_R1158_U446, P2_R1158_U447, P2_R1158_U448, P2_R1158_U449, P2_R1158_U45, P2_R1158_U450, P2_R1158_U451, P2_R1158_U452, P2_R1158_U453, P2_R1158_U454, P2_R1158_U455, P2_R1158_U456, P2_R1158_U457, P2_R1158_U458, P2_R1158_U459, P2_R1158_U46, P2_R1158_U460, P2_R1158_U461, P2_R1158_U462, P2_R1158_U463, P2_R1158_U464, P2_R1158_U465, P2_R1158_U466, P2_R1158_U467, P2_R1158_U468, P2_R1158_U469, P2_R1158_U47, P2_R1158_U470, P2_R1158_U471, P2_R1158_U472, P2_R1158_U473, P2_R1158_U474, P2_R1158_U475, P2_R1158_U476, P2_R1158_U477, P2_R1158_U478, P2_R1158_U479, P2_R1158_U48, P2_R1158_U480, P2_R1158_U481, P2_R1158_U482, P2_R1158_U483, P2_R1158_U484, P2_R1158_U485, P2_R1158_U486, P2_R1158_U487, P2_R1158_U488, P2_R1158_U489, P2_R1158_U49, P2_R1158_U490, P2_R1158_U491, P2_R1158_U492, P2_R1158_U493, P2_R1158_U494, P2_R1158_U495, P2_R1158_U496, P2_R1158_U497, P2_R1158_U498, P2_R1158_U499, P2_R1158_U5, P2_R1158_U50, P2_R1158_U500, P2_R1158_U501, P2_R1158_U502, P2_R1158_U503, P2_R1158_U504, P2_R1158_U505, P2_R1158_U506, P2_R1158_U507, P2_R1158_U508, P2_R1158_U509, P2_R1158_U51, P2_R1158_U510, P2_R1158_U511, P2_R1158_U512, P2_R1158_U513, P2_R1158_U514, P2_R1158_U515, P2_R1158_U516, P2_R1158_U517, P2_R1158_U518, P2_R1158_U519, P2_R1158_U52, P2_R1158_U520, P2_R1158_U521, P2_R1158_U522, P2_R1158_U523, P2_R1158_U524, P2_R1158_U525, P2_R1158_U526, P2_R1158_U527, P2_R1158_U528, P2_R1158_U529, P2_R1158_U53, P2_R1158_U530, P2_R1158_U531, P2_R1158_U532, P2_R1158_U533, P2_R1158_U534, P2_R1158_U535, P2_R1158_U536, P2_R1158_U537, P2_R1158_U538, P2_R1158_U539, P2_R1158_U54, P2_R1158_U540, P2_R1158_U541, P2_R1158_U542, P2_R1158_U543, P2_R1158_U544, P2_R1158_U545, P2_R1158_U546, P2_R1158_U547, P2_R1158_U548, P2_R1158_U549, P2_R1158_U55, P2_R1158_U550, P2_R1158_U551, P2_R1158_U552, P2_R1158_U553, P2_R1158_U554, P2_R1158_U555, P2_R1158_U556, P2_R1158_U557, P2_R1158_U558, P2_R1158_U559, P2_R1158_U56, P2_R1158_U560, P2_R1158_U561, P2_R1158_U562, P2_R1158_U563, P2_R1158_U564, P2_R1158_U565, P2_R1158_U566, P2_R1158_U567, P2_R1158_U568, P2_R1158_U569, P2_R1158_U57, P2_R1158_U570, P2_R1158_U571, P2_R1158_U572, P2_R1158_U573, P2_R1158_U574, P2_R1158_U575, P2_R1158_U576, P2_R1158_U577, P2_R1158_U578, P2_R1158_U579, P2_R1158_U58, P2_R1158_U580, P2_R1158_U581, P2_R1158_U582, P2_R1158_U583, P2_R1158_U584, P2_R1158_U585, P2_R1158_U586, P2_R1158_U587, P2_R1158_U588, P2_R1158_U589, P2_R1158_U59, P2_R1158_U590, P2_R1158_U591, P2_R1158_U592, P2_R1158_U593, P2_R1158_U594, P2_R1158_U595, P2_R1158_U596, P2_R1158_U597, P2_R1158_U598, P2_R1158_U599, P2_R1158_U6, P2_R1158_U60, P2_R1158_U600, P2_R1158_U601, P2_R1158_U602, P2_R1158_U603, P2_R1158_U604, P2_R1158_U605, P2_R1158_U606, P2_R1158_U607, P2_R1158_U608, P2_R1158_U609, P2_R1158_U61, P2_R1158_U610, P2_R1158_U611, P2_R1158_U612, P2_R1158_U613, P2_R1158_U614, P2_R1158_U615, P2_R1158_U616, P2_R1158_U617, P2_R1158_U618, P2_R1158_U619, P2_R1158_U62, P2_R1158_U620, P2_R1158_U621, P2_R1158_U622, P2_R1158_U623, P2_R1158_U624, P2_R1158_U625, P2_R1158_U626, P2_R1158_U627, P2_R1158_U628, P2_R1158_U629, P2_R1158_U63, P2_R1158_U630, P2_R1158_U631, P2_R1158_U632, P2_R1158_U633, P2_R1158_U634, P2_R1158_U64, P2_R1158_U65, P2_R1158_U66, P2_R1158_U67, P2_R1158_U68, P2_R1158_U69, P2_R1158_U7, P2_R1158_U70, P2_R1158_U71, P2_R1158_U72, P2_R1158_U73, P2_R1158_U74, P2_R1158_U75, P2_R1158_U76, P2_R1158_U77, P2_R1158_U78, P2_R1158_U79, P2_R1158_U8, P2_R1158_U80, P2_R1158_U81, P2_R1158_U82, P2_R1158_U83, P2_R1158_U84, P2_R1158_U85, P2_R1158_U86, P2_R1158_U87, P2_R1158_U88, P2_R1158_U89, P2_R1158_U9, P2_R1158_U90, P2_R1158_U91, P2_R1158_U92, P2_R1158_U93, P2_R1158_U94, P2_R1158_U95, P2_R1158_U96, P2_R1158_U97, P2_R1158_U98, P2_R1158_U99, P2_R1161_U10, P2_R1161_U100, P2_R1161_U101, P2_R1161_U102, P2_R1161_U103, P2_R1161_U104, P2_R1161_U105, P2_R1161_U106, P2_R1161_U107, P2_R1161_U108, P2_R1161_U109, P2_R1161_U11, P2_R1161_U110, P2_R1161_U111, P2_R1161_U112, P2_R1161_U113, P2_R1161_U114, P2_R1161_U115, P2_R1161_U116, P2_R1161_U117, P2_R1161_U118, P2_R1161_U119, P2_R1161_U12, P2_R1161_U120, P2_R1161_U121, P2_R1161_U122, P2_R1161_U123, P2_R1161_U124, P2_R1161_U125, P2_R1161_U126, P2_R1161_U127, P2_R1161_U128, P2_R1161_U129, P2_R1161_U13, P2_R1161_U130, P2_R1161_U131, P2_R1161_U132, P2_R1161_U133, P2_R1161_U134, P2_R1161_U135, P2_R1161_U136, P2_R1161_U137, P2_R1161_U138, P2_R1161_U139, P2_R1161_U14, P2_R1161_U140, P2_R1161_U141, P2_R1161_U142, P2_R1161_U143, P2_R1161_U144, P2_R1161_U145, P2_R1161_U146, P2_R1161_U147, P2_R1161_U148, P2_R1161_U149, P2_R1161_U15, P2_R1161_U150, P2_R1161_U151, P2_R1161_U152, P2_R1161_U153, P2_R1161_U154, P2_R1161_U155, P2_R1161_U156, P2_R1161_U157, P2_R1161_U158, P2_R1161_U159, P2_R1161_U16, P2_R1161_U160, P2_R1161_U161, P2_R1161_U162, P2_R1161_U163, P2_R1161_U164, P2_R1161_U165, P2_R1161_U166, P2_R1161_U167, P2_R1161_U168, P2_R1161_U169, P2_R1161_U17, P2_R1161_U170, P2_R1161_U171, P2_R1161_U172, P2_R1161_U173, P2_R1161_U174, P2_R1161_U175, P2_R1161_U176, P2_R1161_U177, P2_R1161_U178, P2_R1161_U179, P2_R1161_U18, P2_R1161_U180, P2_R1161_U181, P2_R1161_U182, P2_R1161_U183, P2_R1161_U184, P2_R1161_U185, P2_R1161_U186, P2_R1161_U187, P2_R1161_U188, P2_R1161_U189, P2_R1161_U19, P2_R1161_U190, P2_R1161_U191, P2_R1161_U192, P2_R1161_U193, P2_R1161_U194, P2_R1161_U195, P2_R1161_U196, P2_R1161_U197, P2_R1161_U198, P2_R1161_U199, P2_R1161_U20, P2_R1161_U200, P2_R1161_U201, P2_R1161_U202, P2_R1161_U203, P2_R1161_U204, P2_R1161_U205, P2_R1161_U206, P2_R1161_U207, P2_R1161_U208, P2_R1161_U209, P2_R1161_U21, P2_R1161_U210, P2_R1161_U211, P2_R1161_U212, P2_R1161_U213, P2_R1161_U214, P2_R1161_U215, P2_R1161_U216, P2_R1161_U217, P2_R1161_U218, P2_R1161_U219, P2_R1161_U22, P2_R1161_U220, P2_R1161_U221, P2_R1161_U222, P2_R1161_U223, P2_R1161_U224, P2_R1161_U225, P2_R1161_U226, P2_R1161_U227, P2_R1161_U228, P2_R1161_U229, P2_R1161_U23, P2_R1161_U230, P2_R1161_U231, P2_R1161_U232, P2_R1161_U233, P2_R1161_U234, P2_R1161_U235, P2_R1161_U236, P2_R1161_U237, P2_R1161_U238, P2_R1161_U239, P2_R1161_U24, P2_R1161_U240, P2_R1161_U241, P2_R1161_U242, P2_R1161_U243, P2_R1161_U244, P2_R1161_U245, P2_R1161_U246, P2_R1161_U247, P2_R1161_U248, P2_R1161_U249, P2_R1161_U25, P2_R1161_U250, P2_R1161_U251, P2_R1161_U252, P2_R1161_U253, P2_R1161_U254, P2_R1161_U255, P2_R1161_U256, P2_R1161_U257, P2_R1161_U258, P2_R1161_U259, P2_R1161_U26, P2_R1161_U260, P2_R1161_U261, P2_R1161_U262, P2_R1161_U263, P2_R1161_U264, P2_R1161_U265, P2_R1161_U266, P2_R1161_U267, P2_R1161_U268, P2_R1161_U269, P2_R1161_U27, P2_R1161_U270, P2_R1161_U271, P2_R1161_U272, P2_R1161_U273, P2_R1161_U274, P2_R1161_U275, P2_R1161_U276, P2_R1161_U277, P2_R1161_U278, P2_R1161_U279, P2_R1161_U28, P2_R1161_U280, P2_R1161_U281, P2_R1161_U282, P2_R1161_U283, P2_R1161_U284, P2_R1161_U285, P2_R1161_U286, P2_R1161_U287, P2_R1161_U288, P2_R1161_U289, P2_R1161_U29, P2_R1161_U290, P2_R1161_U291, P2_R1161_U292, P2_R1161_U293, P2_R1161_U294, P2_R1161_U295, P2_R1161_U296, P2_R1161_U297, P2_R1161_U298, P2_R1161_U299, P2_R1161_U30, P2_R1161_U300, P2_R1161_U301, P2_R1161_U302, P2_R1161_U303, P2_R1161_U304, P2_R1161_U305, P2_R1161_U306, P2_R1161_U307, P2_R1161_U308, P2_R1161_U309, P2_R1161_U31, P2_R1161_U310, P2_R1161_U311, P2_R1161_U312, P2_R1161_U313, P2_R1161_U314, P2_R1161_U315, P2_R1161_U316, P2_R1161_U317, P2_R1161_U318, P2_R1161_U319, P2_R1161_U32, P2_R1161_U320, P2_R1161_U321, P2_R1161_U322, P2_R1161_U323, P2_R1161_U324, P2_R1161_U325, P2_R1161_U326, P2_R1161_U327, P2_R1161_U328, P2_R1161_U329, P2_R1161_U33, P2_R1161_U330, P2_R1161_U331, P2_R1161_U332, P2_R1161_U333, P2_R1161_U334, P2_R1161_U335, P2_R1161_U336, P2_R1161_U337, P2_R1161_U338, P2_R1161_U339, P2_R1161_U34, P2_R1161_U340, P2_R1161_U341, P2_R1161_U342, P2_R1161_U343, P2_R1161_U344, P2_R1161_U345, P2_R1161_U346, P2_R1161_U347, P2_R1161_U348, P2_R1161_U349, P2_R1161_U35, P2_R1161_U350, P2_R1161_U351, P2_R1161_U352, P2_R1161_U353, P2_R1161_U354, P2_R1161_U355, P2_R1161_U356, P2_R1161_U357, P2_R1161_U358, P2_R1161_U359, P2_R1161_U36, P2_R1161_U360, P2_R1161_U361, P2_R1161_U362, P2_R1161_U363, P2_R1161_U364, P2_R1161_U365, P2_R1161_U366, P2_R1161_U367, P2_R1161_U368, P2_R1161_U369, P2_R1161_U37, P2_R1161_U370, P2_R1161_U371, P2_R1161_U372, P2_R1161_U373, P2_R1161_U374, P2_R1161_U375, P2_R1161_U376, P2_R1161_U377, P2_R1161_U378, P2_R1161_U379, P2_R1161_U38, P2_R1161_U380, P2_R1161_U381, P2_R1161_U382, P2_R1161_U383, P2_R1161_U384, P2_R1161_U385, P2_R1161_U386, P2_R1161_U387, P2_R1161_U388, P2_R1161_U389, P2_R1161_U39, P2_R1161_U390, P2_R1161_U391, P2_R1161_U392, P2_R1161_U393, P2_R1161_U394, P2_R1161_U395, P2_R1161_U396, P2_R1161_U397, P2_R1161_U398, P2_R1161_U399, P2_R1161_U4, P2_R1161_U40, P2_R1161_U400, P2_R1161_U401, P2_R1161_U402, P2_R1161_U403, P2_R1161_U404, P2_R1161_U405, P2_R1161_U406, P2_R1161_U407, P2_R1161_U408, P2_R1161_U409, P2_R1161_U41, P2_R1161_U410, P2_R1161_U411, P2_R1161_U412, P2_R1161_U413, P2_R1161_U414, P2_R1161_U415, P2_R1161_U416, P2_R1161_U417, P2_R1161_U418, P2_R1161_U419, P2_R1161_U42, P2_R1161_U420, P2_R1161_U421, P2_R1161_U422, P2_R1161_U423, P2_R1161_U424, P2_R1161_U425, P2_R1161_U426, P2_R1161_U427, P2_R1161_U428, P2_R1161_U429, P2_R1161_U43, P2_R1161_U430, P2_R1161_U431, P2_R1161_U432, P2_R1161_U433, P2_R1161_U434, P2_R1161_U435, P2_R1161_U436, P2_R1161_U437, P2_R1161_U438, P2_R1161_U439, P2_R1161_U44, P2_R1161_U440, P2_R1161_U441, P2_R1161_U442, P2_R1161_U443, P2_R1161_U444, P2_R1161_U445, P2_R1161_U446, P2_R1161_U447, P2_R1161_U448, P2_R1161_U449, P2_R1161_U45, P2_R1161_U450, P2_R1161_U451, P2_R1161_U452, P2_R1161_U453, P2_R1161_U454, P2_R1161_U455, P2_R1161_U456, P2_R1161_U457, P2_R1161_U458, P2_R1161_U459, P2_R1161_U46, P2_R1161_U460, P2_R1161_U461, P2_R1161_U462, P2_R1161_U463, P2_R1161_U464, P2_R1161_U465, P2_R1161_U466, P2_R1161_U467, P2_R1161_U468, P2_R1161_U469, P2_R1161_U47, P2_R1161_U470, P2_R1161_U471, P2_R1161_U472, P2_R1161_U473, P2_R1161_U474, P2_R1161_U475, P2_R1161_U476, P2_R1161_U477, P2_R1161_U478, P2_R1161_U479, P2_R1161_U48, P2_R1161_U480, P2_R1161_U481, P2_R1161_U482, P2_R1161_U483, P2_R1161_U484, P2_R1161_U485, P2_R1161_U486, P2_R1161_U487, P2_R1161_U488, P2_R1161_U489, P2_R1161_U49, P2_R1161_U490, P2_R1161_U491, P2_R1161_U492, P2_R1161_U493, P2_R1161_U494, P2_R1161_U495, P2_R1161_U496, P2_R1161_U497, P2_R1161_U498, P2_R1161_U499, P2_R1161_U5, P2_R1161_U50, P2_R1161_U500, P2_R1161_U501, P2_R1161_U502, P2_R1161_U503, P2_R1161_U504, P2_R1161_U51, P2_R1161_U52, P2_R1161_U53, P2_R1161_U54, P2_R1161_U55, P2_R1161_U56, P2_R1161_U57, P2_R1161_U58, P2_R1161_U59, P2_R1161_U6, P2_R1161_U60, P2_R1161_U61, P2_R1161_U62, P2_R1161_U63, P2_R1161_U64, P2_R1161_U65, P2_R1161_U66, P2_R1161_U67, P2_R1161_U68, P2_R1161_U69, P2_R1161_U7, P2_R1161_U70, P2_R1161_U71, P2_R1161_U72, P2_R1161_U73, P2_R1161_U74, P2_R1161_U75, P2_R1161_U76, P2_R1161_U77, P2_R1161_U78, P2_R1161_U79, P2_R1161_U8, P2_R1161_U80, P2_R1161_U81, P2_R1161_U82, P2_R1161_U83, P2_R1161_U84, P2_R1161_U85, P2_R1161_U86, P2_R1161_U87, P2_R1161_U88, P2_R1161_U89, P2_R1161_U9, P2_R1161_U90, P2_R1161_U91, P2_R1161_U92, P2_R1161_U93, P2_R1161_U94, P2_R1161_U95, P2_R1161_U96, P2_R1161_U97, P2_R1161_U98, P2_R1161_U99, P2_R1179_U10, P2_R1179_U100, P2_R1179_U101, P2_R1179_U102, P2_R1179_U103, P2_R1179_U104, P2_R1179_U105, P2_R1179_U106, P2_R1179_U107, P2_R1179_U108, P2_R1179_U109, P2_R1179_U11, P2_R1179_U110, P2_R1179_U111, P2_R1179_U112, P2_R1179_U113, P2_R1179_U114, P2_R1179_U115, P2_R1179_U116, P2_R1179_U117, P2_R1179_U118, P2_R1179_U119, P2_R1179_U12, P2_R1179_U120, P2_R1179_U121, P2_R1179_U122, P2_R1179_U123, P2_R1179_U124, P2_R1179_U125, P2_R1179_U126, P2_R1179_U127, P2_R1179_U128, P2_R1179_U129, P2_R1179_U13, P2_R1179_U130, P2_R1179_U131, P2_R1179_U132, P2_R1179_U133, P2_R1179_U134, P2_R1179_U135, P2_R1179_U136, P2_R1179_U137, P2_R1179_U138, P2_R1179_U139, P2_R1179_U14, P2_R1179_U140, P2_R1179_U141, P2_R1179_U142, P2_R1179_U143, P2_R1179_U144, P2_R1179_U145, P2_R1179_U146, P2_R1179_U147, P2_R1179_U148, P2_R1179_U149, P2_R1179_U15, P2_R1179_U150, P2_R1179_U151, P2_R1179_U152, P2_R1179_U153, P2_R1179_U154, P2_R1179_U155, P2_R1179_U156, P2_R1179_U157, P2_R1179_U158, P2_R1179_U159, P2_R1179_U16, P2_R1179_U160, P2_R1179_U161, P2_R1179_U162, P2_R1179_U163, P2_R1179_U164, P2_R1179_U165, P2_R1179_U166, P2_R1179_U167, P2_R1179_U168, P2_R1179_U169, P2_R1179_U17, P2_R1179_U170, P2_R1179_U171, P2_R1179_U172, P2_R1179_U173, P2_R1179_U174, P2_R1179_U175, P2_R1179_U176, P2_R1179_U177, P2_R1179_U178, P2_R1179_U179, P2_R1179_U18, P2_R1179_U180, P2_R1179_U181, P2_R1179_U182, P2_R1179_U183, P2_R1179_U184, P2_R1179_U185, P2_R1179_U186, P2_R1179_U187, P2_R1179_U188, P2_R1179_U189, P2_R1179_U19, P2_R1179_U190, P2_R1179_U191, P2_R1179_U192, P2_R1179_U193, P2_R1179_U194, P2_R1179_U195, P2_R1179_U196, P2_R1179_U197, P2_R1179_U198, P2_R1179_U199, P2_R1179_U20, P2_R1179_U200, P2_R1179_U201, P2_R1179_U202, P2_R1179_U203, P2_R1179_U204, P2_R1179_U205, P2_R1179_U206, P2_R1179_U207, P2_R1179_U208, P2_R1179_U209, P2_R1179_U21, P2_R1179_U210, P2_R1179_U211, P2_R1179_U212, P2_R1179_U213, P2_R1179_U214, P2_R1179_U215, P2_R1179_U216, P2_R1179_U217, P2_R1179_U218, P2_R1179_U219, P2_R1179_U22, P2_R1179_U220, P2_R1179_U221, P2_R1179_U222, P2_R1179_U223, P2_R1179_U224, P2_R1179_U225, P2_R1179_U226, P2_R1179_U227, P2_R1179_U228, P2_R1179_U229, P2_R1179_U23, P2_R1179_U230, P2_R1179_U231, P2_R1179_U232, P2_R1179_U233, P2_R1179_U234, P2_R1179_U235, P2_R1179_U236, P2_R1179_U237, P2_R1179_U238, P2_R1179_U239, P2_R1179_U24, P2_R1179_U240, P2_R1179_U241, P2_R1179_U242, P2_R1179_U243, P2_R1179_U244, P2_R1179_U245, P2_R1179_U246, P2_R1179_U247, P2_R1179_U248, P2_R1179_U249, P2_R1179_U25, P2_R1179_U250, P2_R1179_U251, P2_R1179_U252, P2_R1179_U253, P2_R1179_U254, P2_R1179_U255, P2_R1179_U256, P2_R1179_U257, P2_R1179_U258, P2_R1179_U259, P2_R1179_U26, P2_R1179_U260, P2_R1179_U261, P2_R1179_U262, P2_R1179_U263, P2_R1179_U264, P2_R1179_U265, P2_R1179_U266, P2_R1179_U267, P2_R1179_U268, P2_R1179_U269, P2_R1179_U27, P2_R1179_U270, P2_R1179_U271, P2_R1179_U272, P2_R1179_U273, P2_R1179_U274, P2_R1179_U275, P2_R1179_U276, P2_R1179_U277, P2_R1179_U278, P2_R1179_U279, P2_R1179_U28, P2_R1179_U280, P2_R1179_U281, P2_R1179_U282, P2_R1179_U283, P2_R1179_U284, P2_R1179_U285, P2_R1179_U286, P2_R1179_U287, P2_R1179_U288, P2_R1179_U289, P2_R1179_U29, P2_R1179_U290, P2_R1179_U291, P2_R1179_U292, P2_R1179_U293, P2_R1179_U294, P2_R1179_U295, P2_R1179_U296, P2_R1179_U297, P2_R1179_U298, P2_R1179_U299, P2_R1179_U30, P2_R1179_U300, P2_R1179_U301, P2_R1179_U302, P2_R1179_U303, P2_R1179_U304, P2_R1179_U305, P2_R1179_U306, P2_R1179_U307, P2_R1179_U308, P2_R1179_U309, P2_R1179_U31, P2_R1179_U310, P2_R1179_U311, P2_R1179_U312, P2_R1179_U313, P2_R1179_U314, P2_R1179_U315, P2_R1179_U316, P2_R1179_U317, P2_R1179_U318, P2_R1179_U319, P2_R1179_U32, P2_R1179_U320, P2_R1179_U321, P2_R1179_U322, P2_R1179_U323, P2_R1179_U324, P2_R1179_U325, P2_R1179_U326, P2_R1179_U327, P2_R1179_U328, P2_R1179_U329, P2_R1179_U33, P2_R1179_U330, P2_R1179_U331, P2_R1179_U332, P2_R1179_U333, P2_R1179_U334, P2_R1179_U335, P2_R1179_U336, P2_R1179_U337, P2_R1179_U338, P2_R1179_U339, P2_R1179_U34, P2_R1179_U340, P2_R1179_U341, P2_R1179_U342, P2_R1179_U343, P2_R1179_U344, P2_R1179_U345, P2_R1179_U346, P2_R1179_U347, P2_R1179_U348, P2_R1179_U349, P2_R1179_U35, P2_R1179_U350, P2_R1179_U351, P2_R1179_U352, P2_R1179_U353, P2_R1179_U354, P2_R1179_U355, P2_R1179_U356, P2_R1179_U357, P2_R1179_U358, P2_R1179_U359, P2_R1179_U36, P2_R1179_U360, P2_R1179_U361, P2_R1179_U362, P2_R1179_U363, P2_R1179_U364, P2_R1179_U365, P2_R1179_U366, P2_R1179_U367, P2_R1179_U368, P2_R1179_U369, P2_R1179_U37, P2_R1179_U370, P2_R1179_U371, P2_R1179_U372, P2_R1179_U373, P2_R1179_U374, P2_R1179_U375, P2_R1179_U376, P2_R1179_U377, P2_R1179_U378, P2_R1179_U379, P2_R1179_U38, P2_R1179_U380, P2_R1179_U381, P2_R1179_U382, P2_R1179_U383, P2_R1179_U384, P2_R1179_U385, P2_R1179_U386, P2_R1179_U387, P2_R1179_U388, P2_R1179_U389, P2_R1179_U39, P2_R1179_U390, P2_R1179_U391, P2_R1179_U392, P2_R1179_U393, P2_R1179_U394, P2_R1179_U395, P2_R1179_U396, P2_R1179_U397, P2_R1179_U398, P2_R1179_U399, P2_R1179_U40, P2_R1179_U400, P2_R1179_U401, P2_R1179_U402, P2_R1179_U403, P2_R1179_U404, P2_R1179_U405, P2_R1179_U406, P2_R1179_U407, P2_R1179_U408, P2_R1179_U409, P2_R1179_U41, P2_R1179_U410, P2_R1179_U411, P2_R1179_U412, P2_R1179_U413, P2_R1179_U414, P2_R1179_U415, P2_R1179_U416, P2_R1179_U417, P2_R1179_U418, P2_R1179_U419, P2_R1179_U42, P2_R1179_U420, P2_R1179_U421, P2_R1179_U422, P2_R1179_U423, P2_R1179_U424, P2_R1179_U425, P2_R1179_U426, P2_R1179_U427, P2_R1179_U428, P2_R1179_U429, P2_R1179_U43, P2_R1179_U430, P2_R1179_U431, P2_R1179_U432, P2_R1179_U433, P2_R1179_U434, P2_R1179_U435, P2_R1179_U436, P2_R1179_U437, P2_R1179_U438, P2_R1179_U439, P2_R1179_U44, P2_R1179_U440, P2_R1179_U441, P2_R1179_U442, P2_R1179_U443, P2_R1179_U444, P2_R1179_U445, P2_R1179_U446, P2_R1179_U447, P2_R1179_U448, P2_R1179_U449, P2_R1179_U45, P2_R1179_U450, P2_R1179_U451, P2_R1179_U452, P2_R1179_U453, P2_R1179_U454, P2_R1179_U455, P2_R1179_U456, P2_R1179_U457, P2_R1179_U458, P2_R1179_U459, P2_R1179_U46, P2_R1179_U460, P2_R1179_U461, P2_R1179_U462, P2_R1179_U463, P2_R1179_U464, P2_R1179_U465, P2_R1179_U466, P2_R1179_U467, P2_R1179_U468, P2_R1179_U469, P2_R1179_U47, P2_R1179_U470, P2_R1179_U471, P2_R1179_U472, P2_R1179_U473, P2_R1179_U474, P2_R1179_U475, P2_R1179_U476, P2_R1179_U477, P2_R1179_U478, P2_R1179_U479, P2_R1179_U48, P2_R1179_U480, P2_R1179_U481, P2_R1179_U482, P2_R1179_U483, P2_R1179_U484, P2_R1179_U485, P2_R1179_U486, P2_R1179_U487, P2_R1179_U488, P2_R1179_U489, P2_R1179_U49, P2_R1179_U50, P2_R1179_U51, P2_R1179_U52, P2_R1179_U53, P2_R1179_U54, P2_R1179_U55, P2_R1179_U56, P2_R1179_U57, P2_R1179_U58, P2_R1179_U59, P2_R1179_U6, P2_R1179_U60, P2_R1179_U61, P2_R1179_U62, P2_R1179_U63, P2_R1179_U64, P2_R1179_U65, P2_R1179_U66, P2_R1179_U67, P2_R1179_U68, P2_R1179_U69, P2_R1179_U7, P2_R1179_U70, P2_R1179_U71, P2_R1179_U72, P2_R1179_U73, P2_R1179_U74, P2_R1179_U75, P2_R1179_U76, P2_R1179_U77, P2_R1179_U78, P2_R1179_U79, P2_R1179_U8, P2_R1179_U80, P2_R1179_U81, P2_R1179_U82, P2_R1179_U83, P2_R1179_U84, P2_R1179_U85, P2_R1179_U86, P2_R1179_U87, P2_R1179_U88, P2_R1179_U89, P2_R1179_U9, P2_R1179_U90, P2_R1179_U91, P2_R1179_U92, P2_R1179_U93, P2_R1179_U94, P2_R1179_U95, P2_R1179_U96, P2_R1179_U97, P2_R1179_U98, P2_R1179_U99, P2_R1200_U10, P2_R1200_U100, P2_R1200_U101, P2_R1200_U102, P2_R1200_U103, P2_R1200_U104, P2_R1200_U105, P2_R1200_U106, P2_R1200_U107, P2_R1200_U108, P2_R1200_U109, P2_R1200_U11, P2_R1200_U110, P2_R1200_U111, P2_R1200_U112, P2_R1200_U113, P2_R1200_U114, P2_R1200_U115, P2_R1200_U116, P2_R1200_U117, P2_R1200_U118, P2_R1200_U119, P2_R1200_U12, P2_R1200_U120, P2_R1200_U121, P2_R1200_U122, P2_R1200_U123, P2_R1200_U124, P2_R1200_U125, P2_R1200_U126, P2_R1200_U127, P2_R1200_U128, P2_R1200_U129, P2_R1200_U13, P2_R1200_U130, P2_R1200_U131, P2_R1200_U132, P2_R1200_U133, P2_R1200_U134, P2_R1200_U135, P2_R1200_U136, P2_R1200_U137, P2_R1200_U138, P2_R1200_U139, P2_R1200_U14, P2_R1200_U140, P2_R1200_U141, P2_R1200_U142, P2_R1200_U143, P2_R1200_U144, P2_R1200_U145, P2_R1200_U146, P2_R1200_U147, P2_R1200_U148, P2_R1200_U149, P2_R1200_U15, P2_R1200_U150, P2_R1200_U151, P2_R1200_U152, P2_R1200_U153, P2_R1200_U154, P2_R1200_U155, P2_R1200_U156, P2_R1200_U157, P2_R1200_U158, P2_R1200_U159, P2_R1200_U16, P2_R1200_U160, P2_R1200_U161, P2_R1200_U162, P2_R1200_U163, P2_R1200_U164, P2_R1200_U165, P2_R1200_U166, P2_R1200_U167, P2_R1200_U168, P2_R1200_U169, P2_R1200_U17, P2_R1200_U170, P2_R1200_U171, P2_R1200_U172, P2_R1200_U173, P2_R1200_U174, P2_R1200_U175, P2_R1200_U176, P2_R1200_U177, P2_R1200_U178, P2_R1200_U179, P2_R1200_U18, P2_R1200_U180, P2_R1200_U181, P2_R1200_U182, P2_R1200_U183, P2_R1200_U184, P2_R1200_U185, P2_R1200_U186, P2_R1200_U187, P2_R1200_U188, P2_R1200_U189, P2_R1200_U19, P2_R1200_U190, P2_R1200_U191, P2_R1200_U192, P2_R1200_U193, P2_R1200_U194, P2_R1200_U195, P2_R1200_U196, P2_R1200_U197, P2_R1200_U198, P2_R1200_U199, P2_R1200_U20, P2_R1200_U200, P2_R1200_U201, P2_R1200_U202, P2_R1200_U203, P2_R1200_U204, P2_R1200_U205, P2_R1200_U206, P2_R1200_U207, P2_R1200_U208, P2_R1200_U209, P2_R1200_U21, P2_R1200_U210, P2_R1200_U211, P2_R1200_U212, P2_R1200_U213, P2_R1200_U214, P2_R1200_U215, P2_R1200_U216, P2_R1200_U217, P2_R1200_U218, P2_R1200_U219, P2_R1200_U22, P2_R1200_U220, P2_R1200_U221, P2_R1200_U222, P2_R1200_U223, P2_R1200_U224, P2_R1200_U225, P2_R1200_U226, P2_R1200_U227, P2_R1200_U228, P2_R1200_U229, P2_R1200_U23, P2_R1200_U230, P2_R1200_U231, P2_R1200_U232, P2_R1200_U233, P2_R1200_U234, P2_R1200_U235, P2_R1200_U236, P2_R1200_U237, P2_R1200_U238, P2_R1200_U239, P2_R1200_U24, P2_R1200_U240, P2_R1200_U241, P2_R1200_U242, P2_R1200_U243, P2_R1200_U244, P2_R1200_U245, P2_R1200_U246, P2_R1200_U247, P2_R1200_U248, P2_R1200_U249, P2_R1200_U25, P2_R1200_U250, P2_R1200_U251, P2_R1200_U252, P2_R1200_U253, P2_R1200_U254, P2_R1200_U255, P2_R1200_U256, P2_R1200_U257, P2_R1200_U258, P2_R1200_U259, P2_R1200_U26, P2_R1200_U260, P2_R1200_U261, P2_R1200_U262, P2_R1200_U263, P2_R1200_U264, P2_R1200_U265, P2_R1200_U266, P2_R1200_U267, P2_R1200_U268, P2_R1200_U269, P2_R1200_U27, P2_R1200_U270, P2_R1200_U271, P2_R1200_U272, P2_R1200_U273, P2_R1200_U274, P2_R1200_U275, P2_R1200_U276, P2_R1200_U277, P2_R1200_U278, P2_R1200_U279, P2_R1200_U28, P2_R1200_U280, P2_R1200_U281, P2_R1200_U282, P2_R1200_U283, P2_R1200_U284, P2_R1200_U285, P2_R1200_U286, P2_R1200_U287, P2_R1200_U288, P2_R1200_U289, P2_R1200_U29, P2_R1200_U290, P2_R1200_U291, P2_R1200_U292, P2_R1200_U293, P2_R1200_U294, P2_R1200_U295, P2_R1200_U296, P2_R1200_U297, P2_R1200_U298, P2_R1200_U299, P2_R1200_U30, P2_R1200_U300, P2_R1200_U301, P2_R1200_U302, P2_R1200_U303, P2_R1200_U304, P2_R1200_U305, P2_R1200_U306, P2_R1200_U307, P2_R1200_U308, P2_R1200_U309, P2_R1200_U31, P2_R1200_U310, P2_R1200_U311, P2_R1200_U312, P2_R1200_U313, P2_R1200_U314, P2_R1200_U315, P2_R1200_U316, P2_R1200_U317, P2_R1200_U318, P2_R1200_U319, P2_R1200_U32, P2_R1200_U320, P2_R1200_U321, P2_R1200_U322, P2_R1200_U323, P2_R1200_U324, P2_R1200_U325, P2_R1200_U326, P2_R1200_U327, P2_R1200_U328, P2_R1200_U329, P2_R1200_U33, P2_R1200_U330, P2_R1200_U331, P2_R1200_U332, P2_R1200_U333, P2_R1200_U334, P2_R1200_U335, P2_R1200_U336, P2_R1200_U337, P2_R1200_U338, P2_R1200_U339, P2_R1200_U34, P2_R1200_U340, P2_R1200_U341, P2_R1200_U342, P2_R1200_U343, P2_R1200_U344, P2_R1200_U345, P2_R1200_U346, P2_R1200_U347, P2_R1200_U348, P2_R1200_U349, P2_R1200_U35, P2_R1200_U350, P2_R1200_U351, P2_R1200_U352, P2_R1200_U353, P2_R1200_U354, P2_R1200_U355, P2_R1200_U356, P2_R1200_U357, P2_R1200_U358, P2_R1200_U359, P2_R1200_U36, P2_R1200_U360, P2_R1200_U361, P2_R1200_U362, P2_R1200_U363, P2_R1200_U364, P2_R1200_U365, P2_R1200_U366, P2_R1200_U367, P2_R1200_U368, P2_R1200_U369, P2_R1200_U37, P2_R1200_U370, P2_R1200_U371, P2_R1200_U372, P2_R1200_U373, P2_R1200_U374, P2_R1200_U375, P2_R1200_U376, P2_R1200_U377, P2_R1200_U378, P2_R1200_U379, P2_R1200_U38, P2_R1200_U380, P2_R1200_U381, P2_R1200_U382, P2_R1200_U383, P2_R1200_U384, P2_R1200_U385, P2_R1200_U386, P2_R1200_U387, P2_R1200_U388, P2_R1200_U389, P2_R1200_U39, P2_R1200_U390, P2_R1200_U391, P2_R1200_U392, P2_R1200_U393, P2_R1200_U394, P2_R1200_U395, P2_R1200_U396, P2_R1200_U397, P2_R1200_U398, P2_R1200_U399, P2_R1200_U40, P2_R1200_U400, P2_R1200_U401, P2_R1200_U402, P2_R1200_U403, P2_R1200_U404, P2_R1200_U405, P2_R1200_U406, P2_R1200_U407, P2_R1200_U408, P2_R1200_U409, P2_R1200_U41, P2_R1200_U410, P2_R1200_U411, P2_R1200_U412, P2_R1200_U413, P2_R1200_U414, P2_R1200_U415, P2_R1200_U416, P2_R1200_U417, P2_R1200_U418, P2_R1200_U419, P2_R1200_U42, P2_R1200_U420, P2_R1200_U421, P2_R1200_U422, P2_R1200_U423, P2_R1200_U424, P2_R1200_U425, P2_R1200_U426, P2_R1200_U427, P2_R1200_U428, P2_R1200_U429, P2_R1200_U43, P2_R1200_U430, P2_R1200_U431, P2_R1200_U432, P2_R1200_U433, P2_R1200_U434, P2_R1200_U435, P2_R1200_U436, P2_R1200_U437, P2_R1200_U438, P2_R1200_U439, P2_R1200_U44, P2_R1200_U440, P2_R1200_U441, P2_R1200_U442, P2_R1200_U443, P2_R1200_U444, P2_R1200_U445, P2_R1200_U446, P2_R1200_U447, P2_R1200_U448, P2_R1200_U449, P2_R1200_U45, P2_R1200_U450, P2_R1200_U451, P2_R1200_U452, P2_R1200_U453, P2_R1200_U454, P2_R1200_U455, P2_R1200_U456, P2_R1200_U457, P2_R1200_U458, P2_R1200_U459, P2_R1200_U46, P2_R1200_U460, P2_R1200_U461, P2_R1200_U462, P2_R1200_U463, P2_R1200_U464, P2_R1200_U465, P2_R1200_U466, P2_R1200_U467, P2_R1200_U468, P2_R1200_U469, P2_R1200_U47, P2_R1200_U470, P2_R1200_U471, P2_R1200_U472, P2_R1200_U473, P2_R1200_U474, P2_R1200_U475, P2_R1200_U476, P2_R1200_U477, P2_R1200_U478, P2_R1200_U479, P2_R1200_U48, P2_R1200_U480, P2_R1200_U481, P2_R1200_U482, P2_R1200_U483, P2_R1200_U484, P2_R1200_U485, P2_R1200_U486, P2_R1200_U487, P2_R1200_U488, P2_R1200_U489, P2_R1200_U49, P2_R1200_U50, P2_R1200_U51, P2_R1200_U52, P2_R1200_U53, P2_R1200_U54, P2_R1200_U55, P2_R1200_U56, P2_R1200_U57, P2_R1200_U58, P2_R1200_U59, P2_R1200_U6, P2_R1200_U60, P2_R1200_U61, P2_R1200_U62, P2_R1200_U63, P2_R1200_U64, P2_R1200_U65, P2_R1200_U66, P2_R1200_U67, P2_R1200_U68, P2_R1200_U69, P2_R1200_U7, P2_R1200_U70, P2_R1200_U71, P2_R1200_U72, P2_R1200_U73, P2_R1200_U74, P2_R1200_U75, P2_R1200_U76, P2_R1200_U77, P2_R1200_U78, P2_R1200_U79, P2_R1200_U8, P2_R1200_U80, P2_R1200_U81, P2_R1200_U82, P2_R1200_U83, P2_R1200_U84, P2_R1200_U85, P2_R1200_U86, P2_R1200_U87, P2_R1200_U88, P2_R1200_U89, P2_R1200_U9, P2_R1200_U90, P2_R1200_U91, P2_R1200_U92, P2_R1200_U93, P2_R1200_U94, P2_R1200_U95, P2_R1200_U96, P2_R1200_U97, P2_R1200_U98, P2_R1200_U99, P2_R1209_U10, P2_R1209_U100, P2_R1209_U101, P2_R1209_U102, P2_R1209_U103, P2_R1209_U104, P2_R1209_U105, P2_R1209_U106, P2_R1209_U107, P2_R1209_U108, P2_R1209_U109, P2_R1209_U11, P2_R1209_U110, P2_R1209_U111, P2_R1209_U112, P2_R1209_U113, P2_R1209_U114, P2_R1209_U115, P2_R1209_U116, P2_R1209_U117, P2_R1209_U118, P2_R1209_U119, P2_R1209_U12, P2_R1209_U120, P2_R1209_U121, P2_R1209_U122, P2_R1209_U123, P2_R1209_U124, P2_R1209_U125, P2_R1209_U126, P2_R1209_U127, P2_R1209_U128, P2_R1209_U129, P2_R1209_U13, P2_R1209_U130, P2_R1209_U131, P2_R1209_U132, P2_R1209_U133, P2_R1209_U134, P2_R1209_U135, P2_R1209_U136, P2_R1209_U137, P2_R1209_U138, P2_R1209_U139, P2_R1209_U14, P2_R1209_U140, P2_R1209_U141, P2_R1209_U142, P2_R1209_U143, P2_R1209_U144, P2_R1209_U145, P2_R1209_U146, P2_R1209_U147, P2_R1209_U148, P2_R1209_U149, P2_R1209_U15, P2_R1209_U150, P2_R1209_U151, P2_R1209_U152, P2_R1209_U153, P2_R1209_U154, P2_R1209_U155, P2_R1209_U156, P2_R1209_U157, P2_R1209_U158, P2_R1209_U159, P2_R1209_U16, P2_R1209_U160, P2_R1209_U161, P2_R1209_U162, P2_R1209_U163, P2_R1209_U164, P2_R1209_U165, P2_R1209_U166, P2_R1209_U167, P2_R1209_U168, P2_R1209_U169, P2_R1209_U17, P2_R1209_U170, P2_R1209_U171, P2_R1209_U172, P2_R1209_U173, P2_R1209_U174, P2_R1209_U175, P2_R1209_U176, P2_R1209_U177, P2_R1209_U178, P2_R1209_U179, P2_R1209_U18, P2_R1209_U180, P2_R1209_U181, P2_R1209_U182, P2_R1209_U183, P2_R1209_U184, P2_R1209_U185, P2_R1209_U186, P2_R1209_U187, P2_R1209_U188, P2_R1209_U189, P2_R1209_U19, P2_R1209_U190, P2_R1209_U191, P2_R1209_U192, P2_R1209_U193, P2_R1209_U194, P2_R1209_U195, P2_R1209_U196, P2_R1209_U197, P2_R1209_U198, P2_R1209_U199, P2_R1209_U20, P2_R1209_U200, P2_R1209_U201, P2_R1209_U202, P2_R1209_U203, P2_R1209_U204, P2_R1209_U205, P2_R1209_U206, P2_R1209_U207, P2_R1209_U208, P2_R1209_U209, P2_R1209_U21, P2_R1209_U210, P2_R1209_U211, P2_R1209_U212, P2_R1209_U213, P2_R1209_U214, P2_R1209_U215, P2_R1209_U216, P2_R1209_U217, P2_R1209_U218, P2_R1209_U219, P2_R1209_U22, P2_R1209_U220, P2_R1209_U221, P2_R1209_U222, P2_R1209_U223, P2_R1209_U224, P2_R1209_U225, P2_R1209_U226, P2_R1209_U227, P2_R1209_U228, P2_R1209_U229, P2_R1209_U23, P2_R1209_U230, P2_R1209_U231, P2_R1209_U232, P2_R1209_U233, P2_R1209_U234, P2_R1209_U235, P2_R1209_U236, P2_R1209_U237, P2_R1209_U238, P2_R1209_U239, P2_R1209_U24, P2_R1209_U240, P2_R1209_U241, P2_R1209_U242, P2_R1209_U243, P2_R1209_U244, P2_R1209_U245, P2_R1209_U246, P2_R1209_U247, P2_R1209_U248, P2_R1209_U249, P2_R1209_U25, P2_R1209_U250, P2_R1209_U251, P2_R1209_U252, P2_R1209_U253, P2_R1209_U254, P2_R1209_U255, P2_R1209_U256, P2_R1209_U257, P2_R1209_U258, P2_R1209_U259, P2_R1209_U26, P2_R1209_U260, P2_R1209_U261, P2_R1209_U262, P2_R1209_U263, P2_R1209_U264, P2_R1209_U265, P2_R1209_U266, P2_R1209_U267, P2_R1209_U268, P2_R1209_U269, P2_R1209_U27, P2_R1209_U270, P2_R1209_U271, P2_R1209_U272, P2_R1209_U273, P2_R1209_U274, P2_R1209_U275, P2_R1209_U276, P2_R1209_U28, P2_R1209_U29, P2_R1209_U30, P2_R1209_U31, P2_R1209_U32, P2_R1209_U33, P2_R1209_U34, P2_R1209_U35, P2_R1209_U36, P2_R1209_U37, P2_R1209_U38, P2_R1209_U39, P2_R1209_U40, P2_R1209_U41, P2_R1209_U42, P2_R1209_U43, P2_R1209_U44, P2_R1209_U45, P2_R1209_U46, P2_R1209_U47, P2_R1209_U48, P2_R1209_U49, P2_R1209_U50, P2_R1209_U51, P2_R1209_U52, P2_R1209_U53, P2_R1209_U54, P2_R1209_U55, P2_R1209_U56, P2_R1209_U57, P2_R1209_U58, P2_R1209_U59, P2_R1209_U6, P2_R1209_U60, P2_R1209_U61, P2_R1209_U62, P2_R1209_U63, P2_R1209_U64, P2_R1209_U65, P2_R1209_U66, P2_R1209_U67, P2_R1209_U68, P2_R1209_U69, P2_R1209_U7, P2_R1209_U70, P2_R1209_U71, P2_R1209_U72, P2_R1209_U73, P2_R1209_U74, P2_R1209_U75, P2_R1209_U76, P2_R1209_U77, P2_R1209_U78, P2_R1209_U79, P2_R1209_U8, P2_R1209_U80, P2_R1209_U81, P2_R1209_U82, P2_R1209_U83, P2_R1209_U84, P2_R1209_U85, P2_R1209_U86, P2_R1209_U87, P2_R1209_U88, P2_R1209_U89, P2_R1209_U9, P2_R1209_U90, P2_R1209_U91, P2_R1209_U92, P2_R1209_U93, P2_R1209_U94, P2_R1209_U95, P2_R1209_U96, P2_R1209_U97, P2_R1209_U98, P2_R1209_U99, P2_R1212_U10, P2_R1212_U100, P2_R1212_U101, P2_R1212_U102, P2_R1212_U103, P2_R1212_U104, P2_R1212_U105, P2_R1212_U106, P2_R1212_U107, P2_R1212_U108, P2_R1212_U109, P2_R1212_U11, P2_R1212_U110, P2_R1212_U111, P2_R1212_U112, P2_R1212_U113, P2_R1212_U114, P2_R1212_U115, P2_R1212_U116, P2_R1212_U117, P2_R1212_U118, P2_R1212_U119, P2_R1212_U12, P2_R1212_U120, P2_R1212_U121, P2_R1212_U122, P2_R1212_U123, P2_R1212_U124, P2_R1212_U125, P2_R1212_U126, P2_R1212_U127, P2_R1212_U128, P2_R1212_U129, P2_R1212_U13, P2_R1212_U130, P2_R1212_U131, P2_R1212_U132, P2_R1212_U133, P2_R1212_U134, P2_R1212_U135, P2_R1212_U136, P2_R1212_U137, P2_R1212_U138, P2_R1212_U139, P2_R1212_U14, P2_R1212_U140, P2_R1212_U141, P2_R1212_U142, P2_R1212_U143, P2_R1212_U144, P2_R1212_U145, P2_R1212_U146, P2_R1212_U147, P2_R1212_U148, P2_R1212_U149, P2_R1212_U15, P2_R1212_U150, P2_R1212_U151, P2_R1212_U152, P2_R1212_U153, P2_R1212_U154, P2_R1212_U155, P2_R1212_U156, P2_R1212_U157, P2_R1212_U158, P2_R1212_U159, P2_R1212_U16, P2_R1212_U160, P2_R1212_U161, P2_R1212_U162, P2_R1212_U163, P2_R1212_U164, P2_R1212_U165, P2_R1212_U166, P2_R1212_U167, P2_R1212_U168, P2_R1212_U169, P2_R1212_U17, P2_R1212_U170, P2_R1212_U171, P2_R1212_U172, P2_R1212_U173, P2_R1212_U174, P2_R1212_U175, P2_R1212_U176, P2_R1212_U177, P2_R1212_U178, P2_R1212_U179, P2_R1212_U18, P2_R1212_U180, P2_R1212_U181, P2_R1212_U182, P2_R1212_U183, P2_R1212_U184, P2_R1212_U185, P2_R1212_U186, P2_R1212_U187, P2_R1212_U188, P2_R1212_U189, P2_R1212_U19, P2_R1212_U190, P2_R1212_U191, P2_R1212_U192, P2_R1212_U193, P2_R1212_U194, P2_R1212_U195, P2_R1212_U196, P2_R1212_U197, P2_R1212_U198, P2_R1212_U199, P2_R1212_U20, P2_R1212_U200, P2_R1212_U201, P2_R1212_U202, P2_R1212_U203, P2_R1212_U204, P2_R1212_U205, P2_R1212_U206, P2_R1212_U207, P2_R1212_U208, P2_R1212_U209, P2_R1212_U21, P2_R1212_U210, P2_R1212_U211, P2_R1212_U212, P2_R1212_U213, P2_R1212_U214, P2_R1212_U215, P2_R1212_U216, P2_R1212_U217, P2_R1212_U218, P2_R1212_U219, P2_R1212_U22, P2_R1212_U220, P2_R1212_U221, P2_R1212_U222, P2_R1212_U223, P2_R1212_U224, P2_R1212_U225, P2_R1212_U226, P2_R1212_U227, P2_R1212_U228, P2_R1212_U229, P2_R1212_U23, P2_R1212_U230, P2_R1212_U231, P2_R1212_U232, P2_R1212_U233, P2_R1212_U234, P2_R1212_U235, P2_R1212_U236, P2_R1212_U237, P2_R1212_U238, P2_R1212_U239, P2_R1212_U24, P2_R1212_U240, P2_R1212_U241, P2_R1212_U242, P2_R1212_U243, P2_R1212_U244, P2_R1212_U245, P2_R1212_U246, P2_R1212_U247, P2_R1212_U248, P2_R1212_U249, P2_R1212_U25, P2_R1212_U250, P2_R1212_U251, P2_R1212_U252, P2_R1212_U253, P2_R1212_U254, P2_R1212_U255, P2_R1212_U256, P2_R1212_U257, P2_R1212_U258, P2_R1212_U259, P2_R1212_U26, P2_R1212_U260, P2_R1212_U261, P2_R1212_U262, P2_R1212_U263, P2_R1212_U264, P2_R1212_U265, P2_R1212_U266, P2_R1212_U267, P2_R1212_U268, P2_R1212_U269, P2_R1212_U27, P2_R1212_U270, P2_R1212_U271, P2_R1212_U272, P2_R1212_U273, P2_R1212_U274, P2_R1212_U275, P2_R1212_U276, P2_R1212_U28, P2_R1212_U29, P2_R1212_U30, P2_R1212_U31, P2_R1212_U32, P2_R1212_U33, P2_R1212_U34, P2_R1212_U35, P2_R1212_U36, P2_R1212_U37, P2_R1212_U38, P2_R1212_U39, P2_R1212_U40, P2_R1212_U41, P2_R1212_U42, P2_R1212_U43, P2_R1212_U44, P2_R1212_U45, P2_R1212_U46, P2_R1212_U47, P2_R1212_U48, P2_R1212_U49, P2_R1212_U50, P2_R1212_U51, P2_R1212_U52, P2_R1212_U53, P2_R1212_U54, P2_R1212_U55, P2_R1212_U56, P2_R1212_U57, P2_R1212_U58, P2_R1212_U59, P2_R1212_U6, P2_R1212_U60, P2_R1212_U61, P2_R1212_U62, P2_R1212_U63, P2_R1212_U64, P2_R1212_U65, P2_R1212_U66, P2_R1212_U67, P2_R1212_U68, P2_R1212_U69, P2_R1212_U7, P2_R1212_U70, P2_R1212_U71, P2_R1212_U72, P2_R1212_U73, P2_R1212_U74, P2_R1212_U75, P2_R1212_U76, P2_R1212_U77, P2_R1212_U78, P2_R1212_U79, P2_R1212_U8, P2_R1212_U80, P2_R1212_U81, P2_R1212_U82, P2_R1212_U83, P2_R1212_U84, P2_R1212_U85, P2_R1212_U86, P2_R1212_U87, P2_R1212_U88, P2_R1212_U89, P2_R1212_U9, P2_R1212_U90, P2_R1212_U91, P2_R1212_U92, P2_R1212_U93, P2_R1212_U94, P2_R1212_U95, P2_R1212_U96, P2_R1212_U97, P2_R1212_U98, P2_R1212_U99, P2_R1269_U10, P2_R1269_U100, P2_R1269_U101, P2_R1269_U102, P2_R1269_U103, P2_R1269_U104, P2_R1269_U105, P2_R1269_U106, P2_R1269_U107, P2_R1269_U108, P2_R1269_U109, P2_R1269_U11, P2_R1269_U110, P2_R1269_U111, P2_R1269_U112, P2_R1269_U113, P2_R1269_U114, P2_R1269_U115, P2_R1269_U116, P2_R1269_U117, P2_R1269_U118, P2_R1269_U119, P2_R1269_U12, P2_R1269_U120, P2_R1269_U121, P2_R1269_U122, P2_R1269_U123, P2_R1269_U124, P2_R1269_U125, P2_R1269_U126, P2_R1269_U127, P2_R1269_U128, P2_R1269_U129, P2_R1269_U13, P2_R1269_U130, P2_R1269_U131, P2_R1269_U132, P2_R1269_U133, P2_R1269_U134, P2_R1269_U135, P2_R1269_U136, P2_R1269_U137, P2_R1269_U138, P2_R1269_U139, P2_R1269_U14, P2_R1269_U140, P2_R1269_U141, P2_R1269_U142, P2_R1269_U143, P2_R1269_U144, P2_R1269_U145, P2_R1269_U146, P2_R1269_U147, P2_R1269_U148, P2_R1269_U149, P2_R1269_U15, P2_R1269_U150, P2_R1269_U151, P2_R1269_U152, P2_R1269_U153, P2_R1269_U154, P2_R1269_U155, P2_R1269_U156, P2_R1269_U157, P2_R1269_U158, P2_R1269_U159, P2_R1269_U16, P2_R1269_U160, P2_R1269_U161, P2_R1269_U162, P2_R1269_U163, P2_R1269_U164, P2_R1269_U165, P2_R1269_U166, P2_R1269_U167, P2_R1269_U168, P2_R1269_U169, P2_R1269_U17, P2_R1269_U170, P2_R1269_U171, P2_R1269_U172, P2_R1269_U173, P2_R1269_U174, P2_R1269_U175, P2_R1269_U176, P2_R1269_U177, P2_R1269_U178, P2_R1269_U179, P2_R1269_U18, P2_R1269_U180, P2_R1269_U181, P2_R1269_U182, P2_R1269_U183, P2_R1269_U184, P2_R1269_U185, P2_R1269_U186, P2_R1269_U187, P2_R1269_U188, P2_R1269_U189, P2_R1269_U19, P2_R1269_U190, P2_R1269_U191, P2_R1269_U192, P2_R1269_U193, P2_R1269_U194, P2_R1269_U195, P2_R1269_U196, P2_R1269_U197, P2_R1269_U198, P2_R1269_U199, P2_R1269_U20, P2_R1269_U200, P2_R1269_U201, P2_R1269_U202, P2_R1269_U203, P2_R1269_U204, P2_R1269_U205, P2_R1269_U206, P2_R1269_U207, P2_R1269_U208, P2_R1269_U209, P2_R1269_U21, P2_R1269_U22, P2_R1269_U23, P2_R1269_U24, P2_R1269_U25, P2_R1269_U26, P2_R1269_U27, P2_R1269_U28, P2_R1269_U29, P2_R1269_U30, P2_R1269_U31, P2_R1269_U32, P2_R1269_U33, P2_R1269_U34, P2_R1269_U35, P2_R1269_U36, P2_R1269_U37, P2_R1269_U38, P2_R1269_U39, P2_R1269_U40, P2_R1269_U41, P2_R1269_U42, P2_R1269_U43, P2_R1269_U44, P2_R1269_U45, P2_R1269_U46, P2_R1269_U47, P2_R1269_U48, P2_R1269_U49, P2_R1269_U50, P2_R1269_U51, P2_R1269_U52, P2_R1269_U53, P2_R1269_U54, P2_R1269_U55, P2_R1269_U56, P2_R1269_U57, P2_R1269_U58, P2_R1269_U59, P2_R1269_U6, P2_R1269_U60, P2_R1269_U61, P2_R1269_U62, P2_R1269_U63, P2_R1269_U64, P2_R1269_U65, P2_R1269_U66, P2_R1269_U67, P2_R1269_U68, P2_R1269_U69, P2_R1269_U7, P2_R1269_U70, P2_R1269_U71, P2_R1269_U72, P2_R1269_U73, P2_R1269_U74, P2_R1269_U75, P2_R1269_U76, P2_R1269_U77, P2_R1269_U78, P2_R1269_U79, P2_R1269_U8, P2_R1269_U80, P2_R1269_U81, P2_R1269_U82, P2_R1269_U83, P2_R1269_U84, P2_R1269_U85, P2_R1269_U86, P2_R1269_U87, P2_R1269_U88, P2_R1269_U89, P2_R1269_U9, P2_R1269_U90, P2_R1269_U91, P2_R1269_U92, P2_R1269_U93, P2_R1269_U94, P2_R1269_U95, P2_R1269_U96, P2_R1269_U97, P2_R1269_U98, P2_R1269_U99, P2_R1297_U6, P2_R1297_U7, P2_R1300_U10, P2_R1300_U6, P2_R1300_U7, P2_R1300_U8, P2_R1300_U9, P2_R693_U10, P2_R693_U100, P2_R693_U101, P2_R693_U102, P2_R693_U103, P2_R693_U104, P2_R693_U105, P2_R693_U106, P2_R693_U107, P2_R693_U108, P2_R693_U109, P2_R693_U11, P2_R693_U110, P2_R693_U111, P2_R693_U112, P2_R693_U113, P2_R693_U114, P2_R693_U115, P2_R693_U116, P2_R693_U117, P2_R693_U118, P2_R693_U119, P2_R693_U12, P2_R693_U120, P2_R693_U121, P2_R693_U122, P2_R693_U123, P2_R693_U124, P2_R693_U125, P2_R693_U126, P2_R693_U127, P2_R693_U128, P2_R693_U129, P2_R693_U13, P2_R693_U130, P2_R693_U131, P2_R693_U132, P2_R693_U133, P2_R693_U134, P2_R693_U135, P2_R693_U136, P2_R693_U137, P2_R693_U138, P2_R693_U139, P2_R693_U14, P2_R693_U140, P2_R693_U141, P2_R693_U142, P2_R693_U143, P2_R693_U144, P2_R693_U145, P2_R693_U146, P2_R693_U147, P2_R693_U148, P2_R693_U149, P2_R693_U15, P2_R693_U150, P2_R693_U151, P2_R693_U152, P2_R693_U153, P2_R693_U154, P2_R693_U155, P2_R693_U156, P2_R693_U157, P2_R693_U158, P2_R693_U159, P2_R693_U16, P2_R693_U160, P2_R693_U161, P2_R693_U162, P2_R693_U163, P2_R693_U164, P2_R693_U165, P2_R693_U166, P2_R693_U167, P2_R693_U168, P2_R693_U169, P2_R693_U17, P2_R693_U170, P2_R693_U171, P2_R693_U172, P2_R693_U173, P2_R693_U174, P2_R693_U175, P2_R693_U176, P2_R693_U177, P2_R693_U178, P2_R693_U179, P2_R693_U18, P2_R693_U180, P2_R693_U181, P2_R693_U182, P2_R693_U183, P2_R693_U184, P2_R693_U185, P2_R693_U186, P2_R693_U187, P2_R693_U188, P2_R693_U189, P2_R693_U19, P2_R693_U190, P2_R693_U191, P2_R693_U192, P2_R693_U193, P2_R693_U20, P2_R693_U21, P2_R693_U22, P2_R693_U23, P2_R693_U24, P2_R693_U25, P2_R693_U26, P2_R693_U27, P2_R693_U28, P2_R693_U29, P2_R693_U30, P2_R693_U31, P2_R693_U32, P2_R693_U33, P2_R693_U34, P2_R693_U35, P2_R693_U36, P2_R693_U37, P2_R693_U38, P2_R693_U39, P2_R693_U40, P2_R693_U41, P2_R693_U42, P2_R693_U43, P2_R693_U44, P2_R693_U45, P2_R693_U46, P2_R693_U47, P2_R693_U48, P2_R693_U49, P2_R693_U50, P2_R693_U51, P2_R693_U52, P2_R693_U53, P2_R693_U54, P2_R693_U55, P2_R693_U56, P2_R693_U57, P2_R693_U58, P2_R693_U59, P2_R693_U6, P2_R693_U60, P2_R693_U61, P2_R693_U62, P2_R693_U63, P2_R693_U64, P2_R693_U65, P2_R693_U66, P2_R693_U67, P2_R693_U68, P2_R693_U69, P2_R693_U7, P2_R693_U70, P2_R693_U71, P2_R693_U72, P2_R693_U73, P2_R693_U74, P2_R693_U75, P2_R693_U76, P2_R693_U77, P2_R693_U78, P2_R693_U79, P2_R693_U8, P2_R693_U80, P2_R693_U81, P2_R693_U82, P2_R693_U83, P2_R693_U84, P2_R693_U85, P2_R693_U86, P2_R693_U87, P2_R693_U88, P2_R693_U89, P2_R693_U9, P2_R693_U90, P2_R693_U91, P2_R693_U92, P2_R693_U93, P2_R693_U94, P2_R693_U95, P2_R693_U96, P2_R693_U97, P2_R693_U98, P2_R693_U99, P2_SUB_594_U10, P2_SUB_594_U100, P2_SUB_594_U101, P2_SUB_594_U102, P2_SUB_594_U103, P2_SUB_594_U104, P2_SUB_594_U105, P2_SUB_594_U106, P2_SUB_594_U107, P2_SUB_594_U108, P2_SUB_594_U109, P2_SUB_594_U11, P2_SUB_594_U110, P2_SUB_594_U111, P2_SUB_594_U112, P2_SUB_594_U113, P2_SUB_594_U114, P2_SUB_594_U115, P2_SUB_594_U116, P2_SUB_594_U117, P2_SUB_594_U118, P2_SUB_594_U119, P2_SUB_594_U12, P2_SUB_594_U120, P2_SUB_594_U121, P2_SUB_594_U122, P2_SUB_594_U123, P2_SUB_594_U124, P2_SUB_594_U125, P2_SUB_594_U126, P2_SUB_594_U127, P2_SUB_594_U128, P2_SUB_594_U129, P2_SUB_594_U13, P2_SUB_594_U130, P2_SUB_594_U131, P2_SUB_594_U132, P2_SUB_594_U133, P2_SUB_594_U134, P2_SUB_594_U135, P2_SUB_594_U136, P2_SUB_594_U137, P2_SUB_594_U138, P2_SUB_594_U139, P2_SUB_594_U14, P2_SUB_594_U140, P2_SUB_594_U141, P2_SUB_594_U142, P2_SUB_594_U143, P2_SUB_594_U144, P2_SUB_594_U145, P2_SUB_594_U146, P2_SUB_594_U147, P2_SUB_594_U148, P2_SUB_594_U149, P2_SUB_594_U15, P2_SUB_594_U150, P2_SUB_594_U151, P2_SUB_594_U152, P2_SUB_594_U153, P2_SUB_594_U154, P2_SUB_594_U155, P2_SUB_594_U156, P2_SUB_594_U157, P2_SUB_594_U158, P2_SUB_594_U16, P2_SUB_594_U17, P2_SUB_594_U18, P2_SUB_594_U19, P2_SUB_594_U20, P2_SUB_594_U21, P2_SUB_594_U22, P2_SUB_594_U23, P2_SUB_594_U24, P2_SUB_594_U25, P2_SUB_594_U26, P2_SUB_594_U27, P2_SUB_594_U28, P2_SUB_594_U29, P2_SUB_594_U30, P2_SUB_594_U31, P2_SUB_594_U32, P2_SUB_594_U33, P2_SUB_594_U34, P2_SUB_594_U35, P2_SUB_594_U36, P2_SUB_594_U37, P2_SUB_594_U38, P2_SUB_594_U39, P2_SUB_594_U40, P2_SUB_594_U41, P2_SUB_594_U42, P2_SUB_594_U43, P2_SUB_594_U44, P2_SUB_594_U45, P2_SUB_594_U46, P2_SUB_594_U47, P2_SUB_594_U48, P2_SUB_594_U49, P2_SUB_594_U50, P2_SUB_594_U51, P2_SUB_594_U52, P2_SUB_594_U53, P2_SUB_594_U54, P2_SUB_594_U55, P2_SUB_594_U56, P2_SUB_594_U57, P2_SUB_594_U58, P2_SUB_594_U59, P2_SUB_594_U6, P2_SUB_594_U60, P2_SUB_594_U61, P2_SUB_594_U62, P2_SUB_594_U63, P2_SUB_594_U64, P2_SUB_594_U65, P2_SUB_594_U66, P2_SUB_594_U67, P2_SUB_594_U68, P2_SUB_594_U69, P2_SUB_594_U7, P2_SUB_594_U70, P2_SUB_594_U71, P2_SUB_594_U72, P2_SUB_594_U73, P2_SUB_594_U74, P2_SUB_594_U75, P2_SUB_594_U76, P2_SUB_594_U77, P2_SUB_594_U78, P2_SUB_594_U79, P2_SUB_594_U8, P2_SUB_594_U80, P2_SUB_594_U81, P2_SUB_594_U82, P2_SUB_594_U83, P2_SUB_594_U84, P2_SUB_594_U85, P2_SUB_594_U86, P2_SUB_594_U87, P2_SUB_594_U88, P2_SUB_594_U89, P2_SUB_594_U9, P2_SUB_594_U90, P2_SUB_594_U91, P2_SUB_594_U92, P2_SUB_594_U93, P2_SUB_594_U94, P2_SUB_594_U95, P2_SUB_594_U96, P2_SUB_594_U97, P2_SUB_594_U98, P2_SUB_594_U99, P2_SUB_605_U10, P2_SUB_605_U100, P2_SUB_605_U101, P2_SUB_605_U102, P2_SUB_605_U103, P2_SUB_605_U104, P2_SUB_605_U105, P2_SUB_605_U106, P2_SUB_605_U107, P2_SUB_605_U108, P2_SUB_605_U109, P2_SUB_605_U11, P2_SUB_605_U110, P2_SUB_605_U111, P2_SUB_605_U112, P2_SUB_605_U113, P2_SUB_605_U12, P2_SUB_605_U13, P2_SUB_605_U14, P2_SUB_605_U15, P2_SUB_605_U16, P2_SUB_605_U17, P2_SUB_605_U18, P2_SUB_605_U19, P2_SUB_605_U20, P2_SUB_605_U21, P2_SUB_605_U22, P2_SUB_605_U23, P2_SUB_605_U24, P2_SUB_605_U25, P2_SUB_605_U26, P2_SUB_605_U27, P2_SUB_605_U28, P2_SUB_605_U29, P2_SUB_605_U30, P2_SUB_605_U31, P2_SUB_605_U32, P2_SUB_605_U33, P2_SUB_605_U34, P2_SUB_605_U35, P2_SUB_605_U36, P2_SUB_605_U37, P2_SUB_605_U38, P2_SUB_605_U39, P2_SUB_605_U40, P2_SUB_605_U41, P2_SUB_605_U42, P2_SUB_605_U43, P2_SUB_605_U44, P2_SUB_605_U45, P2_SUB_605_U46, P2_SUB_605_U47, P2_SUB_605_U48, P2_SUB_605_U49, P2_SUB_605_U50, P2_SUB_605_U51, P2_SUB_605_U52, P2_SUB_605_U53, P2_SUB_605_U54, P2_SUB_605_U55, P2_SUB_605_U56, P2_SUB_605_U57, P2_SUB_605_U58, P2_SUB_605_U59, P2_SUB_605_U6, P2_SUB_605_U60, P2_SUB_605_U61, P2_SUB_605_U62, P2_SUB_605_U63, P2_SUB_605_U64, P2_SUB_605_U65, P2_SUB_605_U66, P2_SUB_605_U67, P2_SUB_605_U68, P2_SUB_605_U69, P2_SUB_605_U7, P2_SUB_605_U70, P2_SUB_605_U71, P2_SUB_605_U72, P2_SUB_605_U73, P2_SUB_605_U74, P2_SUB_605_U75, P2_SUB_605_U76, P2_SUB_605_U77, P2_SUB_605_U78, P2_SUB_605_U79, P2_SUB_605_U8, P2_SUB_605_U80, P2_SUB_605_U81, P2_SUB_605_U82, P2_SUB_605_U83, P2_SUB_605_U84, P2_SUB_605_U85, P2_SUB_605_U86, P2_SUB_605_U87, P2_SUB_605_U88, P2_SUB_605_U89, P2_SUB_605_U9, P2_SUB_605_U90, P2_SUB_605_U91, P2_SUB_605_U92, P2_SUB_605_U93, P2_SUB_605_U94, P2_SUB_605_U95, P2_SUB_605_U96, P2_SUB_605_U97, P2_SUB_605_U98, P2_SUB_605_U99, P2_U3013, P2_U3014, P2_U3015, P2_U3016, P2_U3017, P2_U3018, P2_U3019, P2_U3020, P2_U3021, P2_U3022, P2_U3023, P2_U3024, P2_U3025, P2_U3026, P2_U3027, P2_U3028, P2_U3029, P2_U3030, P2_U3031, P2_U3032, P2_U3033, P2_U3034, P2_U3035, P2_U3036, P2_U3037, P2_U3038, P2_U3039, P2_U3040, P2_U3041, P2_U3042, P2_U3043, P2_U3044, P2_U3045, P2_U3046, P2_U3047, P2_U3048, P2_U3049, P2_U3050, P2_U3051, P2_U3052, P2_U3053, P2_U3054, P2_U3055, P2_U3056, P2_U3057, P2_U3058, P2_U3059, P2_U3060, P2_U3061, P2_U3062, P2_U3063, P2_U3064, P2_U3065, P2_U3066, P2_U3067, P2_U3068, P2_U3069, P2_U3070, P2_U3071, P2_U3072, P2_U3073, P2_U3074, P2_U3075, P2_U3076, P2_U3077, P2_U3078, P2_U3079, P2_U3080, P2_U3081, P2_U3082, P2_U3083, P2_U3084, P2_U3085, P2_U3086, P2_U3087, P2_U3088, P2_U3089, P2_U3090, P2_U3091, P2_U3092, P2_U3093, P2_U3094, P2_U3095, P2_U3096, P2_U3097, P2_U3098, P2_U3099, P2_U3100, P2_U3101, P2_U3102, P2_U3103, P2_U3104, P2_U3105, P2_U3106, P2_U3107, P2_U3108, P2_U3109, P2_U3110, P2_U3111, P2_U3112, P2_U3113, P2_U3114, P2_U3115, P2_U3116, P2_U3117, P2_U3118, P2_U3119, P2_U3120, P2_U3121, P2_U3122, P2_U3123, P2_U3124, P2_U3125, P2_U3126, P2_U3127, P2_U3128, P2_U3129, P2_U3130, P2_U3131, P2_U3132, P2_U3133, P2_U3134, P2_U3135, P2_U3136, P2_U3137, P2_U3138, P2_U3139, P2_U3140, P2_U3141, P2_U3142, P2_U3143, P2_U3144, P2_U3145, P2_U3146, P2_U3147, P2_U3148, P2_U3149, P2_U3152, P2_U3297, P2_U3298, P2_U3299, P2_U3300, P2_U3301, P2_U3302, P2_U3303, P2_U3304, P2_U3305, P2_U3306, P2_U3307, P2_U3308, P2_U3309, P2_U3310, P2_U3311, P2_U3312, P2_U3313, P2_U3314, P2_U3315, P2_U3316, P2_U3317, P2_U3318, P2_U3319, P2_U3320, P2_U3321, P2_U3322, P2_U3323, P2_U3324, P2_U3325, P2_U3326, P2_U3327, P2_U3328, P2_U3329, P2_U3330, P2_U3331, P2_U3332, P2_U3333, P2_U3334, P2_U3335, P2_U3336, P2_U3337, P2_U3338, P2_U3339, P2_U3340, P2_U3341, P2_U3342, P2_U3343, P2_U3344, P2_U3345, P2_U3346, P2_U3347, P2_U3348, P2_U3349, P2_U3350, P2_U3351, P2_U3352, P2_U3353, P2_U3354, P2_U3355, P2_U3356, P2_U3357, P2_U3358, P2_U3359, P2_U3360, P2_U3361, P2_U3362, P2_U3363, P2_U3364, P2_U3365, P2_U3366, P2_U3367, P2_U3368, P2_U3369, P2_U3370, P2_U3371, P2_U3372, P2_U3373, P2_U3374, P2_U3375, P2_U3378, P2_U3379, P2_U3380, P2_U3381, P2_U3382, P2_U3383, P2_U3384, P2_U3385, P2_U3386, P2_U3387, P2_U3388, P2_U3389, P2_U3391, P2_U3392, P2_U3394, P2_U3395, P2_U3397, P2_U3398, P2_U3400, P2_U3401, P2_U3403, P2_U3404, P2_U3406, P2_U3407, P2_U3409, P2_U3410, P2_U3412, P2_U3413, P2_U3415, P2_U3416, P2_U3418, P2_U3419, P2_U3421, P2_U3422, P2_U3424, P2_U3425, P2_U3427, P2_U3428, P2_U3430, P2_U3431, P2_U3433, P2_U3434, P2_U3436, P2_U3437, P2_U3439, P2_U3440, P2_U3442, P2_U3443, P2_U3445, P2_U3523, P2_U3524, P2_U3525, P2_U3526, P2_U3527, P2_U3528, P2_U3529, P2_U3530, P2_U3531, P2_U3532, P2_U3533, P2_U3534, P2_U3535, P2_U3536, P2_U3537, P2_U3538, P2_U3539, P2_U3540, P2_U3541, P2_U3542, P2_U3543, P2_U3544, P2_U3545, P2_U3546, P2_U3547, P2_U3548, P2_U3549, P2_U3550, P2_U3551, P2_U3552, P2_U3553, P2_U3554, P2_U3555, P2_U3556, P2_U3557, P2_U3558, P2_U3559, P2_U3560, P2_U3561, P2_U3562, P2_U3563, P2_U3564, P2_U3565, P2_U3566, P2_U3567, P2_U3568, P2_U3569, P2_U3570, P2_U3571, P2_U3572, P2_U3573, P2_U3574, P2_U3575, P2_U3576, P2_U3577, P2_U3578, P2_U3579, P2_U3580, P2_U3581, P2_U3582, P2_U3583, P2_U3584, P2_U3585, P2_U3586, P2_U3587, P2_U3588, P2_U3589, P2_U3590, P2_U3591, P2_U3592, P2_U3593, P2_U3594, P2_U3595, P2_U3596, P2_U3597, P2_U3598, P2_U3599, P2_U3600, P2_U3601, P2_U3602, P2_U3603, P2_U3604, P2_U3605, P2_U3606, P2_U3607, P2_U3608, P2_U3609, P2_U3610, P2_U3611, P2_U3612, P2_U3613, P2_U3614, P2_U3615, P2_U3616, P2_U3617, P2_U3618, P2_U3619, P2_U3620, P2_U3621, P2_U3622, P2_U3623, P2_U3624, P2_U3625, P2_U3626, P2_U3627, P2_U3628, P2_U3629, P2_U3630, P2_U3631, P2_U3632, P2_U3633, P2_U3634, P2_U3635, P2_U3636, P2_U3637, P2_U3638, P2_U3639, P2_U3640, P2_U3641, P2_U3642, P2_U3643, P2_U3644, P2_U3645, P2_U3646, P2_U3647, P2_U3648, P2_U3649, P2_U3650, P2_U3651, P2_U3652, P2_U3653, P2_U3654, P2_U3655, P2_U3656, P2_U3657, P2_U3658, P2_U3659, P2_U3660, P2_U3661, P2_U3662, P2_U3663, P2_U3664, P2_U3665, P2_U3666, P2_U3667, P2_U3668, P2_U3669, P2_U3670, P2_U3671, P2_U3672, P2_U3673, P2_U3674, P2_U3675, P2_U3676, P2_U3677, P2_U3678, P2_U3679, P2_U3680, P2_U3681, P2_U3682, P2_U3683, P2_U3684, P2_U3685, P2_U3686, P2_U3687, P2_U3688, P2_U3689, P2_U3690, P2_U3691, P2_U3692, P2_U3693, P2_U3694, P2_U3695, P2_U3696, P2_U3697, P2_U3698, P2_U3699, P2_U3700, P2_U3701, P2_U3702, P2_U3703, P2_U3704, P2_U3705, P2_U3706, P2_U3707, P2_U3708, P2_U3709, P2_U3710, P2_U3711, P2_U3712, P2_U3713, P2_U3714, P2_U3715, P2_U3716, P2_U3717, P2_U3718, P2_U3719, P2_U3720, P2_U3721, P2_U3722, P2_U3723, P2_U3724, P2_U3725, P2_U3726, P2_U3727, P2_U3728, P2_U3729, P2_U3730, P2_U3731, P2_U3732, P2_U3733, P2_U3734, P2_U3735, P2_U3736, P2_U3737, P2_U3738, P2_U3739, P2_U3740, P2_U3741, P2_U3742, P2_U3743, P2_U3744, P2_U3745, P2_U3746, P2_U3747, P2_U3748, P2_U3749, P2_U3750, P2_U3751, P2_U3752, P2_U3753, P2_U3754, P2_U3755, P2_U3756, P2_U3757, P2_U3758, P2_U3759, P2_U3760, P2_U3761, P2_U3762, P2_U3763, P2_U3764, P2_U3765, P2_U3766, P2_U3767, P2_U3768, P2_U3769, P2_U3770, P2_U3771, P2_U3772, P2_U3773, P2_U3774, P2_U3775, P2_U3776, P2_U3777, P2_U3778, P2_U3779, P2_U3780, P2_U3781, P2_U3782, P2_U3783, P2_U3784, P2_U3785, P2_U3786, P2_U3787, P2_U3788, P2_U3789, P2_U3790, P2_U3791, P2_U3792, P2_U3793, P2_U3794, P2_U3795, P2_U3796, P2_U3797, P2_U3798, P2_U3799, P2_U3800, P2_U3801, P2_U3802, P2_U3803, P2_U3804, P2_U3805, P2_U3806, P2_U3807, P2_U3808, P2_U3809, P2_U3810, P2_U3811, P2_U3812, P2_U3813, P2_U3814, P2_U3815, P2_U3816, P2_U3817, P2_U3818, P2_U3819, P2_U3820, P2_U3821, P2_U3822, P2_U3823, P2_U3824, P2_U3825, P2_U3826, P2_U3827, P2_U3828, P2_U3829, P2_U3830, P2_U3831, P2_U3832, P2_U3833, P2_U3834, P2_U3835, P2_U3836, P2_U3837, P2_U3838, P2_U3839, P2_U3840, P2_U3841, P2_U3842, P2_U3843, P2_U3844, P2_U3845, P2_U3846, P2_U3847, P2_U3848, P2_U3849, P2_U3850, P2_U3851, P2_U3852, P2_U3853, P2_U3854, P2_U3855, P2_U3856, P2_U3857, P2_U3858, P2_U3859, P2_U3860, P2_U3861, P2_U3862, P2_U3863, P2_U3864, P2_U3865, P2_U3866, P2_U3867, P2_U3868, P2_U3869, P2_U3870, P2_U3871, P2_U3872, P2_U3873, P2_U3874, P2_U3875, P2_U3876, P2_U3877, P2_U3878, P2_U3879, P2_U3880, P2_U3881, P2_U3882, P2_U3883, P2_U3884, P2_U3885, P2_U3886, P2_U3887, P2_U3888, P2_U3889, P2_U3890, P2_U3891, P2_U3892, P2_U3894, P2_U3895, P2_U3896, P2_U3897, P2_U3898, P2_U3899, P2_U3900, P2_U3901, P2_U3902, P2_U3903, P2_U3904, P2_U3905, P2_U3906, P2_U3907, P2_U3908, P2_U3909, P2_U3910, P2_U3911, P2_U3912, P2_U3913, P2_U3914, P2_U3915, P2_U3916, P2_U3917, P2_U3918, P2_U3919, P2_U3920, P2_U3921, P2_U3922, P2_U3923, P2_U3924, P2_U3925, P2_U3926, P2_U3927, P2_U3928, P2_U3929, P2_U3930, P2_U3931, P2_U3932, P2_U3933, P2_U3934, P2_U3935, P2_U3936, P2_U3937, P2_U3938, P2_U3939, P2_U3940, P2_U3941, P2_U3942, P2_U3943, P2_U3944, P2_U3945, P2_U3946, P2_U3947, P2_U3948, P2_U3949, P2_U3950, P2_U3951, P2_U3952, P2_U3953, P2_U3954, P2_U3955, P2_U3956, P2_U3957, P2_U3958, P2_U3959, P2_U3960, P2_U3961, P2_U3962, P2_U3963, P2_U3964, P2_U3965, P2_U3966, P2_U3967, P2_U3968, P2_U3969, P2_U3970, P2_U3971, P2_U3972, P2_U3973, P2_U3974, P2_U3975, P2_U3976, P2_U3977, P2_U3978, P2_U3979, P2_U3980, P2_U3981, P2_U3982, P2_U3983, P2_U3984, P2_U3985, P2_U3986, P2_U3987, P2_U3988, P2_U3989, P2_U3990, P2_U3991, P2_U3992, P2_U3993, P2_U3994, P2_U3995, P2_U3996, P2_U3997, P2_U3998, P2_U3999, P2_U4000, P2_U4001, P2_U4002, P2_U4003, P2_U4004, P2_U4005, P2_U4006, P2_U4007, P2_U4008, P2_U4009, P2_U4010, P2_U4011, P2_U4012, P2_U4013, P2_U4014, P2_U4015, P2_U4016, P2_U4017, P2_U4018, P2_U4019, P2_U4020, P2_U4021, P2_U4022, P2_U4023, P2_U4024, P2_U4025, P2_U4026, P2_U4027, P2_U4028, P2_U4029, P2_U4030, P2_U4031, P2_U4032, P2_U4033, P2_U4034, P2_U4035, P2_U4036, P2_U4037, P2_U4038, P2_U4039, P2_U4040, P2_U4041, P2_U4042, P2_U4043, P2_U4044, P2_U4045, P2_U4046, P2_U4047, P2_U4048, P2_U4049, P2_U4050, P2_U4051, P2_U4052, P2_U4053, P2_U4054, P2_U4055, P2_U4056, P2_U4057, P2_U4058, P2_U4059, P2_U4060, P2_U4061, P2_U4062, P2_U4063, P2_U4064, P2_U4065, P2_U4066, P2_U4067, P2_U4068, P2_U4069, P2_U4070, P2_U4071, P2_U4072, P2_U4073, P2_U4074, P2_U4075, P2_U4076, P2_U4077, P2_U4078, P2_U4079, P2_U4080, P2_U4081, P2_U4082, P2_U4083, P2_U4084, P2_U4085, P2_U4086, P2_U4087, P2_U4088, P2_U4089, P2_U4090, P2_U4091, P2_U4092, P2_U4093, P2_U4094, P2_U4095, P2_U4096, P2_U4097, P2_U4098, P2_U4099, P2_U4100, P2_U4101, P2_U4102, P2_U4103, P2_U4104, P2_U4105, P2_U4106, P2_U4107, P2_U4108, P2_U4109, P2_U4110, P2_U4111, P2_U4112, P2_U4113, P2_U4114, P2_U4115, P2_U4116, P2_U4117, P2_U4118, P2_U4119, P2_U4120, P2_U4121, P2_U4122, P2_U4123, P2_U4124, P2_U4125, P2_U4126, P2_U4127, P2_U4128, P2_U4129, P2_U4130, P2_U4131, P2_U4132, P2_U4133, P2_U4134, P2_U4135, P2_U4136, P2_U4137, P2_U4138, P2_U4139, P2_U4140, P2_U4141, P2_U4142, P2_U4143, P2_U4144, P2_U4145, P2_U4146, P2_U4147, P2_U4148, P2_U4149, P2_U4150, P2_U4151, P2_U4152, P2_U4153, P2_U4154, P2_U4155, P2_U4156, P2_U4157, P2_U4158, P2_U4159, P2_U4160, P2_U4161, P2_U4162, P2_U4163, P2_U4164, P2_U4165, P2_U4166, P2_U4167, P2_U4168, P2_U4169, P2_U4170, P2_U4171, P2_U4172, P2_U4173, P2_U4174, P2_U4175, P2_U4176, P2_U4177, P2_U4178, P2_U4179, P2_U4180, P2_U4181, P2_U4182, P2_U4183, P2_U4184, P2_U4185, P2_U4186, P2_U4187, P2_U4188, P2_U4189, P2_U4190, P2_U4191, P2_U4192, P2_U4193, P2_U4194, P2_U4195, P2_U4196, P2_U4197, P2_U4198, P2_U4199, P2_U4200, P2_U4201, P2_U4202, P2_U4203, P2_U4204, P2_U4205, P2_U4206, P2_U4207, P2_U4208, P2_U4209, P2_U4210, P2_U4211, P2_U4212, P2_U4213, P2_U4214, P2_U4215, P2_U4216, P2_U4217, P2_U4218, P2_U4219, P2_U4220, P2_U4221, P2_U4222, P2_U4223, P2_U4224, P2_U4225, P2_U4226, P2_U4227, P2_U4228, P2_U4229, P2_U4230, P2_U4231, P2_U4232, P2_U4233, P2_U4234, P2_U4235, P2_U4236, P2_U4237, P2_U4238, P2_U4239, P2_U4240, P2_U4241, P2_U4242, P2_U4243, P2_U4244, P2_U4245, P2_U4246, P2_U4247, P2_U4248, P2_U4249, P2_U4250, P2_U4251, P2_U4252, P2_U4253, P2_U4254, P2_U4255, P2_U4256, P2_U4257, P2_U4258, P2_U4259, P2_U4260, P2_U4261, P2_U4262, P2_U4263, P2_U4264, P2_U4265, P2_U4266, P2_U4267, P2_U4268, P2_U4269, P2_U4270, P2_U4271, P2_U4272, P2_U4273, P2_U4274, P2_U4275, P2_U4276, P2_U4277, P2_U4278, P2_U4279, P2_U4280, P2_U4281, P2_U4282, P2_U4283, P2_U4284, P2_U4285, P2_U4286, P2_U4287, P2_U4288, P2_U4289, P2_U4290, P2_U4291, P2_U4292, P2_U4293, P2_U4294, P2_U4295, P2_U4296, P2_U4297, P2_U4298, P2_U4299, P2_U4300, P2_U4301, P2_U4302, P2_U4303, P2_U4304, P2_U4305, P2_U4306, P2_U4307, P2_U4308, P2_U4309, P2_U4310, P2_U4311, P2_U4312, P2_U4313, P2_U4314, P2_U4315, P2_U4316, P2_U4317, P2_U4318, P2_U4319, P2_U4320, P2_U4321, P2_U4322, P2_U4323, P2_U4324, P2_U4325, P2_U4326, P2_U4327, P2_U4328, P2_U4329, P2_U4330, P2_U4331, P2_U4332, P2_U4333, P2_U4334, P2_U4335, P2_U4336, P2_U4337, P2_U4338, P2_U4339, P2_U4340, P2_U4341, P2_U4342, P2_U4343, P2_U4344, P2_U4345, P2_U4346, P2_U4347, P2_U4348, P2_U4349, P2_U4350, P2_U4351, P2_U4352, P2_U4353, P2_U4354, P2_U4355, P2_U4356, P2_U4357, P2_U4358, P2_U4359, P2_U4360, P2_U4361, P2_U4362, P2_U4363, P2_U4364, P2_U4365, P2_U4366, P2_U4367, P2_U4368, P2_U4369, P2_U4370, P2_U4371, P2_U4372, P2_U4373, P2_U4374, P2_U4375, P2_U4376, P2_U4377, P2_U4378, P2_U4379, P2_U4380, P2_U4381, P2_U4382, P2_U4383, P2_U4384, P2_U4385, P2_U4386, P2_U4387, P2_U4388, P2_U4389, P2_U4390, P2_U4391, P2_U4392, P2_U4393, P2_U4394, P2_U4395, P2_U4396, P2_U4397, P2_U4398, P2_U4399, P2_U4400, P2_U4401, P2_U4402, P2_U4403, P2_U4404, P2_U4405, P2_U4406, P2_U4407, P2_U4408, P2_U4409, P2_U4410, P2_U4411, P2_U4412, P2_U4413, P2_U4414, P2_U4415, P2_U4416, P2_U4417, P2_U4418, P2_U4419, P2_U4420, P2_U4421, P2_U4422, P2_U4423, P2_U4424, P2_U4425, P2_U4426, P2_U4427, P2_U4428, P2_U4429, P2_U4430, P2_U4431, P2_U4432, P2_U4433, P2_U4434, P2_U4435, P2_U4436, P2_U4437, P2_U4438, P2_U4439, P2_U4440, P2_U4441, P2_U4442, P2_U4443, P2_U4444, P2_U4445, P2_U4446, P2_U4447, P2_U4448, P2_U4449, P2_U4450, P2_U4451, P2_U4452, P2_U4453, P2_U4454, P2_U4455, P2_U4456, P2_U4457, P2_U4458, P2_U4459, P2_U4460, P2_U4461, P2_U4462, P2_U4463, P2_U4464, P2_U4465, P2_U4466, P2_U4467, P2_U4468, P2_U4469, P2_U4470, P2_U4471, P2_U4472, P2_U4473, P2_U4474, P2_U4475, P2_U4476, P2_U4477, P2_U4478, P2_U4479, P2_U4480, P2_U4481, P2_U4482, P2_U4483, P2_U4484, P2_U4485, P2_U4486, P2_U4487, P2_U4488, P2_U4489, P2_U4490, P2_U4491, P2_U4492, P2_U4493, P2_U4494, P2_U4495, P2_U4496, P2_U4497, P2_U4498, P2_U4499, P2_U4500, P2_U4501, P2_U4502, P2_U4503, P2_U4504, P2_U4505, P2_U4506, P2_U4507, P2_U4508, P2_U4509, P2_U4510, P2_U4511, P2_U4512, P2_U4513, P2_U4514, P2_U4515, P2_U4516, P2_U4517, P2_U4518, P2_U4519, P2_U4520, P2_U4521, P2_U4522, P2_U4523, P2_U4524, P2_U4525, P2_U4526, P2_U4527, P2_U4528, P2_U4529, P2_U4530, P2_U4531, P2_U4532, P2_U4533, P2_U4534, P2_U4535, P2_U4536, P2_U4537, P2_U4538, P2_U4539, P2_U4540, P2_U4541, P2_U4542, P2_U4543, P2_U4544, P2_U4545, P2_U4546, P2_U4547, P2_U4548, P2_U4549, P2_U4550, P2_U4551, P2_U4552, P2_U4553, P2_U4554, P2_U4555, P2_U4556, P2_U4557, P2_U4558, P2_U4559, P2_U4560, P2_U4561, P2_U4562, P2_U4563, P2_U4564, P2_U4565, P2_U4566, P2_U4567, P2_U4568, P2_U4569, P2_U4570, P2_U4571, P2_U4572, P2_U4573, P2_U4574, P2_U4575, P2_U4576, P2_U4577, P2_U4578, P2_U4579, P2_U4580, P2_U4581, P2_U4582, P2_U4583, P2_U4584, P2_U4585, P2_U4586, P2_U4587, P2_U4588, P2_U4589, P2_U4590, P2_U4591, P2_U4592, P2_U4593, P2_U4594, P2_U4595, P2_U4596, P2_U4597, P2_U4598, P2_U4599, P2_U4600, P2_U4601, P2_U4602, P2_U4603, P2_U4604, P2_U4605, P2_U4606, P2_U4607, P2_U4608, P2_U4609, P2_U4610, P2_U4611, P2_U4612, P2_U4613, P2_U4614, P2_U4615, P2_U4616, P2_U4617, P2_U4618, P2_U4619, P2_U4620, P2_U4621, P2_U4622, P2_U4623, P2_U4624, P2_U4625, P2_U4626, P2_U4627, P2_U4628, P2_U4629, P2_U4630, P2_U4631, P2_U4632, P2_U4633, P2_U4634, P2_U4635, P2_U4636, P2_U4637, P2_U4638, P2_U4639, P2_U4640, P2_U4641, P2_U4642, P2_U4643, P2_U4644, P2_U4645, P2_U4646, P2_U4647, P2_U4648, P2_U4649, P2_U4650, P2_U4651, P2_U4652, P2_U4653, P2_U4654, P2_U4655, P2_U4656, P2_U4657, P2_U4658, P2_U4659, P2_U4660, P2_U4661, P2_U4662, P2_U4663, P2_U4664, P2_U4665, P2_U4666, P2_U4667, P2_U4668, P2_U4669, P2_U4670, P2_U4671, P2_U4672, P2_U4673, P2_U4674, P2_U4675, P2_U4676, P2_U4677, P2_U4678, P2_U4679, P2_U4680, P2_U4681, P2_U4682, P2_U4683, P2_U4684, P2_U4685, P2_U4686, P2_U4687, P2_U4688, P2_U4689, P2_U4690, P2_U4691, P2_U4692, P2_U4693, P2_U4694, P2_U4695, P2_U4696, P2_U4697, P2_U4698, P2_U4699, P2_U4700, P2_U4701, P2_U4702, P2_U4703, P2_U4704, P2_U4705, P2_U4706, P2_U4707, P2_U4708, P2_U4709, P2_U4710, P2_U4711, P2_U4712, P2_U4713, P2_U4714, P2_U4715, P2_U4716, P2_U4717, P2_U4718, P2_U4719, P2_U4720, P2_U4721, P2_U4722, P2_U4723, P2_U4724, P2_U4725, P2_U4726, P2_U4727, P2_U4728, P2_U4729, P2_U4730, P2_U4731, P2_U4732, P2_U4733, P2_U4734, P2_U4735, P2_U4736, P2_U4737, P2_U4738, P2_U4739, P2_U4740, P2_U4741, P2_U4742, P2_U4743, P2_U4744, P2_U4745, P2_U4746, P2_U4747, P2_U4748, P2_U4749, P2_U4750, P2_U4751, P2_U4752, P2_U4753, P2_U4754, P2_U4755, P2_U4756, P2_U4757, P2_U4758, P2_U4759, P2_U4760, P2_U4761, P2_U4762, P2_U4763, P2_U4764, P2_U4765, P2_U4766, P2_U4767, P2_U4768, P2_U4769, P2_U4770, P2_U4771, P2_U4772, P2_U4773, P2_U4774, P2_U4775, P2_U4776, P2_U4777, P2_U4778, P2_U4779, P2_U4780, P2_U4781, P2_U4782, P2_U4783, P2_U4784, P2_U4785, P2_U4786, P2_U4787, P2_U4788, P2_U4789, P2_U4790, P2_U4791, P2_U4792, P2_U4793, P2_U4794, P2_U4795, P2_U4796, P2_U4797, P2_U4798, P2_U4799, P2_U4800, P2_U4801, P2_U4802, P2_U4803, P2_U4804, P2_U4805, P2_U4806, P2_U4807, P2_U4808, P2_U4809, P2_U4810, P2_U4811, P2_U4812, P2_U4813, P2_U4814, P2_U4815, P2_U4816, P2_U4817, P2_U4818, P2_U4819, P2_U4820, P2_U4821, P2_U4822, P2_U4823, P2_U4824, P2_U4825, P2_U4826, P2_U4827, P2_U4828, P2_U4829, P2_U4830, P2_U4831, P2_U4832, P2_U4833, P2_U4834, P2_U4835, P2_U4836, P2_U4837, P2_U4838, P2_U4839, P2_U4840, P2_U4841, P2_U4842, P2_U4843, P2_U4844, P2_U4845, P2_U4846, P2_U4847, P2_U4848, P2_U4849, P2_U4850, P2_U4851, P2_U4852, P2_U4853, P2_U4854, P2_U4855, P2_U4856, P2_U4857, P2_U4858, P2_U4859, P2_U4860, P2_U4861, P2_U4862, P2_U4863, P2_U4864, P2_U4865, P2_U4866, P2_U4867, P2_U4868, P2_U4869, P2_U4870, P2_U4871, P2_U4872, P2_U4873, P2_U4874, P2_U4875, P2_U4876, P2_U4877, P2_U4878, P2_U4879, P2_U4880, P2_U4881, P2_U4882, P2_U4883, P2_U4884, P2_U4885, P2_U4886, P2_U4887, P2_U4888, P2_U4889, P2_U4890, P2_U4891, P2_U4892, P2_U4893, P2_U4894, P2_U4895, P2_U4896, P2_U4897, P2_U4898, P2_U4899, P2_U4900, P2_U4901, P2_U4902, P2_U4903, P2_U4904, P2_U4905, P2_U4906, P2_U4907, P2_U4908, P2_U4909, P2_U4910, P2_U4911, P2_U4912, P2_U4913, P2_U4914, P2_U4915, P2_U4916, P2_U4917, P2_U4918, P2_U4919, P2_U4920, P2_U4921, P2_U4922, P2_U4923, P2_U4924, P2_U4925, P2_U4926, P2_U4927, P2_U4928, P2_U4929, P2_U4930, P2_U4931, P2_U4932, P2_U4933, P2_U4934, P2_U4935, P2_U4936, P2_U4937, P2_U4938, P2_U4939, P2_U4940, P2_U4941, P2_U4942, P2_U4943, P2_U4944, P2_U4945, P2_U4946, P2_U4947, P2_U4948, P2_U4949, P2_U4950, P2_U4951, P2_U4952, P2_U4953, P2_U4954, P2_U4955, P2_U4956, P2_U4957, P2_U4958, P2_U4959, P2_U4960, P2_U4961, P2_U4962, P2_U4963, P2_U4964, P2_U4965, P2_U4966, P2_U4967, P2_U4968, P2_U4969, P2_U4970, P2_U4971, P2_U4972, P2_U4973, P2_U4974, P2_U4975, P2_U4976, P2_U4977, P2_U4978, P2_U4979, P2_U4980, P2_U4981, P2_U4982, P2_U4983, P2_U4984, P2_U4985, P2_U4986, P2_U4987, P2_U4988, P2_U4989, P2_U4990, P2_U4991, P2_U4992, P2_U4993, P2_U4994, P2_U4995, P2_U4996, P2_U4997, P2_U4998, P2_U4999, P2_U5000, P2_U5001, P2_U5002, P2_U5003, P2_U5004, P2_U5005, P2_U5006, P2_U5007, P2_U5008, P2_U5009, P2_U5010, P2_U5011, P2_U5012, P2_U5013, P2_U5014, P2_U5015, P2_U5016, P2_U5017, P2_U5018, P2_U5019, P2_U5020, P2_U5021, P2_U5022, P2_U5023, P2_U5024, P2_U5025, P2_U5026, P2_U5027, P2_U5028, P2_U5029, P2_U5030, P2_U5031, P2_U5032, P2_U5033, P2_U5034, P2_U5035, P2_U5036, P2_U5037, P2_U5038, P2_U5039, P2_U5040, P2_U5041, P2_U5042, P2_U5043, P2_U5044, P2_U5045, P2_U5046, P2_U5047, P2_U5048, P2_U5049, P2_U5050, P2_U5051, P2_U5052, P2_U5053, P2_U5054, P2_U5055, P2_U5056, P2_U5057, P2_U5058, P2_U5059, P2_U5060, P2_U5061, P2_U5062, P2_U5063, P2_U5064, P2_U5065, P2_U5066, P2_U5067, P2_U5068, P2_U5069, P2_U5070, P2_U5071, P2_U5072, P2_U5073, P2_U5074, P2_U5075, P2_U5076, P2_U5077, P2_U5078, P2_U5079, P2_U5080, P2_U5081, P2_U5082, P2_U5083, P2_U5084, P2_U5085, P2_U5086, P2_U5087, P2_U5088, P2_U5089, P2_U5090, P2_U5091, P2_U5092, P2_U5093, P2_U5094, P2_U5095, P2_U5096, P2_U5097, P2_U5098, P2_U5099, P2_U5100, P2_U5101, P2_U5102, P2_U5103, P2_U5104, P2_U5105, P2_U5106, P2_U5107, P2_U5108, P2_U5109, P2_U5110, P2_U5111, P2_U5112, P2_U5113, P2_U5114, P2_U5115, P2_U5116, P2_U5117, P2_U5118, P2_U5119, P2_U5120, P2_U5121, P2_U5122, P2_U5123, P2_U5124, P2_U5125, P2_U5126, P2_U5127, P2_U5128, P2_U5129, P2_U5130, P2_U5131, P2_U5132, P2_U5133, P2_U5134, P2_U5135, P2_U5136, P2_U5137, P2_U5138, P2_U5139, P2_U5140, P2_U5141, P2_U5142, P2_U5143, P2_U5144, P2_U5145, P2_U5146, P2_U5147, P2_U5148, P2_U5149, P2_U5150, P2_U5151, P2_U5152, P2_U5153, P2_U5154, P2_U5155, P2_U5156, P2_U5157, P2_U5158, P2_U5159, P2_U5160, P2_U5161, P2_U5162, P2_U5163, P2_U5164, P2_U5165, P2_U5166, P2_U5167, P2_U5168, P2_U5169, P2_U5170, P2_U5171, P2_U5172, P2_U5173, P2_U5174, P2_U5175, P2_U5176, P2_U5177, P2_U5178, P2_U5179, P2_U5180, P2_U5181, P2_U5182, P2_U5183, P2_U5184, P2_U5185, P2_U5186, P2_U5187, P2_U5188, P2_U5189, P2_U5190, P2_U5191, P2_U5192, P2_U5193, P2_U5194, P2_U5195, P2_U5196, P2_U5197, P2_U5198, P2_U5199, P2_U5200, P2_U5201, P2_U5202, P2_U5203, P2_U5204, P2_U5205, P2_U5206, P2_U5207, P2_U5208, P2_U5209, P2_U5210, P2_U5211, P2_U5212, P2_U5213, P2_U5214, P2_U5215, P2_U5216, P2_U5217, P2_U5218, P2_U5219, P2_U5220, P2_U5221, P2_U5222, P2_U5223, P2_U5224, P2_U5225, P2_U5226, P2_U5227, P2_U5228, P2_U5229, P2_U5230, P2_U5231, P2_U5232, P2_U5233, P2_U5234, P2_U5235, P2_U5236, P2_U5237, P2_U5238, P2_U5239, P2_U5240, P2_U5241, P2_U5242, P2_U5243, P2_U5244, P2_U5245, P2_U5246, P2_U5247, P2_U5248, P2_U5249, P2_U5250, P2_U5251, P2_U5252, P2_U5253, P2_U5254, P2_U5255, P2_U5256, P2_U5257, P2_U5258, P2_U5259, P2_U5260, P2_U5261, P2_U5262, P2_U5263, P2_U5264, P2_U5265, P2_U5266, P2_U5267, P2_U5268, P2_U5269, P2_U5270, P2_U5271, P2_U5272, P2_U5273, P2_U5274, P2_U5275, P2_U5276, P2_U5277, P2_U5278, P2_U5279, P2_U5280, P2_U5281, P2_U5282, P2_U5283, P2_U5284, P2_U5285, P2_U5286, P2_U5287, P2_U5288, P2_U5289, P2_U5290, P2_U5291, P2_U5292, P2_U5293, P2_U5294, P2_U5295, P2_U5296, P2_U5297, P2_U5298, P2_U5299, P2_U5300, P2_U5301, P2_U5302, P2_U5303, P2_U5304, P2_U5305, P2_U5306, P2_U5307, P2_U5308, P2_U5309, P2_U5310, P2_U5311, P2_U5312, P2_U5313, P2_U5314, P2_U5315, P2_U5316, P2_U5317, P2_U5318, P2_U5319, P2_U5320, P2_U5321, P2_U5322, P2_U5323, P2_U5324, P2_U5325, P2_U5326, P2_U5327, P2_U5328, P2_U5329, P2_U5330, P2_U5331, P2_U5332, P2_U5333, P2_U5334, P2_U5335, P2_U5336, P2_U5337, P2_U5338, P2_U5339, P2_U5340, P2_U5341, P2_U5342, P2_U5343, P2_U5344, P2_U5345, P2_U5346, P2_U5347, P2_U5348, P2_U5349, P2_U5350, P2_U5351, P2_U5352, P2_U5353, P2_U5354, P2_U5355, P2_U5356, P2_U5357, P2_U5358, P2_U5359, P2_U5360, P2_U5361, P2_U5362, P2_U5363, P2_U5364, P2_U5365, P2_U5366, P2_U5367, P2_U5368, P2_U5369, P2_U5370, P2_U5371, P2_U5372, P2_U5373, P2_U5374, P2_U5375, P2_U5376, P2_U5377, P2_U5378, P2_U5379, P2_U5380, P2_U5381, P2_U5382, P2_U5383, P2_U5384, P2_U5385, P2_U5386, P2_U5387, P2_U5388, P2_U5389, P2_U5390, P2_U5391, P2_U5392, P2_U5393, P2_U5394, P2_U5395, P2_U5396, P2_U5397, P2_U5398, P2_U5399, P2_U5400, P2_U5401, P2_U5402, P2_U5403, P2_U5404, P2_U5405, P2_U5406, P2_U5407, P2_U5408, P2_U5409, P2_U5410, P2_U5411, P2_U5412, P2_U5413, P2_U5414, P2_U5415, P2_U5416, P2_U5417, P2_U5418, P2_U5419, P2_U5420, P2_U5421, P2_U5422, P2_U5423, P2_U5424, P2_U5425, P2_U5426, P2_U5427, P2_U5428, P2_U5429, P2_U5430, P2_U5431, P2_U5432, P2_U5433, P2_U5434, P2_U5435, P2_U5436, P2_U5437, P2_U5438, P2_U5439, P2_U5440, P2_U5441, P2_U5442, P2_U5443, P2_U5444, P2_U5445, P2_U5446, P2_U5447, P2_U5448, P2_U5449, P2_U5450, P2_U5451, P2_U5452, P2_U5453, P2_U5454, P2_U5455, P2_U5456, P2_U5457, P2_U5458, P2_U5459, P2_U5460, P2_U5461, P2_U5462, P2_U5463, P2_U5464, P2_U5465, P2_U5466, P2_U5467, P2_U5468, P2_U5469, P2_U5470, P2_U5471, P2_U5472, P2_U5473, P2_U5474, P2_U5475, P2_U5476, P2_U5477, P2_U5478, P2_U5479, P2_U5480, P2_U5481, P2_U5482, P2_U5483, P2_U5484, P2_U5485, P2_U5486, P2_U5487, P2_U5488, P2_U5489, P2_U5490, P2_U5491, P2_U5492, P2_U5493, P2_U5494, P2_U5495, P2_U5496, P2_U5497, P2_U5498, P2_U5499, P2_U5500, P2_U5501, P2_U5502, P2_U5503, P2_U5504, P2_U5505, P2_U5506, P2_U5507, P2_U5508, P2_U5509, P2_U5510, P2_U5511, P2_U5512, P2_U5513, P2_U5514, P2_U5515, P2_U5516, P2_U5517, P2_U5518, P2_U5519, P2_U5520, P2_U5521, P2_U5522, P2_U5523, P2_U5524, P2_U5525, P2_U5526, P2_U5527, P2_U5528, P2_U5529, P2_U5530, P2_U5531, P2_U5532, P2_U5533, P2_U5534, P2_U5535, P2_U5536, P2_U5537, P2_U5538, P2_U5539, P2_U5540, P2_U5541, P2_U5542, P2_U5543, P2_U5544, P2_U5545, P2_U5546, P2_U5547, P2_U5548, P2_U5549, P2_U5550, P2_U5551, P2_U5552, P2_U5553, P2_U5554, P2_U5555, P2_U5556, P2_U5557, P2_U5558, P2_U5559, P2_U5560, P2_U5561, P2_U5562, P2_U5563, P2_U5564, P2_U5565, P2_U5566, P2_U5567, P2_U5568, P2_U5569, P2_U5570, P2_U5571, P2_U5572, P2_U5573, P2_U5574, P2_U5575, P2_U5576, P2_U5577, P2_U5578, P2_U5579, P2_U5580, P2_U5581, P2_U5582, P2_U5583, P2_U5584, P2_U5585, P2_U5586, P2_U5587, P2_U5588, P2_U5589, P2_U5590, P2_U5591, P2_U5592, P2_U5593, P2_U5594, P2_U5595, P2_U5596, P2_U5597, P2_U5598, P2_U5599, P2_U5600, P2_U5601, P2_U5602, P2_U5603, P2_U5604, P2_U5605, P2_U5606, P2_U5607, P2_U5608, P2_U5609, P2_U5610, P2_U5611, P2_U5612, P2_U5613, P2_U5614, P2_U5615, P2_U5616, P2_U5617, P2_U5618, P2_U5619, P2_U5620, P2_U5621, P2_U5622, P2_U5623, P2_U5624, P2_U5625, P2_U5626, P2_U5627, P2_U5628, P2_U5629, P2_U5630, P2_U5631, P2_U5632, P2_U5633, P2_U5634, P2_U5635, P2_U5636, P2_U5637, P2_U5638, P2_U5639, P2_U5640, P2_U5641, P2_U5642, P2_U5643, P2_U5644, P2_U5645, P2_U5646, P2_U5647, P2_U5648, P2_U5649, P2_U5650, P2_U5651, P2_U5652, P2_U5653, P2_U5654, P2_U5655, P2_U5656, P2_U5657, P2_U5658, P2_U5659, P2_U5660, P2_U5661, P2_U5662, P2_U5663, P2_U5664, P2_U5665, P2_U5666, P2_U5667, P2_U5668, P2_U5669, P2_U5670, P2_U5671, P2_U5672, P2_U5673, P2_U5674, P2_U5675, P2_U5676, P2_U5677, P2_U5678, P2_U5679, P2_U5680, P2_U5681, P2_U5682, P2_U5683, P2_U5684, P2_U5685, P2_U5686, P2_U5687, P2_U5688, P2_U5689, P2_U5690, P2_U5691, P2_U5692, P2_U5693, P2_U5694, P2_U5695, P2_U5696, P2_U5697, P2_U5698, P2_U5699, P2_U5700, P2_U5701, P2_U5702, P2_U5703, P2_U5704, P2_U5705, P2_U5706, P2_U5707, P2_U5708, P2_U5709, P2_U5710, P2_U5711, P2_U5712, P2_U5713, P2_U5714, P2_U5715, P2_U5716, P2_U5717, P2_U5718, P2_U5719, P2_U5720, P2_U5721, P2_U5722, P2_U5723, P2_U5724, P2_U5725, P2_U5726, P2_U5727, P2_U5728, P2_U5729, P2_U5730, P2_U5731, P2_U5732, P2_U5733, P2_U5734, P2_U5735, P2_U5736, P2_U5737, P2_U5738, P2_U5739, P2_U5740, P2_U5741, P2_U5742, P2_U5743, P2_U5744, P2_U5745, P2_U5746, P2_U5747, P2_U5748, P2_U5749, P2_U5750, P2_U5751, P2_U5752, P2_U5753, P2_U5754, P2_U5755, P2_U5756, P2_U5757, P2_U5758, P2_U5759, P2_U5760, P2_U5761, P2_U5762, P2_U5763, P2_U5764, P2_U5765, P2_U5766, P2_U5767, P2_U5768, P2_U5769, P2_U5770, P2_U5771, P2_U5772, P2_U5773, P2_U5774, P2_U5775, P2_U5776, P2_U5777, P2_U5778, P2_U5779, P2_U5780, P2_U5781, P2_U5782, P2_U5783, P2_U5784, P2_U5785, P2_U5786, P2_U5787, P2_U5788, P2_U5789, P2_U5790, P2_U5791, P2_U5792, P2_U5793, P2_U5794, P2_U5795, P2_U5796, P2_U5797, P2_U5798, P2_U5799, P2_U5800, P2_U5801, P2_U5802, P2_U5803, P2_U5804, P2_U5805, P2_U5806, P2_U5807, P2_U5808, P2_U5809, P2_U5810, P2_U5811, P2_U5812, P2_U5813, P2_U5814, P2_U5815, P2_U5816, P2_U5817, P2_U5818, P2_U5819, P2_U5820, P2_U5821, P2_U5822, P2_U5823, P2_U5824, P2_U5825, P2_U5826, P2_U5827, P2_U5828, P2_U5829, P2_U5830, P2_U5831, P2_U5832, P2_U5833, P2_U5834, P2_U5835, P2_U5836, P2_U5837, P2_U5838, P2_U5839, P2_U5840, P2_U5841, P2_U5842, P2_U5843, P2_U5844, P2_U5845, P2_U5846, P2_U5847, P2_U5848, P2_U5849, P2_U5850, P2_U5851, P2_U5852, P2_U5853, P2_U5854, P2_U5855, P2_U5856, P2_U5857, P2_U5858, P2_U5859, P2_U5860, P2_U5861, P2_U5862, P2_U5863, P2_U5864, P2_U5865, P2_U5866, P2_U5867, P2_U5868, P2_U5869, P2_U5870, P2_U5871, P2_U5872, P2_U5873, P2_U5874, P2_U5875, P2_U5876, P2_U5877, P2_U5878, P2_U5879, P2_U5880, P2_U5881, P2_U5882, P2_U5883, P2_U5884, P2_U5885, P2_U5886, P2_U5887, P2_U5888, P2_U5889, P2_U5890, P2_U5891, P2_U5892, P2_U5893, P2_U5894, P2_U5895, P2_U5896, P2_U5897, P2_U5898, P2_U5899, P2_U5900, P2_U5901, P2_U5902, P2_U5903, P2_U5904, P2_U5905, P2_U5906, P2_U5907, P2_U5908, P2_U5909, P2_U5910, P2_U5911, P2_U5912, P2_U5913, P2_U5914, P2_U5915, P2_U5916, P2_U5917, P2_U5918, P2_U5919, P2_U5920, P2_U5921, P2_U5922, P2_U5923, P2_U5924, P2_U5925, P2_U5926, P2_U5927, P2_U5928, P2_U5929, P2_U5930, P2_U5931, P2_U5932, P2_U5933, P2_U5934, P2_U5935, P2_U5936, P2_U5937, P2_U5938, P2_U5939, P2_U5940, P2_U5941, P2_U5942, P2_U5943, P2_U5944, P2_U5945, P2_U5946, P2_U5947, P2_U5948, P2_U5949, P2_U5950, P2_U5951, P2_U5952, P2_U5953, P2_U5954, P2_U5955, P2_U5956, P2_U5957, P2_U5958, P2_U5959, P2_U5960, P2_U5961, P2_U5962, P2_U5963, P2_U5964, P2_U5965, P2_U5966, P2_U5967, P2_U5968, P2_U5969, P2_U5970, P2_U5971, P2_U5972, P2_U5973, P2_U5974, P2_U5975, P2_U5976, P2_U5977, P2_U5978, P2_U5979, P2_U5980, P2_U5981, P2_U5982, P2_U5983, P2_U5984, P2_U5985, P2_U5986, P2_U5987, P2_U5988, P2_U5989, P2_U5990, P2_U5991, P2_U5992, P2_U5993, P2_U5994, P2_U5995, P2_U5996, P2_U5997, P2_U5998, P2_U5999, P2_U6000, P2_U6001, P2_U6002, P2_U6003, P2_U6004, P2_U6005, P2_U6006, P2_U6007, P2_U6008, P2_U6009, P2_U6010, P2_U6011, P2_U6012, P2_U6013, P2_U6014, P2_U6015, P2_U6016, P2_U6017, P2_U6018, P2_U6019, P2_U6020, P2_U6021, P2_U6022, P2_U6023, P2_U6024, P2_U6025, P2_U6026, P2_U6027, P2_U6028, P2_U6029, P2_U6030, P2_U6031, P2_U6032, P2_U6033, P2_U6034, P2_U6035, P2_U6036, P2_U6037, P2_U6038, P2_U6039, P2_U6040, P2_U6041, P2_U6042, P2_U6043, P2_U6044, R140_U10, R140_U100, R140_U101, R140_U102, R140_U103, R140_U104, R140_U105, R140_U106, R140_U107, R140_U108, R140_U109, R140_U11, R140_U110, R140_U111, R140_U112, R140_U113, R140_U114, R140_U115, R140_U116, R140_U117, R140_U118, R140_U119, R140_U12, R140_U120, R140_U121, R140_U122, R140_U123, R140_U124, R140_U125, R140_U126, R140_U127, R140_U128, R140_U129, R140_U13, R140_U130, R140_U131, R140_U132, R140_U133, R140_U134, R140_U135, R140_U136, R140_U137, R140_U138, R140_U139, R140_U14, R140_U140, R140_U141, R140_U142, R140_U143, R140_U144, R140_U145, R140_U146, R140_U147, R140_U148, R140_U149, R140_U15, R140_U150, R140_U151, R140_U152, R140_U153, R140_U154, R140_U155, R140_U156, R140_U157, R140_U158, R140_U159, R140_U16, R140_U160, R140_U161, R140_U162, R140_U163, R140_U164, R140_U165, R140_U166, R140_U167, R140_U168, R140_U169, R140_U17, R140_U170, R140_U171, R140_U172, R140_U173, R140_U174, R140_U175, R140_U176, R140_U177, R140_U178, R140_U179, R140_U18, R140_U180, R140_U181, R140_U182, R140_U183, R140_U184, R140_U185, R140_U186, R140_U187, R140_U188, R140_U189, R140_U19, R140_U190, R140_U191, R140_U192, R140_U193, R140_U194, R140_U195, R140_U196, R140_U197, R140_U198, R140_U199, R140_U20, R140_U200, R140_U201, R140_U202, R140_U203, R140_U204, R140_U205, R140_U206, R140_U207, R140_U208, R140_U209, R140_U21, R140_U210, R140_U211, R140_U212, R140_U213, R140_U214, R140_U215, R140_U216, R140_U217, R140_U218, R140_U219, R140_U22, R140_U220, R140_U221, R140_U222, R140_U223, R140_U224, R140_U225, R140_U226, R140_U227, R140_U228, R140_U229, R140_U23, R140_U230, R140_U231, R140_U232, R140_U233, R140_U234, R140_U235, R140_U236, R140_U237, R140_U238, R140_U239, R140_U24, R140_U240, R140_U241, R140_U242, R140_U243, R140_U244, R140_U245, R140_U246, R140_U247, R140_U248, R140_U249, R140_U25, R140_U250, R140_U251, R140_U252, R140_U253, R140_U254, R140_U255, R140_U256, R140_U257, R140_U258, R140_U259, R140_U26, R140_U260, R140_U261, R140_U262, R140_U263, R140_U264, R140_U265, R140_U266, R140_U267, R140_U268, R140_U269, R140_U27, R140_U270, R140_U271, R140_U272, R140_U273, R140_U274, R140_U275, R140_U276, R140_U277, R140_U278, R140_U279, R140_U28, R140_U280, R140_U281, R140_U282, R140_U283, R140_U284, R140_U285, R140_U286, R140_U287, R140_U288, R140_U289, R140_U29, R140_U290, R140_U291, R140_U292, R140_U293, R140_U294, R140_U295, R140_U296, R140_U297, R140_U298, R140_U299, R140_U30, R140_U300, R140_U301, R140_U302, R140_U303, R140_U304, R140_U305, R140_U306, R140_U307, R140_U308, R140_U309, R140_U31, R140_U310, R140_U311, R140_U312, R140_U313, R140_U314, R140_U315, R140_U316, R140_U317, R140_U318, R140_U319, R140_U32, R140_U320, R140_U321, R140_U322, R140_U323, R140_U324, R140_U325, R140_U326, R140_U327, R140_U328, R140_U329, R140_U33, R140_U330, R140_U331, R140_U332, R140_U333, R140_U334, R140_U335, R140_U336, R140_U337, R140_U338, R140_U339, R140_U34, R140_U340, R140_U341, R140_U342, R140_U343, R140_U344, R140_U345, R140_U346, R140_U347, R140_U348, R140_U349, R140_U35, R140_U350, R140_U351, R140_U352, R140_U353, R140_U354, R140_U355, R140_U356, R140_U357, R140_U358, R140_U359, R140_U36, R140_U360, R140_U361, R140_U362, R140_U363, R140_U364, R140_U365, R140_U366, R140_U367, R140_U368, R140_U369, R140_U37, R140_U370, R140_U371, R140_U372, R140_U373, R140_U374, R140_U375, R140_U376, R140_U377, R140_U378, R140_U379, R140_U38, R140_U380, R140_U381, R140_U382, R140_U383, R140_U384, R140_U385, R140_U386, R140_U387, R140_U388, R140_U389, R140_U39, R140_U390, R140_U391, R140_U392, R140_U393, R140_U394, R140_U395, R140_U396, R140_U397, R140_U398, R140_U399, R140_U4, R140_U40, R140_U400, R140_U401, R140_U402, R140_U403, R140_U404, R140_U405, R140_U406, R140_U407, R140_U408, R140_U409, R140_U41, R140_U410, R140_U411, R140_U412, R140_U413, R140_U414, R140_U415, R140_U416, R140_U417, R140_U418, R140_U419, R140_U42, R140_U420, R140_U421, R140_U422, R140_U423, R140_U424, R140_U425, R140_U426, R140_U427, R140_U428, R140_U429, R140_U43, R140_U430, R140_U431, R140_U432, R140_U433, R140_U434, R140_U435, R140_U436, R140_U437, R140_U438, R140_U439, R140_U44, R140_U440, R140_U441, R140_U442, R140_U443, R140_U444, R140_U445, R140_U446, R140_U447, R140_U448, R140_U449, R140_U45, R140_U450, R140_U451, R140_U452, R140_U453, R140_U454, R140_U455, R140_U456, R140_U457, R140_U458, R140_U459, R140_U46, R140_U460, R140_U461, R140_U462, R140_U463, R140_U464, R140_U465, R140_U466, R140_U467, R140_U468, R140_U469, R140_U47, R140_U470, R140_U471, R140_U472, R140_U473, R140_U474, R140_U475, R140_U476, R140_U477, R140_U478, R140_U479, R140_U48, R140_U480, R140_U481, R140_U482, R140_U483, R140_U484, R140_U485, R140_U486, R140_U487, R140_U488, R140_U489, R140_U49, R140_U490, R140_U491, R140_U492, R140_U493, R140_U494, R140_U495, R140_U496, R140_U497, R140_U498, R140_U499, R140_U5, R140_U50, R140_U500, R140_U501, R140_U502, R140_U503, R140_U504, R140_U505, R140_U506, R140_U507, R140_U508, R140_U509, R140_U51, R140_U510, R140_U511, R140_U512, R140_U513, R140_U514, R140_U515, R140_U516, R140_U517, R140_U518, R140_U519, R140_U52, R140_U520, R140_U521, R140_U522, R140_U523, R140_U524, R140_U525, R140_U526, R140_U527, R140_U528, R140_U529, R140_U53, R140_U530, R140_U531, R140_U532, R140_U533, R140_U534, R140_U535, R140_U536, R140_U537, R140_U538, R140_U539, R140_U54, R140_U540, R140_U541, R140_U55, R140_U56, R140_U57, R140_U58, R140_U59, R140_U6, R140_U60, R140_U61, R140_U62, R140_U63, R140_U64, R140_U65, R140_U66, R140_U67, R140_U68, R140_U69, R140_U7, R140_U70, R140_U71, R140_U72, R140_U73, R140_U74, R140_U75, R140_U76, R140_U77, R140_U78, R140_U79, R140_U8, R140_U80, R140_U81, R140_U82, R140_U83, R140_U84, R140_U85, R140_U86, R140_U87, R140_U88, R140_U89, R140_U9, R140_U90, R140_U91, R140_U92, R140_U93, R140_U94, R140_U95, R140_U96, R140_U97, R140_U98, R140_U99, U100, U101, U102, U103, U104, U105, U106, U107, U108, U109, U110, U111, U112, U113, U114, U115, U116, U117, U118, U119, U120, U121, U122, U124, U125, U127, U128, U129, U130, U131, U132, U133, U134, U135, U136, U137, U138, U139, U140, U141, U142, U143, U144, U145, U146, U147, U148, U149, U150, U151, U152, U153, U154, U155, U156, U157, U158, U159, U160, U161, U162, U163, U164, U165, U166, U167, U168, U169, U170, U171, U172, U173, U174, U175, U176, U177, U178, U179, U180, U181, U182, U183, U184, U185, U186, U187, U188, U189, U190, U191, U192, U193, U194, U195, U196, U197, U198, U199, U200, U201, U202, U203, U204, U205, U206, U207, U208, U209, U210, U211, U212, U213, U214, U215, U216, U217, U218, U219, U220, U221, U222, U223, U224, U225, U226, U227, U228, U229, U230, U231, U232, U233, U234, U235, U236, U237, U238, U239, U240, U241, U242, U243, U244, U245, U246, U247, U248, U249, U25, U250, U251, U252, U253, U254, U255, U256, U257, U258, U259, U26, U260, U261, U262, U263, U264, U265, U266, U267, U268, U269, U27, U270, U271, U272, U273, U274, U275, U276, U277, U278, U279, U28, U280, U281, U282, U283, U284, U285, U286, U287, U288, U289, U29, U290, U291, U292, U293, U294, U295, U296, U297, U298, U299, U30, U300, U301, U302, U303, U304, U305, U306, U307, U308, U309, U31, U310, U311, U312, U313, U314, U315, U316, U317, U318, U319, U32, U320, U321, U322, U323, U324, U325, U326, U33, U34, U35, U36, U37, U38, U39, U40, U41, U42, U43, U44, U45, U46, U47, U48, U49, U50, U51, U52, U53, U54, U55, U56, U57, U58, U59, U60, U61, U62, U63, U64, U65, U66, U67, U68, U69, U70, U71, U72, U73, U74, U75, U76, U77, U78, U79, U80, U81, U82, U83, U84, U85, U86, U87, U88, U89, U90, U91, U92, U93, U94, U95, U96, U97, U98, U99, P1_U3279_in, flip_signal;

  not ginst1 (ADD_1068_U10, P1_ADDR_REG_1__SCAN_IN);
  or ginst2 (ADD_1068_U100, P1_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_5__SCAN_IN);
  nand ginst3 (ADD_1068_U101, ADD_1068_U100, ADD_1068_U68);
  nand ginst4 (ADD_1068_U102, P1_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_5__SCAN_IN);
  not ginst5 (ADD_1068_U103, ADD_1068_U67);
  or ginst6 (ADD_1068_U104, P1_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_6__SCAN_IN);
  nand ginst7 (ADD_1068_U105, ADD_1068_U104, ADD_1068_U67);
  nand ginst8 (ADD_1068_U106, P1_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_6__SCAN_IN);
  not ginst9 (ADD_1068_U107, ADD_1068_U66);
  or ginst10 (ADD_1068_U108, P1_ADDR_REG_7__SCAN_IN, P2_ADDR_REG_7__SCAN_IN);
  nand ginst11 (ADD_1068_U109, ADD_1068_U108, ADD_1068_U66);
  not ginst12 (ADD_1068_U11, P1_ADDR_REG_2__SCAN_IN);
  nand ginst13 (ADD_1068_U110, P1_ADDR_REG_7__SCAN_IN, P2_ADDR_REG_7__SCAN_IN);
  not ginst14 (ADD_1068_U111, ADD_1068_U65);
  or ginst15 (ADD_1068_U112, P1_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_8__SCAN_IN);
  nand ginst16 (ADD_1068_U113, ADD_1068_U112, ADD_1068_U65);
  nand ginst17 (ADD_1068_U114, P1_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_8__SCAN_IN);
  not ginst18 (ADD_1068_U115, ADD_1068_U64);
  or ginst19 (ADD_1068_U116, P1_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_9__SCAN_IN);
  nand ginst20 (ADD_1068_U117, ADD_1068_U116, ADD_1068_U64);
  nand ginst21 (ADD_1068_U118, P1_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_9__SCAN_IN);
  not ginst22 (ADD_1068_U119, ADD_1068_U82);
  not ginst23 (ADD_1068_U12, P2_ADDR_REG_2__SCAN_IN);
  or ginst24 (ADD_1068_U120, P1_ADDR_REG_10__SCAN_IN, P2_ADDR_REG_10__SCAN_IN);
  nand ginst25 (ADD_1068_U121, ADD_1068_U120, ADD_1068_U82);
  nand ginst26 (ADD_1068_U122, P1_ADDR_REG_10__SCAN_IN, P2_ADDR_REG_10__SCAN_IN);
  not ginst27 (ADD_1068_U123, ADD_1068_U81);
  or ginst28 (ADD_1068_U124, P1_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_11__SCAN_IN);
  nand ginst29 (ADD_1068_U125, ADD_1068_U124, ADD_1068_U81);
  nand ginst30 (ADD_1068_U126, P1_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_11__SCAN_IN);
  not ginst31 (ADD_1068_U127, ADD_1068_U80);
  or ginst32 (ADD_1068_U128, P1_ADDR_REG_12__SCAN_IN, P2_ADDR_REG_12__SCAN_IN);
  nand ginst33 (ADD_1068_U129, ADD_1068_U128, ADD_1068_U80);
  not ginst34 (ADD_1068_U13, P1_ADDR_REG_3__SCAN_IN);
  nand ginst35 (ADD_1068_U130, P1_ADDR_REG_12__SCAN_IN, P2_ADDR_REG_12__SCAN_IN);
  not ginst36 (ADD_1068_U131, ADD_1068_U79);
  or ginst37 (ADD_1068_U132, P1_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_13__SCAN_IN);
  nand ginst38 (ADD_1068_U133, ADD_1068_U132, ADD_1068_U79);
  nand ginst39 (ADD_1068_U134, P1_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_13__SCAN_IN);
  not ginst40 (ADD_1068_U135, ADD_1068_U78);
  or ginst41 (ADD_1068_U136, P1_ADDR_REG_14__SCAN_IN, P2_ADDR_REG_14__SCAN_IN);
  nand ginst42 (ADD_1068_U137, ADD_1068_U136, ADD_1068_U78);
  nand ginst43 (ADD_1068_U138, P1_ADDR_REG_14__SCAN_IN, P2_ADDR_REG_14__SCAN_IN);
  not ginst44 (ADD_1068_U139, ADD_1068_U77);
  not ginst45 (ADD_1068_U14, P2_ADDR_REG_3__SCAN_IN);
  or ginst46 (ADD_1068_U140, P1_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_15__SCAN_IN);
  nand ginst47 (ADD_1068_U141, ADD_1068_U140, ADD_1068_U77);
  nand ginst48 (ADD_1068_U142, P1_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_15__SCAN_IN);
  not ginst49 (ADD_1068_U143, ADD_1068_U76);
  or ginst50 (ADD_1068_U144, P1_ADDR_REG_16__SCAN_IN, P2_ADDR_REG_16__SCAN_IN);
  nand ginst51 (ADD_1068_U145, ADD_1068_U144, ADD_1068_U76);
  nand ginst52 (ADD_1068_U146, P1_ADDR_REG_16__SCAN_IN, P2_ADDR_REG_16__SCAN_IN);
  not ginst53 (ADD_1068_U147, ADD_1068_U75);
  or ginst54 (ADD_1068_U148, P1_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_17__SCAN_IN);
  nand ginst55 (ADD_1068_U149, ADD_1068_U148, ADD_1068_U75);
  not ginst56 (ADD_1068_U15, P1_ADDR_REG_4__SCAN_IN);
  nand ginst57 (ADD_1068_U150, P1_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_17__SCAN_IN);
  not ginst58 (ADD_1068_U151, ADD_1068_U45);
  or ginst59 (ADD_1068_U152, P1_ADDR_REG_18__SCAN_IN, P2_ADDR_REG_18__SCAN_IN);
  nand ginst60 (ADD_1068_U153, ADD_1068_U152, ADD_1068_U45);
  nand ginst61 (ADD_1068_U154, P1_ADDR_REG_18__SCAN_IN, P2_ADDR_REG_18__SCAN_IN);
  nand ginst62 (ADD_1068_U155, ADD_1068_U153, ADD_1068_U154, ADD_1068_U222, ADD_1068_U223);
  nand ginst63 (ADD_1068_U156, P1_ADDR_REG_18__SCAN_IN, P2_ADDR_REG_18__SCAN_IN);
  nand ginst64 (ADD_1068_U157, ADD_1068_U151, ADD_1068_U156);
  or ginst65 (ADD_1068_U158, P1_ADDR_REG_18__SCAN_IN, P2_ADDR_REG_18__SCAN_IN);
  nand ginst66 (ADD_1068_U159, ADD_1068_U157, ADD_1068_U158, ADD_1068_U226);
  not ginst67 (ADD_1068_U16, P2_ADDR_REG_4__SCAN_IN);
  nand ginst68 (ADD_1068_U160, ADD_1068_U10, ADD_1068_U219);
  nand ginst69 (ADD_1068_U161, P2_ADDR_REG_9__SCAN_IN, ADD_1068_U26);
  nand ginst70 (ADD_1068_U162, P1_ADDR_REG_9__SCAN_IN, ADD_1068_U25);
  nand ginst71 (ADD_1068_U163, P2_ADDR_REG_9__SCAN_IN, ADD_1068_U26);
  nand ginst72 (ADD_1068_U164, P1_ADDR_REG_9__SCAN_IN, ADD_1068_U25);
  nand ginst73 (ADD_1068_U165, ADD_1068_U163, ADD_1068_U164);
  nand ginst74 (ADD_1068_U166, ADD_1068_U161, ADD_1068_U162, ADD_1068_U64);
  nand ginst75 (ADD_1068_U167, ADD_1068_U115, ADD_1068_U165);
  nand ginst76 (ADD_1068_U168, P2_ADDR_REG_8__SCAN_IN, ADD_1068_U23);
  nand ginst77 (ADD_1068_U169, P1_ADDR_REG_8__SCAN_IN, ADD_1068_U24);
  not ginst78 (ADD_1068_U17, P1_ADDR_REG_5__SCAN_IN);
  nand ginst79 (ADD_1068_U170, P2_ADDR_REG_8__SCAN_IN, ADD_1068_U23);
  nand ginst80 (ADD_1068_U171, P1_ADDR_REG_8__SCAN_IN, ADD_1068_U24);
  nand ginst81 (ADD_1068_U172, ADD_1068_U170, ADD_1068_U171);
  nand ginst82 (ADD_1068_U173, ADD_1068_U168, ADD_1068_U169, ADD_1068_U65);
  nand ginst83 (ADD_1068_U174, ADD_1068_U111, ADD_1068_U172);
  nand ginst84 (ADD_1068_U175, P2_ADDR_REG_7__SCAN_IN, ADD_1068_U21);
  nand ginst85 (ADD_1068_U176, P1_ADDR_REG_7__SCAN_IN, ADD_1068_U22);
  nand ginst86 (ADD_1068_U177, P2_ADDR_REG_7__SCAN_IN, ADD_1068_U21);
  nand ginst87 (ADD_1068_U178, P1_ADDR_REG_7__SCAN_IN, ADD_1068_U22);
  nand ginst88 (ADD_1068_U179, ADD_1068_U177, ADD_1068_U178);
  not ginst89 (ADD_1068_U18, P2_ADDR_REG_5__SCAN_IN);
  nand ginst90 (ADD_1068_U180, ADD_1068_U175, ADD_1068_U176, ADD_1068_U66);
  nand ginst91 (ADD_1068_U181, ADD_1068_U107, ADD_1068_U179);
  nand ginst92 (ADD_1068_U182, P2_ADDR_REG_6__SCAN_IN, ADD_1068_U19);
  nand ginst93 (ADD_1068_U183, P1_ADDR_REG_6__SCAN_IN, ADD_1068_U20);
  nand ginst94 (ADD_1068_U184, P2_ADDR_REG_6__SCAN_IN, ADD_1068_U19);
  nand ginst95 (ADD_1068_U185, P1_ADDR_REG_6__SCAN_IN, ADD_1068_U20);
  nand ginst96 (ADD_1068_U186, ADD_1068_U184, ADD_1068_U185);
  nand ginst97 (ADD_1068_U187, ADD_1068_U182, ADD_1068_U183, ADD_1068_U67);
  nand ginst98 (ADD_1068_U188, ADD_1068_U103, ADD_1068_U186);
  nand ginst99 (ADD_1068_U189, P2_ADDR_REG_5__SCAN_IN, ADD_1068_U17);
  not ginst100 (ADD_1068_U19, P1_ADDR_REG_6__SCAN_IN);
  nand ginst101 (ADD_1068_U190, P1_ADDR_REG_5__SCAN_IN, ADD_1068_U18);
  nand ginst102 (ADD_1068_U191, P2_ADDR_REG_5__SCAN_IN, ADD_1068_U17);
  nand ginst103 (ADD_1068_U192, P1_ADDR_REG_5__SCAN_IN, ADD_1068_U18);
  nand ginst104 (ADD_1068_U193, ADD_1068_U191, ADD_1068_U192);
  nand ginst105 (ADD_1068_U194, ADD_1068_U189, ADD_1068_U190, ADD_1068_U68);
  nand ginst106 (ADD_1068_U195, ADD_1068_U193, ADD_1068_U99);
  nand ginst107 (ADD_1068_U196, P2_ADDR_REG_4__SCAN_IN, ADD_1068_U15);
  nand ginst108 (ADD_1068_U197, P1_ADDR_REG_4__SCAN_IN, ADD_1068_U16);
  nand ginst109 (ADD_1068_U198, P2_ADDR_REG_4__SCAN_IN, ADD_1068_U15);
  nand ginst110 (ADD_1068_U199, P1_ADDR_REG_4__SCAN_IN, ADD_1068_U16);
  not ginst111 (ADD_1068_U20, P2_ADDR_REG_6__SCAN_IN);
  nand ginst112 (ADD_1068_U200, ADD_1068_U198, ADD_1068_U199);
  nand ginst113 (ADD_1068_U201, ADD_1068_U196, ADD_1068_U197, ADD_1068_U69);
  nand ginst114 (ADD_1068_U202, ADD_1068_U200, ADD_1068_U95);
  nand ginst115 (ADD_1068_U203, P2_ADDR_REG_3__SCAN_IN, ADD_1068_U13);
  nand ginst116 (ADD_1068_U204, P1_ADDR_REG_3__SCAN_IN, ADD_1068_U14);
  nand ginst117 (ADD_1068_U205, P2_ADDR_REG_3__SCAN_IN, ADD_1068_U13);
  nand ginst118 (ADD_1068_U206, P1_ADDR_REG_3__SCAN_IN, ADD_1068_U14);
  nand ginst119 (ADD_1068_U207, ADD_1068_U205, ADD_1068_U206);
  nand ginst120 (ADD_1068_U208, ADD_1068_U203, ADD_1068_U204, ADD_1068_U70);
  nand ginst121 (ADD_1068_U209, ADD_1068_U207, ADD_1068_U91);
  not ginst122 (ADD_1068_U21, P1_ADDR_REG_7__SCAN_IN);
  nand ginst123 (ADD_1068_U210, P2_ADDR_REG_2__SCAN_IN, ADD_1068_U11);
  nand ginst124 (ADD_1068_U211, P1_ADDR_REG_2__SCAN_IN, ADD_1068_U12);
  nand ginst125 (ADD_1068_U212, P2_ADDR_REG_2__SCAN_IN, ADD_1068_U11);
  nand ginst126 (ADD_1068_U213, P1_ADDR_REG_2__SCAN_IN, ADD_1068_U12);
  nand ginst127 (ADD_1068_U214, ADD_1068_U212, ADD_1068_U213);
  nand ginst128 (ADD_1068_U215, ADD_1068_U210, ADD_1068_U211, ADD_1068_U71);
  nand ginst129 (ADD_1068_U216, ADD_1068_U214, ADD_1068_U87);
  nand ginst130 (ADD_1068_U217, P2_ADDR_REG_1__SCAN_IN, ADD_1068_U9);
  nand ginst131 (ADD_1068_U218, ADD_1068_U8, ADD_1068_U84);
  nand ginst132 (ADD_1068_U219, ADD_1068_U217, ADD_1068_U218);
  not ginst133 (ADD_1068_U22, P2_ADDR_REG_7__SCAN_IN);
  nand ginst134 (ADD_1068_U220, P1_ADDR_REG_1__SCAN_IN, ADD_1068_U8, ADD_1068_U9);
  nand ginst135 (ADD_1068_U221, P2_ADDR_REG_1__SCAN_IN, ADD_1068_U83);
  nand ginst136 (ADD_1068_U222, P2_ADDR_REG_19__SCAN_IN, ADD_1068_U74);
  nand ginst137 (ADD_1068_U223, P1_ADDR_REG_19__SCAN_IN, ADD_1068_U73);
  nand ginst138 (ADD_1068_U224, P2_ADDR_REG_19__SCAN_IN, ADD_1068_U74);
  nand ginst139 (ADD_1068_U225, P1_ADDR_REG_19__SCAN_IN, ADD_1068_U73);
  nand ginst140 (ADD_1068_U226, ADD_1068_U224, ADD_1068_U225);
  nand ginst141 (ADD_1068_U227, P2_ADDR_REG_18__SCAN_IN, ADD_1068_U43);
  nand ginst142 (ADD_1068_U228, P1_ADDR_REG_18__SCAN_IN, ADD_1068_U44);
  nand ginst143 (ADD_1068_U229, P2_ADDR_REG_18__SCAN_IN, ADD_1068_U43);
  not ginst144 (ADD_1068_U23, P1_ADDR_REG_8__SCAN_IN);
  nand ginst145 (ADD_1068_U230, P1_ADDR_REG_18__SCAN_IN, ADD_1068_U44);
  nand ginst146 (ADD_1068_U231, ADD_1068_U229, ADD_1068_U230);
  nand ginst147 (ADD_1068_U232, ADD_1068_U227, ADD_1068_U228, ADD_1068_U45);
  nand ginst148 (ADD_1068_U233, ADD_1068_U151, ADD_1068_U231);
  nand ginst149 (ADD_1068_U234, P2_ADDR_REG_17__SCAN_IN, ADD_1068_U41);
  nand ginst150 (ADD_1068_U235, P1_ADDR_REG_17__SCAN_IN, ADD_1068_U42);
  nand ginst151 (ADD_1068_U236, P2_ADDR_REG_17__SCAN_IN, ADD_1068_U41);
  nand ginst152 (ADD_1068_U237, P1_ADDR_REG_17__SCAN_IN, ADD_1068_U42);
  nand ginst153 (ADD_1068_U238, ADD_1068_U236, ADD_1068_U237);
  nand ginst154 (ADD_1068_U239, ADD_1068_U234, ADD_1068_U235, ADD_1068_U75);
  not ginst155 (ADD_1068_U24, P2_ADDR_REG_8__SCAN_IN);
  nand ginst156 (ADD_1068_U240, ADD_1068_U147, ADD_1068_U238);
  nand ginst157 (ADD_1068_U241, P2_ADDR_REG_16__SCAN_IN, ADD_1068_U39);
  nand ginst158 (ADD_1068_U242, P1_ADDR_REG_16__SCAN_IN, ADD_1068_U40);
  nand ginst159 (ADD_1068_U243, P2_ADDR_REG_16__SCAN_IN, ADD_1068_U39);
  nand ginst160 (ADD_1068_U244, P1_ADDR_REG_16__SCAN_IN, ADD_1068_U40);
  nand ginst161 (ADD_1068_U245, ADD_1068_U243, ADD_1068_U244);
  nand ginst162 (ADD_1068_U246, ADD_1068_U241, ADD_1068_U242, ADD_1068_U76);
  nand ginst163 (ADD_1068_U247, ADD_1068_U143, ADD_1068_U245);
  nand ginst164 (ADD_1068_U248, P2_ADDR_REG_15__SCAN_IN, ADD_1068_U37);
  nand ginst165 (ADD_1068_U249, P1_ADDR_REG_15__SCAN_IN, ADD_1068_U38);
  not ginst166 (ADD_1068_U25, P2_ADDR_REG_9__SCAN_IN);
  nand ginst167 (ADD_1068_U250, P2_ADDR_REG_15__SCAN_IN, ADD_1068_U37);
  nand ginst168 (ADD_1068_U251, P1_ADDR_REG_15__SCAN_IN, ADD_1068_U38);
  nand ginst169 (ADD_1068_U252, ADD_1068_U250, ADD_1068_U251);
  nand ginst170 (ADD_1068_U253, ADD_1068_U248, ADD_1068_U249, ADD_1068_U77);
  nand ginst171 (ADD_1068_U254, ADD_1068_U139, ADD_1068_U252);
  nand ginst172 (ADD_1068_U255, P2_ADDR_REG_14__SCAN_IN, ADD_1068_U35);
  nand ginst173 (ADD_1068_U256, P1_ADDR_REG_14__SCAN_IN, ADD_1068_U36);
  nand ginst174 (ADD_1068_U257, P2_ADDR_REG_14__SCAN_IN, ADD_1068_U35);
  nand ginst175 (ADD_1068_U258, P1_ADDR_REG_14__SCAN_IN, ADD_1068_U36);
  nand ginst176 (ADD_1068_U259, ADD_1068_U257, ADD_1068_U258);
  not ginst177 (ADD_1068_U26, P1_ADDR_REG_9__SCAN_IN);
  nand ginst178 (ADD_1068_U260, ADD_1068_U255, ADD_1068_U256, ADD_1068_U78);
  nand ginst179 (ADD_1068_U261, ADD_1068_U135, ADD_1068_U259);
  nand ginst180 (ADD_1068_U262, P2_ADDR_REG_13__SCAN_IN, ADD_1068_U33);
  nand ginst181 (ADD_1068_U263, P1_ADDR_REG_13__SCAN_IN, ADD_1068_U34);
  nand ginst182 (ADD_1068_U264, P2_ADDR_REG_13__SCAN_IN, ADD_1068_U33);
  nand ginst183 (ADD_1068_U265, P1_ADDR_REG_13__SCAN_IN, ADD_1068_U34);
  nand ginst184 (ADD_1068_U266, ADD_1068_U264, ADD_1068_U265);
  nand ginst185 (ADD_1068_U267, ADD_1068_U262, ADD_1068_U263, ADD_1068_U79);
  nand ginst186 (ADD_1068_U268, ADD_1068_U131, ADD_1068_U266);
  nand ginst187 (ADD_1068_U269, P2_ADDR_REG_12__SCAN_IN, ADD_1068_U31);
  not ginst188 (ADD_1068_U27, P1_ADDR_REG_10__SCAN_IN);
  nand ginst189 (ADD_1068_U270, P1_ADDR_REG_12__SCAN_IN, ADD_1068_U32);
  nand ginst190 (ADD_1068_U271, P2_ADDR_REG_12__SCAN_IN, ADD_1068_U31);
  nand ginst191 (ADD_1068_U272, P1_ADDR_REG_12__SCAN_IN, ADD_1068_U32);
  nand ginst192 (ADD_1068_U273, ADD_1068_U271, ADD_1068_U272);
  nand ginst193 (ADD_1068_U274, ADD_1068_U269, ADD_1068_U270, ADD_1068_U80);
  nand ginst194 (ADD_1068_U275, ADD_1068_U127, ADD_1068_U273);
  nand ginst195 (ADD_1068_U276, P2_ADDR_REG_11__SCAN_IN, ADD_1068_U29);
  nand ginst196 (ADD_1068_U277, P1_ADDR_REG_11__SCAN_IN, ADD_1068_U30);
  nand ginst197 (ADD_1068_U278, P2_ADDR_REG_11__SCAN_IN, ADD_1068_U29);
  nand ginst198 (ADD_1068_U279, P1_ADDR_REG_11__SCAN_IN, ADD_1068_U30);
  not ginst199 (ADD_1068_U28, P2_ADDR_REG_10__SCAN_IN);
  nand ginst200 (ADD_1068_U280, ADD_1068_U278, ADD_1068_U279);
  nand ginst201 (ADD_1068_U281, ADD_1068_U276, ADD_1068_U277, ADD_1068_U81);
  nand ginst202 (ADD_1068_U282, ADD_1068_U123, ADD_1068_U280);
  nand ginst203 (ADD_1068_U283, P2_ADDR_REG_10__SCAN_IN, ADD_1068_U27);
  nand ginst204 (ADD_1068_U284, P1_ADDR_REG_10__SCAN_IN, ADD_1068_U28);
  nand ginst205 (ADD_1068_U285, P2_ADDR_REG_10__SCAN_IN, ADD_1068_U27);
  nand ginst206 (ADD_1068_U286, P1_ADDR_REG_10__SCAN_IN, ADD_1068_U28);
  nand ginst207 (ADD_1068_U287, ADD_1068_U285, ADD_1068_U286);
  nand ginst208 (ADD_1068_U288, ADD_1068_U283, ADD_1068_U284, ADD_1068_U82);
  nand ginst209 (ADD_1068_U289, ADD_1068_U119, ADD_1068_U287);
  not ginst210 (ADD_1068_U29, P1_ADDR_REG_11__SCAN_IN);
  nand ginst211 (ADD_1068_U290, P2_ADDR_REG_0__SCAN_IN, ADD_1068_U6);
  nand ginst212 (ADD_1068_U291, P1_ADDR_REG_0__SCAN_IN, ADD_1068_U7);
  not ginst213 (ADD_1068_U30, P2_ADDR_REG_11__SCAN_IN);
  not ginst214 (ADD_1068_U31, P1_ADDR_REG_12__SCAN_IN);
  not ginst215 (ADD_1068_U32, P2_ADDR_REG_12__SCAN_IN);
  not ginst216 (ADD_1068_U33, P1_ADDR_REG_13__SCAN_IN);
  not ginst217 (ADD_1068_U34, P2_ADDR_REG_13__SCAN_IN);
  not ginst218 (ADD_1068_U35, P1_ADDR_REG_14__SCAN_IN);
  not ginst219 (ADD_1068_U36, P2_ADDR_REG_14__SCAN_IN);
  not ginst220 (ADD_1068_U37, P1_ADDR_REG_15__SCAN_IN);
  not ginst221 (ADD_1068_U38, P2_ADDR_REG_15__SCAN_IN);
  not ginst222 (ADD_1068_U39, P1_ADDR_REG_16__SCAN_IN);
  and ginst223 (ADD_1068_U4, ADD_1068_U155, ADD_1068_U159);
  not ginst224 (ADD_1068_U40, P2_ADDR_REG_16__SCAN_IN);
  not ginst225 (ADD_1068_U41, P1_ADDR_REG_17__SCAN_IN);
  not ginst226 (ADD_1068_U42, P2_ADDR_REG_17__SCAN_IN);
  not ginst227 (ADD_1068_U43, P1_ADDR_REG_18__SCAN_IN);
  not ginst228 (ADD_1068_U44, P2_ADDR_REG_18__SCAN_IN);
  nand ginst229 (ADD_1068_U45, ADD_1068_U149, ADD_1068_U150);
  nand ginst230 (ADD_1068_U46, ADD_1068_U290, ADD_1068_U291);
  nand ginst231 (ADD_1068_U47, ADD_1068_U166, ADD_1068_U167);
  nand ginst232 (ADD_1068_U48, ADD_1068_U173, ADD_1068_U174);
  nand ginst233 (ADD_1068_U49, ADD_1068_U180, ADD_1068_U181);
  nand ginst234 (ADD_1068_U5, ADD_1068_U160, ADD_1068_U220, ADD_1068_U221);
  nand ginst235 (ADD_1068_U50, ADD_1068_U187, ADD_1068_U188);
  nand ginst236 (ADD_1068_U51, ADD_1068_U194, ADD_1068_U195);
  nand ginst237 (ADD_1068_U52, ADD_1068_U201, ADD_1068_U202);
  nand ginst238 (ADD_1068_U53, ADD_1068_U208, ADD_1068_U209);
  nand ginst239 (ADD_1068_U54, ADD_1068_U215, ADD_1068_U216);
  nand ginst240 (ADD_1068_U55, ADD_1068_U232, ADD_1068_U233);
  nand ginst241 (ADD_1068_U56, ADD_1068_U239, ADD_1068_U240);
  nand ginst242 (ADD_1068_U57, ADD_1068_U246, ADD_1068_U247);
  nand ginst243 (ADD_1068_U58, ADD_1068_U253, ADD_1068_U254);
  nand ginst244 (ADD_1068_U59, ADD_1068_U260, ADD_1068_U261);
  not ginst245 (ADD_1068_U6, P1_ADDR_REG_0__SCAN_IN);
  nand ginst246 (ADD_1068_U60, ADD_1068_U267, ADD_1068_U268);
  nand ginst247 (ADD_1068_U61, ADD_1068_U274, ADD_1068_U275);
  nand ginst248 (ADD_1068_U62, ADD_1068_U281, ADD_1068_U282);
  nand ginst249 (ADD_1068_U63, ADD_1068_U288, ADD_1068_U289);
  nand ginst250 (ADD_1068_U64, ADD_1068_U113, ADD_1068_U114);
  nand ginst251 (ADD_1068_U65, ADD_1068_U109, ADD_1068_U110);
  nand ginst252 (ADD_1068_U66, ADD_1068_U105, ADD_1068_U106);
  nand ginst253 (ADD_1068_U67, ADD_1068_U101, ADD_1068_U102);
  nand ginst254 (ADD_1068_U68, ADD_1068_U97, ADD_1068_U98);
  nand ginst255 (ADD_1068_U69, ADD_1068_U93, ADD_1068_U94);
  not ginst256 (ADD_1068_U7, P2_ADDR_REG_0__SCAN_IN);
  nand ginst257 (ADD_1068_U70, ADD_1068_U89, ADD_1068_U90);
  nand ginst258 (ADD_1068_U71, ADD_1068_U72, ADD_1068_U86);
  nand ginst259 (ADD_1068_U72, P1_ADDR_REG_1__SCAN_IN, ADD_1068_U84);
  not ginst260 (ADD_1068_U73, P2_ADDR_REG_19__SCAN_IN);
  not ginst261 (ADD_1068_U74, P1_ADDR_REG_19__SCAN_IN);
  nand ginst262 (ADD_1068_U75, ADD_1068_U145, ADD_1068_U146);
  nand ginst263 (ADD_1068_U76, ADD_1068_U141, ADD_1068_U142);
  nand ginst264 (ADD_1068_U77, ADD_1068_U137, ADD_1068_U138);
  nand ginst265 (ADD_1068_U78, ADD_1068_U133, ADD_1068_U134);
  nand ginst266 (ADD_1068_U79, ADD_1068_U129, ADD_1068_U130);
  not ginst267 (ADD_1068_U8, P2_ADDR_REG_1__SCAN_IN);
  nand ginst268 (ADD_1068_U80, ADD_1068_U125, ADD_1068_U126);
  nand ginst269 (ADD_1068_U81, ADD_1068_U121, ADD_1068_U122);
  nand ginst270 (ADD_1068_U82, ADD_1068_U117, ADD_1068_U118);
  not ginst271 (ADD_1068_U83, ADD_1068_U72);
  not ginst272 (ADD_1068_U84, ADD_1068_U9);
  nand ginst273 (ADD_1068_U85, ADD_1068_U10, ADD_1068_U9);
  nand ginst274 (ADD_1068_U86, P2_ADDR_REG_1__SCAN_IN, ADD_1068_U85);
  not ginst275 (ADD_1068_U87, ADD_1068_U71);
  or ginst276 (ADD_1068_U88, P1_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_2__SCAN_IN);
  nand ginst277 (ADD_1068_U89, ADD_1068_U71, ADD_1068_U88);
  nand ginst278 (ADD_1068_U9, P1_ADDR_REG_0__SCAN_IN, P2_ADDR_REG_0__SCAN_IN);
  nand ginst279 (ADD_1068_U90, P1_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_2__SCAN_IN);
  not ginst280 (ADD_1068_U91, ADD_1068_U70);
  or ginst281 (ADD_1068_U92, P1_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_3__SCAN_IN);
  nand ginst282 (ADD_1068_U93, ADD_1068_U70, ADD_1068_U92);
  nand ginst283 (ADD_1068_U94, P1_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_3__SCAN_IN);
  not ginst284 (ADD_1068_U95, ADD_1068_U69);
  or ginst285 (ADD_1068_U96, P1_ADDR_REG_4__SCAN_IN, P2_ADDR_REG_4__SCAN_IN);
  nand ginst286 (ADD_1068_U97, ADD_1068_U69, ADD_1068_U96);
  nand ginst287 (ADD_1068_U98, P1_ADDR_REG_4__SCAN_IN, P2_ADDR_REG_4__SCAN_IN);
  not ginst288 (ADD_1068_U99, ADD_1068_U68);
  not ginst289 (LT_1075_19_U6, P2_ADDR_REG_19__SCAN_IN);
  not ginst290 (LT_1075_U6, P1_ADDR_REG_19__SCAN_IN);
  not ginst291 (P1_ADD_95_U10, P1_REG3_REG_6__SCAN_IN);
  not ginst292 (P1_ADD_95_U100, P1_ADD_95_U47);
  not ginst293 (P1_ADD_95_U101, P1_ADD_95_U49);
  not ginst294 (P1_ADD_95_U102, P1_ADD_95_U51);
  not ginst295 (P1_ADD_95_U103, P1_ADD_95_U79);
  nand ginst296 (P1_ADD_95_U104, P1_REG3_REG_9__SCAN_IN, P1_ADD_95_U16);
  nand ginst297 (P1_ADD_95_U105, P1_ADD_95_U15, P1_ADD_95_U84);
  nand ginst298 (P1_ADD_95_U106, P1_REG3_REG_8__SCAN_IN, P1_ADD_95_U13);
  nand ginst299 (P1_ADD_95_U107, P1_ADD_95_U14, P1_ADD_95_U83);
  nand ginst300 (P1_ADD_95_U108, P1_REG3_REG_7__SCAN_IN, P1_ADD_95_U11);
  nand ginst301 (P1_ADD_95_U109, P1_ADD_95_U12, P1_ADD_95_U82);
  nand ginst302 (P1_ADD_95_U11, P1_REG3_REG_6__SCAN_IN, P1_ADD_95_U81);
  nand ginst303 (P1_ADD_95_U110, P1_REG3_REG_6__SCAN_IN, P1_ADD_95_U9);
  nand ginst304 (P1_ADD_95_U111, P1_ADD_95_U10, P1_ADD_95_U81);
  nand ginst305 (P1_ADD_95_U112, P1_REG3_REG_5__SCAN_IN, P1_ADD_95_U7);
  nand ginst306 (P1_ADD_95_U113, P1_ADD_95_U8, P1_ADD_95_U80);
  nand ginst307 (P1_ADD_95_U114, P1_REG3_REG_4__SCAN_IN, P1_ADD_95_U4);
  nand ginst308 (P1_ADD_95_U115, P1_REG3_REG_3__SCAN_IN, P1_ADD_95_U6);
  nand ginst309 (P1_ADD_95_U116, P1_REG3_REG_28__SCAN_IN, P1_ADD_95_U79);
  nand ginst310 (P1_ADD_95_U117, P1_ADD_95_U103, P1_ADD_95_U52);
  nand ginst311 (P1_ADD_95_U118, P1_REG3_REG_27__SCAN_IN, P1_ADD_95_U51);
  nand ginst312 (P1_ADD_95_U119, P1_ADD_95_U102, P1_ADD_95_U53);
  not ginst313 (P1_ADD_95_U12, P1_REG3_REG_7__SCAN_IN);
  nand ginst314 (P1_ADD_95_U120, P1_REG3_REG_26__SCAN_IN, P1_ADD_95_U49);
  nand ginst315 (P1_ADD_95_U121, P1_ADD_95_U101, P1_ADD_95_U50);
  nand ginst316 (P1_ADD_95_U122, P1_REG3_REG_25__SCAN_IN, P1_ADD_95_U47);
  nand ginst317 (P1_ADD_95_U123, P1_ADD_95_U100, P1_ADD_95_U48);
  nand ginst318 (P1_ADD_95_U124, P1_REG3_REG_24__SCAN_IN, P1_ADD_95_U45);
  nand ginst319 (P1_ADD_95_U125, P1_ADD_95_U46, P1_ADD_95_U99);
  nand ginst320 (P1_ADD_95_U126, P1_REG3_REG_23__SCAN_IN, P1_ADD_95_U43);
  nand ginst321 (P1_ADD_95_U127, P1_ADD_95_U44, P1_ADD_95_U98);
  nand ginst322 (P1_ADD_95_U128, P1_REG3_REG_22__SCAN_IN, P1_ADD_95_U41);
  nand ginst323 (P1_ADD_95_U129, P1_ADD_95_U42, P1_ADD_95_U97);
  nand ginst324 (P1_ADD_95_U13, P1_REG3_REG_7__SCAN_IN, P1_ADD_95_U82);
  nand ginst325 (P1_ADD_95_U130, P1_REG3_REG_21__SCAN_IN, P1_ADD_95_U39);
  nand ginst326 (P1_ADD_95_U131, P1_ADD_95_U40, P1_ADD_95_U96);
  nand ginst327 (P1_ADD_95_U132, P1_REG3_REG_20__SCAN_IN, P1_ADD_95_U37);
  nand ginst328 (P1_ADD_95_U133, P1_ADD_95_U38, P1_ADD_95_U95);
  nand ginst329 (P1_ADD_95_U134, P1_REG3_REG_19__SCAN_IN, P1_ADD_95_U35);
  nand ginst330 (P1_ADD_95_U135, P1_ADD_95_U36, P1_ADD_95_U94);
  nand ginst331 (P1_ADD_95_U136, P1_REG3_REG_18__SCAN_IN, P1_ADD_95_U33);
  nand ginst332 (P1_ADD_95_U137, P1_ADD_95_U34, P1_ADD_95_U93);
  nand ginst333 (P1_ADD_95_U138, P1_REG3_REG_17__SCAN_IN, P1_ADD_95_U31);
  nand ginst334 (P1_ADD_95_U139, P1_ADD_95_U32, P1_ADD_95_U92);
  not ginst335 (P1_ADD_95_U14, P1_REG3_REG_8__SCAN_IN);
  nand ginst336 (P1_ADD_95_U140, P1_REG3_REG_16__SCAN_IN, P1_ADD_95_U29);
  nand ginst337 (P1_ADD_95_U141, P1_ADD_95_U30, P1_ADD_95_U91);
  nand ginst338 (P1_ADD_95_U142, P1_REG3_REG_15__SCAN_IN, P1_ADD_95_U27);
  nand ginst339 (P1_ADD_95_U143, P1_ADD_95_U28, P1_ADD_95_U90);
  nand ginst340 (P1_ADD_95_U144, P1_REG3_REG_14__SCAN_IN, P1_ADD_95_U25);
  nand ginst341 (P1_ADD_95_U145, P1_ADD_95_U26, P1_ADD_95_U89);
  nand ginst342 (P1_ADD_95_U146, P1_REG3_REG_13__SCAN_IN, P1_ADD_95_U23);
  nand ginst343 (P1_ADD_95_U147, P1_ADD_95_U24, P1_ADD_95_U88);
  nand ginst344 (P1_ADD_95_U148, P1_REG3_REG_12__SCAN_IN, P1_ADD_95_U21);
  nand ginst345 (P1_ADD_95_U149, P1_ADD_95_U22, P1_ADD_95_U87);
  not ginst346 (P1_ADD_95_U15, P1_REG3_REG_9__SCAN_IN);
  nand ginst347 (P1_ADD_95_U150, P1_REG3_REG_11__SCAN_IN, P1_ADD_95_U19);
  nand ginst348 (P1_ADD_95_U151, P1_ADD_95_U20, P1_ADD_95_U86);
  nand ginst349 (P1_ADD_95_U152, P1_REG3_REG_10__SCAN_IN, P1_ADD_95_U17);
  nand ginst350 (P1_ADD_95_U153, P1_ADD_95_U18, P1_ADD_95_U85);
  nand ginst351 (P1_ADD_95_U16, P1_REG3_REG_8__SCAN_IN, P1_ADD_95_U83);
  nand ginst352 (P1_ADD_95_U17, P1_REG3_REG_9__SCAN_IN, P1_ADD_95_U84);
  not ginst353 (P1_ADD_95_U18, P1_REG3_REG_10__SCAN_IN);
  nand ginst354 (P1_ADD_95_U19, P1_REG3_REG_10__SCAN_IN, P1_ADD_95_U85);
  not ginst355 (P1_ADD_95_U20, P1_REG3_REG_11__SCAN_IN);
  nand ginst356 (P1_ADD_95_U21, P1_REG3_REG_11__SCAN_IN, P1_ADD_95_U86);
  not ginst357 (P1_ADD_95_U22, P1_REG3_REG_12__SCAN_IN);
  nand ginst358 (P1_ADD_95_U23, P1_REG3_REG_12__SCAN_IN, P1_ADD_95_U87);
  not ginst359 (P1_ADD_95_U24, P1_REG3_REG_13__SCAN_IN);
  nand ginst360 (P1_ADD_95_U25, P1_REG3_REG_13__SCAN_IN, P1_ADD_95_U88);
  not ginst361 (P1_ADD_95_U26, P1_REG3_REG_14__SCAN_IN);
  nand ginst362 (P1_ADD_95_U27, P1_REG3_REG_14__SCAN_IN, P1_ADD_95_U89);
  not ginst363 (P1_ADD_95_U28, P1_REG3_REG_15__SCAN_IN);
  nand ginst364 (P1_ADD_95_U29, P1_REG3_REG_15__SCAN_IN, P1_ADD_95_U90);
  not ginst365 (P1_ADD_95_U30, P1_REG3_REG_16__SCAN_IN);
  nand ginst366 (P1_ADD_95_U31, P1_REG3_REG_16__SCAN_IN, P1_ADD_95_U91);
  not ginst367 (P1_ADD_95_U32, P1_REG3_REG_17__SCAN_IN);
  nand ginst368 (P1_ADD_95_U33, P1_REG3_REG_17__SCAN_IN, P1_ADD_95_U92);
  not ginst369 (P1_ADD_95_U34, P1_REG3_REG_18__SCAN_IN);
  nand ginst370 (P1_ADD_95_U35, P1_REG3_REG_18__SCAN_IN, P1_ADD_95_U93);
  not ginst371 (P1_ADD_95_U36, P1_REG3_REG_19__SCAN_IN);
  nand ginst372 (P1_ADD_95_U37, P1_REG3_REG_19__SCAN_IN, P1_ADD_95_U94);
  not ginst373 (P1_ADD_95_U38, P1_REG3_REG_20__SCAN_IN);
  nand ginst374 (P1_ADD_95_U39, P1_REG3_REG_20__SCAN_IN, P1_ADD_95_U95);
  not ginst375 (P1_ADD_95_U4, P1_REG3_REG_3__SCAN_IN);
  not ginst376 (P1_ADD_95_U40, P1_REG3_REG_21__SCAN_IN);
  nand ginst377 (P1_ADD_95_U41, P1_REG3_REG_21__SCAN_IN, P1_ADD_95_U96);
  not ginst378 (P1_ADD_95_U42, P1_REG3_REG_22__SCAN_IN);
  nand ginst379 (P1_ADD_95_U43, P1_REG3_REG_22__SCAN_IN, P1_ADD_95_U97);
  not ginst380 (P1_ADD_95_U44, P1_REG3_REG_23__SCAN_IN);
  nand ginst381 (P1_ADD_95_U45, P1_REG3_REG_23__SCAN_IN, P1_ADD_95_U98);
  not ginst382 (P1_ADD_95_U46, P1_REG3_REG_24__SCAN_IN);
  nand ginst383 (P1_ADD_95_U47, P1_REG3_REG_24__SCAN_IN, P1_ADD_95_U99);
  not ginst384 (P1_ADD_95_U48, P1_REG3_REG_25__SCAN_IN);
  nand ginst385 (P1_ADD_95_U49, P1_REG3_REG_25__SCAN_IN, P1_ADD_95_U100);
  and ginst386 (P1_ADD_95_U5, P1_REG3_REG_28__SCAN_IN, P1_REG3_REG_27__SCAN_IN, P1_ADD_95_U102);
  not ginst387 (P1_ADD_95_U50, P1_REG3_REG_26__SCAN_IN);
  nand ginst388 (P1_ADD_95_U51, P1_REG3_REG_26__SCAN_IN, P1_ADD_95_U101);
  not ginst389 (P1_ADD_95_U52, P1_REG3_REG_28__SCAN_IN);
  not ginst390 (P1_ADD_95_U53, P1_REG3_REG_27__SCAN_IN);
  nand ginst391 (P1_ADD_95_U54, P1_ADD_95_U104, P1_ADD_95_U105);
  nand ginst392 (P1_ADD_95_U55, P1_ADD_95_U106, P1_ADD_95_U107);
  nand ginst393 (P1_ADD_95_U56, P1_ADD_95_U108, P1_ADD_95_U109);
  nand ginst394 (P1_ADD_95_U57, P1_ADD_95_U110, P1_ADD_95_U111);
  nand ginst395 (P1_ADD_95_U58, P1_ADD_95_U112, P1_ADD_95_U113);
  nand ginst396 (P1_ADD_95_U59, P1_ADD_95_U114, P1_ADD_95_U115);
  not ginst397 (P1_ADD_95_U6, P1_REG3_REG_4__SCAN_IN);
  nand ginst398 (P1_ADD_95_U60, P1_ADD_95_U116, P1_ADD_95_U117);
  nand ginst399 (P1_ADD_95_U61, P1_ADD_95_U118, P1_ADD_95_U119);
  nand ginst400 (P1_ADD_95_U62, P1_ADD_95_U120, P1_ADD_95_U121);
  nand ginst401 (P1_ADD_95_U63, P1_ADD_95_U122, P1_ADD_95_U123);
  nand ginst402 (P1_ADD_95_U64, P1_ADD_95_U124, P1_ADD_95_U125);
  nand ginst403 (P1_ADD_95_U65, P1_ADD_95_U126, P1_ADD_95_U127);
  nand ginst404 (P1_ADD_95_U66, P1_ADD_95_U128, P1_ADD_95_U129);
  nand ginst405 (P1_ADD_95_U67, P1_ADD_95_U130, P1_ADD_95_U131);
  nand ginst406 (P1_ADD_95_U68, P1_ADD_95_U132, P1_ADD_95_U133);
  nand ginst407 (P1_ADD_95_U69, P1_ADD_95_U134, P1_ADD_95_U135);
  nand ginst408 (P1_ADD_95_U7, P1_REG3_REG_4__SCAN_IN, P1_REG3_REG_3__SCAN_IN);
  nand ginst409 (P1_ADD_95_U70, P1_ADD_95_U136, P1_ADD_95_U137);
  nand ginst410 (P1_ADD_95_U71, P1_ADD_95_U138, P1_ADD_95_U139);
  nand ginst411 (P1_ADD_95_U72, P1_ADD_95_U140, P1_ADD_95_U141);
  nand ginst412 (P1_ADD_95_U73, P1_ADD_95_U142, P1_ADD_95_U143);
  nand ginst413 (P1_ADD_95_U74, P1_ADD_95_U144, P1_ADD_95_U145);
  nand ginst414 (P1_ADD_95_U75, P1_ADD_95_U146, P1_ADD_95_U147);
  nand ginst415 (P1_ADD_95_U76, P1_ADD_95_U148, P1_ADD_95_U149);
  nand ginst416 (P1_ADD_95_U77, P1_ADD_95_U150, P1_ADD_95_U151);
  nand ginst417 (P1_ADD_95_U78, P1_ADD_95_U152, P1_ADD_95_U153);
  nand ginst418 (P1_ADD_95_U79, P1_REG3_REG_27__SCAN_IN, P1_ADD_95_U102);
  not ginst419 (P1_ADD_95_U8, P1_REG3_REG_5__SCAN_IN);
  not ginst420 (P1_ADD_95_U80, P1_ADD_95_U7);
  not ginst421 (P1_ADD_95_U81, P1_ADD_95_U9);
  not ginst422 (P1_ADD_95_U82, P1_ADD_95_U11);
  not ginst423 (P1_ADD_95_U83, P1_ADD_95_U13);
  not ginst424 (P1_ADD_95_U84, P1_ADD_95_U16);
  not ginst425 (P1_ADD_95_U85, P1_ADD_95_U17);
  not ginst426 (P1_ADD_95_U86, P1_ADD_95_U19);
  not ginst427 (P1_ADD_95_U87, P1_ADD_95_U21);
  not ginst428 (P1_ADD_95_U88, P1_ADD_95_U23);
  not ginst429 (P1_ADD_95_U89, P1_ADD_95_U25);
  nand ginst430 (P1_ADD_95_U9, P1_REG3_REG_5__SCAN_IN, P1_ADD_95_U80);
  not ginst431 (P1_ADD_95_U90, P1_ADD_95_U27);
  not ginst432 (P1_ADD_95_U91, P1_ADD_95_U29);
  not ginst433 (P1_ADD_95_U92, P1_ADD_95_U31);
  not ginst434 (P1_ADD_95_U93, P1_ADD_95_U33);
  not ginst435 (P1_ADD_95_U94, P1_ADD_95_U35);
  not ginst436 (P1_ADD_95_U95, P1_ADD_95_U37);
  not ginst437 (P1_ADD_95_U96, P1_ADD_95_U39);
  not ginst438 (P1_ADD_95_U97, P1_ADD_95_U41);
  not ginst439 (P1_ADD_95_U98, P1_ADD_95_U43);
  not ginst440 (P1_ADD_95_U99, P1_ADD_95_U45);
  and ginst441 (P1_LT_197_U10, P1_LT_197_U128, P1_LT_197_U131, P1_LT_197_U84, P1_LT_197_U85);
  and ginst442 (P1_LT_197_U100, P1_LT_197_U178, P1_LT_197_U179);
  and ginst443 (P1_LT_197_U101, P1_LT_197_U181, P1_LT_197_U182);
  and ginst444 (P1_LT_197_U102, P1_LT_197_U65, P1_U3602);
  and ginst445 (P1_LT_197_U103, P1_LT_197_U185, P1_LT_197_U186);
  and ginst446 (P1_LT_197_U104, P1_LT_197_U125, P1_LT_197_U189);
  and ginst447 (P1_LT_197_U105, P1_LT_197_U195, P1_LT_197_U196);
  and ginst448 (P1_LT_197_U106, P1_LT_197_U73, P1_U3596);
  and ginst449 (P1_LT_197_U107, P1_LT_197_U112, P1_LT_197_U198);
  not ginst450 (P1_LT_197_U108, P1_U3617);
  nand ginst451 (P1_LT_197_U109, P1_LT_197_U107, P1_LT_197_U197);
  and ginst452 (P1_LT_197_U11, P1_LT_197_U144, P1_LT_197_U145);
  nand ginst453 (P1_LT_197_U110, P1_LT_197_U16, P1_U3984);
  nand ginst454 (P1_LT_197_U111, P1_LT_197_U14, P1_U3593);
  nand ginst455 (P1_LT_197_U112, P1_LT_197_U111, P1_LT_197_U75, P1_U3594);
  nand ginst456 (P1_LT_197_U113, P1_LT_197_U14, P1_U3593);
  nand ginst457 (P1_LT_197_U114, P1_LT_197_U70, P1_U3598);
  nand ginst458 (P1_LT_197_U115, P1_LT_197_U29, P1_U3508);
  nand ginst459 (P1_LT_197_U116, P1_LT_197_U26, P1_U3506);
  nand ginst460 (P1_LT_197_U117, P1_LT_197_U64, P1_U3603);
  nand ginst461 (P1_LT_197_U118, P1_LT_197_U22, P1_U3604);
  nand ginst462 (P1_LT_197_U119, P1_LT_197_U115, P1_LT_197_U79);
  and ginst463 (P1_LT_197_U12, P1_LT_197_U193, P1_LT_197_U72);
  nand ginst464 (P1_LT_197_U120, P1_LT_197_U6, P1_LT_197_U80);
  nand ginst465 (P1_LT_197_U121, P1_LT_197_U25, P1_U3607);
  nand ginst466 (P1_LT_197_U122, P1_LT_197_U24, P1_U3605);
  nand ginst467 (P1_LT_197_U123, P1_LT_197_U32, P1_U3610);
  nand ginst468 (P1_LT_197_U124, P1_LT_197_U67, P1_U3978);
  nand ginst469 (P1_LT_197_U125, P1_LT_197_U68, P1_U3977);
  nand ginst470 (P1_LT_197_U126, P1_LT_197_U63, P1_U3611);
  nand ginst471 (P1_LT_197_U127, P1_LT_197_U42, P1_U3473);
  nand ginst472 (P1_LT_197_U128, P1_LT_197_U127, P1_LT_197_U82);
  nand ginst473 (P1_LT_197_U129, P1_LT_197_U36, P1_U3470);
  and ginst474 (P1_LT_197_U13, P1_LT_197_U199, P1_LT_197_U200);
  nand ginst475 (P1_LT_197_U130, P1_LT_197_U42, P1_U3473);
  nand ginst476 (P1_LT_197_U131, P1_LT_197_U83, P1_LT_197_U9);
  nand ginst477 (P1_LT_197_U132, P1_LT_197_U55, P1_U3586);
  nand ginst478 (P1_LT_197_U133, P1_LT_197_U56, P1_U3616);
  nand ginst479 (P1_LT_197_U134, P1_LT_197_U54, P1_U3587);
  nand ginst480 (P1_LT_197_U135, P1_LT_197_U35, P1_U3588);
  nand ginst481 (P1_LT_197_U136, P1_LT_197_U52, P1_U3591);
  nand ginst482 (P1_LT_197_U137, P1_LT_197_U51, P1_U3592);
  not ginst483 (P1_LT_197_U138, P1_LT_197_U45);
  nand ginst484 (P1_LT_197_U139, P1_LT_197_U138, P1_U3455);
  not ginst485 (P1_LT_197_U14, P1_U3983);
  nand ginst486 (P1_LT_197_U140, P1_LT_197_U139, P1_U3606);
  nand ginst487 (P1_LT_197_U141, P1_LT_197_U45, P1_LT_197_U46);
  nand ginst488 (P1_LT_197_U142, P1_LT_197_U50, P1_U3595);
  nand ginst489 (P1_LT_197_U143, P1_LT_197_U10, P1_LT_197_U87);
  nand ginst490 (P1_LT_197_U144, P1_LT_197_U58, P1_U3488);
  nand ginst491 (P1_LT_197_U145, P1_LT_197_U61, P1_U3491);
  nand ginst492 (P1_LT_197_U146, P1_LT_197_U136, P1_LT_197_U89);
  nand ginst493 (P1_LT_197_U147, P1_LT_197_U43, P1_U3464);
  nand ginst494 (P1_LT_197_U148, P1_LT_197_U146, P1_LT_197_U147, P1_LT_197_U9);
  nand ginst495 (P1_LT_197_U149, P1_LT_197_U131, P1_LT_197_U148);
  not ginst496 (P1_LT_197_U15, P1_U3593);
  nand ginst497 (P1_LT_197_U150, P1_LT_197_U38, P1_U3467);
  nand ginst498 (P1_LT_197_U151, P1_LT_197_U149, P1_LT_197_U150);
  nand ginst499 (P1_LT_197_U152, P1_LT_197_U151, P1_LT_197_U90);
  nand ginst500 (P1_LT_197_U153, P1_LT_197_U41, P1_U3476);
  nand ginst501 (P1_LT_197_U154, P1_LT_197_U152, P1_LT_197_U153);
  nand ginst502 (P1_LT_197_U155, P1_LT_197_U132, P1_LT_197_U154);
  nand ginst503 (P1_LT_197_U156, P1_LT_197_U39, P1_U3479);
  nand ginst504 (P1_LT_197_U157, P1_LT_197_U155, P1_LT_197_U156);
  nand ginst505 (P1_LT_197_U158, P1_LT_197_U10, P1_LT_197_U88);
  nand ginst506 (P1_LT_197_U159, P1_LT_197_U133, P1_LT_197_U157);
  not ginst507 (P1_LT_197_U16, P1_U3594);
  nand ginst508 (P1_LT_197_U160, P1_LT_197_U40, P1_U3482);
  nand ginst509 (P1_LT_197_U161, P1_LT_197_U59, P1_U3485);
  nand ginst510 (P1_LT_197_U162, P1_LT_197_U159, P1_LT_197_U91);
  nand ginst511 (P1_LT_197_U163, P1_LT_197_U61, P1_U3491);
  nand ginst512 (P1_LT_197_U164, P1_LT_197_U163, P1_LT_197_U94);
  nand ginst513 (P1_LT_197_U165, P1_LT_197_U11, P1_LT_197_U95);
  nand ginst514 (P1_LT_197_U166, P1_LT_197_U62, P1_U3612);
  nand ginst515 (P1_LT_197_U167, P1_LT_197_U49, P1_U3613);
  nand ginst516 (P1_LT_197_U168, P1_LT_197_U162, P1_LT_197_U97);
  nand ginst517 (P1_LT_197_U169, P1_LT_197_U60, P1_U3494);
  not ginst518 (P1_LT_197_U17, P1_U3598);
  nand ginst519 (P1_LT_197_U170, P1_LT_197_U168, P1_LT_197_U169);
  nand ginst520 (P1_LT_197_U171, P1_LT_197_U126, P1_LT_197_U170);
  nand ginst521 (P1_LT_197_U172, P1_LT_197_U34, P1_U3497);
  nand ginst522 (P1_LT_197_U173, P1_LT_197_U171, P1_LT_197_U172);
  nand ginst523 (P1_LT_197_U174, P1_LT_197_U28, P1_U3503);
  nand ginst524 (P1_LT_197_U175, P1_LT_197_U33, P1_U3500);
  nand ginst525 (P1_LT_197_U176, P1_LT_197_U6, P1_LT_197_U78);
  nand ginst526 (P1_LT_197_U177, P1_LT_197_U117, P1_LT_197_U76);
  nand ginst527 (P1_LT_197_U178, P1_LT_197_U7, P1_LT_197_U77);
  nand ginst528 (P1_LT_197_U179, P1_LT_197_U176, P1_LT_197_U8);
  not ginst529 (P1_LT_197_U18, P1_U3599);
  nand ginst530 (P1_LT_197_U180, P1_LT_197_U123, P1_LT_197_U173, P1_LT_197_U8);
  nand ginst531 (P1_LT_197_U181, P1_LT_197_U21, P1_U3980);
  nand ginst532 (P1_LT_197_U182, P1_LT_197_U66, P1_U3979);
  nand ginst533 (P1_LT_197_U183, P1_LT_197_U100, P1_LT_197_U101, P1_LT_197_U180, P1_LT_197_U99);
  nand ginst534 (P1_LT_197_U184, P1_LT_197_U102, P1_LT_197_U124);
  nand ginst535 (P1_LT_197_U185, P1_LT_197_U20, P1_U3601);
  nand ginst536 (P1_LT_197_U186, P1_LT_197_U19, P1_U3600);
  nand ginst537 (P1_LT_197_U187, P1_LT_197_U69, P1_U3599);
  nand ginst538 (P1_LT_197_U188, P1_LT_197_U103, P1_LT_197_U183, P1_LT_197_U184);
  nand ginst539 (P1_LT_197_U189, P1_LT_197_U18, P1_U3976);
  not ginst540 (P1_LT_197_U19, P1_U3977);
  nand ginst541 (P1_LT_197_U190, P1_LT_197_U104, P1_LT_197_U188);
  nand ginst542 (P1_LT_197_U191, P1_LT_197_U114, P1_LT_197_U187, P1_LT_197_U190);
  nand ginst543 (P1_LT_197_U192, P1_LT_197_U17, P1_U3975);
  not ginst544 (P1_LT_197_U193, P1_LT_197_U71);
  or ginst545 (P1_LT_197_U194, P1_LT_197_U12, P1_U3597);
  nand ginst546 (P1_LT_197_U195, P1_LT_197_U71, P1_U3974);
  nand ginst547 (P1_LT_197_U196, P1_LT_197_U74, P1_U3985);
  nand ginst548 (P1_LT_197_U197, P1_LT_197_U105, P1_LT_197_U113, P1_LT_197_U194);
  nand ginst549 (P1_LT_197_U198, P1_LT_197_U106, P1_LT_197_U113);
  nand ginst550 (P1_LT_197_U199, P1_LT_197_U15, P1_U3983);
  not ginst551 (P1_LT_197_U20, P1_U3978);
  nand ginst552 (P1_LT_197_U200, P1_LT_197_U109, P1_LT_197_U110);
  not ginst553 (P1_LT_197_U21, P1_U3603);
  not ginst554 (P1_LT_197_U22, P1_U3981);
  not ginst555 (P1_LT_197_U23, P1_U3604);
  not ginst556 (P1_LT_197_U24, P1_U3982);
  not ginst557 (P1_LT_197_U25, P1_U3508);
  not ginst558 (P1_LT_197_U26, P1_U3608);
  not ginst559 (P1_LT_197_U27, P1_U3506);
  not ginst560 (P1_LT_197_U28, P1_U3609);
  not ginst561 (P1_LT_197_U29, P1_U3607);
  not ginst562 (P1_LT_197_U30, P1_U3605);
  not ginst563 (P1_LT_197_U31, P1_U3503);
  not ginst564 (P1_LT_197_U32, P1_U3500);
  not ginst565 (P1_LT_197_U33, P1_U3610);
  not ginst566 (P1_LT_197_U34, P1_U3611);
  not ginst567 (P1_LT_197_U35, P1_U3473);
  not ginst568 (P1_LT_197_U36, P1_U3589);
  not ginst569 (P1_LT_197_U37, P1_U3470);
  not ginst570 (P1_LT_197_U38, P1_U3590);
  not ginst571 (P1_LT_197_U39, P1_U3586);
  not ginst572 (P1_LT_197_U40, P1_U3616);
  not ginst573 (P1_LT_197_U41, P1_U3587);
  not ginst574 (P1_LT_197_U42, P1_U3588);
  not ginst575 (P1_LT_197_U43, P1_U3591);
  not ginst576 (P1_LT_197_U44, P1_U3592);
  nand ginst577 (P1_LT_197_U45, P1_LT_197_U108, P1_U3450);
  not ginst578 (P1_LT_197_U46, P1_U3455);
  not ginst579 (P1_LT_197_U47, P1_U3595);
  not ginst580 (P1_LT_197_U48, P1_U3488);
  not ginst581 (P1_LT_197_U49, P1_U3491);
  not ginst582 (P1_LT_197_U50, P1_U3458);
  not ginst583 (P1_LT_197_U51, P1_U3461);
  not ginst584 (P1_LT_197_U52, P1_U3464);
  not ginst585 (P1_LT_197_U53, P1_U3467);
  not ginst586 (P1_LT_197_U54, P1_U3476);
  not ginst587 (P1_LT_197_U55, P1_U3479);
  not ginst588 (P1_LT_197_U56, P1_U3482);
  not ginst589 (P1_LT_197_U57, P1_U3485);
  not ginst590 (P1_LT_197_U58, P1_U3614);
  not ginst591 (P1_LT_197_U59, P1_U3615);
  and ginst592 (P1_LT_197_U6, P1_LT_197_U115, P1_LT_197_U116);
  not ginst593 (P1_LT_197_U60, P1_U3612);
  not ginst594 (P1_LT_197_U61, P1_U3613);
  not ginst595 (P1_LT_197_U62, P1_U3494);
  not ginst596 (P1_LT_197_U63, P1_U3497);
  not ginst597 (P1_LT_197_U64, P1_U3980);
  not ginst598 (P1_LT_197_U65, P1_U3979);
  not ginst599 (P1_LT_197_U66, P1_U3602);
  not ginst600 (P1_LT_197_U67, P1_U3601);
  not ginst601 (P1_LT_197_U68, P1_U3600);
  not ginst602 (P1_LT_197_U69, P1_U3976);
  and ginst603 (P1_LT_197_U7, P1_LT_197_U117, P1_LT_197_U118);
  not ginst604 (P1_LT_197_U70, P1_U3975);
  nand ginst605 (P1_LT_197_U71, P1_LT_197_U191, P1_LT_197_U192);
  not ginst606 (P1_LT_197_U72, P1_U3974);
  not ginst607 (P1_LT_197_U73, P1_U3985);
  not ginst608 (P1_LT_197_U74, P1_U3596);
  not ginst609 (P1_LT_197_U75, P1_U3984);
  and ginst610 (P1_LT_197_U76, P1_LT_197_U23, P1_U3981);
  and ginst611 (P1_LT_197_U77, P1_LT_197_U30, P1_U3982);
  and ginst612 (P1_LT_197_U78, P1_LT_197_U174, P1_LT_197_U175);
  and ginst613 (P1_LT_197_U79, P1_LT_197_U27, P1_U3608);
  and ginst614 (P1_LT_197_U8, P1_LT_197_U120, P1_LT_197_U122, P1_LT_197_U7, P1_LT_197_U81);
  and ginst615 (P1_LT_197_U80, P1_LT_197_U31, P1_U3609);
  and ginst616 (P1_LT_197_U81, P1_LT_197_U119, P1_LT_197_U121);
  and ginst617 (P1_LT_197_U82, P1_LT_197_U37, P1_U3589);
  and ginst618 (P1_LT_197_U83, P1_LT_197_U53, P1_U3590);
  and ginst619 (P1_LT_197_U84, P1_LT_197_U132, P1_LT_197_U133);
  and ginst620 (P1_LT_197_U85, P1_LT_197_U134, P1_LT_197_U135, P1_LT_197_U136, P1_LT_197_U137);
  and ginst621 (P1_LT_197_U86, P1_LT_197_U141, P1_LT_197_U142);
  and ginst622 (P1_LT_197_U87, P1_LT_197_U140, P1_LT_197_U86);
  and ginst623 (P1_LT_197_U88, P1_LT_197_U47, P1_U3458);
  and ginst624 (P1_LT_197_U89, P1_LT_197_U44, P1_U3461);
  and ginst625 (P1_LT_197_U9, P1_LT_197_U129, P1_LT_197_U130);
  and ginst626 (P1_LT_197_U90, P1_LT_197_U128, P1_LT_197_U134, P1_LT_197_U135);
  and ginst627 (P1_LT_197_U91, P1_LT_197_U143, P1_LT_197_U158, P1_LT_197_U93);
  and ginst628 (P1_LT_197_U92, P1_LT_197_U160, P1_LT_197_U161);
  and ginst629 (P1_LT_197_U93, P1_LT_197_U11, P1_LT_197_U92);
  and ginst630 (P1_LT_197_U94, P1_LT_197_U48, P1_U3614);
  and ginst631 (P1_LT_197_U95, P1_LT_197_U57, P1_U3615);
  and ginst632 (P1_LT_197_U96, P1_LT_197_U164, P1_LT_197_U98);
  and ginst633 (P1_LT_197_U97, P1_LT_197_U165, P1_LT_197_U96);
  and ginst634 (P1_LT_197_U98, P1_LT_197_U166, P1_LT_197_U167);
  and ginst635 (P1_LT_197_U99, P1_LT_197_U124, P1_LT_197_U177);
  and ginst636 (P1_R1105_U10, P1_R1105_U215, P1_R1105_U218);
  not ginst637 (P1_R1105_U100, P1_R1105_U40);
  not ginst638 (P1_R1105_U101, P1_R1105_U41);
  nand ginst639 (P1_R1105_U102, P1_R1105_U40, P1_R1105_U41);
  nand ginst640 (P1_R1105_U103, P1_REG2_REG_2__SCAN_IN, P1_R1105_U96, P1_U3457);
  nand ginst641 (P1_R1105_U104, P1_R1105_U102, P1_R1105_U5);
  nand ginst642 (P1_R1105_U105, P1_REG2_REG_3__SCAN_IN, P1_U3460);
  nand ginst643 (P1_R1105_U106, P1_R1105_U103, P1_R1105_U104, P1_R1105_U105);
  nand ginst644 (P1_R1105_U107, P1_R1105_U32, P1_R1105_U33);
  nand ginst645 (P1_R1105_U108, P1_R1105_U107, P1_U3466);
  nand ginst646 (P1_R1105_U109, P1_R1105_U106, P1_R1105_U4);
  and ginst647 (P1_R1105_U11, P1_R1105_U208, P1_R1105_U211);
  nand ginst648 (P1_R1105_U110, P1_REG2_REG_5__SCAN_IN, P1_R1105_U89);
  not ginst649 (P1_R1105_U111, P1_R1105_U39);
  or ginst650 (P1_R1105_U112, P1_REG2_REG_7__SCAN_IN, P1_U3472);
  or ginst651 (P1_R1105_U113, P1_REG2_REG_6__SCAN_IN, P1_U3469);
  not ginst652 (P1_R1105_U114, P1_R1105_U20);
  nand ginst653 (P1_R1105_U115, P1_R1105_U20, P1_R1105_U21);
  nand ginst654 (P1_R1105_U116, P1_R1105_U115, P1_U3472);
  nand ginst655 (P1_R1105_U117, P1_REG2_REG_7__SCAN_IN, P1_R1105_U114);
  nand ginst656 (P1_R1105_U118, P1_R1105_U39, P1_R1105_U6);
  not ginst657 (P1_R1105_U119, P1_R1105_U81);
  and ginst658 (P1_R1105_U12, P1_R1105_U199, P1_R1105_U202);
  or ginst659 (P1_R1105_U120, P1_REG2_REG_8__SCAN_IN, P1_U3475);
  nand ginst660 (P1_R1105_U121, P1_R1105_U120, P1_R1105_U81);
  not ginst661 (P1_R1105_U122, P1_R1105_U38);
  or ginst662 (P1_R1105_U123, P1_REG2_REG_9__SCAN_IN, P1_U3478);
  or ginst663 (P1_R1105_U124, P1_REG2_REG_6__SCAN_IN, P1_U3469);
  nand ginst664 (P1_R1105_U125, P1_R1105_U124, P1_R1105_U39);
  nand ginst665 (P1_R1105_U126, P1_R1105_U125, P1_R1105_U20, P1_R1105_U237, P1_R1105_U238);
  nand ginst666 (P1_R1105_U127, P1_R1105_U111, P1_R1105_U20);
  nand ginst667 (P1_R1105_U128, P1_REG2_REG_7__SCAN_IN, P1_U3472);
  nand ginst668 (P1_R1105_U129, P1_R1105_U127, P1_R1105_U128, P1_R1105_U6);
  and ginst669 (P1_R1105_U13, P1_R1105_U192, P1_R1105_U196);
  or ginst670 (P1_R1105_U130, P1_REG2_REG_6__SCAN_IN, P1_U3469);
  nand ginst671 (P1_R1105_U131, P1_R1105_U101, P1_R1105_U97);
  nand ginst672 (P1_R1105_U132, P1_REG2_REG_2__SCAN_IN, P1_U3457);
  not ginst673 (P1_R1105_U133, P1_R1105_U43);
  nand ginst674 (P1_R1105_U134, P1_R1105_U100, P1_R1105_U5);
  nand ginst675 (P1_R1105_U135, P1_R1105_U43, P1_R1105_U96);
  nand ginst676 (P1_R1105_U136, P1_REG2_REG_3__SCAN_IN, P1_U3460);
  not ginst677 (P1_R1105_U137, P1_R1105_U42);
  or ginst678 (P1_R1105_U138, P1_REG2_REG_4__SCAN_IN, P1_U3463);
  nand ginst679 (P1_R1105_U139, P1_R1105_U138, P1_R1105_U42);
  and ginst680 (P1_R1105_U14, P1_R1105_U148, P1_R1105_U151);
  nand ginst681 (P1_R1105_U140, P1_R1105_U139, P1_R1105_U244, P1_R1105_U245, P1_R1105_U32);
  nand ginst682 (P1_R1105_U141, P1_R1105_U137, P1_R1105_U32);
  nand ginst683 (P1_R1105_U142, P1_REG2_REG_5__SCAN_IN, P1_U3466);
  nand ginst684 (P1_R1105_U143, P1_R1105_U141, P1_R1105_U142, P1_R1105_U4);
  or ginst685 (P1_R1105_U144, P1_REG2_REG_4__SCAN_IN, P1_U3463);
  nand ginst686 (P1_R1105_U145, P1_R1105_U100, P1_R1105_U97);
  not ginst687 (P1_R1105_U146, P1_R1105_U82);
  nand ginst688 (P1_R1105_U147, P1_REG2_REG_3__SCAN_IN, P1_U3460);
  nand ginst689 (P1_R1105_U148, P1_R1105_U256, P1_R1105_U257, P1_R1105_U40, P1_R1105_U41);
  nand ginst690 (P1_R1105_U149, P1_R1105_U40, P1_R1105_U41);
  and ginst691 (P1_R1105_U15, P1_R1105_U140, P1_R1105_U143);
  nand ginst692 (P1_R1105_U150, P1_REG2_REG_2__SCAN_IN, P1_U3457);
  nand ginst693 (P1_R1105_U151, P1_R1105_U149, P1_R1105_U150, P1_R1105_U97);
  or ginst694 (P1_R1105_U152, P1_REG2_REG_1__SCAN_IN, P1_U3454);
  not ginst695 (P1_R1105_U153, P1_R1105_U83);
  or ginst696 (P1_R1105_U154, P1_REG2_REG_9__SCAN_IN, P1_U3478);
  or ginst697 (P1_R1105_U155, P1_REG2_REG_10__SCAN_IN, P1_U3481);
  nand ginst698 (P1_R1105_U156, P1_R1105_U7, P1_R1105_U93);
  nand ginst699 (P1_R1105_U157, P1_REG2_REG_10__SCAN_IN, P1_U3481);
  nand ginst700 (P1_R1105_U158, P1_R1105_U156, P1_R1105_U157, P1_R1105_U90);
  or ginst701 (P1_R1105_U159, P1_REG2_REG_10__SCAN_IN, P1_U3481);
  and ginst702 (P1_R1105_U16, P1_R1105_U126, P1_R1105_U129);
  nand ginst703 (P1_R1105_U160, P1_R1105_U120, P1_R1105_U7, P1_R1105_U81);
  nand ginst704 (P1_R1105_U161, P1_R1105_U158, P1_R1105_U159);
  not ginst705 (P1_R1105_U162, P1_R1105_U88);
  or ginst706 (P1_R1105_U163, P1_REG2_REG_13__SCAN_IN, P1_U3490);
  or ginst707 (P1_R1105_U164, P1_REG2_REG_12__SCAN_IN, P1_U3487);
  nand ginst708 (P1_R1105_U165, P1_R1105_U8, P1_R1105_U92);
  nand ginst709 (P1_R1105_U166, P1_REG2_REG_13__SCAN_IN, P1_U3490);
  nand ginst710 (P1_R1105_U167, P1_R1105_U165, P1_R1105_U166, P1_R1105_U91);
  or ginst711 (P1_R1105_U168, P1_REG2_REG_11__SCAN_IN, P1_U3484);
  or ginst712 (P1_R1105_U169, P1_REG2_REG_13__SCAN_IN, P1_U3490);
  not ginst713 (P1_R1105_U17, P1_REG2_REG_6__SCAN_IN);
  nand ginst714 (P1_R1105_U170, P1_R1105_U168, P1_R1105_U8, P1_R1105_U88);
  nand ginst715 (P1_R1105_U171, P1_R1105_U167, P1_R1105_U169);
  not ginst716 (P1_R1105_U172, P1_R1105_U87);
  or ginst717 (P1_R1105_U173, P1_REG2_REG_14__SCAN_IN, P1_U3493);
  nand ginst718 (P1_R1105_U174, P1_R1105_U173, P1_R1105_U87);
  nand ginst719 (P1_R1105_U175, P1_REG2_REG_14__SCAN_IN, P1_U3493);
  not ginst720 (P1_R1105_U176, P1_R1105_U86);
  or ginst721 (P1_R1105_U177, P1_REG2_REG_15__SCAN_IN, P1_U3496);
  nand ginst722 (P1_R1105_U178, P1_R1105_U177, P1_R1105_U86);
  nand ginst723 (P1_R1105_U179, P1_REG2_REG_15__SCAN_IN, P1_U3496);
  not ginst724 (P1_R1105_U18, P1_U3469);
  not ginst725 (P1_R1105_U180, P1_R1105_U66);
  or ginst726 (P1_R1105_U181, P1_REG2_REG_17__SCAN_IN, P1_U3502);
  or ginst727 (P1_R1105_U182, P1_REG2_REG_16__SCAN_IN, P1_U3499);
  not ginst728 (P1_R1105_U183, P1_R1105_U47);
  nand ginst729 (P1_R1105_U184, P1_R1105_U47, P1_R1105_U48);
  nand ginst730 (P1_R1105_U185, P1_R1105_U184, P1_U3502);
  nand ginst731 (P1_R1105_U186, P1_REG2_REG_17__SCAN_IN, P1_R1105_U183);
  nand ginst732 (P1_R1105_U187, P1_R1105_U66, P1_R1105_U9);
  not ginst733 (P1_R1105_U188, P1_R1105_U65);
  or ginst734 (P1_R1105_U189, P1_REG2_REG_18__SCAN_IN, P1_U3505);
  not ginst735 (P1_R1105_U19, P1_U3472);
  nand ginst736 (P1_R1105_U190, P1_R1105_U189, P1_R1105_U65);
  nand ginst737 (P1_R1105_U191, P1_REG2_REG_18__SCAN_IN, P1_U3505);
  nand ginst738 (P1_R1105_U192, P1_R1105_U190, P1_R1105_U191, P1_R1105_U260, P1_R1105_U261);
  nand ginst739 (P1_R1105_U193, P1_REG2_REG_18__SCAN_IN, P1_U3505);
  nand ginst740 (P1_R1105_U194, P1_R1105_U188, P1_R1105_U193);
  or ginst741 (P1_R1105_U195, P1_REG2_REG_18__SCAN_IN, P1_U3505);
  nand ginst742 (P1_R1105_U196, P1_R1105_U194, P1_R1105_U195, P1_R1105_U264);
  or ginst743 (P1_R1105_U197, P1_REG2_REG_16__SCAN_IN, P1_U3499);
  nand ginst744 (P1_R1105_U198, P1_R1105_U197, P1_R1105_U66);
  nand ginst745 (P1_R1105_U199, P1_R1105_U198, P1_R1105_U272, P1_R1105_U273, P1_R1105_U47);
  nand ginst746 (P1_R1105_U20, P1_REG2_REG_6__SCAN_IN, P1_U3469);
  nand ginst747 (P1_R1105_U200, P1_R1105_U180, P1_R1105_U47);
  nand ginst748 (P1_R1105_U201, P1_REG2_REG_17__SCAN_IN, P1_U3502);
  nand ginst749 (P1_R1105_U202, P1_R1105_U200, P1_R1105_U201, P1_R1105_U9);
  or ginst750 (P1_R1105_U203, P1_REG2_REG_16__SCAN_IN, P1_U3499);
  nand ginst751 (P1_R1105_U204, P1_R1105_U168, P1_R1105_U88);
  not ginst752 (P1_R1105_U205, P1_R1105_U67);
  or ginst753 (P1_R1105_U206, P1_REG2_REG_12__SCAN_IN, P1_U3487);
  nand ginst754 (P1_R1105_U207, P1_R1105_U206, P1_R1105_U67);
  nand ginst755 (P1_R1105_U208, P1_R1105_U207, P1_R1105_U293, P1_R1105_U294, P1_R1105_U91);
  nand ginst756 (P1_R1105_U209, P1_R1105_U205, P1_R1105_U91);
  not ginst757 (P1_R1105_U21, P1_REG2_REG_7__SCAN_IN);
  nand ginst758 (P1_R1105_U210, P1_REG2_REG_13__SCAN_IN, P1_U3490);
  nand ginst759 (P1_R1105_U211, P1_R1105_U209, P1_R1105_U210, P1_R1105_U8);
  or ginst760 (P1_R1105_U212, P1_REG2_REG_12__SCAN_IN, P1_U3487);
  or ginst761 (P1_R1105_U213, P1_REG2_REG_9__SCAN_IN, P1_U3478);
  nand ginst762 (P1_R1105_U214, P1_R1105_U213, P1_R1105_U38);
  nand ginst763 (P1_R1105_U215, P1_R1105_U214, P1_R1105_U305, P1_R1105_U306, P1_R1105_U90);
  nand ginst764 (P1_R1105_U216, P1_R1105_U122, P1_R1105_U90);
  nand ginst765 (P1_R1105_U217, P1_REG2_REG_10__SCAN_IN, P1_U3481);
  nand ginst766 (P1_R1105_U218, P1_R1105_U216, P1_R1105_U217, P1_R1105_U7);
  nand ginst767 (P1_R1105_U219, P1_R1105_U123, P1_R1105_U90);
  not ginst768 (P1_R1105_U22, P1_REG2_REG_4__SCAN_IN);
  nand ginst769 (P1_R1105_U220, P1_R1105_U120, P1_R1105_U49);
  nand ginst770 (P1_R1105_U221, P1_R1105_U130, P1_R1105_U20);
  nand ginst771 (P1_R1105_U222, P1_R1105_U144, P1_R1105_U32);
  nand ginst772 (P1_R1105_U223, P1_R1105_U147, P1_R1105_U96);
  nand ginst773 (P1_R1105_U224, P1_R1105_U203, P1_R1105_U47);
  nand ginst774 (P1_R1105_U225, P1_R1105_U212, P1_R1105_U91);
  nand ginst775 (P1_R1105_U226, P1_R1105_U168, P1_R1105_U56);
  nand ginst776 (P1_R1105_U227, P1_R1105_U37, P1_U3478);
  nand ginst777 (P1_R1105_U228, P1_REG2_REG_9__SCAN_IN, P1_R1105_U36);
  nand ginst778 (P1_R1105_U229, P1_R1105_U227, P1_R1105_U228);
  not ginst779 (P1_R1105_U23, P1_U3463);
  nand ginst780 (P1_R1105_U230, P1_R1105_U219, P1_R1105_U38);
  nand ginst781 (P1_R1105_U231, P1_R1105_U122, P1_R1105_U229);
  nand ginst782 (P1_R1105_U232, P1_R1105_U34, P1_U3475);
  nand ginst783 (P1_R1105_U233, P1_REG2_REG_8__SCAN_IN, P1_R1105_U35);
  nand ginst784 (P1_R1105_U234, P1_R1105_U232, P1_R1105_U233);
  nand ginst785 (P1_R1105_U235, P1_R1105_U220, P1_R1105_U81);
  nand ginst786 (P1_R1105_U236, P1_R1105_U119, P1_R1105_U234);
  nand ginst787 (P1_R1105_U237, P1_R1105_U21, P1_U3472);
  nand ginst788 (P1_R1105_U238, P1_REG2_REG_7__SCAN_IN, P1_R1105_U19);
  nand ginst789 (P1_R1105_U239, P1_R1105_U17, P1_U3469);
  not ginst790 (P1_R1105_U24, P1_U3466);
  nand ginst791 (P1_R1105_U240, P1_REG2_REG_6__SCAN_IN, P1_R1105_U18);
  nand ginst792 (P1_R1105_U241, P1_R1105_U239, P1_R1105_U240);
  nand ginst793 (P1_R1105_U242, P1_R1105_U221, P1_R1105_U39);
  nand ginst794 (P1_R1105_U243, P1_R1105_U111, P1_R1105_U241);
  nand ginst795 (P1_R1105_U244, P1_R1105_U33, P1_U3466);
  nand ginst796 (P1_R1105_U245, P1_REG2_REG_5__SCAN_IN, P1_R1105_U24);
  nand ginst797 (P1_R1105_U246, P1_R1105_U22, P1_U3463);
  nand ginst798 (P1_R1105_U247, P1_REG2_REG_4__SCAN_IN, P1_R1105_U23);
  nand ginst799 (P1_R1105_U248, P1_R1105_U246, P1_R1105_U247);
  nand ginst800 (P1_R1105_U249, P1_R1105_U222, P1_R1105_U42);
  not ginst801 (P1_R1105_U25, P1_REG2_REG_2__SCAN_IN);
  nand ginst802 (P1_R1105_U250, P1_R1105_U137, P1_R1105_U248);
  nand ginst803 (P1_R1105_U251, P1_R1105_U30, P1_U3460);
  nand ginst804 (P1_R1105_U252, P1_REG2_REG_3__SCAN_IN, P1_R1105_U31);
  nand ginst805 (P1_R1105_U253, P1_R1105_U251, P1_R1105_U252);
  nand ginst806 (P1_R1105_U254, P1_R1105_U223, P1_R1105_U82);
  nand ginst807 (P1_R1105_U255, P1_R1105_U146, P1_R1105_U253);
  nand ginst808 (P1_R1105_U256, P1_R1105_U25, P1_U3457);
  nand ginst809 (P1_R1105_U257, P1_REG2_REG_2__SCAN_IN, P1_R1105_U26);
  nand ginst810 (P1_R1105_U258, P1_R1105_U83, P1_R1105_U98);
  nand ginst811 (P1_R1105_U259, P1_R1105_U153, P1_R1105_U29);
  not ginst812 (P1_R1105_U26, P1_U3457);
  nand ginst813 (P1_R1105_U260, P1_R1105_U85, P1_U3442);
  nand ginst814 (P1_R1105_U261, P1_REG2_REG_19__SCAN_IN, P1_R1105_U84);
  nand ginst815 (P1_R1105_U262, P1_R1105_U85, P1_U3442);
  nand ginst816 (P1_R1105_U263, P1_REG2_REG_19__SCAN_IN, P1_R1105_U84);
  nand ginst817 (P1_R1105_U264, P1_R1105_U262, P1_R1105_U263);
  nand ginst818 (P1_R1105_U265, P1_R1105_U63, P1_U3505);
  nand ginst819 (P1_R1105_U266, P1_REG2_REG_18__SCAN_IN, P1_R1105_U64);
  nand ginst820 (P1_R1105_U267, P1_R1105_U63, P1_U3505);
  nand ginst821 (P1_R1105_U268, P1_REG2_REG_18__SCAN_IN, P1_R1105_U64);
  nand ginst822 (P1_R1105_U269, P1_R1105_U267, P1_R1105_U268);
  not ginst823 (P1_R1105_U27, P1_REG2_REG_0__SCAN_IN);
  nand ginst824 (P1_R1105_U270, P1_R1105_U265, P1_R1105_U266, P1_R1105_U65);
  nand ginst825 (P1_R1105_U271, P1_R1105_U188, P1_R1105_U269);
  nand ginst826 (P1_R1105_U272, P1_R1105_U48, P1_U3502);
  nand ginst827 (P1_R1105_U273, P1_REG2_REG_17__SCAN_IN, P1_R1105_U46);
  nand ginst828 (P1_R1105_U274, P1_R1105_U44, P1_U3499);
  nand ginst829 (P1_R1105_U275, P1_REG2_REG_16__SCAN_IN, P1_R1105_U45);
  nand ginst830 (P1_R1105_U276, P1_R1105_U274, P1_R1105_U275);
  nand ginst831 (P1_R1105_U277, P1_R1105_U224, P1_R1105_U66);
  nand ginst832 (P1_R1105_U278, P1_R1105_U180, P1_R1105_U276);
  nand ginst833 (P1_R1105_U279, P1_R1105_U61, P1_U3496);
  not ginst834 (P1_R1105_U28, P1_U3448);
  nand ginst835 (P1_R1105_U280, P1_REG2_REG_15__SCAN_IN, P1_R1105_U62);
  nand ginst836 (P1_R1105_U281, P1_R1105_U61, P1_U3496);
  nand ginst837 (P1_R1105_U282, P1_REG2_REG_15__SCAN_IN, P1_R1105_U62);
  nand ginst838 (P1_R1105_U283, P1_R1105_U281, P1_R1105_U282);
  nand ginst839 (P1_R1105_U284, P1_R1105_U279, P1_R1105_U280, P1_R1105_U86);
  nand ginst840 (P1_R1105_U285, P1_R1105_U176, P1_R1105_U283);
  nand ginst841 (P1_R1105_U286, P1_R1105_U59, P1_U3493);
  nand ginst842 (P1_R1105_U287, P1_REG2_REG_14__SCAN_IN, P1_R1105_U60);
  nand ginst843 (P1_R1105_U288, P1_R1105_U59, P1_U3493);
  nand ginst844 (P1_R1105_U289, P1_REG2_REG_14__SCAN_IN, P1_R1105_U60);
  nand ginst845 (P1_R1105_U29, P1_REG2_REG_0__SCAN_IN, P1_U3448);
  nand ginst846 (P1_R1105_U290, P1_R1105_U288, P1_R1105_U289);
  nand ginst847 (P1_R1105_U291, P1_R1105_U286, P1_R1105_U287, P1_R1105_U87);
  nand ginst848 (P1_R1105_U292, P1_R1105_U172, P1_R1105_U290);
  nand ginst849 (P1_R1105_U293, P1_R1105_U57, P1_U3490);
  nand ginst850 (P1_R1105_U294, P1_REG2_REG_13__SCAN_IN, P1_R1105_U58);
  nand ginst851 (P1_R1105_U295, P1_R1105_U52, P1_U3487);
  nand ginst852 (P1_R1105_U296, P1_REG2_REG_12__SCAN_IN, P1_R1105_U53);
  nand ginst853 (P1_R1105_U297, P1_R1105_U295, P1_R1105_U296);
  nand ginst854 (P1_R1105_U298, P1_R1105_U225, P1_R1105_U67);
  nand ginst855 (P1_R1105_U299, P1_R1105_U205, P1_R1105_U297);
  not ginst856 (P1_R1105_U30, P1_REG2_REG_3__SCAN_IN);
  nand ginst857 (P1_R1105_U300, P1_R1105_U54, P1_U3484);
  nand ginst858 (P1_R1105_U301, P1_REG2_REG_11__SCAN_IN, P1_R1105_U55);
  nand ginst859 (P1_R1105_U302, P1_R1105_U300, P1_R1105_U301);
  nand ginst860 (P1_R1105_U303, P1_R1105_U226, P1_R1105_U88);
  nand ginst861 (P1_R1105_U304, P1_R1105_U162, P1_R1105_U302);
  nand ginst862 (P1_R1105_U305, P1_R1105_U50, P1_U3481);
  nand ginst863 (P1_R1105_U306, P1_REG2_REG_10__SCAN_IN, P1_R1105_U51);
  nand ginst864 (P1_R1105_U307, P1_R1105_U27, P1_U3448);
  nand ginst865 (P1_R1105_U308, P1_REG2_REG_0__SCAN_IN, P1_R1105_U28);
  not ginst866 (P1_R1105_U31, P1_U3460);
  nand ginst867 (P1_R1105_U32, P1_REG2_REG_4__SCAN_IN, P1_U3463);
  not ginst868 (P1_R1105_U33, P1_REG2_REG_5__SCAN_IN);
  not ginst869 (P1_R1105_U34, P1_REG2_REG_8__SCAN_IN);
  not ginst870 (P1_R1105_U35, P1_U3475);
  not ginst871 (P1_R1105_U36, P1_U3478);
  not ginst872 (P1_R1105_U37, P1_REG2_REG_9__SCAN_IN);
  nand ginst873 (P1_R1105_U38, P1_R1105_U121, P1_R1105_U49);
  nand ginst874 (P1_R1105_U39, P1_R1105_U108, P1_R1105_U109, P1_R1105_U110);
  and ginst875 (P1_R1105_U4, P1_R1105_U94, P1_R1105_U95);
  nand ginst876 (P1_R1105_U40, P1_R1105_U98, P1_R1105_U99);
  nand ginst877 (P1_R1105_U41, P1_REG2_REG_1__SCAN_IN, P1_U3454);
  nand ginst878 (P1_R1105_U42, P1_R1105_U134, P1_R1105_U135, P1_R1105_U136);
  nand ginst879 (P1_R1105_U43, P1_R1105_U131, P1_R1105_U132);
  not ginst880 (P1_R1105_U44, P1_REG2_REG_16__SCAN_IN);
  not ginst881 (P1_R1105_U45, P1_U3499);
  not ginst882 (P1_R1105_U46, P1_U3502);
  nand ginst883 (P1_R1105_U47, P1_REG2_REG_16__SCAN_IN, P1_U3499);
  not ginst884 (P1_R1105_U48, P1_REG2_REG_17__SCAN_IN);
  nand ginst885 (P1_R1105_U49, P1_REG2_REG_8__SCAN_IN, P1_U3475);
  and ginst886 (P1_R1105_U5, P1_R1105_U96, P1_R1105_U97);
  not ginst887 (P1_R1105_U50, P1_REG2_REG_10__SCAN_IN);
  not ginst888 (P1_R1105_U51, P1_U3481);
  not ginst889 (P1_R1105_U52, P1_REG2_REG_12__SCAN_IN);
  not ginst890 (P1_R1105_U53, P1_U3487);
  not ginst891 (P1_R1105_U54, P1_REG2_REG_11__SCAN_IN);
  not ginst892 (P1_R1105_U55, P1_U3484);
  nand ginst893 (P1_R1105_U56, P1_REG2_REG_11__SCAN_IN, P1_U3484);
  not ginst894 (P1_R1105_U57, P1_REG2_REG_13__SCAN_IN);
  not ginst895 (P1_R1105_U58, P1_U3490);
  not ginst896 (P1_R1105_U59, P1_REG2_REG_14__SCAN_IN);
  and ginst897 (P1_R1105_U6, P1_R1105_U112, P1_R1105_U113);
  not ginst898 (P1_R1105_U60, P1_U3493);
  not ginst899 (P1_R1105_U61, P1_REG2_REG_15__SCAN_IN);
  not ginst900 (P1_R1105_U62, P1_U3496);
  not ginst901 (P1_R1105_U63, P1_REG2_REG_18__SCAN_IN);
  not ginst902 (P1_R1105_U64, P1_U3505);
  nand ginst903 (P1_R1105_U65, P1_R1105_U185, P1_R1105_U186, P1_R1105_U187);
  nand ginst904 (P1_R1105_U66, P1_R1105_U178, P1_R1105_U179);
  nand ginst905 (P1_R1105_U67, P1_R1105_U204, P1_R1105_U56);
  nand ginst906 (P1_R1105_U68, P1_R1105_U258, P1_R1105_U259);
  nand ginst907 (P1_R1105_U69, P1_R1105_U307, P1_R1105_U308);
  and ginst908 (P1_R1105_U7, P1_R1105_U154, P1_R1105_U155);
  nand ginst909 (P1_R1105_U70, P1_R1105_U230, P1_R1105_U231);
  nand ginst910 (P1_R1105_U71, P1_R1105_U235, P1_R1105_U236);
  nand ginst911 (P1_R1105_U72, P1_R1105_U242, P1_R1105_U243);
  nand ginst912 (P1_R1105_U73, P1_R1105_U249, P1_R1105_U250);
  nand ginst913 (P1_R1105_U74, P1_R1105_U254, P1_R1105_U255);
  nand ginst914 (P1_R1105_U75, P1_R1105_U270, P1_R1105_U271);
  nand ginst915 (P1_R1105_U76, P1_R1105_U277, P1_R1105_U278);
  nand ginst916 (P1_R1105_U77, P1_R1105_U284, P1_R1105_U285);
  nand ginst917 (P1_R1105_U78, P1_R1105_U291, P1_R1105_U292);
  nand ginst918 (P1_R1105_U79, P1_R1105_U298, P1_R1105_U299);
  and ginst919 (P1_R1105_U8, P1_R1105_U163, P1_R1105_U164);
  nand ginst920 (P1_R1105_U80, P1_R1105_U303, P1_R1105_U304);
  nand ginst921 (P1_R1105_U81, P1_R1105_U116, P1_R1105_U117, P1_R1105_U118);
  nand ginst922 (P1_R1105_U82, P1_R1105_U133, P1_R1105_U145);
  nand ginst923 (P1_R1105_U83, P1_R1105_U152, P1_R1105_U41);
  not ginst924 (P1_R1105_U84, P1_U3442);
  not ginst925 (P1_R1105_U85, P1_REG2_REG_19__SCAN_IN);
  nand ginst926 (P1_R1105_U86, P1_R1105_U174, P1_R1105_U175);
  nand ginst927 (P1_R1105_U87, P1_R1105_U170, P1_R1105_U171);
  nand ginst928 (P1_R1105_U88, P1_R1105_U160, P1_R1105_U161);
  not ginst929 (P1_R1105_U89, P1_R1105_U32);
  and ginst930 (P1_R1105_U9, P1_R1105_U181, P1_R1105_U182);
  nand ginst931 (P1_R1105_U90, P1_REG2_REG_9__SCAN_IN, P1_U3478);
  nand ginst932 (P1_R1105_U91, P1_REG2_REG_12__SCAN_IN, P1_U3487);
  not ginst933 (P1_R1105_U92, P1_R1105_U56);
  not ginst934 (P1_R1105_U93, P1_R1105_U49);
  or ginst935 (P1_R1105_U94, P1_REG2_REG_5__SCAN_IN, P1_U3466);
  or ginst936 (P1_R1105_U95, P1_REG2_REG_4__SCAN_IN, P1_U3463);
  or ginst937 (P1_R1105_U96, P1_REG2_REG_3__SCAN_IN, P1_U3460);
  or ginst938 (P1_R1105_U97, P1_REG2_REG_2__SCAN_IN, P1_U3457);
  not ginst939 (P1_R1105_U98, P1_R1105_U29);
  or ginst940 (P1_R1105_U99, P1_REG2_REG_1__SCAN_IN, P1_U3454);
  nand ginst941 (P1_R1117_U10, P1_R1117_U340, P1_R1117_U343);
  nand ginst942 (P1_R1117_U100, P1_R1117_U460, P1_R1117_U461);
  nand ginst943 (P1_R1117_U101, P1_R1117_U465, P1_R1117_U466);
  nand ginst944 (P1_R1117_U102, P1_R1117_U350, P1_R1117_U351);
  nand ginst945 (P1_R1117_U103, P1_R1117_U359, P1_R1117_U360);
  nand ginst946 (P1_R1117_U104, P1_R1117_U366, P1_R1117_U367);
  nand ginst947 (P1_R1117_U105, P1_R1117_U370, P1_R1117_U371);
  nand ginst948 (P1_R1117_U106, P1_R1117_U379, P1_R1117_U380);
  nand ginst949 (P1_R1117_U107, P1_R1117_U398, P1_R1117_U399);
  nand ginst950 (P1_R1117_U108, P1_R1117_U415, P1_R1117_U416);
  nand ginst951 (P1_R1117_U109, P1_R1117_U419, P1_R1117_U420);
  nand ginst952 (P1_R1117_U11, P1_R1117_U329, P1_R1117_U332);
  nand ginst953 (P1_R1117_U110, P1_R1117_U451, P1_R1117_U452);
  nand ginst954 (P1_R1117_U111, P1_R1117_U455, P1_R1117_U456);
  nand ginst955 (P1_R1117_U112, P1_R1117_U472, P1_R1117_U473);
  and ginst956 (P1_R1117_U113, P1_R1117_U193, P1_R1117_U194);
  and ginst957 (P1_R1117_U114, P1_R1117_U196, P1_R1117_U201);
  and ginst958 (P1_R1117_U115, P1_R1117_U180, P1_R1117_U206);
  and ginst959 (P1_R1117_U116, P1_R1117_U209, P1_R1117_U210);
  and ginst960 (P1_R1117_U117, P1_R1117_U352, P1_R1117_U353, P1_R1117_U37);
  and ginst961 (P1_R1117_U118, P1_R1117_U180, P1_R1117_U356);
  and ginst962 (P1_R1117_U119, P1_R1117_U225, P1_R1117_U6);
  nand ginst963 (P1_R1117_U12, P1_R1117_U318, P1_R1117_U321);
  and ginst964 (P1_R1117_U120, P1_R1117_U179, P1_R1117_U363);
  and ginst965 (P1_R1117_U121, P1_R1117_U27, P1_R1117_U372, P1_R1117_U373);
  and ginst966 (P1_R1117_U122, P1_R1117_U178, P1_R1117_U376);
  and ginst967 (P1_R1117_U123, P1_R1117_U174, P1_R1117_U212, P1_R1117_U235);
  and ginst968 (P1_R1117_U124, P1_R1117_U175, P1_R1117_U252, P1_R1117_U257);
  and ginst969 (P1_R1117_U125, P1_R1117_U176, P1_R1117_U283);
  and ginst970 (P1_R1117_U126, P1_R1117_U299, P1_R1117_U300);
  nand ginst971 (P1_R1117_U127, P1_R1117_U386, P1_R1117_U387);
  and ginst972 (P1_R1117_U128, P1_R1117_U391, P1_R1117_U392, P1_R1117_U82);
  and ginst973 (P1_R1117_U129, P1_R1117_U177, P1_R1117_U395);
  nand ginst974 (P1_R1117_U13, P1_R1117_U310, P1_R1117_U312);
  nand ginst975 (P1_R1117_U130, P1_R1117_U400, P1_R1117_U401);
  nand ginst976 (P1_R1117_U131, P1_R1117_U405, P1_R1117_U406);
  and ginst977 (P1_R1117_U132, P1_R1117_U176, P1_R1117_U412);
  nand ginst978 (P1_R1117_U133, P1_R1117_U421, P1_R1117_U422);
  nand ginst979 (P1_R1117_U134, P1_R1117_U426, P1_R1117_U427);
  nand ginst980 (P1_R1117_U135, P1_R1117_U431, P1_R1117_U432);
  nand ginst981 (P1_R1117_U136, P1_R1117_U436, P1_R1117_U437);
  nand ginst982 (P1_R1117_U137, P1_R1117_U441, P1_R1117_U442);
  and ginst983 (P1_R1117_U138, P1_R1117_U331, P1_R1117_U8);
  and ginst984 (P1_R1117_U139, P1_R1117_U175, P1_R1117_U448);
  nand ginst985 (P1_R1117_U14, P1_R1117_U308, P1_R1117_U347);
  nand ginst986 (P1_R1117_U140, P1_R1117_U457, P1_R1117_U458);
  nand ginst987 (P1_R1117_U141, P1_R1117_U462, P1_R1117_U463);
  and ginst988 (P1_R1117_U142, P1_R1117_U342, P1_R1117_U7);
  and ginst989 (P1_R1117_U143, P1_R1117_U174, P1_R1117_U469);
  and ginst990 (P1_R1117_U144, P1_R1117_U348, P1_R1117_U349);
  nand ginst991 (P1_R1117_U145, P1_R1117_U116, P1_R1117_U207);
  and ginst992 (P1_R1117_U146, P1_R1117_U357, P1_R1117_U358);
  and ginst993 (P1_R1117_U147, P1_R1117_U364, P1_R1117_U365);
  and ginst994 (P1_R1117_U148, P1_R1117_U368, P1_R1117_U369);
  nand ginst995 (P1_R1117_U149, P1_R1117_U113, P1_R1117_U191);
  nand ginst996 (P1_R1117_U15, P1_R1117_U231, P1_R1117_U233);
  and ginst997 (P1_R1117_U150, P1_R1117_U377, P1_R1117_U378);
  not ginst998 (P1_R1117_U151, P1_U3985);
  not ginst999 (P1_R1117_U152, P1_U3055);
  and ginst1000 (P1_R1117_U153, P1_R1117_U381, P1_R1117_U382);
  and ginst1001 (P1_R1117_U154, P1_R1117_U396, P1_R1117_U397);
  nand ginst1002 (P1_R1117_U155, P1_R1117_U289, P1_R1117_U290);
  nand ginst1003 (P1_R1117_U156, P1_R1117_U285, P1_R1117_U286);
  and ginst1004 (P1_R1117_U157, P1_R1117_U413, P1_R1117_U414);
  and ginst1005 (P1_R1117_U158, P1_R1117_U417, P1_R1117_U418);
  nand ginst1006 (P1_R1117_U159, P1_R1117_U275, P1_R1117_U276);
  nand ginst1007 (P1_R1117_U16, P1_R1117_U223, P1_R1117_U226);
  nand ginst1008 (P1_R1117_U160, P1_R1117_U271, P1_R1117_U272);
  not ginst1009 (P1_R1117_U161, P1_U3455);
  nand ginst1010 (P1_R1117_U162, P1_R1117_U267, P1_R1117_U268);
  not ginst1011 (P1_R1117_U163, P1_U3506);
  nand ginst1012 (P1_R1117_U164, P1_R1117_U259, P1_R1117_U260);
  and ginst1013 (P1_R1117_U165, P1_R1117_U449, P1_R1117_U450);
  and ginst1014 (P1_R1117_U166, P1_R1117_U453, P1_R1117_U454);
  nand ginst1015 (P1_R1117_U167, P1_R1117_U249, P1_R1117_U250);
  nand ginst1016 (P1_R1117_U168, P1_R1117_U245, P1_R1117_U246);
  nand ginst1017 (P1_R1117_U169, P1_R1117_U241, P1_R1117_U242);
  nand ginst1018 (P1_R1117_U17, P1_R1117_U215, P1_R1117_U217);
  and ginst1019 (P1_R1117_U170, P1_R1117_U470, P1_R1117_U471);
  not ginst1020 (P1_R1117_U171, P1_R1117_U82);
  not ginst1021 (P1_R1117_U172, P1_R1117_U27);
  not ginst1022 (P1_R1117_U173, P1_R1117_U37);
  nand ginst1023 (P1_R1117_U174, P1_R1117_U50, P1_U3482);
  nand ginst1024 (P1_R1117_U175, P1_R1117_U59, P1_U3497);
  nand ginst1025 (P1_R1117_U176, P1_R1117_U73, P1_U3980);
  nand ginst1026 (P1_R1117_U177, P1_R1117_U81, P1_U3976);
  nand ginst1027 (P1_R1117_U178, P1_R1117_U26, P1_U3458);
  nand ginst1028 (P1_R1117_U179, P1_R1117_U32, P1_U3467);
  nand ginst1029 (P1_R1117_U18, P1_R1117_U23, P1_R1117_U346);
  nand ginst1030 (P1_R1117_U180, P1_R1117_U36, P1_U3473);
  not ginst1031 (P1_R1117_U181, P1_R1117_U61);
  not ginst1032 (P1_R1117_U182, P1_R1117_U75);
  not ginst1033 (P1_R1117_U183, P1_R1117_U34);
  not ginst1034 (P1_R1117_U184, P1_R1117_U51);
  not ginst1035 (P1_R1117_U185, P1_R1117_U23);
  nand ginst1036 (P1_R1117_U186, P1_R1117_U185, P1_R1117_U24);
  nand ginst1037 (P1_R1117_U187, P1_R1117_U161, P1_R1117_U186);
  nand ginst1038 (P1_R1117_U188, P1_R1117_U23, P1_U3078);
  not ginst1039 (P1_R1117_U189, P1_R1117_U43);
  not ginst1040 (P1_R1117_U19, P1_U3473);
  nand ginst1041 (P1_R1117_U190, P1_R1117_U28, P1_U3461);
  nand ginst1042 (P1_R1117_U191, P1_R1117_U178, P1_R1117_U190, P1_R1117_U43);
  nand ginst1043 (P1_R1117_U192, P1_R1117_U27, P1_R1117_U28);
  nand ginst1044 (P1_R1117_U193, P1_R1117_U192, P1_R1117_U25);
  nand ginst1045 (P1_R1117_U194, P1_R1117_U172, P1_U3064);
  not ginst1046 (P1_R1117_U195, P1_R1117_U149);
  nand ginst1047 (P1_R1117_U196, P1_R1117_U31, P1_U3470);
  nand ginst1048 (P1_R1117_U197, P1_R1117_U29, P1_U3071);
  nand ginst1049 (P1_R1117_U198, P1_R1117_U20, P1_U3067);
  nand ginst1050 (P1_R1117_U199, P1_R1117_U179, P1_R1117_U183);
  not ginst1051 (P1_R1117_U20, P1_U3467);
  nand ginst1052 (P1_R1117_U200, P1_R1117_U199, P1_R1117_U6);
  nand ginst1053 (P1_R1117_U201, P1_R1117_U33, P1_U3464);
  nand ginst1054 (P1_R1117_U202, P1_R1117_U31, P1_U3470);
  nand ginst1055 (P1_R1117_U203, P1_R1117_U114, P1_R1117_U149, P1_R1117_U179);
  nand ginst1056 (P1_R1117_U204, P1_R1117_U200, P1_R1117_U202);
  not ginst1057 (P1_R1117_U205, P1_R1117_U41);
  nand ginst1058 (P1_R1117_U206, P1_R1117_U38, P1_U3476);
  nand ginst1059 (P1_R1117_U207, P1_R1117_U115, P1_R1117_U41);
  nand ginst1060 (P1_R1117_U208, P1_R1117_U37, P1_R1117_U38);
  nand ginst1061 (P1_R1117_U209, P1_R1117_U208, P1_R1117_U35);
  not ginst1062 (P1_R1117_U21, P1_U3458);
  nand ginst1063 (P1_R1117_U210, P1_R1117_U173, P1_U3084);
  not ginst1064 (P1_R1117_U211, P1_R1117_U145);
  nand ginst1065 (P1_R1117_U212, P1_R1117_U40, P1_U3479);
  nand ginst1066 (P1_R1117_U213, P1_R1117_U212, P1_R1117_U51);
  nand ginst1067 (P1_R1117_U214, P1_R1117_U205, P1_R1117_U37);
  nand ginst1068 (P1_R1117_U215, P1_R1117_U118, P1_R1117_U214);
  nand ginst1069 (P1_R1117_U216, P1_R1117_U180, P1_R1117_U41);
  nand ginst1070 (P1_R1117_U217, P1_R1117_U117, P1_R1117_U216);
  nand ginst1071 (P1_R1117_U218, P1_R1117_U180, P1_R1117_U37);
  nand ginst1072 (P1_R1117_U219, P1_R1117_U149, P1_R1117_U201);
  not ginst1073 (P1_R1117_U22, P1_U3450);
  not ginst1074 (P1_R1117_U220, P1_R1117_U42);
  nand ginst1075 (P1_R1117_U221, P1_R1117_U20, P1_U3067);
  nand ginst1076 (P1_R1117_U222, P1_R1117_U220, P1_R1117_U221);
  nand ginst1077 (P1_R1117_U223, P1_R1117_U120, P1_R1117_U222);
  nand ginst1078 (P1_R1117_U224, P1_R1117_U179, P1_R1117_U42);
  nand ginst1079 (P1_R1117_U225, P1_R1117_U31, P1_U3470);
  nand ginst1080 (P1_R1117_U226, P1_R1117_U119, P1_R1117_U224);
  nand ginst1081 (P1_R1117_U227, P1_R1117_U20, P1_U3067);
  nand ginst1082 (P1_R1117_U228, P1_R1117_U179, P1_R1117_U227);
  nand ginst1083 (P1_R1117_U229, P1_R1117_U201, P1_R1117_U34);
  nand ginst1084 (P1_R1117_U23, P1_R1117_U91, P1_U3450);
  nand ginst1085 (P1_R1117_U230, P1_R1117_U189, P1_R1117_U27);
  nand ginst1086 (P1_R1117_U231, P1_R1117_U122, P1_R1117_U230);
  nand ginst1087 (P1_R1117_U232, P1_R1117_U178, P1_R1117_U43);
  nand ginst1088 (P1_R1117_U233, P1_R1117_U121, P1_R1117_U232);
  nand ginst1089 (P1_R1117_U234, P1_R1117_U178, P1_R1117_U27);
  nand ginst1090 (P1_R1117_U235, P1_R1117_U49, P1_U3485);
  nand ginst1091 (P1_R1117_U236, P1_R1117_U48, P1_U3063);
  nand ginst1092 (P1_R1117_U237, P1_R1117_U47, P1_U3062);
  nand ginst1093 (P1_R1117_U238, P1_R1117_U174, P1_R1117_U184);
  nand ginst1094 (P1_R1117_U239, P1_R1117_U238, P1_R1117_U7);
  not ginst1095 (P1_R1117_U24, P1_U3078);
  nand ginst1096 (P1_R1117_U240, P1_R1117_U49, P1_U3485);
  nand ginst1097 (P1_R1117_U241, P1_R1117_U123, P1_R1117_U145);
  nand ginst1098 (P1_R1117_U242, P1_R1117_U239, P1_R1117_U240);
  not ginst1099 (P1_R1117_U243, P1_R1117_U169);
  nand ginst1100 (P1_R1117_U244, P1_R1117_U53, P1_U3488);
  nand ginst1101 (P1_R1117_U245, P1_R1117_U169, P1_R1117_U244);
  nand ginst1102 (P1_R1117_U246, P1_R1117_U52, P1_U3072);
  not ginst1103 (P1_R1117_U247, P1_R1117_U168);
  nand ginst1104 (P1_R1117_U248, P1_R1117_U55, P1_U3491);
  nand ginst1105 (P1_R1117_U249, P1_R1117_U168, P1_R1117_U248);
  not ginst1106 (P1_R1117_U25, P1_U3461);
  nand ginst1107 (P1_R1117_U250, P1_R1117_U54, P1_U3080);
  not ginst1108 (P1_R1117_U251, P1_R1117_U167);
  nand ginst1109 (P1_R1117_U252, P1_R1117_U58, P1_U3500);
  nand ginst1110 (P1_R1117_U253, P1_R1117_U56, P1_U3073);
  nand ginst1111 (P1_R1117_U254, P1_R1117_U46, P1_U3074);
  nand ginst1112 (P1_R1117_U255, P1_R1117_U175, P1_R1117_U181);
  nand ginst1113 (P1_R1117_U256, P1_R1117_U255, P1_R1117_U8);
  nand ginst1114 (P1_R1117_U257, P1_R1117_U60, P1_U3494);
  nand ginst1115 (P1_R1117_U258, P1_R1117_U58, P1_U3500);
  nand ginst1116 (P1_R1117_U259, P1_R1117_U124, P1_R1117_U167);
  not ginst1117 (P1_R1117_U26, P1_U3068);
  nand ginst1118 (P1_R1117_U260, P1_R1117_U256, P1_R1117_U258);
  not ginst1119 (P1_R1117_U261, P1_R1117_U164);
  nand ginst1120 (P1_R1117_U262, P1_R1117_U63, P1_U3503);
  nand ginst1121 (P1_R1117_U263, P1_R1117_U164, P1_R1117_U262);
  nand ginst1122 (P1_R1117_U264, P1_R1117_U62, P1_U3069);
  not ginst1123 (P1_R1117_U265, P1_R1117_U64);
  nand ginst1124 (P1_R1117_U266, P1_R1117_U265, P1_R1117_U65);
  nand ginst1125 (P1_R1117_U267, P1_R1117_U163, P1_R1117_U266);
  nand ginst1126 (P1_R1117_U268, P1_R1117_U64, P1_U3082);
  not ginst1127 (P1_R1117_U269, P1_R1117_U162);
  nand ginst1128 (P1_R1117_U27, P1_R1117_U21, P1_U3068);
  nand ginst1129 (P1_R1117_U270, P1_R1117_U67, P1_U3508);
  nand ginst1130 (P1_R1117_U271, P1_R1117_U162, P1_R1117_U270);
  nand ginst1131 (P1_R1117_U272, P1_R1117_U66, P1_U3081);
  not ginst1132 (P1_R1117_U273, P1_R1117_U160);
  nand ginst1133 (P1_R1117_U274, P1_R1117_U69, P1_U3982);
  nand ginst1134 (P1_R1117_U275, P1_R1117_U160, P1_R1117_U274);
  nand ginst1135 (P1_R1117_U276, P1_R1117_U68, P1_U3076);
  not ginst1136 (P1_R1117_U277, P1_R1117_U159);
  nand ginst1137 (P1_R1117_U278, P1_R1117_U72, P1_U3979);
  nand ginst1138 (P1_R1117_U279, P1_R1117_U70, P1_U3066);
  not ginst1139 (P1_R1117_U28, P1_U3064);
  nand ginst1140 (P1_R1117_U280, P1_R1117_U45, P1_U3061);
  nand ginst1141 (P1_R1117_U281, P1_R1117_U176, P1_R1117_U182);
  nand ginst1142 (P1_R1117_U282, P1_R1117_U281, P1_R1117_U9);
  nand ginst1143 (P1_R1117_U283, P1_R1117_U74, P1_U3981);
  nand ginst1144 (P1_R1117_U284, P1_R1117_U72, P1_U3979);
  nand ginst1145 (P1_R1117_U285, P1_R1117_U125, P1_R1117_U159, P1_R1117_U278);
  nand ginst1146 (P1_R1117_U286, P1_R1117_U282, P1_R1117_U284);
  not ginst1147 (P1_R1117_U287, P1_R1117_U156);
  nand ginst1148 (P1_R1117_U288, P1_R1117_U77, P1_U3978);
  nand ginst1149 (P1_R1117_U289, P1_R1117_U156, P1_R1117_U288);
  not ginst1150 (P1_R1117_U29, P1_U3470);
  nand ginst1151 (P1_R1117_U290, P1_R1117_U76, P1_U3065);
  not ginst1152 (P1_R1117_U291, P1_R1117_U155);
  nand ginst1153 (P1_R1117_U292, P1_R1117_U79, P1_U3977);
  nand ginst1154 (P1_R1117_U293, P1_R1117_U155, P1_R1117_U292);
  nand ginst1155 (P1_R1117_U294, P1_R1117_U78, P1_U3058);
  not ginst1156 (P1_R1117_U295, P1_R1117_U87);
  nand ginst1157 (P1_R1117_U296, P1_R1117_U83, P1_U3975);
  nand ginst1158 (P1_R1117_U297, P1_R1117_U177, P1_R1117_U296, P1_R1117_U87);
  nand ginst1159 (P1_R1117_U298, P1_R1117_U82, P1_R1117_U83);
  nand ginst1160 (P1_R1117_U299, P1_R1117_U298, P1_R1117_U80);
  not ginst1161 (P1_R1117_U30, P1_U3464);
  nand ginst1162 (P1_R1117_U300, P1_R1117_U171, P1_U3053);
  not ginst1163 (P1_R1117_U301, P1_R1117_U86);
  nand ginst1164 (P1_R1117_U302, P1_R1117_U84, P1_U3054);
  nand ginst1165 (P1_R1117_U303, P1_R1117_U301, P1_R1117_U302);
  nand ginst1166 (P1_R1117_U304, P1_R1117_U85, P1_U3974);
  nand ginst1167 (P1_R1117_U305, P1_R1117_U85, P1_U3974);
  nand ginst1168 (P1_R1117_U306, P1_R1117_U305, P1_R1117_U86);
  nand ginst1169 (P1_R1117_U307, P1_R1117_U84, P1_U3054);
  nand ginst1170 (P1_R1117_U308, P1_R1117_U153, P1_R1117_U306, P1_R1117_U307);
  nand ginst1171 (P1_R1117_U309, P1_R1117_U295, P1_R1117_U82);
  not ginst1172 (P1_R1117_U31, P1_U3071);
  nand ginst1173 (P1_R1117_U310, P1_R1117_U129, P1_R1117_U309);
  nand ginst1174 (P1_R1117_U311, P1_R1117_U177, P1_R1117_U87);
  nand ginst1175 (P1_R1117_U312, P1_R1117_U128, P1_R1117_U311);
  nand ginst1176 (P1_R1117_U313, P1_R1117_U177, P1_R1117_U82);
  nand ginst1177 (P1_R1117_U314, P1_R1117_U159, P1_R1117_U283);
  not ginst1178 (P1_R1117_U315, P1_R1117_U88);
  nand ginst1179 (P1_R1117_U316, P1_R1117_U45, P1_U3061);
  nand ginst1180 (P1_R1117_U317, P1_R1117_U315, P1_R1117_U316);
  nand ginst1181 (P1_R1117_U318, P1_R1117_U132, P1_R1117_U317);
  nand ginst1182 (P1_R1117_U319, P1_R1117_U176, P1_R1117_U88);
  not ginst1183 (P1_R1117_U32, P1_U3067);
  nand ginst1184 (P1_R1117_U320, P1_R1117_U72, P1_U3979);
  nand ginst1185 (P1_R1117_U321, P1_R1117_U319, P1_R1117_U320, P1_R1117_U9);
  nand ginst1186 (P1_R1117_U322, P1_R1117_U45, P1_U3061);
  nand ginst1187 (P1_R1117_U323, P1_R1117_U176, P1_R1117_U322);
  nand ginst1188 (P1_R1117_U324, P1_R1117_U283, P1_R1117_U75);
  nand ginst1189 (P1_R1117_U325, P1_R1117_U167, P1_R1117_U257);
  not ginst1190 (P1_R1117_U326, P1_R1117_U89);
  nand ginst1191 (P1_R1117_U327, P1_R1117_U46, P1_U3074);
  nand ginst1192 (P1_R1117_U328, P1_R1117_U326, P1_R1117_U327);
  nand ginst1193 (P1_R1117_U329, P1_R1117_U139, P1_R1117_U328);
  not ginst1194 (P1_R1117_U33, P1_U3060);
  nand ginst1195 (P1_R1117_U330, P1_R1117_U175, P1_R1117_U89);
  nand ginst1196 (P1_R1117_U331, P1_R1117_U58, P1_U3500);
  nand ginst1197 (P1_R1117_U332, P1_R1117_U138, P1_R1117_U330);
  nand ginst1198 (P1_R1117_U333, P1_R1117_U46, P1_U3074);
  nand ginst1199 (P1_R1117_U334, P1_R1117_U175, P1_R1117_U333);
  nand ginst1200 (P1_R1117_U335, P1_R1117_U257, P1_R1117_U61);
  nand ginst1201 (P1_R1117_U336, P1_R1117_U145, P1_R1117_U212);
  not ginst1202 (P1_R1117_U337, P1_R1117_U90);
  nand ginst1203 (P1_R1117_U338, P1_R1117_U47, P1_U3062);
  nand ginst1204 (P1_R1117_U339, P1_R1117_U337, P1_R1117_U338);
  nand ginst1205 (P1_R1117_U34, P1_R1117_U30, P1_U3060);
  nand ginst1206 (P1_R1117_U340, P1_R1117_U143, P1_R1117_U339);
  nand ginst1207 (P1_R1117_U341, P1_R1117_U174, P1_R1117_U90);
  nand ginst1208 (P1_R1117_U342, P1_R1117_U49, P1_U3485);
  nand ginst1209 (P1_R1117_U343, P1_R1117_U142, P1_R1117_U341);
  nand ginst1210 (P1_R1117_U344, P1_R1117_U47, P1_U3062);
  nand ginst1211 (P1_R1117_U345, P1_R1117_U174, P1_R1117_U344);
  nand ginst1212 (P1_R1117_U346, P1_R1117_U22, P1_U3077);
  nand ginst1213 (P1_R1117_U347, P1_R1117_U303, P1_R1117_U304, P1_R1117_U385);
  nand ginst1214 (P1_R1117_U348, P1_R1117_U40, P1_U3479);
  nand ginst1215 (P1_R1117_U349, P1_R1117_U39, P1_U3083);
  not ginst1216 (P1_R1117_U35, P1_U3476);
  nand ginst1217 (P1_R1117_U350, P1_R1117_U145, P1_R1117_U213);
  nand ginst1218 (P1_R1117_U351, P1_R1117_U144, P1_R1117_U211);
  nand ginst1219 (P1_R1117_U352, P1_R1117_U38, P1_U3476);
  nand ginst1220 (P1_R1117_U353, P1_R1117_U35, P1_U3084);
  nand ginst1221 (P1_R1117_U354, P1_R1117_U38, P1_U3476);
  nand ginst1222 (P1_R1117_U355, P1_R1117_U35, P1_U3084);
  nand ginst1223 (P1_R1117_U356, P1_R1117_U354, P1_R1117_U355);
  nand ginst1224 (P1_R1117_U357, P1_R1117_U36, P1_U3473);
  nand ginst1225 (P1_R1117_U358, P1_R1117_U19, P1_U3070);
  nand ginst1226 (P1_R1117_U359, P1_R1117_U218, P1_R1117_U41);
  not ginst1227 (P1_R1117_U36, P1_U3070);
  nand ginst1228 (P1_R1117_U360, P1_R1117_U146, P1_R1117_U205);
  nand ginst1229 (P1_R1117_U361, P1_R1117_U31, P1_U3470);
  nand ginst1230 (P1_R1117_U362, P1_R1117_U29, P1_U3071);
  nand ginst1231 (P1_R1117_U363, P1_R1117_U361, P1_R1117_U362);
  nand ginst1232 (P1_R1117_U364, P1_R1117_U32, P1_U3467);
  nand ginst1233 (P1_R1117_U365, P1_R1117_U20, P1_U3067);
  nand ginst1234 (P1_R1117_U366, P1_R1117_U228, P1_R1117_U42);
  nand ginst1235 (P1_R1117_U367, P1_R1117_U147, P1_R1117_U220);
  nand ginst1236 (P1_R1117_U368, P1_R1117_U33, P1_U3464);
  nand ginst1237 (P1_R1117_U369, P1_R1117_U30, P1_U3060);
  nand ginst1238 (P1_R1117_U37, P1_R1117_U19, P1_U3070);
  nand ginst1239 (P1_R1117_U370, P1_R1117_U149, P1_R1117_U229);
  nand ginst1240 (P1_R1117_U371, P1_R1117_U148, P1_R1117_U195);
  nand ginst1241 (P1_R1117_U372, P1_R1117_U28, P1_U3461);
  nand ginst1242 (P1_R1117_U373, P1_R1117_U25, P1_U3064);
  nand ginst1243 (P1_R1117_U374, P1_R1117_U28, P1_U3461);
  nand ginst1244 (P1_R1117_U375, P1_R1117_U25, P1_U3064);
  nand ginst1245 (P1_R1117_U376, P1_R1117_U374, P1_R1117_U375);
  nand ginst1246 (P1_R1117_U377, P1_R1117_U26, P1_U3458);
  nand ginst1247 (P1_R1117_U378, P1_R1117_U21, P1_U3068);
  nand ginst1248 (P1_R1117_U379, P1_R1117_U234, P1_R1117_U43);
  not ginst1249 (P1_R1117_U38, P1_U3084);
  nand ginst1250 (P1_R1117_U380, P1_R1117_U150, P1_R1117_U189);
  nand ginst1251 (P1_R1117_U381, P1_R1117_U152, P1_U3985);
  nand ginst1252 (P1_R1117_U382, P1_R1117_U151, P1_U3055);
  nand ginst1253 (P1_R1117_U383, P1_R1117_U152, P1_U3985);
  nand ginst1254 (P1_R1117_U384, P1_R1117_U151, P1_U3055);
  nand ginst1255 (P1_R1117_U385, P1_R1117_U383, P1_R1117_U384);
  nand ginst1256 (P1_R1117_U386, P1_R1117_U85, P1_U3974);
  nand ginst1257 (P1_R1117_U387, P1_R1117_U84, P1_U3054);
  not ginst1258 (P1_R1117_U388, P1_R1117_U127);
  nand ginst1259 (P1_R1117_U389, P1_R1117_U301, P1_R1117_U388);
  not ginst1260 (P1_R1117_U39, P1_U3479);
  nand ginst1261 (P1_R1117_U390, P1_R1117_U127, P1_R1117_U86);
  nand ginst1262 (P1_R1117_U391, P1_R1117_U83, P1_U3975);
  nand ginst1263 (P1_R1117_U392, P1_R1117_U80, P1_U3053);
  nand ginst1264 (P1_R1117_U393, P1_R1117_U83, P1_U3975);
  nand ginst1265 (P1_R1117_U394, P1_R1117_U80, P1_U3053);
  nand ginst1266 (P1_R1117_U395, P1_R1117_U393, P1_R1117_U394);
  nand ginst1267 (P1_R1117_U396, P1_R1117_U81, P1_U3976);
  nand ginst1268 (P1_R1117_U397, P1_R1117_U44, P1_U3057);
  nand ginst1269 (P1_R1117_U398, P1_R1117_U313, P1_R1117_U87);
  nand ginst1270 (P1_R1117_U399, P1_R1117_U154, P1_R1117_U295);
  not ginst1271 (P1_R1117_U40, P1_U3083);
  nand ginst1272 (P1_R1117_U400, P1_R1117_U79, P1_U3977);
  nand ginst1273 (P1_R1117_U401, P1_R1117_U78, P1_U3058);
  not ginst1274 (P1_R1117_U402, P1_R1117_U130);
  nand ginst1275 (P1_R1117_U403, P1_R1117_U291, P1_R1117_U402);
  nand ginst1276 (P1_R1117_U404, P1_R1117_U130, P1_R1117_U155);
  nand ginst1277 (P1_R1117_U405, P1_R1117_U77, P1_U3978);
  nand ginst1278 (P1_R1117_U406, P1_R1117_U76, P1_U3065);
  not ginst1279 (P1_R1117_U407, P1_R1117_U131);
  nand ginst1280 (P1_R1117_U408, P1_R1117_U287, P1_R1117_U407);
  nand ginst1281 (P1_R1117_U409, P1_R1117_U131, P1_R1117_U156);
  nand ginst1282 (P1_R1117_U41, P1_R1117_U203, P1_R1117_U204);
  nand ginst1283 (P1_R1117_U410, P1_R1117_U72, P1_U3979);
  nand ginst1284 (P1_R1117_U411, P1_R1117_U70, P1_U3066);
  nand ginst1285 (P1_R1117_U412, P1_R1117_U410, P1_R1117_U411);
  nand ginst1286 (P1_R1117_U413, P1_R1117_U73, P1_U3980);
  nand ginst1287 (P1_R1117_U414, P1_R1117_U45, P1_U3061);
  nand ginst1288 (P1_R1117_U415, P1_R1117_U323, P1_R1117_U88);
  nand ginst1289 (P1_R1117_U416, P1_R1117_U157, P1_R1117_U315);
  nand ginst1290 (P1_R1117_U417, P1_R1117_U74, P1_U3981);
  nand ginst1291 (P1_R1117_U418, P1_R1117_U71, P1_U3075);
  nand ginst1292 (P1_R1117_U419, P1_R1117_U159, P1_R1117_U324);
  nand ginst1293 (P1_R1117_U42, P1_R1117_U219, P1_R1117_U34);
  nand ginst1294 (P1_R1117_U420, P1_R1117_U158, P1_R1117_U277);
  nand ginst1295 (P1_R1117_U421, P1_R1117_U69, P1_U3982);
  nand ginst1296 (P1_R1117_U422, P1_R1117_U68, P1_U3076);
  not ginst1297 (P1_R1117_U423, P1_R1117_U133);
  nand ginst1298 (P1_R1117_U424, P1_R1117_U273, P1_R1117_U423);
  nand ginst1299 (P1_R1117_U425, P1_R1117_U133, P1_R1117_U160);
  nand ginst1300 (P1_R1117_U426, P1_R1117_U185, P1_R1117_U24);
  nand ginst1301 (P1_R1117_U427, P1_R1117_U23, P1_U3078);
  not ginst1302 (P1_R1117_U428, P1_R1117_U134);
  nand ginst1303 (P1_R1117_U429, P1_R1117_U428, P1_U3455);
  nand ginst1304 (P1_R1117_U43, P1_R1117_U187, P1_R1117_U188);
  nand ginst1305 (P1_R1117_U430, P1_R1117_U134, P1_R1117_U161);
  nand ginst1306 (P1_R1117_U431, P1_R1117_U67, P1_U3508);
  nand ginst1307 (P1_R1117_U432, P1_R1117_U66, P1_U3081);
  not ginst1308 (P1_R1117_U433, P1_R1117_U135);
  nand ginst1309 (P1_R1117_U434, P1_R1117_U269, P1_R1117_U433);
  nand ginst1310 (P1_R1117_U435, P1_R1117_U135, P1_R1117_U162);
  nand ginst1311 (P1_R1117_U436, P1_R1117_U65, P1_U3506);
  nand ginst1312 (P1_R1117_U437, P1_R1117_U163, P1_U3082);
  not ginst1313 (P1_R1117_U438, P1_R1117_U136);
  nand ginst1314 (P1_R1117_U439, P1_R1117_U265, P1_R1117_U438);
  not ginst1315 (P1_R1117_U44, P1_U3976);
  nand ginst1316 (P1_R1117_U440, P1_R1117_U136, P1_R1117_U64);
  nand ginst1317 (P1_R1117_U441, P1_R1117_U63, P1_U3503);
  nand ginst1318 (P1_R1117_U442, P1_R1117_U62, P1_U3069);
  not ginst1319 (P1_R1117_U443, P1_R1117_U137);
  nand ginst1320 (P1_R1117_U444, P1_R1117_U261, P1_R1117_U443);
  nand ginst1321 (P1_R1117_U445, P1_R1117_U137, P1_R1117_U164);
  nand ginst1322 (P1_R1117_U446, P1_R1117_U58, P1_U3500);
  nand ginst1323 (P1_R1117_U447, P1_R1117_U56, P1_U3073);
  nand ginst1324 (P1_R1117_U448, P1_R1117_U446, P1_R1117_U447);
  nand ginst1325 (P1_R1117_U449, P1_R1117_U59, P1_U3497);
  not ginst1326 (P1_R1117_U45, P1_U3980);
  nand ginst1327 (P1_R1117_U450, P1_R1117_U46, P1_U3074);
  nand ginst1328 (P1_R1117_U451, P1_R1117_U334, P1_R1117_U89);
  nand ginst1329 (P1_R1117_U452, P1_R1117_U165, P1_R1117_U326);
  nand ginst1330 (P1_R1117_U453, P1_R1117_U60, P1_U3494);
  nand ginst1331 (P1_R1117_U454, P1_R1117_U57, P1_U3079);
  nand ginst1332 (P1_R1117_U455, P1_R1117_U167, P1_R1117_U335);
  nand ginst1333 (P1_R1117_U456, P1_R1117_U166, P1_R1117_U251);
  nand ginst1334 (P1_R1117_U457, P1_R1117_U55, P1_U3491);
  nand ginst1335 (P1_R1117_U458, P1_R1117_U54, P1_U3080);
  not ginst1336 (P1_R1117_U459, P1_R1117_U140);
  not ginst1337 (P1_R1117_U46, P1_U3497);
  nand ginst1338 (P1_R1117_U460, P1_R1117_U247, P1_R1117_U459);
  nand ginst1339 (P1_R1117_U461, P1_R1117_U140, P1_R1117_U168);
  nand ginst1340 (P1_R1117_U462, P1_R1117_U53, P1_U3488);
  nand ginst1341 (P1_R1117_U463, P1_R1117_U52, P1_U3072);
  not ginst1342 (P1_R1117_U464, P1_R1117_U141);
  nand ginst1343 (P1_R1117_U465, P1_R1117_U243, P1_R1117_U464);
  nand ginst1344 (P1_R1117_U466, P1_R1117_U141, P1_R1117_U169);
  nand ginst1345 (P1_R1117_U467, P1_R1117_U49, P1_U3485);
  nand ginst1346 (P1_R1117_U468, P1_R1117_U48, P1_U3063);
  nand ginst1347 (P1_R1117_U469, P1_R1117_U467, P1_R1117_U468);
  not ginst1348 (P1_R1117_U47, P1_U3482);
  nand ginst1349 (P1_R1117_U470, P1_R1117_U50, P1_U3482);
  nand ginst1350 (P1_R1117_U471, P1_R1117_U47, P1_U3062);
  nand ginst1351 (P1_R1117_U472, P1_R1117_U345, P1_R1117_U90);
  nand ginst1352 (P1_R1117_U473, P1_R1117_U170, P1_R1117_U337);
  not ginst1353 (P1_R1117_U48, P1_U3485);
  not ginst1354 (P1_R1117_U49, P1_U3063);
  not ginst1355 (P1_R1117_U50, P1_U3062);
  nand ginst1356 (P1_R1117_U51, P1_R1117_U39, P1_U3083);
  not ginst1357 (P1_R1117_U52, P1_U3488);
  not ginst1358 (P1_R1117_U53, P1_U3072);
  not ginst1359 (P1_R1117_U54, P1_U3491);
  not ginst1360 (P1_R1117_U55, P1_U3080);
  not ginst1361 (P1_R1117_U56, P1_U3500);
  not ginst1362 (P1_R1117_U57, P1_U3494);
  not ginst1363 (P1_R1117_U58, P1_U3073);
  not ginst1364 (P1_R1117_U59, P1_U3074);
  and ginst1365 (P1_R1117_U6, P1_R1117_U197, P1_R1117_U198);
  not ginst1366 (P1_R1117_U60, P1_U3079);
  nand ginst1367 (P1_R1117_U61, P1_R1117_U57, P1_U3079);
  not ginst1368 (P1_R1117_U62, P1_U3503);
  not ginst1369 (P1_R1117_U63, P1_U3069);
  nand ginst1370 (P1_R1117_U64, P1_R1117_U263, P1_R1117_U264);
  not ginst1371 (P1_R1117_U65, P1_U3082);
  not ginst1372 (P1_R1117_U66, P1_U3508);
  not ginst1373 (P1_R1117_U67, P1_U3081);
  not ginst1374 (P1_R1117_U68, P1_U3982);
  not ginst1375 (P1_R1117_U69, P1_U3076);
  and ginst1376 (P1_R1117_U7, P1_R1117_U236, P1_R1117_U237);
  not ginst1377 (P1_R1117_U70, P1_U3979);
  not ginst1378 (P1_R1117_U71, P1_U3981);
  not ginst1379 (P1_R1117_U72, P1_U3066);
  not ginst1380 (P1_R1117_U73, P1_U3061);
  not ginst1381 (P1_R1117_U74, P1_U3075);
  nand ginst1382 (P1_R1117_U75, P1_R1117_U71, P1_U3075);
  not ginst1383 (P1_R1117_U76, P1_U3978);
  not ginst1384 (P1_R1117_U77, P1_U3065);
  not ginst1385 (P1_R1117_U78, P1_U3977);
  not ginst1386 (P1_R1117_U79, P1_U3058);
  and ginst1387 (P1_R1117_U8, P1_R1117_U253, P1_R1117_U254);
  not ginst1388 (P1_R1117_U80, P1_U3975);
  not ginst1389 (P1_R1117_U81, P1_U3057);
  nand ginst1390 (P1_R1117_U82, P1_R1117_U44, P1_U3057);
  not ginst1391 (P1_R1117_U83, P1_U3053);
  not ginst1392 (P1_R1117_U84, P1_U3974);
  not ginst1393 (P1_R1117_U85, P1_U3054);
  nand ginst1394 (P1_R1117_U86, P1_R1117_U126, P1_R1117_U297);
  nand ginst1395 (P1_R1117_U87, P1_R1117_U293, P1_R1117_U294);
  nand ginst1396 (P1_R1117_U88, P1_R1117_U314, P1_R1117_U75);
  nand ginst1397 (P1_R1117_U89, P1_R1117_U325, P1_R1117_U61);
  and ginst1398 (P1_R1117_U9, P1_R1117_U279, P1_R1117_U280);
  nand ginst1399 (P1_R1117_U90, P1_R1117_U336, P1_R1117_U51);
  not ginst1400 (P1_R1117_U91, P1_U3077);
  nand ginst1401 (P1_R1117_U92, P1_R1117_U389, P1_R1117_U390);
  nand ginst1402 (P1_R1117_U93, P1_R1117_U403, P1_R1117_U404);
  nand ginst1403 (P1_R1117_U94, P1_R1117_U408, P1_R1117_U409);
  nand ginst1404 (P1_R1117_U95, P1_R1117_U424, P1_R1117_U425);
  nand ginst1405 (P1_R1117_U96, P1_R1117_U429, P1_R1117_U430);
  nand ginst1406 (P1_R1117_U97, P1_R1117_U434, P1_R1117_U435);
  nand ginst1407 (P1_R1117_U98, P1_R1117_U439, P1_R1117_U440);
  nand ginst1408 (P1_R1117_U99, P1_R1117_U444, P1_R1117_U445);
  and ginst1409 (P1_R1138_U10, P1_R1138_U270, P1_R1138_U271);
  nand ginst1410 (P1_R1138_U100, P1_R1138_U392, P1_R1138_U393);
  nand ginst1411 (P1_R1138_U101, P1_R1138_U397, P1_R1138_U398);
  nand ginst1412 (P1_R1138_U102, P1_R1138_U406, P1_R1138_U407);
  nand ginst1413 (P1_R1138_U103, P1_R1138_U413, P1_R1138_U414);
  nand ginst1414 (P1_R1138_U104, P1_R1138_U420, P1_R1138_U421);
  nand ginst1415 (P1_R1138_U105, P1_R1138_U427, P1_R1138_U428);
  nand ginst1416 (P1_R1138_U106, P1_R1138_U432, P1_R1138_U433);
  nand ginst1417 (P1_R1138_U107, P1_R1138_U439, P1_R1138_U440);
  nand ginst1418 (P1_R1138_U108, P1_R1138_U446, P1_R1138_U447);
  nand ginst1419 (P1_R1138_U109, P1_R1138_U460, P1_R1138_U461);
  and ginst1420 (P1_R1138_U11, P1_R1138_U347, P1_R1138_U350);
  nand ginst1421 (P1_R1138_U110, P1_R1138_U465, P1_R1138_U466);
  nand ginst1422 (P1_R1138_U111, P1_R1138_U472, P1_R1138_U473);
  nand ginst1423 (P1_R1138_U112, P1_R1138_U479, P1_R1138_U480);
  nand ginst1424 (P1_R1138_U113, P1_R1138_U486, P1_R1138_U487);
  nand ginst1425 (P1_R1138_U114, P1_R1138_U493, P1_R1138_U494);
  nand ginst1426 (P1_R1138_U115, P1_R1138_U498, P1_R1138_U499);
  and ginst1427 (P1_R1138_U116, P1_U3068, P1_U3458);
  and ginst1428 (P1_R1138_U117, P1_R1138_U186, P1_R1138_U188);
  and ginst1429 (P1_R1138_U118, P1_R1138_U191, P1_R1138_U193);
  and ginst1430 (P1_R1138_U119, P1_R1138_U199, P1_R1138_U200);
  and ginst1431 (P1_R1138_U12, P1_R1138_U340, P1_R1138_U343);
  and ginst1432 (P1_R1138_U120, P1_R1138_U23, P1_R1138_U380, P1_R1138_U381);
  and ginst1433 (P1_R1138_U121, P1_R1138_U211, P1_R1138_U6);
  and ginst1434 (P1_R1138_U122, P1_R1138_U217, P1_R1138_U219);
  and ginst1435 (P1_R1138_U123, P1_R1138_U35, P1_R1138_U387, P1_R1138_U388);
  and ginst1436 (P1_R1138_U124, P1_R1138_U225, P1_R1138_U4);
  and ginst1437 (P1_R1138_U125, P1_R1138_U180, P1_R1138_U233);
  and ginst1438 (P1_R1138_U126, P1_R1138_U203, P1_R1138_U7);
  and ginst1439 (P1_R1138_U127, P1_R1138_U170, P1_R1138_U238);
  and ginst1440 (P1_R1138_U128, P1_R1138_U249, P1_R1138_U8);
  and ginst1441 (P1_R1138_U129, P1_R1138_U171, P1_R1138_U247);
  and ginst1442 (P1_R1138_U13, P1_R1138_U331, P1_R1138_U334);
  and ginst1443 (P1_R1138_U130, P1_R1138_U266, P1_R1138_U267);
  and ginst1444 (P1_R1138_U131, P1_R1138_U10, P1_R1138_U281);
  and ginst1445 (P1_R1138_U132, P1_R1138_U279, P1_R1138_U284);
  and ginst1446 (P1_R1138_U133, P1_R1138_U297, P1_R1138_U300);
  and ginst1447 (P1_R1138_U134, P1_R1138_U301, P1_R1138_U367);
  and ginst1448 (P1_R1138_U135, P1_R1138_U159, P1_R1138_U277);
  and ginst1449 (P1_R1138_U136, P1_R1138_U453, P1_R1138_U454, P1_R1138_U81);
  and ginst1450 (P1_R1138_U137, P1_R1138_U467, P1_R1138_U468, P1_R1138_U60);
  and ginst1451 (P1_R1138_U138, P1_R1138_U333, P1_R1138_U9);
  and ginst1452 (P1_R1138_U139, P1_R1138_U171, P1_R1138_U488, P1_R1138_U489);
  and ginst1453 (P1_R1138_U14, P1_R1138_U322, P1_R1138_U325);
  and ginst1454 (P1_R1138_U140, P1_R1138_U342, P1_R1138_U8);
  and ginst1455 (P1_R1138_U141, P1_R1138_U170, P1_R1138_U500, P1_R1138_U501);
  and ginst1456 (P1_R1138_U142, P1_R1138_U349, P1_R1138_U7);
  nand ginst1457 (P1_R1138_U143, P1_R1138_U119, P1_R1138_U201);
  nand ginst1458 (P1_R1138_U144, P1_R1138_U216, P1_R1138_U228);
  not ginst1459 (P1_R1138_U145, P1_U3055);
  not ginst1460 (P1_R1138_U146, P1_U3985);
  and ginst1461 (P1_R1138_U147, P1_R1138_U401, P1_R1138_U402);
  nand ginst1462 (P1_R1138_U148, P1_R1138_U168, P1_R1138_U303, P1_R1138_U363);
  and ginst1463 (P1_R1138_U149, P1_R1138_U408, P1_R1138_U409);
  and ginst1464 (P1_R1138_U15, P1_R1138_U317, P1_R1138_U319);
  nand ginst1465 (P1_R1138_U150, P1_R1138_U134, P1_R1138_U368, P1_R1138_U369);
  and ginst1466 (P1_R1138_U151, P1_R1138_U415, P1_R1138_U416);
  nand ginst1467 (P1_R1138_U152, P1_R1138_U298, P1_R1138_U364, P1_R1138_U87);
  and ginst1468 (P1_R1138_U153, P1_R1138_U422, P1_R1138_U423);
  nand ginst1469 (P1_R1138_U154, P1_R1138_U291, P1_R1138_U292);
  and ginst1470 (P1_R1138_U155, P1_R1138_U434, P1_R1138_U435);
  nand ginst1471 (P1_R1138_U156, P1_R1138_U287, P1_R1138_U288);
  and ginst1472 (P1_R1138_U157, P1_R1138_U441, P1_R1138_U442);
  nand ginst1473 (P1_R1138_U158, P1_R1138_U132, P1_R1138_U283);
  and ginst1474 (P1_R1138_U159, P1_R1138_U448, P1_R1138_U449);
  and ginst1475 (P1_R1138_U16, P1_R1138_U309, P1_R1138_U312);
  nand ginst1476 (P1_R1138_U160, P1_R1138_U326, P1_R1138_U44);
  nand ginst1477 (P1_R1138_U161, P1_R1138_U130, P1_R1138_U268);
  and ginst1478 (P1_R1138_U162, P1_R1138_U474, P1_R1138_U475);
  nand ginst1479 (P1_R1138_U163, P1_R1138_U255, P1_R1138_U256);
  and ginst1480 (P1_R1138_U164, P1_R1138_U481, P1_R1138_U482);
  nand ginst1481 (P1_R1138_U165, P1_R1138_U251, P1_R1138_U252);
  nand ginst1482 (P1_R1138_U166, P1_R1138_U241, P1_R1138_U242);
  nand ginst1483 (P1_R1138_U167, P1_R1138_U365, P1_R1138_U366);
  nand ginst1484 (P1_R1138_U168, P1_R1138_U150, P1_U3054);
  not ginst1485 (P1_R1138_U169, P1_R1138_U35);
  and ginst1486 (P1_R1138_U17, P1_R1138_U231, P1_R1138_U234);
  nand ginst1487 (P1_R1138_U170, P1_U3083, P1_U3479);
  nand ginst1488 (P1_R1138_U171, P1_U3072, P1_U3488);
  nand ginst1489 (P1_R1138_U172, P1_U3058, P1_U3977);
  not ginst1490 (P1_R1138_U173, P1_R1138_U69);
  not ginst1491 (P1_R1138_U174, P1_R1138_U78);
  nand ginst1492 (P1_R1138_U175, P1_U3065, P1_U3978);
  not ginst1493 (P1_R1138_U176, P1_R1138_U62);
  or ginst1494 (P1_R1138_U177, P1_U3067, P1_U3467);
  or ginst1495 (P1_R1138_U178, P1_U3060, P1_U3464);
  or ginst1496 (P1_R1138_U179, P1_U3064, P1_U3461);
  and ginst1497 (P1_R1138_U18, P1_R1138_U223, P1_R1138_U226);
  or ginst1498 (P1_R1138_U180, P1_U3068, P1_U3458);
  not ginst1499 (P1_R1138_U181, P1_R1138_U32);
  or ginst1500 (P1_R1138_U182, P1_U3078, P1_U3455);
  not ginst1501 (P1_R1138_U183, P1_R1138_U43);
  not ginst1502 (P1_R1138_U184, P1_R1138_U44);
  nand ginst1503 (P1_R1138_U185, P1_R1138_U43, P1_R1138_U44);
  nand ginst1504 (P1_R1138_U186, P1_R1138_U116, P1_R1138_U179);
  nand ginst1505 (P1_R1138_U187, P1_R1138_U185, P1_R1138_U5);
  nand ginst1506 (P1_R1138_U188, P1_U3064, P1_U3461);
  nand ginst1507 (P1_R1138_U189, P1_R1138_U117, P1_R1138_U187);
  and ginst1508 (P1_R1138_U19, P1_R1138_U209, P1_R1138_U212);
  nand ginst1509 (P1_R1138_U190, P1_R1138_U35, P1_R1138_U36);
  nand ginst1510 (P1_R1138_U191, P1_R1138_U190, P1_U3067);
  nand ginst1511 (P1_R1138_U192, P1_R1138_U189, P1_R1138_U4);
  nand ginst1512 (P1_R1138_U193, P1_R1138_U169, P1_U3467);
  not ginst1513 (P1_R1138_U194, P1_R1138_U42);
  or ginst1514 (P1_R1138_U195, P1_U3070, P1_U3473);
  or ginst1515 (P1_R1138_U196, P1_U3071, P1_U3470);
  not ginst1516 (P1_R1138_U197, P1_R1138_U23);
  nand ginst1517 (P1_R1138_U198, P1_R1138_U23, P1_R1138_U24);
  nand ginst1518 (P1_R1138_U199, P1_R1138_U198, P1_U3070);
  not ginst1519 (P1_R1138_U20, P1_U3470);
  nand ginst1520 (P1_R1138_U200, P1_R1138_U197, P1_U3473);
  nand ginst1521 (P1_R1138_U201, P1_R1138_U42, P1_R1138_U6);
  not ginst1522 (P1_R1138_U202, P1_R1138_U143);
  or ginst1523 (P1_R1138_U203, P1_U3084, P1_U3476);
  nand ginst1524 (P1_R1138_U204, P1_R1138_U143, P1_R1138_U203);
  not ginst1525 (P1_R1138_U205, P1_R1138_U41);
  or ginst1526 (P1_R1138_U206, P1_U3083, P1_U3479);
  or ginst1527 (P1_R1138_U207, P1_U3071, P1_U3470);
  nand ginst1528 (P1_R1138_U208, P1_R1138_U207, P1_R1138_U42);
  nand ginst1529 (P1_R1138_U209, P1_R1138_U120, P1_R1138_U208);
  not ginst1530 (P1_R1138_U21, P1_U3071);
  nand ginst1531 (P1_R1138_U210, P1_R1138_U194, P1_R1138_U23);
  nand ginst1532 (P1_R1138_U211, P1_U3070, P1_U3473);
  nand ginst1533 (P1_R1138_U212, P1_R1138_U121, P1_R1138_U210);
  or ginst1534 (P1_R1138_U213, P1_U3071, P1_U3470);
  nand ginst1535 (P1_R1138_U214, P1_R1138_U180, P1_R1138_U184);
  nand ginst1536 (P1_R1138_U215, P1_U3068, P1_U3458);
  not ginst1537 (P1_R1138_U216, P1_R1138_U46);
  nand ginst1538 (P1_R1138_U217, P1_R1138_U183, P1_R1138_U5);
  nand ginst1539 (P1_R1138_U218, P1_R1138_U179, P1_R1138_U46);
  nand ginst1540 (P1_R1138_U219, P1_U3064, P1_U3461);
  not ginst1541 (P1_R1138_U22, P1_U3070);
  not ginst1542 (P1_R1138_U220, P1_R1138_U45);
  or ginst1543 (P1_R1138_U221, P1_U3060, P1_U3464);
  nand ginst1544 (P1_R1138_U222, P1_R1138_U221, P1_R1138_U45);
  nand ginst1545 (P1_R1138_U223, P1_R1138_U123, P1_R1138_U222);
  nand ginst1546 (P1_R1138_U224, P1_R1138_U220, P1_R1138_U35);
  nand ginst1547 (P1_R1138_U225, P1_U3067, P1_U3467);
  nand ginst1548 (P1_R1138_U226, P1_R1138_U124, P1_R1138_U224);
  or ginst1549 (P1_R1138_U227, P1_U3060, P1_U3464);
  nand ginst1550 (P1_R1138_U228, P1_R1138_U180, P1_R1138_U183);
  not ginst1551 (P1_R1138_U229, P1_R1138_U144);
  nand ginst1552 (P1_R1138_U23, P1_U3071, P1_U3470);
  nand ginst1553 (P1_R1138_U230, P1_U3064, P1_U3461);
  nand ginst1554 (P1_R1138_U231, P1_R1138_U399, P1_R1138_U400, P1_R1138_U43, P1_R1138_U44);
  nand ginst1555 (P1_R1138_U232, P1_R1138_U43, P1_R1138_U44);
  nand ginst1556 (P1_R1138_U233, P1_U3068, P1_U3458);
  nand ginst1557 (P1_R1138_U234, P1_R1138_U125, P1_R1138_U232);
  or ginst1558 (P1_R1138_U235, P1_U3083, P1_U3479);
  or ginst1559 (P1_R1138_U236, P1_U3062, P1_U3482);
  nand ginst1560 (P1_R1138_U237, P1_R1138_U176, P1_R1138_U7);
  nand ginst1561 (P1_R1138_U238, P1_U3062, P1_U3482);
  nand ginst1562 (P1_R1138_U239, P1_R1138_U127, P1_R1138_U237);
  not ginst1563 (P1_R1138_U24, P1_U3473);
  or ginst1564 (P1_R1138_U240, P1_U3062, P1_U3482);
  nand ginst1565 (P1_R1138_U241, P1_R1138_U126, P1_R1138_U143);
  nand ginst1566 (P1_R1138_U242, P1_R1138_U239, P1_R1138_U240);
  not ginst1567 (P1_R1138_U243, P1_R1138_U166);
  or ginst1568 (P1_R1138_U244, P1_U3080, P1_U3491);
  or ginst1569 (P1_R1138_U245, P1_U3072, P1_U3488);
  nand ginst1570 (P1_R1138_U246, P1_R1138_U173, P1_R1138_U8);
  nand ginst1571 (P1_R1138_U247, P1_U3080, P1_U3491);
  nand ginst1572 (P1_R1138_U248, P1_R1138_U129, P1_R1138_U246);
  or ginst1573 (P1_R1138_U249, P1_U3063, P1_U3485);
  not ginst1574 (P1_R1138_U25, P1_U3464);
  or ginst1575 (P1_R1138_U250, P1_U3080, P1_U3491);
  nand ginst1576 (P1_R1138_U251, P1_R1138_U128, P1_R1138_U166);
  nand ginst1577 (P1_R1138_U252, P1_R1138_U248, P1_R1138_U250);
  not ginst1578 (P1_R1138_U253, P1_R1138_U165);
  or ginst1579 (P1_R1138_U254, P1_U3079, P1_U3494);
  nand ginst1580 (P1_R1138_U255, P1_R1138_U165, P1_R1138_U254);
  nand ginst1581 (P1_R1138_U256, P1_U3079, P1_U3494);
  not ginst1582 (P1_R1138_U257, P1_R1138_U163);
  or ginst1583 (P1_R1138_U258, P1_U3074, P1_U3497);
  nand ginst1584 (P1_R1138_U259, P1_R1138_U163, P1_R1138_U258);
  not ginst1585 (P1_R1138_U26, P1_U3060);
  nand ginst1586 (P1_R1138_U260, P1_U3074, P1_U3497);
  not ginst1587 (P1_R1138_U261, P1_R1138_U93);
  or ginst1588 (P1_R1138_U262, P1_U3069, P1_U3503);
  or ginst1589 (P1_R1138_U263, P1_U3073, P1_U3500);
  not ginst1590 (P1_R1138_U264, P1_R1138_U60);
  nand ginst1591 (P1_R1138_U265, P1_R1138_U60, P1_R1138_U61);
  nand ginst1592 (P1_R1138_U266, P1_R1138_U265, P1_U3069);
  nand ginst1593 (P1_R1138_U267, P1_R1138_U264, P1_U3503);
  nand ginst1594 (P1_R1138_U268, P1_R1138_U9, P1_R1138_U93);
  not ginst1595 (P1_R1138_U269, P1_R1138_U161);
  not ginst1596 (P1_R1138_U27, P1_U3067);
  or ginst1597 (P1_R1138_U270, P1_U3076, P1_U3982);
  or ginst1598 (P1_R1138_U271, P1_U3081, P1_U3508);
  or ginst1599 (P1_R1138_U272, P1_U3075, P1_U3981);
  not ginst1600 (P1_R1138_U273, P1_R1138_U81);
  nand ginst1601 (P1_R1138_U274, P1_R1138_U273, P1_U3982);
  nand ginst1602 (P1_R1138_U275, P1_R1138_U274, P1_R1138_U91);
  nand ginst1603 (P1_R1138_U276, P1_R1138_U81, P1_R1138_U82);
  nand ginst1604 (P1_R1138_U277, P1_R1138_U275, P1_R1138_U276);
  nand ginst1605 (P1_R1138_U278, P1_R1138_U10, P1_R1138_U174);
  nand ginst1606 (P1_R1138_U279, P1_U3075, P1_U3981);
  not ginst1607 (P1_R1138_U28, P1_U3458);
  nand ginst1608 (P1_R1138_U280, P1_R1138_U277, P1_R1138_U278);
  or ginst1609 (P1_R1138_U281, P1_U3082, P1_U3506);
  or ginst1610 (P1_R1138_U282, P1_U3075, P1_U3981);
  nand ginst1611 (P1_R1138_U283, P1_R1138_U131, P1_R1138_U161, P1_R1138_U272);
  nand ginst1612 (P1_R1138_U284, P1_R1138_U280, P1_R1138_U282);
  not ginst1613 (P1_R1138_U285, P1_R1138_U158);
  or ginst1614 (P1_R1138_U286, P1_U3061, P1_U3980);
  nand ginst1615 (P1_R1138_U287, P1_R1138_U158, P1_R1138_U286);
  nand ginst1616 (P1_R1138_U288, P1_U3061, P1_U3980);
  not ginst1617 (P1_R1138_U289, P1_R1138_U156);
  not ginst1618 (P1_R1138_U29, P1_U3068);
  or ginst1619 (P1_R1138_U290, P1_U3066, P1_U3979);
  nand ginst1620 (P1_R1138_U291, P1_R1138_U156, P1_R1138_U290);
  nand ginst1621 (P1_R1138_U292, P1_U3066, P1_U3979);
  not ginst1622 (P1_R1138_U293, P1_R1138_U154);
  or ginst1623 (P1_R1138_U294, P1_U3058, P1_U3977);
  nand ginst1624 (P1_R1138_U295, P1_R1138_U172, P1_R1138_U175);
  not ginst1625 (P1_R1138_U296, P1_R1138_U87);
  or ginst1626 (P1_R1138_U297, P1_U3065, P1_U3978);
  nand ginst1627 (P1_R1138_U298, P1_R1138_U154, P1_R1138_U167, P1_R1138_U297);
  not ginst1628 (P1_R1138_U299, P1_R1138_U152);
  not ginst1629 (P1_R1138_U30, P1_U3450);
  or ginst1630 (P1_R1138_U300, P1_U3053, P1_U3975);
  nand ginst1631 (P1_R1138_U301, P1_U3053, P1_U3975);
  not ginst1632 (P1_R1138_U302, P1_R1138_U150);
  nand ginst1633 (P1_R1138_U303, P1_R1138_U150, P1_U3974);
  not ginst1634 (P1_R1138_U304, P1_R1138_U148);
  nand ginst1635 (P1_R1138_U305, P1_R1138_U154, P1_R1138_U297);
  not ginst1636 (P1_R1138_U306, P1_R1138_U90);
  or ginst1637 (P1_R1138_U307, P1_U3058, P1_U3977);
  nand ginst1638 (P1_R1138_U308, P1_R1138_U307, P1_R1138_U90);
  nand ginst1639 (P1_R1138_U309, P1_R1138_U153, P1_R1138_U172, P1_R1138_U308);
  not ginst1640 (P1_R1138_U31, P1_U3077);
  nand ginst1641 (P1_R1138_U310, P1_R1138_U172, P1_R1138_U306);
  nand ginst1642 (P1_R1138_U311, P1_U3057, P1_U3976);
  nand ginst1643 (P1_R1138_U312, P1_R1138_U167, P1_R1138_U310, P1_R1138_U311);
  or ginst1644 (P1_R1138_U313, P1_U3058, P1_U3977);
  nand ginst1645 (P1_R1138_U314, P1_R1138_U161, P1_R1138_U281);
  not ginst1646 (P1_R1138_U315, P1_R1138_U92);
  nand ginst1647 (P1_R1138_U316, P1_R1138_U10, P1_R1138_U92);
  nand ginst1648 (P1_R1138_U317, P1_R1138_U135, P1_R1138_U316);
  nand ginst1649 (P1_R1138_U318, P1_R1138_U277, P1_R1138_U316);
  nand ginst1650 (P1_R1138_U319, P1_R1138_U318, P1_R1138_U452);
  nand ginst1651 (P1_R1138_U32, P1_U3077, P1_U3450);
  or ginst1652 (P1_R1138_U320, P1_U3081, P1_U3508);
  nand ginst1653 (P1_R1138_U321, P1_R1138_U320, P1_R1138_U92);
  nand ginst1654 (P1_R1138_U322, P1_R1138_U136, P1_R1138_U321);
  nand ginst1655 (P1_R1138_U323, P1_R1138_U315, P1_R1138_U81);
  nand ginst1656 (P1_R1138_U324, P1_U3076, P1_U3982);
  nand ginst1657 (P1_R1138_U325, P1_R1138_U10, P1_R1138_U323, P1_R1138_U324);
  or ginst1658 (P1_R1138_U326, P1_U3078, P1_U3455);
  not ginst1659 (P1_R1138_U327, P1_R1138_U160);
  or ginst1660 (P1_R1138_U328, P1_U3081, P1_U3508);
  or ginst1661 (P1_R1138_U329, P1_U3073, P1_U3500);
  not ginst1662 (P1_R1138_U33, P1_U3461);
  nand ginst1663 (P1_R1138_U330, P1_R1138_U329, P1_R1138_U93);
  nand ginst1664 (P1_R1138_U331, P1_R1138_U137, P1_R1138_U330);
  nand ginst1665 (P1_R1138_U332, P1_R1138_U261, P1_R1138_U60);
  nand ginst1666 (P1_R1138_U333, P1_U3069, P1_U3503);
  nand ginst1667 (P1_R1138_U334, P1_R1138_U138, P1_R1138_U332);
  or ginst1668 (P1_R1138_U335, P1_U3073, P1_U3500);
  nand ginst1669 (P1_R1138_U336, P1_R1138_U166, P1_R1138_U249);
  not ginst1670 (P1_R1138_U337, P1_R1138_U94);
  or ginst1671 (P1_R1138_U338, P1_U3072, P1_U3488);
  nand ginst1672 (P1_R1138_U339, P1_R1138_U338, P1_R1138_U94);
  not ginst1673 (P1_R1138_U34, P1_U3064);
  nand ginst1674 (P1_R1138_U340, P1_R1138_U139, P1_R1138_U339);
  nand ginst1675 (P1_R1138_U341, P1_R1138_U171, P1_R1138_U337);
  nand ginst1676 (P1_R1138_U342, P1_U3080, P1_U3491);
  nand ginst1677 (P1_R1138_U343, P1_R1138_U140, P1_R1138_U341);
  or ginst1678 (P1_R1138_U344, P1_U3072, P1_U3488);
  or ginst1679 (P1_R1138_U345, P1_U3083, P1_U3479);
  nand ginst1680 (P1_R1138_U346, P1_R1138_U345, P1_R1138_U41);
  nand ginst1681 (P1_R1138_U347, P1_R1138_U141, P1_R1138_U346);
  nand ginst1682 (P1_R1138_U348, P1_R1138_U170, P1_R1138_U205);
  nand ginst1683 (P1_R1138_U349, P1_U3062, P1_U3482);
  nand ginst1684 (P1_R1138_U35, P1_U3060, P1_U3464);
  nand ginst1685 (P1_R1138_U350, P1_R1138_U142, P1_R1138_U348);
  nand ginst1686 (P1_R1138_U351, P1_R1138_U170, P1_R1138_U206);
  nand ginst1687 (P1_R1138_U352, P1_R1138_U203, P1_R1138_U62);
  nand ginst1688 (P1_R1138_U353, P1_R1138_U213, P1_R1138_U23);
  nand ginst1689 (P1_R1138_U354, P1_R1138_U227, P1_R1138_U35);
  nand ginst1690 (P1_R1138_U355, P1_R1138_U179, P1_R1138_U230);
  nand ginst1691 (P1_R1138_U356, P1_R1138_U172, P1_R1138_U313);
  nand ginst1692 (P1_R1138_U357, P1_R1138_U175, P1_R1138_U297);
  nand ginst1693 (P1_R1138_U358, P1_R1138_U328, P1_R1138_U81);
  nand ginst1694 (P1_R1138_U359, P1_R1138_U281, P1_R1138_U78);
  not ginst1695 (P1_R1138_U36, P1_U3467);
  nand ginst1696 (P1_R1138_U360, P1_R1138_U335, P1_R1138_U60);
  nand ginst1697 (P1_R1138_U361, P1_R1138_U171, P1_R1138_U344);
  nand ginst1698 (P1_R1138_U362, P1_R1138_U249, P1_R1138_U69);
  nand ginst1699 (P1_R1138_U363, P1_U3054, P1_U3974);
  nand ginst1700 (P1_R1138_U364, P1_R1138_U167, P1_R1138_U295);
  nand ginst1701 (P1_R1138_U365, P1_R1138_U294, P1_U3057);
  nand ginst1702 (P1_R1138_U366, P1_R1138_U294, P1_U3976);
  nand ginst1703 (P1_R1138_U367, P1_R1138_U167, P1_R1138_U295, P1_R1138_U300);
  nand ginst1704 (P1_R1138_U368, P1_R1138_U133, P1_R1138_U154, P1_R1138_U167);
  nand ginst1705 (P1_R1138_U369, P1_R1138_U296, P1_R1138_U300);
  not ginst1706 (P1_R1138_U37, P1_U3476);
  nand ginst1707 (P1_R1138_U370, P1_R1138_U40, P1_U3083);
  nand ginst1708 (P1_R1138_U371, P1_R1138_U39, P1_U3479);
  nand ginst1709 (P1_R1138_U372, P1_R1138_U370, P1_R1138_U371);
  nand ginst1710 (P1_R1138_U373, P1_R1138_U351, P1_R1138_U41);
  nand ginst1711 (P1_R1138_U374, P1_R1138_U205, P1_R1138_U372);
  nand ginst1712 (P1_R1138_U375, P1_R1138_U37, P1_U3084);
  nand ginst1713 (P1_R1138_U376, P1_R1138_U38, P1_U3476);
  nand ginst1714 (P1_R1138_U377, P1_R1138_U375, P1_R1138_U376);
  nand ginst1715 (P1_R1138_U378, P1_R1138_U143, P1_R1138_U352);
  nand ginst1716 (P1_R1138_U379, P1_R1138_U202, P1_R1138_U377);
  not ginst1717 (P1_R1138_U38, P1_U3084);
  nand ginst1718 (P1_R1138_U380, P1_R1138_U24, P1_U3070);
  nand ginst1719 (P1_R1138_U381, P1_R1138_U22, P1_U3473);
  nand ginst1720 (P1_R1138_U382, P1_R1138_U20, P1_U3071);
  nand ginst1721 (P1_R1138_U383, P1_R1138_U21, P1_U3470);
  nand ginst1722 (P1_R1138_U384, P1_R1138_U382, P1_R1138_U383);
  nand ginst1723 (P1_R1138_U385, P1_R1138_U353, P1_R1138_U42);
  nand ginst1724 (P1_R1138_U386, P1_R1138_U194, P1_R1138_U384);
  nand ginst1725 (P1_R1138_U387, P1_R1138_U36, P1_U3067);
  nand ginst1726 (P1_R1138_U388, P1_R1138_U27, P1_U3467);
  nand ginst1727 (P1_R1138_U389, P1_R1138_U25, P1_U3060);
  not ginst1728 (P1_R1138_U39, P1_U3083);
  nand ginst1729 (P1_R1138_U390, P1_R1138_U26, P1_U3464);
  nand ginst1730 (P1_R1138_U391, P1_R1138_U389, P1_R1138_U390);
  nand ginst1731 (P1_R1138_U392, P1_R1138_U354, P1_R1138_U45);
  nand ginst1732 (P1_R1138_U393, P1_R1138_U220, P1_R1138_U391);
  nand ginst1733 (P1_R1138_U394, P1_R1138_U33, P1_U3064);
  nand ginst1734 (P1_R1138_U395, P1_R1138_U34, P1_U3461);
  nand ginst1735 (P1_R1138_U396, P1_R1138_U394, P1_R1138_U395);
  nand ginst1736 (P1_R1138_U397, P1_R1138_U144, P1_R1138_U355);
  nand ginst1737 (P1_R1138_U398, P1_R1138_U229, P1_R1138_U396);
  nand ginst1738 (P1_R1138_U399, P1_R1138_U28, P1_U3068);
  and ginst1739 (P1_R1138_U4, P1_R1138_U177, P1_R1138_U178);
  not ginst1740 (P1_R1138_U40, P1_U3479);
  nand ginst1741 (P1_R1138_U400, P1_R1138_U29, P1_U3458);
  nand ginst1742 (P1_R1138_U401, P1_R1138_U146, P1_U3055);
  nand ginst1743 (P1_R1138_U402, P1_R1138_U145, P1_U3985);
  nand ginst1744 (P1_R1138_U403, P1_R1138_U146, P1_U3055);
  nand ginst1745 (P1_R1138_U404, P1_R1138_U145, P1_U3985);
  nand ginst1746 (P1_R1138_U405, P1_R1138_U403, P1_R1138_U404);
  nand ginst1747 (P1_R1138_U406, P1_R1138_U147, P1_R1138_U148);
  nand ginst1748 (P1_R1138_U407, P1_R1138_U304, P1_R1138_U405);
  nand ginst1749 (P1_R1138_U408, P1_R1138_U89, P1_U3054);
  nand ginst1750 (P1_R1138_U409, P1_R1138_U88, P1_U3974);
  nand ginst1751 (P1_R1138_U41, P1_R1138_U204, P1_R1138_U62);
  nand ginst1752 (P1_R1138_U410, P1_R1138_U89, P1_U3054);
  nand ginst1753 (P1_R1138_U411, P1_R1138_U88, P1_U3974);
  nand ginst1754 (P1_R1138_U412, P1_R1138_U410, P1_R1138_U411);
  nand ginst1755 (P1_R1138_U413, P1_R1138_U149, P1_R1138_U150);
  nand ginst1756 (P1_R1138_U414, P1_R1138_U302, P1_R1138_U412);
  nand ginst1757 (P1_R1138_U415, P1_R1138_U47, P1_U3053);
  nand ginst1758 (P1_R1138_U416, P1_R1138_U48, P1_U3975);
  nand ginst1759 (P1_R1138_U417, P1_R1138_U47, P1_U3053);
  nand ginst1760 (P1_R1138_U418, P1_R1138_U48, P1_U3975);
  nand ginst1761 (P1_R1138_U419, P1_R1138_U417, P1_R1138_U418);
  nand ginst1762 (P1_R1138_U42, P1_R1138_U118, P1_R1138_U192);
  nand ginst1763 (P1_R1138_U420, P1_R1138_U151, P1_R1138_U152);
  nand ginst1764 (P1_R1138_U421, P1_R1138_U299, P1_R1138_U419);
  nand ginst1765 (P1_R1138_U422, P1_R1138_U50, P1_U3057);
  nand ginst1766 (P1_R1138_U423, P1_R1138_U49, P1_U3976);
  nand ginst1767 (P1_R1138_U424, P1_R1138_U51, P1_U3058);
  nand ginst1768 (P1_R1138_U425, P1_R1138_U52, P1_U3977);
  nand ginst1769 (P1_R1138_U426, P1_R1138_U424, P1_R1138_U425);
  nand ginst1770 (P1_R1138_U427, P1_R1138_U356, P1_R1138_U90);
  nand ginst1771 (P1_R1138_U428, P1_R1138_U306, P1_R1138_U426);
  nand ginst1772 (P1_R1138_U429, P1_R1138_U53, P1_U3065);
  nand ginst1773 (P1_R1138_U43, P1_R1138_U181, P1_R1138_U182);
  nand ginst1774 (P1_R1138_U430, P1_R1138_U54, P1_U3978);
  nand ginst1775 (P1_R1138_U431, P1_R1138_U429, P1_R1138_U430);
  nand ginst1776 (P1_R1138_U432, P1_R1138_U154, P1_R1138_U357);
  nand ginst1777 (P1_R1138_U433, P1_R1138_U293, P1_R1138_U431);
  nand ginst1778 (P1_R1138_U434, P1_R1138_U85, P1_U3066);
  nand ginst1779 (P1_R1138_U435, P1_R1138_U86, P1_U3979);
  nand ginst1780 (P1_R1138_U436, P1_R1138_U85, P1_U3066);
  nand ginst1781 (P1_R1138_U437, P1_R1138_U86, P1_U3979);
  nand ginst1782 (P1_R1138_U438, P1_R1138_U436, P1_R1138_U437);
  nand ginst1783 (P1_R1138_U439, P1_R1138_U155, P1_R1138_U156);
  nand ginst1784 (P1_R1138_U44, P1_U3078, P1_U3455);
  nand ginst1785 (P1_R1138_U440, P1_R1138_U289, P1_R1138_U438);
  nand ginst1786 (P1_R1138_U441, P1_R1138_U83, P1_U3061);
  nand ginst1787 (P1_R1138_U442, P1_R1138_U84, P1_U3980);
  nand ginst1788 (P1_R1138_U443, P1_R1138_U83, P1_U3061);
  nand ginst1789 (P1_R1138_U444, P1_R1138_U84, P1_U3980);
  nand ginst1790 (P1_R1138_U445, P1_R1138_U443, P1_R1138_U444);
  nand ginst1791 (P1_R1138_U446, P1_R1138_U157, P1_R1138_U158);
  nand ginst1792 (P1_R1138_U447, P1_R1138_U285, P1_R1138_U445);
  nand ginst1793 (P1_R1138_U448, P1_R1138_U55, P1_U3075);
  nand ginst1794 (P1_R1138_U449, P1_R1138_U56, P1_U3981);
  nand ginst1795 (P1_R1138_U45, P1_R1138_U122, P1_R1138_U218);
  nand ginst1796 (P1_R1138_U450, P1_R1138_U55, P1_U3075);
  nand ginst1797 (P1_R1138_U451, P1_R1138_U56, P1_U3981);
  nand ginst1798 (P1_R1138_U452, P1_R1138_U450, P1_R1138_U451);
  nand ginst1799 (P1_R1138_U453, P1_R1138_U82, P1_U3076);
  nand ginst1800 (P1_R1138_U454, P1_R1138_U91, P1_U3982);
  nand ginst1801 (P1_R1138_U455, P1_R1138_U160, P1_R1138_U181);
  nand ginst1802 (P1_R1138_U456, P1_R1138_U32, P1_R1138_U327);
  nand ginst1803 (P1_R1138_U457, P1_R1138_U79, P1_U3081);
  nand ginst1804 (P1_R1138_U458, P1_R1138_U80, P1_U3508);
  nand ginst1805 (P1_R1138_U459, P1_R1138_U457, P1_R1138_U458);
  nand ginst1806 (P1_R1138_U46, P1_R1138_U214, P1_R1138_U215);
  nand ginst1807 (P1_R1138_U460, P1_R1138_U358, P1_R1138_U92);
  nand ginst1808 (P1_R1138_U461, P1_R1138_U315, P1_R1138_U459);
  nand ginst1809 (P1_R1138_U462, P1_R1138_U76, P1_U3082);
  nand ginst1810 (P1_R1138_U463, P1_R1138_U77, P1_U3506);
  nand ginst1811 (P1_R1138_U464, P1_R1138_U462, P1_R1138_U463);
  nand ginst1812 (P1_R1138_U465, P1_R1138_U161, P1_R1138_U359);
  nand ginst1813 (P1_R1138_U466, P1_R1138_U269, P1_R1138_U464);
  nand ginst1814 (P1_R1138_U467, P1_R1138_U61, P1_U3069);
  nand ginst1815 (P1_R1138_U468, P1_R1138_U59, P1_U3503);
  nand ginst1816 (P1_R1138_U469, P1_R1138_U57, P1_U3073);
  not ginst1817 (P1_R1138_U47, P1_U3975);
  nand ginst1818 (P1_R1138_U470, P1_R1138_U58, P1_U3500);
  nand ginst1819 (P1_R1138_U471, P1_R1138_U469, P1_R1138_U470);
  nand ginst1820 (P1_R1138_U472, P1_R1138_U360, P1_R1138_U93);
  nand ginst1821 (P1_R1138_U473, P1_R1138_U261, P1_R1138_U471);
  nand ginst1822 (P1_R1138_U474, P1_R1138_U74, P1_U3074);
  nand ginst1823 (P1_R1138_U475, P1_R1138_U75, P1_U3497);
  nand ginst1824 (P1_R1138_U476, P1_R1138_U74, P1_U3074);
  nand ginst1825 (P1_R1138_U477, P1_R1138_U75, P1_U3497);
  nand ginst1826 (P1_R1138_U478, P1_R1138_U476, P1_R1138_U477);
  nand ginst1827 (P1_R1138_U479, P1_R1138_U162, P1_R1138_U163);
  not ginst1828 (P1_R1138_U48, P1_U3053);
  nand ginst1829 (P1_R1138_U480, P1_R1138_U257, P1_R1138_U478);
  nand ginst1830 (P1_R1138_U481, P1_R1138_U72, P1_U3079);
  nand ginst1831 (P1_R1138_U482, P1_R1138_U73, P1_U3494);
  nand ginst1832 (P1_R1138_U483, P1_R1138_U72, P1_U3079);
  nand ginst1833 (P1_R1138_U484, P1_R1138_U73, P1_U3494);
  nand ginst1834 (P1_R1138_U485, P1_R1138_U483, P1_R1138_U484);
  nand ginst1835 (P1_R1138_U486, P1_R1138_U164, P1_R1138_U165);
  nand ginst1836 (P1_R1138_U487, P1_R1138_U253, P1_R1138_U485);
  nand ginst1837 (P1_R1138_U488, P1_R1138_U70, P1_U3080);
  nand ginst1838 (P1_R1138_U489, P1_R1138_U71, P1_U3491);
  not ginst1839 (P1_R1138_U49, P1_U3057);
  nand ginst1840 (P1_R1138_U490, P1_R1138_U65, P1_U3072);
  nand ginst1841 (P1_R1138_U491, P1_R1138_U66, P1_U3488);
  nand ginst1842 (P1_R1138_U492, P1_R1138_U490, P1_R1138_U491);
  nand ginst1843 (P1_R1138_U493, P1_R1138_U361, P1_R1138_U94);
  nand ginst1844 (P1_R1138_U494, P1_R1138_U337, P1_R1138_U492);
  nand ginst1845 (P1_R1138_U495, P1_R1138_U67, P1_U3063);
  nand ginst1846 (P1_R1138_U496, P1_R1138_U68, P1_U3485);
  nand ginst1847 (P1_R1138_U497, P1_R1138_U495, P1_R1138_U496);
  nand ginst1848 (P1_R1138_U498, P1_R1138_U166, P1_R1138_U362);
  nand ginst1849 (P1_R1138_U499, P1_R1138_U243, P1_R1138_U497);
  and ginst1850 (P1_R1138_U5, P1_R1138_U179, P1_R1138_U180);
  not ginst1851 (P1_R1138_U50, P1_U3976);
  nand ginst1852 (P1_R1138_U500, P1_R1138_U63, P1_U3062);
  nand ginst1853 (P1_R1138_U501, P1_R1138_U64, P1_U3482);
  nand ginst1854 (P1_R1138_U502, P1_R1138_U30, P1_U3077);
  nand ginst1855 (P1_R1138_U503, P1_R1138_U31, P1_U3450);
  not ginst1856 (P1_R1138_U51, P1_U3977);
  not ginst1857 (P1_R1138_U52, P1_U3058);
  not ginst1858 (P1_R1138_U53, P1_U3978);
  not ginst1859 (P1_R1138_U54, P1_U3065);
  not ginst1860 (P1_R1138_U55, P1_U3981);
  not ginst1861 (P1_R1138_U56, P1_U3075);
  not ginst1862 (P1_R1138_U57, P1_U3500);
  not ginst1863 (P1_R1138_U58, P1_U3073);
  not ginst1864 (P1_R1138_U59, P1_U3069);
  and ginst1865 (P1_R1138_U6, P1_R1138_U195, P1_R1138_U196);
  nand ginst1866 (P1_R1138_U60, P1_U3073, P1_U3500);
  not ginst1867 (P1_R1138_U61, P1_U3503);
  nand ginst1868 (P1_R1138_U62, P1_U3084, P1_U3476);
  not ginst1869 (P1_R1138_U63, P1_U3482);
  not ginst1870 (P1_R1138_U64, P1_U3062);
  not ginst1871 (P1_R1138_U65, P1_U3488);
  not ginst1872 (P1_R1138_U66, P1_U3072);
  not ginst1873 (P1_R1138_U67, P1_U3485);
  not ginst1874 (P1_R1138_U68, P1_U3063);
  nand ginst1875 (P1_R1138_U69, P1_U3063, P1_U3485);
  and ginst1876 (P1_R1138_U7, P1_R1138_U235, P1_R1138_U236);
  not ginst1877 (P1_R1138_U70, P1_U3491);
  not ginst1878 (P1_R1138_U71, P1_U3080);
  not ginst1879 (P1_R1138_U72, P1_U3494);
  not ginst1880 (P1_R1138_U73, P1_U3079);
  not ginst1881 (P1_R1138_U74, P1_U3497);
  not ginst1882 (P1_R1138_U75, P1_U3074);
  not ginst1883 (P1_R1138_U76, P1_U3506);
  not ginst1884 (P1_R1138_U77, P1_U3082);
  nand ginst1885 (P1_R1138_U78, P1_U3082, P1_U3506);
  not ginst1886 (P1_R1138_U79, P1_U3508);
  and ginst1887 (P1_R1138_U8, P1_R1138_U244, P1_R1138_U245);
  not ginst1888 (P1_R1138_U80, P1_U3081);
  nand ginst1889 (P1_R1138_U81, P1_U3081, P1_U3508);
  not ginst1890 (P1_R1138_U82, P1_U3982);
  not ginst1891 (P1_R1138_U83, P1_U3980);
  not ginst1892 (P1_R1138_U84, P1_U3061);
  not ginst1893 (P1_R1138_U85, P1_U3979);
  not ginst1894 (P1_R1138_U86, P1_U3066);
  nand ginst1895 (P1_R1138_U87, P1_U3057, P1_U3976);
  not ginst1896 (P1_R1138_U88, P1_U3054);
  not ginst1897 (P1_R1138_U89, P1_U3974);
  and ginst1898 (P1_R1138_U9, P1_R1138_U262, P1_R1138_U263);
  nand ginst1899 (P1_R1138_U90, P1_R1138_U175, P1_R1138_U305);
  not ginst1900 (P1_R1138_U91, P1_U3076);
  nand ginst1901 (P1_R1138_U92, P1_R1138_U314, P1_R1138_U78);
  nand ginst1902 (P1_R1138_U93, P1_R1138_U259, P1_R1138_U260);
  nand ginst1903 (P1_R1138_U94, P1_R1138_U336, P1_R1138_U69);
  nand ginst1904 (P1_R1138_U95, P1_R1138_U455, P1_R1138_U456);
  nand ginst1905 (P1_R1138_U96, P1_R1138_U502, P1_R1138_U503);
  nand ginst1906 (P1_R1138_U97, P1_R1138_U373, P1_R1138_U374);
  nand ginst1907 (P1_R1138_U98, P1_R1138_U378, P1_R1138_U379);
  nand ginst1908 (P1_R1138_U99, P1_R1138_U385, P1_R1138_U386);
  nand ginst1909 (P1_R1150_U10, P1_R1150_U340, P1_R1150_U343);
  nand ginst1910 (P1_R1150_U100, P1_R1150_U460, P1_R1150_U461);
  nand ginst1911 (P1_R1150_U101, P1_R1150_U465, P1_R1150_U466);
  nand ginst1912 (P1_R1150_U102, P1_R1150_U350, P1_R1150_U351);
  nand ginst1913 (P1_R1150_U103, P1_R1150_U359, P1_R1150_U360);
  nand ginst1914 (P1_R1150_U104, P1_R1150_U366, P1_R1150_U367);
  nand ginst1915 (P1_R1150_U105, P1_R1150_U370, P1_R1150_U371);
  nand ginst1916 (P1_R1150_U106, P1_R1150_U379, P1_R1150_U380);
  nand ginst1917 (P1_R1150_U107, P1_R1150_U398, P1_R1150_U399);
  nand ginst1918 (P1_R1150_U108, P1_R1150_U415, P1_R1150_U416);
  nand ginst1919 (P1_R1150_U109, P1_R1150_U419, P1_R1150_U420);
  nand ginst1920 (P1_R1150_U11, P1_R1150_U329, P1_R1150_U332);
  nand ginst1921 (P1_R1150_U110, P1_R1150_U451, P1_R1150_U452);
  nand ginst1922 (P1_R1150_U111, P1_R1150_U455, P1_R1150_U456);
  nand ginst1923 (P1_R1150_U112, P1_R1150_U472, P1_R1150_U473);
  and ginst1924 (P1_R1150_U113, P1_R1150_U193, P1_R1150_U194);
  and ginst1925 (P1_R1150_U114, P1_R1150_U196, P1_R1150_U201);
  and ginst1926 (P1_R1150_U115, P1_R1150_U180, P1_R1150_U206);
  and ginst1927 (P1_R1150_U116, P1_R1150_U209, P1_R1150_U210);
  and ginst1928 (P1_R1150_U117, P1_R1150_U352, P1_R1150_U353, P1_R1150_U37);
  and ginst1929 (P1_R1150_U118, P1_R1150_U180, P1_R1150_U356);
  and ginst1930 (P1_R1150_U119, P1_R1150_U225, P1_R1150_U6);
  nand ginst1931 (P1_R1150_U12, P1_R1150_U318, P1_R1150_U321);
  and ginst1932 (P1_R1150_U120, P1_R1150_U179, P1_R1150_U363);
  and ginst1933 (P1_R1150_U121, P1_R1150_U27, P1_R1150_U372, P1_R1150_U373);
  and ginst1934 (P1_R1150_U122, P1_R1150_U178, P1_R1150_U376);
  and ginst1935 (P1_R1150_U123, P1_R1150_U174, P1_R1150_U212, P1_R1150_U235);
  and ginst1936 (P1_R1150_U124, P1_R1150_U175, P1_R1150_U252, P1_R1150_U257);
  and ginst1937 (P1_R1150_U125, P1_R1150_U176, P1_R1150_U283);
  and ginst1938 (P1_R1150_U126, P1_R1150_U299, P1_R1150_U300);
  nand ginst1939 (P1_R1150_U127, P1_R1150_U386, P1_R1150_U387);
  and ginst1940 (P1_R1150_U128, P1_R1150_U391, P1_R1150_U392, P1_R1150_U82);
  and ginst1941 (P1_R1150_U129, P1_R1150_U177, P1_R1150_U395);
  nand ginst1942 (P1_R1150_U13, P1_R1150_U310, P1_R1150_U312);
  nand ginst1943 (P1_R1150_U130, P1_R1150_U400, P1_R1150_U401);
  nand ginst1944 (P1_R1150_U131, P1_R1150_U405, P1_R1150_U406);
  and ginst1945 (P1_R1150_U132, P1_R1150_U176, P1_R1150_U412);
  nand ginst1946 (P1_R1150_U133, P1_R1150_U421, P1_R1150_U422);
  nand ginst1947 (P1_R1150_U134, P1_R1150_U426, P1_R1150_U427);
  nand ginst1948 (P1_R1150_U135, P1_R1150_U431, P1_R1150_U432);
  nand ginst1949 (P1_R1150_U136, P1_R1150_U436, P1_R1150_U437);
  nand ginst1950 (P1_R1150_U137, P1_R1150_U441, P1_R1150_U442);
  and ginst1951 (P1_R1150_U138, P1_R1150_U331, P1_R1150_U8);
  and ginst1952 (P1_R1150_U139, P1_R1150_U175, P1_R1150_U448);
  nand ginst1953 (P1_R1150_U14, P1_R1150_U308, P1_R1150_U347);
  nand ginst1954 (P1_R1150_U140, P1_R1150_U457, P1_R1150_U458);
  nand ginst1955 (P1_R1150_U141, P1_R1150_U462, P1_R1150_U463);
  and ginst1956 (P1_R1150_U142, P1_R1150_U342, P1_R1150_U7);
  and ginst1957 (P1_R1150_U143, P1_R1150_U174, P1_R1150_U469);
  and ginst1958 (P1_R1150_U144, P1_R1150_U348, P1_R1150_U349);
  nand ginst1959 (P1_R1150_U145, P1_R1150_U116, P1_R1150_U207);
  and ginst1960 (P1_R1150_U146, P1_R1150_U357, P1_R1150_U358);
  and ginst1961 (P1_R1150_U147, P1_R1150_U364, P1_R1150_U365);
  and ginst1962 (P1_R1150_U148, P1_R1150_U368, P1_R1150_U369);
  nand ginst1963 (P1_R1150_U149, P1_R1150_U113, P1_R1150_U191);
  nand ginst1964 (P1_R1150_U15, P1_R1150_U231, P1_R1150_U233);
  and ginst1965 (P1_R1150_U150, P1_R1150_U377, P1_R1150_U378);
  not ginst1966 (P1_R1150_U151, P1_U3985);
  not ginst1967 (P1_R1150_U152, P1_U3055);
  and ginst1968 (P1_R1150_U153, P1_R1150_U381, P1_R1150_U382);
  and ginst1969 (P1_R1150_U154, P1_R1150_U396, P1_R1150_U397);
  nand ginst1970 (P1_R1150_U155, P1_R1150_U289, P1_R1150_U290);
  nand ginst1971 (P1_R1150_U156, P1_R1150_U285, P1_R1150_U286);
  and ginst1972 (P1_R1150_U157, P1_R1150_U413, P1_R1150_U414);
  and ginst1973 (P1_R1150_U158, P1_R1150_U417, P1_R1150_U418);
  nand ginst1974 (P1_R1150_U159, P1_R1150_U275, P1_R1150_U276);
  nand ginst1975 (P1_R1150_U16, P1_R1150_U223, P1_R1150_U226);
  nand ginst1976 (P1_R1150_U160, P1_R1150_U271, P1_R1150_U272);
  not ginst1977 (P1_R1150_U161, P1_U3455);
  nand ginst1978 (P1_R1150_U162, P1_R1150_U267, P1_R1150_U268);
  not ginst1979 (P1_R1150_U163, P1_U3506);
  nand ginst1980 (P1_R1150_U164, P1_R1150_U259, P1_R1150_U260);
  and ginst1981 (P1_R1150_U165, P1_R1150_U449, P1_R1150_U450);
  and ginst1982 (P1_R1150_U166, P1_R1150_U453, P1_R1150_U454);
  nand ginst1983 (P1_R1150_U167, P1_R1150_U249, P1_R1150_U250);
  nand ginst1984 (P1_R1150_U168, P1_R1150_U245, P1_R1150_U246);
  nand ginst1985 (P1_R1150_U169, P1_R1150_U241, P1_R1150_U242);
  nand ginst1986 (P1_R1150_U17, P1_R1150_U215, P1_R1150_U217);
  and ginst1987 (P1_R1150_U170, P1_R1150_U470, P1_R1150_U471);
  not ginst1988 (P1_R1150_U171, P1_R1150_U82);
  not ginst1989 (P1_R1150_U172, P1_R1150_U27);
  not ginst1990 (P1_R1150_U173, P1_R1150_U37);
  nand ginst1991 (P1_R1150_U174, P1_R1150_U50, P1_U3482);
  nand ginst1992 (P1_R1150_U175, P1_R1150_U59, P1_U3497);
  nand ginst1993 (P1_R1150_U176, P1_R1150_U73, P1_U3980);
  nand ginst1994 (P1_R1150_U177, P1_R1150_U81, P1_U3976);
  nand ginst1995 (P1_R1150_U178, P1_R1150_U26, P1_U3458);
  nand ginst1996 (P1_R1150_U179, P1_R1150_U32, P1_U3467);
  nand ginst1997 (P1_R1150_U18, P1_R1150_U23, P1_R1150_U346);
  nand ginst1998 (P1_R1150_U180, P1_R1150_U36, P1_U3473);
  not ginst1999 (P1_R1150_U181, P1_R1150_U61);
  not ginst2000 (P1_R1150_U182, P1_R1150_U75);
  not ginst2001 (P1_R1150_U183, P1_R1150_U34);
  not ginst2002 (P1_R1150_U184, P1_R1150_U51);
  not ginst2003 (P1_R1150_U185, P1_R1150_U23);
  nand ginst2004 (P1_R1150_U186, P1_R1150_U185, P1_R1150_U24);
  nand ginst2005 (P1_R1150_U187, P1_R1150_U161, P1_R1150_U186);
  nand ginst2006 (P1_R1150_U188, P1_R1150_U23, P1_U3078);
  not ginst2007 (P1_R1150_U189, P1_R1150_U43);
  not ginst2008 (P1_R1150_U19, P1_U3473);
  nand ginst2009 (P1_R1150_U190, P1_R1150_U28, P1_U3461);
  nand ginst2010 (P1_R1150_U191, P1_R1150_U178, P1_R1150_U190, P1_R1150_U43);
  nand ginst2011 (P1_R1150_U192, P1_R1150_U27, P1_R1150_U28);
  nand ginst2012 (P1_R1150_U193, P1_R1150_U192, P1_R1150_U25);
  nand ginst2013 (P1_R1150_U194, P1_R1150_U172, P1_U3064);
  not ginst2014 (P1_R1150_U195, P1_R1150_U149);
  nand ginst2015 (P1_R1150_U196, P1_R1150_U31, P1_U3470);
  nand ginst2016 (P1_R1150_U197, P1_R1150_U29, P1_U3071);
  nand ginst2017 (P1_R1150_U198, P1_R1150_U20, P1_U3067);
  nand ginst2018 (P1_R1150_U199, P1_R1150_U179, P1_R1150_U183);
  not ginst2019 (P1_R1150_U20, P1_U3467);
  nand ginst2020 (P1_R1150_U200, P1_R1150_U199, P1_R1150_U6);
  nand ginst2021 (P1_R1150_U201, P1_R1150_U33, P1_U3464);
  nand ginst2022 (P1_R1150_U202, P1_R1150_U31, P1_U3470);
  nand ginst2023 (P1_R1150_U203, P1_R1150_U114, P1_R1150_U149, P1_R1150_U179);
  nand ginst2024 (P1_R1150_U204, P1_R1150_U200, P1_R1150_U202);
  not ginst2025 (P1_R1150_U205, P1_R1150_U41);
  nand ginst2026 (P1_R1150_U206, P1_R1150_U38, P1_U3476);
  nand ginst2027 (P1_R1150_U207, P1_R1150_U115, P1_R1150_U41);
  nand ginst2028 (P1_R1150_U208, P1_R1150_U37, P1_R1150_U38);
  nand ginst2029 (P1_R1150_U209, P1_R1150_U208, P1_R1150_U35);
  not ginst2030 (P1_R1150_U21, P1_U3458);
  nand ginst2031 (P1_R1150_U210, P1_R1150_U173, P1_U3084);
  not ginst2032 (P1_R1150_U211, P1_R1150_U145);
  nand ginst2033 (P1_R1150_U212, P1_R1150_U40, P1_U3479);
  nand ginst2034 (P1_R1150_U213, P1_R1150_U212, P1_R1150_U51);
  nand ginst2035 (P1_R1150_U214, P1_R1150_U205, P1_R1150_U37);
  nand ginst2036 (P1_R1150_U215, P1_R1150_U118, P1_R1150_U214);
  nand ginst2037 (P1_R1150_U216, P1_R1150_U180, P1_R1150_U41);
  nand ginst2038 (P1_R1150_U217, P1_R1150_U117, P1_R1150_U216);
  nand ginst2039 (P1_R1150_U218, P1_R1150_U180, P1_R1150_U37);
  nand ginst2040 (P1_R1150_U219, P1_R1150_U149, P1_R1150_U201);
  not ginst2041 (P1_R1150_U22, P1_U3450);
  not ginst2042 (P1_R1150_U220, P1_R1150_U42);
  nand ginst2043 (P1_R1150_U221, P1_R1150_U20, P1_U3067);
  nand ginst2044 (P1_R1150_U222, P1_R1150_U220, P1_R1150_U221);
  nand ginst2045 (P1_R1150_U223, P1_R1150_U120, P1_R1150_U222);
  nand ginst2046 (P1_R1150_U224, P1_R1150_U179, P1_R1150_U42);
  nand ginst2047 (P1_R1150_U225, P1_R1150_U31, P1_U3470);
  nand ginst2048 (P1_R1150_U226, P1_R1150_U119, P1_R1150_U224);
  nand ginst2049 (P1_R1150_U227, P1_R1150_U20, P1_U3067);
  nand ginst2050 (P1_R1150_U228, P1_R1150_U179, P1_R1150_U227);
  nand ginst2051 (P1_R1150_U229, P1_R1150_U201, P1_R1150_U34);
  nand ginst2052 (P1_R1150_U23, P1_R1150_U91, P1_U3450);
  nand ginst2053 (P1_R1150_U230, P1_R1150_U189, P1_R1150_U27);
  nand ginst2054 (P1_R1150_U231, P1_R1150_U122, P1_R1150_U230);
  nand ginst2055 (P1_R1150_U232, P1_R1150_U178, P1_R1150_U43);
  nand ginst2056 (P1_R1150_U233, P1_R1150_U121, P1_R1150_U232);
  nand ginst2057 (P1_R1150_U234, P1_R1150_U178, P1_R1150_U27);
  nand ginst2058 (P1_R1150_U235, P1_R1150_U49, P1_U3485);
  nand ginst2059 (P1_R1150_U236, P1_R1150_U48, P1_U3063);
  nand ginst2060 (P1_R1150_U237, P1_R1150_U47, P1_U3062);
  nand ginst2061 (P1_R1150_U238, P1_R1150_U174, P1_R1150_U184);
  nand ginst2062 (P1_R1150_U239, P1_R1150_U238, P1_R1150_U7);
  not ginst2063 (P1_R1150_U24, P1_U3078);
  nand ginst2064 (P1_R1150_U240, P1_R1150_U49, P1_U3485);
  nand ginst2065 (P1_R1150_U241, P1_R1150_U123, P1_R1150_U145);
  nand ginst2066 (P1_R1150_U242, P1_R1150_U239, P1_R1150_U240);
  not ginst2067 (P1_R1150_U243, P1_R1150_U169);
  nand ginst2068 (P1_R1150_U244, P1_R1150_U53, P1_U3488);
  nand ginst2069 (P1_R1150_U245, P1_R1150_U169, P1_R1150_U244);
  nand ginst2070 (P1_R1150_U246, P1_R1150_U52, P1_U3072);
  not ginst2071 (P1_R1150_U247, P1_R1150_U168);
  nand ginst2072 (P1_R1150_U248, P1_R1150_U55, P1_U3491);
  nand ginst2073 (P1_R1150_U249, P1_R1150_U168, P1_R1150_U248);
  not ginst2074 (P1_R1150_U25, P1_U3461);
  nand ginst2075 (P1_R1150_U250, P1_R1150_U54, P1_U3080);
  not ginst2076 (P1_R1150_U251, P1_R1150_U167);
  nand ginst2077 (P1_R1150_U252, P1_R1150_U58, P1_U3500);
  nand ginst2078 (P1_R1150_U253, P1_R1150_U56, P1_U3073);
  nand ginst2079 (P1_R1150_U254, P1_R1150_U46, P1_U3074);
  nand ginst2080 (P1_R1150_U255, P1_R1150_U175, P1_R1150_U181);
  nand ginst2081 (P1_R1150_U256, P1_R1150_U255, P1_R1150_U8);
  nand ginst2082 (P1_R1150_U257, P1_R1150_U60, P1_U3494);
  nand ginst2083 (P1_R1150_U258, P1_R1150_U58, P1_U3500);
  nand ginst2084 (P1_R1150_U259, P1_R1150_U124, P1_R1150_U167);
  not ginst2085 (P1_R1150_U26, P1_U3068);
  nand ginst2086 (P1_R1150_U260, P1_R1150_U256, P1_R1150_U258);
  not ginst2087 (P1_R1150_U261, P1_R1150_U164);
  nand ginst2088 (P1_R1150_U262, P1_R1150_U63, P1_U3503);
  nand ginst2089 (P1_R1150_U263, P1_R1150_U164, P1_R1150_U262);
  nand ginst2090 (P1_R1150_U264, P1_R1150_U62, P1_U3069);
  not ginst2091 (P1_R1150_U265, P1_R1150_U64);
  nand ginst2092 (P1_R1150_U266, P1_R1150_U265, P1_R1150_U65);
  nand ginst2093 (P1_R1150_U267, P1_R1150_U163, P1_R1150_U266);
  nand ginst2094 (P1_R1150_U268, P1_R1150_U64, P1_U3082);
  not ginst2095 (P1_R1150_U269, P1_R1150_U162);
  nand ginst2096 (P1_R1150_U27, P1_R1150_U21, P1_U3068);
  nand ginst2097 (P1_R1150_U270, P1_R1150_U67, P1_U3508);
  nand ginst2098 (P1_R1150_U271, P1_R1150_U162, P1_R1150_U270);
  nand ginst2099 (P1_R1150_U272, P1_R1150_U66, P1_U3081);
  not ginst2100 (P1_R1150_U273, P1_R1150_U160);
  nand ginst2101 (P1_R1150_U274, P1_R1150_U69, P1_U3982);
  nand ginst2102 (P1_R1150_U275, P1_R1150_U160, P1_R1150_U274);
  nand ginst2103 (P1_R1150_U276, P1_R1150_U68, P1_U3076);
  not ginst2104 (P1_R1150_U277, P1_R1150_U159);
  nand ginst2105 (P1_R1150_U278, P1_R1150_U72, P1_U3979);
  nand ginst2106 (P1_R1150_U279, P1_R1150_U70, P1_U3066);
  not ginst2107 (P1_R1150_U28, P1_U3064);
  nand ginst2108 (P1_R1150_U280, P1_R1150_U45, P1_U3061);
  nand ginst2109 (P1_R1150_U281, P1_R1150_U176, P1_R1150_U182);
  nand ginst2110 (P1_R1150_U282, P1_R1150_U281, P1_R1150_U9);
  nand ginst2111 (P1_R1150_U283, P1_R1150_U74, P1_U3981);
  nand ginst2112 (P1_R1150_U284, P1_R1150_U72, P1_U3979);
  nand ginst2113 (P1_R1150_U285, P1_R1150_U125, P1_R1150_U159, P1_R1150_U278);
  nand ginst2114 (P1_R1150_U286, P1_R1150_U282, P1_R1150_U284);
  not ginst2115 (P1_R1150_U287, P1_R1150_U156);
  nand ginst2116 (P1_R1150_U288, P1_R1150_U77, P1_U3978);
  nand ginst2117 (P1_R1150_U289, P1_R1150_U156, P1_R1150_U288);
  not ginst2118 (P1_R1150_U29, P1_U3470);
  nand ginst2119 (P1_R1150_U290, P1_R1150_U76, P1_U3065);
  not ginst2120 (P1_R1150_U291, P1_R1150_U155);
  nand ginst2121 (P1_R1150_U292, P1_R1150_U79, P1_U3977);
  nand ginst2122 (P1_R1150_U293, P1_R1150_U155, P1_R1150_U292);
  nand ginst2123 (P1_R1150_U294, P1_R1150_U78, P1_U3058);
  not ginst2124 (P1_R1150_U295, P1_R1150_U87);
  nand ginst2125 (P1_R1150_U296, P1_R1150_U83, P1_U3975);
  nand ginst2126 (P1_R1150_U297, P1_R1150_U177, P1_R1150_U296, P1_R1150_U87);
  nand ginst2127 (P1_R1150_U298, P1_R1150_U82, P1_R1150_U83);
  nand ginst2128 (P1_R1150_U299, P1_R1150_U298, P1_R1150_U80);
  not ginst2129 (P1_R1150_U30, P1_U3464);
  nand ginst2130 (P1_R1150_U300, P1_R1150_U171, P1_U3053);
  not ginst2131 (P1_R1150_U301, P1_R1150_U86);
  nand ginst2132 (P1_R1150_U302, P1_R1150_U84, P1_U3054);
  nand ginst2133 (P1_R1150_U303, P1_R1150_U301, P1_R1150_U302);
  nand ginst2134 (P1_R1150_U304, P1_R1150_U85, P1_U3974);
  nand ginst2135 (P1_R1150_U305, P1_R1150_U85, P1_U3974);
  nand ginst2136 (P1_R1150_U306, P1_R1150_U305, P1_R1150_U86);
  nand ginst2137 (P1_R1150_U307, P1_R1150_U84, P1_U3054);
  nand ginst2138 (P1_R1150_U308, P1_R1150_U153, P1_R1150_U306, P1_R1150_U307);
  nand ginst2139 (P1_R1150_U309, P1_R1150_U295, P1_R1150_U82);
  not ginst2140 (P1_R1150_U31, P1_U3071);
  nand ginst2141 (P1_R1150_U310, P1_R1150_U129, P1_R1150_U309);
  nand ginst2142 (P1_R1150_U311, P1_R1150_U177, P1_R1150_U87);
  nand ginst2143 (P1_R1150_U312, P1_R1150_U128, P1_R1150_U311);
  nand ginst2144 (P1_R1150_U313, P1_R1150_U177, P1_R1150_U82);
  nand ginst2145 (P1_R1150_U314, P1_R1150_U159, P1_R1150_U283);
  not ginst2146 (P1_R1150_U315, P1_R1150_U88);
  nand ginst2147 (P1_R1150_U316, P1_R1150_U45, P1_U3061);
  nand ginst2148 (P1_R1150_U317, P1_R1150_U315, P1_R1150_U316);
  nand ginst2149 (P1_R1150_U318, P1_R1150_U132, P1_R1150_U317);
  nand ginst2150 (P1_R1150_U319, P1_R1150_U176, P1_R1150_U88);
  not ginst2151 (P1_R1150_U32, P1_U3067);
  nand ginst2152 (P1_R1150_U320, P1_R1150_U72, P1_U3979);
  nand ginst2153 (P1_R1150_U321, P1_R1150_U319, P1_R1150_U320, P1_R1150_U9);
  nand ginst2154 (P1_R1150_U322, P1_R1150_U45, P1_U3061);
  nand ginst2155 (P1_R1150_U323, P1_R1150_U176, P1_R1150_U322);
  nand ginst2156 (P1_R1150_U324, P1_R1150_U283, P1_R1150_U75);
  nand ginst2157 (P1_R1150_U325, P1_R1150_U167, P1_R1150_U257);
  not ginst2158 (P1_R1150_U326, P1_R1150_U89);
  nand ginst2159 (P1_R1150_U327, P1_R1150_U46, P1_U3074);
  nand ginst2160 (P1_R1150_U328, P1_R1150_U326, P1_R1150_U327);
  nand ginst2161 (P1_R1150_U329, P1_R1150_U139, P1_R1150_U328);
  not ginst2162 (P1_R1150_U33, P1_U3060);
  nand ginst2163 (P1_R1150_U330, P1_R1150_U175, P1_R1150_U89);
  nand ginst2164 (P1_R1150_U331, P1_R1150_U58, P1_U3500);
  nand ginst2165 (P1_R1150_U332, P1_R1150_U138, P1_R1150_U330);
  nand ginst2166 (P1_R1150_U333, P1_R1150_U46, P1_U3074);
  nand ginst2167 (P1_R1150_U334, P1_R1150_U175, P1_R1150_U333);
  nand ginst2168 (P1_R1150_U335, P1_R1150_U257, P1_R1150_U61);
  nand ginst2169 (P1_R1150_U336, P1_R1150_U145, P1_R1150_U212);
  not ginst2170 (P1_R1150_U337, P1_R1150_U90);
  nand ginst2171 (P1_R1150_U338, P1_R1150_U47, P1_U3062);
  nand ginst2172 (P1_R1150_U339, P1_R1150_U337, P1_R1150_U338);
  nand ginst2173 (P1_R1150_U34, P1_R1150_U30, P1_U3060);
  nand ginst2174 (P1_R1150_U340, P1_R1150_U143, P1_R1150_U339);
  nand ginst2175 (P1_R1150_U341, P1_R1150_U174, P1_R1150_U90);
  nand ginst2176 (P1_R1150_U342, P1_R1150_U49, P1_U3485);
  nand ginst2177 (P1_R1150_U343, P1_R1150_U142, P1_R1150_U341);
  nand ginst2178 (P1_R1150_U344, P1_R1150_U47, P1_U3062);
  nand ginst2179 (P1_R1150_U345, P1_R1150_U174, P1_R1150_U344);
  nand ginst2180 (P1_R1150_U346, P1_R1150_U22, P1_U3077);
  nand ginst2181 (P1_R1150_U347, P1_R1150_U303, P1_R1150_U304, P1_R1150_U385);
  nand ginst2182 (P1_R1150_U348, P1_R1150_U40, P1_U3479);
  nand ginst2183 (P1_R1150_U349, P1_R1150_U39, P1_U3083);
  not ginst2184 (P1_R1150_U35, P1_U3476);
  nand ginst2185 (P1_R1150_U350, P1_R1150_U145, P1_R1150_U213);
  nand ginst2186 (P1_R1150_U351, P1_R1150_U144, P1_R1150_U211);
  nand ginst2187 (P1_R1150_U352, P1_R1150_U38, P1_U3476);
  nand ginst2188 (P1_R1150_U353, P1_R1150_U35, P1_U3084);
  nand ginst2189 (P1_R1150_U354, P1_R1150_U38, P1_U3476);
  nand ginst2190 (P1_R1150_U355, P1_R1150_U35, P1_U3084);
  nand ginst2191 (P1_R1150_U356, P1_R1150_U354, P1_R1150_U355);
  nand ginst2192 (P1_R1150_U357, P1_R1150_U36, P1_U3473);
  nand ginst2193 (P1_R1150_U358, P1_R1150_U19, P1_U3070);
  nand ginst2194 (P1_R1150_U359, P1_R1150_U218, P1_R1150_U41);
  not ginst2195 (P1_R1150_U36, P1_U3070);
  nand ginst2196 (P1_R1150_U360, P1_R1150_U146, P1_R1150_U205);
  nand ginst2197 (P1_R1150_U361, P1_R1150_U31, P1_U3470);
  nand ginst2198 (P1_R1150_U362, P1_R1150_U29, P1_U3071);
  nand ginst2199 (P1_R1150_U363, P1_R1150_U361, P1_R1150_U362);
  nand ginst2200 (P1_R1150_U364, P1_R1150_U32, P1_U3467);
  nand ginst2201 (P1_R1150_U365, P1_R1150_U20, P1_U3067);
  nand ginst2202 (P1_R1150_U366, P1_R1150_U228, P1_R1150_U42);
  nand ginst2203 (P1_R1150_U367, P1_R1150_U147, P1_R1150_U220);
  nand ginst2204 (P1_R1150_U368, P1_R1150_U33, P1_U3464);
  nand ginst2205 (P1_R1150_U369, P1_R1150_U30, P1_U3060);
  nand ginst2206 (P1_R1150_U37, P1_R1150_U19, P1_U3070);
  nand ginst2207 (P1_R1150_U370, P1_R1150_U149, P1_R1150_U229);
  nand ginst2208 (P1_R1150_U371, P1_R1150_U148, P1_R1150_U195);
  nand ginst2209 (P1_R1150_U372, P1_R1150_U28, P1_U3461);
  nand ginst2210 (P1_R1150_U373, P1_R1150_U25, P1_U3064);
  nand ginst2211 (P1_R1150_U374, P1_R1150_U28, P1_U3461);
  nand ginst2212 (P1_R1150_U375, P1_R1150_U25, P1_U3064);
  nand ginst2213 (P1_R1150_U376, P1_R1150_U374, P1_R1150_U375);
  nand ginst2214 (P1_R1150_U377, P1_R1150_U26, P1_U3458);
  nand ginst2215 (P1_R1150_U378, P1_R1150_U21, P1_U3068);
  nand ginst2216 (P1_R1150_U379, P1_R1150_U234, P1_R1150_U43);
  not ginst2217 (P1_R1150_U38, P1_U3084);
  nand ginst2218 (P1_R1150_U380, P1_R1150_U150, P1_R1150_U189);
  nand ginst2219 (P1_R1150_U381, P1_R1150_U152, P1_U3985);
  nand ginst2220 (P1_R1150_U382, P1_R1150_U151, P1_U3055);
  nand ginst2221 (P1_R1150_U383, P1_R1150_U152, P1_U3985);
  nand ginst2222 (P1_R1150_U384, P1_R1150_U151, P1_U3055);
  nand ginst2223 (P1_R1150_U385, P1_R1150_U383, P1_R1150_U384);
  nand ginst2224 (P1_R1150_U386, P1_R1150_U85, P1_U3974);
  nand ginst2225 (P1_R1150_U387, P1_R1150_U84, P1_U3054);
  not ginst2226 (P1_R1150_U388, P1_R1150_U127);
  nand ginst2227 (P1_R1150_U389, P1_R1150_U301, P1_R1150_U388);
  not ginst2228 (P1_R1150_U39, P1_U3479);
  nand ginst2229 (P1_R1150_U390, P1_R1150_U127, P1_R1150_U86);
  nand ginst2230 (P1_R1150_U391, P1_R1150_U83, P1_U3975);
  nand ginst2231 (P1_R1150_U392, P1_R1150_U80, P1_U3053);
  nand ginst2232 (P1_R1150_U393, P1_R1150_U83, P1_U3975);
  nand ginst2233 (P1_R1150_U394, P1_R1150_U80, P1_U3053);
  nand ginst2234 (P1_R1150_U395, P1_R1150_U393, P1_R1150_U394);
  nand ginst2235 (P1_R1150_U396, P1_R1150_U81, P1_U3976);
  nand ginst2236 (P1_R1150_U397, P1_R1150_U44, P1_U3057);
  nand ginst2237 (P1_R1150_U398, P1_R1150_U313, P1_R1150_U87);
  nand ginst2238 (P1_R1150_U399, P1_R1150_U154, P1_R1150_U295);
  not ginst2239 (P1_R1150_U40, P1_U3083);
  nand ginst2240 (P1_R1150_U400, P1_R1150_U79, P1_U3977);
  nand ginst2241 (P1_R1150_U401, P1_R1150_U78, P1_U3058);
  not ginst2242 (P1_R1150_U402, P1_R1150_U130);
  nand ginst2243 (P1_R1150_U403, P1_R1150_U291, P1_R1150_U402);
  nand ginst2244 (P1_R1150_U404, P1_R1150_U130, P1_R1150_U155);
  nand ginst2245 (P1_R1150_U405, P1_R1150_U77, P1_U3978);
  nand ginst2246 (P1_R1150_U406, P1_R1150_U76, P1_U3065);
  not ginst2247 (P1_R1150_U407, P1_R1150_U131);
  nand ginst2248 (P1_R1150_U408, P1_R1150_U287, P1_R1150_U407);
  nand ginst2249 (P1_R1150_U409, P1_R1150_U131, P1_R1150_U156);
  nand ginst2250 (P1_R1150_U41, P1_R1150_U203, P1_R1150_U204);
  nand ginst2251 (P1_R1150_U410, P1_R1150_U72, P1_U3979);
  nand ginst2252 (P1_R1150_U411, P1_R1150_U70, P1_U3066);
  nand ginst2253 (P1_R1150_U412, P1_R1150_U410, P1_R1150_U411);
  nand ginst2254 (P1_R1150_U413, P1_R1150_U73, P1_U3980);
  nand ginst2255 (P1_R1150_U414, P1_R1150_U45, P1_U3061);
  nand ginst2256 (P1_R1150_U415, P1_R1150_U323, P1_R1150_U88);
  nand ginst2257 (P1_R1150_U416, P1_R1150_U157, P1_R1150_U315);
  nand ginst2258 (P1_R1150_U417, P1_R1150_U74, P1_U3981);
  nand ginst2259 (P1_R1150_U418, P1_R1150_U71, P1_U3075);
  nand ginst2260 (P1_R1150_U419, P1_R1150_U159, P1_R1150_U324);
  nand ginst2261 (P1_R1150_U42, P1_R1150_U219, P1_R1150_U34);
  nand ginst2262 (P1_R1150_U420, P1_R1150_U158, P1_R1150_U277);
  nand ginst2263 (P1_R1150_U421, P1_R1150_U69, P1_U3982);
  nand ginst2264 (P1_R1150_U422, P1_R1150_U68, P1_U3076);
  not ginst2265 (P1_R1150_U423, P1_R1150_U133);
  nand ginst2266 (P1_R1150_U424, P1_R1150_U273, P1_R1150_U423);
  nand ginst2267 (P1_R1150_U425, P1_R1150_U133, P1_R1150_U160);
  nand ginst2268 (P1_R1150_U426, P1_R1150_U185, P1_R1150_U24);
  nand ginst2269 (P1_R1150_U427, P1_R1150_U23, P1_U3078);
  not ginst2270 (P1_R1150_U428, P1_R1150_U134);
  nand ginst2271 (P1_R1150_U429, P1_R1150_U428, P1_U3455);
  nand ginst2272 (P1_R1150_U43, P1_R1150_U187, P1_R1150_U188);
  nand ginst2273 (P1_R1150_U430, P1_R1150_U134, P1_R1150_U161);
  nand ginst2274 (P1_R1150_U431, P1_R1150_U67, P1_U3508);
  nand ginst2275 (P1_R1150_U432, P1_R1150_U66, P1_U3081);
  not ginst2276 (P1_R1150_U433, P1_R1150_U135);
  nand ginst2277 (P1_R1150_U434, P1_R1150_U269, P1_R1150_U433);
  nand ginst2278 (P1_R1150_U435, P1_R1150_U135, P1_R1150_U162);
  nand ginst2279 (P1_R1150_U436, P1_R1150_U65, P1_U3506);
  nand ginst2280 (P1_R1150_U437, P1_R1150_U163, P1_U3082);
  not ginst2281 (P1_R1150_U438, P1_R1150_U136);
  nand ginst2282 (P1_R1150_U439, P1_R1150_U265, P1_R1150_U438);
  not ginst2283 (P1_R1150_U44, P1_U3976);
  nand ginst2284 (P1_R1150_U440, P1_R1150_U136, P1_R1150_U64);
  nand ginst2285 (P1_R1150_U441, P1_R1150_U63, P1_U3503);
  nand ginst2286 (P1_R1150_U442, P1_R1150_U62, P1_U3069);
  not ginst2287 (P1_R1150_U443, P1_R1150_U137);
  nand ginst2288 (P1_R1150_U444, P1_R1150_U261, P1_R1150_U443);
  nand ginst2289 (P1_R1150_U445, P1_R1150_U137, P1_R1150_U164);
  nand ginst2290 (P1_R1150_U446, P1_R1150_U58, P1_U3500);
  nand ginst2291 (P1_R1150_U447, P1_R1150_U56, P1_U3073);
  nand ginst2292 (P1_R1150_U448, P1_R1150_U446, P1_R1150_U447);
  nand ginst2293 (P1_R1150_U449, P1_R1150_U59, P1_U3497);
  not ginst2294 (P1_R1150_U45, P1_U3980);
  nand ginst2295 (P1_R1150_U450, P1_R1150_U46, P1_U3074);
  nand ginst2296 (P1_R1150_U451, P1_R1150_U334, P1_R1150_U89);
  nand ginst2297 (P1_R1150_U452, P1_R1150_U165, P1_R1150_U326);
  nand ginst2298 (P1_R1150_U453, P1_R1150_U60, P1_U3494);
  nand ginst2299 (P1_R1150_U454, P1_R1150_U57, P1_U3079);
  nand ginst2300 (P1_R1150_U455, P1_R1150_U167, P1_R1150_U335);
  nand ginst2301 (P1_R1150_U456, P1_R1150_U166, P1_R1150_U251);
  nand ginst2302 (P1_R1150_U457, P1_R1150_U55, P1_U3491);
  nand ginst2303 (P1_R1150_U458, P1_R1150_U54, P1_U3080);
  not ginst2304 (P1_R1150_U459, P1_R1150_U140);
  not ginst2305 (P1_R1150_U46, P1_U3497);
  nand ginst2306 (P1_R1150_U460, P1_R1150_U247, P1_R1150_U459);
  nand ginst2307 (P1_R1150_U461, P1_R1150_U140, P1_R1150_U168);
  nand ginst2308 (P1_R1150_U462, P1_R1150_U53, P1_U3488);
  nand ginst2309 (P1_R1150_U463, P1_R1150_U52, P1_U3072);
  not ginst2310 (P1_R1150_U464, P1_R1150_U141);
  nand ginst2311 (P1_R1150_U465, P1_R1150_U243, P1_R1150_U464);
  nand ginst2312 (P1_R1150_U466, P1_R1150_U141, P1_R1150_U169);
  nand ginst2313 (P1_R1150_U467, P1_R1150_U49, P1_U3485);
  nand ginst2314 (P1_R1150_U468, P1_R1150_U48, P1_U3063);
  nand ginst2315 (P1_R1150_U469, P1_R1150_U467, P1_R1150_U468);
  not ginst2316 (P1_R1150_U47, P1_U3482);
  nand ginst2317 (P1_R1150_U470, P1_R1150_U50, P1_U3482);
  nand ginst2318 (P1_R1150_U471, P1_R1150_U47, P1_U3062);
  nand ginst2319 (P1_R1150_U472, P1_R1150_U345, P1_R1150_U90);
  nand ginst2320 (P1_R1150_U473, P1_R1150_U170, P1_R1150_U337);
  not ginst2321 (P1_R1150_U48, P1_U3485);
  not ginst2322 (P1_R1150_U49, P1_U3063);
  not ginst2323 (P1_R1150_U50, P1_U3062);
  nand ginst2324 (P1_R1150_U51, P1_R1150_U39, P1_U3083);
  not ginst2325 (P1_R1150_U52, P1_U3488);
  not ginst2326 (P1_R1150_U53, P1_U3072);
  not ginst2327 (P1_R1150_U54, P1_U3491);
  not ginst2328 (P1_R1150_U55, P1_U3080);
  not ginst2329 (P1_R1150_U56, P1_U3500);
  not ginst2330 (P1_R1150_U57, P1_U3494);
  not ginst2331 (P1_R1150_U58, P1_U3073);
  not ginst2332 (P1_R1150_U59, P1_U3074);
  and ginst2333 (P1_R1150_U6, P1_R1150_U197, P1_R1150_U198);
  not ginst2334 (P1_R1150_U60, P1_U3079);
  nand ginst2335 (P1_R1150_U61, P1_R1150_U57, P1_U3079);
  not ginst2336 (P1_R1150_U62, P1_U3503);
  not ginst2337 (P1_R1150_U63, P1_U3069);
  nand ginst2338 (P1_R1150_U64, P1_R1150_U263, P1_R1150_U264);
  not ginst2339 (P1_R1150_U65, P1_U3082);
  not ginst2340 (P1_R1150_U66, P1_U3508);
  not ginst2341 (P1_R1150_U67, P1_U3081);
  not ginst2342 (P1_R1150_U68, P1_U3982);
  not ginst2343 (P1_R1150_U69, P1_U3076);
  and ginst2344 (P1_R1150_U7, P1_R1150_U236, P1_R1150_U237);
  not ginst2345 (P1_R1150_U70, P1_U3979);
  not ginst2346 (P1_R1150_U71, P1_U3981);
  not ginst2347 (P1_R1150_U72, P1_U3066);
  not ginst2348 (P1_R1150_U73, P1_U3061);
  not ginst2349 (P1_R1150_U74, P1_U3075);
  nand ginst2350 (P1_R1150_U75, P1_R1150_U71, P1_U3075);
  not ginst2351 (P1_R1150_U76, P1_U3978);
  not ginst2352 (P1_R1150_U77, P1_U3065);
  not ginst2353 (P1_R1150_U78, P1_U3977);
  not ginst2354 (P1_R1150_U79, P1_U3058);
  and ginst2355 (P1_R1150_U8, P1_R1150_U253, P1_R1150_U254);
  not ginst2356 (P1_R1150_U80, P1_U3975);
  not ginst2357 (P1_R1150_U81, P1_U3057);
  nand ginst2358 (P1_R1150_U82, P1_R1150_U44, P1_U3057);
  not ginst2359 (P1_R1150_U83, P1_U3053);
  not ginst2360 (P1_R1150_U84, P1_U3974);
  not ginst2361 (P1_R1150_U85, P1_U3054);
  nand ginst2362 (P1_R1150_U86, P1_R1150_U126, P1_R1150_U297);
  nand ginst2363 (P1_R1150_U87, P1_R1150_U293, P1_R1150_U294);
  nand ginst2364 (P1_R1150_U88, P1_R1150_U314, P1_R1150_U75);
  nand ginst2365 (P1_R1150_U89, P1_R1150_U325, P1_R1150_U61);
  and ginst2366 (P1_R1150_U9, P1_R1150_U279, P1_R1150_U280);
  nand ginst2367 (P1_R1150_U90, P1_R1150_U336, P1_R1150_U51);
  not ginst2368 (P1_R1150_U91, P1_U3077);
  nand ginst2369 (P1_R1150_U92, P1_R1150_U389, P1_R1150_U390);
  nand ginst2370 (P1_R1150_U93, P1_R1150_U403, P1_R1150_U404);
  nand ginst2371 (P1_R1150_U94, P1_R1150_U408, P1_R1150_U409);
  nand ginst2372 (P1_R1150_U95, P1_R1150_U424, P1_R1150_U425);
  nand ginst2373 (P1_R1150_U96, P1_R1150_U429, P1_R1150_U430);
  nand ginst2374 (P1_R1150_U97, P1_R1150_U434, P1_R1150_U435);
  nand ginst2375 (P1_R1150_U98, P1_R1150_U439, P1_R1150_U440);
  nand ginst2376 (P1_R1150_U99, P1_R1150_U444, P1_R1150_U445);
  and ginst2377 (P1_R1162_U10, P1_R1162_U215, P1_R1162_U218);
  not ginst2378 (P1_R1162_U100, P1_R1162_U40);
  not ginst2379 (P1_R1162_U101, P1_R1162_U41);
  nand ginst2380 (P1_R1162_U102, P1_R1162_U40, P1_R1162_U41);
  nand ginst2381 (P1_R1162_U103, P1_REG1_REG_2__SCAN_IN, P1_R1162_U96, P1_U3457);
  nand ginst2382 (P1_R1162_U104, P1_R1162_U102, P1_R1162_U5);
  nand ginst2383 (P1_R1162_U105, P1_REG1_REG_3__SCAN_IN, P1_U3460);
  nand ginst2384 (P1_R1162_U106, P1_R1162_U103, P1_R1162_U104, P1_R1162_U105);
  nand ginst2385 (P1_R1162_U107, P1_R1162_U32, P1_R1162_U33);
  nand ginst2386 (P1_R1162_U108, P1_R1162_U107, P1_U3466);
  nand ginst2387 (P1_R1162_U109, P1_R1162_U106, P1_R1162_U4);
  and ginst2388 (P1_R1162_U11, P1_R1162_U208, P1_R1162_U211);
  nand ginst2389 (P1_R1162_U110, P1_REG1_REG_5__SCAN_IN, P1_R1162_U89);
  not ginst2390 (P1_R1162_U111, P1_R1162_U39);
  or ginst2391 (P1_R1162_U112, P1_REG1_REG_7__SCAN_IN, P1_U3472);
  or ginst2392 (P1_R1162_U113, P1_REG1_REG_6__SCAN_IN, P1_U3469);
  not ginst2393 (P1_R1162_U114, P1_R1162_U20);
  nand ginst2394 (P1_R1162_U115, P1_R1162_U20, P1_R1162_U21);
  nand ginst2395 (P1_R1162_U116, P1_R1162_U115, P1_U3472);
  nand ginst2396 (P1_R1162_U117, P1_REG1_REG_7__SCAN_IN, P1_R1162_U114);
  nand ginst2397 (P1_R1162_U118, P1_R1162_U39, P1_R1162_U6);
  not ginst2398 (P1_R1162_U119, P1_R1162_U81);
  and ginst2399 (P1_R1162_U12, P1_R1162_U199, P1_R1162_U202);
  or ginst2400 (P1_R1162_U120, P1_REG1_REG_8__SCAN_IN, P1_U3475);
  nand ginst2401 (P1_R1162_U121, P1_R1162_U120, P1_R1162_U81);
  not ginst2402 (P1_R1162_U122, P1_R1162_U38);
  or ginst2403 (P1_R1162_U123, P1_REG1_REG_9__SCAN_IN, P1_U3478);
  or ginst2404 (P1_R1162_U124, P1_REG1_REG_6__SCAN_IN, P1_U3469);
  nand ginst2405 (P1_R1162_U125, P1_R1162_U124, P1_R1162_U39);
  nand ginst2406 (P1_R1162_U126, P1_R1162_U125, P1_R1162_U20, P1_R1162_U237, P1_R1162_U238);
  nand ginst2407 (P1_R1162_U127, P1_R1162_U111, P1_R1162_U20);
  nand ginst2408 (P1_R1162_U128, P1_REG1_REG_7__SCAN_IN, P1_U3472);
  nand ginst2409 (P1_R1162_U129, P1_R1162_U127, P1_R1162_U128, P1_R1162_U6);
  and ginst2410 (P1_R1162_U13, P1_R1162_U192, P1_R1162_U196);
  or ginst2411 (P1_R1162_U130, P1_REG1_REG_6__SCAN_IN, P1_U3469);
  nand ginst2412 (P1_R1162_U131, P1_R1162_U101, P1_R1162_U97);
  nand ginst2413 (P1_R1162_U132, P1_REG1_REG_2__SCAN_IN, P1_U3457);
  not ginst2414 (P1_R1162_U133, P1_R1162_U43);
  nand ginst2415 (P1_R1162_U134, P1_R1162_U100, P1_R1162_U5);
  nand ginst2416 (P1_R1162_U135, P1_R1162_U43, P1_R1162_U96);
  nand ginst2417 (P1_R1162_U136, P1_REG1_REG_3__SCAN_IN, P1_U3460);
  not ginst2418 (P1_R1162_U137, P1_R1162_U42);
  or ginst2419 (P1_R1162_U138, P1_REG1_REG_4__SCAN_IN, P1_U3463);
  nand ginst2420 (P1_R1162_U139, P1_R1162_U138, P1_R1162_U42);
  and ginst2421 (P1_R1162_U14, P1_R1162_U148, P1_R1162_U151);
  nand ginst2422 (P1_R1162_U140, P1_R1162_U139, P1_R1162_U244, P1_R1162_U245, P1_R1162_U32);
  nand ginst2423 (P1_R1162_U141, P1_R1162_U137, P1_R1162_U32);
  nand ginst2424 (P1_R1162_U142, P1_REG1_REG_5__SCAN_IN, P1_U3466);
  nand ginst2425 (P1_R1162_U143, P1_R1162_U141, P1_R1162_U142, P1_R1162_U4);
  or ginst2426 (P1_R1162_U144, P1_REG1_REG_4__SCAN_IN, P1_U3463);
  nand ginst2427 (P1_R1162_U145, P1_R1162_U100, P1_R1162_U97);
  not ginst2428 (P1_R1162_U146, P1_R1162_U82);
  nand ginst2429 (P1_R1162_U147, P1_REG1_REG_3__SCAN_IN, P1_U3460);
  nand ginst2430 (P1_R1162_U148, P1_R1162_U256, P1_R1162_U257, P1_R1162_U40, P1_R1162_U41);
  nand ginst2431 (P1_R1162_U149, P1_R1162_U40, P1_R1162_U41);
  and ginst2432 (P1_R1162_U15, P1_R1162_U140, P1_R1162_U143);
  nand ginst2433 (P1_R1162_U150, P1_REG1_REG_2__SCAN_IN, P1_U3457);
  nand ginst2434 (P1_R1162_U151, P1_R1162_U149, P1_R1162_U150, P1_R1162_U97);
  or ginst2435 (P1_R1162_U152, P1_REG1_REG_1__SCAN_IN, P1_U3454);
  not ginst2436 (P1_R1162_U153, P1_R1162_U83);
  or ginst2437 (P1_R1162_U154, P1_REG1_REG_9__SCAN_IN, P1_U3478);
  or ginst2438 (P1_R1162_U155, P1_REG1_REG_10__SCAN_IN, P1_U3481);
  nand ginst2439 (P1_R1162_U156, P1_R1162_U7, P1_R1162_U93);
  nand ginst2440 (P1_R1162_U157, P1_REG1_REG_10__SCAN_IN, P1_U3481);
  nand ginst2441 (P1_R1162_U158, P1_R1162_U156, P1_R1162_U157, P1_R1162_U90);
  or ginst2442 (P1_R1162_U159, P1_REG1_REG_10__SCAN_IN, P1_U3481);
  and ginst2443 (P1_R1162_U16, P1_R1162_U126, P1_R1162_U129);
  nand ginst2444 (P1_R1162_U160, P1_R1162_U120, P1_R1162_U7, P1_R1162_U81);
  nand ginst2445 (P1_R1162_U161, P1_R1162_U158, P1_R1162_U159);
  not ginst2446 (P1_R1162_U162, P1_R1162_U88);
  or ginst2447 (P1_R1162_U163, P1_REG1_REG_13__SCAN_IN, P1_U3490);
  or ginst2448 (P1_R1162_U164, P1_REG1_REG_12__SCAN_IN, P1_U3487);
  nand ginst2449 (P1_R1162_U165, P1_R1162_U8, P1_R1162_U92);
  nand ginst2450 (P1_R1162_U166, P1_REG1_REG_13__SCAN_IN, P1_U3490);
  nand ginst2451 (P1_R1162_U167, P1_R1162_U165, P1_R1162_U166, P1_R1162_U91);
  or ginst2452 (P1_R1162_U168, P1_REG1_REG_11__SCAN_IN, P1_U3484);
  or ginst2453 (P1_R1162_U169, P1_REG1_REG_13__SCAN_IN, P1_U3490);
  not ginst2454 (P1_R1162_U17, P1_REG1_REG_6__SCAN_IN);
  nand ginst2455 (P1_R1162_U170, P1_R1162_U168, P1_R1162_U8, P1_R1162_U88);
  nand ginst2456 (P1_R1162_U171, P1_R1162_U167, P1_R1162_U169);
  not ginst2457 (P1_R1162_U172, P1_R1162_U87);
  or ginst2458 (P1_R1162_U173, P1_REG1_REG_14__SCAN_IN, P1_U3493);
  nand ginst2459 (P1_R1162_U174, P1_R1162_U173, P1_R1162_U87);
  nand ginst2460 (P1_R1162_U175, P1_REG1_REG_14__SCAN_IN, P1_U3493);
  not ginst2461 (P1_R1162_U176, P1_R1162_U86);
  or ginst2462 (P1_R1162_U177, P1_REG1_REG_15__SCAN_IN, P1_U3496);
  nand ginst2463 (P1_R1162_U178, P1_R1162_U177, P1_R1162_U86);
  nand ginst2464 (P1_R1162_U179, P1_REG1_REG_15__SCAN_IN, P1_U3496);
  not ginst2465 (P1_R1162_U18, P1_U3469);
  not ginst2466 (P1_R1162_U180, P1_R1162_U66);
  or ginst2467 (P1_R1162_U181, P1_REG1_REG_17__SCAN_IN, P1_U3502);
  or ginst2468 (P1_R1162_U182, P1_REG1_REG_16__SCAN_IN, P1_U3499);
  not ginst2469 (P1_R1162_U183, P1_R1162_U47);
  nand ginst2470 (P1_R1162_U184, P1_R1162_U47, P1_R1162_U48);
  nand ginst2471 (P1_R1162_U185, P1_R1162_U184, P1_U3502);
  nand ginst2472 (P1_R1162_U186, P1_REG1_REG_17__SCAN_IN, P1_R1162_U183);
  nand ginst2473 (P1_R1162_U187, P1_R1162_U66, P1_R1162_U9);
  not ginst2474 (P1_R1162_U188, P1_R1162_U65);
  or ginst2475 (P1_R1162_U189, P1_REG1_REG_18__SCAN_IN, P1_U3505);
  not ginst2476 (P1_R1162_U19, P1_U3472);
  nand ginst2477 (P1_R1162_U190, P1_R1162_U189, P1_R1162_U65);
  nand ginst2478 (P1_R1162_U191, P1_REG1_REG_18__SCAN_IN, P1_U3505);
  nand ginst2479 (P1_R1162_U192, P1_R1162_U190, P1_R1162_U191, P1_R1162_U260, P1_R1162_U261);
  nand ginst2480 (P1_R1162_U193, P1_REG1_REG_18__SCAN_IN, P1_U3505);
  nand ginst2481 (P1_R1162_U194, P1_R1162_U188, P1_R1162_U193);
  or ginst2482 (P1_R1162_U195, P1_REG1_REG_18__SCAN_IN, P1_U3505);
  nand ginst2483 (P1_R1162_U196, P1_R1162_U194, P1_R1162_U195, P1_R1162_U264);
  or ginst2484 (P1_R1162_U197, P1_REG1_REG_16__SCAN_IN, P1_U3499);
  nand ginst2485 (P1_R1162_U198, P1_R1162_U197, P1_R1162_U66);
  nand ginst2486 (P1_R1162_U199, P1_R1162_U198, P1_R1162_U272, P1_R1162_U273, P1_R1162_U47);
  nand ginst2487 (P1_R1162_U20, P1_REG1_REG_6__SCAN_IN, P1_U3469);
  nand ginst2488 (P1_R1162_U200, P1_R1162_U180, P1_R1162_U47);
  nand ginst2489 (P1_R1162_U201, P1_REG1_REG_17__SCAN_IN, P1_U3502);
  nand ginst2490 (P1_R1162_U202, P1_R1162_U200, P1_R1162_U201, P1_R1162_U9);
  or ginst2491 (P1_R1162_U203, P1_REG1_REG_16__SCAN_IN, P1_U3499);
  nand ginst2492 (P1_R1162_U204, P1_R1162_U168, P1_R1162_U88);
  not ginst2493 (P1_R1162_U205, P1_R1162_U67);
  or ginst2494 (P1_R1162_U206, P1_REG1_REG_12__SCAN_IN, P1_U3487);
  nand ginst2495 (P1_R1162_U207, P1_R1162_U206, P1_R1162_U67);
  nand ginst2496 (P1_R1162_U208, P1_R1162_U207, P1_R1162_U293, P1_R1162_U294, P1_R1162_U91);
  nand ginst2497 (P1_R1162_U209, P1_R1162_U205, P1_R1162_U91);
  not ginst2498 (P1_R1162_U21, P1_REG1_REG_7__SCAN_IN);
  nand ginst2499 (P1_R1162_U210, P1_REG1_REG_13__SCAN_IN, P1_U3490);
  nand ginst2500 (P1_R1162_U211, P1_R1162_U209, P1_R1162_U210, P1_R1162_U8);
  or ginst2501 (P1_R1162_U212, P1_REG1_REG_12__SCAN_IN, P1_U3487);
  or ginst2502 (P1_R1162_U213, P1_REG1_REG_9__SCAN_IN, P1_U3478);
  nand ginst2503 (P1_R1162_U214, P1_R1162_U213, P1_R1162_U38);
  nand ginst2504 (P1_R1162_U215, P1_R1162_U214, P1_R1162_U305, P1_R1162_U306, P1_R1162_U90);
  nand ginst2505 (P1_R1162_U216, P1_R1162_U122, P1_R1162_U90);
  nand ginst2506 (P1_R1162_U217, P1_REG1_REG_10__SCAN_IN, P1_U3481);
  nand ginst2507 (P1_R1162_U218, P1_R1162_U216, P1_R1162_U217, P1_R1162_U7);
  nand ginst2508 (P1_R1162_U219, P1_R1162_U123, P1_R1162_U90);
  not ginst2509 (P1_R1162_U22, P1_REG1_REG_4__SCAN_IN);
  nand ginst2510 (P1_R1162_U220, P1_R1162_U120, P1_R1162_U49);
  nand ginst2511 (P1_R1162_U221, P1_R1162_U130, P1_R1162_U20);
  nand ginst2512 (P1_R1162_U222, P1_R1162_U144, P1_R1162_U32);
  nand ginst2513 (P1_R1162_U223, P1_R1162_U147, P1_R1162_U96);
  nand ginst2514 (P1_R1162_U224, P1_R1162_U203, P1_R1162_U47);
  nand ginst2515 (P1_R1162_U225, P1_R1162_U212, P1_R1162_U91);
  nand ginst2516 (P1_R1162_U226, P1_R1162_U168, P1_R1162_U56);
  nand ginst2517 (P1_R1162_U227, P1_R1162_U37, P1_U3478);
  nand ginst2518 (P1_R1162_U228, P1_REG1_REG_9__SCAN_IN, P1_R1162_U36);
  nand ginst2519 (P1_R1162_U229, P1_R1162_U227, P1_R1162_U228);
  not ginst2520 (P1_R1162_U23, P1_U3463);
  nand ginst2521 (P1_R1162_U230, P1_R1162_U219, P1_R1162_U38);
  nand ginst2522 (P1_R1162_U231, P1_R1162_U122, P1_R1162_U229);
  nand ginst2523 (P1_R1162_U232, P1_R1162_U34, P1_U3475);
  nand ginst2524 (P1_R1162_U233, P1_REG1_REG_8__SCAN_IN, P1_R1162_U35);
  nand ginst2525 (P1_R1162_U234, P1_R1162_U232, P1_R1162_U233);
  nand ginst2526 (P1_R1162_U235, P1_R1162_U220, P1_R1162_U81);
  nand ginst2527 (P1_R1162_U236, P1_R1162_U119, P1_R1162_U234);
  nand ginst2528 (P1_R1162_U237, P1_R1162_U21, P1_U3472);
  nand ginst2529 (P1_R1162_U238, P1_REG1_REG_7__SCAN_IN, P1_R1162_U19);
  nand ginst2530 (P1_R1162_U239, P1_R1162_U17, P1_U3469);
  not ginst2531 (P1_R1162_U24, P1_U3466);
  nand ginst2532 (P1_R1162_U240, P1_REG1_REG_6__SCAN_IN, P1_R1162_U18);
  nand ginst2533 (P1_R1162_U241, P1_R1162_U239, P1_R1162_U240);
  nand ginst2534 (P1_R1162_U242, P1_R1162_U221, P1_R1162_U39);
  nand ginst2535 (P1_R1162_U243, P1_R1162_U111, P1_R1162_U241);
  nand ginst2536 (P1_R1162_U244, P1_R1162_U33, P1_U3466);
  nand ginst2537 (P1_R1162_U245, P1_REG1_REG_5__SCAN_IN, P1_R1162_U24);
  nand ginst2538 (P1_R1162_U246, P1_R1162_U22, P1_U3463);
  nand ginst2539 (P1_R1162_U247, P1_REG1_REG_4__SCAN_IN, P1_R1162_U23);
  nand ginst2540 (P1_R1162_U248, P1_R1162_U246, P1_R1162_U247);
  nand ginst2541 (P1_R1162_U249, P1_R1162_U222, P1_R1162_U42);
  not ginst2542 (P1_R1162_U25, P1_REG1_REG_2__SCAN_IN);
  nand ginst2543 (P1_R1162_U250, P1_R1162_U137, P1_R1162_U248);
  nand ginst2544 (P1_R1162_U251, P1_R1162_U30, P1_U3460);
  nand ginst2545 (P1_R1162_U252, P1_REG1_REG_3__SCAN_IN, P1_R1162_U31);
  nand ginst2546 (P1_R1162_U253, P1_R1162_U251, P1_R1162_U252);
  nand ginst2547 (P1_R1162_U254, P1_R1162_U223, P1_R1162_U82);
  nand ginst2548 (P1_R1162_U255, P1_R1162_U146, P1_R1162_U253);
  nand ginst2549 (P1_R1162_U256, P1_R1162_U25, P1_U3457);
  nand ginst2550 (P1_R1162_U257, P1_REG1_REG_2__SCAN_IN, P1_R1162_U26);
  nand ginst2551 (P1_R1162_U258, P1_R1162_U83, P1_R1162_U98);
  nand ginst2552 (P1_R1162_U259, P1_R1162_U153, P1_R1162_U29);
  not ginst2553 (P1_R1162_U26, P1_U3457);
  nand ginst2554 (P1_R1162_U260, P1_R1162_U85, P1_U3442);
  nand ginst2555 (P1_R1162_U261, P1_REG1_REG_19__SCAN_IN, P1_R1162_U84);
  nand ginst2556 (P1_R1162_U262, P1_R1162_U85, P1_U3442);
  nand ginst2557 (P1_R1162_U263, P1_REG1_REG_19__SCAN_IN, P1_R1162_U84);
  nand ginst2558 (P1_R1162_U264, P1_R1162_U262, P1_R1162_U263);
  nand ginst2559 (P1_R1162_U265, P1_R1162_U63, P1_U3505);
  nand ginst2560 (P1_R1162_U266, P1_REG1_REG_18__SCAN_IN, P1_R1162_U64);
  nand ginst2561 (P1_R1162_U267, P1_R1162_U63, P1_U3505);
  nand ginst2562 (P1_R1162_U268, P1_REG1_REG_18__SCAN_IN, P1_R1162_U64);
  nand ginst2563 (P1_R1162_U269, P1_R1162_U267, P1_R1162_U268);
  not ginst2564 (P1_R1162_U27, P1_REG1_REG_0__SCAN_IN);
  nand ginst2565 (P1_R1162_U270, P1_R1162_U265, P1_R1162_U266, P1_R1162_U65);
  nand ginst2566 (P1_R1162_U271, P1_R1162_U188, P1_R1162_U269);
  nand ginst2567 (P1_R1162_U272, P1_R1162_U48, P1_U3502);
  nand ginst2568 (P1_R1162_U273, P1_REG1_REG_17__SCAN_IN, P1_R1162_U46);
  nand ginst2569 (P1_R1162_U274, P1_R1162_U44, P1_U3499);
  nand ginst2570 (P1_R1162_U275, P1_REG1_REG_16__SCAN_IN, P1_R1162_U45);
  nand ginst2571 (P1_R1162_U276, P1_R1162_U274, P1_R1162_U275);
  nand ginst2572 (P1_R1162_U277, P1_R1162_U224, P1_R1162_U66);
  nand ginst2573 (P1_R1162_U278, P1_R1162_U180, P1_R1162_U276);
  nand ginst2574 (P1_R1162_U279, P1_R1162_U61, P1_U3496);
  not ginst2575 (P1_R1162_U28, P1_U3448);
  nand ginst2576 (P1_R1162_U280, P1_REG1_REG_15__SCAN_IN, P1_R1162_U62);
  nand ginst2577 (P1_R1162_U281, P1_R1162_U61, P1_U3496);
  nand ginst2578 (P1_R1162_U282, P1_REG1_REG_15__SCAN_IN, P1_R1162_U62);
  nand ginst2579 (P1_R1162_U283, P1_R1162_U281, P1_R1162_U282);
  nand ginst2580 (P1_R1162_U284, P1_R1162_U279, P1_R1162_U280, P1_R1162_U86);
  nand ginst2581 (P1_R1162_U285, P1_R1162_U176, P1_R1162_U283);
  nand ginst2582 (P1_R1162_U286, P1_R1162_U59, P1_U3493);
  nand ginst2583 (P1_R1162_U287, P1_REG1_REG_14__SCAN_IN, P1_R1162_U60);
  nand ginst2584 (P1_R1162_U288, P1_R1162_U59, P1_U3493);
  nand ginst2585 (P1_R1162_U289, P1_REG1_REG_14__SCAN_IN, P1_R1162_U60);
  nand ginst2586 (P1_R1162_U29, P1_REG1_REG_0__SCAN_IN, P1_U3448);
  nand ginst2587 (P1_R1162_U290, P1_R1162_U288, P1_R1162_U289);
  nand ginst2588 (P1_R1162_U291, P1_R1162_U286, P1_R1162_U287, P1_R1162_U87);
  nand ginst2589 (P1_R1162_U292, P1_R1162_U172, P1_R1162_U290);
  nand ginst2590 (P1_R1162_U293, P1_R1162_U57, P1_U3490);
  nand ginst2591 (P1_R1162_U294, P1_REG1_REG_13__SCAN_IN, P1_R1162_U58);
  nand ginst2592 (P1_R1162_U295, P1_R1162_U52, P1_U3487);
  nand ginst2593 (P1_R1162_U296, P1_REG1_REG_12__SCAN_IN, P1_R1162_U53);
  nand ginst2594 (P1_R1162_U297, P1_R1162_U295, P1_R1162_U296);
  nand ginst2595 (P1_R1162_U298, P1_R1162_U225, P1_R1162_U67);
  nand ginst2596 (P1_R1162_U299, P1_R1162_U205, P1_R1162_U297);
  not ginst2597 (P1_R1162_U30, P1_REG1_REG_3__SCAN_IN);
  nand ginst2598 (P1_R1162_U300, P1_R1162_U54, P1_U3484);
  nand ginst2599 (P1_R1162_U301, P1_REG1_REG_11__SCAN_IN, P1_R1162_U55);
  nand ginst2600 (P1_R1162_U302, P1_R1162_U300, P1_R1162_U301);
  nand ginst2601 (P1_R1162_U303, P1_R1162_U226, P1_R1162_U88);
  nand ginst2602 (P1_R1162_U304, P1_R1162_U162, P1_R1162_U302);
  nand ginst2603 (P1_R1162_U305, P1_R1162_U50, P1_U3481);
  nand ginst2604 (P1_R1162_U306, P1_REG1_REG_10__SCAN_IN, P1_R1162_U51);
  nand ginst2605 (P1_R1162_U307, P1_R1162_U27, P1_U3448);
  nand ginst2606 (P1_R1162_U308, P1_REG1_REG_0__SCAN_IN, P1_R1162_U28);
  not ginst2607 (P1_R1162_U31, P1_U3460);
  nand ginst2608 (P1_R1162_U32, P1_REG1_REG_4__SCAN_IN, P1_U3463);
  not ginst2609 (P1_R1162_U33, P1_REG1_REG_5__SCAN_IN);
  not ginst2610 (P1_R1162_U34, P1_REG1_REG_8__SCAN_IN);
  not ginst2611 (P1_R1162_U35, P1_U3475);
  not ginst2612 (P1_R1162_U36, P1_U3478);
  not ginst2613 (P1_R1162_U37, P1_REG1_REG_9__SCAN_IN);
  nand ginst2614 (P1_R1162_U38, P1_R1162_U121, P1_R1162_U49);
  nand ginst2615 (P1_R1162_U39, P1_R1162_U108, P1_R1162_U109, P1_R1162_U110);
  and ginst2616 (P1_R1162_U4, P1_R1162_U94, P1_R1162_U95);
  nand ginst2617 (P1_R1162_U40, P1_R1162_U98, P1_R1162_U99);
  nand ginst2618 (P1_R1162_U41, P1_REG1_REG_1__SCAN_IN, P1_U3454);
  nand ginst2619 (P1_R1162_U42, P1_R1162_U134, P1_R1162_U135, P1_R1162_U136);
  nand ginst2620 (P1_R1162_U43, P1_R1162_U131, P1_R1162_U132);
  not ginst2621 (P1_R1162_U44, P1_REG1_REG_16__SCAN_IN);
  not ginst2622 (P1_R1162_U45, P1_U3499);
  not ginst2623 (P1_R1162_U46, P1_U3502);
  nand ginst2624 (P1_R1162_U47, P1_REG1_REG_16__SCAN_IN, P1_U3499);
  not ginst2625 (P1_R1162_U48, P1_REG1_REG_17__SCAN_IN);
  nand ginst2626 (P1_R1162_U49, P1_REG1_REG_8__SCAN_IN, P1_U3475);
  and ginst2627 (P1_R1162_U5, P1_R1162_U96, P1_R1162_U97);
  not ginst2628 (P1_R1162_U50, P1_REG1_REG_10__SCAN_IN);
  not ginst2629 (P1_R1162_U51, P1_U3481);
  not ginst2630 (P1_R1162_U52, P1_REG1_REG_12__SCAN_IN);
  not ginst2631 (P1_R1162_U53, P1_U3487);
  not ginst2632 (P1_R1162_U54, P1_REG1_REG_11__SCAN_IN);
  not ginst2633 (P1_R1162_U55, P1_U3484);
  nand ginst2634 (P1_R1162_U56, P1_REG1_REG_11__SCAN_IN, P1_U3484);
  not ginst2635 (P1_R1162_U57, P1_REG1_REG_13__SCAN_IN);
  not ginst2636 (P1_R1162_U58, P1_U3490);
  not ginst2637 (P1_R1162_U59, P1_REG1_REG_14__SCAN_IN);
  and ginst2638 (P1_R1162_U6, P1_R1162_U112, P1_R1162_U113);
  not ginst2639 (P1_R1162_U60, P1_U3493);
  not ginst2640 (P1_R1162_U61, P1_REG1_REG_15__SCAN_IN);
  not ginst2641 (P1_R1162_U62, P1_U3496);
  not ginst2642 (P1_R1162_U63, P1_REG1_REG_18__SCAN_IN);
  not ginst2643 (P1_R1162_U64, P1_U3505);
  nand ginst2644 (P1_R1162_U65, P1_R1162_U185, P1_R1162_U186, P1_R1162_U187);
  nand ginst2645 (P1_R1162_U66, P1_R1162_U178, P1_R1162_U179);
  nand ginst2646 (P1_R1162_U67, P1_R1162_U204, P1_R1162_U56);
  nand ginst2647 (P1_R1162_U68, P1_R1162_U258, P1_R1162_U259);
  nand ginst2648 (P1_R1162_U69, P1_R1162_U307, P1_R1162_U308);
  and ginst2649 (P1_R1162_U7, P1_R1162_U154, P1_R1162_U155);
  nand ginst2650 (P1_R1162_U70, P1_R1162_U230, P1_R1162_U231);
  nand ginst2651 (P1_R1162_U71, P1_R1162_U235, P1_R1162_U236);
  nand ginst2652 (P1_R1162_U72, P1_R1162_U242, P1_R1162_U243);
  nand ginst2653 (P1_R1162_U73, P1_R1162_U249, P1_R1162_U250);
  nand ginst2654 (P1_R1162_U74, P1_R1162_U254, P1_R1162_U255);
  nand ginst2655 (P1_R1162_U75, P1_R1162_U270, P1_R1162_U271);
  nand ginst2656 (P1_R1162_U76, P1_R1162_U277, P1_R1162_U278);
  nand ginst2657 (P1_R1162_U77, P1_R1162_U284, P1_R1162_U285);
  nand ginst2658 (P1_R1162_U78, P1_R1162_U291, P1_R1162_U292);
  nand ginst2659 (P1_R1162_U79, P1_R1162_U298, P1_R1162_U299);
  and ginst2660 (P1_R1162_U8, P1_R1162_U163, P1_R1162_U164);
  nand ginst2661 (P1_R1162_U80, P1_R1162_U303, P1_R1162_U304);
  nand ginst2662 (P1_R1162_U81, P1_R1162_U116, P1_R1162_U117, P1_R1162_U118);
  nand ginst2663 (P1_R1162_U82, P1_R1162_U133, P1_R1162_U145);
  nand ginst2664 (P1_R1162_U83, P1_R1162_U152, P1_R1162_U41);
  not ginst2665 (P1_R1162_U84, P1_U3442);
  not ginst2666 (P1_R1162_U85, P1_REG1_REG_19__SCAN_IN);
  nand ginst2667 (P1_R1162_U86, P1_R1162_U174, P1_R1162_U175);
  nand ginst2668 (P1_R1162_U87, P1_R1162_U170, P1_R1162_U171);
  nand ginst2669 (P1_R1162_U88, P1_R1162_U160, P1_R1162_U161);
  not ginst2670 (P1_R1162_U89, P1_R1162_U32);
  and ginst2671 (P1_R1162_U9, P1_R1162_U181, P1_R1162_U182);
  nand ginst2672 (P1_R1162_U90, P1_REG1_REG_9__SCAN_IN, P1_U3478);
  nand ginst2673 (P1_R1162_U91, P1_REG1_REG_12__SCAN_IN, P1_U3487);
  not ginst2674 (P1_R1162_U92, P1_R1162_U56);
  not ginst2675 (P1_R1162_U93, P1_R1162_U49);
  or ginst2676 (P1_R1162_U94, P1_REG1_REG_5__SCAN_IN, P1_U3466);
  or ginst2677 (P1_R1162_U95, P1_REG1_REG_4__SCAN_IN, P1_U3463);
  or ginst2678 (P1_R1162_U96, P1_REG1_REG_3__SCAN_IN, P1_U3460);
  or ginst2679 (P1_R1162_U97, P1_REG1_REG_2__SCAN_IN, P1_U3457);
  not ginst2680 (P1_R1162_U98, P1_R1162_U29);
  or ginst2681 (P1_R1162_U99, P1_REG1_REG_1__SCAN_IN, P1_U3454);
  and ginst2682 (P1_R1165_U10, P1_R1165_U336, P1_R1165_U339);
  nand ginst2683 (P1_R1165_U100, P1_R1165_U544, P1_R1165_U545);
  nand ginst2684 (P1_R1165_U101, P1_R1165_U549, P1_R1165_U550);
  nand ginst2685 (P1_R1165_U102, P1_R1165_U556, P1_R1165_U557);
  nand ginst2686 (P1_R1165_U103, P1_R1165_U563, P1_R1165_U564);
  nand ginst2687 (P1_R1165_U104, P1_R1165_U570, P1_R1165_U571);
  nand ginst2688 (P1_R1165_U105, P1_R1165_U577, P1_R1165_U578);
  nand ginst2689 (P1_R1165_U106, P1_R1165_U584, P1_R1165_U585);
  nand ginst2690 (P1_R1165_U107, P1_R1165_U589, P1_R1165_U590);
  nand ginst2691 (P1_R1165_U108, P1_R1165_U596, P1_R1165_U597);
  and ginst2692 (P1_R1165_U109, P1_R1165_U212, P1_R1165_U213);
  and ginst2693 (P1_R1165_U11, P1_R1165_U327, P1_R1165_U330);
  and ginst2694 (P1_R1165_U110, P1_R1165_U225, P1_R1165_U226);
  and ginst2695 (P1_R1165_U111, P1_R1165_U18, P1_R1165_U409, P1_R1165_U410);
  and ginst2696 (P1_R1165_U112, P1_R1165_U237, P1_R1165_U5);
  and ginst2697 (P1_R1165_U113, P1_R1165_U22, P1_R1165_U430, P1_R1165_U431);
  and ginst2698 (P1_R1165_U114, P1_R1165_U244, P1_R1165_U4);
  and ginst2699 (P1_R1165_U115, P1_R1165_U257, P1_R1165_U6);
  and ginst2700 (P1_R1165_U116, P1_R1165_U195, P1_R1165_U255);
  and ginst2701 (P1_R1165_U117, P1_R1165_U274, P1_R1165_U275);
  and ginst2702 (P1_R1165_U118, P1_R1165_U287, P1_R1165_U8);
  and ginst2703 (P1_R1165_U119, P1_R1165_U196, P1_R1165_U285);
  and ginst2704 (P1_R1165_U12, P1_R1165_U320, P1_R1165_U323);
  and ginst2705 (P1_R1165_U120, P1_R1165_U359, P1_R1165_U52);
  and ginst2706 (P1_R1165_U121, P1_R1165_U303, P1_R1165_U308);
  and ginst2707 (P1_R1165_U122, P1_R1165_U307, P1_R1165_U356);
  nand ginst2708 (P1_R1165_U123, P1_R1165_U491, P1_R1165_U492);
  and ginst2709 (P1_R1165_U124, P1_R1165_U352, P1_R1165_U52);
  and ginst2710 (P1_R1165_U125, P1_R1165_U33, P1_R1165_U442);
  and ginst2711 (P1_R1165_U126, P1_R1165_U197, P1_R1165_U200);
  and ginst2712 (P1_R1165_U127, P1_R1165_U193, P1_R1165_U313);
  and ginst2713 (P1_R1165_U128, P1_R1165_U197, P1_R1165_U9);
  and ginst2714 (P1_R1165_U129, P1_R1165_U196, P1_R1165_U532, P1_R1165_U533);
  and ginst2715 (P1_R1165_U13, P1_R1165_U311, P1_R1165_U314, P1_R1165_U360);
  and ginst2716 (P1_R1165_U130, P1_R1165_U322, P1_R1165_U8);
  and ginst2717 (P1_R1165_U131, P1_R1165_U36, P1_R1165_U558, P1_R1165_U559);
  and ginst2718 (P1_R1165_U132, P1_R1165_U329, P1_R1165_U7);
  and ginst2719 (P1_R1165_U133, P1_R1165_U195, P1_R1165_U579, P1_R1165_U580);
  and ginst2720 (P1_R1165_U134, P1_R1165_U338, P1_R1165_U6);
  nand ginst2721 (P1_R1165_U135, P1_R1165_U598, P1_R1165_U599);
  not ginst2722 (P1_R1165_U136, P1_U3201);
  and ginst2723 (P1_R1165_U137, P1_R1165_U368, P1_R1165_U369);
  not ginst2724 (P1_R1165_U138, P1_U3206);
  not ginst2725 (P1_R1165_U139, P1_U3210);
  and ginst2726 (P1_R1165_U14, P1_R1165_U242, P1_R1165_U245);
  not ginst2727 (P1_R1165_U140, P1_U3209);
  not ginst2728 (P1_R1165_U141, P1_U3207);
  not ginst2729 (P1_R1165_U142, P1_U3208);
  not ginst2730 (P1_R1165_U143, P1_U3205);
  not ginst2731 (P1_R1165_U144, P1_U3203);
  not ginst2732 (P1_R1165_U145, P1_U3204);
  not ginst2733 (P1_R1165_U146, P1_U3202);
  nand ginst2734 (P1_R1165_U147, P1_R1165_U230, P1_R1165_U231);
  and ginst2735 (P1_R1165_U148, P1_R1165_U402, P1_R1165_U403);
  nand ginst2736 (P1_R1165_U149, P1_R1165_U110, P1_R1165_U227);
  and ginst2737 (P1_R1165_U15, P1_R1165_U235, P1_R1165_U238);
  and ginst2738 (P1_R1165_U150, P1_R1165_U416, P1_R1165_U417);
  nand ginst2739 (P1_R1165_U151, P1_R1165_U350, P1_R1165_U361);
  and ginst2740 (P1_R1165_U152, P1_R1165_U423, P1_R1165_U424);
  nand ginst2741 (P1_R1165_U153, P1_R1165_U109, P1_R1165_U214);
  not ginst2742 (P1_R1165_U154, P1_U3183);
  not ginst2743 (P1_R1165_U155, P1_U3185);
  not ginst2744 (P1_R1165_U156, P1_U3184);
  not ginst2745 (P1_R1165_U157, P1_U3186);
  not ginst2746 (P1_R1165_U158, P1_U3200);
  not ginst2747 (P1_R1165_U159, P1_U3197);
  not ginst2748 (P1_R1165_U16, P1_U3211);
  not ginst2749 (P1_R1165_U160, P1_U3198);
  not ginst2750 (P1_R1165_U161, P1_U3199);
  not ginst2751 (P1_R1165_U162, P1_U3196);
  not ginst2752 (P1_R1165_U163, P1_U3195);
  not ginst2753 (P1_R1165_U164, P1_U3193);
  not ginst2754 (P1_R1165_U165, P1_U3194);
  not ginst2755 (P1_R1165_U166, P1_U3192);
  not ginst2756 (P1_R1165_U167, P1_U3189);
  not ginst2757 (P1_R1165_U168, P1_U3190);
  not ginst2758 (P1_R1165_U169, P1_U3191);
  not ginst2759 (P1_R1165_U17, P1_U3175);
  not ginst2760 (P1_R1165_U170, P1_U3188);
  not ginst2761 (P1_R1165_U171, P1_U3187);
  not ginst2762 (P1_R1165_U172, P1_U3153);
  not ginst2763 (P1_R1165_U173, P1_U3182);
  and ginst2764 (P1_R1165_U174, P1_R1165_U499, P1_R1165_U500);
  nand ginst2765 (P1_R1165_U175, P1_R1165_U124, P1_R1165_U304);
  nand ginst2766 (P1_R1165_U176, P1_R1165_U297, P1_R1165_U298);
  and ginst2767 (P1_R1165_U177, P1_R1165_U518, P1_R1165_U519);
  nand ginst2768 (P1_R1165_U178, P1_R1165_U293, P1_R1165_U294);
  and ginst2769 (P1_R1165_U179, P1_R1165_U525, P1_R1165_U526);
  nand ginst2770 (P1_R1165_U18, P1_R1165_U58, P1_U3175);
  nand ginst2771 (P1_R1165_U180, P1_R1165_U289, P1_R1165_U290);
  and ginst2772 (P1_R1165_U181, P1_R1165_U539, P1_R1165_U540);
  nand ginst2773 (P1_R1165_U182, P1_R1165_U202, P1_R1165_U203);
  nand ginst2774 (P1_R1165_U183, P1_R1165_U279, P1_R1165_U280);
  and ginst2775 (P1_R1165_U184, P1_R1165_U551, P1_R1165_U552);
  nand ginst2776 (P1_R1165_U185, P1_R1165_U117, P1_R1165_U276);
  and ginst2777 (P1_R1165_U186, P1_R1165_U565, P1_R1165_U566);
  nand ginst2778 (P1_R1165_U187, P1_R1165_U263, P1_R1165_U264);
  and ginst2779 (P1_R1165_U188, P1_R1165_U572, P1_R1165_U573);
  nand ginst2780 (P1_R1165_U189, P1_R1165_U259, P1_R1165_U260);
  not ginst2781 (P1_R1165_U19, P1_U3174);
  nand ginst2782 (P1_R1165_U190, P1_R1165_U249, P1_R1165_U250);
  and ginst2783 (P1_R1165_U191, P1_R1165_U591, P1_R1165_U592);
  nand ginst2784 (P1_R1165_U192, P1_R1165_U353, P1_R1165_U363);
  nand ginst2785 (P1_R1165_U193, P1_R1165_U354, P1_R1165_U355);
  not ginst2786 (P1_R1165_U194, P1_R1165_U22);
  nand ginst2787 (P1_R1165_U195, P1_R1165_U76, P1_U3169);
  nand ginst2788 (P1_R1165_U196, P1_R1165_U82, P1_U3161);
  nand ginst2789 (P1_R1165_U197, P1_R1165_U68, P1_U3156);
  not ginst2790 (P1_R1165_U198, P1_R1165_U41);
  not ginst2791 (P1_R1165_U199, P1_R1165_U48);
  not ginst2792 (P1_R1165_U20, P1_U3177);
  nand ginst2793 (P1_R1165_U200, P1_R1165_U70, P1_U3157);
  or ginst2794 (P1_R1165_U201, P1_U3181, P1_U3211);
  nand ginst2795 (P1_R1165_U202, P1_R1165_U201, P1_R1165_U63);
  nand ginst2796 (P1_R1165_U203, P1_U3181, P1_U3211);
  not ginst2797 (P1_R1165_U204, P1_R1165_U182);
  nand ginst2798 (P1_R1165_U205, P1_R1165_U25, P1_R1165_U381);
  nand ginst2799 (P1_R1165_U206, P1_R1165_U182, P1_R1165_U205);
  nand ginst2800 (P1_R1165_U207, P1_R1165_U64, P1_U3180);
  not ginst2801 (P1_R1165_U208, P1_R1165_U30);
  nand ginst2802 (P1_R1165_U209, P1_R1165_U23, P1_R1165_U384);
  not ginst2803 (P1_R1165_U21, P1_U3179);
  nand ginst2804 (P1_R1165_U210, P1_R1165_U21, P1_R1165_U387);
  nand ginst2805 (P1_R1165_U211, P1_R1165_U22, P1_R1165_U23);
  nand ginst2806 (P1_R1165_U212, P1_R1165_U211, P1_R1165_U62);
  nand ginst2807 (P1_R1165_U213, P1_R1165_U194, P1_U3178);
  nand ginst2808 (P1_R1165_U214, P1_R1165_U30, P1_R1165_U4);
  not ginst2809 (P1_R1165_U215, P1_R1165_U153);
  nand ginst2810 (P1_R1165_U216, P1_R1165_U20, P1_R1165_U375);
  nand ginst2811 (P1_R1165_U217, P1_R1165_U26, P1_R1165_U390);
  nand ginst2812 (P1_R1165_U218, P1_R1165_U151, P1_R1165_U217);
  nand ginst2813 (P1_R1165_U219, P1_R1165_U65, P1_U3176);
  nand ginst2814 (P1_R1165_U22, P1_R1165_U61, P1_U3179);
  not ginst2815 (P1_R1165_U220, P1_R1165_U29);
  nand ginst2816 (P1_R1165_U221, P1_R1165_U19, P1_R1165_U393);
  nand ginst2817 (P1_R1165_U222, P1_R1165_U17, P1_R1165_U396);
  not ginst2818 (P1_R1165_U223, P1_R1165_U18);
  nand ginst2819 (P1_R1165_U224, P1_R1165_U18, P1_R1165_U19);
  nand ginst2820 (P1_R1165_U225, P1_R1165_U224, P1_R1165_U59);
  nand ginst2821 (P1_R1165_U226, P1_R1165_U223, P1_U3174);
  nand ginst2822 (P1_R1165_U227, P1_R1165_U29, P1_R1165_U5);
  not ginst2823 (P1_R1165_U228, P1_R1165_U149);
  nand ginst2824 (P1_R1165_U229, P1_R1165_U27, P1_R1165_U399);
  not ginst2825 (P1_R1165_U23, P1_U3178);
  nand ginst2826 (P1_R1165_U230, P1_R1165_U149, P1_R1165_U229);
  nand ginst2827 (P1_R1165_U231, P1_R1165_U66, P1_U3173);
  not ginst2828 (P1_R1165_U232, P1_R1165_U147);
  nand ginst2829 (P1_R1165_U233, P1_R1165_U17, P1_R1165_U396);
  nand ginst2830 (P1_R1165_U234, P1_R1165_U233, P1_R1165_U29);
  nand ginst2831 (P1_R1165_U235, P1_R1165_U111, P1_R1165_U234);
  nand ginst2832 (P1_R1165_U236, P1_R1165_U18, P1_R1165_U220);
  nand ginst2833 (P1_R1165_U237, P1_R1165_U59, P1_U3174);
  nand ginst2834 (P1_R1165_U238, P1_R1165_U112, P1_R1165_U236);
  nand ginst2835 (P1_R1165_U239, P1_R1165_U17, P1_R1165_U396);
  not ginst2836 (P1_R1165_U24, P1_U3181);
  nand ginst2837 (P1_R1165_U240, P1_R1165_U21, P1_R1165_U387);
  nand ginst2838 (P1_R1165_U241, P1_R1165_U240, P1_R1165_U30);
  nand ginst2839 (P1_R1165_U242, P1_R1165_U113, P1_R1165_U241);
  nand ginst2840 (P1_R1165_U243, P1_R1165_U208, P1_R1165_U22);
  nand ginst2841 (P1_R1165_U244, P1_R1165_U62, P1_U3178);
  nand ginst2842 (P1_R1165_U245, P1_R1165_U114, P1_R1165_U243);
  nand ginst2843 (P1_R1165_U246, P1_R1165_U21, P1_R1165_U387);
  nand ginst2844 (P1_R1165_U247, P1_R1165_U28, P1_R1165_U367);
  nand ginst2845 (P1_R1165_U248, P1_R1165_U38, P1_R1165_U451);
  nand ginst2846 (P1_R1165_U249, P1_R1165_U192, P1_R1165_U248);
  not ginst2847 (P1_R1165_U25, P1_U3180);
  nand ginst2848 (P1_R1165_U250, P1_R1165_U73, P1_U3171);
  not ginst2849 (P1_R1165_U251, P1_R1165_U190);
  nand ginst2850 (P1_R1165_U252, P1_R1165_U42, P1_R1165_U454);
  nand ginst2851 (P1_R1165_U253, P1_R1165_U39, P1_R1165_U457);
  nand ginst2852 (P1_R1165_U254, P1_R1165_U198, P1_R1165_U6);
  nand ginst2853 (P1_R1165_U255, P1_R1165_U75, P1_U3168);
  nand ginst2854 (P1_R1165_U256, P1_R1165_U116, P1_R1165_U254);
  nand ginst2855 (P1_R1165_U257, P1_R1165_U40, P1_R1165_U460);
  nand ginst2856 (P1_R1165_U258, P1_R1165_U42, P1_R1165_U454);
  nand ginst2857 (P1_R1165_U259, P1_R1165_U115, P1_R1165_U190);
  not ginst2858 (P1_R1165_U26, P1_U3176);
  nand ginst2859 (P1_R1165_U260, P1_R1165_U256, P1_R1165_U258);
  not ginst2860 (P1_R1165_U261, P1_R1165_U189);
  nand ginst2861 (P1_R1165_U262, P1_R1165_U43, P1_R1165_U463);
  nand ginst2862 (P1_R1165_U263, P1_R1165_U189, P1_R1165_U262);
  nand ginst2863 (P1_R1165_U264, P1_R1165_U77, P1_U3167);
  not ginst2864 (P1_R1165_U265, P1_R1165_U187);
  nand ginst2865 (P1_R1165_U266, P1_R1165_U44, P1_R1165_U466);
  nand ginst2866 (P1_R1165_U267, P1_R1165_U187, P1_R1165_U266);
  nand ginst2867 (P1_R1165_U268, P1_R1165_U78, P1_U3166);
  not ginst2868 (P1_R1165_U269, P1_R1165_U55);
  not ginst2869 (P1_R1165_U27, P1_U3173);
  nand ginst2870 (P1_R1165_U270, P1_R1165_U37, P1_R1165_U469);
  nand ginst2871 (P1_R1165_U271, P1_R1165_U35, P1_R1165_U472);
  not ginst2872 (P1_R1165_U272, P1_R1165_U36);
  nand ginst2873 (P1_R1165_U273, P1_R1165_U36, P1_R1165_U37);
  nand ginst2874 (P1_R1165_U274, P1_R1165_U273, P1_R1165_U72);
  nand ginst2875 (P1_R1165_U275, P1_R1165_U272, P1_U3164);
  nand ginst2876 (P1_R1165_U276, P1_R1165_U55, P1_R1165_U7);
  not ginst2877 (P1_R1165_U277, P1_R1165_U185);
  nand ginst2878 (P1_R1165_U278, P1_R1165_U45, P1_R1165_U475);
  nand ginst2879 (P1_R1165_U279, P1_R1165_U185, P1_R1165_U278);
  not ginst2880 (P1_R1165_U28, P1_U3172);
  nand ginst2881 (P1_R1165_U280, P1_R1165_U79, P1_U3163);
  not ginst2882 (P1_R1165_U281, P1_R1165_U183);
  nand ginst2883 (P1_R1165_U282, P1_R1165_U478, P1_R1165_U49);
  nand ginst2884 (P1_R1165_U283, P1_R1165_U46, P1_R1165_U481);
  nand ginst2885 (P1_R1165_U284, P1_R1165_U199, P1_R1165_U8);
  nand ginst2886 (P1_R1165_U285, P1_R1165_U81, P1_U3160);
  nand ginst2887 (P1_R1165_U286, P1_R1165_U119, P1_R1165_U284);
  nand ginst2888 (P1_R1165_U287, P1_R1165_U47, P1_R1165_U484);
  nand ginst2889 (P1_R1165_U288, P1_R1165_U478, P1_R1165_U49);
  nand ginst2890 (P1_R1165_U289, P1_R1165_U118, P1_R1165_U183);
  nand ginst2891 (P1_R1165_U29, P1_R1165_U218, P1_R1165_U219);
  nand ginst2892 (P1_R1165_U290, P1_R1165_U286, P1_R1165_U288);
  not ginst2893 (P1_R1165_U291, P1_R1165_U180);
  nand ginst2894 (P1_R1165_U292, P1_R1165_U487, P1_R1165_U50);
  nand ginst2895 (P1_R1165_U293, P1_R1165_U180, P1_R1165_U292);
  nand ginst2896 (P1_R1165_U294, P1_R1165_U83, P1_U3159);
  not ginst2897 (P1_R1165_U295, P1_R1165_U178);
  nand ginst2898 (P1_R1165_U296, P1_R1165_U490, P1_R1165_U51);
  nand ginst2899 (P1_R1165_U297, P1_R1165_U178, P1_R1165_U296);
  nand ginst2900 (P1_R1165_U298, P1_R1165_U84, P1_U3158);
  not ginst2901 (P1_R1165_U299, P1_R1165_U176);
  nand ginst2902 (P1_R1165_U30, P1_R1165_U206, P1_R1165_U207);
  nand ginst2903 (P1_R1165_U300, P1_R1165_U33, P1_R1165_U442);
  nand ginst2904 (P1_R1165_U301, P1_R1165_U197, P1_R1165_U200);
  not ginst2905 (P1_R1165_U302, P1_R1165_U52);
  nand ginst2906 (P1_R1165_U303, P1_R1165_U34, P1_R1165_U448);
  nand ginst2907 (P1_R1165_U304, P1_R1165_U176, P1_R1165_U193, P1_R1165_U303);
  not ginst2908 (P1_R1165_U305, P1_R1165_U175);
  nand ginst2909 (P1_R1165_U306, P1_R1165_U31, P1_R1165_U439);
  nand ginst2910 (P1_R1165_U307, P1_R1165_U67, P1_U3154);
  nand ginst2911 (P1_R1165_U308, P1_R1165_U31, P1_R1165_U439);
  nand ginst2912 (P1_R1165_U309, P1_R1165_U176, P1_R1165_U303);
  not ginst2913 (P1_R1165_U31, P1_U3154);
  not ginst2914 (P1_R1165_U310, P1_R1165_U53);
  nand ginst2915 (P1_R1165_U311, P1_R1165_U125, P1_R1165_U9);
  nand ginst2916 (P1_R1165_U312, P1_R1165_U126, P1_R1165_U309);
  nand ginst2917 (P1_R1165_U313, P1_R1165_U69, P1_U3155);
  nand ginst2918 (P1_R1165_U314, P1_R1165_U127, P1_R1165_U312);
  nand ginst2919 (P1_R1165_U315, P1_R1165_U33, P1_R1165_U442);
  nand ginst2920 (P1_R1165_U316, P1_R1165_U183, P1_R1165_U287);
  not ginst2921 (P1_R1165_U317, P1_R1165_U54);
  nand ginst2922 (P1_R1165_U318, P1_R1165_U46, P1_R1165_U481);
  nand ginst2923 (P1_R1165_U319, P1_R1165_U318, P1_R1165_U54);
  not ginst2924 (P1_R1165_U32, P1_U3155);
  nand ginst2925 (P1_R1165_U320, P1_R1165_U129, P1_R1165_U319);
  nand ginst2926 (P1_R1165_U321, P1_R1165_U196, P1_R1165_U317);
  nand ginst2927 (P1_R1165_U322, P1_R1165_U81, P1_U3160);
  nand ginst2928 (P1_R1165_U323, P1_R1165_U130, P1_R1165_U321);
  nand ginst2929 (P1_R1165_U324, P1_R1165_U46, P1_R1165_U481);
  nand ginst2930 (P1_R1165_U325, P1_R1165_U35, P1_R1165_U472);
  nand ginst2931 (P1_R1165_U326, P1_R1165_U325, P1_R1165_U55);
  nand ginst2932 (P1_R1165_U327, P1_R1165_U131, P1_R1165_U326);
  nand ginst2933 (P1_R1165_U328, P1_R1165_U269, P1_R1165_U36);
  nand ginst2934 (P1_R1165_U329, P1_R1165_U72, P1_U3164);
  not ginst2935 (P1_R1165_U33, P1_U3156);
  nand ginst2936 (P1_R1165_U330, P1_R1165_U132, P1_R1165_U328);
  nand ginst2937 (P1_R1165_U331, P1_R1165_U35, P1_R1165_U472);
  nand ginst2938 (P1_R1165_U332, P1_R1165_U190, P1_R1165_U257);
  not ginst2939 (P1_R1165_U333, P1_R1165_U56);
  nand ginst2940 (P1_R1165_U334, P1_R1165_U39, P1_R1165_U457);
  nand ginst2941 (P1_R1165_U335, P1_R1165_U334, P1_R1165_U56);
  nand ginst2942 (P1_R1165_U336, P1_R1165_U133, P1_R1165_U335);
  nand ginst2943 (P1_R1165_U337, P1_R1165_U195, P1_R1165_U333);
  nand ginst2944 (P1_R1165_U338, P1_R1165_U75, P1_U3168);
  nand ginst2945 (P1_R1165_U339, P1_R1165_U134, P1_R1165_U337);
  not ginst2946 (P1_R1165_U34, P1_U3157);
  nand ginst2947 (P1_R1165_U340, P1_R1165_U39, P1_R1165_U457);
  nand ginst2948 (P1_R1165_U341, P1_R1165_U18, P1_R1165_U239);
  nand ginst2949 (P1_R1165_U342, P1_R1165_U22, P1_R1165_U246);
  nand ginst2950 (P1_R1165_U343, P1_R1165_U197, P1_R1165_U315);
  nand ginst2951 (P1_R1165_U344, P1_R1165_U200, P1_R1165_U303);
  nand ginst2952 (P1_R1165_U345, P1_R1165_U196, P1_R1165_U324);
  nand ginst2953 (P1_R1165_U346, P1_R1165_U287, P1_R1165_U48);
  nand ginst2954 (P1_R1165_U347, P1_R1165_U331, P1_R1165_U36);
  nand ginst2955 (P1_R1165_U348, P1_R1165_U195, P1_R1165_U340);
  nand ginst2956 (P1_R1165_U349, P1_R1165_U257, P1_R1165_U41);
  not ginst2957 (P1_R1165_U35, P1_U3165);
  nand ginst2958 (P1_R1165_U350, P1_R1165_U60, P1_U3177);
  nand ginst2959 (P1_R1165_U351, P1_R1165_U120, P1_R1165_U304, P1_R1165_U352);
  nand ginst2960 (P1_R1165_U352, P1_R1165_U193, P1_R1165_U301);
  nand ginst2961 (P1_R1165_U353, P1_R1165_U57, P1_U3172);
  nand ginst2962 (P1_R1165_U354, P1_R1165_U300, P1_R1165_U69);
  nand ginst2963 (P1_R1165_U355, P1_R1165_U300, P1_U3155);
  nand ginst2964 (P1_R1165_U356, P1_R1165_U193, P1_R1165_U301, P1_R1165_U308);
  nand ginst2965 (P1_R1165_U357, P1_R1165_U121, P1_R1165_U176, P1_R1165_U193);
  nand ginst2966 (P1_R1165_U358, P1_R1165_U302, P1_R1165_U308);
  nand ginst2967 (P1_R1165_U359, P1_R1165_U67, P1_U3154);
  nand ginst2968 (P1_R1165_U36, P1_R1165_U71, P1_U3165);
  nand ginst2969 (P1_R1165_U360, P1_R1165_U128, P1_R1165_U310);
  nand ginst2970 (P1_R1165_U361, P1_R1165_U153, P1_R1165_U216);
  not ginst2971 (P1_R1165_U362, P1_R1165_U151);
  nand ginst2972 (P1_R1165_U363, P1_R1165_U147, P1_R1165_U247);
  not ginst2973 (P1_R1165_U364, P1_R1165_U192);
  nand ginst2974 (P1_R1165_U365, P1_R1165_U136, P1_U3211);
  nand ginst2975 (P1_R1165_U366, P1_R1165_U16, P1_U3201);
  not ginst2976 (P1_R1165_U367, P1_R1165_U57);
  nand ginst2977 (P1_R1165_U368, P1_R1165_U367, P1_U3172);
  nand ginst2978 (P1_R1165_U369, P1_R1165_U28, P1_R1165_U57);
  not ginst2979 (P1_R1165_U37, P1_U3164);
  nand ginst2980 (P1_R1165_U370, P1_R1165_U367, P1_U3172);
  nand ginst2981 (P1_R1165_U371, P1_R1165_U28, P1_R1165_U57);
  nand ginst2982 (P1_R1165_U372, P1_R1165_U370, P1_R1165_U371);
  nand ginst2983 (P1_R1165_U373, P1_R1165_U138, P1_U3211);
  nand ginst2984 (P1_R1165_U374, P1_R1165_U16, P1_U3206);
  not ginst2985 (P1_R1165_U375, P1_R1165_U60);
  nand ginst2986 (P1_R1165_U376, P1_R1165_U139, P1_U3211);
  nand ginst2987 (P1_R1165_U377, P1_R1165_U16, P1_U3210);
  not ginst2988 (P1_R1165_U378, P1_R1165_U63);
  nand ginst2989 (P1_R1165_U379, P1_R1165_U140, P1_U3211);
  not ginst2990 (P1_R1165_U38, P1_U3171);
  nand ginst2991 (P1_R1165_U380, P1_R1165_U16, P1_U3209);
  not ginst2992 (P1_R1165_U381, P1_R1165_U64);
  nand ginst2993 (P1_R1165_U382, P1_R1165_U141, P1_U3211);
  nand ginst2994 (P1_R1165_U383, P1_R1165_U16, P1_U3207);
  not ginst2995 (P1_R1165_U384, P1_R1165_U62);
  nand ginst2996 (P1_R1165_U385, P1_R1165_U142, P1_U3211);
  nand ginst2997 (P1_R1165_U386, P1_R1165_U16, P1_U3208);
  not ginst2998 (P1_R1165_U387, P1_R1165_U61);
  nand ginst2999 (P1_R1165_U388, P1_R1165_U143, P1_U3211);
  nand ginst3000 (P1_R1165_U389, P1_R1165_U16, P1_U3205);
  not ginst3001 (P1_R1165_U39, P1_U3169);
  not ginst3002 (P1_R1165_U390, P1_R1165_U65);
  nand ginst3003 (P1_R1165_U391, P1_R1165_U144, P1_U3211);
  nand ginst3004 (P1_R1165_U392, P1_R1165_U16, P1_U3203);
  not ginst3005 (P1_R1165_U393, P1_R1165_U59);
  nand ginst3006 (P1_R1165_U394, P1_R1165_U145, P1_U3211);
  nand ginst3007 (P1_R1165_U395, P1_R1165_U16, P1_U3204);
  not ginst3008 (P1_R1165_U396, P1_R1165_U58);
  nand ginst3009 (P1_R1165_U397, P1_R1165_U146, P1_U3211);
  nand ginst3010 (P1_R1165_U398, P1_R1165_U16, P1_U3202);
  not ginst3011 (P1_R1165_U399, P1_R1165_U66);
  and ginst3012 (P1_R1165_U4, P1_R1165_U209, P1_R1165_U210);
  not ginst3013 (P1_R1165_U40, P1_U3170);
  nand ginst3014 (P1_R1165_U400, P1_R1165_U137, P1_R1165_U147);
  nand ginst3015 (P1_R1165_U401, P1_R1165_U232, P1_R1165_U372);
  nand ginst3016 (P1_R1165_U402, P1_R1165_U399, P1_U3173);
  nand ginst3017 (P1_R1165_U403, P1_R1165_U27, P1_R1165_U66);
  nand ginst3018 (P1_R1165_U404, P1_R1165_U399, P1_U3173);
  nand ginst3019 (P1_R1165_U405, P1_R1165_U27, P1_R1165_U66);
  nand ginst3020 (P1_R1165_U406, P1_R1165_U404, P1_R1165_U405);
  nand ginst3021 (P1_R1165_U407, P1_R1165_U148, P1_R1165_U149);
  nand ginst3022 (P1_R1165_U408, P1_R1165_U228, P1_R1165_U406);
  nand ginst3023 (P1_R1165_U409, P1_R1165_U393, P1_U3174);
  nand ginst3024 (P1_R1165_U41, P1_R1165_U74, P1_U3170);
  nand ginst3025 (P1_R1165_U410, P1_R1165_U19, P1_R1165_U59);
  nand ginst3026 (P1_R1165_U411, P1_R1165_U396, P1_U3175);
  nand ginst3027 (P1_R1165_U412, P1_R1165_U17, P1_R1165_U58);
  nand ginst3028 (P1_R1165_U413, P1_R1165_U411, P1_R1165_U412);
  nand ginst3029 (P1_R1165_U414, P1_R1165_U29, P1_R1165_U341);
  nand ginst3030 (P1_R1165_U415, P1_R1165_U220, P1_R1165_U413);
  nand ginst3031 (P1_R1165_U416, P1_R1165_U390, P1_U3176);
  nand ginst3032 (P1_R1165_U417, P1_R1165_U26, P1_R1165_U65);
  nand ginst3033 (P1_R1165_U418, P1_R1165_U390, P1_U3176);
  nand ginst3034 (P1_R1165_U419, P1_R1165_U26, P1_R1165_U65);
  not ginst3035 (P1_R1165_U42, P1_U3168);
  nand ginst3036 (P1_R1165_U420, P1_R1165_U418, P1_R1165_U419);
  nand ginst3037 (P1_R1165_U421, P1_R1165_U150, P1_R1165_U151);
  nand ginst3038 (P1_R1165_U422, P1_R1165_U362, P1_R1165_U420);
  nand ginst3039 (P1_R1165_U423, P1_R1165_U375, P1_U3177);
  nand ginst3040 (P1_R1165_U424, P1_R1165_U20, P1_R1165_U60);
  nand ginst3041 (P1_R1165_U425, P1_R1165_U375, P1_U3177);
  nand ginst3042 (P1_R1165_U426, P1_R1165_U20, P1_R1165_U60);
  nand ginst3043 (P1_R1165_U427, P1_R1165_U425, P1_R1165_U426);
  nand ginst3044 (P1_R1165_U428, P1_R1165_U152, P1_R1165_U153);
  nand ginst3045 (P1_R1165_U429, P1_R1165_U215, P1_R1165_U427);
  not ginst3046 (P1_R1165_U43, P1_U3167);
  nand ginst3047 (P1_R1165_U430, P1_R1165_U384, P1_U3178);
  nand ginst3048 (P1_R1165_U431, P1_R1165_U23, P1_R1165_U62);
  nand ginst3049 (P1_R1165_U432, P1_R1165_U387, P1_U3179);
  nand ginst3050 (P1_R1165_U433, P1_R1165_U21, P1_R1165_U61);
  nand ginst3051 (P1_R1165_U434, P1_R1165_U432, P1_R1165_U433);
  nand ginst3052 (P1_R1165_U435, P1_R1165_U30, P1_R1165_U342);
  nand ginst3053 (P1_R1165_U436, P1_R1165_U208, P1_R1165_U434);
  nand ginst3054 (P1_R1165_U437, P1_R1165_U154, P1_U3211);
  nand ginst3055 (P1_R1165_U438, P1_R1165_U16, P1_U3183);
  not ginst3056 (P1_R1165_U439, P1_R1165_U67);
  not ginst3057 (P1_R1165_U44, P1_U3166);
  nand ginst3058 (P1_R1165_U440, P1_R1165_U155, P1_U3211);
  nand ginst3059 (P1_R1165_U441, P1_R1165_U16, P1_U3185);
  not ginst3060 (P1_R1165_U442, P1_R1165_U68);
  nand ginst3061 (P1_R1165_U443, P1_R1165_U156, P1_U3211);
  nand ginst3062 (P1_R1165_U444, P1_R1165_U16, P1_U3184);
  not ginst3063 (P1_R1165_U445, P1_R1165_U69);
  nand ginst3064 (P1_R1165_U446, P1_R1165_U157, P1_U3211);
  nand ginst3065 (P1_R1165_U447, P1_R1165_U16, P1_U3186);
  not ginst3066 (P1_R1165_U448, P1_R1165_U70);
  nand ginst3067 (P1_R1165_U449, P1_R1165_U158, P1_U3211);
  not ginst3068 (P1_R1165_U45, P1_U3163);
  nand ginst3069 (P1_R1165_U450, P1_R1165_U16, P1_U3200);
  not ginst3070 (P1_R1165_U451, P1_R1165_U73);
  nand ginst3071 (P1_R1165_U452, P1_R1165_U159, P1_U3211);
  nand ginst3072 (P1_R1165_U453, P1_R1165_U16, P1_U3197);
  not ginst3073 (P1_R1165_U454, P1_R1165_U75);
  nand ginst3074 (P1_R1165_U455, P1_R1165_U160, P1_U3211);
  nand ginst3075 (P1_R1165_U456, P1_R1165_U16, P1_U3198);
  not ginst3076 (P1_R1165_U457, P1_R1165_U76);
  nand ginst3077 (P1_R1165_U458, P1_R1165_U161, P1_U3211);
  nand ginst3078 (P1_R1165_U459, P1_R1165_U16, P1_U3199);
  not ginst3079 (P1_R1165_U46, P1_U3161);
  not ginst3080 (P1_R1165_U460, P1_R1165_U74);
  nand ginst3081 (P1_R1165_U461, P1_R1165_U162, P1_U3211);
  nand ginst3082 (P1_R1165_U462, P1_R1165_U16, P1_U3196);
  not ginst3083 (P1_R1165_U463, P1_R1165_U77);
  nand ginst3084 (P1_R1165_U464, P1_R1165_U163, P1_U3211);
  nand ginst3085 (P1_R1165_U465, P1_R1165_U16, P1_U3195);
  not ginst3086 (P1_R1165_U466, P1_R1165_U78);
  nand ginst3087 (P1_R1165_U467, P1_R1165_U164, P1_U3211);
  nand ginst3088 (P1_R1165_U468, P1_R1165_U16, P1_U3193);
  not ginst3089 (P1_R1165_U469, P1_R1165_U72);
  not ginst3090 (P1_R1165_U47, P1_U3162);
  nand ginst3091 (P1_R1165_U470, P1_R1165_U165, P1_U3211);
  nand ginst3092 (P1_R1165_U471, P1_R1165_U16, P1_U3194);
  not ginst3093 (P1_R1165_U472, P1_R1165_U71);
  nand ginst3094 (P1_R1165_U473, P1_R1165_U166, P1_U3211);
  nand ginst3095 (P1_R1165_U474, P1_R1165_U16, P1_U3192);
  not ginst3096 (P1_R1165_U475, P1_R1165_U79);
  nand ginst3097 (P1_R1165_U476, P1_R1165_U167, P1_U3211);
  nand ginst3098 (P1_R1165_U477, P1_R1165_U16, P1_U3189);
  not ginst3099 (P1_R1165_U478, P1_R1165_U81);
  nand ginst3100 (P1_R1165_U479, P1_R1165_U168, P1_U3211);
  nand ginst3101 (P1_R1165_U48, P1_R1165_U80, P1_U3162);
  nand ginst3102 (P1_R1165_U480, P1_R1165_U16, P1_U3190);
  not ginst3103 (P1_R1165_U481, P1_R1165_U82);
  nand ginst3104 (P1_R1165_U482, P1_R1165_U169, P1_U3211);
  nand ginst3105 (P1_R1165_U483, P1_R1165_U16, P1_U3191);
  not ginst3106 (P1_R1165_U484, P1_R1165_U80);
  nand ginst3107 (P1_R1165_U485, P1_R1165_U170, P1_U3211);
  nand ginst3108 (P1_R1165_U486, P1_R1165_U16, P1_U3188);
  not ginst3109 (P1_R1165_U487, P1_R1165_U83);
  nand ginst3110 (P1_R1165_U488, P1_R1165_U171, P1_U3211);
  nand ginst3111 (P1_R1165_U489, P1_R1165_U16, P1_U3187);
  not ginst3112 (P1_R1165_U49, P1_U3160);
  not ginst3113 (P1_R1165_U490, P1_R1165_U84);
  nand ginst3114 (P1_R1165_U491, P1_R1165_U172, P1_U3211);
  nand ginst3115 (P1_R1165_U492, P1_R1165_U16, P1_U3153);
  not ginst3116 (P1_R1165_U493, P1_R1165_U123);
  nand ginst3117 (P1_R1165_U494, P1_R1165_U493, P1_U3182);
  nand ginst3118 (P1_R1165_U495, P1_R1165_U123, P1_R1165_U173);
  not ginst3119 (P1_R1165_U496, P1_R1165_U85);
  nand ginst3120 (P1_R1165_U497, P1_R1165_U306, P1_R1165_U351, P1_R1165_U496);
  nand ginst3121 (P1_R1165_U498, P1_R1165_U122, P1_R1165_U357, P1_R1165_U358, P1_R1165_U85);
  nand ginst3122 (P1_R1165_U499, P1_R1165_U439, P1_U3154);
  and ginst3123 (P1_R1165_U5, P1_R1165_U221, P1_R1165_U222);
  not ginst3124 (P1_R1165_U50, P1_U3159);
  nand ginst3125 (P1_R1165_U500, P1_R1165_U31, P1_R1165_U67);
  nand ginst3126 (P1_R1165_U501, P1_R1165_U439, P1_U3154);
  nand ginst3127 (P1_R1165_U502, P1_R1165_U31, P1_R1165_U67);
  nand ginst3128 (P1_R1165_U503, P1_R1165_U501, P1_R1165_U502);
  nand ginst3129 (P1_R1165_U504, P1_R1165_U174, P1_R1165_U175);
  nand ginst3130 (P1_R1165_U505, P1_R1165_U305, P1_R1165_U503);
  nand ginst3131 (P1_R1165_U506, P1_R1165_U445, P1_U3155);
  nand ginst3132 (P1_R1165_U507, P1_R1165_U32, P1_R1165_U69);
  nand ginst3133 (P1_R1165_U508, P1_R1165_U442, P1_U3156);
  nand ginst3134 (P1_R1165_U509, P1_R1165_U33, P1_R1165_U68);
  not ginst3135 (P1_R1165_U51, P1_U3158);
  nand ginst3136 (P1_R1165_U510, P1_R1165_U508, P1_R1165_U509);
  nand ginst3137 (P1_R1165_U511, P1_R1165_U343, P1_R1165_U53);
  nand ginst3138 (P1_R1165_U512, P1_R1165_U310, P1_R1165_U510);
  nand ginst3139 (P1_R1165_U513, P1_R1165_U448, P1_U3157);
  nand ginst3140 (P1_R1165_U514, P1_R1165_U34, P1_R1165_U70);
  nand ginst3141 (P1_R1165_U515, P1_R1165_U513, P1_R1165_U514);
  nand ginst3142 (P1_R1165_U516, P1_R1165_U176, P1_R1165_U344);
  nand ginst3143 (P1_R1165_U517, P1_R1165_U299, P1_R1165_U515);
  nand ginst3144 (P1_R1165_U518, P1_R1165_U490, P1_U3158);
  nand ginst3145 (P1_R1165_U519, P1_R1165_U51, P1_R1165_U84);
  nand ginst3146 (P1_R1165_U52, P1_R1165_U69, P1_U3155);
  nand ginst3147 (P1_R1165_U520, P1_R1165_U490, P1_U3158);
  nand ginst3148 (P1_R1165_U521, P1_R1165_U51, P1_R1165_U84);
  nand ginst3149 (P1_R1165_U522, P1_R1165_U520, P1_R1165_U521);
  nand ginst3150 (P1_R1165_U523, P1_R1165_U177, P1_R1165_U178);
  nand ginst3151 (P1_R1165_U524, P1_R1165_U295, P1_R1165_U522);
  nand ginst3152 (P1_R1165_U525, P1_R1165_U487, P1_U3159);
  nand ginst3153 (P1_R1165_U526, P1_R1165_U50, P1_R1165_U83);
  nand ginst3154 (P1_R1165_U527, P1_R1165_U487, P1_U3159);
  nand ginst3155 (P1_R1165_U528, P1_R1165_U50, P1_R1165_U83);
  nand ginst3156 (P1_R1165_U529, P1_R1165_U527, P1_R1165_U528);
  nand ginst3157 (P1_R1165_U53, P1_R1165_U200, P1_R1165_U309);
  nand ginst3158 (P1_R1165_U530, P1_R1165_U179, P1_R1165_U180);
  nand ginst3159 (P1_R1165_U531, P1_R1165_U291, P1_R1165_U529);
  nand ginst3160 (P1_R1165_U532, P1_R1165_U478, P1_U3160);
  nand ginst3161 (P1_R1165_U533, P1_R1165_U49, P1_R1165_U81);
  nand ginst3162 (P1_R1165_U534, P1_R1165_U481, P1_U3161);
  nand ginst3163 (P1_R1165_U535, P1_R1165_U46, P1_R1165_U82);
  nand ginst3164 (P1_R1165_U536, P1_R1165_U534, P1_R1165_U535);
  nand ginst3165 (P1_R1165_U537, P1_R1165_U345, P1_R1165_U54);
  nand ginst3166 (P1_R1165_U538, P1_R1165_U317, P1_R1165_U536);
  nand ginst3167 (P1_R1165_U539, P1_R1165_U381, P1_U3180);
  nand ginst3168 (P1_R1165_U54, P1_R1165_U316, P1_R1165_U48);
  nand ginst3169 (P1_R1165_U540, P1_R1165_U25, P1_R1165_U64);
  nand ginst3170 (P1_R1165_U541, P1_R1165_U381, P1_U3180);
  nand ginst3171 (P1_R1165_U542, P1_R1165_U25, P1_R1165_U64);
  nand ginst3172 (P1_R1165_U543, P1_R1165_U541, P1_R1165_U542);
  nand ginst3173 (P1_R1165_U544, P1_R1165_U181, P1_R1165_U182);
  nand ginst3174 (P1_R1165_U545, P1_R1165_U204, P1_R1165_U543);
  nand ginst3175 (P1_R1165_U546, P1_R1165_U484, P1_U3162);
  nand ginst3176 (P1_R1165_U547, P1_R1165_U47, P1_R1165_U80);
  nand ginst3177 (P1_R1165_U548, P1_R1165_U546, P1_R1165_U547);
  nand ginst3178 (P1_R1165_U549, P1_R1165_U183, P1_R1165_U346);
  nand ginst3179 (P1_R1165_U55, P1_R1165_U267, P1_R1165_U268);
  nand ginst3180 (P1_R1165_U550, P1_R1165_U281, P1_R1165_U548);
  nand ginst3181 (P1_R1165_U551, P1_R1165_U475, P1_U3163);
  nand ginst3182 (P1_R1165_U552, P1_R1165_U45, P1_R1165_U79);
  nand ginst3183 (P1_R1165_U553, P1_R1165_U475, P1_U3163);
  nand ginst3184 (P1_R1165_U554, P1_R1165_U45, P1_R1165_U79);
  nand ginst3185 (P1_R1165_U555, P1_R1165_U553, P1_R1165_U554);
  nand ginst3186 (P1_R1165_U556, P1_R1165_U184, P1_R1165_U185);
  nand ginst3187 (P1_R1165_U557, P1_R1165_U277, P1_R1165_U555);
  nand ginst3188 (P1_R1165_U558, P1_R1165_U469, P1_U3164);
  nand ginst3189 (P1_R1165_U559, P1_R1165_U37, P1_R1165_U72);
  nand ginst3190 (P1_R1165_U56, P1_R1165_U332, P1_R1165_U41);
  nand ginst3191 (P1_R1165_U560, P1_R1165_U472, P1_U3165);
  nand ginst3192 (P1_R1165_U561, P1_R1165_U35, P1_R1165_U71);
  nand ginst3193 (P1_R1165_U562, P1_R1165_U560, P1_R1165_U561);
  nand ginst3194 (P1_R1165_U563, P1_R1165_U347, P1_R1165_U55);
  nand ginst3195 (P1_R1165_U564, P1_R1165_U269, P1_R1165_U562);
  nand ginst3196 (P1_R1165_U565, P1_R1165_U466, P1_U3166);
  nand ginst3197 (P1_R1165_U566, P1_R1165_U44, P1_R1165_U78);
  nand ginst3198 (P1_R1165_U567, P1_R1165_U466, P1_U3166);
  nand ginst3199 (P1_R1165_U568, P1_R1165_U44, P1_R1165_U78);
  nand ginst3200 (P1_R1165_U569, P1_R1165_U567, P1_R1165_U568);
  nand ginst3201 (P1_R1165_U57, P1_R1165_U365, P1_R1165_U366);
  nand ginst3202 (P1_R1165_U570, P1_R1165_U186, P1_R1165_U187);
  nand ginst3203 (P1_R1165_U571, P1_R1165_U265, P1_R1165_U569);
  nand ginst3204 (P1_R1165_U572, P1_R1165_U463, P1_U3167);
  nand ginst3205 (P1_R1165_U573, P1_R1165_U43, P1_R1165_U77);
  nand ginst3206 (P1_R1165_U574, P1_R1165_U463, P1_U3167);
  nand ginst3207 (P1_R1165_U575, P1_R1165_U43, P1_R1165_U77);
  nand ginst3208 (P1_R1165_U576, P1_R1165_U574, P1_R1165_U575);
  nand ginst3209 (P1_R1165_U577, P1_R1165_U188, P1_R1165_U189);
  nand ginst3210 (P1_R1165_U578, P1_R1165_U261, P1_R1165_U576);
  nand ginst3211 (P1_R1165_U579, P1_R1165_U454, P1_U3168);
  nand ginst3212 (P1_R1165_U58, P1_R1165_U394, P1_R1165_U395);
  nand ginst3213 (P1_R1165_U580, P1_R1165_U42, P1_R1165_U75);
  nand ginst3214 (P1_R1165_U581, P1_R1165_U457, P1_U3169);
  nand ginst3215 (P1_R1165_U582, P1_R1165_U39, P1_R1165_U76);
  nand ginst3216 (P1_R1165_U583, P1_R1165_U581, P1_R1165_U582);
  nand ginst3217 (P1_R1165_U584, P1_R1165_U348, P1_R1165_U56);
  nand ginst3218 (P1_R1165_U585, P1_R1165_U333, P1_R1165_U583);
  nand ginst3219 (P1_R1165_U586, P1_R1165_U460, P1_U3170);
  nand ginst3220 (P1_R1165_U587, P1_R1165_U40, P1_R1165_U74);
  nand ginst3221 (P1_R1165_U588, P1_R1165_U586, P1_R1165_U587);
  nand ginst3222 (P1_R1165_U589, P1_R1165_U190, P1_R1165_U349);
  nand ginst3223 (P1_R1165_U59, P1_R1165_U391, P1_R1165_U392);
  nand ginst3224 (P1_R1165_U590, P1_R1165_U251, P1_R1165_U588);
  nand ginst3225 (P1_R1165_U591, P1_R1165_U451, P1_U3171);
  nand ginst3226 (P1_R1165_U592, P1_R1165_U38, P1_R1165_U73);
  nand ginst3227 (P1_R1165_U593, P1_R1165_U451, P1_U3171);
  nand ginst3228 (P1_R1165_U594, P1_R1165_U38, P1_R1165_U73);
  nand ginst3229 (P1_R1165_U595, P1_R1165_U593, P1_R1165_U594);
  nand ginst3230 (P1_R1165_U596, P1_R1165_U191, P1_R1165_U192);
  nand ginst3231 (P1_R1165_U597, P1_R1165_U364, P1_R1165_U595);
  nand ginst3232 (P1_R1165_U598, P1_R1165_U16, P1_U3181);
  nand ginst3233 (P1_R1165_U599, P1_R1165_U24, P1_U3211);
  and ginst3234 (P1_R1165_U6, P1_R1165_U252, P1_R1165_U253);
  nand ginst3235 (P1_R1165_U60, P1_R1165_U373, P1_R1165_U374);
  not ginst3236 (P1_R1165_U600, P1_R1165_U135);
  nand ginst3237 (P1_R1165_U601, P1_R1165_U600, P1_R1165_U63);
  nand ginst3238 (P1_R1165_U602, P1_R1165_U135, P1_R1165_U378);
  nand ginst3239 (P1_R1165_U61, P1_R1165_U385, P1_R1165_U386);
  nand ginst3240 (P1_R1165_U62, P1_R1165_U382, P1_R1165_U383);
  nand ginst3241 (P1_R1165_U63, P1_R1165_U376, P1_R1165_U377);
  nand ginst3242 (P1_R1165_U64, P1_R1165_U379, P1_R1165_U380);
  nand ginst3243 (P1_R1165_U65, P1_R1165_U388, P1_R1165_U389);
  nand ginst3244 (P1_R1165_U66, P1_R1165_U397, P1_R1165_U398);
  nand ginst3245 (P1_R1165_U67, P1_R1165_U437, P1_R1165_U438);
  nand ginst3246 (P1_R1165_U68, P1_R1165_U440, P1_R1165_U441);
  nand ginst3247 (P1_R1165_U69, P1_R1165_U443, P1_R1165_U444);
  and ginst3248 (P1_R1165_U7, P1_R1165_U270, P1_R1165_U271);
  nand ginst3249 (P1_R1165_U70, P1_R1165_U446, P1_R1165_U447);
  nand ginst3250 (P1_R1165_U71, P1_R1165_U470, P1_R1165_U471);
  nand ginst3251 (P1_R1165_U72, P1_R1165_U467, P1_R1165_U468);
  nand ginst3252 (P1_R1165_U73, P1_R1165_U449, P1_R1165_U450);
  nand ginst3253 (P1_R1165_U74, P1_R1165_U458, P1_R1165_U459);
  nand ginst3254 (P1_R1165_U75, P1_R1165_U452, P1_R1165_U453);
  nand ginst3255 (P1_R1165_U76, P1_R1165_U455, P1_R1165_U456);
  nand ginst3256 (P1_R1165_U77, P1_R1165_U461, P1_R1165_U462);
  nand ginst3257 (P1_R1165_U78, P1_R1165_U464, P1_R1165_U465);
  nand ginst3258 (P1_R1165_U79, P1_R1165_U473, P1_R1165_U474);
  and ginst3259 (P1_R1165_U8, P1_R1165_U282, P1_R1165_U283);
  nand ginst3260 (P1_R1165_U80, P1_R1165_U482, P1_R1165_U483);
  nand ginst3261 (P1_R1165_U81, P1_R1165_U476, P1_R1165_U477);
  nand ginst3262 (P1_R1165_U82, P1_R1165_U479, P1_R1165_U480);
  nand ginst3263 (P1_R1165_U83, P1_R1165_U485, P1_R1165_U486);
  nand ginst3264 (P1_R1165_U84, P1_R1165_U488, P1_R1165_U489);
  nand ginst3265 (P1_R1165_U85, P1_R1165_U494, P1_R1165_U495);
  nand ginst3266 (P1_R1165_U86, P1_R1165_U601, P1_R1165_U602);
  nand ginst3267 (P1_R1165_U87, P1_R1165_U400, P1_R1165_U401);
  nand ginst3268 (P1_R1165_U88, P1_R1165_U407, P1_R1165_U408);
  nand ginst3269 (P1_R1165_U89, P1_R1165_U414, P1_R1165_U415);
  and ginst3270 (P1_R1165_U9, P1_R1165_U506, P1_R1165_U507);
  nand ginst3271 (P1_R1165_U90, P1_R1165_U421, P1_R1165_U422);
  nand ginst3272 (P1_R1165_U91, P1_R1165_U428, P1_R1165_U429);
  nand ginst3273 (P1_R1165_U92, P1_R1165_U435, P1_R1165_U436);
  nand ginst3274 (P1_R1165_U93, P1_R1165_U497, P1_R1165_U498);
  nand ginst3275 (P1_R1165_U94, P1_R1165_U504, P1_R1165_U505);
  nand ginst3276 (P1_R1165_U95, P1_R1165_U511, P1_R1165_U512);
  nand ginst3277 (P1_R1165_U96, P1_R1165_U516, P1_R1165_U517);
  nand ginst3278 (P1_R1165_U97, P1_R1165_U523, P1_R1165_U524);
  nand ginst3279 (P1_R1165_U98, P1_R1165_U530, P1_R1165_U531);
  nand ginst3280 (P1_R1165_U99, P1_R1165_U537, P1_R1165_U538);
  and ginst3281 (P1_R1171_U10, P1_R1171_U270, P1_R1171_U271);
  nand ginst3282 (P1_R1171_U100, P1_R1171_U392, P1_R1171_U393);
  nand ginst3283 (P1_R1171_U101, P1_R1171_U397, P1_R1171_U398);
  nand ginst3284 (P1_R1171_U102, P1_R1171_U406, P1_R1171_U407);
  nand ginst3285 (P1_R1171_U103, P1_R1171_U413, P1_R1171_U414);
  nand ginst3286 (P1_R1171_U104, P1_R1171_U420, P1_R1171_U421);
  nand ginst3287 (P1_R1171_U105, P1_R1171_U427, P1_R1171_U428);
  nand ginst3288 (P1_R1171_U106, P1_R1171_U432, P1_R1171_U433);
  nand ginst3289 (P1_R1171_U107, P1_R1171_U439, P1_R1171_U440);
  nand ginst3290 (P1_R1171_U108, P1_R1171_U446, P1_R1171_U447);
  nand ginst3291 (P1_R1171_U109, P1_R1171_U460, P1_R1171_U461);
  and ginst3292 (P1_R1171_U11, P1_R1171_U347, P1_R1171_U350);
  nand ginst3293 (P1_R1171_U110, P1_R1171_U465, P1_R1171_U466);
  nand ginst3294 (P1_R1171_U111, P1_R1171_U472, P1_R1171_U473);
  nand ginst3295 (P1_R1171_U112, P1_R1171_U479, P1_R1171_U480);
  nand ginst3296 (P1_R1171_U113, P1_R1171_U486, P1_R1171_U487);
  nand ginst3297 (P1_R1171_U114, P1_R1171_U493, P1_R1171_U494);
  nand ginst3298 (P1_R1171_U115, P1_R1171_U498, P1_R1171_U499);
  and ginst3299 (P1_R1171_U116, P1_U3068, P1_U3458);
  and ginst3300 (P1_R1171_U117, P1_R1171_U186, P1_R1171_U188);
  and ginst3301 (P1_R1171_U118, P1_R1171_U191, P1_R1171_U193);
  and ginst3302 (P1_R1171_U119, P1_R1171_U199, P1_R1171_U200);
  and ginst3303 (P1_R1171_U12, P1_R1171_U340, P1_R1171_U343);
  and ginst3304 (P1_R1171_U120, P1_R1171_U23, P1_R1171_U380, P1_R1171_U381);
  and ginst3305 (P1_R1171_U121, P1_R1171_U211, P1_R1171_U6);
  and ginst3306 (P1_R1171_U122, P1_R1171_U217, P1_R1171_U219);
  and ginst3307 (P1_R1171_U123, P1_R1171_U35, P1_R1171_U387, P1_R1171_U388);
  and ginst3308 (P1_R1171_U124, P1_R1171_U225, P1_R1171_U4);
  and ginst3309 (P1_R1171_U125, P1_R1171_U180, P1_R1171_U233);
  and ginst3310 (P1_R1171_U126, P1_R1171_U203, P1_R1171_U7);
  and ginst3311 (P1_R1171_U127, P1_R1171_U170, P1_R1171_U238);
  and ginst3312 (P1_R1171_U128, P1_R1171_U249, P1_R1171_U8);
  and ginst3313 (P1_R1171_U129, P1_R1171_U171, P1_R1171_U247);
  and ginst3314 (P1_R1171_U13, P1_R1171_U331, P1_R1171_U334);
  and ginst3315 (P1_R1171_U130, P1_R1171_U266, P1_R1171_U267);
  and ginst3316 (P1_R1171_U131, P1_R1171_U10, P1_R1171_U281);
  and ginst3317 (P1_R1171_U132, P1_R1171_U279, P1_R1171_U284);
  and ginst3318 (P1_R1171_U133, P1_R1171_U297, P1_R1171_U300);
  and ginst3319 (P1_R1171_U134, P1_R1171_U301, P1_R1171_U367);
  and ginst3320 (P1_R1171_U135, P1_R1171_U159, P1_R1171_U277);
  and ginst3321 (P1_R1171_U136, P1_R1171_U453, P1_R1171_U454, P1_R1171_U81);
  and ginst3322 (P1_R1171_U137, P1_R1171_U467, P1_R1171_U468, P1_R1171_U60);
  and ginst3323 (P1_R1171_U138, P1_R1171_U333, P1_R1171_U9);
  and ginst3324 (P1_R1171_U139, P1_R1171_U171, P1_R1171_U488, P1_R1171_U489);
  and ginst3325 (P1_R1171_U14, P1_R1171_U322, P1_R1171_U325);
  and ginst3326 (P1_R1171_U140, P1_R1171_U342, P1_R1171_U8);
  and ginst3327 (P1_R1171_U141, P1_R1171_U170, P1_R1171_U500, P1_R1171_U501);
  and ginst3328 (P1_R1171_U142, P1_R1171_U349, P1_R1171_U7);
  nand ginst3329 (P1_R1171_U143, P1_R1171_U119, P1_R1171_U201);
  nand ginst3330 (P1_R1171_U144, P1_R1171_U216, P1_R1171_U228);
  not ginst3331 (P1_R1171_U145, P1_U3055);
  not ginst3332 (P1_R1171_U146, P1_U3985);
  and ginst3333 (P1_R1171_U147, P1_R1171_U401, P1_R1171_U402);
  nand ginst3334 (P1_R1171_U148, P1_R1171_U168, P1_R1171_U303, P1_R1171_U363);
  and ginst3335 (P1_R1171_U149, P1_R1171_U408, P1_R1171_U409);
  and ginst3336 (P1_R1171_U15, P1_R1171_U317, P1_R1171_U319);
  nand ginst3337 (P1_R1171_U150, P1_R1171_U134, P1_R1171_U368, P1_R1171_U369);
  and ginst3338 (P1_R1171_U151, P1_R1171_U415, P1_R1171_U416);
  nand ginst3339 (P1_R1171_U152, P1_R1171_U298, P1_R1171_U364, P1_R1171_U87);
  and ginst3340 (P1_R1171_U153, P1_R1171_U422, P1_R1171_U423);
  nand ginst3341 (P1_R1171_U154, P1_R1171_U291, P1_R1171_U292);
  and ginst3342 (P1_R1171_U155, P1_R1171_U434, P1_R1171_U435);
  nand ginst3343 (P1_R1171_U156, P1_R1171_U287, P1_R1171_U288);
  and ginst3344 (P1_R1171_U157, P1_R1171_U441, P1_R1171_U442);
  nand ginst3345 (P1_R1171_U158, P1_R1171_U132, P1_R1171_U283);
  and ginst3346 (P1_R1171_U159, P1_R1171_U448, P1_R1171_U449);
  and ginst3347 (P1_R1171_U16, P1_R1171_U309, P1_R1171_U312);
  nand ginst3348 (P1_R1171_U160, P1_R1171_U326, P1_R1171_U44);
  nand ginst3349 (P1_R1171_U161, P1_R1171_U130, P1_R1171_U268);
  and ginst3350 (P1_R1171_U162, P1_R1171_U474, P1_R1171_U475);
  nand ginst3351 (P1_R1171_U163, P1_R1171_U255, P1_R1171_U256);
  and ginst3352 (P1_R1171_U164, P1_R1171_U481, P1_R1171_U482);
  nand ginst3353 (P1_R1171_U165, P1_R1171_U251, P1_R1171_U252);
  nand ginst3354 (P1_R1171_U166, P1_R1171_U241, P1_R1171_U242);
  nand ginst3355 (P1_R1171_U167, P1_R1171_U365, P1_R1171_U366);
  nand ginst3356 (P1_R1171_U168, P1_R1171_U150, P1_U3054);
  not ginst3357 (P1_R1171_U169, P1_R1171_U35);
  and ginst3358 (P1_R1171_U17, P1_R1171_U231, P1_R1171_U234);
  nand ginst3359 (P1_R1171_U170, P1_U3083, P1_U3479);
  nand ginst3360 (P1_R1171_U171, P1_U3072, P1_U3488);
  nand ginst3361 (P1_R1171_U172, P1_U3058, P1_U3977);
  not ginst3362 (P1_R1171_U173, P1_R1171_U69);
  not ginst3363 (P1_R1171_U174, P1_R1171_U78);
  nand ginst3364 (P1_R1171_U175, P1_U3065, P1_U3978);
  not ginst3365 (P1_R1171_U176, P1_R1171_U62);
  or ginst3366 (P1_R1171_U177, P1_U3067, P1_U3467);
  or ginst3367 (P1_R1171_U178, P1_U3060, P1_U3464);
  or ginst3368 (P1_R1171_U179, P1_U3064, P1_U3461);
  and ginst3369 (P1_R1171_U18, P1_R1171_U223, P1_R1171_U226);
  or ginst3370 (P1_R1171_U180, P1_U3068, P1_U3458);
  not ginst3371 (P1_R1171_U181, P1_R1171_U32);
  or ginst3372 (P1_R1171_U182, P1_U3078, P1_U3455);
  not ginst3373 (P1_R1171_U183, P1_R1171_U43);
  not ginst3374 (P1_R1171_U184, P1_R1171_U44);
  nand ginst3375 (P1_R1171_U185, P1_R1171_U43, P1_R1171_U44);
  nand ginst3376 (P1_R1171_U186, P1_R1171_U116, P1_R1171_U179);
  nand ginst3377 (P1_R1171_U187, P1_R1171_U185, P1_R1171_U5);
  nand ginst3378 (P1_R1171_U188, P1_U3064, P1_U3461);
  nand ginst3379 (P1_R1171_U189, P1_R1171_U117, P1_R1171_U187);
  and ginst3380 (P1_R1171_U19, P1_R1171_U209, P1_R1171_U212);
  nand ginst3381 (P1_R1171_U190, P1_R1171_U35, P1_R1171_U36);
  nand ginst3382 (P1_R1171_U191, P1_R1171_U190, P1_U3067);
  nand ginst3383 (P1_R1171_U192, P1_R1171_U189, P1_R1171_U4);
  nand ginst3384 (P1_R1171_U193, P1_R1171_U169, P1_U3467);
  not ginst3385 (P1_R1171_U194, P1_R1171_U42);
  or ginst3386 (P1_R1171_U195, P1_U3070, P1_U3473);
  or ginst3387 (P1_R1171_U196, P1_U3071, P1_U3470);
  not ginst3388 (P1_R1171_U197, P1_R1171_U23);
  nand ginst3389 (P1_R1171_U198, P1_R1171_U23, P1_R1171_U24);
  nand ginst3390 (P1_R1171_U199, P1_R1171_U198, P1_U3070);
  not ginst3391 (P1_R1171_U20, P1_U3470);
  nand ginst3392 (P1_R1171_U200, P1_R1171_U197, P1_U3473);
  nand ginst3393 (P1_R1171_U201, P1_R1171_U42, P1_R1171_U6);
  not ginst3394 (P1_R1171_U202, P1_R1171_U143);
  or ginst3395 (P1_R1171_U203, P1_U3084, P1_U3476);
  nand ginst3396 (P1_R1171_U204, P1_R1171_U143, P1_R1171_U203);
  not ginst3397 (P1_R1171_U205, P1_R1171_U41);
  or ginst3398 (P1_R1171_U206, P1_U3083, P1_U3479);
  or ginst3399 (P1_R1171_U207, P1_U3071, P1_U3470);
  nand ginst3400 (P1_R1171_U208, P1_R1171_U207, P1_R1171_U42);
  nand ginst3401 (P1_R1171_U209, P1_R1171_U120, P1_R1171_U208);
  not ginst3402 (P1_R1171_U21, P1_U3071);
  nand ginst3403 (P1_R1171_U210, P1_R1171_U194, P1_R1171_U23);
  nand ginst3404 (P1_R1171_U211, P1_U3070, P1_U3473);
  nand ginst3405 (P1_R1171_U212, P1_R1171_U121, P1_R1171_U210);
  or ginst3406 (P1_R1171_U213, P1_U3071, P1_U3470);
  nand ginst3407 (P1_R1171_U214, P1_R1171_U180, P1_R1171_U184);
  nand ginst3408 (P1_R1171_U215, P1_U3068, P1_U3458);
  not ginst3409 (P1_R1171_U216, P1_R1171_U46);
  nand ginst3410 (P1_R1171_U217, P1_R1171_U183, P1_R1171_U5);
  nand ginst3411 (P1_R1171_U218, P1_R1171_U179, P1_R1171_U46);
  nand ginst3412 (P1_R1171_U219, P1_U3064, P1_U3461);
  not ginst3413 (P1_R1171_U22, P1_U3070);
  not ginst3414 (P1_R1171_U220, P1_R1171_U45);
  or ginst3415 (P1_R1171_U221, P1_U3060, P1_U3464);
  nand ginst3416 (P1_R1171_U222, P1_R1171_U221, P1_R1171_U45);
  nand ginst3417 (P1_R1171_U223, P1_R1171_U123, P1_R1171_U222);
  nand ginst3418 (P1_R1171_U224, P1_R1171_U220, P1_R1171_U35);
  nand ginst3419 (P1_R1171_U225, P1_U3067, P1_U3467);
  nand ginst3420 (P1_R1171_U226, P1_R1171_U124, P1_R1171_U224);
  or ginst3421 (P1_R1171_U227, P1_U3060, P1_U3464);
  nand ginst3422 (P1_R1171_U228, P1_R1171_U180, P1_R1171_U183);
  not ginst3423 (P1_R1171_U229, P1_R1171_U144);
  nand ginst3424 (P1_R1171_U23, P1_U3071, P1_U3470);
  nand ginst3425 (P1_R1171_U230, P1_U3064, P1_U3461);
  nand ginst3426 (P1_R1171_U231, P1_R1171_U399, P1_R1171_U400, P1_R1171_U43, P1_R1171_U44);
  nand ginst3427 (P1_R1171_U232, P1_R1171_U43, P1_R1171_U44);
  nand ginst3428 (P1_R1171_U233, P1_U3068, P1_U3458);
  nand ginst3429 (P1_R1171_U234, P1_R1171_U125, P1_R1171_U232);
  or ginst3430 (P1_R1171_U235, P1_U3083, P1_U3479);
  or ginst3431 (P1_R1171_U236, P1_U3062, P1_U3482);
  nand ginst3432 (P1_R1171_U237, P1_R1171_U176, P1_R1171_U7);
  nand ginst3433 (P1_R1171_U238, P1_U3062, P1_U3482);
  nand ginst3434 (P1_R1171_U239, P1_R1171_U127, P1_R1171_U237);
  not ginst3435 (P1_R1171_U24, P1_U3473);
  or ginst3436 (P1_R1171_U240, P1_U3062, P1_U3482);
  nand ginst3437 (P1_R1171_U241, P1_R1171_U126, P1_R1171_U143);
  nand ginst3438 (P1_R1171_U242, P1_R1171_U239, P1_R1171_U240);
  not ginst3439 (P1_R1171_U243, P1_R1171_U166);
  or ginst3440 (P1_R1171_U244, P1_U3080, P1_U3491);
  or ginst3441 (P1_R1171_U245, P1_U3072, P1_U3488);
  nand ginst3442 (P1_R1171_U246, P1_R1171_U173, P1_R1171_U8);
  nand ginst3443 (P1_R1171_U247, P1_U3080, P1_U3491);
  nand ginst3444 (P1_R1171_U248, P1_R1171_U129, P1_R1171_U246);
  or ginst3445 (P1_R1171_U249, P1_U3063, P1_U3485);
  not ginst3446 (P1_R1171_U25, P1_U3464);
  or ginst3447 (P1_R1171_U250, P1_U3080, P1_U3491);
  nand ginst3448 (P1_R1171_U251, P1_R1171_U128, P1_R1171_U166);
  nand ginst3449 (P1_R1171_U252, P1_R1171_U248, P1_R1171_U250);
  not ginst3450 (P1_R1171_U253, P1_R1171_U165);
  or ginst3451 (P1_R1171_U254, P1_U3079, P1_U3494);
  nand ginst3452 (P1_R1171_U255, P1_R1171_U165, P1_R1171_U254);
  nand ginst3453 (P1_R1171_U256, P1_U3079, P1_U3494);
  not ginst3454 (P1_R1171_U257, P1_R1171_U163);
  or ginst3455 (P1_R1171_U258, P1_U3074, P1_U3497);
  nand ginst3456 (P1_R1171_U259, P1_R1171_U163, P1_R1171_U258);
  not ginst3457 (P1_R1171_U26, P1_U3060);
  nand ginst3458 (P1_R1171_U260, P1_U3074, P1_U3497);
  not ginst3459 (P1_R1171_U261, P1_R1171_U93);
  or ginst3460 (P1_R1171_U262, P1_U3069, P1_U3503);
  or ginst3461 (P1_R1171_U263, P1_U3073, P1_U3500);
  not ginst3462 (P1_R1171_U264, P1_R1171_U60);
  nand ginst3463 (P1_R1171_U265, P1_R1171_U60, P1_R1171_U61);
  nand ginst3464 (P1_R1171_U266, P1_R1171_U265, P1_U3069);
  nand ginst3465 (P1_R1171_U267, P1_R1171_U264, P1_U3503);
  nand ginst3466 (P1_R1171_U268, P1_R1171_U9, P1_R1171_U93);
  not ginst3467 (P1_R1171_U269, P1_R1171_U161);
  not ginst3468 (P1_R1171_U27, P1_U3067);
  or ginst3469 (P1_R1171_U270, P1_U3076, P1_U3982);
  or ginst3470 (P1_R1171_U271, P1_U3081, P1_U3508);
  or ginst3471 (P1_R1171_U272, P1_U3075, P1_U3981);
  not ginst3472 (P1_R1171_U273, P1_R1171_U81);
  nand ginst3473 (P1_R1171_U274, P1_R1171_U273, P1_U3982);
  nand ginst3474 (P1_R1171_U275, P1_R1171_U274, P1_R1171_U91);
  nand ginst3475 (P1_R1171_U276, P1_R1171_U81, P1_R1171_U82);
  nand ginst3476 (P1_R1171_U277, P1_R1171_U275, P1_R1171_U276);
  nand ginst3477 (P1_R1171_U278, P1_R1171_U10, P1_R1171_U174);
  nand ginst3478 (P1_R1171_U279, P1_U3075, P1_U3981);
  not ginst3479 (P1_R1171_U28, P1_U3458);
  nand ginst3480 (P1_R1171_U280, P1_R1171_U277, P1_R1171_U278);
  or ginst3481 (P1_R1171_U281, P1_U3082, P1_U3506);
  or ginst3482 (P1_R1171_U282, P1_U3075, P1_U3981);
  nand ginst3483 (P1_R1171_U283, P1_R1171_U131, P1_R1171_U161, P1_R1171_U272);
  nand ginst3484 (P1_R1171_U284, P1_R1171_U280, P1_R1171_U282);
  not ginst3485 (P1_R1171_U285, P1_R1171_U158);
  or ginst3486 (P1_R1171_U286, P1_U3061, P1_U3980);
  nand ginst3487 (P1_R1171_U287, P1_R1171_U158, P1_R1171_U286);
  nand ginst3488 (P1_R1171_U288, P1_U3061, P1_U3980);
  not ginst3489 (P1_R1171_U289, P1_R1171_U156);
  not ginst3490 (P1_R1171_U29, P1_U3068);
  or ginst3491 (P1_R1171_U290, P1_U3066, P1_U3979);
  nand ginst3492 (P1_R1171_U291, P1_R1171_U156, P1_R1171_U290);
  nand ginst3493 (P1_R1171_U292, P1_U3066, P1_U3979);
  not ginst3494 (P1_R1171_U293, P1_R1171_U154);
  or ginst3495 (P1_R1171_U294, P1_U3058, P1_U3977);
  nand ginst3496 (P1_R1171_U295, P1_R1171_U172, P1_R1171_U175);
  not ginst3497 (P1_R1171_U296, P1_R1171_U87);
  or ginst3498 (P1_R1171_U297, P1_U3065, P1_U3978);
  nand ginst3499 (P1_R1171_U298, P1_R1171_U154, P1_R1171_U167, P1_R1171_U297);
  not ginst3500 (P1_R1171_U299, P1_R1171_U152);
  not ginst3501 (P1_R1171_U30, P1_U3450);
  or ginst3502 (P1_R1171_U300, P1_U3053, P1_U3975);
  nand ginst3503 (P1_R1171_U301, P1_U3053, P1_U3975);
  not ginst3504 (P1_R1171_U302, P1_R1171_U150);
  nand ginst3505 (P1_R1171_U303, P1_R1171_U150, P1_U3974);
  not ginst3506 (P1_R1171_U304, P1_R1171_U148);
  nand ginst3507 (P1_R1171_U305, P1_R1171_U154, P1_R1171_U297);
  not ginst3508 (P1_R1171_U306, P1_R1171_U90);
  or ginst3509 (P1_R1171_U307, P1_U3058, P1_U3977);
  nand ginst3510 (P1_R1171_U308, P1_R1171_U307, P1_R1171_U90);
  nand ginst3511 (P1_R1171_U309, P1_R1171_U153, P1_R1171_U172, P1_R1171_U308);
  not ginst3512 (P1_R1171_U31, P1_U3077);
  nand ginst3513 (P1_R1171_U310, P1_R1171_U172, P1_R1171_U306);
  nand ginst3514 (P1_R1171_U311, P1_U3057, P1_U3976);
  nand ginst3515 (P1_R1171_U312, P1_R1171_U167, P1_R1171_U310, P1_R1171_U311);
  or ginst3516 (P1_R1171_U313, P1_U3058, P1_U3977);
  nand ginst3517 (P1_R1171_U314, P1_R1171_U161, P1_R1171_U281);
  not ginst3518 (P1_R1171_U315, P1_R1171_U92);
  nand ginst3519 (P1_R1171_U316, P1_R1171_U10, P1_R1171_U92);
  nand ginst3520 (P1_R1171_U317, P1_R1171_U135, P1_R1171_U316);
  nand ginst3521 (P1_R1171_U318, P1_R1171_U277, P1_R1171_U316);
  nand ginst3522 (P1_R1171_U319, P1_R1171_U318, P1_R1171_U452);
  nand ginst3523 (P1_R1171_U32, P1_U3077, P1_U3450);
  or ginst3524 (P1_R1171_U320, P1_U3081, P1_U3508);
  nand ginst3525 (P1_R1171_U321, P1_R1171_U320, P1_R1171_U92);
  nand ginst3526 (P1_R1171_U322, P1_R1171_U136, P1_R1171_U321);
  nand ginst3527 (P1_R1171_U323, P1_R1171_U315, P1_R1171_U81);
  nand ginst3528 (P1_R1171_U324, P1_U3076, P1_U3982);
  nand ginst3529 (P1_R1171_U325, P1_R1171_U10, P1_R1171_U323, P1_R1171_U324);
  or ginst3530 (P1_R1171_U326, P1_U3078, P1_U3455);
  not ginst3531 (P1_R1171_U327, P1_R1171_U160);
  or ginst3532 (P1_R1171_U328, P1_U3081, P1_U3508);
  or ginst3533 (P1_R1171_U329, P1_U3073, P1_U3500);
  not ginst3534 (P1_R1171_U33, P1_U3461);
  nand ginst3535 (P1_R1171_U330, P1_R1171_U329, P1_R1171_U93);
  nand ginst3536 (P1_R1171_U331, P1_R1171_U137, P1_R1171_U330);
  nand ginst3537 (P1_R1171_U332, P1_R1171_U261, P1_R1171_U60);
  nand ginst3538 (P1_R1171_U333, P1_U3069, P1_U3503);
  nand ginst3539 (P1_R1171_U334, P1_R1171_U138, P1_R1171_U332);
  or ginst3540 (P1_R1171_U335, P1_U3073, P1_U3500);
  nand ginst3541 (P1_R1171_U336, P1_R1171_U166, P1_R1171_U249);
  not ginst3542 (P1_R1171_U337, P1_R1171_U94);
  or ginst3543 (P1_R1171_U338, P1_U3072, P1_U3488);
  nand ginst3544 (P1_R1171_U339, P1_R1171_U338, P1_R1171_U94);
  not ginst3545 (P1_R1171_U34, P1_U3064);
  nand ginst3546 (P1_R1171_U340, P1_R1171_U139, P1_R1171_U339);
  nand ginst3547 (P1_R1171_U341, P1_R1171_U171, P1_R1171_U337);
  nand ginst3548 (P1_R1171_U342, P1_U3080, P1_U3491);
  nand ginst3549 (P1_R1171_U343, P1_R1171_U140, P1_R1171_U341);
  or ginst3550 (P1_R1171_U344, P1_U3072, P1_U3488);
  or ginst3551 (P1_R1171_U345, P1_U3083, P1_U3479);
  nand ginst3552 (P1_R1171_U346, P1_R1171_U345, P1_R1171_U41);
  nand ginst3553 (P1_R1171_U347, P1_R1171_U141, P1_R1171_U346);
  nand ginst3554 (P1_R1171_U348, P1_R1171_U170, P1_R1171_U205);
  nand ginst3555 (P1_R1171_U349, P1_U3062, P1_U3482);
  nand ginst3556 (P1_R1171_U35, P1_U3060, P1_U3464);
  nand ginst3557 (P1_R1171_U350, P1_R1171_U142, P1_R1171_U348);
  nand ginst3558 (P1_R1171_U351, P1_R1171_U170, P1_R1171_U206);
  nand ginst3559 (P1_R1171_U352, P1_R1171_U203, P1_R1171_U62);
  nand ginst3560 (P1_R1171_U353, P1_R1171_U213, P1_R1171_U23);
  nand ginst3561 (P1_R1171_U354, P1_R1171_U227, P1_R1171_U35);
  nand ginst3562 (P1_R1171_U355, P1_R1171_U179, P1_R1171_U230);
  nand ginst3563 (P1_R1171_U356, P1_R1171_U172, P1_R1171_U313);
  nand ginst3564 (P1_R1171_U357, P1_R1171_U175, P1_R1171_U297);
  nand ginst3565 (P1_R1171_U358, P1_R1171_U328, P1_R1171_U81);
  nand ginst3566 (P1_R1171_U359, P1_R1171_U281, P1_R1171_U78);
  not ginst3567 (P1_R1171_U36, P1_U3467);
  nand ginst3568 (P1_R1171_U360, P1_R1171_U335, P1_R1171_U60);
  nand ginst3569 (P1_R1171_U361, P1_R1171_U171, P1_R1171_U344);
  nand ginst3570 (P1_R1171_U362, P1_R1171_U249, P1_R1171_U69);
  nand ginst3571 (P1_R1171_U363, P1_U3054, P1_U3974);
  nand ginst3572 (P1_R1171_U364, P1_R1171_U167, P1_R1171_U295);
  nand ginst3573 (P1_R1171_U365, P1_R1171_U294, P1_U3057);
  nand ginst3574 (P1_R1171_U366, P1_R1171_U294, P1_U3976);
  nand ginst3575 (P1_R1171_U367, P1_R1171_U167, P1_R1171_U295, P1_R1171_U300);
  nand ginst3576 (P1_R1171_U368, P1_R1171_U133, P1_R1171_U154, P1_R1171_U167);
  nand ginst3577 (P1_R1171_U369, P1_R1171_U296, P1_R1171_U300);
  not ginst3578 (P1_R1171_U37, P1_U3476);
  nand ginst3579 (P1_R1171_U370, P1_R1171_U40, P1_U3083);
  nand ginst3580 (P1_R1171_U371, P1_R1171_U39, P1_U3479);
  nand ginst3581 (P1_R1171_U372, P1_R1171_U370, P1_R1171_U371);
  nand ginst3582 (P1_R1171_U373, P1_R1171_U351, P1_R1171_U41);
  nand ginst3583 (P1_R1171_U374, P1_R1171_U205, P1_R1171_U372);
  nand ginst3584 (P1_R1171_U375, P1_R1171_U37, P1_U3084);
  nand ginst3585 (P1_R1171_U376, P1_R1171_U38, P1_U3476);
  nand ginst3586 (P1_R1171_U377, P1_R1171_U375, P1_R1171_U376);
  nand ginst3587 (P1_R1171_U378, P1_R1171_U143, P1_R1171_U352);
  nand ginst3588 (P1_R1171_U379, P1_R1171_U202, P1_R1171_U377);
  not ginst3589 (P1_R1171_U38, P1_U3084);
  nand ginst3590 (P1_R1171_U380, P1_R1171_U24, P1_U3070);
  nand ginst3591 (P1_R1171_U381, P1_R1171_U22, P1_U3473);
  nand ginst3592 (P1_R1171_U382, P1_R1171_U20, P1_U3071);
  nand ginst3593 (P1_R1171_U383, P1_R1171_U21, P1_U3470);
  nand ginst3594 (P1_R1171_U384, P1_R1171_U382, P1_R1171_U383);
  nand ginst3595 (P1_R1171_U385, P1_R1171_U353, P1_R1171_U42);
  nand ginst3596 (P1_R1171_U386, P1_R1171_U194, P1_R1171_U384);
  nand ginst3597 (P1_R1171_U387, P1_R1171_U36, P1_U3067);
  nand ginst3598 (P1_R1171_U388, P1_R1171_U27, P1_U3467);
  nand ginst3599 (P1_R1171_U389, P1_R1171_U25, P1_U3060);
  not ginst3600 (P1_R1171_U39, P1_U3083);
  nand ginst3601 (P1_R1171_U390, P1_R1171_U26, P1_U3464);
  nand ginst3602 (P1_R1171_U391, P1_R1171_U389, P1_R1171_U390);
  nand ginst3603 (P1_R1171_U392, P1_R1171_U354, P1_R1171_U45);
  nand ginst3604 (P1_R1171_U393, P1_R1171_U220, P1_R1171_U391);
  nand ginst3605 (P1_R1171_U394, P1_R1171_U33, P1_U3064);
  nand ginst3606 (P1_R1171_U395, P1_R1171_U34, P1_U3461);
  nand ginst3607 (P1_R1171_U396, P1_R1171_U394, P1_R1171_U395);
  nand ginst3608 (P1_R1171_U397, P1_R1171_U144, P1_R1171_U355);
  nand ginst3609 (P1_R1171_U398, P1_R1171_U229, P1_R1171_U396);
  nand ginst3610 (P1_R1171_U399, P1_R1171_U28, P1_U3068);
  and ginst3611 (P1_R1171_U4, P1_R1171_U177, P1_R1171_U178);
  not ginst3612 (P1_R1171_U40, P1_U3479);
  nand ginst3613 (P1_R1171_U400, P1_R1171_U29, P1_U3458);
  nand ginst3614 (P1_R1171_U401, P1_R1171_U146, P1_U3055);
  nand ginst3615 (P1_R1171_U402, P1_R1171_U145, P1_U3985);
  nand ginst3616 (P1_R1171_U403, P1_R1171_U146, P1_U3055);
  nand ginst3617 (P1_R1171_U404, P1_R1171_U145, P1_U3985);
  nand ginst3618 (P1_R1171_U405, P1_R1171_U403, P1_R1171_U404);
  nand ginst3619 (P1_R1171_U406, P1_R1171_U147, P1_R1171_U148);
  nand ginst3620 (P1_R1171_U407, P1_R1171_U304, P1_R1171_U405);
  nand ginst3621 (P1_R1171_U408, P1_R1171_U89, P1_U3054);
  nand ginst3622 (P1_R1171_U409, P1_R1171_U88, P1_U3974);
  nand ginst3623 (P1_R1171_U41, P1_R1171_U204, P1_R1171_U62);
  nand ginst3624 (P1_R1171_U410, P1_R1171_U89, P1_U3054);
  nand ginst3625 (P1_R1171_U411, P1_R1171_U88, P1_U3974);
  nand ginst3626 (P1_R1171_U412, P1_R1171_U410, P1_R1171_U411);
  nand ginst3627 (P1_R1171_U413, P1_R1171_U149, P1_R1171_U150);
  nand ginst3628 (P1_R1171_U414, P1_R1171_U302, P1_R1171_U412);
  nand ginst3629 (P1_R1171_U415, P1_R1171_U47, P1_U3053);
  nand ginst3630 (P1_R1171_U416, P1_R1171_U48, P1_U3975);
  nand ginst3631 (P1_R1171_U417, P1_R1171_U47, P1_U3053);
  nand ginst3632 (P1_R1171_U418, P1_R1171_U48, P1_U3975);
  nand ginst3633 (P1_R1171_U419, P1_R1171_U417, P1_R1171_U418);
  nand ginst3634 (P1_R1171_U42, P1_R1171_U118, P1_R1171_U192);
  nand ginst3635 (P1_R1171_U420, P1_R1171_U151, P1_R1171_U152);
  nand ginst3636 (P1_R1171_U421, P1_R1171_U299, P1_R1171_U419);
  nand ginst3637 (P1_R1171_U422, P1_R1171_U50, P1_U3057);
  nand ginst3638 (P1_R1171_U423, P1_R1171_U49, P1_U3976);
  nand ginst3639 (P1_R1171_U424, P1_R1171_U51, P1_U3058);
  nand ginst3640 (P1_R1171_U425, P1_R1171_U52, P1_U3977);
  nand ginst3641 (P1_R1171_U426, P1_R1171_U424, P1_R1171_U425);
  nand ginst3642 (P1_R1171_U427, P1_R1171_U356, P1_R1171_U90);
  nand ginst3643 (P1_R1171_U428, P1_R1171_U306, P1_R1171_U426);
  nand ginst3644 (P1_R1171_U429, P1_R1171_U53, P1_U3065);
  nand ginst3645 (P1_R1171_U43, P1_R1171_U181, P1_R1171_U182);
  nand ginst3646 (P1_R1171_U430, P1_R1171_U54, P1_U3978);
  nand ginst3647 (P1_R1171_U431, P1_R1171_U429, P1_R1171_U430);
  nand ginst3648 (P1_R1171_U432, P1_R1171_U154, P1_R1171_U357);
  nand ginst3649 (P1_R1171_U433, P1_R1171_U293, P1_R1171_U431);
  nand ginst3650 (P1_R1171_U434, P1_R1171_U85, P1_U3066);
  nand ginst3651 (P1_R1171_U435, P1_R1171_U86, P1_U3979);
  nand ginst3652 (P1_R1171_U436, P1_R1171_U85, P1_U3066);
  nand ginst3653 (P1_R1171_U437, P1_R1171_U86, P1_U3979);
  nand ginst3654 (P1_R1171_U438, P1_R1171_U436, P1_R1171_U437);
  nand ginst3655 (P1_R1171_U439, P1_R1171_U155, P1_R1171_U156);
  nand ginst3656 (P1_R1171_U44, P1_U3078, P1_U3455);
  nand ginst3657 (P1_R1171_U440, P1_R1171_U289, P1_R1171_U438);
  nand ginst3658 (P1_R1171_U441, P1_R1171_U83, P1_U3061);
  nand ginst3659 (P1_R1171_U442, P1_R1171_U84, P1_U3980);
  nand ginst3660 (P1_R1171_U443, P1_R1171_U83, P1_U3061);
  nand ginst3661 (P1_R1171_U444, P1_R1171_U84, P1_U3980);
  nand ginst3662 (P1_R1171_U445, P1_R1171_U443, P1_R1171_U444);
  nand ginst3663 (P1_R1171_U446, P1_R1171_U157, P1_R1171_U158);
  nand ginst3664 (P1_R1171_U447, P1_R1171_U285, P1_R1171_U445);
  nand ginst3665 (P1_R1171_U448, P1_R1171_U55, P1_U3075);
  nand ginst3666 (P1_R1171_U449, P1_R1171_U56, P1_U3981);
  nand ginst3667 (P1_R1171_U45, P1_R1171_U122, P1_R1171_U218);
  nand ginst3668 (P1_R1171_U450, P1_R1171_U55, P1_U3075);
  nand ginst3669 (P1_R1171_U451, P1_R1171_U56, P1_U3981);
  nand ginst3670 (P1_R1171_U452, P1_R1171_U450, P1_R1171_U451);
  nand ginst3671 (P1_R1171_U453, P1_R1171_U82, P1_U3076);
  nand ginst3672 (P1_R1171_U454, P1_R1171_U91, P1_U3982);
  nand ginst3673 (P1_R1171_U455, P1_R1171_U160, P1_R1171_U181);
  nand ginst3674 (P1_R1171_U456, P1_R1171_U32, P1_R1171_U327);
  nand ginst3675 (P1_R1171_U457, P1_R1171_U79, P1_U3081);
  nand ginst3676 (P1_R1171_U458, P1_R1171_U80, P1_U3508);
  nand ginst3677 (P1_R1171_U459, P1_R1171_U457, P1_R1171_U458);
  nand ginst3678 (P1_R1171_U46, P1_R1171_U214, P1_R1171_U215);
  nand ginst3679 (P1_R1171_U460, P1_R1171_U358, P1_R1171_U92);
  nand ginst3680 (P1_R1171_U461, P1_R1171_U315, P1_R1171_U459);
  nand ginst3681 (P1_R1171_U462, P1_R1171_U76, P1_U3082);
  nand ginst3682 (P1_R1171_U463, P1_R1171_U77, P1_U3506);
  nand ginst3683 (P1_R1171_U464, P1_R1171_U462, P1_R1171_U463);
  nand ginst3684 (P1_R1171_U465, P1_R1171_U161, P1_R1171_U359);
  nand ginst3685 (P1_R1171_U466, P1_R1171_U269, P1_R1171_U464);
  nand ginst3686 (P1_R1171_U467, P1_R1171_U61, P1_U3069);
  nand ginst3687 (P1_R1171_U468, P1_R1171_U59, P1_U3503);
  nand ginst3688 (P1_R1171_U469, P1_R1171_U57, P1_U3073);
  not ginst3689 (P1_R1171_U47, P1_U3975);
  nand ginst3690 (P1_R1171_U470, P1_R1171_U58, P1_U3500);
  nand ginst3691 (P1_R1171_U471, P1_R1171_U469, P1_R1171_U470);
  nand ginst3692 (P1_R1171_U472, P1_R1171_U360, P1_R1171_U93);
  nand ginst3693 (P1_R1171_U473, P1_R1171_U261, P1_R1171_U471);
  nand ginst3694 (P1_R1171_U474, P1_R1171_U74, P1_U3074);
  nand ginst3695 (P1_R1171_U475, P1_R1171_U75, P1_U3497);
  nand ginst3696 (P1_R1171_U476, P1_R1171_U74, P1_U3074);
  nand ginst3697 (P1_R1171_U477, P1_R1171_U75, P1_U3497);
  nand ginst3698 (P1_R1171_U478, P1_R1171_U476, P1_R1171_U477);
  nand ginst3699 (P1_R1171_U479, P1_R1171_U162, P1_R1171_U163);
  not ginst3700 (P1_R1171_U48, P1_U3053);
  nand ginst3701 (P1_R1171_U480, P1_R1171_U257, P1_R1171_U478);
  nand ginst3702 (P1_R1171_U481, P1_R1171_U72, P1_U3079);
  nand ginst3703 (P1_R1171_U482, P1_R1171_U73, P1_U3494);
  nand ginst3704 (P1_R1171_U483, P1_R1171_U72, P1_U3079);
  nand ginst3705 (P1_R1171_U484, P1_R1171_U73, P1_U3494);
  nand ginst3706 (P1_R1171_U485, P1_R1171_U483, P1_R1171_U484);
  nand ginst3707 (P1_R1171_U486, P1_R1171_U164, P1_R1171_U165);
  nand ginst3708 (P1_R1171_U487, P1_R1171_U253, P1_R1171_U485);
  nand ginst3709 (P1_R1171_U488, P1_R1171_U70, P1_U3080);
  nand ginst3710 (P1_R1171_U489, P1_R1171_U71, P1_U3491);
  not ginst3711 (P1_R1171_U49, P1_U3057);
  nand ginst3712 (P1_R1171_U490, P1_R1171_U65, P1_U3072);
  nand ginst3713 (P1_R1171_U491, P1_R1171_U66, P1_U3488);
  nand ginst3714 (P1_R1171_U492, P1_R1171_U490, P1_R1171_U491);
  nand ginst3715 (P1_R1171_U493, P1_R1171_U361, P1_R1171_U94);
  nand ginst3716 (P1_R1171_U494, P1_R1171_U337, P1_R1171_U492);
  nand ginst3717 (P1_R1171_U495, P1_R1171_U67, P1_U3063);
  nand ginst3718 (P1_R1171_U496, P1_R1171_U68, P1_U3485);
  nand ginst3719 (P1_R1171_U497, P1_R1171_U495, P1_R1171_U496);
  nand ginst3720 (P1_R1171_U498, P1_R1171_U166, P1_R1171_U362);
  nand ginst3721 (P1_R1171_U499, P1_R1171_U243, P1_R1171_U497);
  and ginst3722 (P1_R1171_U5, P1_R1171_U179, P1_R1171_U180);
  not ginst3723 (P1_R1171_U50, P1_U3976);
  nand ginst3724 (P1_R1171_U500, P1_R1171_U63, P1_U3062);
  nand ginst3725 (P1_R1171_U501, P1_R1171_U64, P1_U3482);
  nand ginst3726 (P1_R1171_U502, P1_R1171_U30, P1_U3077);
  nand ginst3727 (P1_R1171_U503, P1_R1171_U31, P1_U3450);
  not ginst3728 (P1_R1171_U51, P1_U3977);
  not ginst3729 (P1_R1171_U52, P1_U3058);
  not ginst3730 (P1_R1171_U53, P1_U3978);
  not ginst3731 (P1_R1171_U54, P1_U3065);
  not ginst3732 (P1_R1171_U55, P1_U3981);
  not ginst3733 (P1_R1171_U56, P1_U3075);
  not ginst3734 (P1_R1171_U57, P1_U3500);
  not ginst3735 (P1_R1171_U58, P1_U3073);
  not ginst3736 (P1_R1171_U59, P1_U3069);
  and ginst3737 (P1_R1171_U6, P1_R1171_U195, P1_R1171_U196);
  nand ginst3738 (P1_R1171_U60, P1_U3073, P1_U3500);
  not ginst3739 (P1_R1171_U61, P1_U3503);
  nand ginst3740 (P1_R1171_U62, P1_U3084, P1_U3476);
  not ginst3741 (P1_R1171_U63, P1_U3482);
  not ginst3742 (P1_R1171_U64, P1_U3062);
  not ginst3743 (P1_R1171_U65, P1_U3488);
  not ginst3744 (P1_R1171_U66, P1_U3072);
  not ginst3745 (P1_R1171_U67, P1_U3485);
  not ginst3746 (P1_R1171_U68, P1_U3063);
  nand ginst3747 (P1_R1171_U69, P1_U3063, P1_U3485);
  and ginst3748 (P1_R1171_U7, P1_R1171_U235, P1_R1171_U236);
  not ginst3749 (P1_R1171_U70, P1_U3491);
  not ginst3750 (P1_R1171_U71, P1_U3080);
  not ginst3751 (P1_R1171_U72, P1_U3494);
  not ginst3752 (P1_R1171_U73, P1_U3079);
  not ginst3753 (P1_R1171_U74, P1_U3497);
  not ginst3754 (P1_R1171_U75, P1_U3074);
  not ginst3755 (P1_R1171_U76, P1_U3506);
  not ginst3756 (P1_R1171_U77, P1_U3082);
  nand ginst3757 (P1_R1171_U78, P1_U3082, P1_U3506);
  not ginst3758 (P1_R1171_U79, P1_U3508);
  and ginst3759 (P1_R1171_U8, P1_R1171_U244, P1_R1171_U245);
  not ginst3760 (P1_R1171_U80, P1_U3081);
  nand ginst3761 (P1_R1171_U81, P1_U3081, P1_U3508);
  not ginst3762 (P1_R1171_U82, P1_U3982);
  not ginst3763 (P1_R1171_U83, P1_U3980);
  not ginst3764 (P1_R1171_U84, P1_U3061);
  not ginst3765 (P1_R1171_U85, P1_U3979);
  not ginst3766 (P1_R1171_U86, P1_U3066);
  nand ginst3767 (P1_R1171_U87, P1_U3057, P1_U3976);
  not ginst3768 (P1_R1171_U88, P1_U3054);
  not ginst3769 (P1_R1171_U89, P1_U3974);
  and ginst3770 (P1_R1171_U9, P1_R1171_U262, P1_R1171_U263);
  nand ginst3771 (P1_R1171_U90, P1_R1171_U175, P1_R1171_U305);
  not ginst3772 (P1_R1171_U91, P1_U3076);
  nand ginst3773 (P1_R1171_U92, P1_R1171_U314, P1_R1171_U78);
  nand ginst3774 (P1_R1171_U93, P1_R1171_U259, P1_R1171_U260);
  nand ginst3775 (P1_R1171_U94, P1_R1171_U336, P1_R1171_U69);
  nand ginst3776 (P1_R1171_U95, P1_R1171_U455, P1_R1171_U456);
  nand ginst3777 (P1_R1171_U96, P1_R1171_U502, P1_R1171_U503);
  nand ginst3778 (P1_R1171_U97, P1_R1171_U373, P1_R1171_U374);
  nand ginst3779 (P1_R1171_U98, P1_R1171_U378, P1_R1171_U379);
  nand ginst3780 (P1_R1171_U99, P1_R1171_U385, P1_R1171_U386);
  nand ginst3781 (P1_R1192_U10, P1_R1192_U340, P1_R1192_U343);
  nand ginst3782 (P1_R1192_U100, P1_R1192_U460, P1_R1192_U461);
  nand ginst3783 (P1_R1192_U101, P1_R1192_U465, P1_R1192_U466);
  nand ginst3784 (P1_R1192_U102, P1_R1192_U350, P1_R1192_U351);
  nand ginst3785 (P1_R1192_U103, P1_R1192_U359, P1_R1192_U360);
  nand ginst3786 (P1_R1192_U104, P1_R1192_U366, P1_R1192_U367);
  nand ginst3787 (P1_R1192_U105, P1_R1192_U370, P1_R1192_U371);
  nand ginst3788 (P1_R1192_U106, P1_R1192_U379, P1_R1192_U380);
  nand ginst3789 (P1_R1192_U107, P1_R1192_U398, P1_R1192_U399);
  nand ginst3790 (P1_R1192_U108, P1_R1192_U415, P1_R1192_U416);
  nand ginst3791 (P1_R1192_U109, P1_R1192_U419, P1_R1192_U420);
  nand ginst3792 (P1_R1192_U11, P1_R1192_U329, P1_R1192_U332);
  nand ginst3793 (P1_R1192_U110, P1_R1192_U451, P1_R1192_U452);
  nand ginst3794 (P1_R1192_U111, P1_R1192_U455, P1_R1192_U456);
  nand ginst3795 (P1_R1192_U112, P1_R1192_U472, P1_R1192_U473);
  and ginst3796 (P1_R1192_U113, P1_R1192_U193, P1_R1192_U194);
  and ginst3797 (P1_R1192_U114, P1_R1192_U196, P1_R1192_U201);
  and ginst3798 (P1_R1192_U115, P1_R1192_U180, P1_R1192_U206);
  and ginst3799 (P1_R1192_U116, P1_R1192_U209, P1_R1192_U210);
  and ginst3800 (P1_R1192_U117, P1_R1192_U352, P1_R1192_U353, P1_R1192_U37);
  and ginst3801 (P1_R1192_U118, P1_R1192_U180, P1_R1192_U356);
  and ginst3802 (P1_R1192_U119, P1_R1192_U225, P1_R1192_U6);
  nand ginst3803 (P1_R1192_U12, P1_R1192_U318, P1_R1192_U321);
  and ginst3804 (P1_R1192_U120, P1_R1192_U179, P1_R1192_U363);
  and ginst3805 (P1_R1192_U121, P1_R1192_U27, P1_R1192_U372, P1_R1192_U373);
  and ginst3806 (P1_R1192_U122, P1_R1192_U178, P1_R1192_U376);
  and ginst3807 (P1_R1192_U123, P1_R1192_U174, P1_R1192_U212, P1_R1192_U235);
  and ginst3808 (P1_R1192_U124, P1_R1192_U175, P1_R1192_U252, P1_R1192_U257);
  and ginst3809 (P1_R1192_U125, P1_R1192_U176, P1_R1192_U283);
  and ginst3810 (P1_R1192_U126, P1_R1192_U299, P1_R1192_U300);
  nand ginst3811 (P1_R1192_U127, P1_R1192_U386, P1_R1192_U387);
  and ginst3812 (P1_R1192_U128, P1_R1192_U391, P1_R1192_U392, P1_R1192_U82);
  and ginst3813 (P1_R1192_U129, P1_R1192_U177, P1_R1192_U395);
  nand ginst3814 (P1_R1192_U13, P1_R1192_U310, P1_R1192_U312);
  nand ginst3815 (P1_R1192_U130, P1_R1192_U400, P1_R1192_U401);
  nand ginst3816 (P1_R1192_U131, P1_R1192_U405, P1_R1192_U406);
  and ginst3817 (P1_R1192_U132, P1_R1192_U176, P1_R1192_U412);
  nand ginst3818 (P1_R1192_U133, P1_R1192_U421, P1_R1192_U422);
  nand ginst3819 (P1_R1192_U134, P1_R1192_U426, P1_R1192_U427);
  nand ginst3820 (P1_R1192_U135, P1_R1192_U431, P1_R1192_U432);
  nand ginst3821 (P1_R1192_U136, P1_R1192_U436, P1_R1192_U437);
  nand ginst3822 (P1_R1192_U137, P1_R1192_U441, P1_R1192_U442);
  and ginst3823 (P1_R1192_U138, P1_R1192_U331, P1_R1192_U8);
  and ginst3824 (P1_R1192_U139, P1_R1192_U175, P1_R1192_U448);
  nand ginst3825 (P1_R1192_U14, P1_R1192_U308, P1_R1192_U347);
  nand ginst3826 (P1_R1192_U140, P1_R1192_U457, P1_R1192_U458);
  nand ginst3827 (P1_R1192_U141, P1_R1192_U462, P1_R1192_U463);
  and ginst3828 (P1_R1192_U142, P1_R1192_U342, P1_R1192_U7);
  and ginst3829 (P1_R1192_U143, P1_R1192_U174, P1_R1192_U469);
  and ginst3830 (P1_R1192_U144, P1_R1192_U348, P1_R1192_U349);
  nand ginst3831 (P1_R1192_U145, P1_R1192_U116, P1_R1192_U207);
  and ginst3832 (P1_R1192_U146, P1_R1192_U357, P1_R1192_U358);
  and ginst3833 (P1_R1192_U147, P1_R1192_U364, P1_R1192_U365);
  and ginst3834 (P1_R1192_U148, P1_R1192_U368, P1_R1192_U369);
  nand ginst3835 (P1_R1192_U149, P1_R1192_U113, P1_R1192_U191);
  nand ginst3836 (P1_R1192_U15, P1_R1192_U231, P1_R1192_U233);
  and ginst3837 (P1_R1192_U150, P1_R1192_U377, P1_R1192_U378);
  not ginst3838 (P1_R1192_U151, P1_U3985);
  not ginst3839 (P1_R1192_U152, P1_U3055);
  and ginst3840 (P1_R1192_U153, P1_R1192_U381, P1_R1192_U382);
  and ginst3841 (P1_R1192_U154, P1_R1192_U396, P1_R1192_U397);
  nand ginst3842 (P1_R1192_U155, P1_R1192_U289, P1_R1192_U290);
  nand ginst3843 (P1_R1192_U156, P1_R1192_U285, P1_R1192_U286);
  and ginst3844 (P1_R1192_U157, P1_R1192_U413, P1_R1192_U414);
  and ginst3845 (P1_R1192_U158, P1_R1192_U417, P1_R1192_U418);
  nand ginst3846 (P1_R1192_U159, P1_R1192_U275, P1_R1192_U276);
  nand ginst3847 (P1_R1192_U16, P1_R1192_U223, P1_R1192_U226);
  nand ginst3848 (P1_R1192_U160, P1_R1192_U271, P1_R1192_U272);
  not ginst3849 (P1_R1192_U161, P1_U3455);
  nand ginst3850 (P1_R1192_U162, P1_R1192_U267, P1_R1192_U268);
  not ginst3851 (P1_R1192_U163, P1_U3506);
  nand ginst3852 (P1_R1192_U164, P1_R1192_U259, P1_R1192_U260);
  and ginst3853 (P1_R1192_U165, P1_R1192_U449, P1_R1192_U450);
  and ginst3854 (P1_R1192_U166, P1_R1192_U453, P1_R1192_U454);
  nand ginst3855 (P1_R1192_U167, P1_R1192_U249, P1_R1192_U250);
  nand ginst3856 (P1_R1192_U168, P1_R1192_U245, P1_R1192_U246);
  nand ginst3857 (P1_R1192_U169, P1_R1192_U241, P1_R1192_U242);
  nand ginst3858 (P1_R1192_U17, P1_R1192_U215, P1_R1192_U217);
  and ginst3859 (P1_R1192_U170, P1_R1192_U470, P1_R1192_U471);
  not ginst3860 (P1_R1192_U171, P1_R1192_U82);
  not ginst3861 (P1_R1192_U172, P1_R1192_U27);
  not ginst3862 (P1_R1192_U173, P1_R1192_U37);
  nand ginst3863 (P1_R1192_U174, P1_R1192_U50, P1_U3482);
  nand ginst3864 (P1_R1192_U175, P1_R1192_U59, P1_U3497);
  nand ginst3865 (P1_R1192_U176, P1_R1192_U73, P1_U3980);
  nand ginst3866 (P1_R1192_U177, P1_R1192_U81, P1_U3976);
  nand ginst3867 (P1_R1192_U178, P1_R1192_U26, P1_U3458);
  nand ginst3868 (P1_R1192_U179, P1_R1192_U32, P1_U3467);
  nand ginst3869 (P1_R1192_U18, P1_R1192_U23, P1_R1192_U346);
  nand ginst3870 (P1_R1192_U180, P1_R1192_U36, P1_U3473);
  not ginst3871 (P1_R1192_U181, P1_R1192_U61);
  not ginst3872 (P1_R1192_U182, P1_R1192_U75);
  not ginst3873 (P1_R1192_U183, P1_R1192_U34);
  not ginst3874 (P1_R1192_U184, P1_R1192_U51);
  not ginst3875 (P1_R1192_U185, P1_R1192_U23);
  nand ginst3876 (P1_R1192_U186, P1_R1192_U185, P1_R1192_U24);
  nand ginst3877 (P1_R1192_U187, P1_R1192_U161, P1_R1192_U186);
  nand ginst3878 (P1_R1192_U188, P1_R1192_U23, P1_U3078);
  not ginst3879 (P1_R1192_U189, P1_R1192_U43);
  not ginst3880 (P1_R1192_U19, P1_U3473);
  nand ginst3881 (P1_R1192_U190, P1_R1192_U28, P1_U3461);
  nand ginst3882 (P1_R1192_U191, P1_R1192_U178, P1_R1192_U190, P1_R1192_U43);
  nand ginst3883 (P1_R1192_U192, P1_R1192_U27, P1_R1192_U28);
  nand ginst3884 (P1_R1192_U193, P1_R1192_U192, P1_R1192_U25);
  nand ginst3885 (P1_R1192_U194, P1_R1192_U172, P1_U3064);
  not ginst3886 (P1_R1192_U195, P1_R1192_U149);
  nand ginst3887 (P1_R1192_U196, P1_R1192_U31, P1_U3470);
  nand ginst3888 (P1_R1192_U197, P1_R1192_U29, P1_U3071);
  nand ginst3889 (P1_R1192_U198, P1_R1192_U20, P1_U3067);
  nand ginst3890 (P1_R1192_U199, P1_R1192_U179, P1_R1192_U183);
  not ginst3891 (P1_R1192_U20, P1_U3467);
  nand ginst3892 (P1_R1192_U200, P1_R1192_U199, P1_R1192_U6);
  nand ginst3893 (P1_R1192_U201, P1_R1192_U33, P1_U3464);
  nand ginst3894 (P1_R1192_U202, P1_R1192_U31, P1_U3470);
  nand ginst3895 (P1_R1192_U203, P1_R1192_U114, P1_R1192_U149, P1_R1192_U179);
  nand ginst3896 (P1_R1192_U204, P1_R1192_U200, P1_R1192_U202);
  not ginst3897 (P1_R1192_U205, P1_R1192_U41);
  nand ginst3898 (P1_R1192_U206, P1_R1192_U38, P1_U3476);
  nand ginst3899 (P1_R1192_U207, P1_R1192_U115, P1_R1192_U41);
  nand ginst3900 (P1_R1192_U208, P1_R1192_U37, P1_R1192_U38);
  nand ginst3901 (P1_R1192_U209, P1_R1192_U208, P1_R1192_U35);
  not ginst3902 (P1_R1192_U21, P1_U3458);
  nand ginst3903 (P1_R1192_U210, P1_R1192_U173, P1_U3084);
  not ginst3904 (P1_R1192_U211, P1_R1192_U145);
  nand ginst3905 (P1_R1192_U212, P1_R1192_U40, P1_U3479);
  nand ginst3906 (P1_R1192_U213, P1_R1192_U212, P1_R1192_U51);
  nand ginst3907 (P1_R1192_U214, P1_R1192_U205, P1_R1192_U37);
  nand ginst3908 (P1_R1192_U215, P1_R1192_U118, P1_R1192_U214);
  nand ginst3909 (P1_R1192_U216, P1_R1192_U180, P1_R1192_U41);
  nand ginst3910 (P1_R1192_U217, P1_R1192_U117, P1_R1192_U216);
  nand ginst3911 (P1_R1192_U218, P1_R1192_U180, P1_R1192_U37);
  nand ginst3912 (P1_R1192_U219, P1_R1192_U149, P1_R1192_U201);
  not ginst3913 (P1_R1192_U22, P1_U3450);
  not ginst3914 (P1_R1192_U220, P1_R1192_U42);
  nand ginst3915 (P1_R1192_U221, P1_R1192_U20, P1_U3067);
  nand ginst3916 (P1_R1192_U222, P1_R1192_U220, P1_R1192_U221);
  nand ginst3917 (P1_R1192_U223, P1_R1192_U120, P1_R1192_U222);
  nand ginst3918 (P1_R1192_U224, P1_R1192_U179, P1_R1192_U42);
  nand ginst3919 (P1_R1192_U225, P1_R1192_U31, P1_U3470);
  nand ginst3920 (P1_R1192_U226, P1_R1192_U119, P1_R1192_U224);
  nand ginst3921 (P1_R1192_U227, P1_R1192_U20, P1_U3067);
  nand ginst3922 (P1_R1192_U228, P1_R1192_U179, P1_R1192_U227);
  nand ginst3923 (P1_R1192_U229, P1_R1192_U201, P1_R1192_U34);
  nand ginst3924 (P1_R1192_U23, P1_R1192_U91, P1_U3450);
  nand ginst3925 (P1_R1192_U230, P1_R1192_U189, P1_R1192_U27);
  nand ginst3926 (P1_R1192_U231, P1_R1192_U122, P1_R1192_U230);
  nand ginst3927 (P1_R1192_U232, P1_R1192_U178, P1_R1192_U43);
  nand ginst3928 (P1_R1192_U233, P1_R1192_U121, P1_R1192_U232);
  nand ginst3929 (P1_R1192_U234, P1_R1192_U178, P1_R1192_U27);
  nand ginst3930 (P1_R1192_U235, P1_R1192_U49, P1_U3485);
  nand ginst3931 (P1_R1192_U236, P1_R1192_U48, P1_U3063);
  nand ginst3932 (P1_R1192_U237, P1_R1192_U47, P1_U3062);
  nand ginst3933 (P1_R1192_U238, P1_R1192_U174, P1_R1192_U184);
  nand ginst3934 (P1_R1192_U239, P1_R1192_U238, P1_R1192_U7);
  not ginst3935 (P1_R1192_U24, P1_U3078);
  nand ginst3936 (P1_R1192_U240, P1_R1192_U49, P1_U3485);
  nand ginst3937 (P1_R1192_U241, P1_R1192_U123, P1_R1192_U145);
  nand ginst3938 (P1_R1192_U242, P1_R1192_U239, P1_R1192_U240);
  not ginst3939 (P1_R1192_U243, P1_R1192_U169);
  nand ginst3940 (P1_R1192_U244, P1_R1192_U53, P1_U3488);
  nand ginst3941 (P1_R1192_U245, P1_R1192_U169, P1_R1192_U244);
  nand ginst3942 (P1_R1192_U246, P1_R1192_U52, P1_U3072);
  not ginst3943 (P1_R1192_U247, P1_R1192_U168);
  nand ginst3944 (P1_R1192_U248, P1_R1192_U55, P1_U3491);
  nand ginst3945 (P1_R1192_U249, P1_R1192_U168, P1_R1192_U248);
  not ginst3946 (P1_R1192_U25, P1_U3461);
  nand ginst3947 (P1_R1192_U250, P1_R1192_U54, P1_U3080);
  not ginst3948 (P1_R1192_U251, P1_R1192_U167);
  nand ginst3949 (P1_R1192_U252, P1_R1192_U58, P1_U3500);
  nand ginst3950 (P1_R1192_U253, P1_R1192_U56, P1_U3073);
  nand ginst3951 (P1_R1192_U254, P1_R1192_U46, P1_U3074);
  nand ginst3952 (P1_R1192_U255, P1_R1192_U175, P1_R1192_U181);
  nand ginst3953 (P1_R1192_U256, P1_R1192_U255, P1_R1192_U8);
  nand ginst3954 (P1_R1192_U257, P1_R1192_U60, P1_U3494);
  nand ginst3955 (P1_R1192_U258, P1_R1192_U58, P1_U3500);
  nand ginst3956 (P1_R1192_U259, P1_R1192_U124, P1_R1192_U167);
  not ginst3957 (P1_R1192_U26, P1_U3068);
  nand ginst3958 (P1_R1192_U260, P1_R1192_U256, P1_R1192_U258);
  not ginst3959 (P1_R1192_U261, P1_R1192_U164);
  nand ginst3960 (P1_R1192_U262, P1_R1192_U63, P1_U3503);
  nand ginst3961 (P1_R1192_U263, P1_R1192_U164, P1_R1192_U262);
  nand ginst3962 (P1_R1192_U264, P1_R1192_U62, P1_U3069);
  not ginst3963 (P1_R1192_U265, P1_R1192_U64);
  nand ginst3964 (P1_R1192_U266, P1_R1192_U265, P1_R1192_U65);
  nand ginst3965 (P1_R1192_U267, P1_R1192_U163, P1_R1192_U266);
  nand ginst3966 (P1_R1192_U268, P1_R1192_U64, P1_U3082);
  not ginst3967 (P1_R1192_U269, P1_R1192_U162);
  nand ginst3968 (P1_R1192_U27, P1_R1192_U21, P1_U3068);
  nand ginst3969 (P1_R1192_U270, P1_R1192_U67, P1_U3508);
  nand ginst3970 (P1_R1192_U271, P1_R1192_U162, P1_R1192_U270);
  nand ginst3971 (P1_R1192_U272, P1_R1192_U66, P1_U3081);
  not ginst3972 (P1_R1192_U273, P1_R1192_U160);
  nand ginst3973 (P1_R1192_U274, P1_R1192_U69, P1_U3982);
  nand ginst3974 (P1_R1192_U275, P1_R1192_U160, P1_R1192_U274);
  nand ginst3975 (P1_R1192_U276, P1_R1192_U68, P1_U3076);
  not ginst3976 (P1_R1192_U277, P1_R1192_U159);
  nand ginst3977 (P1_R1192_U278, P1_R1192_U72, P1_U3979);
  nand ginst3978 (P1_R1192_U279, P1_R1192_U70, P1_U3066);
  not ginst3979 (P1_R1192_U28, P1_U3064);
  nand ginst3980 (P1_R1192_U280, P1_R1192_U45, P1_U3061);
  nand ginst3981 (P1_R1192_U281, P1_R1192_U176, P1_R1192_U182);
  nand ginst3982 (P1_R1192_U282, P1_R1192_U281, P1_R1192_U9);
  nand ginst3983 (P1_R1192_U283, P1_R1192_U74, P1_U3981);
  nand ginst3984 (P1_R1192_U284, P1_R1192_U72, P1_U3979);
  nand ginst3985 (P1_R1192_U285, P1_R1192_U125, P1_R1192_U159, P1_R1192_U278);
  nand ginst3986 (P1_R1192_U286, P1_R1192_U282, P1_R1192_U284);
  not ginst3987 (P1_R1192_U287, P1_R1192_U156);
  nand ginst3988 (P1_R1192_U288, P1_R1192_U77, P1_U3978);
  nand ginst3989 (P1_R1192_U289, P1_R1192_U156, P1_R1192_U288);
  not ginst3990 (P1_R1192_U29, P1_U3470);
  nand ginst3991 (P1_R1192_U290, P1_R1192_U76, P1_U3065);
  not ginst3992 (P1_R1192_U291, P1_R1192_U155);
  nand ginst3993 (P1_R1192_U292, P1_R1192_U79, P1_U3977);
  nand ginst3994 (P1_R1192_U293, P1_R1192_U155, P1_R1192_U292);
  nand ginst3995 (P1_R1192_U294, P1_R1192_U78, P1_U3058);
  not ginst3996 (P1_R1192_U295, P1_R1192_U87);
  nand ginst3997 (P1_R1192_U296, P1_R1192_U83, P1_U3975);
  nand ginst3998 (P1_R1192_U297, P1_R1192_U177, P1_R1192_U296, P1_R1192_U87);
  nand ginst3999 (P1_R1192_U298, P1_R1192_U82, P1_R1192_U83);
  nand ginst4000 (P1_R1192_U299, P1_R1192_U298, P1_R1192_U80);
  not ginst4001 (P1_R1192_U30, P1_U3464);
  nand ginst4002 (P1_R1192_U300, P1_R1192_U171, P1_U3053);
  not ginst4003 (P1_R1192_U301, P1_R1192_U86);
  nand ginst4004 (P1_R1192_U302, P1_R1192_U84, P1_U3054);
  nand ginst4005 (P1_R1192_U303, P1_R1192_U301, P1_R1192_U302);
  nand ginst4006 (P1_R1192_U304, P1_R1192_U85, P1_U3974);
  nand ginst4007 (P1_R1192_U305, P1_R1192_U85, P1_U3974);
  nand ginst4008 (P1_R1192_U306, P1_R1192_U305, P1_R1192_U86);
  nand ginst4009 (P1_R1192_U307, P1_R1192_U84, P1_U3054);
  nand ginst4010 (P1_R1192_U308, P1_R1192_U153, P1_R1192_U306, P1_R1192_U307);
  nand ginst4011 (P1_R1192_U309, P1_R1192_U295, P1_R1192_U82);
  not ginst4012 (P1_R1192_U31, P1_U3071);
  nand ginst4013 (P1_R1192_U310, P1_R1192_U129, P1_R1192_U309);
  nand ginst4014 (P1_R1192_U311, P1_R1192_U177, P1_R1192_U87);
  nand ginst4015 (P1_R1192_U312, P1_R1192_U128, P1_R1192_U311);
  nand ginst4016 (P1_R1192_U313, P1_R1192_U177, P1_R1192_U82);
  nand ginst4017 (P1_R1192_U314, P1_R1192_U159, P1_R1192_U283);
  not ginst4018 (P1_R1192_U315, P1_R1192_U88);
  nand ginst4019 (P1_R1192_U316, P1_R1192_U45, P1_U3061);
  nand ginst4020 (P1_R1192_U317, P1_R1192_U315, P1_R1192_U316);
  nand ginst4021 (P1_R1192_U318, P1_R1192_U132, P1_R1192_U317);
  nand ginst4022 (P1_R1192_U319, P1_R1192_U176, P1_R1192_U88);
  not ginst4023 (P1_R1192_U32, P1_U3067);
  nand ginst4024 (P1_R1192_U320, P1_R1192_U72, P1_U3979);
  nand ginst4025 (P1_R1192_U321, P1_R1192_U319, P1_R1192_U320, P1_R1192_U9);
  nand ginst4026 (P1_R1192_U322, P1_R1192_U45, P1_U3061);
  nand ginst4027 (P1_R1192_U323, P1_R1192_U176, P1_R1192_U322);
  nand ginst4028 (P1_R1192_U324, P1_R1192_U283, P1_R1192_U75);
  nand ginst4029 (P1_R1192_U325, P1_R1192_U167, P1_R1192_U257);
  not ginst4030 (P1_R1192_U326, P1_R1192_U89);
  nand ginst4031 (P1_R1192_U327, P1_R1192_U46, P1_U3074);
  nand ginst4032 (P1_R1192_U328, P1_R1192_U326, P1_R1192_U327);
  nand ginst4033 (P1_R1192_U329, P1_R1192_U139, P1_R1192_U328);
  not ginst4034 (P1_R1192_U33, P1_U3060);
  nand ginst4035 (P1_R1192_U330, P1_R1192_U175, P1_R1192_U89);
  nand ginst4036 (P1_R1192_U331, P1_R1192_U58, P1_U3500);
  nand ginst4037 (P1_R1192_U332, P1_R1192_U138, P1_R1192_U330);
  nand ginst4038 (P1_R1192_U333, P1_R1192_U46, P1_U3074);
  nand ginst4039 (P1_R1192_U334, P1_R1192_U175, P1_R1192_U333);
  nand ginst4040 (P1_R1192_U335, P1_R1192_U257, P1_R1192_U61);
  nand ginst4041 (P1_R1192_U336, P1_R1192_U145, P1_R1192_U212);
  not ginst4042 (P1_R1192_U337, P1_R1192_U90);
  nand ginst4043 (P1_R1192_U338, P1_R1192_U47, P1_U3062);
  nand ginst4044 (P1_R1192_U339, P1_R1192_U337, P1_R1192_U338);
  nand ginst4045 (P1_R1192_U34, P1_R1192_U30, P1_U3060);
  nand ginst4046 (P1_R1192_U340, P1_R1192_U143, P1_R1192_U339);
  nand ginst4047 (P1_R1192_U341, P1_R1192_U174, P1_R1192_U90);
  nand ginst4048 (P1_R1192_U342, P1_R1192_U49, P1_U3485);
  nand ginst4049 (P1_R1192_U343, P1_R1192_U142, P1_R1192_U341);
  nand ginst4050 (P1_R1192_U344, P1_R1192_U47, P1_U3062);
  nand ginst4051 (P1_R1192_U345, P1_R1192_U174, P1_R1192_U344);
  nand ginst4052 (P1_R1192_U346, P1_R1192_U22, P1_U3077);
  nand ginst4053 (P1_R1192_U347, P1_R1192_U303, P1_R1192_U304, P1_R1192_U385);
  nand ginst4054 (P1_R1192_U348, P1_R1192_U40, P1_U3479);
  nand ginst4055 (P1_R1192_U349, P1_R1192_U39, P1_U3083);
  not ginst4056 (P1_R1192_U35, P1_U3476);
  nand ginst4057 (P1_R1192_U350, P1_R1192_U145, P1_R1192_U213);
  nand ginst4058 (P1_R1192_U351, P1_R1192_U144, P1_R1192_U211);
  nand ginst4059 (P1_R1192_U352, P1_R1192_U38, P1_U3476);
  nand ginst4060 (P1_R1192_U353, P1_R1192_U35, P1_U3084);
  nand ginst4061 (P1_R1192_U354, P1_R1192_U38, P1_U3476);
  nand ginst4062 (P1_R1192_U355, P1_R1192_U35, P1_U3084);
  nand ginst4063 (P1_R1192_U356, P1_R1192_U354, P1_R1192_U355);
  nand ginst4064 (P1_R1192_U357, P1_R1192_U36, P1_U3473);
  nand ginst4065 (P1_R1192_U358, P1_R1192_U19, P1_U3070);
  nand ginst4066 (P1_R1192_U359, P1_R1192_U218, P1_R1192_U41);
  not ginst4067 (P1_R1192_U36, P1_U3070);
  nand ginst4068 (P1_R1192_U360, P1_R1192_U146, P1_R1192_U205);
  nand ginst4069 (P1_R1192_U361, P1_R1192_U31, P1_U3470);
  nand ginst4070 (P1_R1192_U362, P1_R1192_U29, P1_U3071);
  nand ginst4071 (P1_R1192_U363, P1_R1192_U361, P1_R1192_U362);
  nand ginst4072 (P1_R1192_U364, P1_R1192_U32, P1_U3467);
  nand ginst4073 (P1_R1192_U365, P1_R1192_U20, P1_U3067);
  nand ginst4074 (P1_R1192_U366, P1_R1192_U228, P1_R1192_U42);
  nand ginst4075 (P1_R1192_U367, P1_R1192_U147, P1_R1192_U220);
  nand ginst4076 (P1_R1192_U368, P1_R1192_U33, P1_U3464);
  nand ginst4077 (P1_R1192_U369, P1_R1192_U30, P1_U3060);
  nand ginst4078 (P1_R1192_U37, P1_R1192_U19, P1_U3070);
  nand ginst4079 (P1_R1192_U370, P1_R1192_U149, P1_R1192_U229);
  nand ginst4080 (P1_R1192_U371, P1_R1192_U148, P1_R1192_U195);
  nand ginst4081 (P1_R1192_U372, P1_R1192_U28, P1_U3461);
  nand ginst4082 (P1_R1192_U373, P1_R1192_U25, P1_U3064);
  nand ginst4083 (P1_R1192_U374, P1_R1192_U28, P1_U3461);
  nand ginst4084 (P1_R1192_U375, P1_R1192_U25, P1_U3064);
  nand ginst4085 (P1_R1192_U376, P1_R1192_U374, P1_R1192_U375);
  nand ginst4086 (P1_R1192_U377, P1_R1192_U26, P1_U3458);
  nand ginst4087 (P1_R1192_U378, P1_R1192_U21, P1_U3068);
  nand ginst4088 (P1_R1192_U379, P1_R1192_U234, P1_R1192_U43);
  not ginst4089 (P1_R1192_U38, P1_U3084);
  nand ginst4090 (P1_R1192_U380, P1_R1192_U150, P1_R1192_U189);
  nand ginst4091 (P1_R1192_U381, P1_R1192_U152, P1_U3985);
  nand ginst4092 (P1_R1192_U382, P1_R1192_U151, P1_U3055);
  nand ginst4093 (P1_R1192_U383, P1_R1192_U152, P1_U3985);
  nand ginst4094 (P1_R1192_U384, P1_R1192_U151, P1_U3055);
  nand ginst4095 (P1_R1192_U385, P1_R1192_U383, P1_R1192_U384);
  nand ginst4096 (P1_R1192_U386, P1_R1192_U85, P1_U3974);
  nand ginst4097 (P1_R1192_U387, P1_R1192_U84, P1_U3054);
  not ginst4098 (P1_R1192_U388, P1_R1192_U127);
  nand ginst4099 (P1_R1192_U389, P1_R1192_U301, P1_R1192_U388);
  not ginst4100 (P1_R1192_U39, P1_U3479);
  nand ginst4101 (P1_R1192_U390, P1_R1192_U127, P1_R1192_U86);
  nand ginst4102 (P1_R1192_U391, P1_R1192_U83, P1_U3975);
  nand ginst4103 (P1_R1192_U392, P1_R1192_U80, P1_U3053);
  nand ginst4104 (P1_R1192_U393, P1_R1192_U83, P1_U3975);
  nand ginst4105 (P1_R1192_U394, P1_R1192_U80, P1_U3053);
  nand ginst4106 (P1_R1192_U395, P1_R1192_U393, P1_R1192_U394);
  nand ginst4107 (P1_R1192_U396, P1_R1192_U81, P1_U3976);
  nand ginst4108 (P1_R1192_U397, P1_R1192_U44, P1_U3057);
  nand ginst4109 (P1_R1192_U398, P1_R1192_U313, P1_R1192_U87);
  nand ginst4110 (P1_R1192_U399, P1_R1192_U154, P1_R1192_U295);
  not ginst4111 (P1_R1192_U40, P1_U3083);
  nand ginst4112 (P1_R1192_U400, P1_R1192_U79, P1_U3977);
  nand ginst4113 (P1_R1192_U401, P1_R1192_U78, P1_U3058);
  not ginst4114 (P1_R1192_U402, P1_R1192_U130);
  nand ginst4115 (P1_R1192_U403, P1_R1192_U291, P1_R1192_U402);
  nand ginst4116 (P1_R1192_U404, P1_R1192_U130, P1_R1192_U155);
  nand ginst4117 (P1_R1192_U405, P1_R1192_U77, P1_U3978);
  nand ginst4118 (P1_R1192_U406, P1_R1192_U76, P1_U3065);
  not ginst4119 (P1_R1192_U407, P1_R1192_U131);
  nand ginst4120 (P1_R1192_U408, P1_R1192_U287, P1_R1192_U407);
  nand ginst4121 (P1_R1192_U409, P1_R1192_U131, P1_R1192_U156);
  nand ginst4122 (P1_R1192_U41, P1_R1192_U203, P1_R1192_U204);
  nand ginst4123 (P1_R1192_U410, P1_R1192_U72, P1_U3979);
  nand ginst4124 (P1_R1192_U411, P1_R1192_U70, P1_U3066);
  nand ginst4125 (P1_R1192_U412, P1_R1192_U410, P1_R1192_U411);
  nand ginst4126 (P1_R1192_U413, P1_R1192_U73, P1_U3980);
  nand ginst4127 (P1_R1192_U414, P1_R1192_U45, P1_U3061);
  nand ginst4128 (P1_R1192_U415, P1_R1192_U323, P1_R1192_U88);
  nand ginst4129 (P1_R1192_U416, P1_R1192_U157, P1_R1192_U315);
  nand ginst4130 (P1_R1192_U417, P1_R1192_U74, P1_U3981);
  nand ginst4131 (P1_R1192_U418, P1_R1192_U71, P1_U3075);
  nand ginst4132 (P1_R1192_U419, P1_R1192_U159, P1_R1192_U324);
  nand ginst4133 (P1_R1192_U42, P1_R1192_U219, P1_R1192_U34);
  nand ginst4134 (P1_R1192_U420, P1_R1192_U158, P1_R1192_U277);
  nand ginst4135 (P1_R1192_U421, P1_R1192_U69, P1_U3982);
  nand ginst4136 (P1_R1192_U422, P1_R1192_U68, P1_U3076);
  not ginst4137 (P1_R1192_U423, P1_R1192_U133);
  nand ginst4138 (P1_R1192_U424, P1_R1192_U273, P1_R1192_U423);
  nand ginst4139 (P1_R1192_U425, P1_R1192_U133, P1_R1192_U160);
  nand ginst4140 (P1_R1192_U426, P1_R1192_U185, P1_R1192_U24);
  nand ginst4141 (P1_R1192_U427, P1_R1192_U23, P1_U3078);
  not ginst4142 (P1_R1192_U428, P1_R1192_U134);
  nand ginst4143 (P1_R1192_U429, P1_R1192_U428, P1_U3455);
  nand ginst4144 (P1_R1192_U43, P1_R1192_U187, P1_R1192_U188);
  nand ginst4145 (P1_R1192_U430, P1_R1192_U134, P1_R1192_U161);
  nand ginst4146 (P1_R1192_U431, P1_R1192_U67, P1_U3508);
  nand ginst4147 (P1_R1192_U432, P1_R1192_U66, P1_U3081);
  not ginst4148 (P1_R1192_U433, P1_R1192_U135);
  nand ginst4149 (P1_R1192_U434, P1_R1192_U269, P1_R1192_U433);
  nand ginst4150 (P1_R1192_U435, P1_R1192_U135, P1_R1192_U162);
  nand ginst4151 (P1_R1192_U436, P1_R1192_U65, P1_U3506);
  nand ginst4152 (P1_R1192_U437, P1_R1192_U163, P1_U3082);
  not ginst4153 (P1_R1192_U438, P1_R1192_U136);
  nand ginst4154 (P1_R1192_U439, P1_R1192_U265, P1_R1192_U438);
  not ginst4155 (P1_R1192_U44, P1_U3976);
  nand ginst4156 (P1_R1192_U440, P1_R1192_U136, P1_R1192_U64);
  nand ginst4157 (P1_R1192_U441, P1_R1192_U63, P1_U3503);
  nand ginst4158 (P1_R1192_U442, P1_R1192_U62, P1_U3069);
  not ginst4159 (P1_R1192_U443, P1_R1192_U137);
  nand ginst4160 (P1_R1192_U444, P1_R1192_U261, P1_R1192_U443);
  nand ginst4161 (P1_R1192_U445, P1_R1192_U137, P1_R1192_U164);
  nand ginst4162 (P1_R1192_U446, P1_R1192_U58, P1_U3500);
  nand ginst4163 (P1_R1192_U447, P1_R1192_U56, P1_U3073);
  nand ginst4164 (P1_R1192_U448, P1_R1192_U446, P1_R1192_U447);
  nand ginst4165 (P1_R1192_U449, P1_R1192_U59, P1_U3497);
  not ginst4166 (P1_R1192_U45, P1_U3980);
  nand ginst4167 (P1_R1192_U450, P1_R1192_U46, P1_U3074);
  nand ginst4168 (P1_R1192_U451, P1_R1192_U334, P1_R1192_U89);
  nand ginst4169 (P1_R1192_U452, P1_R1192_U165, P1_R1192_U326);
  nand ginst4170 (P1_R1192_U453, P1_R1192_U60, P1_U3494);
  nand ginst4171 (P1_R1192_U454, P1_R1192_U57, P1_U3079);
  nand ginst4172 (P1_R1192_U455, P1_R1192_U167, P1_R1192_U335);
  nand ginst4173 (P1_R1192_U456, P1_R1192_U166, P1_R1192_U251);
  nand ginst4174 (P1_R1192_U457, P1_R1192_U55, P1_U3491);
  nand ginst4175 (P1_R1192_U458, P1_R1192_U54, P1_U3080);
  not ginst4176 (P1_R1192_U459, P1_R1192_U140);
  not ginst4177 (P1_R1192_U46, P1_U3497);
  nand ginst4178 (P1_R1192_U460, P1_R1192_U247, P1_R1192_U459);
  nand ginst4179 (P1_R1192_U461, P1_R1192_U140, P1_R1192_U168);
  nand ginst4180 (P1_R1192_U462, P1_R1192_U53, P1_U3488);
  nand ginst4181 (P1_R1192_U463, P1_R1192_U52, P1_U3072);
  not ginst4182 (P1_R1192_U464, P1_R1192_U141);
  nand ginst4183 (P1_R1192_U465, P1_R1192_U243, P1_R1192_U464);
  nand ginst4184 (P1_R1192_U466, P1_R1192_U141, P1_R1192_U169);
  nand ginst4185 (P1_R1192_U467, P1_R1192_U49, P1_U3485);
  nand ginst4186 (P1_R1192_U468, P1_R1192_U48, P1_U3063);
  nand ginst4187 (P1_R1192_U469, P1_R1192_U467, P1_R1192_U468);
  not ginst4188 (P1_R1192_U47, P1_U3482);
  nand ginst4189 (P1_R1192_U470, P1_R1192_U50, P1_U3482);
  nand ginst4190 (P1_R1192_U471, P1_R1192_U47, P1_U3062);
  nand ginst4191 (P1_R1192_U472, P1_R1192_U345, P1_R1192_U90);
  nand ginst4192 (P1_R1192_U473, P1_R1192_U170, P1_R1192_U337);
  not ginst4193 (P1_R1192_U48, P1_U3485);
  not ginst4194 (P1_R1192_U49, P1_U3063);
  not ginst4195 (P1_R1192_U50, P1_U3062);
  nand ginst4196 (P1_R1192_U51, P1_R1192_U39, P1_U3083);
  not ginst4197 (P1_R1192_U52, P1_U3488);
  not ginst4198 (P1_R1192_U53, P1_U3072);
  not ginst4199 (P1_R1192_U54, P1_U3491);
  not ginst4200 (P1_R1192_U55, P1_U3080);
  not ginst4201 (P1_R1192_U56, P1_U3500);
  not ginst4202 (P1_R1192_U57, P1_U3494);
  not ginst4203 (P1_R1192_U58, P1_U3073);
  not ginst4204 (P1_R1192_U59, P1_U3074);
  and ginst4205 (P1_R1192_U6, P1_R1192_U197, P1_R1192_U198);
  not ginst4206 (P1_R1192_U60, P1_U3079);
  nand ginst4207 (P1_R1192_U61, P1_R1192_U57, P1_U3079);
  not ginst4208 (P1_R1192_U62, P1_U3503);
  not ginst4209 (P1_R1192_U63, P1_U3069);
  nand ginst4210 (P1_R1192_U64, P1_R1192_U263, P1_R1192_U264);
  not ginst4211 (P1_R1192_U65, P1_U3082);
  not ginst4212 (P1_R1192_U66, P1_U3508);
  not ginst4213 (P1_R1192_U67, P1_U3081);
  not ginst4214 (P1_R1192_U68, P1_U3982);
  not ginst4215 (P1_R1192_U69, P1_U3076);
  and ginst4216 (P1_R1192_U7, P1_R1192_U236, P1_R1192_U237);
  not ginst4217 (P1_R1192_U70, P1_U3979);
  not ginst4218 (P1_R1192_U71, P1_U3981);
  not ginst4219 (P1_R1192_U72, P1_U3066);
  not ginst4220 (P1_R1192_U73, P1_U3061);
  not ginst4221 (P1_R1192_U74, P1_U3075);
  nand ginst4222 (P1_R1192_U75, P1_R1192_U71, P1_U3075);
  not ginst4223 (P1_R1192_U76, P1_U3978);
  not ginst4224 (P1_R1192_U77, P1_U3065);
  not ginst4225 (P1_R1192_U78, P1_U3977);
  not ginst4226 (P1_R1192_U79, P1_U3058);
  and ginst4227 (P1_R1192_U8, P1_R1192_U253, P1_R1192_U254);
  not ginst4228 (P1_R1192_U80, P1_U3975);
  not ginst4229 (P1_R1192_U81, P1_U3057);
  nand ginst4230 (P1_R1192_U82, P1_R1192_U44, P1_U3057);
  not ginst4231 (P1_R1192_U83, P1_U3053);
  not ginst4232 (P1_R1192_U84, P1_U3974);
  not ginst4233 (P1_R1192_U85, P1_U3054);
  nand ginst4234 (P1_R1192_U86, P1_R1192_U126, P1_R1192_U297);
  nand ginst4235 (P1_R1192_U87, P1_R1192_U293, P1_R1192_U294);
  nand ginst4236 (P1_R1192_U88, P1_R1192_U314, P1_R1192_U75);
  nand ginst4237 (P1_R1192_U89, P1_R1192_U325, P1_R1192_U61);
  and ginst4238 (P1_R1192_U9, P1_R1192_U279, P1_R1192_U280);
  nand ginst4239 (P1_R1192_U90, P1_R1192_U336, P1_R1192_U51);
  not ginst4240 (P1_R1192_U91, P1_U3077);
  nand ginst4241 (P1_R1192_U92, P1_R1192_U389, P1_R1192_U390);
  nand ginst4242 (P1_R1192_U93, P1_R1192_U403, P1_R1192_U404);
  nand ginst4243 (P1_R1192_U94, P1_R1192_U408, P1_R1192_U409);
  nand ginst4244 (P1_R1192_U95, P1_R1192_U424, P1_R1192_U425);
  nand ginst4245 (P1_R1192_U96, P1_R1192_U429, P1_R1192_U430);
  nand ginst4246 (P1_R1192_U97, P1_R1192_U434, P1_R1192_U435);
  nand ginst4247 (P1_R1192_U98, P1_R1192_U439, P1_R1192_U440);
  nand ginst4248 (P1_R1192_U99, P1_R1192_U444, P1_R1192_U445);
  nand ginst4249 (P1_R1207_U10, P1_R1207_U340, P1_R1207_U343);
  nand ginst4250 (P1_R1207_U100, P1_R1207_U460, P1_R1207_U461);
  nand ginst4251 (P1_R1207_U101, P1_R1207_U465, P1_R1207_U466);
  nand ginst4252 (P1_R1207_U102, P1_R1207_U350, P1_R1207_U351);
  nand ginst4253 (P1_R1207_U103, P1_R1207_U359, P1_R1207_U360);
  nand ginst4254 (P1_R1207_U104, P1_R1207_U366, P1_R1207_U367);
  nand ginst4255 (P1_R1207_U105, P1_R1207_U370, P1_R1207_U371);
  nand ginst4256 (P1_R1207_U106, P1_R1207_U379, P1_R1207_U380);
  nand ginst4257 (P1_R1207_U107, P1_R1207_U398, P1_R1207_U399);
  nand ginst4258 (P1_R1207_U108, P1_R1207_U415, P1_R1207_U416);
  nand ginst4259 (P1_R1207_U109, P1_R1207_U419, P1_R1207_U420);
  nand ginst4260 (P1_R1207_U11, P1_R1207_U329, P1_R1207_U332);
  nand ginst4261 (P1_R1207_U110, P1_R1207_U451, P1_R1207_U452);
  nand ginst4262 (P1_R1207_U111, P1_R1207_U455, P1_R1207_U456);
  nand ginst4263 (P1_R1207_U112, P1_R1207_U472, P1_R1207_U473);
  and ginst4264 (P1_R1207_U113, P1_R1207_U193, P1_R1207_U194);
  and ginst4265 (P1_R1207_U114, P1_R1207_U196, P1_R1207_U201);
  and ginst4266 (P1_R1207_U115, P1_R1207_U180, P1_R1207_U206);
  and ginst4267 (P1_R1207_U116, P1_R1207_U209, P1_R1207_U210);
  and ginst4268 (P1_R1207_U117, P1_R1207_U352, P1_R1207_U353, P1_R1207_U37);
  and ginst4269 (P1_R1207_U118, P1_R1207_U180, P1_R1207_U356);
  and ginst4270 (P1_R1207_U119, P1_R1207_U225, P1_R1207_U6);
  nand ginst4271 (P1_R1207_U12, P1_R1207_U318, P1_R1207_U321);
  and ginst4272 (P1_R1207_U120, P1_R1207_U179, P1_R1207_U363);
  and ginst4273 (P1_R1207_U121, P1_R1207_U27, P1_R1207_U372, P1_R1207_U373);
  and ginst4274 (P1_R1207_U122, P1_R1207_U178, P1_R1207_U376);
  and ginst4275 (P1_R1207_U123, P1_R1207_U174, P1_R1207_U212, P1_R1207_U235);
  and ginst4276 (P1_R1207_U124, P1_R1207_U175, P1_R1207_U252, P1_R1207_U257);
  and ginst4277 (P1_R1207_U125, P1_R1207_U176, P1_R1207_U283);
  and ginst4278 (P1_R1207_U126, P1_R1207_U299, P1_R1207_U300);
  nand ginst4279 (P1_R1207_U127, P1_R1207_U386, P1_R1207_U387);
  and ginst4280 (P1_R1207_U128, P1_R1207_U391, P1_R1207_U392, P1_R1207_U82);
  and ginst4281 (P1_R1207_U129, P1_R1207_U177, P1_R1207_U395);
  nand ginst4282 (P1_R1207_U13, P1_R1207_U310, P1_R1207_U312);
  nand ginst4283 (P1_R1207_U130, P1_R1207_U400, P1_R1207_U401);
  nand ginst4284 (P1_R1207_U131, P1_R1207_U405, P1_R1207_U406);
  and ginst4285 (P1_R1207_U132, P1_R1207_U176, P1_R1207_U412);
  nand ginst4286 (P1_R1207_U133, P1_R1207_U421, P1_R1207_U422);
  nand ginst4287 (P1_R1207_U134, P1_R1207_U426, P1_R1207_U427);
  nand ginst4288 (P1_R1207_U135, P1_R1207_U431, P1_R1207_U432);
  nand ginst4289 (P1_R1207_U136, P1_R1207_U436, P1_R1207_U437);
  nand ginst4290 (P1_R1207_U137, P1_R1207_U441, P1_R1207_U442);
  and ginst4291 (P1_R1207_U138, P1_R1207_U331, P1_R1207_U8);
  and ginst4292 (P1_R1207_U139, P1_R1207_U175, P1_R1207_U448);
  nand ginst4293 (P1_R1207_U14, P1_R1207_U308, P1_R1207_U347);
  nand ginst4294 (P1_R1207_U140, P1_R1207_U457, P1_R1207_U458);
  nand ginst4295 (P1_R1207_U141, P1_R1207_U462, P1_R1207_U463);
  and ginst4296 (P1_R1207_U142, P1_R1207_U342, P1_R1207_U7);
  and ginst4297 (P1_R1207_U143, P1_R1207_U174, P1_R1207_U469);
  and ginst4298 (P1_R1207_U144, P1_R1207_U348, P1_R1207_U349);
  nand ginst4299 (P1_R1207_U145, P1_R1207_U116, P1_R1207_U207);
  and ginst4300 (P1_R1207_U146, P1_R1207_U357, P1_R1207_U358);
  and ginst4301 (P1_R1207_U147, P1_R1207_U364, P1_R1207_U365);
  and ginst4302 (P1_R1207_U148, P1_R1207_U368, P1_R1207_U369);
  nand ginst4303 (P1_R1207_U149, P1_R1207_U113, P1_R1207_U191);
  nand ginst4304 (P1_R1207_U15, P1_R1207_U231, P1_R1207_U233);
  and ginst4305 (P1_R1207_U150, P1_R1207_U377, P1_R1207_U378);
  not ginst4306 (P1_R1207_U151, P1_U3985);
  not ginst4307 (P1_R1207_U152, P1_U3055);
  and ginst4308 (P1_R1207_U153, P1_R1207_U381, P1_R1207_U382);
  and ginst4309 (P1_R1207_U154, P1_R1207_U396, P1_R1207_U397);
  nand ginst4310 (P1_R1207_U155, P1_R1207_U289, P1_R1207_U290);
  nand ginst4311 (P1_R1207_U156, P1_R1207_U285, P1_R1207_U286);
  and ginst4312 (P1_R1207_U157, P1_R1207_U413, P1_R1207_U414);
  and ginst4313 (P1_R1207_U158, P1_R1207_U417, P1_R1207_U418);
  nand ginst4314 (P1_R1207_U159, P1_R1207_U275, P1_R1207_U276);
  nand ginst4315 (P1_R1207_U16, P1_R1207_U223, P1_R1207_U226);
  nand ginst4316 (P1_R1207_U160, P1_R1207_U271, P1_R1207_U272);
  not ginst4317 (P1_R1207_U161, P1_U3455);
  nand ginst4318 (P1_R1207_U162, P1_R1207_U267, P1_R1207_U268);
  not ginst4319 (P1_R1207_U163, P1_U3506);
  nand ginst4320 (P1_R1207_U164, P1_R1207_U259, P1_R1207_U260);
  and ginst4321 (P1_R1207_U165, P1_R1207_U449, P1_R1207_U450);
  and ginst4322 (P1_R1207_U166, P1_R1207_U453, P1_R1207_U454);
  nand ginst4323 (P1_R1207_U167, P1_R1207_U249, P1_R1207_U250);
  nand ginst4324 (P1_R1207_U168, P1_R1207_U245, P1_R1207_U246);
  nand ginst4325 (P1_R1207_U169, P1_R1207_U241, P1_R1207_U242);
  nand ginst4326 (P1_R1207_U17, P1_R1207_U215, P1_R1207_U217);
  and ginst4327 (P1_R1207_U170, P1_R1207_U470, P1_R1207_U471);
  not ginst4328 (P1_R1207_U171, P1_R1207_U82);
  not ginst4329 (P1_R1207_U172, P1_R1207_U27);
  not ginst4330 (P1_R1207_U173, P1_R1207_U37);
  nand ginst4331 (P1_R1207_U174, P1_R1207_U50, P1_U3482);
  nand ginst4332 (P1_R1207_U175, P1_R1207_U59, P1_U3497);
  nand ginst4333 (P1_R1207_U176, P1_R1207_U73, P1_U3980);
  nand ginst4334 (P1_R1207_U177, P1_R1207_U81, P1_U3976);
  nand ginst4335 (P1_R1207_U178, P1_R1207_U26, P1_U3458);
  nand ginst4336 (P1_R1207_U179, P1_R1207_U32, P1_U3467);
  nand ginst4337 (P1_R1207_U18, P1_R1207_U23, P1_R1207_U346);
  nand ginst4338 (P1_R1207_U180, P1_R1207_U36, P1_U3473);
  not ginst4339 (P1_R1207_U181, P1_R1207_U61);
  not ginst4340 (P1_R1207_U182, P1_R1207_U75);
  not ginst4341 (P1_R1207_U183, P1_R1207_U34);
  not ginst4342 (P1_R1207_U184, P1_R1207_U51);
  not ginst4343 (P1_R1207_U185, P1_R1207_U23);
  nand ginst4344 (P1_R1207_U186, P1_R1207_U185, P1_R1207_U24);
  nand ginst4345 (P1_R1207_U187, P1_R1207_U161, P1_R1207_U186);
  nand ginst4346 (P1_R1207_U188, P1_R1207_U23, P1_U3078);
  not ginst4347 (P1_R1207_U189, P1_R1207_U43);
  not ginst4348 (P1_R1207_U19, P1_U3473);
  nand ginst4349 (P1_R1207_U190, P1_R1207_U28, P1_U3461);
  nand ginst4350 (P1_R1207_U191, P1_R1207_U178, P1_R1207_U190, P1_R1207_U43);
  nand ginst4351 (P1_R1207_U192, P1_R1207_U27, P1_R1207_U28);
  nand ginst4352 (P1_R1207_U193, P1_R1207_U192, P1_R1207_U25);
  nand ginst4353 (P1_R1207_U194, P1_R1207_U172, P1_U3064);
  not ginst4354 (P1_R1207_U195, P1_R1207_U149);
  nand ginst4355 (P1_R1207_U196, P1_R1207_U31, P1_U3470);
  nand ginst4356 (P1_R1207_U197, P1_R1207_U29, P1_U3071);
  nand ginst4357 (P1_R1207_U198, P1_R1207_U20, P1_U3067);
  nand ginst4358 (P1_R1207_U199, P1_R1207_U179, P1_R1207_U183);
  not ginst4359 (P1_R1207_U20, P1_U3467);
  nand ginst4360 (P1_R1207_U200, P1_R1207_U199, P1_R1207_U6);
  nand ginst4361 (P1_R1207_U201, P1_R1207_U33, P1_U3464);
  nand ginst4362 (P1_R1207_U202, P1_R1207_U31, P1_U3470);
  nand ginst4363 (P1_R1207_U203, P1_R1207_U114, P1_R1207_U149, P1_R1207_U179);
  nand ginst4364 (P1_R1207_U204, P1_R1207_U200, P1_R1207_U202);
  not ginst4365 (P1_R1207_U205, P1_R1207_U41);
  nand ginst4366 (P1_R1207_U206, P1_R1207_U38, P1_U3476);
  nand ginst4367 (P1_R1207_U207, P1_R1207_U115, P1_R1207_U41);
  nand ginst4368 (P1_R1207_U208, P1_R1207_U37, P1_R1207_U38);
  nand ginst4369 (P1_R1207_U209, P1_R1207_U208, P1_R1207_U35);
  not ginst4370 (P1_R1207_U21, P1_U3458);
  nand ginst4371 (P1_R1207_U210, P1_R1207_U173, P1_U3084);
  not ginst4372 (P1_R1207_U211, P1_R1207_U145);
  nand ginst4373 (P1_R1207_U212, P1_R1207_U40, P1_U3479);
  nand ginst4374 (P1_R1207_U213, P1_R1207_U212, P1_R1207_U51);
  nand ginst4375 (P1_R1207_U214, P1_R1207_U205, P1_R1207_U37);
  nand ginst4376 (P1_R1207_U215, P1_R1207_U118, P1_R1207_U214);
  nand ginst4377 (P1_R1207_U216, P1_R1207_U180, P1_R1207_U41);
  nand ginst4378 (P1_R1207_U217, P1_R1207_U117, P1_R1207_U216);
  nand ginst4379 (P1_R1207_U218, P1_R1207_U180, P1_R1207_U37);
  nand ginst4380 (P1_R1207_U219, P1_R1207_U149, P1_R1207_U201);
  not ginst4381 (P1_R1207_U22, P1_U3450);
  not ginst4382 (P1_R1207_U220, P1_R1207_U42);
  nand ginst4383 (P1_R1207_U221, P1_R1207_U20, P1_U3067);
  nand ginst4384 (P1_R1207_U222, P1_R1207_U220, P1_R1207_U221);
  nand ginst4385 (P1_R1207_U223, P1_R1207_U120, P1_R1207_U222);
  nand ginst4386 (P1_R1207_U224, P1_R1207_U179, P1_R1207_U42);
  nand ginst4387 (P1_R1207_U225, P1_R1207_U31, P1_U3470);
  nand ginst4388 (P1_R1207_U226, P1_R1207_U119, P1_R1207_U224);
  nand ginst4389 (P1_R1207_U227, P1_R1207_U20, P1_U3067);
  nand ginst4390 (P1_R1207_U228, P1_R1207_U179, P1_R1207_U227);
  nand ginst4391 (P1_R1207_U229, P1_R1207_U201, P1_R1207_U34);
  nand ginst4392 (P1_R1207_U23, P1_R1207_U91, P1_U3450);
  nand ginst4393 (P1_R1207_U230, P1_R1207_U189, P1_R1207_U27);
  nand ginst4394 (P1_R1207_U231, P1_R1207_U122, P1_R1207_U230);
  nand ginst4395 (P1_R1207_U232, P1_R1207_U178, P1_R1207_U43);
  nand ginst4396 (P1_R1207_U233, P1_R1207_U121, P1_R1207_U232);
  nand ginst4397 (P1_R1207_U234, P1_R1207_U178, P1_R1207_U27);
  nand ginst4398 (P1_R1207_U235, P1_R1207_U49, P1_U3485);
  nand ginst4399 (P1_R1207_U236, P1_R1207_U48, P1_U3063);
  nand ginst4400 (P1_R1207_U237, P1_R1207_U47, P1_U3062);
  nand ginst4401 (P1_R1207_U238, P1_R1207_U174, P1_R1207_U184);
  nand ginst4402 (P1_R1207_U239, P1_R1207_U238, P1_R1207_U7);
  not ginst4403 (P1_R1207_U24, P1_U3078);
  nand ginst4404 (P1_R1207_U240, P1_R1207_U49, P1_U3485);
  nand ginst4405 (P1_R1207_U241, P1_R1207_U123, P1_R1207_U145);
  nand ginst4406 (P1_R1207_U242, P1_R1207_U239, P1_R1207_U240);
  not ginst4407 (P1_R1207_U243, P1_R1207_U169);
  nand ginst4408 (P1_R1207_U244, P1_R1207_U53, P1_U3488);
  nand ginst4409 (P1_R1207_U245, P1_R1207_U169, P1_R1207_U244);
  nand ginst4410 (P1_R1207_U246, P1_R1207_U52, P1_U3072);
  not ginst4411 (P1_R1207_U247, P1_R1207_U168);
  nand ginst4412 (P1_R1207_U248, P1_R1207_U55, P1_U3491);
  nand ginst4413 (P1_R1207_U249, P1_R1207_U168, P1_R1207_U248);
  not ginst4414 (P1_R1207_U25, P1_U3461);
  nand ginst4415 (P1_R1207_U250, P1_R1207_U54, P1_U3080);
  not ginst4416 (P1_R1207_U251, P1_R1207_U167);
  nand ginst4417 (P1_R1207_U252, P1_R1207_U58, P1_U3500);
  nand ginst4418 (P1_R1207_U253, P1_R1207_U56, P1_U3073);
  nand ginst4419 (P1_R1207_U254, P1_R1207_U46, P1_U3074);
  nand ginst4420 (P1_R1207_U255, P1_R1207_U175, P1_R1207_U181);
  nand ginst4421 (P1_R1207_U256, P1_R1207_U255, P1_R1207_U8);
  nand ginst4422 (P1_R1207_U257, P1_R1207_U60, P1_U3494);
  nand ginst4423 (P1_R1207_U258, P1_R1207_U58, P1_U3500);
  nand ginst4424 (P1_R1207_U259, P1_R1207_U124, P1_R1207_U167);
  not ginst4425 (P1_R1207_U26, P1_U3068);
  nand ginst4426 (P1_R1207_U260, P1_R1207_U256, P1_R1207_U258);
  not ginst4427 (P1_R1207_U261, P1_R1207_U164);
  nand ginst4428 (P1_R1207_U262, P1_R1207_U63, P1_U3503);
  nand ginst4429 (P1_R1207_U263, P1_R1207_U164, P1_R1207_U262);
  nand ginst4430 (P1_R1207_U264, P1_R1207_U62, P1_U3069);
  not ginst4431 (P1_R1207_U265, P1_R1207_U64);
  nand ginst4432 (P1_R1207_U266, P1_R1207_U265, P1_R1207_U65);
  nand ginst4433 (P1_R1207_U267, P1_R1207_U163, P1_R1207_U266);
  nand ginst4434 (P1_R1207_U268, P1_R1207_U64, P1_U3082);
  not ginst4435 (P1_R1207_U269, P1_R1207_U162);
  nand ginst4436 (P1_R1207_U27, P1_R1207_U21, P1_U3068);
  nand ginst4437 (P1_R1207_U270, P1_R1207_U67, P1_U3508);
  nand ginst4438 (P1_R1207_U271, P1_R1207_U162, P1_R1207_U270);
  nand ginst4439 (P1_R1207_U272, P1_R1207_U66, P1_U3081);
  not ginst4440 (P1_R1207_U273, P1_R1207_U160);
  nand ginst4441 (P1_R1207_U274, P1_R1207_U69, P1_U3982);
  nand ginst4442 (P1_R1207_U275, P1_R1207_U160, P1_R1207_U274);
  nand ginst4443 (P1_R1207_U276, P1_R1207_U68, P1_U3076);
  not ginst4444 (P1_R1207_U277, P1_R1207_U159);
  nand ginst4445 (P1_R1207_U278, P1_R1207_U72, P1_U3979);
  nand ginst4446 (P1_R1207_U279, P1_R1207_U70, P1_U3066);
  not ginst4447 (P1_R1207_U28, P1_U3064);
  nand ginst4448 (P1_R1207_U280, P1_R1207_U45, P1_U3061);
  nand ginst4449 (P1_R1207_U281, P1_R1207_U176, P1_R1207_U182);
  nand ginst4450 (P1_R1207_U282, P1_R1207_U281, P1_R1207_U9);
  nand ginst4451 (P1_R1207_U283, P1_R1207_U74, P1_U3981);
  nand ginst4452 (P1_R1207_U284, P1_R1207_U72, P1_U3979);
  nand ginst4453 (P1_R1207_U285, P1_R1207_U125, P1_R1207_U159, P1_R1207_U278);
  nand ginst4454 (P1_R1207_U286, P1_R1207_U282, P1_R1207_U284);
  not ginst4455 (P1_R1207_U287, P1_R1207_U156);
  nand ginst4456 (P1_R1207_U288, P1_R1207_U77, P1_U3978);
  nand ginst4457 (P1_R1207_U289, P1_R1207_U156, P1_R1207_U288);
  not ginst4458 (P1_R1207_U29, P1_U3470);
  nand ginst4459 (P1_R1207_U290, P1_R1207_U76, P1_U3065);
  not ginst4460 (P1_R1207_U291, P1_R1207_U155);
  nand ginst4461 (P1_R1207_U292, P1_R1207_U79, P1_U3977);
  nand ginst4462 (P1_R1207_U293, P1_R1207_U155, P1_R1207_U292);
  nand ginst4463 (P1_R1207_U294, P1_R1207_U78, P1_U3058);
  not ginst4464 (P1_R1207_U295, P1_R1207_U87);
  nand ginst4465 (P1_R1207_U296, P1_R1207_U83, P1_U3975);
  nand ginst4466 (P1_R1207_U297, P1_R1207_U177, P1_R1207_U296, P1_R1207_U87);
  nand ginst4467 (P1_R1207_U298, P1_R1207_U82, P1_R1207_U83);
  nand ginst4468 (P1_R1207_U299, P1_R1207_U298, P1_R1207_U80);
  not ginst4469 (P1_R1207_U30, P1_U3464);
  nand ginst4470 (P1_R1207_U300, P1_R1207_U171, P1_U3053);
  not ginst4471 (P1_R1207_U301, P1_R1207_U86);
  nand ginst4472 (P1_R1207_U302, P1_R1207_U84, P1_U3054);
  nand ginst4473 (P1_R1207_U303, P1_R1207_U301, P1_R1207_U302);
  nand ginst4474 (P1_R1207_U304, P1_R1207_U85, P1_U3974);
  nand ginst4475 (P1_R1207_U305, P1_R1207_U85, P1_U3974);
  nand ginst4476 (P1_R1207_U306, P1_R1207_U305, P1_R1207_U86);
  nand ginst4477 (P1_R1207_U307, P1_R1207_U84, P1_U3054);
  nand ginst4478 (P1_R1207_U308, P1_R1207_U153, P1_R1207_U306, P1_R1207_U307);
  nand ginst4479 (P1_R1207_U309, P1_R1207_U295, P1_R1207_U82);
  not ginst4480 (P1_R1207_U31, P1_U3071);
  nand ginst4481 (P1_R1207_U310, P1_R1207_U129, P1_R1207_U309);
  nand ginst4482 (P1_R1207_U311, P1_R1207_U177, P1_R1207_U87);
  nand ginst4483 (P1_R1207_U312, P1_R1207_U128, P1_R1207_U311);
  nand ginst4484 (P1_R1207_U313, P1_R1207_U177, P1_R1207_U82);
  nand ginst4485 (P1_R1207_U314, P1_R1207_U159, P1_R1207_U283);
  not ginst4486 (P1_R1207_U315, P1_R1207_U88);
  nand ginst4487 (P1_R1207_U316, P1_R1207_U45, P1_U3061);
  nand ginst4488 (P1_R1207_U317, P1_R1207_U315, P1_R1207_U316);
  nand ginst4489 (P1_R1207_U318, P1_R1207_U132, P1_R1207_U317);
  nand ginst4490 (P1_R1207_U319, P1_R1207_U176, P1_R1207_U88);
  not ginst4491 (P1_R1207_U32, P1_U3067);
  nand ginst4492 (P1_R1207_U320, P1_R1207_U72, P1_U3979);
  nand ginst4493 (P1_R1207_U321, P1_R1207_U319, P1_R1207_U320, P1_R1207_U9);
  nand ginst4494 (P1_R1207_U322, P1_R1207_U45, P1_U3061);
  nand ginst4495 (P1_R1207_U323, P1_R1207_U176, P1_R1207_U322);
  nand ginst4496 (P1_R1207_U324, P1_R1207_U283, P1_R1207_U75);
  nand ginst4497 (P1_R1207_U325, P1_R1207_U167, P1_R1207_U257);
  not ginst4498 (P1_R1207_U326, P1_R1207_U89);
  nand ginst4499 (P1_R1207_U327, P1_R1207_U46, P1_U3074);
  nand ginst4500 (P1_R1207_U328, P1_R1207_U326, P1_R1207_U327);
  nand ginst4501 (P1_R1207_U329, P1_R1207_U139, P1_R1207_U328);
  not ginst4502 (P1_R1207_U33, P1_U3060);
  nand ginst4503 (P1_R1207_U330, P1_R1207_U175, P1_R1207_U89);
  nand ginst4504 (P1_R1207_U331, P1_R1207_U58, P1_U3500);
  nand ginst4505 (P1_R1207_U332, P1_R1207_U138, P1_R1207_U330);
  nand ginst4506 (P1_R1207_U333, P1_R1207_U46, P1_U3074);
  nand ginst4507 (P1_R1207_U334, P1_R1207_U175, P1_R1207_U333);
  nand ginst4508 (P1_R1207_U335, P1_R1207_U257, P1_R1207_U61);
  nand ginst4509 (P1_R1207_U336, P1_R1207_U145, P1_R1207_U212);
  not ginst4510 (P1_R1207_U337, P1_R1207_U90);
  nand ginst4511 (P1_R1207_U338, P1_R1207_U47, P1_U3062);
  nand ginst4512 (P1_R1207_U339, P1_R1207_U337, P1_R1207_U338);
  nand ginst4513 (P1_R1207_U34, P1_R1207_U30, P1_U3060);
  nand ginst4514 (P1_R1207_U340, P1_R1207_U143, P1_R1207_U339);
  nand ginst4515 (P1_R1207_U341, P1_R1207_U174, P1_R1207_U90);
  nand ginst4516 (P1_R1207_U342, P1_R1207_U49, P1_U3485);
  nand ginst4517 (P1_R1207_U343, P1_R1207_U142, P1_R1207_U341);
  nand ginst4518 (P1_R1207_U344, P1_R1207_U47, P1_U3062);
  nand ginst4519 (P1_R1207_U345, P1_R1207_U174, P1_R1207_U344);
  nand ginst4520 (P1_R1207_U346, P1_R1207_U22, P1_U3077);
  nand ginst4521 (P1_R1207_U347, P1_R1207_U303, P1_R1207_U304, P1_R1207_U385);
  nand ginst4522 (P1_R1207_U348, P1_R1207_U40, P1_U3479);
  nand ginst4523 (P1_R1207_U349, P1_R1207_U39, P1_U3083);
  not ginst4524 (P1_R1207_U35, P1_U3476);
  nand ginst4525 (P1_R1207_U350, P1_R1207_U145, P1_R1207_U213);
  nand ginst4526 (P1_R1207_U351, P1_R1207_U144, P1_R1207_U211);
  nand ginst4527 (P1_R1207_U352, P1_R1207_U38, P1_U3476);
  nand ginst4528 (P1_R1207_U353, P1_R1207_U35, P1_U3084);
  nand ginst4529 (P1_R1207_U354, P1_R1207_U38, P1_U3476);
  nand ginst4530 (P1_R1207_U355, P1_R1207_U35, P1_U3084);
  nand ginst4531 (P1_R1207_U356, P1_R1207_U354, P1_R1207_U355);
  nand ginst4532 (P1_R1207_U357, P1_R1207_U36, P1_U3473);
  nand ginst4533 (P1_R1207_U358, P1_R1207_U19, P1_U3070);
  nand ginst4534 (P1_R1207_U359, P1_R1207_U218, P1_R1207_U41);
  not ginst4535 (P1_R1207_U36, P1_U3070);
  nand ginst4536 (P1_R1207_U360, P1_R1207_U146, P1_R1207_U205);
  nand ginst4537 (P1_R1207_U361, P1_R1207_U31, P1_U3470);
  nand ginst4538 (P1_R1207_U362, P1_R1207_U29, P1_U3071);
  nand ginst4539 (P1_R1207_U363, P1_R1207_U361, P1_R1207_U362);
  nand ginst4540 (P1_R1207_U364, P1_R1207_U32, P1_U3467);
  nand ginst4541 (P1_R1207_U365, P1_R1207_U20, P1_U3067);
  nand ginst4542 (P1_R1207_U366, P1_R1207_U228, P1_R1207_U42);
  nand ginst4543 (P1_R1207_U367, P1_R1207_U147, P1_R1207_U220);
  nand ginst4544 (P1_R1207_U368, P1_R1207_U33, P1_U3464);
  nand ginst4545 (P1_R1207_U369, P1_R1207_U30, P1_U3060);
  nand ginst4546 (P1_R1207_U37, P1_R1207_U19, P1_U3070);
  nand ginst4547 (P1_R1207_U370, P1_R1207_U149, P1_R1207_U229);
  nand ginst4548 (P1_R1207_U371, P1_R1207_U148, P1_R1207_U195);
  nand ginst4549 (P1_R1207_U372, P1_R1207_U28, P1_U3461);
  nand ginst4550 (P1_R1207_U373, P1_R1207_U25, P1_U3064);
  nand ginst4551 (P1_R1207_U374, P1_R1207_U28, P1_U3461);
  nand ginst4552 (P1_R1207_U375, P1_R1207_U25, P1_U3064);
  nand ginst4553 (P1_R1207_U376, P1_R1207_U374, P1_R1207_U375);
  nand ginst4554 (P1_R1207_U377, P1_R1207_U26, P1_U3458);
  nand ginst4555 (P1_R1207_U378, P1_R1207_U21, P1_U3068);
  nand ginst4556 (P1_R1207_U379, P1_R1207_U234, P1_R1207_U43);
  not ginst4557 (P1_R1207_U38, P1_U3084);
  nand ginst4558 (P1_R1207_U380, P1_R1207_U150, P1_R1207_U189);
  nand ginst4559 (P1_R1207_U381, P1_R1207_U152, P1_U3985);
  nand ginst4560 (P1_R1207_U382, P1_R1207_U151, P1_U3055);
  nand ginst4561 (P1_R1207_U383, P1_R1207_U152, P1_U3985);
  nand ginst4562 (P1_R1207_U384, P1_R1207_U151, P1_U3055);
  nand ginst4563 (P1_R1207_U385, P1_R1207_U383, P1_R1207_U384);
  nand ginst4564 (P1_R1207_U386, P1_R1207_U85, P1_U3974);
  nand ginst4565 (P1_R1207_U387, P1_R1207_U84, P1_U3054);
  not ginst4566 (P1_R1207_U388, P1_R1207_U127);
  nand ginst4567 (P1_R1207_U389, P1_R1207_U301, P1_R1207_U388);
  not ginst4568 (P1_R1207_U39, P1_U3479);
  nand ginst4569 (P1_R1207_U390, P1_R1207_U127, P1_R1207_U86);
  nand ginst4570 (P1_R1207_U391, P1_R1207_U83, P1_U3975);
  nand ginst4571 (P1_R1207_U392, P1_R1207_U80, P1_U3053);
  nand ginst4572 (P1_R1207_U393, P1_R1207_U83, P1_U3975);
  nand ginst4573 (P1_R1207_U394, P1_R1207_U80, P1_U3053);
  nand ginst4574 (P1_R1207_U395, P1_R1207_U393, P1_R1207_U394);
  nand ginst4575 (P1_R1207_U396, P1_R1207_U81, P1_U3976);
  nand ginst4576 (P1_R1207_U397, P1_R1207_U44, P1_U3057);
  nand ginst4577 (P1_R1207_U398, P1_R1207_U313, P1_R1207_U87);
  nand ginst4578 (P1_R1207_U399, P1_R1207_U154, P1_R1207_U295);
  not ginst4579 (P1_R1207_U40, P1_U3083);
  nand ginst4580 (P1_R1207_U400, P1_R1207_U79, P1_U3977);
  nand ginst4581 (P1_R1207_U401, P1_R1207_U78, P1_U3058);
  not ginst4582 (P1_R1207_U402, P1_R1207_U130);
  nand ginst4583 (P1_R1207_U403, P1_R1207_U291, P1_R1207_U402);
  nand ginst4584 (P1_R1207_U404, P1_R1207_U130, P1_R1207_U155);
  nand ginst4585 (P1_R1207_U405, P1_R1207_U77, P1_U3978);
  nand ginst4586 (P1_R1207_U406, P1_R1207_U76, P1_U3065);
  not ginst4587 (P1_R1207_U407, P1_R1207_U131);
  nand ginst4588 (P1_R1207_U408, P1_R1207_U287, P1_R1207_U407);
  nand ginst4589 (P1_R1207_U409, P1_R1207_U131, P1_R1207_U156);
  nand ginst4590 (P1_R1207_U41, P1_R1207_U203, P1_R1207_U204);
  nand ginst4591 (P1_R1207_U410, P1_R1207_U72, P1_U3979);
  nand ginst4592 (P1_R1207_U411, P1_R1207_U70, P1_U3066);
  nand ginst4593 (P1_R1207_U412, P1_R1207_U410, P1_R1207_U411);
  nand ginst4594 (P1_R1207_U413, P1_R1207_U73, P1_U3980);
  nand ginst4595 (P1_R1207_U414, P1_R1207_U45, P1_U3061);
  nand ginst4596 (P1_R1207_U415, P1_R1207_U323, P1_R1207_U88);
  nand ginst4597 (P1_R1207_U416, P1_R1207_U157, P1_R1207_U315);
  nand ginst4598 (P1_R1207_U417, P1_R1207_U74, P1_U3981);
  nand ginst4599 (P1_R1207_U418, P1_R1207_U71, P1_U3075);
  nand ginst4600 (P1_R1207_U419, P1_R1207_U159, P1_R1207_U324);
  nand ginst4601 (P1_R1207_U42, P1_R1207_U219, P1_R1207_U34);
  nand ginst4602 (P1_R1207_U420, P1_R1207_U158, P1_R1207_U277);
  nand ginst4603 (P1_R1207_U421, P1_R1207_U69, P1_U3982);
  nand ginst4604 (P1_R1207_U422, P1_R1207_U68, P1_U3076);
  not ginst4605 (P1_R1207_U423, P1_R1207_U133);
  nand ginst4606 (P1_R1207_U424, P1_R1207_U273, P1_R1207_U423);
  nand ginst4607 (P1_R1207_U425, P1_R1207_U133, P1_R1207_U160);
  nand ginst4608 (P1_R1207_U426, P1_R1207_U185, P1_R1207_U24);
  nand ginst4609 (P1_R1207_U427, P1_R1207_U23, P1_U3078);
  not ginst4610 (P1_R1207_U428, P1_R1207_U134);
  nand ginst4611 (P1_R1207_U429, P1_R1207_U428, P1_U3455);
  nand ginst4612 (P1_R1207_U43, P1_R1207_U187, P1_R1207_U188);
  nand ginst4613 (P1_R1207_U430, P1_R1207_U134, P1_R1207_U161);
  nand ginst4614 (P1_R1207_U431, P1_R1207_U67, P1_U3508);
  nand ginst4615 (P1_R1207_U432, P1_R1207_U66, P1_U3081);
  not ginst4616 (P1_R1207_U433, P1_R1207_U135);
  nand ginst4617 (P1_R1207_U434, P1_R1207_U269, P1_R1207_U433);
  nand ginst4618 (P1_R1207_U435, P1_R1207_U135, P1_R1207_U162);
  nand ginst4619 (P1_R1207_U436, P1_R1207_U65, P1_U3506);
  nand ginst4620 (P1_R1207_U437, P1_R1207_U163, P1_U3082);
  not ginst4621 (P1_R1207_U438, P1_R1207_U136);
  nand ginst4622 (P1_R1207_U439, P1_R1207_U265, P1_R1207_U438);
  not ginst4623 (P1_R1207_U44, P1_U3976);
  nand ginst4624 (P1_R1207_U440, P1_R1207_U136, P1_R1207_U64);
  nand ginst4625 (P1_R1207_U441, P1_R1207_U63, P1_U3503);
  nand ginst4626 (P1_R1207_U442, P1_R1207_U62, P1_U3069);
  not ginst4627 (P1_R1207_U443, P1_R1207_U137);
  nand ginst4628 (P1_R1207_U444, P1_R1207_U261, P1_R1207_U443);
  nand ginst4629 (P1_R1207_U445, P1_R1207_U137, P1_R1207_U164);
  nand ginst4630 (P1_R1207_U446, P1_R1207_U58, P1_U3500);
  nand ginst4631 (P1_R1207_U447, P1_R1207_U56, P1_U3073);
  nand ginst4632 (P1_R1207_U448, P1_R1207_U446, P1_R1207_U447);
  nand ginst4633 (P1_R1207_U449, P1_R1207_U59, P1_U3497);
  not ginst4634 (P1_R1207_U45, P1_U3980);
  nand ginst4635 (P1_R1207_U450, P1_R1207_U46, P1_U3074);
  nand ginst4636 (P1_R1207_U451, P1_R1207_U334, P1_R1207_U89);
  nand ginst4637 (P1_R1207_U452, P1_R1207_U165, P1_R1207_U326);
  nand ginst4638 (P1_R1207_U453, P1_R1207_U60, P1_U3494);
  nand ginst4639 (P1_R1207_U454, P1_R1207_U57, P1_U3079);
  nand ginst4640 (P1_R1207_U455, P1_R1207_U167, P1_R1207_U335);
  nand ginst4641 (P1_R1207_U456, P1_R1207_U166, P1_R1207_U251);
  nand ginst4642 (P1_R1207_U457, P1_R1207_U55, P1_U3491);
  nand ginst4643 (P1_R1207_U458, P1_R1207_U54, P1_U3080);
  not ginst4644 (P1_R1207_U459, P1_R1207_U140);
  not ginst4645 (P1_R1207_U46, P1_U3497);
  nand ginst4646 (P1_R1207_U460, P1_R1207_U247, P1_R1207_U459);
  nand ginst4647 (P1_R1207_U461, P1_R1207_U140, P1_R1207_U168);
  nand ginst4648 (P1_R1207_U462, P1_R1207_U53, P1_U3488);
  nand ginst4649 (P1_R1207_U463, P1_R1207_U52, P1_U3072);
  not ginst4650 (P1_R1207_U464, P1_R1207_U141);
  nand ginst4651 (P1_R1207_U465, P1_R1207_U243, P1_R1207_U464);
  nand ginst4652 (P1_R1207_U466, P1_R1207_U141, P1_R1207_U169);
  nand ginst4653 (P1_R1207_U467, P1_R1207_U49, P1_U3485);
  nand ginst4654 (P1_R1207_U468, P1_R1207_U48, P1_U3063);
  nand ginst4655 (P1_R1207_U469, P1_R1207_U467, P1_R1207_U468);
  not ginst4656 (P1_R1207_U47, P1_U3482);
  nand ginst4657 (P1_R1207_U470, P1_R1207_U50, P1_U3482);
  nand ginst4658 (P1_R1207_U471, P1_R1207_U47, P1_U3062);
  nand ginst4659 (P1_R1207_U472, P1_R1207_U345, P1_R1207_U90);
  nand ginst4660 (P1_R1207_U473, P1_R1207_U170, P1_R1207_U337);
  not ginst4661 (P1_R1207_U48, P1_U3485);
  not ginst4662 (P1_R1207_U49, P1_U3063);
  not ginst4663 (P1_R1207_U50, P1_U3062);
  nand ginst4664 (P1_R1207_U51, P1_R1207_U39, P1_U3083);
  not ginst4665 (P1_R1207_U52, P1_U3488);
  not ginst4666 (P1_R1207_U53, P1_U3072);
  not ginst4667 (P1_R1207_U54, P1_U3491);
  not ginst4668 (P1_R1207_U55, P1_U3080);
  not ginst4669 (P1_R1207_U56, P1_U3500);
  not ginst4670 (P1_R1207_U57, P1_U3494);
  not ginst4671 (P1_R1207_U58, P1_U3073);
  not ginst4672 (P1_R1207_U59, P1_U3074);
  and ginst4673 (P1_R1207_U6, P1_R1207_U197, P1_R1207_U198);
  not ginst4674 (P1_R1207_U60, P1_U3079);
  nand ginst4675 (P1_R1207_U61, P1_R1207_U57, P1_U3079);
  not ginst4676 (P1_R1207_U62, P1_U3503);
  not ginst4677 (P1_R1207_U63, P1_U3069);
  nand ginst4678 (P1_R1207_U64, P1_R1207_U263, P1_R1207_U264);
  not ginst4679 (P1_R1207_U65, P1_U3082);
  not ginst4680 (P1_R1207_U66, P1_U3508);
  not ginst4681 (P1_R1207_U67, P1_U3081);
  not ginst4682 (P1_R1207_U68, P1_U3982);
  not ginst4683 (P1_R1207_U69, P1_U3076);
  and ginst4684 (P1_R1207_U7, P1_R1207_U236, P1_R1207_U237);
  not ginst4685 (P1_R1207_U70, P1_U3979);
  not ginst4686 (P1_R1207_U71, P1_U3981);
  not ginst4687 (P1_R1207_U72, P1_U3066);
  not ginst4688 (P1_R1207_U73, P1_U3061);
  not ginst4689 (P1_R1207_U74, P1_U3075);
  nand ginst4690 (P1_R1207_U75, P1_R1207_U71, P1_U3075);
  not ginst4691 (P1_R1207_U76, P1_U3978);
  not ginst4692 (P1_R1207_U77, P1_U3065);
  not ginst4693 (P1_R1207_U78, P1_U3977);
  not ginst4694 (P1_R1207_U79, P1_U3058);
  and ginst4695 (P1_R1207_U8, P1_R1207_U253, P1_R1207_U254);
  not ginst4696 (P1_R1207_U80, P1_U3975);
  not ginst4697 (P1_R1207_U81, P1_U3057);
  nand ginst4698 (P1_R1207_U82, P1_R1207_U44, P1_U3057);
  not ginst4699 (P1_R1207_U83, P1_U3053);
  not ginst4700 (P1_R1207_U84, P1_U3974);
  not ginst4701 (P1_R1207_U85, P1_U3054);
  nand ginst4702 (P1_R1207_U86, P1_R1207_U126, P1_R1207_U297);
  nand ginst4703 (P1_R1207_U87, P1_R1207_U293, P1_R1207_U294);
  nand ginst4704 (P1_R1207_U88, P1_R1207_U314, P1_R1207_U75);
  nand ginst4705 (P1_R1207_U89, P1_R1207_U325, P1_R1207_U61);
  and ginst4706 (P1_R1207_U9, P1_R1207_U279, P1_R1207_U280);
  nand ginst4707 (P1_R1207_U90, P1_R1207_U336, P1_R1207_U51);
  not ginst4708 (P1_R1207_U91, P1_U3077);
  nand ginst4709 (P1_R1207_U92, P1_R1207_U389, P1_R1207_U390);
  nand ginst4710 (P1_R1207_U93, P1_R1207_U403, P1_R1207_U404);
  nand ginst4711 (P1_R1207_U94, P1_R1207_U408, P1_R1207_U409);
  nand ginst4712 (P1_R1207_U95, P1_R1207_U424, P1_R1207_U425);
  nand ginst4713 (P1_R1207_U96, P1_R1207_U429, P1_R1207_U430);
  nand ginst4714 (P1_R1207_U97, P1_R1207_U434, P1_R1207_U435);
  nand ginst4715 (P1_R1207_U98, P1_R1207_U439, P1_R1207_U440);
  nand ginst4716 (P1_R1207_U99, P1_R1207_U444, P1_R1207_U445);
  and ginst4717 (P1_R1222_U10, P1_R1222_U270, P1_R1222_U271);
  nand ginst4718 (P1_R1222_U100, P1_R1222_U392, P1_R1222_U393);
  nand ginst4719 (P1_R1222_U101, P1_R1222_U397, P1_R1222_U398);
  nand ginst4720 (P1_R1222_U102, P1_R1222_U406, P1_R1222_U407);
  nand ginst4721 (P1_R1222_U103, P1_R1222_U413, P1_R1222_U414);
  nand ginst4722 (P1_R1222_U104, P1_R1222_U420, P1_R1222_U421);
  nand ginst4723 (P1_R1222_U105, P1_R1222_U427, P1_R1222_U428);
  nand ginst4724 (P1_R1222_U106, P1_R1222_U432, P1_R1222_U433);
  nand ginst4725 (P1_R1222_U107, P1_R1222_U439, P1_R1222_U440);
  nand ginst4726 (P1_R1222_U108, P1_R1222_U446, P1_R1222_U447);
  nand ginst4727 (P1_R1222_U109, P1_R1222_U460, P1_R1222_U461);
  and ginst4728 (P1_R1222_U11, P1_R1222_U347, P1_R1222_U350);
  nand ginst4729 (P1_R1222_U110, P1_R1222_U465, P1_R1222_U466);
  nand ginst4730 (P1_R1222_U111, P1_R1222_U472, P1_R1222_U473);
  nand ginst4731 (P1_R1222_U112, P1_R1222_U479, P1_R1222_U480);
  nand ginst4732 (P1_R1222_U113, P1_R1222_U486, P1_R1222_U487);
  nand ginst4733 (P1_R1222_U114, P1_R1222_U493, P1_R1222_U494);
  nand ginst4734 (P1_R1222_U115, P1_R1222_U498, P1_R1222_U499);
  and ginst4735 (P1_R1222_U116, P1_U3068, P1_U3458);
  and ginst4736 (P1_R1222_U117, P1_R1222_U186, P1_R1222_U188);
  and ginst4737 (P1_R1222_U118, P1_R1222_U191, P1_R1222_U193);
  and ginst4738 (P1_R1222_U119, P1_R1222_U199, P1_R1222_U200);
  and ginst4739 (P1_R1222_U12, P1_R1222_U340, P1_R1222_U343);
  and ginst4740 (P1_R1222_U120, P1_R1222_U23, P1_R1222_U380, P1_R1222_U381);
  and ginst4741 (P1_R1222_U121, P1_R1222_U211, P1_R1222_U6);
  and ginst4742 (P1_R1222_U122, P1_R1222_U217, P1_R1222_U219);
  and ginst4743 (P1_R1222_U123, P1_R1222_U35, P1_R1222_U387, P1_R1222_U388);
  and ginst4744 (P1_R1222_U124, P1_R1222_U225, P1_R1222_U4);
  and ginst4745 (P1_R1222_U125, P1_R1222_U180, P1_R1222_U233);
  and ginst4746 (P1_R1222_U126, P1_R1222_U203, P1_R1222_U7);
  and ginst4747 (P1_R1222_U127, P1_R1222_U170, P1_R1222_U238);
  and ginst4748 (P1_R1222_U128, P1_R1222_U249, P1_R1222_U8);
  and ginst4749 (P1_R1222_U129, P1_R1222_U171, P1_R1222_U247);
  and ginst4750 (P1_R1222_U13, P1_R1222_U331, P1_R1222_U334);
  and ginst4751 (P1_R1222_U130, P1_R1222_U266, P1_R1222_U267);
  and ginst4752 (P1_R1222_U131, P1_R1222_U10, P1_R1222_U281);
  and ginst4753 (P1_R1222_U132, P1_R1222_U279, P1_R1222_U284);
  and ginst4754 (P1_R1222_U133, P1_R1222_U297, P1_R1222_U300);
  and ginst4755 (P1_R1222_U134, P1_R1222_U301, P1_R1222_U367);
  and ginst4756 (P1_R1222_U135, P1_R1222_U159, P1_R1222_U277);
  and ginst4757 (P1_R1222_U136, P1_R1222_U453, P1_R1222_U454, P1_R1222_U81);
  and ginst4758 (P1_R1222_U137, P1_R1222_U467, P1_R1222_U468, P1_R1222_U60);
  and ginst4759 (P1_R1222_U138, P1_R1222_U333, P1_R1222_U9);
  and ginst4760 (P1_R1222_U139, P1_R1222_U171, P1_R1222_U488, P1_R1222_U489);
  and ginst4761 (P1_R1222_U14, P1_R1222_U322, P1_R1222_U325);
  and ginst4762 (P1_R1222_U140, P1_R1222_U342, P1_R1222_U8);
  and ginst4763 (P1_R1222_U141, P1_R1222_U170, P1_R1222_U500, P1_R1222_U501);
  and ginst4764 (P1_R1222_U142, P1_R1222_U349, P1_R1222_U7);
  nand ginst4765 (P1_R1222_U143, P1_R1222_U119, P1_R1222_U201);
  nand ginst4766 (P1_R1222_U144, P1_R1222_U216, P1_R1222_U228);
  not ginst4767 (P1_R1222_U145, P1_U3055);
  not ginst4768 (P1_R1222_U146, P1_U3985);
  and ginst4769 (P1_R1222_U147, P1_R1222_U401, P1_R1222_U402);
  nand ginst4770 (P1_R1222_U148, P1_R1222_U168, P1_R1222_U303, P1_R1222_U363);
  and ginst4771 (P1_R1222_U149, P1_R1222_U408, P1_R1222_U409);
  and ginst4772 (P1_R1222_U15, P1_R1222_U317, P1_R1222_U319);
  nand ginst4773 (P1_R1222_U150, P1_R1222_U134, P1_R1222_U368, P1_R1222_U369);
  and ginst4774 (P1_R1222_U151, P1_R1222_U415, P1_R1222_U416);
  nand ginst4775 (P1_R1222_U152, P1_R1222_U298, P1_R1222_U364, P1_R1222_U87);
  and ginst4776 (P1_R1222_U153, P1_R1222_U422, P1_R1222_U423);
  nand ginst4777 (P1_R1222_U154, P1_R1222_U291, P1_R1222_U292);
  and ginst4778 (P1_R1222_U155, P1_R1222_U434, P1_R1222_U435);
  nand ginst4779 (P1_R1222_U156, P1_R1222_U287, P1_R1222_U288);
  and ginst4780 (P1_R1222_U157, P1_R1222_U441, P1_R1222_U442);
  nand ginst4781 (P1_R1222_U158, P1_R1222_U132, P1_R1222_U283);
  and ginst4782 (P1_R1222_U159, P1_R1222_U448, P1_R1222_U449);
  and ginst4783 (P1_R1222_U16, P1_R1222_U309, P1_R1222_U312);
  nand ginst4784 (P1_R1222_U160, P1_R1222_U326, P1_R1222_U44);
  nand ginst4785 (P1_R1222_U161, P1_R1222_U130, P1_R1222_U268);
  and ginst4786 (P1_R1222_U162, P1_R1222_U474, P1_R1222_U475);
  nand ginst4787 (P1_R1222_U163, P1_R1222_U255, P1_R1222_U256);
  and ginst4788 (P1_R1222_U164, P1_R1222_U481, P1_R1222_U482);
  nand ginst4789 (P1_R1222_U165, P1_R1222_U251, P1_R1222_U252);
  nand ginst4790 (P1_R1222_U166, P1_R1222_U241, P1_R1222_U242);
  nand ginst4791 (P1_R1222_U167, P1_R1222_U365, P1_R1222_U366);
  nand ginst4792 (P1_R1222_U168, P1_R1222_U150, P1_U3054);
  not ginst4793 (P1_R1222_U169, P1_R1222_U35);
  and ginst4794 (P1_R1222_U17, P1_R1222_U231, P1_R1222_U234);
  nand ginst4795 (P1_R1222_U170, P1_U3083, P1_U3479);
  nand ginst4796 (P1_R1222_U171, P1_U3072, P1_U3488);
  nand ginst4797 (P1_R1222_U172, P1_U3058, P1_U3977);
  not ginst4798 (P1_R1222_U173, P1_R1222_U69);
  not ginst4799 (P1_R1222_U174, P1_R1222_U78);
  nand ginst4800 (P1_R1222_U175, P1_U3065, P1_U3978);
  not ginst4801 (P1_R1222_U176, P1_R1222_U62);
  or ginst4802 (P1_R1222_U177, P1_U3067, P1_U3467);
  or ginst4803 (P1_R1222_U178, P1_U3060, P1_U3464);
  or ginst4804 (P1_R1222_U179, P1_U3064, P1_U3461);
  and ginst4805 (P1_R1222_U18, P1_R1222_U223, P1_R1222_U226);
  or ginst4806 (P1_R1222_U180, P1_U3068, P1_U3458);
  not ginst4807 (P1_R1222_U181, P1_R1222_U32);
  or ginst4808 (P1_R1222_U182, P1_U3078, P1_U3455);
  not ginst4809 (P1_R1222_U183, P1_R1222_U43);
  not ginst4810 (P1_R1222_U184, P1_R1222_U44);
  nand ginst4811 (P1_R1222_U185, P1_R1222_U43, P1_R1222_U44);
  nand ginst4812 (P1_R1222_U186, P1_R1222_U116, P1_R1222_U179);
  nand ginst4813 (P1_R1222_U187, P1_R1222_U185, P1_R1222_U5);
  nand ginst4814 (P1_R1222_U188, P1_U3064, P1_U3461);
  nand ginst4815 (P1_R1222_U189, P1_R1222_U117, P1_R1222_U187);
  and ginst4816 (P1_R1222_U19, P1_R1222_U209, P1_R1222_U212);
  nand ginst4817 (P1_R1222_U190, P1_R1222_U35, P1_R1222_U36);
  nand ginst4818 (P1_R1222_U191, P1_R1222_U190, P1_U3067);
  nand ginst4819 (P1_R1222_U192, P1_R1222_U189, P1_R1222_U4);
  nand ginst4820 (P1_R1222_U193, P1_R1222_U169, P1_U3467);
  not ginst4821 (P1_R1222_U194, P1_R1222_U42);
  or ginst4822 (P1_R1222_U195, P1_U3070, P1_U3473);
  or ginst4823 (P1_R1222_U196, P1_U3071, P1_U3470);
  not ginst4824 (P1_R1222_U197, P1_R1222_U23);
  nand ginst4825 (P1_R1222_U198, P1_R1222_U23, P1_R1222_U24);
  nand ginst4826 (P1_R1222_U199, P1_R1222_U198, P1_U3070);
  not ginst4827 (P1_R1222_U20, P1_U3470);
  nand ginst4828 (P1_R1222_U200, P1_R1222_U197, P1_U3473);
  nand ginst4829 (P1_R1222_U201, P1_R1222_U42, P1_R1222_U6);
  not ginst4830 (P1_R1222_U202, P1_R1222_U143);
  or ginst4831 (P1_R1222_U203, P1_U3084, P1_U3476);
  nand ginst4832 (P1_R1222_U204, P1_R1222_U143, P1_R1222_U203);
  not ginst4833 (P1_R1222_U205, P1_R1222_U41);
  or ginst4834 (P1_R1222_U206, P1_U3083, P1_U3479);
  or ginst4835 (P1_R1222_U207, P1_U3071, P1_U3470);
  nand ginst4836 (P1_R1222_U208, P1_R1222_U207, P1_R1222_U42);
  nand ginst4837 (P1_R1222_U209, P1_R1222_U120, P1_R1222_U208);
  not ginst4838 (P1_R1222_U21, P1_U3071);
  nand ginst4839 (P1_R1222_U210, P1_R1222_U194, P1_R1222_U23);
  nand ginst4840 (P1_R1222_U211, P1_U3070, P1_U3473);
  nand ginst4841 (P1_R1222_U212, P1_R1222_U121, P1_R1222_U210);
  or ginst4842 (P1_R1222_U213, P1_U3071, P1_U3470);
  nand ginst4843 (P1_R1222_U214, P1_R1222_U180, P1_R1222_U184);
  nand ginst4844 (P1_R1222_U215, P1_U3068, P1_U3458);
  not ginst4845 (P1_R1222_U216, P1_R1222_U46);
  nand ginst4846 (P1_R1222_U217, P1_R1222_U183, P1_R1222_U5);
  nand ginst4847 (P1_R1222_U218, P1_R1222_U179, P1_R1222_U46);
  nand ginst4848 (P1_R1222_U219, P1_U3064, P1_U3461);
  not ginst4849 (P1_R1222_U22, P1_U3070);
  not ginst4850 (P1_R1222_U220, P1_R1222_U45);
  or ginst4851 (P1_R1222_U221, P1_U3060, P1_U3464);
  nand ginst4852 (P1_R1222_U222, P1_R1222_U221, P1_R1222_U45);
  nand ginst4853 (P1_R1222_U223, P1_R1222_U123, P1_R1222_U222);
  nand ginst4854 (P1_R1222_U224, P1_R1222_U220, P1_R1222_U35);
  nand ginst4855 (P1_R1222_U225, P1_U3067, P1_U3467);
  nand ginst4856 (P1_R1222_U226, P1_R1222_U124, P1_R1222_U224);
  or ginst4857 (P1_R1222_U227, P1_U3060, P1_U3464);
  nand ginst4858 (P1_R1222_U228, P1_R1222_U180, P1_R1222_U183);
  not ginst4859 (P1_R1222_U229, P1_R1222_U144);
  nand ginst4860 (P1_R1222_U23, P1_U3071, P1_U3470);
  nand ginst4861 (P1_R1222_U230, P1_U3064, P1_U3461);
  nand ginst4862 (P1_R1222_U231, P1_R1222_U399, P1_R1222_U400, P1_R1222_U43, P1_R1222_U44);
  nand ginst4863 (P1_R1222_U232, P1_R1222_U43, P1_R1222_U44);
  nand ginst4864 (P1_R1222_U233, P1_U3068, P1_U3458);
  nand ginst4865 (P1_R1222_U234, P1_R1222_U125, P1_R1222_U232);
  or ginst4866 (P1_R1222_U235, P1_U3083, P1_U3479);
  or ginst4867 (P1_R1222_U236, P1_U3062, P1_U3482);
  nand ginst4868 (P1_R1222_U237, P1_R1222_U176, P1_R1222_U7);
  nand ginst4869 (P1_R1222_U238, P1_U3062, P1_U3482);
  nand ginst4870 (P1_R1222_U239, P1_R1222_U127, P1_R1222_U237);
  not ginst4871 (P1_R1222_U24, P1_U3473);
  or ginst4872 (P1_R1222_U240, P1_U3062, P1_U3482);
  nand ginst4873 (P1_R1222_U241, P1_R1222_U126, P1_R1222_U143);
  nand ginst4874 (P1_R1222_U242, P1_R1222_U239, P1_R1222_U240);
  not ginst4875 (P1_R1222_U243, P1_R1222_U166);
  or ginst4876 (P1_R1222_U244, P1_U3080, P1_U3491);
  or ginst4877 (P1_R1222_U245, P1_U3072, P1_U3488);
  nand ginst4878 (P1_R1222_U246, P1_R1222_U173, P1_R1222_U8);
  nand ginst4879 (P1_R1222_U247, P1_U3080, P1_U3491);
  nand ginst4880 (P1_R1222_U248, P1_R1222_U129, P1_R1222_U246);
  or ginst4881 (P1_R1222_U249, P1_U3063, P1_U3485);
  not ginst4882 (P1_R1222_U25, P1_U3464);
  or ginst4883 (P1_R1222_U250, P1_U3080, P1_U3491);
  nand ginst4884 (P1_R1222_U251, P1_R1222_U128, P1_R1222_U166);
  nand ginst4885 (P1_R1222_U252, P1_R1222_U248, P1_R1222_U250);
  not ginst4886 (P1_R1222_U253, P1_R1222_U165);
  or ginst4887 (P1_R1222_U254, P1_U3079, P1_U3494);
  nand ginst4888 (P1_R1222_U255, P1_R1222_U165, P1_R1222_U254);
  nand ginst4889 (P1_R1222_U256, P1_U3079, P1_U3494);
  not ginst4890 (P1_R1222_U257, P1_R1222_U163);
  or ginst4891 (P1_R1222_U258, P1_U3074, P1_U3497);
  nand ginst4892 (P1_R1222_U259, P1_R1222_U163, P1_R1222_U258);
  not ginst4893 (P1_R1222_U26, P1_U3060);
  nand ginst4894 (P1_R1222_U260, P1_U3074, P1_U3497);
  not ginst4895 (P1_R1222_U261, P1_R1222_U93);
  or ginst4896 (P1_R1222_U262, P1_U3069, P1_U3503);
  or ginst4897 (P1_R1222_U263, P1_U3073, P1_U3500);
  not ginst4898 (P1_R1222_U264, P1_R1222_U60);
  nand ginst4899 (P1_R1222_U265, P1_R1222_U60, P1_R1222_U61);
  nand ginst4900 (P1_R1222_U266, P1_R1222_U265, P1_U3069);
  nand ginst4901 (P1_R1222_U267, P1_R1222_U264, P1_U3503);
  nand ginst4902 (P1_R1222_U268, P1_R1222_U9, P1_R1222_U93);
  not ginst4903 (P1_R1222_U269, P1_R1222_U161);
  not ginst4904 (P1_R1222_U27, P1_U3067);
  or ginst4905 (P1_R1222_U270, P1_U3076, P1_U3982);
  or ginst4906 (P1_R1222_U271, P1_U3081, P1_U3508);
  or ginst4907 (P1_R1222_U272, P1_U3075, P1_U3981);
  not ginst4908 (P1_R1222_U273, P1_R1222_U81);
  nand ginst4909 (P1_R1222_U274, P1_R1222_U273, P1_U3982);
  nand ginst4910 (P1_R1222_U275, P1_R1222_U274, P1_R1222_U91);
  nand ginst4911 (P1_R1222_U276, P1_R1222_U81, P1_R1222_U82);
  nand ginst4912 (P1_R1222_U277, P1_R1222_U275, P1_R1222_U276);
  nand ginst4913 (P1_R1222_U278, P1_R1222_U10, P1_R1222_U174);
  nand ginst4914 (P1_R1222_U279, P1_U3075, P1_U3981);
  not ginst4915 (P1_R1222_U28, P1_U3458);
  nand ginst4916 (P1_R1222_U280, P1_R1222_U277, P1_R1222_U278);
  or ginst4917 (P1_R1222_U281, P1_U3082, P1_U3506);
  or ginst4918 (P1_R1222_U282, P1_U3075, P1_U3981);
  nand ginst4919 (P1_R1222_U283, P1_R1222_U131, P1_R1222_U161, P1_R1222_U272);
  nand ginst4920 (P1_R1222_U284, P1_R1222_U280, P1_R1222_U282);
  not ginst4921 (P1_R1222_U285, P1_R1222_U158);
  or ginst4922 (P1_R1222_U286, P1_U3061, P1_U3980);
  nand ginst4923 (P1_R1222_U287, P1_R1222_U158, P1_R1222_U286);
  nand ginst4924 (P1_R1222_U288, P1_U3061, P1_U3980);
  not ginst4925 (P1_R1222_U289, P1_R1222_U156);
  not ginst4926 (P1_R1222_U29, P1_U3068);
  or ginst4927 (P1_R1222_U290, P1_U3066, P1_U3979);
  nand ginst4928 (P1_R1222_U291, P1_R1222_U156, P1_R1222_U290);
  nand ginst4929 (P1_R1222_U292, P1_U3066, P1_U3979);
  not ginst4930 (P1_R1222_U293, P1_R1222_U154);
  or ginst4931 (P1_R1222_U294, P1_U3058, P1_U3977);
  nand ginst4932 (P1_R1222_U295, P1_R1222_U172, P1_R1222_U175);
  not ginst4933 (P1_R1222_U296, P1_R1222_U87);
  or ginst4934 (P1_R1222_U297, P1_U3065, P1_U3978);
  nand ginst4935 (P1_R1222_U298, P1_R1222_U154, P1_R1222_U167, P1_R1222_U297);
  not ginst4936 (P1_R1222_U299, P1_R1222_U152);
  not ginst4937 (P1_R1222_U30, P1_U3450);
  or ginst4938 (P1_R1222_U300, P1_U3053, P1_U3975);
  nand ginst4939 (P1_R1222_U301, P1_U3053, P1_U3975);
  not ginst4940 (P1_R1222_U302, P1_R1222_U150);
  nand ginst4941 (P1_R1222_U303, P1_R1222_U150, P1_U3974);
  not ginst4942 (P1_R1222_U304, P1_R1222_U148);
  nand ginst4943 (P1_R1222_U305, P1_R1222_U154, P1_R1222_U297);
  not ginst4944 (P1_R1222_U306, P1_R1222_U90);
  or ginst4945 (P1_R1222_U307, P1_U3058, P1_U3977);
  nand ginst4946 (P1_R1222_U308, P1_R1222_U307, P1_R1222_U90);
  nand ginst4947 (P1_R1222_U309, P1_R1222_U153, P1_R1222_U172, P1_R1222_U308);
  not ginst4948 (P1_R1222_U31, P1_U3077);
  nand ginst4949 (P1_R1222_U310, P1_R1222_U172, P1_R1222_U306);
  nand ginst4950 (P1_R1222_U311, P1_U3057, P1_U3976);
  nand ginst4951 (P1_R1222_U312, P1_R1222_U167, P1_R1222_U310, P1_R1222_U311);
  or ginst4952 (P1_R1222_U313, P1_U3058, P1_U3977);
  nand ginst4953 (P1_R1222_U314, P1_R1222_U161, P1_R1222_U281);
  not ginst4954 (P1_R1222_U315, P1_R1222_U92);
  nand ginst4955 (P1_R1222_U316, P1_R1222_U10, P1_R1222_U92);
  nand ginst4956 (P1_R1222_U317, P1_R1222_U135, P1_R1222_U316);
  nand ginst4957 (P1_R1222_U318, P1_R1222_U277, P1_R1222_U316);
  nand ginst4958 (P1_R1222_U319, P1_R1222_U318, P1_R1222_U452);
  nand ginst4959 (P1_R1222_U32, P1_U3077, P1_U3450);
  or ginst4960 (P1_R1222_U320, P1_U3081, P1_U3508);
  nand ginst4961 (P1_R1222_U321, P1_R1222_U320, P1_R1222_U92);
  nand ginst4962 (P1_R1222_U322, P1_R1222_U136, P1_R1222_U321);
  nand ginst4963 (P1_R1222_U323, P1_R1222_U315, P1_R1222_U81);
  nand ginst4964 (P1_R1222_U324, P1_U3076, P1_U3982);
  nand ginst4965 (P1_R1222_U325, P1_R1222_U10, P1_R1222_U323, P1_R1222_U324);
  or ginst4966 (P1_R1222_U326, P1_U3078, P1_U3455);
  not ginst4967 (P1_R1222_U327, P1_R1222_U160);
  or ginst4968 (P1_R1222_U328, P1_U3081, P1_U3508);
  or ginst4969 (P1_R1222_U329, P1_U3073, P1_U3500);
  not ginst4970 (P1_R1222_U33, P1_U3461);
  nand ginst4971 (P1_R1222_U330, P1_R1222_U329, P1_R1222_U93);
  nand ginst4972 (P1_R1222_U331, P1_R1222_U137, P1_R1222_U330);
  nand ginst4973 (P1_R1222_U332, P1_R1222_U261, P1_R1222_U60);
  nand ginst4974 (P1_R1222_U333, P1_U3069, P1_U3503);
  nand ginst4975 (P1_R1222_U334, P1_R1222_U138, P1_R1222_U332);
  or ginst4976 (P1_R1222_U335, P1_U3073, P1_U3500);
  nand ginst4977 (P1_R1222_U336, P1_R1222_U166, P1_R1222_U249);
  not ginst4978 (P1_R1222_U337, P1_R1222_U94);
  or ginst4979 (P1_R1222_U338, P1_U3072, P1_U3488);
  nand ginst4980 (P1_R1222_U339, P1_R1222_U338, P1_R1222_U94);
  not ginst4981 (P1_R1222_U34, P1_U3064);
  nand ginst4982 (P1_R1222_U340, P1_R1222_U139, P1_R1222_U339);
  nand ginst4983 (P1_R1222_U341, P1_R1222_U171, P1_R1222_U337);
  nand ginst4984 (P1_R1222_U342, P1_U3080, P1_U3491);
  nand ginst4985 (P1_R1222_U343, P1_R1222_U140, P1_R1222_U341);
  or ginst4986 (P1_R1222_U344, P1_U3072, P1_U3488);
  or ginst4987 (P1_R1222_U345, P1_U3083, P1_U3479);
  nand ginst4988 (P1_R1222_U346, P1_R1222_U345, P1_R1222_U41);
  nand ginst4989 (P1_R1222_U347, P1_R1222_U141, P1_R1222_U346);
  nand ginst4990 (P1_R1222_U348, P1_R1222_U170, P1_R1222_U205);
  nand ginst4991 (P1_R1222_U349, P1_U3062, P1_U3482);
  nand ginst4992 (P1_R1222_U35, P1_U3060, P1_U3464);
  nand ginst4993 (P1_R1222_U350, P1_R1222_U142, P1_R1222_U348);
  nand ginst4994 (P1_R1222_U351, P1_R1222_U170, P1_R1222_U206);
  nand ginst4995 (P1_R1222_U352, P1_R1222_U203, P1_R1222_U62);
  nand ginst4996 (P1_R1222_U353, P1_R1222_U213, P1_R1222_U23);
  nand ginst4997 (P1_R1222_U354, P1_R1222_U227, P1_R1222_U35);
  nand ginst4998 (P1_R1222_U355, P1_R1222_U179, P1_R1222_U230);
  nand ginst4999 (P1_R1222_U356, P1_R1222_U172, P1_R1222_U313);
  nand ginst5000 (P1_R1222_U357, P1_R1222_U175, P1_R1222_U297);
  nand ginst5001 (P1_R1222_U358, P1_R1222_U328, P1_R1222_U81);
  nand ginst5002 (P1_R1222_U359, P1_R1222_U281, P1_R1222_U78);
  not ginst5003 (P1_R1222_U36, P1_U3467);
  nand ginst5004 (P1_R1222_U360, P1_R1222_U335, P1_R1222_U60);
  nand ginst5005 (P1_R1222_U361, P1_R1222_U171, P1_R1222_U344);
  nand ginst5006 (P1_R1222_U362, P1_R1222_U249, P1_R1222_U69);
  nand ginst5007 (P1_R1222_U363, P1_U3054, P1_U3974);
  nand ginst5008 (P1_R1222_U364, P1_R1222_U167, P1_R1222_U295);
  nand ginst5009 (P1_R1222_U365, P1_R1222_U294, P1_U3057);
  nand ginst5010 (P1_R1222_U366, P1_R1222_U294, P1_U3976);
  nand ginst5011 (P1_R1222_U367, P1_R1222_U167, P1_R1222_U295, P1_R1222_U300);
  nand ginst5012 (P1_R1222_U368, P1_R1222_U133, P1_R1222_U154, P1_R1222_U167);
  nand ginst5013 (P1_R1222_U369, P1_R1222_U296, P1_R1222_U300);
  not ginst5014 (P1_R1222_U37, P1_U3476);
  nand ginst5015 (P1_R1222_U370, P1_R1222_U40, P1_U3083);
  nand ginst5016 (P1_R1222_U371, P1_R1222_U39, P1_U3479);
  nand ginst5017 (P1_R1222_U372, P1_R1222_U370, P1_R1222_U371);
  nand ginst5018 (P1_R1222_U373, P1_R1222_U351, P1_R1222_U41);
  nand ginst5019 (P1_R1222_U374, P1_R1222_U205, P1_R1222_U372);
  nand ginst5020 (P1_R1222_U375, P1_R1222_U37, P1_U3084);
  nand ginst5021 (P1_R1222_U376, P1_R1222_U38, P1_U3476);
  nand ginst5022 (P1_R1222_U377, P1_R1222_U375, P1_R1222_U376);
  nand ginst5023 (P1_R1222_U378, P1_R1222_U143, P1_R1222_U352);
  nand ginst5024 (P1_R1222_U379, P1_R1222_U202, P1_R1222_U377);
  not ginst5025 (P1_R1222_U38, P1_U3084);
  nand ginst5026 (P1_R1222_U380, P1_R1222_U24, P1_U3070);
  nand ginst5027 (P1_R1222_U381, P1_R1222_U22, P1_U3473);
  nand ginst5028 (P1_R1222_U382, P1_R1222_U20, P1_U3071);
  nand ginst5029 (P1_R1222_U383, P1_R1222_U21, P1_U3470);
  nand ginst5030 (P1_R1222_U384, P1_R1222_U382, P1_R1222_U383);
  nand ginst5031 (P1_R1222_U385, P1_R1222_U353, P1_R1222_U42);
  nand ginst5032 (P1_R1222_U386, P1_R1222_U194, P1_R1222_U384);
  nand ginst5033 (P1_R1222_U387, P1_R1222_U36, P1_U3067);
  nand ginst5034 (P1_R1222_U388, P1_R1222_U27, P1_U3467);
  nand ginst5035 (P1_R1222_U389, P1_R1222_U25, P1_U3060);
  not ginst5036 (P1_R1222_U39, P1_U3083);
  nand ginst5037 (P1_R1222_U390, P1_R1222_U26, P1_U3464);
  nand ginst5038 (P1_R1222_U391, P1_R1222_U389, P1_R1222_U390);
  nand ginst5039 (P1_R1222_U392, P1_R1222_U354, P1_R1222_U45);
  nand ginst5040 (P1_R1222_U393, P1_R1222_U220, P1_R1222_U391);
  nand ginst5041 (P1_R1222_U394, P1_R1222_U33, P1_U3064);
  nand ginst5042 (P1_R1222_U395, P1_R1222_U34, P1_U3461);
  nand ginst5043 (P1_R1222_U396, P1_R1222_U394, P1_R1222_U395);
  nand ginst5044 (P1_R1222_U397, P1_R1222_U144, P1_R1222_U355);
  nand ginst5045 (P1_R1222_U398, P1_R1222_U229, P1_R1222_U396);
  nand ginst5046 (P1_R1222_U399, P1_R1222_U28, P1_U3068);
  and ginst5047 (P1_R1222_U4, P1_R1222_U177, P1_R1222_U178);
  not ginst5048 (P1_R1222_U40, P1_U3479);
  nand ginst5049 (P1_R1222_U400, P1_R1222_U29, P1_U3458);
  nand ginst5050 (P1_R1222_U401, P1_R1222_U146, P1_U3055);
  nand ginst5051 (P1_R1222_U402, P1_R1222_U145, P1_U3985);
  nand ginst5052 (P1_R1222_U403, P1_R1222_U146, P1_U3055);
  nand ginst5053 (P1_R1222_U404, P1_R1222_U145, P1_U3985);
  nand ginst5054 (P1_R1222_U405, P1_R1222_U403, P1_R1222_U404);
  nand ginst5055 (P1_R1222_U406, P1_R1222_U147, P1_R1222_U148);
  nand ginst5056 (P1_R1222_U407, P1_R1222_U304, P1_R1222_U405);
  nand ginst5057 (P1_R1222_U408, P1_R1222_U89, P1_U3054);
  nand ginst5058 (P1_R1222_U409, P1_R1222_U88, P1_U3974);
  nand ginst5059 (P1_R1222_U41, P1_R1222_U204, P1_R1222_U62);
  nand ginst5060 (P1_R1222_U410, P1_R1222_U89, P1_U3054);
  nand ginst5061 (P1_R1222_U411, P1_R1222_U88, P1_U3974);
  nand ginst5062 (P1_R1222_U412, P1_R1222_U410, P1_R1222_U411);
  nand ginst5063 (P1_R1222_U413, P1_R1222_U149, P1_R1222_U150);
  nand ginst5064 (P1_R1222_U414, P1_R1222_U302, P1_R1222_U412);
  nand ginst5065 (P1_R1222_U415, P1_R1222_U47, P1_U3053);
  nand ginst5066 (P1_R1222_U416, P1_R1222_U48, P1_U3975);
  nand ginst5067 (P1_R1222_U417, P1_R1222_U47, P1_U3053);
  nand ginst5068 (P1_R1222_U418, P1_R1222_U48, P1_U3975);
  nand ginst5069 (P1_R1222_U419, P1_R1222_U417, P1_R1222_U418);
  nand ginst5070 (P1_R1222_U42, P1_R1222_U118, P1_R1222_U192);
  nand ginst5071 (P1_R1222_U420, P1_R1222_U151, P1_R1222_U152);
  nand ginst5072 (P1_R1222_U421, P1_R1222_U299, P1_R1222_U419);
  nand ginst5073 (P1_R1222_U422, P1_R1222_U50, P1_U3057);
  nand ginst5074 (P1_R1222_U423, P1_R1222_U49, P1_U3976);
  nand ginst5075 (P1_R1222_U424, P1_R1222_U51, P1_U3058);
  nand ginst5076 (P1_R1222_U425, P1_R1222_U52, P1_U3977);
  nand ginst5077 (P1_R1222_U426, P1_R1222_U424, P1_R1222_U425);
  nand ginst5078 (P1_R1222_U427, P1_R1222_U356, P1_R1222_U90);
  nand ginst5079 (P1_R1222_U428, P1_R1222_U306, P1_R1222_U426);
  nand ginst5080 (P1_R1222_U429, P1_R1222_U53, P1_U3065);
  nand ginst5081 (P1_R1222_U43, P1_R1222_U181, P1_R1222_U182);
  nand ginst5082 (P1_R1222_U430, P1_R1222_U54, P1_U3978);
  nand ginst5083 (P1_R1222_U431, P1_R1222_U429, P1_R1222_U430);
  nand ginst5084 (P1_R1222_U432, P1_R1222_U154, P1_R1222_U357);
  nand ginst5085 (P1_R1222_U433, P1_R1222_U293, P1_R1222_U431);
  nand ginst5086 (P1_R1222_U434, P1_R1222_U85, P1_U3066);
  nand ginst5087 (P1_R1222_U435, P1_R1222_U86, P1_U3979);
  nand ginst5088 (P1_R1222_U436, P1_R1222_U85, P1_U3066);
  nand ginst5089 (P1_R1222_U437, P1_R1222_U86, P1_U3979);
  nand ginst5090 (P1_R1222_U438, P1_R1222_U436, P1_R1222_U437);
  nand ginst5091 (P1_R1222_U439, P1_R1222_U155, P1_R1222_U156);
  nand ginst5092 (P1_R1222_U44, P1_U3078, P1_U3455);
  nand ginst5093 (P1_R1222_U440, P1_R1222_U289, P1_R1222_U438);
  nand ginst5094 (P1_R1222_U441, P1_R1222_U83, P1_U3061);
  nand ginst5095 (P1_R1222_U442, P1_R1222_U84, P1_U3980);
  nand ginst5096 (P1_R1222_U443, P1_R1222_U83, P1_U3061);
  nand ginst5097 (P1_R1222_U444, P1_R1222_U84, P1_U3980);
  nand ginst5098 (P1_R1222_U445, P1_R1222_U443, P1_R1222_U444);
  nand ginst5099 (P1_R1222_U446, P1_R1222_U157, P1_R1222_U158);
  nand ginst5100 (P1_R1222_U447, P1_R1222_U285, P1_R1222_U445);
  nand ginst5101 (P1_R1222_U448, P1_R1222_U55, P1_U3075);
  nand ginst5102 (P1_R1222_U449, P1_R1222_U56, P1_U3981);
  nand ginst5103 (P1_R1222_U45, P1_R1222_U122, P1_R1222_U218);
  nand ginst5104 (P1_R1222_U450, P1_R1222_U55, P1_U3075);
  nand ginst5105 (P1_R1222_U451, P1_R1222_U56, P1_U3981);
  nand ginst5106 (P1_R1222_U452, P1_R1222_U450, P1_R1222_U451);
  nand ginst5107 (P1_R1222_U453, P1_R1222_U82, P1_U3076);
  nand ginst5108 (P1_R1222_U454, P1_R1222_U91, P1_U3982);
  nand ginst5109 (P1_R1222_U455, P1_R1222_U160, P1_R1222_U181);
  nand ginst5110 (P1_R1222_U456, P1_R1222_U32, P1_R1222_U327);
  nand ginst5111 (P1_R1222_U457, P1_R1222_U79, P1_U3081);
  nand ginst5112 (P1_R1222_U458, P1_R1222_U80, P1_U3508);
  nand ginst5113 (P1_R1222_U459, P1_R1222_U457, P1_R1222_U458);
  nand ginst5114 (P1_R1222_U46, P1_R1222_U214, P1_R1222_U215);
  nand ginst5115 (P1_R1222_U460, P1_R1222_U358, P1_R1222_U92);
  nand ginst5116 (P1_R1222_U461, P1_R1222_U315, P1_R1222_U459);
  nand ginst5117 (P1_R1222_U462, P1_R1222_U76, P1_U3082);
  nand ginst5118 (P1_R1222_U463, P1_R1222_U77, P1_U3506);
  nand ginst5119 (P1_R1222_U464, P1_R1222_U462, P1_R1222_U463);
  nand ginst5120 (P1_R1222_U465, P1_R1222_U161, P1_R1222_U359);
  nand ginst5121 (P1_R1222_U466, P1_R1222_U269, P1_R1222_U464);
  nand ginst5122 (P1_R1222_U467, P1_R1222_U61, P1_U3069);
  nand ginst5123 (P1_R1222_U468, P1_R1222_U59, P1_U3503);
  nand ginst5124 (P1_R1222_U469, P1_R1222_U57, P1_U3073);
  not ginst5125 (P1_R1222_U47, P1_U3975);
  nand ginst5126 (P1_R1222_U470, P1_R1222_U58, P1_U3500);
  nand ginst5127 (P1_R1222_U471, P1_R1222_U469, P1_R1222_U470);
  nand ginst5128 (P1_R1222_U472, P1_R1222_U360, P1_R1222_U93);
  nand ginst5129 (P1_R1222_U473, P1_R1222_U261, P1_R1222_U471);
  nand ginst5130 (P1_R1222_U474, P1_R1222_U74, P1_U3074);
  nand ginst5131 (P1_R1222_U475, P1_R1222_U75, P1_U3497);
  nand ginst5132 (P1_R1222_U476, P1_R1222_U74, P1_U3074);
  nand ginst5133 (P1_R1222_U477, P1_R1222_U75, P1_U3497);
  nand ginst5134 (P1_R1222_U478, P1_R1222_U476, P1_R1222_U477);
  nand ginst5135 (P1_R1222_U479, P1_R1222_U162, P1_R1222_U163);
  not ginst5136 (P1_R1222_U48, P1_U3053);
  nand ginst5137 (P1_R1222_U480, P1_R1222_U257, P1_R1222_U478);
  nand ginst5138 (P1_R1222_U481, P1_R1222_U72, P1_U3079);
  nand ginst5139 (P1_R1222_U482, P1_R1222_U73, P1_U3494);
  nand ginst5140 (P1_R1222_U483, P1_R1222_U72, P1_U3079);
  nand ginst5141 (P1_R1222_U484, P1_R1222_U73, P1_U3494);
  nand ginst5142 (P1_R1222_U485, P1_R1222_U483, P1_R1222_U484);
  nand ginst5143 (P1_R1222_U486, P1_R1222_U164, P1_R1222_U165);
  nand ginst5144 (P1_R1222_U487, P1_R1222_U253, P1_R1222_U485);
  nand ginst5145 (P1_R1222_U488, P1_R1222_U70, P1_U3080);
  nand ginst5146 (P1_R1222_U489, P1_R1222_U71, P1_U3491);
  not ginst5147 (P1_R1222_U49, P1_U3057);
  nand ginst5148 (P1_R1222_U490, P1_R1222_U65, P1_U3072);
  nand ginst5149 (P1_R1222_U491, P1_R1222_U66, P1_U3488);
  nand ginst5150 (P1_R1222_U492, P1_R1222_U490, P1_R1222_U491);
  nand ginst5151 (P1_R1222_U493, P1_R1222_U361, P1_R1222_U94);
  nand ginst5152 (P1_R1222_U494, P1_R1222_U337, P1_R1222_U492);
  nand ginst5153 (P1_R1222_U495, P1_R1222_U67, P1_U3063);
  nand ginst5154 (P1_R1222_U496, P1_R1222_U68, P1_U3485);
  nand ginst5155 (P1_R1222_U497, P1_R1222_U495, P1_R1222_U496);
  nand ginst5156 (P1_R1222_U498, P1_R1222_U166, P1_R1222_U362);
  nand ginst5157 (P1_R1222_U499, P1_R1222_U243, P1_R1222_U497);
  and ginst5158 (P1_R1222_U5, P1_R1222_U179, P1_R1222_U180);
  not ginst5159 (P1_R1222_U50, P1_U3976);
  nand ginst5160 (P1_R1222_U500, P1_R1222_U63, P1_U3062);
  nand ginst5161 (P1_R1222_U501, P1_R1222_U64, P1_U3482);
  nand ginst5162 (P1_R1222_U502, P1_R1222_U30, P1_U3077);
  nand ginst5163 (P1_R1222_U503, P1_R1222_U31, P1_U3450);
  not ginst5164 (P1_R1222_U51, P1_U3977);
  not ginst5165 (P1_R1222_U52, P1_U3058);
  not ginst5166 (P1_R1222_U53, P1_U3978);
  not ginst5167 (P1_R1222_U54, P1_U3065);
  not ginst5168 (P1_R1222_U55, P1_U3981);
  not ginst5169 (P1_R1222_U56, P1_U3075);
  not ginst5170 (P1_R1222_U57, P1_U3500);
  not ginst5171 (P1_R1222_U58, P1_U3073);
  not ginst5172 (P1_R1222_U59, P1_U3069);
  and ginst5173 (P1_R1222_U6, P1_R1222_U195, P1_R1222_U196);
  nand ginst5174 (P1_R1222_U60, P1_U3073, P1_U3500);
  not ginst5175 (P1_R1222_U61, P1_U3503);
  nand ginst5176 (P1_R1222_U62, P1_U3084, P1_U3476);
  not ginst5177 (P1_R1222_U63, P1_U3482);
  not ginst5178 (P1_R1222_U64, P1_U3062);
  not ginst5179 (P1_R1222_U65, P1_U3488);
  not ginst5180 (P1_R1222_U66, P1_U3072);
  not ginst5181 (P1_R1222_U67, P1_U3485);
  not ginst5182 (P1_R1222_U68, P1_U3063);
  nand ginst5183 (P1_R1222_U69, P1_U3063, P1_U3485);
  and ginst5184 (P1_R1222_U7, P1_R1222_U235, P1_R1222_U236);
  not ginst5185 (P1_R1222_U70, P1_U3491);
  not ginst5186 (P1_R1222_U71, P1_U3080);
  not ginst5187 (P1_R1222_U72, P1_U3494);
  not ginst5188 (P1_R1222_U73, P1_U3079);
  not ginst5189 (P1_R1222_U74, P1_U3497);
  not ginst5190 (P1_R1222_U75, P1_U3074);
  not ginst5191 (P1_R1222_U76, P1_U3506);
  not ginst5192 (P1_R1222_U77, P1_U3082);
  nand ginst5193 (P1_R1222_U78, P1_U3082, P1_U3506);
  not ginst5194 (P1_R1222_U79, P1_U3508);
  and ginst5195 (P1_R1222_U8, P1_R1222_U244, P1_R1222_U245);
  not ginst5196 (P1_R1222_U80, P1_U3081);
  nand ginst5197 (P1_R1222_U81, P1_U3081, P1_U3508);
  not ginst5198 (P1_R1222_U82, P1_U3982);
  not ginst5199 (P1_R1222_U83, P1_U3980);
  not ginst5200 (P1_R1222_U84, P1_U3061);
  not ginst5201 (P1_R1222_U85, P1_U3979);
  not ginst5202 (P1_R1222_U86, P1_U3066);
  nand ginst5203 (P1_R1222_U87, P1_U3057, P1_U3976);
  not ginst5204 (P1_R1222_U88, P1_U3054);
  not ginst5205 (P1_R1222_U89, P1_U3974);
  and ginst5206 (P1_R1222_U9, P1_R1222_U262, P1_R1222_U263);
  nand ginst5207 (P1_R1222_U90, P1_R1222_U175, P1_R1222_U305);
  not ginst5208 (P1_R1222_U91, P1_U3076);
  nand ginst5209 (P1_R1222_U92, P1_R1222_U314, P1_R1222_U78);
  nand ginst5210 (P1_R1222_U93, P1_R1222_U259, P1_R1222_U260);
  nand ginst5211 (P1_R1222_U94, P1_R1222_U336, P1_R1222_U69);
  nand ginst5212 (P1_R1222_U95, P1_R1222_U455, P1_R1222_U456);
  nand ginst5213 (P1_R1222_U96, P1_R1222_U502, P1_R1222_U503);
  nand ginst5214 (P1_R1222_U97, P1_R1222_U373, P1_R1222_U374);
  nand ginst5215 (P1_R1222_U98, P1_R1222_U378, P1_R1222_U379);
  nand ginst5216 (P1_R1222_U99, P1_R1222_U385, P1_R1222_U386);
  and ginst5217 (P1_R1240_U10, P1_R1240_U270, P1_R1240_U271);
  nand ginst5218 (P1_R1240_U100, P1_R1240_U392, P1_R1240_U393);
  nand ginst5219 (P1_R1240_U101, P1_R1240_U397, P1_R1240_U398);
  nand ginst5220 (P1_R1240_U102, P1_R1240_U406, P1_R1240_U407);
  nand ginst5221 (P1_R1240_U103, P1_R1240_U413, P1_R1240_U414);
  nand ginst5222 (P1_R1240_U104, P1_R1240_U420, P1_R1240_U421);
  nand ginst5223 (P1_R1240_U105, P1_R1240_U427, P1_R1240_U428);
  nand ginst5224 (P1_R1240_U106, P1_R1240_U432, P1_R1240_U433);
  nand ginst5225 (P1_R1240_U107, P1_R1240_U439, P1_R1240_U440);
  nand ginst5226 (P1_R1240_U108, P1_R1240_U446, P1_R1240_U447);
  nand ginst5227 (P1_R1240_U109, P1_R1240_U460, P1_R1240_U461);
  and ginst5228 (P1_R1240_U11, P1_R1240_U347, P1_R1240_U350);
  nand ginst5229 (P1_R1240_U110, P1_R1240_U465, P1_R1240_U466);
  nand ginst5230 (P1_R1240_U111, P1_R1240_U472, P1_R1240_U473);
  nand ginst5231 (P1_R1240_U112, P1_R1240_U479, P1_R1240_U480);
  nand ginst5232 (P1_R1240_U113, P1_R1240_U486, P1_R1240_U487);
  nand ginst5233 (P1_R1240_U114, P1_R1240_U493, P1_R1240_U494);
  nand ginst5234 (P1_R1240_U115, P1_R1240_U498, P1_R1240_U499);
  and ginst5235 (P1_R1240_U116, P1_U3068, P1_U3458);
  and ginst5236 (P1_R1240_U117, P1_R1240_U186, P1_R1240_U188);
  and ginst5237 (P1_R1240_U118, P1_R1240_U191, P1_R1240_U193);
  and ginst5238 (P1_R1240_U119, P1_R1240_U199, P1_R1240_U200);
  and ginst5239 (P1_R1240_U12, P1_R1240_U340, P1_R1240_U343);
  and ginst5240 (P1_R1240_U120, P1_R1240_U23, P1_R1240_U380, P1_R1240_U381);
  and ginst5241 (P1_R1240_U121, P1_R1240_U211, P1_R1240_U6);
  and ginst5242 (P1_R1240_U122, P1_R1240_U217, P1_R1240_U219);
  and ginst5243 (P1_R1240_U123, P1_R1240_U35, P1_R1240_U387, P1_R1240_U388);
  and ginst5244 (P1_R1240_U124, P1_R1240_U225, P1_R1240_U4);
  and ginst5245 (P1_R1240_U125, P1_R1240_U180, P1_R1240_U233);
  and ginst5246 (P1_R1240_U126, P1_R1240_U203, P1_R1240_U7);
  and ginst5247 (P1_R1240_U127, P1_R1240_U170, P1_R1240_U238);
  and ginst5248 (P1_R1240_U128, P1_R1240_U249, P1_R1240_U8);
  and ginst5249 (P1_R1240_U129, P1_R1240_U171, P1_R1240_U247);
  and ginst5250 (P1_R1240_U13, P1_R1240_U331, P1_R1240_U334);
  and ginst5251 (P1_R1240_U130, P1_R1240_U266, P1_R1240_U267);
  and ginst5252 (P1_R1240_U131, P1_R1240_U10, P1_R1240_U281);
  and ginst5253 (P1_R1240_U132, P1_R1240_U279, P1_R1240_U284);
  and ginst5254 (P1_R1240_U133, P1_R1240_U297, P1_R1240_U300);
  and ginst5255 (P1_R1240_U134, P1_R1240_U301, P1_R1240_U367);
  and ginst5256 (P1_R1240_U135, P1_R1240_U159, P1_R1240_U277);
  and ginst5257 (P1_R1240_U136, P1_R1240_U453, P1_R1240_U454, P1_R1240_U81);
  and ginst5258 (P1_R1240_U137, P1_R1240_U467, P1_R1240_U468, P1_R1240_U60);
  and ginst5259 (P1_R1240_U138, P1_R1240_U333, P1_R1240_U9);
  and ginst5260 (P1_R1240_U139, P1_R1240_U171, P1_R1240_U488, P1_R1240_U489);
  and ginst5261 (P1_R1240_U14, P1_R1240_U322, P1_R1240_U325);
  and ginst5262 (P1_R1240_U140, P1_R1240_U342, P1_R1240_U8);
  and ginst5263 (P1_R1240_U141, P1_R1240_U170, P1_R1240_U500, P1_R1240_U501);
  and ginst5264 (P1_R1240_U142, P1_R1240_U349, P1_R1240_U7);
  nand ginst5265 (P1_R1240_U143, P1_R1240_U119, P1_R1240_U201);
  nand ginst5266 (P1_R1240_U144, P1_R1240_U216, P1_R1240_U228);
  not ginst5267 (P1_R1240_U145, P1_U3055);
  not ginst5268 (P1_R1240_U146, P1_U3985);
  and ginst5269 (P1_R1240_U147, P1_R1240_U401, P1_R1240_U402);
  nand ginst5270 (P1_R1240_U148, P1_R1240_U168, P1_R1240_U303, P1_R1240_U363);
  and ginst5271 (P1_R1240_U149, P1_R1240_U408, P1_R1240_U409);
  and ginst5272 (P1_R1240_U15, P1_R1240_U317, P1_R1240_U319);
  nand ginst5273 (P1_R1240_U150, P1_R1240_U134, P1_R1240_U368, P1_R1240_U369);
  and ginst5274 (P1_R1240_U151, P1_R1240_U415, P1_R1240_U416);
  nand ginst5275 (P1_R1240_U152, P1_R1240_U298, P1_R1240_U364, P1_R1240_U87);
  and ginst5276 (P1_R1240_U153, P1_R1240_U422, P1_R1240_U423);
  nand ginst5277 (P1_R1240_U154, P1_R1240_U291, P1_R1240_U292);
  and ginst5278 (P1_R1240_U155, P1_R1240_U434, P1_R1240_U435);
  nand ginst5279 (P1_R1240_U156, P1_R1240_U287, P1_R1240_U288);
  and ginst5280 (P1_R1240_U157, P1_R1240_U441, P1_R1240_U442);
  nand ginst5281 (P1_R1240_U158, P1_R1240_U132, P1_R1240_U283);
  and ginst5282 (P1_R1240_U159, P1_R1240_U448, P1_R1240_U449);
  and ginst5283 (P1_R1240_U16, P1_R1240_U309, P1_R1240_U312);
  nand ginst5284 (P1_R1240_U160, P1_R1240_U326, P1_R1240_U44);
  nand ginst5285 (P1_R1240_U161, P1_R1240_U130, P1_R1240_U268);
  and ginst5286 (P1_R1240_U162, P1_R1240_U474, P1_R1240_U475);
  nand ginst5287 (P1_R1240_U163, P1_R1240_U255, P1_R1240_U256);
  and ginst5288 (P1_R1240_U164, P1_R1240_U481, P1_R1240_U482);
  nand ginst5289 (P1_R1240_U165, P1_R1240_U251, P1_R1240_U252);
  nand ginst5290 (P1_R1240_U166, P1_R1240_U241, P1_R1240_U242);
  nand ginst5291 (P1_R1240_U167, P1_R1240_U365, P1_R1240_U366);
  nand ginst5292 (P1_R1240_U168, P1_R1240_U150, P1_U3054);
  not ginst5293 (P1_R1240_U169, P1_R1240_U35);
  and ginst5294 (P1_R1240_U17, P1_R1240_U231, P1_R1240_U234);
  nand ginst5295 (P1_R1240_U170, P1_U3083, P1_U3479);
  nand ginst5296 (P1_R1240_U171, P1_U3072, P1_U3488);
  nand ginst5297 (P1_R1240_U172, P1_U3058, P1_U3977);
  not ginst5298 (P1_R1240_U173, P1_R1240_U69);
  not ginst5299 (P1_R1240_U174, P1_R1240_U78);
  nand ginst5300 (P1_R1240_U175, P1_U3065, P1_U3978);
  not ginst5301 (P1_R1240_U176, P1_R1240_U62);
  or ginst5302 (P1_R1240_U177, P1_U3067, P1_U3467);
  or ginst5303 (P1_R1240_U178, P1_U3060, P1_U3464);
  or ginst5304 (P1_R1240_U179, P1_U3064, P1_U3461);
  and ginst5305 (P1_R1240_U18, P1_R1240_U223, P1_R1240_U226);
  or ginst5306 (P1_R1240_U180, P1_U3068, P1_U3458);
  not ginst5307 (P1_R1240_U181, P1_R1240_U32);
  or ginst5308 (P1_R1240_U182, P1_U3078, P1_U3455);
  not ginst5309 (P1_R1240_U183, P1_R1240_U43);
  not ginst5310 (P1_R1240_U184, P1_R1240_U44);
  nand ginst5311 (P1_R1240_U185, P1_R1240_U43, P1_R1240_U44);
  nand ginst5312 (P1_R1240_U186, P1_R1240_U116, P1_R1240_U179);
  nand ginst5313 (P1_R1240_U187, P1_R1240_U185, P1_R1240_U5);
  nand ginst5314 (P1_R1240_U188, P1_U3064, P1_U3461);
  nand ginst5315 (P1_R1240_U189, P1_R1240_U117, P1_R1240_U187);
  and ginst5316 (P1_R1240_U19, P1_R1240_U209, P1_R1240_U212);
  nand ginst5317 (P1_R1240_U190, P1_R1240_U35, P1_R1240_U36);
  nand ginst5318 (P1_R1240_U191, P1_R1240_U190, P1_U3067);
  nand ginst5319 (P1_R1240_U192, P1_R1240_U189, P1_R1240_U4);
  nand ginst5320 (P1_R1240_U193, P1_R1240_U169, P1_U3467);
  not ginst5321 (P1_R1240_U194, P1_R1240_U42);
  or ginst5322 (P1_R1240_U195, P1_U3070, P1_U3473);
  or ginst5323 (P1_R1240_U196, P1_U3071, P1_U3470);
  not ginst5324 (P1_R1240_U197, P1_R1240_U23);
  nand ginst5325 (P1_R1240_U198, P1_R1240_U23, P1_R1240_U24);
  nand ginst5326 (P1_R1240_U199, P1_R1240_U198, P1_U3070);
  not ginst5327 (P1_R1240_U20, P1_U3470);
  nand ginst5328 (P1_R1240_U200, P1_R1240_U197, P1_U3473);
  nand ginst5329 (P1_R1240_U201, P1_R1240_U42, P1_R1240_U6);
  not ginst5330 (P1_R1240_U202, P1_R1240_U143);
  or ginst5331 (P1_R1240_U203, P1_U3084, P1_U3476);
  nand ginst5332 (P1_R1240_U204, P1_R1240_U143, P1_R1240_U203);
  not ginst5333 (P1_R1240_U205, P1_R1240_U41);
  or ginst5334 (P1_R1240_U206, P1_U3083, P1_U3479);
  or ginst5335 (P1_R1240_U207, P1_U3071, P1_U3470);
  nand ginst5336 (P1_R1240_U208, P1_R1240_U207, P1_R1240_U42);
  nand ginst5337 (P1_R1240_U209, P1_R1240_U120, P1_R1240_U208);
  not ginst5338 (P1_R1240_U21, P1_U3071);
  nand ginst5339 (P1_R1240_U210, P1_R1240_U194, P1_R1240_U23);
  nand ginst5340 (P1_R1240_U211, P1_U3070, P1_U3473);
  nand ginst5341 (P1_R1240_U212, P1_R1240_U121, P1_R1240_U210);
  or ginst5342 (P1_R1240_U213, P1_U3071, P1_U3470);
  nand ginst5343 (P1_R1240_U214, P1_R1240_U180, P1_R1240_U184);
  nand ginst5344 (P1_R1240_U215, P1_U3068, P1_U3458);
  not ginst5345 (P1_R1240_U216, P1_R1240_U46);
  nand ginst5346 (P1_R1240_U217, P1_R1240_U183, P1_R1240_U5);
  nand ginst5347 (P1_R1240_U218, P1_R1240_U179, P1_R1240_U46);
  nand ginst5348 (P1_R1240_U219, P1_U3064, P1_U3461);
  not ginst5349 (P1_R1240_U22, P1_U3070);
  not ginst5350 (P1_R1240_U220, P1_R1240_U45);
  or ginst5351 (P1_R1240_U221, P1_U3060, P1_U3464);
  nand ginst5352 (P1_R1240_U222, P1_R1240_U221, P1_R1240_U45);
  nand ginst5353 (P1_R1240_U223, P1_R1240_U123, P1_R1240_U222);
  nand ginst5354 (P1_R1240_U224, P1_R1240_U220, P1_R1240_U35);
  nand ginst5355 (P1_R1240_U225, P1_U3067, P1_U3467);
  nand ginst5356 (P1_R1240_U226, P1_R1240_U124, P1_R1240_U224);
  or ginst5357 (P1_R1240_U227, P1_U3060, P1_U3464);
  nand ginst5358 (P1_R1240_U228, P1_R1240_U180, P1_R1240_U183);
  not ginst5359 (P1_R1240_U229, P1_R1240_U144);
  nand ginst5360 (P1_R1240_U23, P1_U3071, P1_U3470);
  nand ginst5361 (P1_R1240_U230, P1_U3064, P1_U3461);
  nand ginst5362 (P1_R1240_U231, P1_R1240_U399, P1_R1240_U400, P1_R1240_U43, P1_R1240_U44);
  nand ginst5363 (P1_R1240_U232, P1_R1240_U43, P1_R1240_U44);
  nand ginst5364 (P1_R1240_U233, P1_U3068, P1_U3458);
  nand ginst5365 (P1_R1240_U234, P1_R1240_U125, P1_R1240_U232);
  or ginst5366 (P1_R1240_U235, P1_U3083, P1_U3479);
  or ginst5367 (P1_R1240_U236, P1_U3062, P1_U3482);
  nand ginst5368 (P1_R1240_U237, P1_R1240_U176, P1_R1240_U7);
  nand ginst5369 (P1_R1240_U238, P1_U3062, P1_U3482);
  nand ginst5370 (P1_R1240_U239, P1_R1240_U127, P1_R1240_U237);
  not ginst5371 (P1_R1240_U24, P1_U3473);
  or ginst5372 (P1_R1240_U240, P1_U3062, P1_U3482);
  nand ginst5373 (P1_R1240_U241, P1_R1240_U126, P1_R1240_U143);
  nand ginst5374 (P1_R1240_U242, P1_R1240_U239, P1_R1240_U240);
  not ginst5375 (P1_R1240_U243, P1_R1240_U166);
  or ginst5376 (P1_R1240_U244, P1_U3080, P1_U3491);
  or ginst5377 (P1_R1240_U245, P1_U3072, P1_U3488);
  nand ginst5378 (P1_R1240_U246, P1_R1240_U173, P1_R1240_U8);
  nand ginst5379 (P1_R1240_U247, P1_U3080, P1_U3491);
  nand ginst5380 (P1_R1240_U248, P1_R1240_U129, P1_R1240_U246);
  or ginst5381 (P1_R1240_U249, P1_U3063, P1_U3485);
  not ginst5382 (P1_R1240_U25, P1_U3464);
  or ginst5383 (P1_R1240_U250, P1_U3080, P1_U3491);
  nand ginst5384 (P1_R1240_U251, P1_R1240_U128, P1_R1240_U166);
  nand ginst5385 (P1_R1240_U252, P1_R1240_U248, P1_R1240_U250);
  not ginst5386 (P1_R1240_U253, P1_R1240_U165);
  or ginst5387 (P1_R1240_U254, P1_U3079, P1_U3494);
  nand ginst5388 (P1_R1240_U255, P1_R1240_U165, P1_R1240_U254);
  nand ginst5389 (P1_R1240_U256, P1_U3079, P1_U3494);
  not ginst5390 (P1_R1240_U257, P1_R1240_U163);
  or ginst5391 (P1_R1240_U258, P1_U3074, P1_U3497);
  nand ginst5392 (P1_R1240_U259, P1_R1240_U163, P1_R1240_U258);
  not ginst5393 (P1_R1240_U26, P1_U3060);
  nand ginst5394 (P1_R1240_U260, P1_U3074, P1_U3497);
  not ginst5395 (P1_R1240_U261, P1_R1240_U93);
  or ginst5396 (P1_R1240_U262, P1_U3069, P1_U3503);
  or ginst5397 (P1_R1240_U263, P1_U3073, P1_U3500);
  not ginst5398 (P1_R1240_U264, P1_R1240_U60);
  nand ginst5399 (P1_R1240_U265, P1_R1240_U60, P1_R1240_U61);
  nand ginst5400 (P1_R1240_U266, P1_R1240_U265, P1_U3069);
  nand ginst5401 (P1_R1240_U267, P1_R1240_U264, P1_U3503);
  nand ginst5402 (P1_R1240_U268, P1_R1240_U9, P1_R1240_U93);
  not ginst5403 (P1_R1240_U269, P1_R1240_U161);
  not ginst5404 (P1_R1240_U27, P1_U3067);
  or ginst5405 (P1_R1240_U270, P1_U3076, P1_U3982);
  or ginst5406 (P1_R1240_U271, P1_U3081, P1_U3508);
  or ginst5407 (P1_R1240_U272, P1_U3075, P1_U3981);
  not ginst5408 (P1_R1240_U273, P1_R1240_U81);
  nand ginst5409 (P1_R1240_U274, P1_R1240_U273, P1_U3982);
  nand ginst5410 (P1_R1240_U275, P1_R1240_U274, P1_R1240_U91);
  nand ginst5411 (P1_R1240_U276, P1_R1240_U81, P1_R1240_U82);
  nand ginst5412 (P1_R1240_U277, P1_R1240_U275, P1_R1240_U276);
  nand ginst5413 (P1_R1240_U278, P1_R1240_U10, P1_R1240_U174);
  nand ginst5414 (P1_R1240_U279, P1_U3075, P1_U3981);
  not ginst5415 (P1_R1240_U28, P1_U3458);
  nand ginst5416 (P1_R1240_U280, P1_R1240_U277, P1_R1240_U278);
  or ginst5417 (P1_R1240_U281, P1_U3082, P1_U3506);
  or ginst5418 (P1_R1240_U282, P1_U3075, P1_U3981);
  nand ginst5419 (P1_R1240_U283, P1_R1240_U131, P1_R1240_U161, P1_R1240_U272);
  nand ginst5420 (P1_R1240_U284, P1_R1240_U280, P1_R1240_U282);
  not ginst5421 (P1_R1240_U285, P1_R1240_U158);
  or ginst5422 (P1_R1240_U286, P1_U3061, P1_U3980);
  nand ginst5423 (P1_R1240_U287, P1_R1240_U158, P1_R1240_U286);
  nand ginst5424 (P1_R1240_U288, P1_U3061, P1_U3980);
  not ginst5425 (P1_R1240_U289, P1_R1240_U156);
  not ginst5426 (P1_R1240_U29, P1_U3068);
  or ginst5427 (P1_R1240_U290, P1_U3066, P1_U3979);
  nand ginst5428 (P1_R1240_U291, P1_R1240_U156, P1_R1240_U290);
  nand ginst5429 (P1_R1240_U292, P1_U3066, P1_U3979);
  not ginst5430 (P1_R1240_U293, P1_R1240_U154);
  or ginst5431 (P1_R1240_U294, P1_U3058, P1_U3977);
  nand ginst5432 (P1_R1240_U295, P1_R1240_U172, P1_R1240_U175);
  not ginst5433 (P1_R1240_U296, P1_R1240_U87);
  or ginst5434 (P1_R1240_U297, P1_U3065, P1_U3978);
  nand ginst5435 (P1_R1240_U298, P1_R1240_U154, P1_R1240_U167, P1_R1240_U297);
  not ginst5436 (P1_R1240_U299, P1_R1240_U152);
  not ginst5437 (P1_R1240_U30, P1_U3450);
  or ginst5438 (P1_R1240_U300, P1_U3053, P1_U3975);
  nand ginst5439 (P1_R1240_U301, P1_U3053, P1_U3975);
  not ginst5440 (P1_R1240_U302, P1_R1240_U150);
  nand ginst5441 (P1_R1240_U303, P1_R1240_U150, P1_U3974);
  not ginst5442 (P1_R1240_U304, P1_R1240_U148);
  nand ginst5443 (P1_R1240_U305, P1_R1240_U154, P1_R1240_U297);
  not ginst5444 (P1_R1240_U306, P1_R1240_U90);
  or ginst5445 (P1_R1240_U307, P1_U3058, P1_U3977);
  nand ginst5446 (P1_R1240_U308, P1_R1240_U307, P1_R1240_U90);
  nand ginst5447 (P1_R1240_U309, P1_R1240_U153, P1_R1240_U172, P1_R1240_U308);
  not ginst5448 (P1_R1240_U31, P1_U3077);
  nand ginst5449 (P1_R1240_U310, P1_R1240_U172, P1_R1240_U306);
  nand ginst5450 (P1_R1240_U311, P1_U3057, P1_U3976);
  nand ginst5451 (P1_R1240_U312, P1_R1240_U167, P1_R1240_U310, P1_R1240_U311);
  or ginst5452 (P1_R1240_U313, P1_U3058, P1_U3977);
  nand ginst5453 (P1_R1240_U314, P1_R1240_U161, P1_R1240_U281);
  not ginst5454 (P1_R1240_U315, P1_R1240_U92);
  nand ginst5455 (P1_R1240_U316, P1_R1240_U10, P1_R1240_U92);
  nand ginst5456 (P1_R1240_U317, P1_R1240_U135, P1_R1240_U316);
  nand ginst5457 (P1_R1240_U318, P1_R1240_U277, P1_R1240_U316);
  nand ginst5458 (P1_R1240_U319, P1_R1240_U318, P1_R1240_U452);
  nand ginst5459 (P1_R1240_U32, P1_U3077, P1_U3450);
  or ginst5460 (P1_R1240_U320, P1_U3081, P1_U3508);
  nand ginst5461 (P1_R1240_U321, P1_R1240_U320, P1_R1240_U92);
  nand ginst5462 (P1_R1240_U322, P1_R1240_U136, P1_R1240_U321);
  nand ginst5463 (P1_R1240_U323, P1_R1240_U315, P1_R1240_U81);
  nand ginst5464 (P1_R1240_U324, P1_U3076, P1_U3982);
  nand ginst5465 (P1_R1240_U325, P1_R1240_U10, P1_R1240_U323, P1_R1240_U324);
  or ginst5466 (P1_R1240_U326, P1_U3078, P1_U3455);
  not ginst5467 (P1_R1240_U327, P1_R1240_U160);
  or ginst5468 (P1_R1240_U328, P1_U3081, P1_U3508);
  or ginst5469 (P1_R1240_U329, P1_U3073, P1_U3500);
  not ginst5470 (P1_R1240_U33, P1_U3461);
  nand ginst5471 (P1_R1240_U330, P1_R1240_U329, P1_R1240_U93);
  nand ginst5472 (P1_R1240_U331, P1_R1240_U137, P1_R1240_U330);
  nand ginst5473 (P1_R1240_U332, P1_R1240_U261, P1_R1240_U60);
  nand ginst5474 (P1_R1240_U333, P1_U3069, P1_U3503);
  nand ginst5475 (P1_R1240_U334, P1_R1240_U138, P1_R1240_U332);
  or ginst5476 (P1_R1240_U335, P1_U3073, P1_U3500);
  nand ginst5477 (P1_R1240_U336, P1_R1240_U166, P1_R1240_U249);
  not ginst5478 (P1_R1240_U337, P1_R1240_U94);
  or ginst5479 (P1_R1240_U338, P1_U3072, P1_U3488);
  nand ginst5480 (P1_R1240_U339, P1_R1240_U338, P1_R1240_U94);
  not ginst5481 (P1_R1240_U34, P1_U3064);
  nand ginst5482 (P1_R1240_U340, P1_R1240_U139, P1_R1240_U339);
  nand ginst5483 (P1_R1240_U341, P1_R1240_U171, P1_R1240_U337);
  nand ginst5484 (P1_R1240_U342, P1_U3080, P1_U3491);
  nand ginst5485 (P1_R1240_U343, P1_R1240_U140, P1_R1240_U341);
  or ginst5486 (P1_R1240_U344, P1_U3072, P1_U3488);
  or ginst5487 (P1_R1240_U345, P1_U3083, P1_U3479);
  nand ginst5488 (P1_R1240_U346, P1_R1240_U345, P1_R1240_U41);
  nand ginst5489 (P1_R1240_U347, P1_R1240_U141, P1_R1240_U346);
  nand ginst5490 (P1_R1240_U348, P1_R1240_U170, P1_R1240_U205);
  nand ginst5491 (P1_R1240_U349, P1_U3062, P1_U3482);
  nand ginst5492 (P1_R1240_U35, P1_U3060, P1_U3464);
  nand ginst5493 (P1_R1240_U350, P1_R1240_U142, P1_R1240_U348);
  nand ginst5494 (P1_R1240_U351, P1_R1240_U170, P1_R1240_U206);
  nand ginst5495 (P1_R1240_U352, P1_R1240_U203, P1_R1240_U62);
  nand ginst5496 (P1_R1240_U353, P1_R1240_U213, P1_R1240_U23);
  nand ginst5497 (P1_R1240_U354, P1_R1240_U227, P1_R1240_U35);
  nand ginst5498 (P1_R1240_U355, P1_R1240_U179, P1_R1240_U230);
  nand ginst5499 (P1_R1240_U356, P1_R1240_U172, P1_R1240_U313);
  nand ginst5500 (P1_R1240_U357, P1_R1240_U175, P1_R1240_U297);
  nand ginst5501 (P1_R1240_U358, P1_R1240_U328, P1_R1240_U81);
  nand ginst5502 (P1_R1240_U359, P1_R1240_U281, P1_R1240_U78);
  not ginst5503 (P1_R1240_U36, P1_U3467);
  nand ginst5504 (P1_R1240_U360, P1_R1240_U335, P1_R1240_U60);
  nand ginst5505 (P1_R1240_U361, P1_R1240_U171, P1_R1240_U344);
  nand ginst5506 (P1_R1240_U362, P1_R1240_U249, P1_R1240_U69);
  nand ginst5507 (P1_R1240_U363, P1_U3054, P1_U3974);
  nand ginst5508 (P1_R1240_U364, P1_R1240_U167, P1_R1240_U295);
  nand ginst5509 (P1_R1240_U365, P1_R1240_U294, P1_U3057);
  nand ginst5510 (P1_R1240_U366, P1_R1240_U294, P1_U3976);
  nand ginst5511 (P1_R1240_U367, P1_R1240_U167, P1_R1240_U295, P1_R1240_U300);
  nand ginst5512 (P1_R1240_U368, P1_R1240_U133, P1_R1240_U154, P1_R1240_U167);
  nand ginst5513 (P1_R1240_U369, P1_R1240_U296, P1_R1240_U300);
  not ginst5514 (P1_R1240_U37, P1_U3476);
  nand ginst5515 (P1_R1240_U370, P1_R1240_U40, P1_U3083);
  nand ginst5516 (P1_R1240_U371, P1_R1240_U39, P1_U3479);
  nand ginst5517 (P1_R1240_U372, P1_R1240_U370, P1_R1240_U371);
  nand ginst5518 (P1_R1240_U373, P1_R1240_U351, P1_R1240_U41);
  nand ginst5519 (P1_R1240_U374, P1_R1240_U205, P1_R1240_U372);
  nand ginst5520 (P1_R1240_U375, P1_R1240_U37, P1_U3084);
  nand ginst5521 (P1_R1240_U376, P1_R1240_U38, P1_U3476);
  nand ginst5522 (P1_R1240_U377, P1_R1240_U375, P1_R1240_U376);
  nand ginst5523 (P1_R1240_U378, P1_R1240_U143, P1_R1240_U352);
  nand ginst5524 (P1_R1240_U379, P1_R1240_U202, P1_R1240_U377);
  not ginst5525 (P1_R1240_U38, P1_U3084);
  nand ginst5526 (P1_R1240_U380, P1_R1240_U24, P1_U3070);
  nand ginst5527 (P1_R1240_U381, P1_R1240_U22, P1_U3473);
  nand ginst5528 (P1_R1240_U382, P1_R1240_U20, P1_U3071);
  nand ginst5529 (P1_R1240_U383, P1_R1240_U21, P1_U3470);
  nand ginst5530 (P1_R1240_U384, P1_R1240_U382, P1_R1240_U383);
  nand ginst5531 (P1_R1240_U385, P1_R1240_U353, P1_R1240_U42);
  nand ginst5532 (P1_R1240_U386, P1_R1240_U194, P1_R1240_U384);
  nand ginst5533 (P1_R1240_U387, P1_R1240_U36, P1_U3067);
  nand ginst5534 (P1_R1240_U388, P1_R1240_U27, P1_U3467);
  nand ginst5535 (P1_R1240_U389, P1_R1240_U25, P1_U3060);
  not ginst5536 (P1_R1240_U39, P1_U3083);
  nand ginst5537 (P1_R1240_U390, P1_R1240_U26, P1_U3464);
  nand ginst5538 (P1_R1240_U391, P1_R1240_U389, P1_R1240_U390);
  nand ginst5539 (P1_R1240_U392, P1_R1240_U354, P1_R1240_U45);
  nand ginst5540 (P1_R1240_U393, P1_R1240_U220, P1_R1240_U391);
  nand ginst5541 (P1_R1240_U394, P1_R1240_U33, P1_U3064);
  nand ginst5542 (P1_R1240_U395, P1_R1240_U34, P1_U3461);
  nand ginst5543 (P1_R1240_U396, P1_R1240_U394, P1_R1240_U395);
  nand ginst5544 (P1_R1240_U397, P1_R1240_U144, P1_R1240_U355);
  nand ginst5545 (P1_R1240_U398, P1_R1240_U229, P1_R1240_U396);
  nand ginst5546 (P1_R1240_U399, P1_R1240_U28, P1_U3068);
  and ginst5547 (P1_R1240_U4, P1_R1240_U177, P1_R1240_U178);
  not ginst5548 (P1_R1240_U40, P1_U3479);
  nand ginst5549 (P1_R1240_U400, P1_R1240_U29, P1_U3458);
  nand ginst5550 (P1_R1240_U401, P1_R1240_U146, P1_U3055);
  nand ginst5551 (P1_R1240_U402, P1_R1240_U145, P1_U3985);
  nand ginst5552 (P1_R1240_U403, P1_R1240_U146, P1_U3055);
  nand ginst5553 (P1_R1240_U404, P1_R1240_U145, P1_U3985);
  nand ginst5554 (P1_R1240_U405, P1_R1240_U403, P1_R1240_U404);
  nand ginst5555 (P1_R1240_U406, P1_R1240_U147, P1_R1240_U148);
  nand ginst5556 (P1_R1240_U407, P1_R1240_U304, P1_R1240_U405);
  nand ginst5557 (P1_R1240_U408, P1_R1240_U89, P1_U3054);
  nand ginst5558 (P1_R1240_U409, P1_R1240_U88, P1_U3974);
  nand ginst5559 (P1_R1240_U41, P1_R1240_U204, P1_R1240_U62);
  nand ginst5560 (P1_R1240_U410, P1_R1240_U89, P1_U3054);
  nand ginst5561 (P1_R1240_U411, P1_R1240_U88, P1_U3974);
  nand ginst5562 (P1_R1240_U412, P1_R1240_U410, P1_R1240_U411);
  nand ginst5563 (P1_R1240_U413, P1_R1240_U149, P1_R1240_U150);
  nand ginst5564 (P1_R1240_U414, P1_R1240_U302, P1_R1240_U412);
  nand ginst5565 (P1_R1240_U415, P1_R1240_U47, P1_U3053);
  nand ginst5566 (P1_R1240_U416, P1_R1240_U48, P1_U3975);
  nand ginst5567 (P1_R1240_U417, P1_R1240_U47, P1_U3053);
  nand ginst5568 (P1_R1240_U418, P1_R1240_U48, P1_U3975);
  nand ginst5569 (P1_R1240_U419, P1_R1240_U417, P1_R1240_U418);
  nand ginst5570 (P1_R1240_U42, P1_R1240_U118, P1_R1240_U192);
  nand ginst5571 (P1_R1240_U420, P1_R1240_U151, P1_R1240_U152);
  nand ginst5572 (P1_R1240_U421, P1_R1240_U299, P1_R1240_U419);
  nand ginst5573 (P1_R1240_U422, P1_R1240_U50, P1_U3057);
  nand ginst5574 (P1_R1240_U423, P1_R1240_U49, P1_U3976);
  nand ginst5575 (P1_R1240_U424, P1_R1240_U51, P1_U3058);
  nand ginst5576 (P1_R1240_U425, P1_R1240_U52, P1_U3977);
  nand ginst5577 (P1_R1240_U426, P1_R1240_U424, P1_R1240_U425);
  nand ginst5578 (P1_R1240_U427, P1_R1240_U356, P1_R1240_U90);
  nand ginst5579 (P1_R1240_U428, P1_R1240_U306, P1_R1240_U426);
  nand ginst5580 (P1_R1240_U429, P1_R1240_U53, P1_U3065);
  nand ginst5581 (P1_R1240_U43, P1_R1240_U181, P1_R1240_U182);
  nand ginst5582 (P1_R1240_U430, P1_R1240_U54, P1_U3978);
  nand ginst5583 (P1_R1240_U431, P1_R1240_U429, P1_R1240_U430);
  nand ginst5584 (P1_R1240_U432, P1_R1240_U154, P1_R1240_U357);
  nand ginst5585 (P1_R1240_U433, P1_R1240_U293, P1_R1240_U431);
  nand ginst5586 (P1_R1240_U434, P1_R1240_U85, P1_U3066);
  nand ginst5587 (P1_R1240_U435, P1_R1240_U86, P1_U3979);
  nand ginst5588 (P1_R1240_U436, P1_R1240_U85, P1_U3066);
  nand ginst5589 (P1_R1240_U437, P1_R1240_U86, P1_U3979);
  nand ginst5590 (P1_R1240_U438, P1_R1240_U436, P1_R1240_U437);
  nand ginst5591 (P1_R1240_U439, P1_R1240_U155, P1_R1240_U156);
  nand ginst5592 (P1_R1240_U44, P1_U3078, P1_U3455);
  nand ginst5593 (P1_R1240_U440, P1_R1240_U289, P1_R1240_U438);
  nand ginst5594 (P1_R1240_U441, P1_R1240_U83, P1_U3061);
  nand ginst5595 (P1_R1240_U442, P1_R1240_U84, P1_U3980);
  nand ginst5596 (P1_R1240_U443, P1_R1240_U83, P1_U3061);
  nand ginst5597 (P1_R1240_U444, P1_R1240_U84, P1_U3980);
  nand ginst5598 (P1_R1240_U445, P1_R1240_U443, P1_R1240_U444);
  nand ginst5599 (P1_R1240_U446, P1_R1240_U157, P1_R1240_U158);
  nand ginst5600 (P1_R1240_U447, P1_R1240_U285, P1_R1240_U445);
  nand ginst5601 (P1_R1240_U448, P1_R1240_U55, P1_U3075);
  nand ginst5602 (P1_R1240_U449, P1_R1240_U56, P1_U3981);
  nand ginst5603 (P1_R1240_U45, P1_R1240_U122, P1_R1240_U218);
  nand ginst5604 (P1_R1240_U450, P1_R1240_U55, P1_U3075);
  nand ginst5605 (P1_R1240_U451, P1_R1240_U56, P1_U3981);
  nand ginst5606 (P1_R1240_U452, P1_R1240_U450, P1_R1240_U451);
  nand ginst5607 (P1_R1240_U453, P1_R1240_U82, P1_U3076);
  nand ginst5608 (P1_R1240_U454, P1_R1240_U91, P1_U3982);
  nand ginst5609 (P1_R1240_U455, P1_R1240_U160, P1_R1240_U181);
  nand ginst5610 (P1_R1240_U456, P1_R1240_U32, P1_R1240_U327);
  nand ginst5611 (P1_R1240_U457, P1_R1240_U79, P1_U3081);
  nand ginst5612 (P1_R1240_U458, P1_R1240_U80, P1_U3508);
  nand ginst5613 (P1_R1240_U459, P1_R1240_U457, P1_R1240_U458);
  nand ginst5614 (P1_R1240_U46, P1_R1240_U214, P1_R1240_U215);
  nand ginst5615 (P1_R1240_U460, P1_R1240_U358, P1_R1240_U92);
  nand ginst5616 (P1_R1240_U461, P1_R1240_U315, P1_R1240_U459);
  nand ginst5617 (P1_R1240_U462, P1_R1240_U76, P1_U3082);
  nand ginst5618 (P1_R1240_U463, P1_R1240_U77, P1_U3506);
  nand ginst5619 (P1_R1240_U464, P1_R1240_U462, P1_R1240_U463);
  nand ginst5620 (P1_R1240_U465, P1_R1240_U161, P1_R1240_U359);
  nand ginst5621 (P1_R1240_U466, P1_R1240_U269, P1_R1240_U464);
  nand ginst5622 (P1_R1240_U467, P1_R1240_U61, P1_U3069);
  nand ginst5623 (P1_R1240_U468, P1_R1240_U59, P1_U3503);
  nand ginst5624 (P1_R1240_U469, P1_R1240_U57, P1_U3073);
  not ginst5625 (P1_R1240_U47, P1_U3975);
  nand ginst5626 (P1_R1240_U470, P1_R1240_U58, P1_U3500);
  nand ginst5627 (P1_R1240_U471, P1_R1240_U469, P1_R1240_U470);
  nand ginst5628 (P1_R1240_U472, P1_R1240_U360, P1_R1240_U93);
  nand ginst5629 (P1_R1240_U473, P1_R1240_U261, P1_R1240_U471);
  nand ginst5630 (P1_R1240_U474, P1_R1240_U74, P1_U3074);
  nand ginst5631 (P1_R1240_U475, P1_R1240_U75, P1_U3497);
  nand ginst5632 (P1_R1240_U476, P1_R1240_U74, P1_U3074);
  nand ginst5633 (P1_R1240_U477, P1_R1240_U75, P1_U3497);
  nand ginst5634 (P1_R1240_U478, P1_R1240_U476, P1_R1240_U477);
  nand ginst5635 (P1_R1240_U479, P1_R1240_U162, P1_R1240_U163);
  not ginst5636 (P1_R1240_U48, P1_U3053);
  nand ginst5637 (P1_R1240_U480, P1_R1240_U257, P1_R1240_U478);
  nand ginst5638 (P1_R1240_U481, P1_R1240_U72, P1_U3079);
  nand ginst5639 (P1_R1240_U482, P1_R1240_U73, P1_U3494);
  nand ginst5640 (P1_R1240_U483, P1_R1240_U72, P1_U3079);
  nand ginst5641 (P1_R1240_U484, P1_R1240_U73, P1_U3494);
  nand ginst5642 (P1_R1240_U485, P1_R1240_U483, P1_R1240_U484);
  nand ginst5643 (P1_R1240_U486, P1_R1240_U164, P1_R1240_U165);
  nand ginst5644 (P1_R1240_U487, P1_R1240_U253, P1_R1240_U485);
  nand ginst5645 (P1_R1240_U488, P1_R1240_U70, P1_U3080);
  nand ginst5646 (P1_R1240_U489, P1_R1240_U71, P1_U3491);
  not ginst5647 (P1_R1240_U49, P1_U3057);
  nand ginst5648 (P1_R1240_U490, P1_R1240_U65, P1_U3072);
  nand ginst5649 (P1_R1240_U491, P1_R1240_U66, P1_U3488);
  nand ginst5650 (P1_R1240_U492, P1_R1240_U490, P1_R1240_U491);
  nand ginst5651 (P1_R1240_U493, P1_R1240_U361, P1_R1240_U94);
  nand ginst5652 (P1_R1240_U494, P1_R1240_U337, P1_R1240_U492);
  nand ginst5653 (P1_R1240_U495, P1_R1240_U67, P1_U3063);
  nand ginst5654 (P1_R1240_U496, P1_R1240_U68, P1_U3485);
  nand ginst5655 (P1_R1240_U497, P1_R1240_U495, P1_R1240_U496);
  nand ginst5656 (P1_R1240_U498, P1_R1240_U166, P1_R1240_U362);
  nand ginst5657 (P1_R1240_U499, P1_R1240_U243, P1_R1240_U497);
  and ginst5658 (P1_R1240_U5, P1_R1240_U179, P1_R1240_U180);
  not ginst5659 (P1_R1240_U50, P1_U3976);
  nand ginst5660 (P1_R1240_U500, P1_R1240_U63, P1_U3062);
  nand ginst5661 (P1_R1240_U501, P1_R1240_U64, P1_U3482);
  nand ginst5662 (P1_R1240_U502, P1_R1240_U30, P1_U3077);
  nand ginst5663 (P1_R1240_U503, P1_R1240_U31, P1_U3450);
  not ginst5664 (P1_R1240_U51, P1_U3977);
  not ginst5665 (P1_R1240_U52, P1_U3058);
  not ginst5666 (P1_R1240_U53, P1_U3978);
  not ginst5667 (P1_R1240_U54, P1_U3065);
  not ginst5668 (P1_R1240_U55, P1_U3981);
  not ginst5669 (P1_R1240_U56, P1_U3075);
  not ginst5670 (P1_R1240_U57, P1_U3500);
  not ginst5671 (P1_R1240_U58, P1_U3073);
  not ginst5672 (P1_R1240_U59, P1_U3069);
  and ginst5673 (P1_R1240_U6, P1_R1240_U195, P1_R1240_U196);
  nand ginst5674 (P1_R1240_U60, P1_U3073, P1_U3500);
  not ginst5675 (P1_R1240_U61, P1_U3503);
  nand ginst5676 (P1_R1240_U62, P1_U3084, P1_U3476);
  not ginst5677 (P1_R1240_U63, P1_U3482);
  not ginst5678 (P1_R1240_U64, P1_U3062);
  not ginst5679 (P1_R1240_U65, P1_U3488);
  not ginst5680 (P1_R1240_U66, P1_U3072);
  not ginst5681 (P1_R1240_U67, P1_U3485);
  not ginst5682 (P1_R1240_U68, P1_U3063);
  nand ginst5683 (P1_R1240_U69, P1_U3063, P1_U3485);
  and ginst5684 (P1_R1240_U7, P1_R1240_U235, P1_R1240_U236);
  not ginst5685 (P1_R1240_U70, P1_U3491);
  not ginst5686 (P1_R1240_U71, P1_U3080);
  not ginst5687 (P1_R1240_U72, P1_U3494);
  not ginst5688 (P1_R1240_U73, P1_U3079);
  not ginst5689 (P1_R1240_U74, P1_U3497);
  not ginst5690 (P1_R1240_U75, P1_U3074);
  not ginst5691 (P1_R1240_U76, P1_U3506);
  not ginst5692 (P1_R1240_U77, P1_U3082);
  nand ginst5693 (P1_R1240_U78, P1_U3082, P1_U3506);
  not ginst5694 (P1_R1240_U79, P1_U3508);
  and ginst5695 (P1_R1240_U8, P1_R1240_U244, P1_R1240_U245);
  not ginst5696 (P1_R1240_U80, P1_U3081);
  nand ginst5697 (P1_R1240_U81, P1_U3081, P1_U3508);
  not ginst5698 (P1_R1240_U82, P1_U3982);
  not ginst5699 (P1_R1240_U83, P1_U3980);
  not ginst5700 (P1_R1240_U84, P1_U3061);
  not ginst5701 (P1_R1240_U85, P1_U3979);
  not ginst5702 (P1_R1240_U86, P1_U3066);
  nand ginst5703 (P1_R1240_U87, P1_U3057, P1_U3976);
  not ginst5704 (P1_R1240_U88, P1_U3054);
  not ginst5705 (P1_R1240_U89, P1_U3974);
  and ginst5706 (P1_R1240_U9, P1_R1240_U262, P1_R1240_U263);
  nand ginst5707 (P1_R1240_U90, P1_R1240_U175, P1_R1240_U305);
  not ginst5708 (P1_R1240_U91, P1_U3076);
  nand ginst5709 (P1_R1240_U92, P1_R1240_U314, P1_R1240_U78);
  nand ginst5710 (P1_R1240_U93, P1_R1240_U259, P1_R1240_U260);
  nand ginst5711 (P1_R1240_U94, P1_R1240_U336, P1_R1240_U69);
  nand ginst5712 (P1_R1240_U95, P1_R1240_U455, P1_R1240_U456);
  nand ginst5713 (P1_R1240_U96, P1_R1240_U502, P1_R1240_U503);
  nand ginst5714 (P1_R1240_U97, P1_R1240_U373, P1_R1240_U374);
  nand ginst5715 (P1_R1240_U98, P1_R1240_U378, P1_R1240_U379);
  nand ginst5716 (P1_R1240_U99, P1_R1240_U385, P1_R1240_U386);
  and ginst5717 (P1_R1282_U10, P1_R1282_U129, P1_R1282_U39);
  not ginst5718 (P1_R1282_U100, P1_R1282_U36);
  not ginst5719 (P1_R1282_U101, P1_R1282_U37);
  not ginst5720 (P1_R1282_U102, P1_R1282_U38);
  not ginst5721 (P1_R1282_U103, P1_R1282_U39);
  not ginst5722 (P1_R1282_U104, P1_R1282_U40);
  not ginst5723 (P1_R1282_U105, P1_R1282_U41);
  not ginst5724 (P1_R1282_U106, P1_R1282_U42);
  not ginst5725 (P1_R1282_U107, P1_R1282_U43);
  not ginst5726 (P1_R1282_U108, P1_R1282_U44);
  not ginst5727 (P1_R1282_U109, P1_R1282_U45);
  and ginst5728 (P1_R1282_U11, P1_R1282_U128, P1_R1282_U40);
  not ginst5729 (P1_R1282_U110, P1_R1282_U46);
  not ginst5730 (P1_R1282_U111, P1_R1282_U67);
  nand ginst5731 (P1_R1282_U112, P1_R1282_U110, P1_R1282_U69);
  nand ginst5732 (P1_R1282_U113, P1_R1282_U112, P1_U3984);
  or ginst5733 (P1_R1282_U114, P1_U3450, P1_U3455);
  nand ginst5734 (P1_R1282_U115, P1_R1282_U114, P1_U3458);
  nand ginst5735 (P1_R1282_U116, P1_R1282_U109, P1_R1282_U71);
  nand ginst5736 (P1_R1282_U117, P1_R1282_U116, P1_U3974);
  nand ginst5737 (P1_R1282_U118, P1_R1282_U108, P1_R1282_U73);
  nand ginst5738 (P1_R1282_U119, P1_R1282_U118, P1_U3976);
  and ginst5739 (P1_R1282_U12, P1_R1282_U127, P1_R1282_U41);
  nand ginst5740 (P1_R1282_U120, P1_R1282_U107, P1_R1282_U75);
  nand ginst5741 (P1_R1282_U121, P1_R1282_U120, P1_U3978);
  nand ginst5742 (P1_R1282_U122, P1_R1282_U106, P1_R1282_U77);
  nand ginst5743 (P1_R1282_U123, P1_R1282_U122, P1_U3980);
  nand ginst5744 (P1_R1282_U124, P1_R1282_U105, P1_R1282_U81);
  nand ginst5745 (P1_R1282_U125, P1_R1282_U124, P1_U3982);
  nand ginst5746 (P1_R1282_U126, P1_R1282_U104, P1_R1282_U83);
  nand ginst5747 (P1_R1282_U127, P1_R1282_U126, P1_U3506);
  nand ginst5748 (P1_R1282_U128, P1_R1282_U39, P1_U3500);
  nand ginst5749 (P1_R1282_U129, P1_R1282_U38, P1_U3497);
  and ginst5750 (P1_R1282_U13, P1_R1282_U125, P1_R1282_U42);
  nand ginst5751 (P1_R1282_U130, P1_R1282_U101, P1_R1282_U85);
  nand ginst5752 (P1_R1282_U131, P1_R1282_U130, P1_U3494);
  nand ginst5753 (P1_R1282_U132, P1_R1282_U36, P1_U3488);
  nand ginst5754 (P1_R1282_U133, P1_R1282_U35, P1_U3485);
  nand ginst5755 (P1_R1282_U134, P1_R1282_U62, P1_R1282_U92);
  nand ginst5756 (P1_R1282_U135, P1_R1282_U134, P1_U3482);
  nand ginst5757 (P1_R1282_U136, P1_R1282_U30, P1_U3479);
  nand ginst5758 (P1_R1282_U137, P1_R1282_U62, P1_R1282_U92);
  nand ginst5759 (P1_R1282_U138, P1_R1282_U27, P1_U3467);
  nand ginst5760 (P1_R1282_U139, P1_R1282_U64, P1_R1282_U89);
  and ginst5761 (P1_R1282_U14, P1_R1282_U123, P1_R1282_U43);
  nand ginst5762 (P1_R1282_U140, P1_R1282_U67, P1_U3983);
  nand ginst5763 (P1_R1282_U141, P1_R1282_U111, P1_R1282_U66);
  nand ginst5764 (P1_R1282_U142, P1_R1282_U46, P1_U3985);
  nand ginst5765 (P1_R1282_U143, P1_R1282_U110, P1_R1282_U69);
  nand ginst5766 (P1_R1282_U144, P1_R1282_U45, P1_U3975);
  nand ginst5767 (P1_R1282_U145, P1_R1282_U109, P1_R1282_U71);
  nand ginst5768 (P1_R1282_U146, P1_R1282_U44, P1_U3977);
  nand ginst5769 (P1_R1282_U147, P1_R1282_U108, P1_R1282_U73);
  nand ginst5770 (P1_R1282_U148, P1_R1282_U43, P1_U3979);
  nand ginst5771 (P1_R1282_U149, P1_R1282_U107, P1_R1282_U75);
  and ginst5772 (P1_R1282_U15, P1_R1282_U121, P1_R1282_U44);
  nand ginst5773 (P1_R1282_U150, P1_R1282_U42, P1_U3981);
  nand ginst5774 (P1_R1282_U151, P1_R1282_U106, P1_R1282_U77);
  nand ginst5775 (P1_R1282_U152, P1_R1282_U80, P1_U3455);
  nand ginst5776 (P1_R1282_U153, P1_R1282_U79, P1_U3450);
  nand ginst5777 (P1_R1282_U154, P1_R1282_U41, P1_U3508);
  nand ginst5778 (P1_R1282_U155, P1_R1282_U105, P1_R1282_U81);
  nand ginst5779 (P1_R1282_U156, P1_R1282_U40, P1_U3503);
  nand ginst5780 (P1_R1282_U157, P1_R1282_U104, P1_R1282_U83);
  nand ginst5781 (P1_R1282_U158, P1_R1282_U37, P1_U3491);
  nand ginst5782 (P1_R1282_U159, P1_R1282_U101, P1_R1282_U85);
  and ginst5783 (P1_R1282_U16, P1_R1282_U119, P1_R1282_U45);
  and ginst5784 (P1_R1282_U17, P1_R1282_U117, P1_R1282_U46);
  and ginst5785 (P1_R1282_U18, P1_R1282_U115, P1_R1282_U25);
  and ginst5786 (P1_R1282_U19, P1_R1282_U113, P1_R1282_U67);
  and ginst5787 (P1_R1282_U20, P1_R1282_U26, P1_R1282_U98);
  and ginst5788 (P1_R1282_U21, P1_R1282_U27, P1_R1282_U97);
  and ginst5789 (P1_R1282_U22, P1_R1282_U28, P1_R1282_U96);
  and ginst5790 (P1_R1282_U23, P1_R1282_U29, P1_R1282_U94);
  and ginst5791 (P1_R1282_U24, P1_R1282_U30, P1_R1282_U93);
  or ginst5792 (P1_R1282_U25, P1_U3450, P1_U3455, P1_U3458);
  nand ginst5793 (P1_R1282_U26, P1_R1282_U34, P1_R1282_U87);
  nand ginst5794 (P1_R1282_U27, P1_R1282_U33, P1_R1282_U88);
  nand ginst5795 (P1_R1282_U28, P1_R1282_U58, P1_R1282_U89);
  nand ginst5796 (P1_R1282_U29, P1_R1282_U32, P1_R1282_U90);
  nand ginst5797 (P1_R1282_U30, P1_R1282_U31, P1_R1282_U91);
  not ginst5798 (P1_R1282_U31, P1_U3476);
  not ginst5799 (P1_R1282_U32, P1_U3473);
  not ginst5800 (P1_R1282_U33, P1_U3464);
  not ginst5801 (P1_R1282_U34, P1_U3461);
  nand ginst5802 (P1_R1282_U35, P1_R1282_U59, P1_R1282_U92);
  nand ginst5803 (P1_R1282_U36, P1_R1282_U56, P1_R1282_U99);
  nand ginst5804 (P1_R1282_U37, P1_R1282_U100, P1_R1282_U55);
  nand ginst5805 (P1_R1282_U38, P1_R1282_U101, P1_R1282_U60);
  nand ginst5806 (P1_R1282_U39, P1_R1282_U102, P1_R1282_U54);
  nand ginst5807 (P1_R1282_U40, P1_R1282_U103, P1_R1282_U53);
  nand ginst5808 (P1_R1282_U41, P1_R1282_U104, P1_R1282_U61);
  nand ginst5809 (P1_R1282_U42, P1_R1282_U105, P1_R1282_U52, P1_R1282_U81);
  nand ginst5810 (P1_R1282_U43, P1_R1282_U106, P1_R1282_U51, P1_R1282_U77);
  nand ginst5811 (P1_R1282_U44, P1_R1282_U107, P1_R1282_U50, P1_R1282_U75);
  nand ginst5812 (P1_R1282_U45, P1_R1282_U108, P1_R1282_U49, P1_R1282_U73);
  nand ginst5813 (P1_R1282_U46, P1_R1282_U109, P1_R1282_U48, P1_R1282_U71);
  not ginst5814 (P1_R1282_U47, P1_U3984);
  not ginst5815 (P1_R1282_U48, P1_U3974);
  not ginst5816 (P1_R1282_U49, P1_U3976);
  not ginst5817 (P1_R1282_U50, P1_U3978);
  not ginst5818 (P1_R1282_U51, P1_U3980);
  not ginst5819 (P1_R1282_U52, P1_U3982);
  not ginst5820 (P1_R1282_U53, P1_U3500);
  not ginst5821 (P1_R1282_U54, P1_U3497);
  not ginst5822 (P1_R1282_U55, P1_U3488);
  not ginst5823 (P1_R1282_U56, P1_U3485);
  nand ginst5824 (P1_R1282_U57, P1_R1282_U152, P1_R1282_U153);
  nor ginst5825 (P1_R1282_U58, P1_U3467, P1_U3470);
  nor ginst5826 (P1_R1282_U59, P1_U3479, P1_U3482);
  and ginst5827 (P1_R1282_U6, P1_R1282_U135, P1_R1282_U35);
  nor ginst5828 (P1_R1282_U60, P1_U3491, P1_U3494);
  nor ginst5829 (P1_R1282_U61, P1_U3503, P1_U3506);
  not ginst5830 (P1_R1282_U62, P1_U3479);
  and ginst5831 (P1_R1282_U63, P1_R1282_U136, P1_R1282_U137);
  not ginst5832 (P1_R1282_U64, P1_U3467);
  and ginst5833 (P1_R1282_U65, P1_R1282_U138, P1_R1282_U139);
  not ginst5834 (P1_R1282_U66, P1_U3983);
  nand ginst5835 (P1_R1282_U67, P1_R1282_U110, P1_R1282_U47, P1_R1282_U69);
  and ginst5836 (P1_R1282_U68, P1_R1282_U140, P1_R1282_U141);
  not ginst5837 (P1_R1282_U69, P1_U3985);
  and ginst5838 (P1_R1282_U7, P1_R1282_U133, P1_R1282_U36);
  and ginst5839 (P1_R1282_U70, P1_R1282_U142, P1_R1282_U143);
  not ginst5840 (P1_R1282_U71, P1_U3975);
  and ginst5841 (P1_R1282_U72, P1_R1282_U144, P1_R1282_U145);
  not ginst5842 (P1_R1282_U73, P1_U3977);
  and ginst5843 (P1_R1282_U74, P1_R1282_U146, P1_R1282_U147);
  not ginst5844 (P1_R1282_U75, P1_U3979);
  and ginst5845 (P1_R1282_U76, P1_R1282_U148, P1_R1282_U149);
  not ginst5846 (P1_R1282_U77, P1_U3981);
  and ginst5847 (P1_R1282_U78, P1_R1282_U150, P1_R1282_U151);
  not ginst5848 (P1_R1282_U79, P1_U3455);
  and ginst5849 (P1_R1282_U8, P1_R1282_U132, P1_R1282_U37);
  not ginst5850 (P1_R1282_U80, P1_U3450);
  not ginst5851 (P1_R1282_U81, P1_U3508);
  and ginst5852 (P1_R1282_U82, P1_R1282_U154, P1_R1282_U155);
  not ginst5853 (P1_R1282_U83, P1_U3503);
  and ginst5854 (P1_R1282_U84, P1_R1282_U156, P1_R1282_U157);
  not ginst5855 (P1_R1282_U85, P1_U3491);
  and ginst5856 (P1_R1282_U86, P1_R1282_U158, P1_R1282_U159);
  not ginst5857 (P1_R1282_U87, P1_R1282_U25);
  not ginst5858 (P1_R1282_U88, P1_R1282_U26);
  not ginst5859 (P1_R1282_U89, P1_R1282_U27);
  and ginst5860 (P1_R1282_U9, P1_R1282_U131, P1_R1282_U38);
  not ginst5861 (P1_R1282_U90, P1_R1282_U28);
  not ginst5862 (P1_R1282_U91, P1_R1282_U29);
  not ginst5863 (P1_R1282_U92, P1_R1282_U30);
  nand ginst5864 (P1_R1282_U93, P1_R1282_U29, P1_U3476);
  nand ginst5865 (P1_R1282_U94, P1_R1282_U28, P1_U3473);
  nand ginst5866 (P1_R1282_U95, P1_R1282_U64, P1_R1282_U89);
  nand ginst5867 (P1_R1282_U96, P1_R1282_U95, P1_U3470);
  nand ginst5868 (P1_R1282_U97, P1_R1282_U26, P1_U3464);
  nand ginst5869 (P1_R1282_U98, P1_R1282_U25, P1_U3461);
  not ginst5870 (P1_R1282_U99, P1_R1282_U35);
  nand ginst5871 (P1_R1309_U10, P1_R1309_U7, P1_U3059);
  not ginst5872 (P1_R1309_U6, P1_U3059);
  not ginst5873 (P1_R1309_U7, P1_U3056);
  and ginst5874 (P1_R1309_U8, P1_R1309_U10, P1_R1309_U9);
  nand ginst5875 (P1_R1309_U9, P1_R1309_U6, P1_U3056);
  and ginst5876 (P1_R1352_U6, P1_R1352_U7, P1_U3059);
  not ginst5877 (P1_R1352_U7, P1_U3056);
  and ginst5878 (P1_R1360_U10, P1_R1360_U183, P1_R1360_U184, P1_R1360_U185, P1_R1360_U186, P1_R1360_U199);
  and ginst5879 (P1_R1360_U100, P1_R1360_U170, P1_R1360_U171);
  and ginst5880 (P1_R1360_U101, P1_R1360_U179, P1_R1360_U180);
  and ginst5881 (P1_R1360_U102, P1_R1360_U23, P1_U3095);
  and ginst5882 (P1_R1360_U103, P1_R1360_U67, P1_U3096);
  and ginst5883 (P1_R1360_U104, P1_R1360_U106, P1_R1360_U181, P1_R1360_U184, P1_R1360_U185, P1_R1360_U186);
  and ginst5884 (P1_R1360_U105, P1_R1360_U189, P1_R1360_U190);
  and ginst5885 (P1_R1360_U106, P1_R1360_U105, P1_R1360_U187, P1_R1360_U188);
  and ginst5886 (P1_R1360_U107, P1_R1360_U194, P1_R1360_U195, P1_R1360_U196);
  and ginst5887 (P1_R1360_U108, P1_R1360_U13, P1_R1360_U201);
  not ginst5888 (P1_R1360_U109, P1_U3119);
  and ginst5889 (P1_R1360_U11, P1_R1360_U104, P1_R1360_U183);
  nand ginst5890 (P1_R1360_U110, P1_R1360_U66, P1_U3097);
  nand ginst5891 (P1_R1360_U111, P1_R1360_U73, P1_U3126);
  nand ginst5892 (P1_R1360_U112, P1_R1360_U70, P1_U3127);
  nand ginst5893 (P1_R1360_U113, P1_R1360_U65, P1_U3098);
  nand ginst5894 (P1_R1360_U114, P1_R1360_U58, P1_U3103);
  nand ginst5895 (P1_R1360_U115, P1_R1360_U61, P1_U3133);
  nand ginst5896 (P1_R1360_U116, P1_R1360_U62, P1_U3132);
  nand ginst5897 (P1_R1360_U117, P1_R1360_U57, P1_U3104);
  nand ginst5898 (P1_R1360_U118, P1_R1360_U50, P1_U3109);
  nand ginst5899 (P1_R1360_U119, P1_R1360_U34, P1_U3110);
  and ginst5900 (P1_R1360_U12, P1_R1360_U202, P1_R1360_U203);
  nand ginst5901 (P1_R1360_U120, P1_R1360_U49, P1_U3112);
  nand ginst5902 (P1_R1360_U121, P1_R1360_U36, P1_U3111);
  nand ginst5903 (P1_R1360_U122, P1_R1360_U54, P1_U3139);
  nand ginst5904 (P1_R1360_U123, P1_R1360_U53, P1_U3138);
  nand ginst5905 (P1_R1360_U124, P1_R1360_U47, P1_U3114);
  nand ginst5906 (P1_R1360_U125, P1_R1360_U48, P1_U3113);
  nand ginst5907 (P1_R1360_U126, P1_R1360_U45, P1_U3116);
  nand ginst5908 (P1_R1360_U127, P1_R1360_U46, P1_U3115);
  nand ginst5909 (P1_R1360_U128, P1_U3150, P1_U3151);
  nand ginst5910 (P1_R1360_U129, P1_R1360_U128, P1_U3118);
  and ginst5911 (P1_R1360_U13, P1_R1360_U204, P1_R1360_U205);
  or ginst5912 (P1_R1360_U130, P1_U3150, P1_U3151);
  nand ginst5913 (P1_R1360_U131, P1_R1360_U44, P1_U3117);
  nand ginst5914 (P1_R1360_U132, P1_R1360_U81, P1_R1360_U82);
  nand ginst5915 (P1_R1360_U133, P1_R1360_U126, P1_R1360_U83);
  nand ginst5916 (P1_R1360_U134, P1_R1360_U41, P1_U3148);
  nand ginst5917 (P1_R1360_U135, P1_R1360_U133, P1_R1360_U134);
  nand ginst5918 (P1_R1360_U136, P1_R1360_U127, P1_R1360_U135);
  nand ginst5919 (P1_R1360_U137, P1_R1360_U42, P1_U3147);
  nand ginst5920 (P1_R1360_U138, P1_R1360_U136, P1_R1360_U137);
  nand ginst5921 (P1_R1360_U139, P1_R1360_U124, P1_R1360_U138);
  nand ginst5922 (P1_R1360_U14, P1_R1360_U107, P1_R1360_U108, P1_R1360_U200);
  nand ginst5923 (P1_R1360_U140, P1_R1360_U39, P1_U3146);
  nand ginst5924 (P1_R1360_U141, P1_R1360_U139, P1_R1360_U140);
  nand ginst5925 (P1_R1360_U142, P1_R1360_U125, P1_R1360_U141);
  nand ginst5926 (P1_R1360_U143, P1_R1360_U40, P1_U3145);
  nand ginst5927 (P1_R1360_U144, P1_R1360_U37, P1_U3144);
  nand ginst5928 (P1_R1360_U145, P1_R1360_U142, P1_R1360_U84);
  nand ginst5929 (P1_R1360_U146, P1_R1360_U118, P1_R1360_U79);
  nand ginst5930 (P1_R1360_U147, P1_R1360_U8, P1_R1360_U80);
  nand ginst5931 (P1_R1360_U148, P1_R1360_U145, P1_R1360_U87);
  nand ginst5932 (P1_R1360_U149, P1_R1360_U33, P1_U3141);
  not ginst5933 (P1_R1360_U15, P1_U3088);
  nand ginst5934 (P1_R1360_U150, P1_R1360_U52, P1_U3140);
  nand ginst5935 (P1_R1360_U151, P1_R1360_U148, P1_R1360_U88);
  nand ginst5936 (P1_R1360_U152, P1_R1360_U9, P1_R1360_U91);
  nand ginst5937 (P1_R1360_U153, P1_R1360_U32, P1_U3106);
  nand ginst5938 (P1_R1360_U154, P1_R1360_U53, P1_U3138);
  nand ginst5939 (P1_R1360_U155, P1_R1360_U154, P1_R1360_U92);
  nand ginst5940 (P1_R1360_U156, P1_R1360_U56, P1_U3105);
  nand ginst5941 (P1_R1360_U157, P1_R1360_U151, P1_R1360_U93);
  nand ginst5942 (P1_R1360_U158, P1_R1360_U55, P1_U3137);
  nand ginst5943 (P1_R1360_U159, P1_R1360_U157, P1_R1360_U158);
  not ginst5944 (P1_R1360_U16, P1_U3087);
  nand ginst5945 (P1_R1360_U160, P1_R1360_U117, P1_R1360_U159);
  nand ginst5946 (P1_R1360_U161, P1_R1360_U30, P1_U3136);
  nand ginst5947 (P1_R1360_U162, P1_R1360_U160, P1_R1360_U161);
  nand ginst5948 (P1_R1360_U163, P1_R1360_U114, P1_R1360_U162);
  nand ginst5949 (P1_R1360_U164, P1_R1360_U29, P1_U3135);
  nand ginst5950 (P1_R1360_U165, P1_R1360_U60, P1_U3134);
  nand ginst5951 (P1_R1360_U166, P1_R1360_U163, P1_R1360_U95);
  nand ginst5952 (P1_R1360_U167, P1_R1360_U7, P1_R1360_U97);
  nand ginst5953 (P1_R1360_U168, P1_R1360_U62, P1_U3132);
  nand ginst5954 (P1_R1360_U169, P1_R1360_U168, P1_R1360_U98);
  not ginst5955 (P1_R1360_U17, P1_U3121);
  nand ginst5956 (P1_R1360_U170, P1_R1360_U28, P1_U3100);
  nand ginst5957 (P1_R1360_U171, P1_R1360_U64, P1_U3099);
  nand ginst5958 (P1_R1360_U172, P1_R1360_U166, P1_R1360_U99);
  nand ginst5959 (P1_R1360_U173, P1_R1360_U63, P1_U3131);
  nand ginst5960 (P1_R1360_U174, P1_R1360_U172, P1_R1360_U173);
  nand ginst5961 (P1_R1360_U175, P1_R1360_U113, P1_R1360_U174);
  nand ginst5962 (P1_R1360_U176, P1_R1360_U26, P1_U3130);
  nand ginst5963 (P1_R1360_U177, P1_R1360_U175, P1_R1360_U176);
  nand ginst5964 (P1_R1360_U178, P1_R1360_U110, P1_R1360_U177);
  nand ginst5965 (P1_R1360_U179, P1_R1360_U25, P1_U3129);
  not ginst5966 (P1_R1360_U18, P1_U3089);
  nand ginst5967 (P1_R1360_U180, P1_R1360_U71, P1_U3128);
  nand ginst5968 (P1_R1360_U181, P1_R1360_U101, P1_R1360_U178, P1_R1360_U6);
  nand ginst5969 (P1_R1360_U182, P1_R1360_U22, P1_U3088);
  nand ginst5970 (P1_R1360_U183, P1_R1360_U17, P1_U3089);
  nand ginst5971 (P1_R1360_U184, P1_R1360_U21, P1_U3090);
  nand ginst5972 (P1_R1360_U185, P1_R1360_U74, P1_U3092);
  nand ginst5973 (P1_R1360_U186, P1_R1360_U20, P1_U3091);
  nand ginst5974 (P1_R1360_U187, P1_R1360_U102, P1_R1360_U111);
  nand ginst5975 (P1_R1360_U188, P1_R1360_U103, P1_R1360_U6);
  nand ginst5976 (P1_R1360_U189, P1_R1360_U75, P1_U3093);
  not ginst5977 (P1_R1360_U19, P1_U3090);
  nand ginst5978 (P1_R1360_U190, P1_R1360_U24, P1_U3094);
  nand ginst5979 (P1_R1360_U191, P1_R1360_U69, P1_U3123);
  nand ginst5980 (P1_R1360_U192, P1_R1360_U19, P1_U3122);
  nand ginst5981 (P1_R1360_U193, P1_R1360_U191, P1_R1360_U192);
  nand ginst5982 (P1_R1360_U194, P1_R1360_U12, P1_R1360_U182, P1_R1360_U77);
  nand ginst5983 (P1_R1360_U195, P1_R1360_U12, P1_R1360_U182, P1_R1360_U193, P1_R1360_U78);
  nand ginst5984 (P1_R1360_U196, P1_R1360_U12, P1_R1360_U15, P1_U3120);
  nand ginst5985 (P1_R1360_U197, P1_R1360_U68, P1_U3124);
  nand ginst5986 (P1_R1360_U198, P1_R1360_U72, P1_U3125);
  nand ginst5987 (P1_R1360_U199, P1_R1360_U197, P1_R1360_U198);
  not ginst5988 (P1_R1360_U20, P1_U3123);
  nand ginst5989 (P1_R1360_U200, P1_R1360_U11, P1_R1360_U12, P1_R1360_U182);
  nand ginst5990 (P1_R1360_U201, P1_R1360_U10, P1_R1360_U12, P1_R1360_U182);
  nand ginst5991 (P1_R1360_U202, P1_R1360_U109, P1_U3087);
  nand ginst5992 (P1_R1360_U203, P1_R1360_U16, P1_U3119);
  nand ginst5993 (P1_R1360_U204, P1_R1360_U109, P1_U3087, P1_U3152);
  nand ginst5994 (P1_R1360_U205, P1_R1360_U16, P1_R1360_U76, P1_U3119);
  not ginst5995 (P1_R1360_U21, P1_U3122);
  not ginst5996 (P1_R1360_U22, P1_U3120);
  not ginst5997 (P1_R1360_U23, P1_U3127);
  not ginst5998 (P1_R1360_U24, P1_U3126);
  not ginst5999 (P1_R1360_U25, P1_U3097);
  not ginst6000 (P1_R1360_U26, P1_U3098);
  not ginst6001 (P1_R1360_U27, P1_U3133);
  not ginst6002 (P1_R1360_U28, P1_U3132);
  not ginst6003 (P1_R1360_U29, P1_U3103);
  not ginst6004 (P1_R1360_U30, P1_U3104);
  not ginst6005 (P1_R1360_U31, P1_U3139);
  not ginst6006 (P1_R1360_U32, P1_U3138);
  not ginst6007 (P1_R1360_U33, P1_U3109);
  not ginst6008 (P1_R1360_U34, P1_U3142);
  not ginst6009 (P1_R1360_U35, P1_U3110);
  not ginst6010 (P1_R1360_U36, P1_U3143);
  not ginst6011 (P1_R1360_U37, P1_U3112);
  not ginst6012 (P1_R1360_U38, P1_U3111);
  not ginst6013 (P1_R1360_U39, P1_U3114);
  not ginst6014 (P1_R1360_U40, P1_U3113);
  not ginst6015 (P1_R1360_U41, P1_U3116);
  not ginst6016 (P1_R1360_U42, P1_U3115);
  not ginst6017 (P1_R1360_U43, P1_U3117);
  not ginst6018 (P1_R1360_U44, P1_U3149);
  not ginst6019 (P1_R1360_U45, P1_U3148);
  not ginst6020 (P1_R1360_U46, P1_U3147);
  not ginst6021 (P1_R1360_U47, P1_U3146);
  not ginst6022 (P1_R1360_U48, P1_U3145);
  not ginst6023 (P1_R1360_U49, P1_U3144);
  not ginst6024 (P1_R1360_U50, P1_U3141);
  not ginst6025 (P1_R1360_U51, P1_U3140);
  not ginst6026 (P1_R1360_U52, P1_U3108);
  not ginst6027 (P1_R1360_U53, P1_U3106);
  not ginst6028 (P1_R1360_U54, P1_U3107);
  not ginst6029 (P1_R1360_U55, P1_U3105);
  not ginst6030 (P1_R1360_U56, P1_U3137);
  not ginst6031 (P1_R1360_U57, P1_U3136);
  not ginst6032 (P1_R1360_U58, P1_U3135);
  not ginst6033 (P1_R1360_U59, P1_U3134);
  and ginst6034 (P1_R1360_U6, P1_R1360_U111, P1_R1360_U112);
  not ginst6035 (P1_R1360_U60, P1_U3102);
  not ginst6036 (P1_R1360_U61, P1_U3101);
  not ginst6037 (P1_R1360_U62, P1_U3100);
  not ginst6038 (P1_R1360_U63, P1_U3099);
  not ginst6039 (P1_R1360_U64, P1_U3131);
  not ginst6040 (P1_R1360_U65, P1_U3130);
  not ginst6041 (P1_R1360_U66, P1_U3129);
  not ginst6042 (P1_R1360_U67, P1_U3128);
  not ginst6043 (P1_R1360_U68, P1_U3092);
  not ginst6044 (P1_R1360_U69, P1_U3091);
  and ginst6045 (P1_R1360_U7, P1_R1360_U115, P1_R1360_U116);
  not ginst6046 (P1_R1360_U70, P1_U3095);
  not ginst6047 (P1_R1360_U71, P1_U3096);
  not ginst6048 (P1_R1360_U72, P1_U3093);
  not ginst6049 (P1_R1360_U73, P1_U3094);
  not ginst6050 (P1_R1360_U74, P1_U3124);
  not ginst6051 (P1_R1360_U75, P1_U3125);
  not ginst6052 (P1_R1360_U76, P1_U3152);
  and ginst6053 (P1_R1360_U77, P1_R1360_U18, P1_U3121);
  and ginst6054 (P1_R1360_U78, P1_R1360_U183, P1_R1360_U184);
  and ginst6055 (P1_R1360_U79, P1_R1360_U35, P1_U3142);
  and ginst6056 (P1_R1360_U8, P1_R1360_U118, P1_R1360_U119);
  and ginst6057 (P1_R1360_U80, P1_R1360_U38, P1_U3143);
  and ginst6058 (P1_R1360_U81, P1_R1360_U124, P1_R1360_U125, P1_R1360_U126, P1_R1360_U127);
  and ginst6059 (P1_R1360_U82, P1_R1360_U129, P1_R1360_U130, P1_R1360_U131);
  and ginst6060 (P1_R1360_U83, P1_R1360_U43, P1_U3149);
  and ginst6061 (P1_R1360_U84, P1_R1360_U132, P1_R1360_U85);
  and ginst6062 (P1_R1360_U85, P1_R1360_U143, P1_R1360_U144);
  and ginst6063 (P1_R1360_U86, P1_R1360_U120, P1_R1360_U121);
  and ginst6064 (P1_R1360_U87, P1_R1360_U8, P1_R1360_U86);
  and ginst6065 (P1_R1360_U88, P1_R1360_U146, P1_R1360_U147, P1_R1360_U90);
  and ginst6066 (P1_R1360_U89, P1_R1360_U149, P1_R1360_U150);
  and ginst6067 (P1_R1360_U9, P1_R1360_U122, P1_R1360_U123);
  and ginst6068 (P1_R1360_U90, P1_R1360_U89, P1_R1360_U9);
  and ginst6069 (P1_R1360_U91, P1_R1360_U51, P1_U3108);
  and ginst6070 (P1_R1360_U92, P1_R1360_U31, P1_U3107);
  and ginst6071 (P1_R1360_U93, P1_R1360_U152, P1_R1360_U153, P1_R1360_U94);
  and ginst6072 (P1_R1360_U94, P1_R1360_U155, P1_R1360_U156);
  and ginst6073 (P1_R1360_U95, P1_R1360_U7, P1_R1360_U96);
  and ginst6074 (P1_R1360_U96, P1_R1360_U164, P1_R1360_U165);
  and ginst6075 (P1_R1360_U97, P1_R1360_U59, P1_U3102);
  and ginst6076 (P1_R1360_U98, P1_R1360_U27, P1_U3101);
  and ginst6077 (P1_R1360_U99, P1_R1360_U100, P1_R1360_U167, P1_R1360_U169);
  and ginst6078 (P1_R1375_U10, P1_R1375_U196, P1_R1375_U197, P1_R1375_U198, P1_R1375_U6);
  and ginst6079 (P1_R1375_U100, P1_R1375_U52, P1_U3063);
  and ginst6080 (P1_R1375_U101, P1_R1375_U102, P1_R1375_U173, P1_R1375_U174);
  and ginst6081 (P1_R1375_U102, P1_R1375_U176, P1_R1375_U177);
  and ginst6082 (P1_R1375_U103, P1_R1375_U104, P1_R1375_U7);
  and ginst6083 (P1_R1375_U104, P1_R1375_U185, P1_R1375_U186);
  and ginst6084 (P1_R1375_U105, P1_R1375_U69, P1_U3073);
  and ginst6085 (P1_R1375_U106, P1_R1375_U35, P1_U3069);
  and ginst6086 (P1_R1375_U107, P1_R1375_U108, P1_R1375_U188, P1_R1375_U190);
  and ginst6087 (P1_R1375_U108, P1_R1375_U191, P1_R1375_U192);
  and ginst6088 (P1_R1375_U109, P1_R1375_U133, P1_R1375_U134);
  and ginst6089 (P1_R1375_U11, P1_R1375_U20, P1_U3985);
  and ginst6090 (P1_R1375_U110, P1_R1375_U34, P1_U3982);
  and ginst6091 (P1_R1375_U111, P1_R1375_U127, P1_R1375_U128);
  and ginst6092 (P1_R1375_U112, P1_R1375_U10, P1_R1375_U129, P1_R1375_U130, P1_R1375_U131);
  not ginst6093 (P1_R1375_U113, P1_U3053);
  nand ginst6094 (P1_R1375_U114, P1_R1375_U199, P1_R1375_U200);
  nand ginst6095 (P1_R1375_U115, P1_R1375_U17, P1_U3983);
  nand ginst6096 (P1_R1375_U116, P1_R1375_U18, P1_U3055);
  nand ginst6097 (P1_R1375_U117, P1_R1375_U25, P1_U3054);
  nand ginst6098 (P1_R1375_U118, P1_R1375_U26, P1_U3057);
  nand ginst6099 (P1_R1375_U119, P1_R1375_U32, P1_U3978);
  and ginst6100 (P1_R1375_U12, P1_R1375_U117, P1_R1375_U118, P1_R1375_U206, P1_R1375_U207);
  nand ginst6101 (P1_R1375_U120, P1_R1375_U28, P1_U3979);
  nand ginst6102 (P1_R1375_U121, P1_R1375_U119, P1_R1375_U85);
  nand ginst6103 (P1_R1375_U122, P1_R1375_U6, P1_R1375_U86);
  nand ginst6104 (P1_R1375_U123, P1_R1375_U24, P1_U3058);
  nand ginst6105 (P1_R1375_U124, P1_R1375_U27, P1_U3065);
  nand ginst6106 (P1_R1375_U125, P1_R1375_U16, P1_U3059);
  nand ginst6107 (P1_R1375_U126, P1_R1375_U115, P1_R1375_U117, P1_R1375_U81);
  nand ginst6108 (P1_R1375_U127, P1_R1375_U115, P1_R1375_U12, P1_R1375_U82);
  nand ginst6109 (P1_R1375_U128, P1_R1375_U115, P1_R1375_U19, P1_U3984);
  nand ginst6110 (P1_R1375_U129, P1_R1375_U115, P1_R1375_U83);
  and ginst6111 (P1_R1375_U13, P1_R1375_U48, P1_U3450);
  nand ginst6112 (P1_R1375_U130, P1_R1375_U115, P1_R1375_U12, P1_R1375_U84);
  nand ginst6113 (P1_R1375_U131, P1_R1375_U15, P1_U3056);
  nand ginst6114 (P1_R1375_U132, P1_R1375_U127, P1_R1375_U130, P1_R1375_U79, P1_R1375_U88);
  nand ginst6115 (P1_R1375_U133, P1_R1375_U76, P1_U3075);
  nand ginst6116 (P1_R1375_U134, P1_R1375_U75, P1_U3076);
  nand ginst6117 (P1_R1375_U135, P1_R1375_U68, P1_U3074);
  nand ginst6118 (P1_R1375_U136, P1_R1375_U71, P1_U3503);
  nand ginst6119 (P1_R1375_U137, P1_R1375_U72, P1_U3506);
  nand ginst6120 (P1_R1375_U138, P1_R1375_U67, P1_U3079);
  nand ginst6121 (P1_R1375_U139, P1_R1375_U43, P1_U3470);
  and ginst6122 (P1_R1375_U14, P1_R1375_U115, P1_R1375_U204, P1_R1375_U205);
  nand ginst6123 (P1_R1375_U140, P1_R1375_U139, P1_R1375_U90);
  nand ginst6124 (P1_R1375_U141, P1_R1375_U60, P1_U3083);
  nand ginst6125 (P1_R1375_U142, P1_R1375_U59, P1_U3084);
  nand ginst6126 (P1_R1375_U143, P1_R1375_U39, P1_U3071);
  nand ginst6127 (P1_R1375_U144, P1_R1375_U58, P1_U3070);
  nand ginst6128 (P1_R1375_U145, P1_R1375_U57, P1_U3060);
  or ginst6129 (P1_R1375_U146, P1_R1375_U13, P1_U3447);
  nand ginst6130 (P1_R1375_U147, P1_R1375_U47, P1_U3077);
  not ginst6131 (P1_R1375_U148, P1_R1375_U49);
  nand ginst6132 (P1_R1375_U149, P1_R1375_U55, P1_U3064);
  not ginst6133 (P1_R1375_U15, P1_U3983);
  nand ginst6134 (P1_R1375_U150, P1_R1375_U148, P1_U3455);
  nand ginst6135 (P1_R1375_U151, P1_R1375_U150, P1_U3078);
  nand ginst6136 (P1_R1375_U152, P1_R1375_U49, P1_R1375_U50);
  nand ginst6137 (P1_R1375_U153, P1_R1375_U54, P1_U3068);
  nand ginst6138 (P1_R1375_U154, P1_R1375_U151, P1_R1375_U92, P1_R1375_U93);
  nand ginst6139 (P1_R1375_U155, P1_R1375_U149, P1_R1375_U94);
  nand ginst6140 (P1_R1375_U156, P1_R1375_U46, P1_U3461);
  nand ginst6141 (P1_R1375_U157, P1_R1375_U155, P1_R1375_U156);
  nand ginst6142 (P1_R1375_U158, P1_R1375_U145, P1_R1375_U157);
  nand ginst6143 (P1_R1375_U159, P1_R1375_U40, P1_U3467);
  not ginst6144 (P1_R1375_U16, P1_U3984);
  nand ginst6145 (P1_R1375_U160, P1_R1375_U45, P1_U3464);
  nand ginst6146 (P1_R1375_U161, P1_R1375_U43, P1_U3470);
  nand ginst6147 (P1_R1375_U162, P1_R1375_U158, P1_R1375_U95);
  nand ginst6148 (P1_R1375_U163, P1_R1375_U64, P1_U3485);
  nand ginst6149 (P1_R1375_U164, P1_R1375_U63, P1_U3488);
  nand ginst6150 (P1_R1375_U165, P1_R1375_U142, P1_R1375_U96);
  nand ginst6151 (P1_R1375_U166, P1_R1375_U42, P1_U3476);
  nand ginst6152 (P1_R1375_U167, P1_R1375_U165, P1_R1375_U166);
  nand ginst6153 (P1_R1375_U168, P1_R1375_U140, P1_R1375_U162, P1_R1375_U8);
  nand ginst6154 (P1_R1375_U169, P1_R1375_U141, P1_R1375_U167);
  not ginst6155 (P1_R1375_U17, P1_U3056);
  nand ginst6156 (P1_R1375_U170, P1_R1375_U41, P1_U3479);
  nand ginst6157 (P1_R1375_U171, P1_R1375_U62, P1_U3482);
  nand ginst6158 (P1_R1375_U172, P1_R1375_U154, P1_R1375_U168, P1_R1375_U169, P1_R1375_U98);
  nand ginst6159 (P1_R1375_U173, P1_R1375_U9, P1_R1375_U99);
  nand ginst6160 (P1_R1375_U174, P1_R1375_U53, P1_U3072);
  nand ginst6161 (P1_R1375_U175, P1_R1375_U63, P1_U3488);
  nand ginst6162 (P1_R1375_U176, P1_R1375_U100, P1_R1375_U175);
  nand ginst6163 (P1_R1375_U177, P1_R1375_U66, P1_U3080);
  nand ginst6164 (P1_R1375_U178, P1_R1375_U101, P1_R1375_U172);
  nand ginst6165 (P1_R1375_U179, P1_R1375_U65, P1_U3491);
  not ginst6166 (P1_R1375_U18, P1_U3985);
  nand ginst6167 (P1_R1375_U180, P1_R1375_U178, P1_R1375_U179);
  nand ginst6168 (P1_R1375_U181, P1_R1375_U138, P1_R1375_U180);
  nand ginst6169 (P1_R1375_U182, P1_R1375_U38, P1_U3494);
  nand ginst6170 (P1_R1375_U183, P1_R1375_U181, P1_R1375_U182);
  nand ginst6171 (P1_R1375_U184, P1_R1375_U135, P1_R1375_U183);
  nand ginst6172 (P1_R1375_U185, P1_R1375_U37, P1_U3497);
  nand ginst6173 (P1_R1375_U186, P1_R1375_U70, P1_U3500);
  nand ginst6174 (P1_R1375_U187, P1_R1375_U103, P1_R1375_U184);
  nand ginst6175 (P1_R1375_U188, P1_R1375_U105, P1_R1375_U7);
  nand ginst6176 (P1_R1375_U189, P1_R1375_U72, P1_U3506);
  not ginst6177 (P1_R1375_U19, P1_U3059);
  nand ginst6178 (P1_R1375_U190, P1_R1375_U106, P1_R1375_U189);
  nand ginst6179 (P1_R1375_U191, P1_R1375_U36, P1_U3082);
  nand ginst6180 (P1_R1375_U192, P1_R1375_U74, P1_U3081);
  nand ginst6181 (P1_R1375_U193, P1_R1375_U107, P1_R1375_U187);
  nand ginst6182 (P1_R1375_U194, P1_R1375_U73, P1_U3508);
  nand ginst6183 (P1_R1375_U195, P1_R1375_U193, P1_R1375_U194);
  nand ginst6184 (P1_R1375_U196, P1_R1375_U110, P1_R1375_U133);
  nand ginst6185 (P1_R1375_U197, P1_R1375_U33, P1_U3981);
  nand ginst6186 (P1_R1375_U198, P1_R1375_U30, P1_U3980);
  nand ginst6187 (P1_R1375_U199, P1_R1375_U116, P1_U3984);
  not ginst6188 (P1_R1375_U20, P1_U3055);
  nand ginst6189 (P1_R1375_U200, P1_R1375_U116, P1_R1375_U19);
  nand ginst6190 (P1_R1375_U201, P1_R1375_U11, P1_R1375_U202);
  nand ginst6191 (P1_R1375_U202, P1_R1375_U16, P1_U3059);
  nand ginst6192 (P1_R1375_U203, P1_R1375_U114, P1_R1375_U132);
  nand ginst6193 (P1_R1375_U204, P1_R1375_U203, P1_R1375_U89);
  nand ginst6194 (P1_R1375_U205, P1_R1375_U111, P1_R1375_U112, P1_R1375_U126, P1_R1375_U78, P1_R1375_U80);
  nand ginst6195 (P1_R1375_U206, P1_R1375_U22, P1_U3053);
  nand ginst6196 (P1_R1375_U207, P1_R1375_U113, P1_U3975);
  not ginst6197 (P1_R1375_U21, P1_U3054);
  not ginst6198 (P1_R1375_U22, P1_U3975);
  not ginst6199 (P1_R1375_U23, P1_U3057);
  not ginst6200 (P1_R1375_U24, P1_U3977);
  not ginst6201 (P1_R1375_U25, P1_U3974);
  not ginst6202 (P1_R1375_U26, P1_U3976);
  not ginst6203 (P1_R1375_U27, P1_U3978);
  not ginst6204 (P1_R1375_U28, P1_U3066);
  not ginst6205 (P1_R1375_U29, P1_U3979);
  not ginst6206 (P1_R1375_U30, P1_U3061);
  not ginst6207 (P1_R1375_U31, P1_U3058);
  not ginst6208 (P1_R1375_U32, P1_U3065);
  not ginst6209 (P1_R1375_U33, P1_U3075);
  not ginst6210 (P1_R1375_U34, P1_U3076);
  not ginst6211 (P1_R1375_U35, P1_U3503);
  not ginst6212 (P1_R1375_U36, P1_U3506);
  not ginst6213 (P1_R1375_U37, P1_U3074);
  not ginst6214 (P1_R1375_U38, P1_U3079);
  not ginst6215 (P1_R1375_U39, P1_U3470);
  not ginst6216 (P1_R1375_U40, P1_U3067);
  not ginst6217 (P1_R1375_U41, P1_U3083);
  not ginst6218 (P1_R1375_U42, P1_U3084);
  not ginst6219 (P1_R1375_U43, P1_U3071);
  not ginst6220 (P1_R1375_U44, P1_U3070);
  not ginst6221 (P1_R1375_U45, P1_U3060);
  not ginst6222 (P1_R1375_U46, P1_U3064);
  not ginst6223 (P1_R1375_U47, P1_U3450);
  not ginst6224 (P1_R1375_U48, P1_U3077);
  nand ginst6225 (P1_R1375_U49, P1_R1375_U146, P1_R1375_U147);
  not ginst6226 (P1_R1375_U50, P1_U3455);
  not ginst6227 (P1_R1375_U51, P1_U3068);
  not ginst6228 (P1_R1375_U52, P1_U3485);
  not ginst6229 (P1_R1375_U53, P1_U3488);
  not ginst6230 (P1_R1375_U54, P1_U3458);
  not ginst6231 (P1_R1375_U55, P1_U3461);
  not ginst6232 (P1_R1375_U56, P1_U3467);
  not ginst6233 (P1_R1375_U57, P1_U3464);
  not ginst6234 (P1_R1375_U58, P1_U3473);
  not ginst6235 (P1_R1375_U59, P1_U3476);
  and ginst6236 (P1_R1375_U6, P1_R1375_U119, P1_R1375_U120);
  not ginst6237 (P1_R1375_U60, P1_U3479);
  not ginst6238 (P1_R1375_U61, P1_U3482);
  not ginst6239 (P1_R1375_U62, P1_U3062);
  not ginst6240 (P1_R1375_U63, P1_U3072);
  not ginst6241 (P1_R1375_U64, P1_U3063);
  not ginst6242 (P1_R1375_U65, P1_U3080);
  not ginst6243 (P1_R1375_U66, P1_U3491);
  not ginst6244 (P1_R1375_U67, P1_U3494);
  not ginst6245 (P1_R1375_U68, P1_U3497);
  not ginst6246 (P1_R1375_U69, P1_U3500);
  and ginst6247 (P1_R1375_U7, P1_R1375_U136, P1_R1375_U137);
  not ginst6248 (P1_R1375_U70, P1_U3073);
  not ginst6249 (P1_R1375_U71, P1_U3069);
  not ginst6250 (P1_R1375_U72, P1_U3082);
  not ginst6251 (P1_R1375_U73, P1_U3081);
  not ginst6252 (P1_R1375_U74, P1_U3508);
  not ginst6253 (P1_R1375_U75, P1_U3982);
  not ginst6254 (P1_R1375_U76, P1_U3981);
  not ginst6255 (P1_R1375_U77, P1_U3980);
  nand ginst6256 (P1_R1375_U78, P1_R1375_U11, P1_R1375_U125);
  nand ginst6257 (P1_R1375_U79, P1_R1375_U12, P1_R1375_U122, P1_R1375_U124, P1_R1375_U87);
  and ginst6258 (P1_R1375_U8, P1_R1375_U141, P1_R1375_U142, P1_R1375_U143, P1_R1375_U144);
  nand ginst6259 (P1_R1375_U80, P1_R1375_U109, P1_R1375_U195);
  and ginst6260 (P1_R1375_U81, P1_R1375_U113, P1_U3975);
  and ginst6261 (P1_R1375_U82, P1_R1375_U31, P1_U3977);
  and ginst6262 (P1_R1375_U83, P1_R1375_U21, P1_U3974);
  and ginst6263 (P1_R1375_U84, P1_R1375_U23, P1_U3976);
  and ginst6264 (P1_R1375_U85, P1_R1375_U29, P1_U3066);
  and ginst6265 (P1_R1375_U86, P1_R1375_U77, P1_U3061);
  and ginst6266 (P1_R1375_U87, P1_R1375_U121, P1_R1375_U123);
  and ginst6267 (P1_R1375_U88, P1_R1375_U126, P1_R1375_U129);
  and ginst6268 (P1_R1375_U89, P1_R1375_U128, P1_R1375_U131, P1_R1375_U201);
  and ginst6269 (P1_R1375_U9, P1_R1375_U163, P1_R1375_U164);
  and ginst6270 (P1_R1375_U90, P1_R1375_U56, P1_U3067);
  and ginst6271 (P1_R1375_U91, P1_R1375_U145, P1_R1375_U149);
  and ginst6272 (P1_R1375_U92, P1_R1375_U140, P1_R1375_U91);
  and ginst6273 (P1_R1375_U93, P1_R1375_U152, P1_R1375_U153, P1_R1375_U8);
  and ginst6274 (P1_R1375_U94, P1_R1375_U51, P1_U3458);
  and ginst6275 (P1_R1375_U95, P1_R1375_U159, P1_R1375_U160, P1_R1375_U161);
  and ginst6276 (P1_R1375_U96, P1_R1375_U44, P1_U3473);
  and ginst6277 (P1_R1375_U97, P1_R1375_U170, P1_R1375_U171);
  and ginst6278 (P1_R1375_U98, P1_R1375_U9, P1_R1375_U97);
  and ginst6279 (P1_R1375_U99, P1_R1375_U61, P1_U3062);
  and ginst6280 (P1_SUB_84_U10, P1_SUB_84_U195, P1_SUB_84_U221);
  nor ginst6281 (P1_SUB_84_U100, P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN, P1_IR_REG_20__SCAN_IN);
  and ginst6282 (P1_SUB_84_U101, P1_SUB_84_U100, P1_SUB_84_U97, P1_SUB_84_U98, P1_SUB_84_U99);
  nor ginst6283 (P1_SUB_84_U102, P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN);
  nor ginst6284 (P1_SUB_84_U103, P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN, P1_IR_REG_25__SCAN_IN);
  nor ginst6285 (P1_SUB_84_U104, P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN);
  nor ginst6286 (P1_SUB_84_U105, P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN);
  and ginst6287 (P1_SUB_84_U106, P1_SUB_84_U102, P1_SUB_84_U103, P1_SUB_84_U104, P1_SUB_84_U105);
  nor ginst6288 (P1_SUB_84_U107, P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN);
  nor ginst6289 (P1_SUB_84_U108, P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN);
  nor ginst6290 (P1_SUB_84_U109, P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN);
  and ginst6291 (P1_SUB_84_U11, P1_SUB_84_U220, P1_SUB_84_U34);
  nor ginst6292 (P1_SUB_84_U110, P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN, P1_IR_REG_20__SCAN_IN);
  and ginst6293 (P1_SUB_84_U111, P1_SUB_84_U107, P1_SUB_84_U108, P1_SUB_84_U109, P1_SUB_84_U110);
  nor ginst6294 (P1_SUB_84_U112, P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN);
  nor ginst6295 (P1_SUB_84_U113, P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN, P1_IR_REG_24__SCAN_IN);
  nor ginst6296 (P1_SUB_84_U114, P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN);
  nor ginst6297 (P1_SUB_84_U115, P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN);
  and ginst6298 (P1_SUB_84_U116, P1_SUB_84_U112, P1_SUB_84_U113, P1_SUB_84_U114, P1_SUB_84_U115);
  nor ginst6299 (P1_SUB_84_U117, P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN);
  nor ginst6300 (P1_SUB_84_U118, P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN);
  nor ginst6301 (P1_SUB_84_U119, P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN);
  and ginst6302 (P1_SUB_84_U12, P1_SUB_84_U197, P1_SUB_84_U219);
  nor ginst6303 (P1_SUB_84_U120, P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN, P1_IR_REG_19__SCAN_IN);
  and ginst6304 (P1_SUB_84_U121, P1_SUB_84_U117, P1_SUB_84_U118, P1_SUB_84_U119, P1_SUB_84_U120);
  nor ginst6305 (P1_SUB_84_U122, P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN);
  nor ginst6306 (P1_SUB_84_U123, P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN, P1_IR_REG_23__SCAN_IN);
  nor ginst6307 (P1_SUB_84_U124, P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN);
  nor ginst6308 (P1_SUB_84_U125, P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN);
  and ginst6309 (P1_SUB_84_U126, P1_SUB_84_U122, P1_SUB_84_U123, P1_SUB_84_U124, P1_SUB_84_U125);
  nor ginst6310 (P1_SUB_84_U127, P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN);
  nor ginst6311 (P1_SUB_84_U128, P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN, P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN);
  nor ginst6312 (P1_SUB_84_U129, P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN);
  and ginst6313 (P1_SUB_84_U13, P1_SUB_84_U198, P1_SUB_84_U217);
  nor ginst6314 (P1_SUB_84_U130, P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN);
  nor ginst6315 (P1_SUB_84_U131, P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN);
  nor ginst6316 (P1_SUB_84_U132, P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN);
  nor ginst6317 (P1_SUB_84_U133, P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN);
  and ginst6318 (P1_SUB_84_U134, P1_SUB_84_U131, P1_SUB_84_U132, P1_SUB_84_U133);
  nor ginst6319 (P1_SUB_84_U135, P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN);
  nor ginst6320 (P1_SUB_84_U136, P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN);
  and ginst6321 (P1_SUB_84_U137, P1_SUB_84_U135, P1_SUB_84_U136);
  nor ginst6322 (P1_SUB_84_U138, P1_IR_REG_1__SCAN_IN, P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN);
  nor ginst6323 (P1_SUB_84_U139, P1_IR_REG_0__SCAN_IN, P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN);
  and ginst6324 (P1_SUB_84_U14, P1_SUB_84_U172, P1_SUB_84_U216);
  nor ginst6325 (P1_SUB_84_U140, P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN);
  and ginst6326 (P1_SUB_84_U141, P1_SUB_84_U139, P1_SUB_84_U140);
  nor ginst6327 (P1_SUB_84_U142, P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN);
  nor ginst6328 (P1_SUB_84_U143, P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN);
  nor ginst6329 (P1_SUB_84_U144, P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN);
  nor ginst6330 (P1_SUB_84_U145, P1_IR_REG_1__SCAN_IN, P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN);
  nor ginst6331 (P1_SUB_84_U146, P1_IR_REG_0__SCAN_IN, P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN, P1_IR_REG_20__SCAN_IN);
  nor ginst6332 (P1_SUB_84_U147, P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN);
  nor ginst6333 (P1_SUB_84_U148, P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN);
  nor ginst6334 (P1_SUB_84_U149, P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN);
  and ginst6335 (P1_SUB_84_U15, P1_SUB_84_U200, P1_SUB_84_U215);
  nor ginst6336 (P1_SUB_84_U150, P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN);
  nor ginst6337 (P1_SUB_84_U151, P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN);
  nor ginst6338 (P1_SUB_84_U152, P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN);
  nor ginst6339 (P1_SUB_84_U153, P1_IR_REG_1__SCAN_IN, P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN);
  nor ginst6340 (P1_SUB_84_U154, P1_IR_REG_0__SCAN_IN, P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN);
  nor ginst6341 (P1_SUB_84_U155, P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN);
  nor ginst6342 (P1_SUB_84_U156, P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN);
  nor ginst6343 (P1_SUB_84_U157, P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN);
  nor ginst6344 (P1_SUB_84_U158, P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN);
  not ginst6345 (P1_SUB_84_U159, P1_IR_REG_9__SCAN_IN);
  and ginst6346 (P1_SUB_84_U16, P1_SUB_84_U201, P1_SUB_84_U213);
  and ginst6347 (P1_SUB_84_U160, P1_SUB_84_U232, P1_SUB_84_U233);
  not ginst6348 (P1_SUB_84_U161, P1_IR_REG_5__SCAN_IN);
  and ginst6349 (P1_SUB_84_U162, P1_SUB_84_U234, P1_SUB_84_U235);
  not ginst6350 (P1_SUB_84_U163, P1_IR_REG_31__SCAN_IN);
  not ginst6351 (P1_SUB_84_U164, P1_IR_REG_30__SCAN_IN);
  and ginst6352 (P1_SUB_84_U165, P1_SUB_84_U238, P1_SUB_84_U239);
  not ginst6353 (P1_SUB_84_U166, P1_IR_REG_27__SCAN_IN);
  nand ginst6354 (P1_SUB_84_U167, P1_SUB_84_U91, P1_SUB_84_U96);
  not ginst6355 (P1_SUB_84_U168, P1_IR_REG_25__SCAN_IN);
  nand ginst6356 (P1_SUB_84_U169, P1_SUB_84_U111, P1_SUB_84_U116);
  and ginst6357 (P1_SUB_84_U17, P1_SUB_84_U169, P1_SUB_84_U212);
  and ginst6358 (P1_SUB_84_U170, P1_SUB_84_U242, P1_SUB_84_U243);
  not ginst6359 (P1_SUB_84_U171, P1_IR_REG_21__SCAN_IN);
  nand ginst6360 (P1_SUB_84_U172, P1_SUB_84_U143, P1_SUB_84_U144, P1_SUB_84_U145, P1_SUB_84_U146, P1_SUB_84_U147);
  and ginst6361 (P1_SUB_84_U173, P1_SUB_84_U244, P1_SUB_84_U245);
  not ginst6362 (P1_SUB_84_U174, P1_IR_REG_1__SCAN_IN);
  not ginst6363 (P1_SUB_84_U175, P1_IR_REG_0__SCAN_IN);
  not ginst6364 (P1_SUB_84_U176, P1_IR_REG_17__SCAN_IN);
  and ginst6365 (P1_SUB_84_U177, P1_SUB_84_U248, P1_SUB_84_U249);
  not ginst6366 (P1_SUB_84_U178, P1_IR_REG_13__SCAN_IN);
  and ginst6367 (P1_SUB_84_U179, P1_SUB_84_U250, P1_SUB_84_U251);
  and ginst6368 (P1_SUB_84_U18, P1_SUB_84_U167, P1_SUB_84_U211);
  nand ginst6369 (P1_SUB_84_U180, P1_SUB_84_U230, P1_SUB_84_U32);
  not ginst6370 (P1_SUB_84_U181, P1_SUB_84_U29);
  not ginst6371 (P1_SUB_84_U182, P1_SUB_84_U30);
  nand ginst6372 (P1_SUB_84_U183, P1_SUB_84_U182, P1_SUB_84_U31);
  not ginst6373 (P1_SUB_84_U184, P1_SUB_84_U28);
  nand ginst6374 (P1_SUB_84_U185, P1_IR_REG_8__SCAN_IN, P1_SUB_84_U183);
  nand ginst6375 (P1_SUB_84_U186, P1_IR_REG_7__SCAN_IN, P1_SUB_84_U30);
  nand ginst6376 (P1_SUB_84_U187, P1_SUB_84_U161, P1_SUB_84_U181);
  nand ginst6377 (P1_SUB_84_U188, P1_IR_REG_6__SCAN_IN, P1_SUB_84_U187);
  nand ginst6378 (P1_SUB_84_U189, P1_IR_REG_4__SCAN_IN, P1_SUB_84_U180);
  and ginst6379 (P1_SUB_84_U19, P1_SUB_84_U204, P1_SUB_84_U209);
  nand ginst6380 (P1_SUB_84_U190, P1_IR_REG_3__SCAN_IN, P1_SUB_84_U27);
  not ginst6381 (P1_SUB_84_U191, P1_SUB_84_U38);
  nand ginst6382 (P1_SUB_84_U192, P1_SUB_84_U191, P1_SUB_84_U39);
  not ginst6383 (P1_SUB_84_U193, P1_SUB_84_U35);
  not ginst6384 (P1_SUB_84_U194, P1_SUB_84_U36);
  nand ginst6385 (P1_SUB_84_U195, P1_SUB_84_U194, P1_SUB_84_U37);
  not ginst6386 (P1_SUB_84_U196, P1_SUB_84_U34);
  nand ginst6387 (P1_SUB_84_U197, P1_SUB_84_U152, P1_SUB_84_U153, P1_SUB_84_U154, P1_SUB_84_U155);
  nand ginst6388 (P1_SUB_84_U198, P1_SUB_84_U148, P1_SUB_84_U149, P1_SUB_84_U150, P1_SUB_84_U151);
  not ginst6389 (P1_SUB_84_U199, P1_SUB_84_U172);
  and ginst6390 (P1_SUB_84_U20, P1_SUB_84_U208, P1_SUB_84_U33);
  nand ginst6391 (P1_SUB_84_U200, P1_SUB_84_U134, P1_SUB_84_U196);
  nand ginst6392 (P1_SUB_84_U201, P1_SUB_84_U121, P1_SUB_84_U126);
  not ginst6393 (P1_SUB_84_U202, P1_SUB_84_U169);
  not ginst6394 (P1_SUB_84_U203, P1_SUB_84_U167);
  nand ginst6395 (P1_SUB_84_U204, P1_SUB_84_U61, P1_SUB_84_U66);
  not ginst6396 (P1_SUB_84_U205, P1_SUB_84_U33);
  or ginst6397 (P1_SUB_84_U206, P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN);
  nand ginst6398 (P1_SUB_84_U207, P1_IR_REG_2__SCAN_IN, P1_SUB_84_U206);
  nand ginst6399 (P1_SUB_84_U208, P1_IR_REG_29__SCAN_IN, P1_SUB_84_U204);
  nand ginst6400 (P1_SUB_84_U209, P1_IR_REG_28__SCAN_IN, P1_SUB_84_U229);
  and ginst6401 (P1_SUB_84_U21, P1_SUB_84_U207, P1_SUB_84_U27);
  nand ginst6402 (P1_SUB_84_U210, P1_SUB_84_U101, P1_SUB_84_U106);
  nand ginst6403 (P1_SUB_84_U211, P1_IR_REG_26__SCAN_IN, P1_SUB_84_U210);
  nand ginst6404 (P1_SUB_84_U212, P1_IR_REG_24__SCAN_IN, P1_SUB_84_U201);
  nand ginst6405 (P1_SUB_84_U213, P1_IR_REG_23__SCAN_IN, P1_SUB_84_U200);
  nand ginst6406 (P1_SUB_84_U214, P1_SUB_84_U137, P1_SUB_84_U138, P1_SUB_84_U141, P1_SUB_84_U142);
  nand ginst6407 (P1_SUB_84_U215, P1_IR_REG_22__SCAN_IN, P1_SUB_84_U214);
  nand ginst6408 (P1_SUB_84_U216, P1_IR_REG_20__SCAN_IN, P1_SUB_84_U198);
  nand ginst6409 (P1_SUB_84_U217, P1_IR_REG_19__SCAN_IN, P1_SUB_84_U197);
  nand ginst6410 (P1_SUB_84_U218, P1_SUB_84_U176, P1_SUB_84_U196);
  nand ginst6411 (P1_SUB_84_U219, P1_IR_REG_18__SCAN_IN, P1_SUB_84_U218);
  and ginst6412 (P1_SUB_84_U22, P1_SUB_84_U180, P1_SUB_84_U190);
  nand ginst6413 (P1_SUB_84_U220, P1_IR_REG_16__SCAN_IN, P1_SUB_84_U195);
  nand ginst6414 (P1_SUB_84_U221, P1_IR_REG_15__SCAN_IN, P1_SUB_84_U36);
  nand ginst6415 (P1_SUB_84_U222, P1_SUB_84_U178, P1_SUB_84_U193);
  nand ginst6416 (P1_SUB_84_U223, P1_IR_REG_14__SCAN_IN, P1_SUB_84_U222);
  nand ginst6417 (P1_SUB_84_U224, P1_IR_REG_12__SCAN_IN, P1_SUB_84_U192);
  nand ginst6418 (P1_SUB_84_U225, P1_IR_REG_11__SCAN_IN, P1_SUB_84_U38);
  nand ginst6419 (P1_SUB_84_U226, P1_SUB_84_U159, P1_SUB_84_U184);
  nand ginst6420 (P1_SUB_84_U227, P1_IR_REG_10__SCAN_IN, P1_SUB_84_U226);
  nand ginst6421 (P1_SUB_84_U228, P1_SUB_84_U164, P1_SUB_84_U205);
  nand ginst6422 (P1_SUB_84_U229, P1_SUB_84_U71, P1_SUB_84_U76);
  and ginst6423 (P1_SUB_84_U23, P1_SUB_84_U189, P1_SUB_84_U29);
  not ginst6424 (P1_SUB_84_U230, P1_SUB_84_U27);
  nand ginst6425 (P1_SUB_84_U231, P1_SUB_84_U81, P1_SUB_84_U86);
  nand ginst6426 (P1_SUB_84_U232, P1_IR_REG_9__SCAN_IN, P1_SUB_84_U28);
  nand ginst6427 (P1_SUB_84_U233, P1_SUB_84_U159, P1_SUB_84_U184);
  nand ginst6428 (P1_SUB_84_U234, P1_IR_REG_5__SCAN_IN, P1_SUB_84_U29);
  nand ginst6429 (P1_SUB_84_U235, P1_SUB_84_U161, P1_SUB_84_U181);
  nand ginst6430 (P1_SUB_84_U236, P1_SUB_84_U163, P1_SUB_84_U228);
  nand ginst6431 (P1_SUB_84_U237, P1_IR_REG_31__SCAN_IN, P1_SUB_84_U164, P1_SUB_84_U205);
  nand ginst6432 (P1_SUB_84_U238, P1_IR_REG_30__SCAN_IN, P1_SUB_84_U33);
  nand ginst6433 (P1_SUB_84_U239, P1_SUB_84_U164, P1_SUB_84_U205);
  and ginst6434 (P1_SUB_84_U24, P1_SUB_84_U188, P1_SUB_84_U30);
  nand ginst6435 (P1_SUB_84_U240, P1_IR_REG_27__SCAN_IN, P1_SUB_84_U203);
  nand ginst6436 (P1_SUB_84_U241, P1_SUB_84_U166, P1_SUB_84_U231);
  nand ginst6437 (P1_SUB_84_U242, P1_IR_REG_25__SCAN_IN, P1_SUB_84_U169);
  nand ginst6438 (P1_SUB_84_U243, P1_SUB_84_U168, P1_SUB_84_U202);
  nand ginst6439 (P1_SUB_84_U244, P1_IR_REG_21__SCAN_IN, P1_SUB_84_U172);
  nand ginst6440 (P1_SUB_84_U245, P1_SUB_84_U171, P1_SUB_84_U199);
  nand ginst6441 (P1_SUB_84_U246, P1_IR_REG_1__SCAN_IN, P1_SUB_84_U175);
  nand ginst6442 (P1_SUB_84_U247, P1_IR_REG_0__SCAN_IN, P1_SUB_84_U174);
  nand ginst6443 (P1_SUB_84_U248, P1_IR_REG_17__SCAN_IN, P1_SUB_84_U34);
  nand ginst6444 (P1_SUB_84_U249, P1_SUB_84_U176, P1_SUB_84_U196);
  and ginst6445 (P1_SUB_84_U25, P1_SUB_84_U183, P1_SUB_84_U186);
  nand ginst6446 (P1_SUB_84_U250, P1_IR_REG_13__SCAN_IN, P1_SUB_84_U35);
  nand ginst6447 (P1_SUB_84_U251, P1_SUB_84_U178, P1_SUB_84_U193);
  and ginst6448 (P1_SUB_84_U26, P1_SUB_84_U185, P1_SUB_84_U28);
  or ginst6449 (P1_SUB_84_U27, P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN);
  nand ginst6450 (P1_SUB_84_U28, P1_SUB_84_U230, P1_SUB_84_U43, P1_SUB_84_U44);
  nand ginst6451 (P1_SUB_84_U29, P1_SUB_84_U230, P1_SUB_84_U45);
  nand ginst6452 (P1_SUB_84_U30, P1_SUB_84_U181, P1_SUB_84_U46);
  not ginst6453 (P1_SUB_84_U31, P1_IR_REG_7__SCAN_IN);
  not ginst6454 (P1_SUB_84_U32, P1_IR_REG_3__SCAN_IN);
  nand ginst6455 (P1_SUB_84_U33, P1_SUB_84_U51, P1_SUB_84_U56);
  nand ginst6456 (P1_SUB_84_U34, P1_SUB_84_U127, P1_SUB_84_U128, P1_SUB_84_U129, P1_SUB_84_U130);
  nand ginst6457 (P1_SUB_84_U35, P1_SUB_84_U156, P1_SUB_84_U184);
  nand ginst6458 (P1_SUB_84_U36, P1_SUB_84_U157, P1_SUB_84_U193);
  not ginst6459 (P1_SUB_84_U37, P1_IR_REG_15__SCAN_IN);
  nand ginst6460 (P1_SUB_84_U38, P1_SUB_84_U158, P1_SUB_84_U184);
  not ginst6461 (P1_SUB_84_U39, P1_IR_REG_11__SCAN_IN);
  nand ginst6462 (P1_SUB_84_U40, P1_SUB_84_U246, P1_SUB_84_U247);
  nand ginst6463 (P1_SUB_84_U41, P1_SUB_84_U236, P1_SUB_84_U237);
  nand ginst6464 (P1_SUB_84_U42, P1_SUB_84_U240, P1_SUB_84_U241);
  nor ginst6465 (P1_SUB_84_U43, P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN);
  nor ginst6466 (P1_SUB_84_U44, P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN);
  nor ginst6467 (P1_SUB_84_U45, P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN);
  nor ginst6468 (P1_SUB_84_U46, P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN);
  nor ginst6469 (P1_SUB_84_U47, P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN);
  nor ginst6470 (P1_SUB_84_U48, P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN);
  nor ginst6471 (P1_SUB_84_U49, P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN, P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN);
  nor ginst6472 (P1_SUB_84_U50, P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN);
  and ginst6473 (P1_SUB_84_U51, P1_SUB_84_U47, P1_SUB_84_U48, P1_SUB_84_U49, P1_SUB_84_U50);
  nor ginst6474 (P1_SUB_84_U52, P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN);
  nor ginst6475 (P1_SUB_84_U53, P1_IR_REG_2__SCAN_IN, P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN);
  nor ginst6476 (P1_SUB_84_U54, P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN);
  nor ginst6477 (P1_SUB_84_U55, P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN);
  and ginst6478 (P1_SUB_84_U56, P1_SUB_84_U52, P1_SUB_84_U53, P1_SUB_84_U54, P1_SUB_84_U55);
  nor ginst6479 (P1_SUB_84_U57, P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN);
  nor ginst6480 (P1_SUB_84_U58, P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN);
  nor ginst6481 (P1_SUB_84_U59, P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN, P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN);
  and ginst6482 (P1_SUB_84_U6, P1_SUB_84_U227, P1_SUB_84_U38);
  nor ginst6483 (P1_SUB_84_U60, P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN);
  and ginst6484 (P1_SUB_84_U61, P1_SUB_84_U57, P1_SUB_84_U58, P1_SUB_84_U59, P1_SUB_84_U60);
  nor ginst6485 (P1_SUB_84_U62, P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN);
  nor ginst6486 (P1_SUB_84_U63, P1_IR_REG_2__SCAN_IN, P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN);
  nor ginst6487 (P1_SUB_84_U64, P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN);
  nor ginst6488 (P1_SUB_84_U65, P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN);
  and ginst6489 (P1_SUB_84_U66, P1_SUB_84_U62, P1_SUB_84_U63, P1_SUB_84_U64, P1_SUB_84_U65);
  nor ginst6490 (P1_SUB_84_U67, P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN);
  nor ginst6491 (P1_SUB_84_U68, P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN);
  nor ginst6492 (P1_SUB_84_U69, P1_IR_REG_1__SCAN_IN, P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN);
  and ginst6493 (P1_SUB_84_U7, P1_SUB_84_U192, P1_SUB_84_U225);
  nor ginst6494 (P1_SUB_84_U70, P1_IR_REG_0__SCAN_IN, P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN);
  and ginst6495 (P1_SUB_84_U71, P1_SUB_84_U67, P1_SUB_84_U68, P1_SUB_84_U69, P1_SUB_84_U70);
  nor ginst6496 (P1_SUB_84_U72, P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN);
  nor ginst6497 (P1_SUB_84_U73, P1_IR_REG_2__SCAN_IN, P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN);
  nor ginst6498 (P1_SUB_84_U74, P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN);
  nor ginst6499 (P1_SUB_84_U75, P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN);
  and ginst6500 (P1_SUB_84_U76, P1_SUB_84_U72, P1_SUB_84_U73, P1_SUB_84_U74, P1_SUB_84_U75);
  nor ginst6501 (P1_SUB_84_U77, P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN);
  nor ginst6502 (P1_SUB_84_U78, P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN);
  nor ginst6503 (P1_SUB_84_U79, P1_IR_REG_1__SCAN_IN, P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN);
  and ginst6504 (P1_SUB_84_U8, P1_SUB_84_U224, P1_SUB_84_U35);
  nor ginst6505 (P1_SUB_84_U80, P1_IR_REG_0__SCAN_IN, P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN);
  and ginst6506 (P1_SUB_84_U81, P1_SUB_84_U77, P1_SUB_84_U78, P1_SUB_84_U79, P1_SUB_84_U80);
  nor ginst6507 (P1_SUB_84_U82, P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN);
  nor ginst6508 (P1_SUB_84_U83, P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN, P1_IR_REG_26__SCAN_IN);
  nor ginst6509 (P1_SUB_84_U84, P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN);
  nor ginst6510 (P1_SUB_84_U85, P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN);
  and ginst6511 (P1_SUB_84_U86, P1_SUB_84_U82, P1_SUB_84_U83, P1_SUB_84_U84, P1_SUB_84_U85);
  nor ginst6512 (P1_SUB_84_U87, P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN);
  nor ginst6513 (P1_SUB_84_U88, P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN);
  nor ginst6514 (P1_SUB_84_U89, P1_IR_REG_1__SCAN_IN, P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN);
  and ginst6515 (P1_SUB_84_U9, P1_SUB_84_U223, P1_SUB_84_U36);
  nor ginst6516 (P1_SUB_84_U90, P1_IR_REG_0__SCAN_IN, P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN);
  and ginst6517 (P1_SUB_84_U91, P1_SUB_84_U87, P1_SUB_84_U88, P1_SUB_84_U89, P1_SUB_84_U90);
  nor ginst6518 (P1_SUB_84_U92, P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN);
  nor ginst6519 (P1_SUB_84_U93, P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN, P1_IR_REG_26__SCAN_IN);
  nor ginst6520 (P1_SUB_84_U94, P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN);
  nor ginst6521 (P1_SUB_84_U95, P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN);
  and ginst6522 (P1_SUB_84_U96, P1_SUB_84_U92, P1_SUB_84_U93, P1_SUB_84_U94, P1_SUB_84_U95);
  nor ginst6523 (P1_SUB_84_U97, P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN);
  nor ginst6524 (P1_SUB_84_U98, P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN);
  nor ginst6525 (P1_SUB_84_U99, P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN);
  and ginst6526 (P1_U3014, P1_U3443, P1_U3956);
  and ginst6527 (P1_U3015, P1_U3446, P1_U3449);
  and ginst6528 (P1_U3016, P1_U3625, P1_U3630);
  and ginst6529 (P1_U3017, P1_U3444, P1_U3445);
  and ginst6530 (P1_U3018, P1_U3444, P1_U5711);
  and ginst6531 (P1_U3019, P1_U3445, P1_U5708);
  and ginst6532 (P1_U3020, P1_U5708, P1_U5711);
  and ginst6533 (P1_U3021, P1_U3421, P1_U5368);
  and ginst6534 (P1_U3022, P1_STATE_REG_SCAN_IN, P1_U3046);
  and ginst6535 (P1_U3023, P1_U3049, P1_U5690);
  and ginst6536 (P1_U3024, P1_U3423, P1_U3807);
  and ginst6537 (P1_U3025, P1_U3987, P1_U5699);
  and ginst6538 (P1_U3026, P1_U3953, P1_U5690);
  and ginst6539 (P1_U3027, P1_U3871, P1_U3972);
  and ginst6540 (P1_U3028, P1_STATE_REG_SCAN_IN, P1_U3357);
  and ginst6541 (P1_U3029, P1_U3964, P1_U3989);
  and ginst6542 (P1_U3030, P1_U3422, P1_U3989);
  and ginst6543 (P1_U3031, P1_U3957, P1_U3989);
  and ginst6544 (P1_U3032, P1_U3965, P1_U3989);
  and ginst6545 (P1_U3033, P1_U3446, P1_U3987);
  and ginst6546 (P1_U3034, P1_U3972, P1_U5699);
  and ginst6547 (P1_U3035, P1_U3025, P1_U3989);
  and ginst6548 (P1_U3036, P1_U3446, P1_U3972);
  and ginst6549 (P1_U3037, P1_U4880, P1_U5702);
  and ginst6550 (P1_U3038, P1_U3024, P1_U5702);
  and ginst6551 (P1_U3039, P1_U4880, P1_U5699);
  and ginst6552 (P1_U3040, P1_U3024, P1_U5699);
  and ginst6553 (P1_U3041, P1_U3015, P1_U4880);
  and ginst6554 (P1_U3042, P1_U3015, P1_U3024);
  and ginst6555 (P1_U3043, P1_U3022, P1_U3423);
  and ginst6556 (P1_U3044, P1_STATE_REG_SCAN_IN, P1_U5113);
  and ginst6557 (P1_U3045, P1_U3022, P1_U5115);
  and ginst6558 (P1_U3046, P1_U3421, P1_U5677);
  and ginst6559 (P1_U3047, P1_U3016, P1_U3631);
  and ginst6560 (P1_U3048, P1_U3442, P1_U5690);
  and ginst6561 (P1_U3049, P1_U5684, P1_U5693);
  and ginst6562 (P1_U3050, P1_U3435, P1_U3437);
  and ginst6563 (P1_U3051, P1_U4699, P1_U4700, P1_U4703, P1_U4706);
  and ginst6564 (P1_U3052, P1_U6069, P1_U6070);
  nand ginst6565 (P1_U3053, P1_U4636, P1_U4637, P1_U4638, P1_U4639);
  nand ginst6566 (P1_U3054, P1_U4655, P1_U4656, P1_U4657, P1_U4658);
  nand ginst6567 (P1_U3055, P1_U4674, P1_U4675, P1_U4676, P1_U4677);
  nand ginst6568 (P1_U3056, P1_U4713, P1_U4714, P1_U4715);
  nand ginst6569 (P1_U3057, P1_U4617, P1_U4618, P1_U4619, P1_U4620);
  nand ginst6570 (P1_U3058, P1_U4598, P1_U4599, P1_U4600, P1_U4601);
  nand ginst6571 (P1_U3059, P1_U4693, P1_U4694, P1_U4695);
  nand ginst6572 (P1_U3060, P1_U4199, P1_U4200, P1_U4201, P1_U4202);
  nand ginst6573 (P1_U3061, P1_U4541, P1_U4542, P1_U4543, P1_U4544);
  nand ginst6574 (P1_U3062, P1_U4313, P1_U4314, P1_U4315, P1_U4316);
  nand ginst6575 (P1_U3063, P1_U4332, P1_U4333, P1_U4334, P1_U4335);
  nand ginst6576 (P1_U3064, P1_U4180, P1_U4181, P1_U4182, P1_U4183);
  nand ginst6577 (P1_U3065, P1_U4579, P1_U4580, P1_U4581, P1_U4582);
  nand ginst6578 (P1_U3066, P1_U4560, P1_U4561, P1_U4562, P1_U4563);
  nand ginst6579 (P1_U3067, P1_U4218, P1_U4219, P1_U4220, P1_U4221);
  nand ginst6580 (P1_U3068, P1_U4156, P1_U4157, P1_U4158, P1_U4159);
  nand ginst6581 (P1_U3069, P1_U4446, P1_U4447, P1_U4448, P1_U4449);
  nand ginst6582 (P1_U3070, P1_U4256, P1_U4257, P1_U4258, P1_U4259);
  nand ginst6583 (P1_U3071, P1_U4237, P1_U4238, P1_U4239, P1_U4240);
  nand ginst6584 (P1_U3072, P1_U4351, P1_U4352, P1_U4353, P1_U4354);
  nand ginst6585 (P1_U3073, P1_U4427, P1_U4428, P1_U4429, P1_U4430);
  nand ginst6586 (P1_U3074, P1_U4408, P1_U4409, P1_U4410, P1_U4411);
  nand ginst6587 (P1_U3075, P1_U4522, P1_U4523, P1_U4524, P1_U4525);
  nand ginst6588 (P1_U3076, P1_U4503, P1_U4504, P1_U4505, P1_U4506);
  nand ginst6589 (P1_U3077, P1_U4161, P1_U4162, P1_U4163, P1_U4164);
  nand ginst6590 (P1_U3078, P1_U4137, P1_U4138, P1_U4139, P1_U4140);
  nand ginst6591 (P1_U3079, P1_U4389, P1_U4390, P1_U4391, P1_U4392);
  nand ginst6592 (P1_U3080, P1_U4370, P1_U4371, P1_U4372, P1_U4373);
  nand ginst6593 (P1_U3081, P1_U4484, P1_U4485, P1_U4486, P1_U4487);
  nand ginst6594 (P1_U3082, P1_U4465, P1_U4466, P1_U4467, P1_U4468);
  nand ginst6595 (P1_U3083, P1_U4294, P1_U4295, P1_U4296, P1_U4297);
  nand ginst6596 (P1_U3084, P1_U4275, P1_U4276, P1_U4277, P1_U4278);
  nand ginst6597 (P1_U3085, P1_STATE_REG_SCAN_IN, P1_U4887);
  not ginst6598 (P1_U3086, P1_STATE_REG_SCAN_IN);
  nand ginst6599 (P1_U3087, P1_U5575, P1_U5576);
  nand ginst6600 (P1_U3088, P1_U5577, P1_U5578);
  nand ginst6601 (P1_U3089, P1_U5582, P1_U5583, P1_U5584);
  nand ginst6602 (P1_U3090, P1_U3895, P1_U5586);
  nand ginst6603 (P1_U3091, P1_U3896, P1_U5589);
  nand ginst6604 (P1_U3092, P1_U3897, P1_U5592);
  nand ginst6605 (P1_U3093, P1_U3898, P1_U5595);
  nand ginst6606 (P1_U3094, P1_U3899, P1_U5598);
  nand ginst6607 (P1_U3095, P1_U3900, P1_U5601);
  nand ginst6608 (P1_U3096, P1_U3901, P1_U5604);
  nand ginst6609 (P1_U3097, P1_U3902, P1_U5607);
  nand ginst6610 (P1_U3098, P1_U3903, P1_U5610);
  nand ginst6611 (P1_U3099, P1_U3904, P1_U5616);
  nand ginst6612 (P1_U3100, P1_U3905, P1_U5619);
  nand ginst6613 (P1_U3101, P1_U3906, P1_U5622);
  nand ginst6614 (P1_U3102, P1_U3907, P1_U5625);
  nand ginst6615 (P1_U3103, P1_U3908, P1_U5628);
  nand ginst6616 (P1_U3104, P1_U3909, P1_U5631);
  nand ginst6617 (P1_U3105, P1_U5633, P1_U5634, P1_U5635);
  nand ginst6618 (P1_U3106, P1_U5636, P1_U5637, P1_U5638);
  nand ginst6619 (P1_U3107, P1_U5639, P1_U5640, P1_U5641);
  nand ginst6620 (P1_U3108, P1_U5642, P1_U5643, P1_U5644);
  nand ginst6621 (P1_U3109, P1_U5557, P1_U5558, P1_U5559);
  nand ginst6622 (P1_U3110, P1_U5560, P1_U5561, P1_U5562);
  nand ginst6623 (P1_U3111, P1_U5563, P1_U5564, P1_U5565);
  nand ginst6624 (P1_U3112, P1_U5566, P1_U5567, P1_U5568);
  nand ginst6625 (P1_U3113, P1_U5569, P1_U5570, P1_U5571);
  nand ginst6626 (P1_U3114, P1_U5572, P1_U5573, P1_U5574);
  nand ginst6627 (P1_U3115, P1_U5579, P1_U5580, P1_U5581);
  nand ginst6628 (P1_U3116, P1_U5612, P1_U5613, P1_U5614);
  nand ginst6629 (P1_U3117, P1_U5645, P1_U5646, P1_U5647);
  nand ginst6630 (P1_U3118, P1_U5648, P1_U5649);
  nand ginst6631 (P1_U3119, P1_U5505, P1_U5506);
  nand ginst6632 (P1_U3120, P1_U5507, P1_U5508);
  nand ginst6633 (P1_U3121, P1_U3438, P1_U5511, P1_U5512);
  nand ginst6634 (P1_U3122, P1_U3879, P1_U5513);
  nand ginst6635 (P1_U3123, P1_U3880, P1_U5515);
  nand ginst6636 (P1_U3124, P1_U3881, P1_U5517);
  nand ginst6637 (P1_U3125, P1_U3882, P1_U5519);
  nand ginst6638 (P1_U3126, P1_U3883, P1_U5521);
  nand ginst6639 (P1_U3127, P1_U3884, P1_U5523);
  nand ginst6640 (P1_U3128, P1_U3885, P1_U5525);
  nand ginst6641 (P1_U3129, P1_U3886, P1_U5527);
  nand ginst6642 (P1_U3130, P1_U3887, P1_U5529);
  nand ginst6643 (P1_U3131, P1_U3888, P1_U5534);
  nand ginst6644 (P1_U3132, P1_U3889, P1_U5536);
  nand ginst6645 (P1_U3133, P1_U3890, P1_U5538);
  nand ginst6646 (P1_U3134, P1_U3891, P1_U5540);
  nand ginst6647 (P1_U3135, P1_U3892, P1_U5542);
  nand ginst6648 (P1_U3136, P1_U3893, P1_U5544);
  nand ginst6649 (P1_U3137, P1_U3438, P1_U5545, P1_U5546);
  nand ginst6650 (P1_U3138, P1_U3438, P1_U5547, P1_U5548);
  nand ginst6651 (P1_U3139, P1_U3438, P1_U5549, P1_U5550);
  nand ginst6652 (P1_U3140, P1_U3438, P1_U5551, P1_U5552);
  nand ginst6653 (P1_U3141, P1_U3438, P1_U5493, P1_U5494);
  nand ginst6654 (P1_U3142, P1_U3438, P1_U5495, P1_U5496);
  nand ginst6655 (P1_U3143, P1_U3438, P1_U5497, P1_U5498);
  nand ginst6656 (P1_U3144, P1_U3438, P1_U5499, P1_U5500);
  nand ginst6657 (P1_U3145, P1_U3438, P1_U5501, P1_U5502);
  nand ginst6658 (P1_U3146, P1_U3438, P1_U5503, P1_U5504);
  nand ginst6659 (P1_U3147, P1_U3438, P1_U5509, P1_U5510);
  nand ginst6660 (P1_U3148, P1_U3438, P1_U5531, P1_U5532);
  nand ginst6661 (P1_U3149, P1_U3438, P1_U5553, P1_U5554);
  nand ginst6662 (P1_U3150, P1_U3894, P1_U5556);
  nand ginst6663 (P1_U3151, P1_U3438, P1_U3953);
  nand ginst6664 (P1_U3152, P1_U3372, P1_U5677);
  nand ginst6665 (P1_U3153, P1_U5447, P1_U5448);
  nand ginst6666 (P1_U3154, P1_U5449, P1_U5450);
  nand ginst6667 (P1_U3155, P1_U5451, P1_U5452);
  nand ginst6668 (P1_U3156, P1_U5453, P1_U5454);
  nand ginst6669 (P1_U3157, P1_U5455, P1_U5456);
  nand ginst6670 (P1_U3158, P1_U5457, P1_U5458);
  nand ginst6671 (P1_U3159, P1_U5459, P1_U5460);
  nand ginst6672 (P1_U3160, P1_U5461, P1_U5462);
  nand ginst6673 (P1_U3161, P1_U5463, P1_U5464);
  nand ginst6674 (P1_U3162, P1_U5467, P1_U5468);
  nand ginst6675 (P1_U3163, P1_U5469, P1_U5470);
  nand ginst6676 (P1_U3164, P1_U5471, P1_U5472);
  nand ginst6677 (P1_U3165, P1_U5473, P1_U5474);
  nand ginst6678 (P1_U3166, P1_U5475, P1_U5476);
  nand ginst6679 (P1_U3167, P1_U5477, P1_U5478);
  nand ginst6680 (P1_U3168, P1_U5479, P1_U5480);
  nand ginst6681 (P1_U3169, P1_U5481, P1_U5482);
  nand ginst6682 (P1_U3170, P1_U5483, P1_U5484);
  nand ginst6683 (P1_U3171, P1_U5485, P1_U5486);
  nand ginst6684 (P1_U3172, P1_U5433, P1_U5434);
  nand ginst6685 (P1_U3173, P1_U5435, P1_U5436);
  nand ginst6686 (P1_U3174, P1_U5437, P1_U5438);
  nand ginst6687 (P1_U3175, P1_U5439, P1_U5440);
  nand ginst6688 (P1_U3176, P1_U5441, P1_U5442);
  nand ginst6689 (P1_U3177, P1_U5443, P1_U5444);
  nand ginst6690 (P1_U3178, P1_U5445, P1_U5446);
  nand ginst6691 (P1_U3179, P1_U5465, P1_U5466);
  nand ginst6692 (P1_U3180, P1_U5487, P1_U5488);
  nand ginst6693 (P1_U3181, P1_U5489, P1_U5490, P1_U5491);
  nand ginst6694 (P1_U3182, P1_U5388, P1_U5389);
  nand ginst6695 (P1_U3183, P1_U5390, P1_U5391);
  nand ginst6696 (P1_U3184, P1_U5392, P1_U5393);
  nand ginst6697 (P1_U3185, P1_U5394, P1_U5395);
  nand ginst6698 (P1_U3186, P1_U5396, P1_U5397);
  nand ginst6699 (P1_U3187, P1_U5398, P1_U5399);
  nand ginst6700 (P1_U3188, P1_U5400, P1_U5401);
  nand ginst6701 (P1_U3189, P1_U5402, P1_U5403);
  nand ginst6702 (P1_U3190, P1_U5404, P1_U5405);
  nand ginst6703 (P1_U3191, P1_U5408, P1_U5409);
  nand ginst6704 (P1_U3192, P1_U5410, P1_U5411);
  nand ginst6705 (P1_U3193, P1_U5412, P1_U5413);
  nand ginst6706 (P1_U3194, P1_U5414, P1_U5415);
  nand ginst6707 (P1_U3195, P1_U5416, P1_U5417);
  nand ginst6708 (P1_U3196, P1_U5418, P1_U5419);
  nand ginst6709 (P1_U3197, P1_U5420, P1_U5421);
  nand ginst6710 (P1_U3198, P1_U5422, P1_U5423);
  nand ginst6711 (P1_U3199, P1_U5424, P1_U5425);
  nand ginst6712 (P1_U3200, P1_U5426, P1_U5427);
  nand ginst6713 (P1_U3201, P1_U5374, P1_U5375);
  nand ginst6714 (P1_U3202, P1_U5376, P1_U5377);
  nand ginst6715 (P1_U3203, P1_U5378, P1_U5379);
  nand ginst6716 (P1_U3204, P1_U5380, P1_U5381);
  nand ginst6717 (P1_U3205, P1_U5382, P1_U5383);
  nand ginst6718 (P1_U3206, P1_U5384, P1_U5385);
  nand ginst6719 (P1_U3207, P1_U5386, P1_U5387);
  nand ginst6720 (P1_U3208, P1_U5406, P1_U5407);
  nand ginst6721 (P1_U3209, P1_U5428, P1_U5429);
  nand ginst6722 (P1_U3210, P1_U3878, P1_U5430);
  and ginst6723 (P1_U3211, P1_U3421, P1_U5367);
  nand ginst6724 (P1_U3212, P1_U5365, P1_U6235, P1_U6236);
  nand ginst6725 (P1_U3213, P1_U5358, P1_U5359, P1_U5360, P1_U5361, P1_U5362);
  nand ginst6726 (P1_U3214, P1_U5349, P1_U5350, P1_U5351, P1_U5352, P1_U5353);
  nand ginst6727 (P1_U3215, P1_U5340, P1_U5341, P1_U5342, P1_U5343, P1_U5344);
  nand ginst6728 (P1_U3216, P1_U5331, P1_U5332, P1_U5333, P1_U5334, P1_U5335);
  nand ginst6729 (P1_U3217, P1_U5322, P1_U5323, P1_U5324, P1_U5325, P1_U5326);
  nand ginst6730 (P1_U3218, P1_U5313, P1_U5314, P1_U5315, P1_U5316, P1_U5317);
  nand ginst6731 (P1_U3219, P1_U5304, P1_U5305, P1_U5306, P1_U5307, P1_U5308);
  nand ginst6732 (P1_U3220, P1_U5295, P1_U5296, P1_U5297, P1_U5298, P1_U5299);
  nand ginst6733 (P1_U3221, P1_U5286, P1_U5287, P1_U5288, P1_U5289, P1_U5290);
  nand ginst6734 (P1_U3222, P1_U3876, P1_U5277, P1_U5278, P1_U5279);
  nand ginst6735 (P1_U3223, P1_U5268, P1_U5269, P1_U5270, P1_U5271, P1_U5272);
  nand ginst6736 (P1_U3224, P1_U5259, P1_U5260, P1_U5261, P1_U5262, P1_U5263);
  nand ginst6737 (P1_U3225, P1_U5250, P1_U5251, P1_U5252, P1_U5253, P1_U5254);
  nand ginst6738 (P1_U3226, P1_U5241, P1_U5242, P1_U5243, P1_U5244, P1_U5245);
  nand ginst6739 (P1_U3227, P1_U5232, P1_U5233, P1_U5234, P1_U5235, P1_U5236);
  nand ginst6740 (P1_U3228, P1_U5223, P1_U5224, P1_U5225, P1_U5226, P1_U5227);
  nand ginst6741 (P1_U3229, P1_U5214, P1_U5215, P1_U5216, P1_U5217, P1_U5218);
  nand ginst6742 (P1_U3230, P1_U5205, P1_U5206, P1_U5207, P1_U5208, P1_U5209);
  nand ginst6743 (P1_U3231, P1_U5196, P1_U5197, P1_U5198, P1_U5199, P1_U5200);
  nand ginst6744 (P1_U3232, P1_U3874, P1_U3875, P1_U5189);
  nand ginst6745 (P1_U3233, P1_U5179, P1_U5180, P1_U5181, P1_U5182, P1_U5183);
  nand ginst6746 (P1_U3234, P1_U5170, P1_U5171, P1_U5172, P1_U5173, P1_U5174);
  nand ginst6747 (P1_U3235, P1_U5161, P1_U5162, P1_U5163, P1_U5164, P1_U5165);
  nand ginst6748 (P1_U3236, P1_U5152, P1_U5153, P1_U5154, P1_U5155, P1_U5156);
  nand ginst6749 (P1_U3237, P1_U3872, P1_U5143, P1_U5144, P1_U5145);
  nand ginst6750 (P1_U3238, P1_U5134, P1_U5135, P1_U5136, P1_U5137, P1_U5138);
  nand ginst6751 (P1_U3239, P1_U5125, P1_U5126, P1_U5127, P1_U5128, P1_U5129);
  nand ginst6752 (P1_U3240, P1_U5116, P1_U5117, P1_U5118, P1_U5119, P1_U5120);
  nand ginst6753 (P1_U3241, P1_U5103, P1_U5104, P1_U5105, P1_U5106, P1_U5107);
  and ginst6754 (P1_U3242, P1_U3866, P1_U5650);
  nand ginst6755 (P1_U3243, P1_U3848, P1_U3849);
  nand ginst6756 (P1_U3244, P1_U3846, P1_U3847);
  nand ginst6757 (P1_U3245, P1_U3844, P1_U3845);
  nand ginst6758 (P1_U3246, P1_U3841, P1_U3842);
  nand ginst6759 (P1_U3247, P1_U3839, P1_U3840);
  nand ginst6760 (P1_U3248, P1_U3836, P1_U3837);
  nand ginst6761 (P1_U3249, P1_U3834, P1_U3835);
  nand ginst6762 (P1_U3250, P1_U3832, P1_U3833, P1_U5010);
  nand ginst6763 (P1_U3251, P1_U3830, P1_U3831, P1_U5000);
  nand ginst6764 (P1_U3252, P1_U3828, P1_U3829, P1_U4990);
  nand ginst6765 (P1_U3253, P1_U3826, P1_U3827, P1_U4980);
  nand ginst6766 (P1_U3254, P1_U3824, P1_U3825, P1_U4970);
  nand ginst6767 (P1_U3255, P1_U3822, P1_U3823, P1_U4960);
  nand ginst6768 (P1_U3256, P1_U3820, P1_U3821, P1_U4950);
  nand ginst6769 (P1_U3257, P1_U3818, P1_U3819, P1_U4940);
  nand ginst6770 (P1_U3258, P1_U3816, P1_U3817, P1_U4930);
  nand ginst6771 (P1_U3259, P1_U3814, P1_U3815, P1_U4920);
  nand ginst6772 (P1_U3260, P1_U3812, P1_U3813, P1_U4910);
  nand ginst6773 (P1_U3261, P1_U3810, P1_U3811, P1_U4900);
  nand ginst6774 (P1_U3262, P1_U3808, P1_U3809, P1_U4890);
  nand ginst6775 (P1_U3263, P1_U3947, P1_U4878, P1_U4879);
  nand ginst6776 (P1_U3264, P1_U3946, P1_U4876, P1_U4877);
  nand ginst6777 (P1_U3265, P1_U3799, P1_U3800, P1_U3943, P1_U4869);
  nand ginst6778 (P1_U3266, P1_U3797, P1_U3798, P1_U3942, P1_U4864);
  nand ginst6779 (P1_U3267, P1_U3795, P1_U3796, P1_U3941, P1_U4859);
  nand ginst6780 (P1_U3268, P1_U3793, P1_U3794, P1_U3940, P1_U4854);
  nand ginst6781 (P1_U3269, P1_U3791, P1_U3792, P1_U3939, P1_U4849);
  nand ginst6782 (P1_U3270, P1_U3789, P1_U3790, P1_U3938);
  nand ginst6783 (P1_U3271, P1_U3787, P1_U3788, P1_U3937);
  nand ginst6784 (P1_U3272, P1_U3786, P1_U3936);
  nand ginst6785 (P1_U3273, P1_U3784, P1_U3785, P1_U3935);
  nand ginst6786 (P1_U3274, P1_U3783, P1_U3934);
  nand ginst6787 (P1_U3275, P1_U3782, P1_U3933);
  nand ginst6788 (P1_U3276, P1_U3781, P1_U3932);
  nand ginst6789 (P1_U3277, P1_U3780, P1_U3931);
  nand ginst6790 (P1_U3278, P1_U3779, P1_U3930);
  xor ginst6791 (P1_U3279, P1_U3279_in, flip_signal);
  nand ginst6792 (P1_U3279_in, P1_U3778, P1_U3929);
  nand ginst6793 (P1_U3280, P1_U3776, P1_U3777, P1_U3928);
  nand ginst6794 (P1_U3281, P1_U3774, P1_U3775, P1_U3927);
  nand ginst6795 (P1_U3282, P1_U3772, P1_U3773, P1_U3926);
  nand ginst6796 (P1_U3283, P1_U3770, P1_U3771, P1_U3925, P1_U4779);
  nand ginst6797 (P1_U3284, P1_U3768, P1_U3769, P1_U3924, P1_U4774);
  nand ginst6798 (P1_U3285, P1_U3766, P1_U3767, P1_U3923, P1_U4769);
  nand ginst6799 (P1_U3286, P1_U3764, P1_U3765, P1_U3922, P1_U4764);
  nand ginst6800 (P1_U3287, P1_U3762, P1_U3763, P1_U3921, P1_U4759);
  nand ginst6801 (P1_U3288, P1_U3760, P1_U3761, P1_U3920, P1_U4754);
  nand ginst6802 (P1_U3289, P1_U3758, P1_U3759, P1_U3919, P1_U4749);
  nand ginst6803 (P1_U3290, P1_U3756, P1_U3757, P1_U3918);
  nand ginst6804 (P1_U3291, P1_U3754, P1_U3755);
  nand ginst6805 (P1_U3292, P1_U3752, P1_U3753);
  nand ginst6806 (P1_U3293, P1_U3750, P1_U3751);
  and ginst6807 (P1_U3294, P1_D_REG_31__SCAN_IN, P1_U3911);
  and ginst6808 (P1_U3295, P1_D_REG_30__SCAN_IN, P1_U3911);
  and ginst6809 (P1_U3296, P1_D_REG_29__SCAN_IN, P1_U3911);
  and ginst6810 (P1_U3297, P1_D_REG_28__SCAN_IN, P1_U3911);
  and ginst6811 (P1_U3298, P1_D_REG_27__SCAN_IN, P1_U3911);
  and ginst6812 (P1_U3299, P1_D_REG_26__SCAN_IN, P1_U3911);
  and ginst6813 (P1_U3300, P1_D_REG_25__SCAN_IN, P1_U3911);
  and ginst6814 (P1_U3301, P1_D_REG_24__SCAN_IN, P1_U3911);
  and ginst6815 (P1_U3302, P1_D_REG_23__SCAN_IN, P1_U3911);
  and ginst6816 (P1_U3303, P1_D_REG_22__SCAN_IN, P1_U3911);
  and ginst6817 (P1_U3304, P1_D_REG_21__SCAN_IN, P1_U3911);
  and ginst6818 (P1_U3305, P1_D_REG_20__SCAN_IN, P1_U3911);
  and ginst6819 (P1_U3306, P1_D_REG_19__SCAN_IN, P1_U3911);
  and ginst6820 (P1_U3307, P1_D_REG_18__SCAN_IN, P1_U3911);
  and ginst6821 (P1_U3308, P1_D_REG_17__SCAN_IN, P1_U3911);
  and ginst6822 (P1_U3309, P1_D_REG_16__SCAN_IN, P1_U3911);
  and ginst6823 (P1_U3310, P1_D_REG_15__SCAN_IN, P1_U3911);
  and ginst6824 (P1_U3311, P1_D_REG_14__SCAN_IN, P1_U3911);
  and ginst6825 (P1_U3312, P1_D_REG_13__SCAN_IN, P1_U3911);
  and ginst6826 (P1_U3313, P1_D_REG_12__SCAN_IN, P1_U3911);
  and ginst6827 (P1_U3314, P1_D_REG_11__SCAN_IN, P1_U3911);
  and ginst6828 (P1_U3315, P1_D_REG_10__SCAN_IN, P1_U3911);
  and ginst6829 (P1_U3316, P1_D_REG_9__SCAN_IN, P1_U3911);
  and ginst6830 (P1_U3317, P1_D_REG_8__SCAN_IN, P1_U3911);
  and ginst6831 (P1_U3318, P1_D_REG_7__SCAN_IN, P1_U3911);
  and ginst6832 (P1_U3319, P1_D_REG_6__SCAN_IN, P1_U3911);
  and ginst6833 (P1_U3320, P1_D_REG_5__SCAN_IN, P1_U3911);
  and ginst6834 (P1_U3321, P1_D_REG_4__SCAN_IN, P1_U3911);
  and ginst6835 (P1_U3322, P1_D_REG_3__SCAN_IN, P1_U3911);
  and ginst6836 (P1_U3323, P1_D_REG_2__SCAN_IN, P1_U3911);
  nand ginst6837 (P1_U3324, P1_U4098, P1_U4099, P1_U4100);
  nand ginst6838 (P1_U3325, P1_U4095, P1_U4096, P1_U4097);
  nand ginst6839 (P1_U3326, P1_U4092, P1_U4093, P1_U4094);
  nand ginst6840 (P1_U3327, P1_U4089, P1_U4090, P1_U4091);
  nand ginst6841 (P1_U3328, P1_U4086, P1_U4087, P1_U4088);
  nand ginst6842 (P1_U3329, P1_U4083, P1_U4084, P1_U4085);
  nand ginst6843 (P1_U3330, P1_U4080, P1_U4081, P1_U4082);
  nand ginst6844 (P1_U3331, P1_U4077, P1_U4078, P1_U4079);
  nand ginst6845 (P1_U3332, P1_U4074, P1_U4075, P1_U4076);
  nand ginst6846 (P1_U3333, P1_U4071, P1_U4072, P1_U4073);
  nand ginst6847 (P1_U3334, P1_U4068, P1_U4069, P1_U4070);
  nand ginst6848 (P1_U3335, P1_U4065, P1_U4066, P1_U4067);
  nand ginst6849 (P1_U3336, P1_U4062, P1_U4063, P1_U4064);
  nand ginst6850 (P1_U3337, P1_U4059, P1_U4060, P1_U4061);
  nand ginst6851 (P1_U3338, P1_U4056, P1_U4057, P1_U4058);
  nand ginst6852 (P1_U3339, P1_U4053, P1_U4054, P1_U4055);
  nand ginst6853 (P1_U3340, P1_U4050, P1_U4051, P1_U4052);
  nand ginst6854 (P1_U3341, P1_U4047, P1_U4048, P1_U4049);
  nand ginst6855 (P1_U3342, P1_U4044, P1_U4045, P1_U4046);
  nand ginst6856 (P1_U3343, P1_U4041, P1_U4042, P1_U4043);
  nand ginst6857 (P1_U3344, P1_U4038, P1_U4039, P1_U4040);
  nand ginst6858 (P1_U3345, P1_U4035, P1_U4036, P1_U4037);
  nand ginst6859 (P1_U3346, P1_U4032, P1_U4033, P1_U4034);
  nand ginst6860 (P1_U3347, P1_U4029, P1_U4030, P1_U4031);
  nand ginst6861 (P1_U3348, P1_U4026, P1_U4027, P1_U4028);
  nand ginst6862 (P1_U3349, P1_U4023, P1_U4024, P1_U4025);
  nand ginst6863 (P1_U3350, P1_U4020, P1_U4021, P1_U4022);
  nand ginst6864 (P1_U3351, P1_U4017, P1_U4018, P1_U4019);
  nand ginst6865 (P1_U3352, P1_U4014, P1_U4015, P1_U4016);
  nand ginst6866 (P1_U3353, P1_U4011, P1_U4012, P1_U4013);
  nand ginst6867 (P1_U3354, P1_U4008, P1_U4009, P1_U4010);
  nand ginst6868 (P1_U3355, P1_U4005, P1_U4006, P1_U4007);
  nand ginst6869 (P1_U3356, P1_U3944, P1_U4872, P1_U4873, P1_U4874, P1_U4875);
  nand ginst6870 (P1_U3357, P1_STATE_REG_SCAN_IN, P1_U3910);
  nand ginst6871 (P1_U3358, P1_U3437, P1_U5669);
  not ginst6872 (P1_U3359, P1_B_REG_SCAN_IN);
  nand ginst6873 (P1_U3360, P1_U3437, P1_U5673, P1_U5674);
  nand ginst6874 (P1_U3361, P1_U3048, P1_U3443);
  nand ginst6875 (P1_U3362, P1_U3441, P1_U3442, P1_U3443);
  nand ginst6876 (P1_U3363, P1_U3441, P1_U5687);
  nand ginst6877 (P1_U3364, P1_U3443, P1_U4001);
  nand ginst6878 (P1_U3365, P1_U3441, P1_U3442, P1_U3447);
  nand ginst6879 (P1_U3366, P1_U3447, P1_U4001);
  nand ginst6880 (P1_U3367, P1_U5687, P1_U5690);
  nand ginst6881 (P1_U3368, P1_U3443, P1_U4002);
  nand ginst6882 (P1_U3369, P1_U3960, P1_U5693);
  nand ginst6883 (P1_U3370, P1_U3447, P1_U4002);
  nand ginst6884 (P1_U3371, P1_U3956, P1_U5684);
  nand ginst6885 (P1_U3372, P1_U3442, P1_U5684);
  nand ginst6886 (P1_U3373, P1_U3443, P1_U3447);
  nand ginst6887 (P1_U3374, P1_U3618, P1_U3619, P1_U4147, P1_U4148, P1_U4149);
  not ginst6888 (P1_U3375, P1_REG2_REG_0__SCAN_IN);
  nand ginst6889 (P1_U3376, P1_U3633, P1_U3635, P1_U4166, P1_U4167);
  nand ginst6890 (P1_U3377, P1_U3637, P1_U3639, P1_U4185, P1_U4186);
  nand ginst6891 (P1_U3378, P1_U3642, P1_U4204, P1_U4205, P1_U4206, P1_U4207);
  nand ginst6892 (P1_U3379, P1_U3645, P1_U4223, P1_U4224, P1_U4225, P1_U4226);
  nand ginst6893 (P1_U3380, P1_U3647, P1_U3649, P1_U4242, P1_U4243);
  nand ginst6894 (P1_U3381, P1_U3651, P1_U3653, P1_U4261, P1_U4262);
  nand ginst6895 (P1_U3382, P1_U3655, P1_U3657, P1_U4280, P1_U4281);
  nand ginst6896 (P1_U3383, P1_U3659, P1_U3661, P1_U4299, P1_U4300);
  nand ginst6897 (P1_U3384, P1_U3663, P1_U3665, P1_U4318, P1_U4319);
  nand ginst6898 (P1_U3385, P1_U3667, P1_U3669, P1_U4337, P1_U4338);
  nand ginst6899 (P1_U3386, P1_U3671, P1_U3673, P1_U4356, P1_U4357);
  nand ginst6900 (P1_U3387, P1_U3675, P1_U3677, P1_U4375, P1_U4376);
  nand ginst6901 (P1_U3388, P1_U3679, P1_U3681, P1_U4394, P1_U4395);
  nand ginst6902 (P1_U3389, P1_U3683, P1_U3685, P1_U4413, P1_U4414);
  nand ginst6903 (P1_U3390, P1_U3687, P1_U3689, P1_U4432, P1_U4433);
  nand ginst6904 (P1_U3391, P1_U3691, P1_U3693, P1_U4451, P1_U4452);
  nand ginst6905 (P1_U3392, P1_U3695, P1_U3697, P1_U4470, P1_U4471);
  nand ginst6906 (P1_U3393, P1_U3699, P1_U3701, P1_U4489, P1_U4490);
  nand ginst6907 (P1_U3394, P1_U3703, P1_U3705, P1_U4508, P1_U4509);
  nand ginst6908 (P1_U3395, P1_U3912, U76);
  nand ginst6909 (P1_U3396, P1_U3707, P1_U3709, P1_U4527, P1_U4528);
  nand ginst6910 (P1_U3397, P1_U3912, U75);
  nand ginst6911 (P1_U3398, P1_U3711, P1_U3713, P1_U4546, P1_U4547);
  nand ginst6912 (P1_U3399, P1_U3912, U74);
  nand ginst6913 (P1_U3400, P1_U3715, P1_U3717, P1_U4565, P1_U4566);
  nand ginst6914 (P1_U3401, P1_U3912, U73);
  nand ginst6915 (P1_U3402, P1_U3719, P1_U3721, P1_U4584, P1_U4585);
  nand ginst6916 (P1_U3403, P1_U3912, U72);
  nand ginst6917 (P1_U3404, P1_U3723, P1_U3725, P1_U4603, P1_U4604);
  nand ginst6918 (P1_U3405, P1_U3912, U71);
  nand ginst6919 (P1_U3406, P1_U3727, P1_U3729, P1_U4622, P1_U4623);
  nand ginst6920 (P1_U3407, P1_U3912, U70);
  nand ginst6921 (P1_U3408, P1_U3731, P1_U3733, P1_U4641, P1_U4642);
  nand ginst6922 (P1_U3409, P1_U3912, U69);
  nand ginst6923 (P1_U3410, P1_U3735, P1_U3737, P1_U4660, P1_U4661);
  nand ginst6924 (P1_U3411, P1_U3912, U68);
  nand ginst6925 (P1_U3412, P1_U3739, P1_U3741, P1_U4679, P1_U4680);
  nand ginst6926 (P1_U3413, P1_U3912, U67);
  nand ginst6927 (P1_U3414, P1_U3912, U65);
  nand ginst6928 (P1_U3415, P1_U3912, U64);
  nand ginst6929 (P1_U3416, P1_U3953, P1_U5693);
  nand ginst6930 (P1_U3417, P1_U3022, P1_U4724);
  nand ginst6931 (P1_U3418, P1_U3988, P1_U5690);
  nand ginst6932 (P1_U3419, P1_U3048, P1_U3447);
  nand ginst6933 (P1_U3420, P1_U3023, P1_U5687);
  nand ginst6934 (P1_U3421, P1_U3050, P1_U3436);
  nand ginst6935 (P1_U3422, P1_U3966, P1_U4725);
  nand ginst6936 (P1_U3423, P1_U3424, P1_U4888);
  nand ginst6937 (P1_U3424, P1_U4102, P1_U5677);
  nand ginst6938 (P1_U3425, P1_STATE_REG_SCAN_IN, P1_U3999);
  nand ginst6939 (P1_U3426, P1_U3438, P1_U5687);
  nand ginst6940 (P1_U3427, P1_U3014, P1_U3015);
  nand ginst6941 (P1_U3428, P1_U3438, P1_U3443);
  nand ginst6942 (P1_U3429, P1_U3022, P1_U3422);
  nand ginst6943 (P1_U3430, P1_U3016, P1_U3867);
  nand ginst6944 (P1_U3431, P1_U3014, P1_U3022);
  nand ginst6945 (P1_U3432, P1_U3870, P1_U5101);
  nand ginst6946 (P1_U3433, P1_U3442, P1_U5693);
  nand ginst6947 (P1_U3434, P1_U5370, P1_U5371);
  nand ginst6948 (P1_U3435, P1_U5664, P1_U5665);
  nand ginst6949 (P1_U3436, P1_U5667, P1_U5668);
  nand ginst6950 (P1_U3437, P1_U5670, P1_U5671);
  nand ginst6951 (P1_U3438, P1_U5675, P1_U5676);
  nand ginst6952 (P1_U3439, P1_U5678, P1_U5679);
  nand ginst6953 (P1_U3440, P1_U5680, P1_U5681);
  nand ginst6954 (P1_U3441, P1_U5688, P1_U5689);
  nand ginst6955 (P1_U3442, P1_U5685, P1_U5686);
  nand ginst6956 (P1_U3443, P1_U5682, P1_U5683);
  nand ginst6957 (P1_U3444, P1_U5706, P1_U5707);
  nand ginst6958 (P1_U3445, P1_U5709, P1_U5710);
  nand ginst6959 (P1_U3446, P1_U5697, P1_U5698);
  nand ginst6960 (P1_U3447, P1_U5691, P1_U5692);
  nand ginst6961 (P1_U3448, P1_U5694, P1_U5695);
  nand ginst6962 (P1_U3449, P1_U5700, P1_U5701);
  nand ginst6963 (P1_U3450, P1_U5703, P1_U5704);
  nand ginst6964 (P1_U3451, P1_U5717, P1_U5718);
  nand ginst6965 (P1_U3452, P1_U5714, P1_U5715);
  nand ginst6966 (P1_U3453, P1_U5720, P1_U5721);
  nand ginst6967 (P1_U3454, P1_U5722, P1_U5723);
  nand ginst6968 (P1_U3455, P1_U5724, P1_U5725);
  nand ginst6969 (P1_U3456, P1_U5727, P1_U5728);
  nand ginst6970 (P1_U3457, P1_U5729, P1_U5730);
  nand ginst6971 (P1_U3458, P1_U5731, P1_U5732);
  nand ginst6972 (P1_U3459, P1_U5734, P1_U5735);
  nand ginst6973 (P1_U3460, P1_U5736, P1_U5737);
  nand ginst6974 (P1_U3461, P1_U5738, P1_U5739);
  nand ginst6975 (P1_U3462, P1_U5741, P1_U5742);
  nand ginst6976 (P1_U3463, P1_U5743, P1_U5744);
  nand ginst6977 (P1_U3464, P1_U5745, P1_U5746);
  nand ginst6978 (P1_U3465, P1_U5748, P1_U5749);
  nand ginst6979 (P1_U3466, P1_U5750, P1_U5751);
  nand ginst6980 (P1_U3467, P1_U5752, P1_U5753);
  nand ginst6981 (P1_U3468, P1_U5755, P1_U5756);
  nand ginst6982 (P1_U3469, P1_U5757, P1_U5758);
  nand ginst6983 (P1_U3470, P1_U5759, P1_U5760);
  nand ginst6984 (P1_U3471, P1_U5762, P1_U5763);
  nand ginst6985 (P1_U3472, P1_U5764, P1_U5765);
  nand ginst6986 (P1_U3473, P1_U5766, P1_U5767);
  nand ginst6987 (P1_U3474, P1_U5769, P1_U5770);
  nand ginst6988 (P1_U3475, P1_U5771, P1_U5772);
  nand ginst6989 (P1_U3476, P1_U5773, P1_U5774);
  nand ginst6990 (P1_U3477, P1_U5776, P1_U5777);
  nand ginst6991 (P1_U3478, P1_U5778, P1_U5779);
  nand ginst6992 (P1_U3479, P1_U5780, P1_U5781);
  nand ginst6993 (P1_U3480, P1_U5783, P1_U5784);
  nand ginst6994 (P1_U3481, P1_U5785, P1_U5786);
  nand ginst6995 (P1_U3482, P1_U5787, P1_U5788);
  nand ginst6996 (P1_U3483, P1_U5790, P1_U5791);
  nand ginst6997 (P1_U3484, P1_U5792, P1_U5793);
  nand ginst6998 (P1_U3485, P1_U5794, P1_U5795);
  nand ginst6999 (P1_U3486, P1_U5797, P1_U5798);
  nand ginst7000 (P1_U3487, P1_U5799, P1_U5800);
  nand ginst7001 (P1_U3488, P1_U5801, P1_U5802);
  nand ginst7002 (P1_U3489, P1_U5804, P1_U5805);
  nand ginst7003 (P1_U3490, P1_U5806, P1_U5807);
  nand ginst7004 (P1_U3491, P1_U5808, P1_U5809);
  nand ginst7005 (P1_U3492, P1_U5811, P1_U5812);
  nand ginst7006 (P1_U3493, P1_U5813, P1_U5814);
  nand ginst7007 (P1_U3494, P1_U5815, P1_U5816);
  nand ginst7008 (P1_U3495, P1_U5818, P1_U5819);
  nand ginst7009 (P1_U3496, P1_U5820, P1_U5821);
  nand ginst7010 (P1_U3497, P1_U5822, P1_U5823);
  nand ginst7011 (P1_U3498, P1_U5825, P1_U5826);
  nand ginst7012 (P1_U3499, P1_U5827, P1_U5828);
  nand ginst7013 (P1_U3500, P1_U5829, P1_U5830);
  nand ginst7014 (P1_U3501, P1_U5832, P1_U5833);
  nand ginst7015 (P1_U3502, P1_U5834, P1_U5835);
  nand ginst7016 (P1_U3503, P1_U5836, P1_U5837);
  nand ginst7017 (P1_U3504, P1_U5839, P1_U5840);
  nand ginst7018 (P1_U3505, P1_U5841, P1_U5842);
  nand ginst7019 (P1_U3506, P1_U5843, P1_U5844);
  nand ginst7020 (P1_U3507, P1_U5846, P1_U5847);
  nand ginst7021 (P1_U3508, P1_U5848, P1_U5849);
  nand ginst7022 (P1_U3509, P1_U5851, P1_U5852);
  nand ginst7023 (P1_U3510, P1_U5853, P1_U5854);
  nand ginst7024 (P1_U3511, P1_U5855, P1_U5856);
  nand ginst7025 (P1_U3512, P1_U5857, P1_U5858);
  nand ginst7026 (P1_U3513, P1_U5859, P1_U5860);
  nand ginst7027 (P1_U3514, P1_U5861, P1_U5862);
  nand ginst7028 (P1_U3515, P1_U5863, P1_U5864);
  nand ginst7029 (P1_U3516, P1_U5865, P1_U5866);
  nand ginst7030 (P1_U3517, P1_U5867, P1_U5868);
  nand ginst7031 (P1_U3518, P1_U5869, P1_U5870);
  nand ginst7032 (P1_U3519, P1_U5871, P1_U5872);
  nand ginst7033 (P1_U3520, P1_U5873, P1_U5874);
  nand ginst7034 (P1_U3521, P1_U5875, P1_U5876);
  nand ginst7035 (P1_U3522, P1_U5877, P1_U5878);
  nand ginst7036 (P1_U3523, P1_U5879, P1_U5880);
  nand ginst7037 (P1_U3524, P1_U5881, P1_U5882);
  nand ginst7038 (P1_U3525, P1_U5883, P1_U5884);
  nand ginst7039 (P1_U3526, P1_U5885, P1_U5886);
  nand ginst7040 (P1_U3527, P1_U5887, P1_U5888);
  nand ginst7041 (P1_U3528, P1_U5889, P1_U5890);
  nand ginst7042 (P1_U3529, P1_U5891, P1_U5892);
  nand ginst7043 (P1_U3530, P1_U5893, P1_U5894);
  nand ginst7044 (P1_U3531, P1_U5895, P1_U5896);
  nand ginst7045 (P1_U3532, P1_U5897, P1_U5898);
  nand ginst7046 (P1_U3533, P1_U5899, P1_U5900);
  nand ginst7047 (P1_U3534, P1_U5901, P1_U5902);
  nand ginst7048 (P1_U3535, P1_U5903, P1_U5904);
  nand ginst7049 (P1_U3536, P1_U5905, P1_U5906);
  nand ginst7050 (P1_U3537, P1_U5907, P1_U5908);
  nand ginst7051 (P1_U3538, P1_U5909, P1_U5910);
  nand ginst7052 (P1_U3539, P1_U5911, P1_U5912);
  nand ginst7053 (P1_U3540, P1_U5913, P1_U5914);
  nand ginst7054 (P1_U3541, P1_U5915, P1_U5916);
  nand ginst7055 (P1_U3542, P1_U5917, P1_U5918);
  nand ginst7056 (P1_U3543, P1_U5919, P1_U5920);
  nand ginst7057 (P1_U3544, P1_U5921, P1_U5922);
  nand ginst7058 (P1_U3545, P1_U5923, P1_U5924);
  nand ginst7059 (P1_U3546, P1_U5925, P1_U5926);
  nand ginst7060 (P1_U3547, P1_U5927, P1_U5928);
  nand ginst7061 (P1_U3548, P1_U5929, P1_U5930);
  nand ginst7062 (P1_U3549, P1_U5931, P1_U5932);
  nand ginst7063 (P1_U3550, P1_U5933, P1_U5934);
  nand ginst7064 (P1_U3551, P1_U5935, P1_U5936);
  nand ginst7065 (P1_U3552, P1_U5937, P1_U5938);
  nand ginst7066 (P1_U3553, P1_U5939, P1_U5940);
  nand ginst7067 (P1_U3554, P1_U6005, P1_U6006);
  nand ginst7068 (P1_U3555, P1_U6007, P1_U6008);
  nand ginst7069 (P1_U3556, P1_U6009, P1_U6010);
  nand ginst7070 (P1_U3557, P1_U6011, P1_U6012);
  nand ginst7071 (P1_U3558, P1_U6013, P1_U6014);
  nand ginst7072 (P1_U3559, P1_U6015, P1_U6016);
  nand ginst7073 (P1_U3560, P1_U6017, P1_U6018);
  nand ginst7074 (P1_U3561, P1_U6019, P1_U6020);
  nand ginst7075 (P1_U3562, P1_U6021, P1_U6022);
  nand ginst7076 (P1_U3563, P1_U6023, P1_U6024);
  nand ginst7077 (P1_U3564, P1_U6025, P1_U6026);
  nand ginst7078 (P1_U3565, P1_U6027, P1_U6028);
  nand ginst7079 (P1_U3566, P1_U6029, P1_U6030);
  nand ginst7080 (P1_U3567, P1_U6031, P1_U6032);
  nand ginst7081 (P1_U3568, P1_U6033, P1_U6034);
  nand ginst7082 (P1_U3569, P1_U6035, P1_U6036);
  nand ginst7083 (P1_U3570, P1_U6037, P1_U6038);
  nand ginst7084 (P1_U3571, P1_U6039, P1_U6040);
  nand ginst7085 (P1_U3572, P1_U6041, P1_U6042);
  nand ginst7086 (P1_U3573, P1_U6043, P1_U6044);
  nand ginst7087 (P1_U3574, P1_U6045, P1_U6046);
  nand ginst7088 (P1_U3575, P1_U6047, P1_U6048);
  nand ginst7089 (P1_U3576, P1_U6049, P1_U6050);
  nand ginst7090 (P1_U3577, P1_U6051, P1_U6052);
  nand ginst7091 (P1_U3578, P1_U6053, P1_U6054);
  nand ginst7092 (P1_U3579, P1_U6055, P1_U6056);
  nand ginst7093 (P1_U3580, P1_U6057, P1_U6058);
  nand ginst7094 (P1_U3581, P1_U6059, P1_U6060);
  nand ginst7095 (P1_U3582, P1_U6061, P1_U6062);
  nand ginst7096 (P1_U3583, P1_U6063, P1_U6064);
  nand ginst7097 (P1_U3584, P1_U6065, P1_U6066);
  nand ginst7098 (P1_U3585, P1_U6067, P1_U6068);
  nand ginst7099 (P1_U3586, P1_U6171, P1_U6172);
  nand ginst7100 (P1_U3587, P1_U6173, P1_U6174);
  nand ginst7101 (P1_U3588, P1_U6175, P1_U6176);
  nand ginst7102 (P1_U3589, P1_U6177, P1_U6178);
  nand ginst7103 (P1_U3590, P1_U6179, P1_U6180);
  nand ginst7104 (P1_U3591, P1_U6181, P1_U6182);
  nand ginst7105 (P1_U3592, P1_U6183, P1_U6184);
  nand ginst7106 (P1_U3593, P1_U6185, P1_U6186);
  nand ginst7107 (P1_U3594, P1_U6187, P1_U6188);
  nand ginst7108 (P1_U3595, P1_U6189, P1_U6190);
  nand ginst7109 (P1_U3596, P1_U6191, P1_U6192);
  nand ginst7110 (P1_U3597, P1_U6193, P1_U6194);
  nand ginst7111 (P1_U3598, P1_U6195, P1_U6196);
  nand ginst7112 (P1_U3599, P1_U6197, P1_U6198);
  nand ginst7113 (P1_U3600, P1_U6199, P1_U6200);
  nand ginst7114 (P1_U3601, P1_U6201, P1_U6202);
  nand ginst7115 (P1_U3602, P1_U6203, P1_U6204);
  nand ginst7116 (P1_U3603, P1_U6205, P1_U6206);
  nand ginst7117 (P1_U3604, P1_U6207, P1_U6208);
  nand ginst7118 (P1_U3605, P1_U6209, P1_U6210);
  nand ginst7119 (P1_U3606, P1_U6211, P1_U6212);
  nand ginst7120 (P1_U3607, P1_U6213, P1_U6214);
  nand ginst7121 (P1_U3608, P1_U6215, P1_U6216);
  nand ginst7122 (P1_U3609, P1_U6217, P1_U6218);
  nand ginst7123 (P1_U3610, P1_U6219, P1_U6220);
  nand ginst7124 (P1_U3611, P1_U6221, P1_U6222);
  nand ginst7125 (P1_U3612, P1_U6223, P1_U6224);
  nand ginst7126 (P1_U3613, P1_U6225, P1_U6226);
  nand ginst7127 (P1_U3614, P1_U6227, P1_U6228);
  nand ginst7128 (P1_U3615, P1_U6229, P1_U6230);
  nand ginst7129 (P1_U3616, P1_U6231, P1_U6232);
  nand ginst7130 (P1_U3617, P1_U6233, P1_U6234);
  and ginst7131 (P1_U3618, P1_U4143, P1_U4144);
  and ginst7132 (P1_U3619, P1_U4145, P1_U4146);
  and ginst7133 (P1_U3620, P1_U4151, P1_U4152, P1_U4153, P1_U4154);
  and ginst7134 (P1_U3621, P1_U4105, P1_U4106, P1_U4107, P1_U4108);
  and ginst7135 (P1_U3622, P1_U4109, P1_U4110, P1_U4111, P1_U4112);
  and ginst7136 (P1_U3623, P1_U4113, P1_U4114, P1_U4115, P1_U4116);
  and ginst7137 (P1_U3624, P1_U4117, P1_U4118, P1_U4119);
  and ginst7138 (P1_U3625, P1_U3621, P1_U3622, P1_U3623, P1_U3624);
  and ginst7139 (P1_U3626, P1_U4120, P1_U4121, P1_U4122, P1_U4123);
  and ginst7140 (P1_U3627, P1_U4124, P1_U4125, P1_U4126, P1_U4127);
  and ginst7141 (P1_U3628, P1_U4128, P1_U4129, P1_U4130, P1_U4131);
  and ginst7142 (P1_U3629, P1_U4132, P1_U4133, P1_U4134);
  and ginst7143 (P1_U3630, P1_U3626, P1_U3627, P1_U3628, P1_U3629);
  and ginst7144 (P1_U3631, P1_U4136, P1_U5716);
  and ginst7145 (P1_U3632, P1_U3022, P1_U5719);
  and ginst7146 (P1_U3633, P1_U4168, P1_U4169);
  and ginst7147 (P1_U3634, P1_U4170, P1_U4171);
  and ginst7148 (P1_U3635, P1_U3634, P1_U4172, P1_U4173);
  and ginst7149 (P1_U3636, P1_U4175, P1_U4176, P1_U4177, P1_U4178);
  and ginst7150 (P1_U3637, P1_U4187, P1_U4188);
  and ginst7151 (P1_U3638, P1_U4189, P1_U4190);
  and ginst7152 (P1_U3639, P1_U3638, P1_U4191, P1_U4192);
  and ginst7153 (P1_U3640, P1_U4194, P1_U4195, P1_U4196, P1_U4197);
  and ginst7154 (P1_U3641, P1_U4208, P1_U4209);
  and ginst7155 (P1_U3642, P1_U3641, P1_U4210, P1_U4211);
  and ginst7156 (P1_U3643, P1_U4213, P1_U4214, P1_U4215, P1_U4216);
  and ginst7157 (P1_U3644, P1_U4227, P1_U4228);
  and ginst7158 (P1_U3645, P1_U3644, P1_U4229, P1_U4230);
  and ginst7159 (P1_U3646, P1_U4232, P1_U4233, P1_U4234, P1_U4235);
  and ginst7160 (P1_U3647, P1_U4244, P1_U4245);
  and ginst7161 (P1_U3648, P1_U4246, P1_U4247);
  and ginst7162 (P1_U3649, P1_U3648, P1_U4248, P1_U4249);
  and ginst7163 (P1_U3650, P1_U4251, P1_U4252, P1_U4253, P1_U4254);
  and ginst7164 (P1_U3651, P1_U4263, P1_U4264);
  and ginst7165 (P1_U3652, P1_U4265, P1_U4266);
  and ginst7166 (P1_U3653, P1_U3652, P1_U4267, P1_U4268);
  and ginst7167 (P1_U3654, P1_U4270, P1_U4271, P1_U4272, P1_U4273);
  and ginst7168 (P1_U3655, P1_U4282, P1_U4283);
  and ginst7169 (P1_U3656, P1_U4284, P1_U4285);
  and ginst7170 (P1_U3657, P1_U3656, P1_U4286, P1_U4287);
  and ginst7171 (P1_U3658, P1_U4289, P1_U4290, P1_U4291, P1_U4292);
  and ginst7172 (P1_U3659, P1_U4301, P1_U4302);
  and ginst7173 (P1_U3660, P1_U4303, P1_U4304);
  and ginst7174 (P1_U3661, P1_U3660, P1_U4305, P1_U4306);
  and ginst7175 (P1_U3662, P1_U4308, P1_U4309, P1_U4310, P1_U4311);
  and ginst7176 (P1_U3663, P1_U4320, P1_U4321);
  and ginst7177 (P1_U3664, P1_U4322, P1_U4323);
  and ginst7178 (P1_U3665, P1_U3664, P1_U4324, P1_U4325);
  and ginst7179 (P1_U3666, P1_U4327, P1_U4328, P1_U4329, P1_U4330);
  and ginst7180 (P1_U3667, P1_U4339, P1_U4340);
  and ginst7181 (P1_U3668, P1_U4341, P1_U4342);
  and ginst7182 (P1_U3669, P1_U3668, P1_U4343, P1_U4344);
  and ginst7183 (P1_U3670, P1_U4346, P1_U4347, P1_U4348, P1_U4349);
  and ginst7184 (P1_U3671, P1_U4358, P1_U4359);
  and ginst7185 (P1_U3672, P1_U4360, P1_U4361);
  and ginst7186 (P1_U3673, P1_U3672, P1_U4362, P1_U4363);
  and ginst7187 (P1_U3674, P1_U4365, P1_U4366, P1_U4367, P1_U4368);
  and ginst7188 (P1_U3675, P1_U4377, P1_U4378);
  and ginst7189 (P1_U3676, P1_U4379, P1_U4380);
  and ginst7190 (P1_U3677, P1_U3676, P1_U4381, P1_U4382);
  and ginst7191 (P1_U3678, P1_U4384, P1_U4385, P1_U4386, P1_U4387);
  and ginst7192 (P1_U3679, P1_U4396, P1_U4397);
  and ginst7193 (P1_U3680, P1_U4398, P1_U4399);
  and ginst7194 (P1_U3681, P1_U3680, P1_U4400, P1_U4401);
  and ginst7195 (P1_U3682, P1_U4403, P1_U4404, P1_U4405, P1_U4406);
  and ginst7196 (P1_U3683, P1_U4415, P1_U4416);
  and ginst7197 (P1_U3684, P1_U4417, P1_U4418);
  and ginst7198 (P1_U3685, P1_U3684, P1_U4419, P1_U4420);
  and ginst7199 (P1_U3686, P1_U4422, P1_U4423, P1_U4424, P1_U4425);
  and ginst7200 (P1_U3687, P1_U4434, P1_U4435);
  and ginst7201 (P1_U3688, P1_U4436, P1_U4437);
  and ginst7202 (P1_U3689, P1_U3688, P1_U4438, P1_U4439);
  and ginst7203 (P1_U3690, P1_U4441, P1_U4442, P1_U4443, P1_U4444);
  and ginst7204 (P1_U3691, P1_U4453, P1_U4454);
  and ginst7205 (P1_U3692, P1_U4455, P1_U4456);
  and ginst7206 (P1_U3693, P1_U3692, P1_U4457, P1_U4458);
  and ginst7207 (P1_U3694, P1_U4460, P1_U4461, P1_U4462, P1_U4463);
  and ginst7208 (P1_U3695, P1_U4472, P1_U4473);
  and ginst7209 (P1_U3696, P1_U4474, P1_U4475);
  and ginst7210 (P1_U3697, P1_U3696, P1_U4476, P1_U4477);
  and ginst7211 (P1_U3698, P1_U4479, P1_U4480, P1_U4481, P1_U4482);
  and ginst7212 (P1_U3699, P1_U4491, P1_U4492);
  and ginst7213 (P1_U3700, P1_U4493, P1_U4494);
  and ginst7214 (P1_U3701, P1_U3700, P1_U4495, P1_U4496);
  and ginst7215 (P1_U3702, P1_U4498, P1_U4499, P1_U4500, P1_U4501);
  and ginst7216 (P1_U3703, P1_U4510, P1_U4511);
  and ginst7217 (P1_U3704, P1_U4512, P1_U4513);
  and ginst7218 (P1_U3705, P1_U3704, P1_U4514, P1_U4515);
  and ginst7219 (P1_U3706, P1_U4517, P1_U4518, P1_U4519, P1_U4520);
  and ginst7220 (P1_U3707, P1_U4529, P1_U4530);
  and ginst7221 (P1_U3708, P1_U4531, P1_U4532);
  and ginst7222 (P1_U3709, P1_U3708, P1_U4533, P1_U4534);
  and ginst7223 (P1_U3710, P1_U4536, P1_U4537, P1_U4538, P1_U4539);
  and ginst7224 (P1_U3711, P1_U4548, P1_U4549);
  and ginst7225 (P1_U3712, P1_U4550, P1_U4551);
  and ginst7226 (P1_U3713, P1_U3712, P1_U4552, P1_U4553);
  and ginst7227 (P1_U3714, P1_U4555, P1_U4556, P1_U4557, P1_U4558);
  and ginst7228 (P1_U3715, P1_U4567, P1_U4568);
  and ginst7229 (P1_U3716, P1_U4569, P1_U4570);
  and ginst7230 (P1_U3717, P1_U3716, P1_U4571, P1_U4572);
  and ginst7231 (P1_U3718, P1_U4574, P1_U4575, P1_U4576, P1_U4577);
  and ginst7232 (P1_U3719, P1_U4586, P1_U4587);
  and ginst7233 (P1_U3720, P1_U4588, P1_U4589);
  and ginst7234 (P1_U3721, P1_U3720, P1_U4590, P1_U4591);
  and ginst7235 (P1_U3722, P1_U4593, P1_U4594, P1_U4595, P1_U4596);
  and ginst7236 (P1_U3723, P1_U4605, P1_U4606);
  and ginst7237 (P1_U3724, P1_U4607, P1_U4608);
  and ginst7238 (P1_U3725, P1_U3724, P1_U4609, P1_U4610);
  and ginst7239 (P1_U3726, P1_U4612, P1_U4613, P1_U4614, P1_U4615);
  and ginst7240 (P1_U3727, P1_U4624, P1_U4625);
  and ginst7241 (P1_U3728, P1_U4626, P1_U4627);
  and ginst7242 (P1_U3729, P1_U3728, P1_U4628, P1_U4629);
  and ginst7243 (P1_U3730, P1_U4631, P1_U4632, P1_U4633, P1_U4634);
  and ginst7244 (P1_U3731, P1_U4643, P1_U4644);
  and ginst7245 (P1_U3732, P1_U4645, P1_U4646);
  and ginst7246 (P1_U3733, P1_U3732, P1_U4647, P1_U4648);
  and ginst7247 (P1_U3734, P1_U4650, P1_U4651, P1_U4652, P1_U4653);
  and ginst7248 (P1_U3735, P1_U4662, P1_U4663);
  and ginst7249 (P1_U3736, P1_U4664, P1_U4665);
  and ginst7250 (P1_U3737, P1_U3736, P1_U4666, P1_U4667);
  and ginst7251 (P1_U3738, P1_U4669, P1_U4670, P1_U4671, P1_U4672);
  and ginst7252 (P1_U3739, P1_U4681, P1_U4682);
  and ginst7253 (P1_U3740, P1_U4683, P1_U4684);
  and ginst7254 (P1_U3741, P1_U3740, P1_U4685, P1_U4686);
  and ginst7255 (P1_U3742, P1_U4688, P1_U4689, P1_U4690, P1_U4691);
  and ginst7256 (P1_U3743, P1_U3987, P1_U4698);
  and ginst7257 (P1_U3744, P1_U4701, P1_U4702, P1_U4704);
  and ginst7258 (P1_U3745, P1_U4705, P1_U4707);
  and ginst7259 (P1_U3746, P1_U4709, P1_U4710, P1_U4711);
  and ginst7260 (P1_U3747, P1_U3987, P1_U4698);
  and ginst7261 (P1_U3748, P1_U3022, P1_U3451);
  and ginst7262 (P1_U3749, P1_U3452, P1_U3969, P1_U5719);
  and ginst7263 (P1_U3750, P1_U4727, P1_U4728, P1_U4729);
  and ginst7264 (P1_U3751, P1_U3915, P1_U4730, P1_U4731);
  and ginst7265 (P1_U3752, P1_U4732, P1_U4733, P1_U4734);
  and ginst7266 (P1_U3753, P1_U3916, P1_U4735, P1_U4736);
  and ginst7267 (P1_U3754, P1_U4737, P1_U4738, P1_U4739);
  and ginst7268 (P1_U3755, P1_U3917, P1_U4740, P1_U4741);
  and ginst7269 (P1_U3756, P1_U4742, P1_U4743, P1_U4744);
  and ginst7270 (P1_U3757, P1_U4745, P1_U4746);
  and ginst7271 (P1_U3758, P1_U4747, P1_U4748);
  and ginst7272 (P1_U3759, P1_U4750, P1_U4751);
  and ginst7273 (P1_U3760, P1_U4752, P1_U4753);
  and ginst7274 (P1_U3761, P1_U4755, P1_U4756);
  and ginst7275 (P1_U3762, P1_U4757, P1_U4758);
  and ginst7276 (P1_U3763, P1_U4760, P1_U4761);
  and ginst7277 (P1_U3764, P1_U4762, P1_U4763);
  and ginst7278 (P1_U3765, P1_U4765, P1_U4766);
  and ginst7279 (P1_U3766, P1_U4767, P1_U4768);
  and ginst7280 (P1_U3767, P1_U4770, P1_U4771);
  and ginst7281 (P1_U3768, P1_U4772, P1_U4773);
  and ginst7282 (P1_U3769, P1_U4775, P1_U4776);
  and ginst7283 (P1_U3770, P1_U4777, P1_U4778);
  and ginst7284 (P1_U3771, P1_U4780, P1_U4781);
  and ginst7285 (P1_U3772, P1_U4782, P1_U4783, P1_U4784);
  and ginst7286 (P1_U3773, P1_U4785, P1_U4786);
  and ginst7287 (P1_U3774, P1_U4787, P1_U4788, P1_U4789);
  and ginst7288 (P1_U3775, P1_U4790, P1_U4791);
  and ginst7289 (P1_U3776, P1_U4792, P1_U4793, P1_U4794);
  and ginst7290 (P1_U3777, P1_U4795, P1_U4796);
  and ginst7291 (P1_U3778, P1_U4797, P1_U4798, P1_U4799, P1_U4800, P1_U4801);
  and ginst7292 (P1_U3779, P1_U4802, P1_U4803, P1_U4804, P1_U4805, P1_U4806);
  and ginst7293 (P1_U3780, P1_U4807, P1_U4808, P1_U4809, P1_U4810, P1_U4811);
  and ginst7294 (P1_U3781, P1_U4812, P1_U4813, P1_U4814, P1_U4815, P1_U4816);
  and ginst7295 (P1_U3782, P1_U4817, P1_U4818, P1_U4819, P1_U4820, P1_U4821);
  and ginst7296 (P1_U3783, P1_U4822, P1_U4823, P1_U4824, P1_U4825, P1_U4826);
  and ginst7297 (P1_U3784, P1_U4827, P1_U4828, P1_U4829);
  and ginst7298 (P1_U3785, P1_U4830, P1_U4831);
  and ginst7299 (P1_U3786, P1_U4832, P1_U4833, P1_U4834, P1_U4835, P1_U4836);
  and ginst7300 (P1_U3787, P1_U4837, P1_U4838, P1_U4839);
  and ginst7301 (P1_U3788, P1_U4840, P1_U4841);
  and ginst7302 (P1_U3789, P1_U4842, P1_U4843, P1_U4844);
  and ginst7303 (P1_U3790, P1_U4845, P1_U4846);
  and ginst7304 (P1_U3791, P1_U4847, P1_U4848);
  and ginst7305 (P1_U3792, P1_U4850, P1_U4851);
  and ginst7306 (P1_U3793, P1_U4852, P1_U4853);
  and ginst7307 (P1_U3794, P1_U4855, P1_U4856);
  and ginst7308 (P1_U3795, P1_U4857, P1_U4858);
  and ginst7309 (P1_U3796, P1_U4860, P1_U4861);
  and ginst7310 (P1_U3797, P1_U4862, P1_U4863);
  and ginst7311 (P1_U3798, P1_U4865, P1_U4866);
  and ginst7312 (P1_U3799, P1_U4867, P1_U4868);
  and ginst7313 (P1_U3800, P1_U4870, P1_U4871);
  and ginst7314 (P1_U3801, P1_U4707, P1_U5657, P1_U5658);
  and ginst7315 (P1_U3802, P1_U5659, P1_U5660);
  and ginst7316 (P1_U3803, P1_U3366, P1_U3370, P1_U3419);
  and ginst7317 (P1_U3804, P1_U3361, P1_U3365, P1_U3368);
  and ginst7318 (P1_U3805, P1_U3362, P1_U3364);
  and ginst7319 (P1_U3806, P1_U3420, P1_U3805);
  and ginst7320 (P1_U3807, P1_STATE_REG_SCAN_IN, P1_U3438);
  and ginst7321 (P1_U3808, P1_U4891, P1_U4892);
  and ginst7322 (P1_U3809, P1_U4893, P1_U4894, P1_U4895);
  and ginst7323 (P1_U3810, P1_U4901, P1_U4902);
  and ginst7324 (P1_U3811, P1_U4903, P1_U4904, P1_U4905);
  and ginst7325 (P1_U3812, P1_U4911, P1_U4912);
  and ginst7326 (P1_U3813, P1_U4913, P1_U4914, P1_U4915);
  and ginst7327 (P1_U3814, P1_U4921, P1_U4922);
  and ginst7328 (P1_U3815, P1_U4923, P1_U4924, P1_U4925);
  and ginst7329 (P1_U3816, P1_U4931, P1_U4932);
  and ginst7330 (P1_U3817, P1_U4933, P1_U4934, P1_U4935);
  and ginst7331 (P1_U3818, P1_U4941, P1_U4942);
  and ginst7332 (P1_U3819, P1_U4943, P1_U4944, P1_U4945);
  and ginst7333 (P1_U3820, P1_U4951, P1_U4952);
  and ginst7334 (P1_U3821, P1_U4953, P1_U4954, P1_U4955);
  and ginst7335 (P1_U3822, P1_U4961, P1_U4962);
  and ginst7336 (P1_U3823, P1_U4963, P1_U4964, P1_U4965);
  and ginst7337 (P1_U3824, P1_U4971, P1_U4972);
  and ginst7338 (P1_U3825, P1_U4973, P1_U4974, P1_U4975);
  and ginst7339 (P1_U3826, P1_U4981, P1_U4982);
  and ginst7340 (P1_U3827, P1_U4983, P1_U4984, P1_U4985);
  and ginst7341 (P1_U3828, P1_U4991, P1_U4992);
  and ginst7342 (P1_U3829, P1_U4993, P1_U4994, P1_U4995);
  and ginst7343 (P1_U3830, P1_U5001, P1_U5002);
  and ginst7344 (P1_U3831, P1_U5003, P1_U5004, P1_U5005);
  and ginst7345 (P1_U3832, P1_U5011, P1_U5012);
  and ginst7346 (P1_U3833, P1_U5013, P1_U5014, P1_U5015);
  and ginst7347 (P1_U3834, P1_U5020, P1_U5021, P1_U5022);
  and ginst7348 (P1_U3835, P1_U5023, P1_U5024, P1_U5025);
  and ginst7349 (P1_U3836, P1_U5030, P1_U5031, P1_U5032);
  and ginst7350 (P1_U3837, P1_U5033, P1_U5034, P1_U5035);
  and ginst7351 (P1_U3838, P1_U3998, P1_U5040);
  and ginst7352 (P1_U3839, P1_U3838, P1_U5041, P1_U5042);
  and ginst7353 (P1_U3840, P1_U5043, P1_U5044, P1_U5045);
  and ginst7354 (P1_U3841, P1_U5050, P1_U5051, P1_U5052);
  and ginst7355 (P1_U3842, P1_U5053, P1_U5054, P1_U5055);
  and ginst7356 (P1_U3843, P1_U3998, P1_U5060);
  and ginst7357 (P1_U3844, P1_U3843, P1_U5061, P1_U5062);
  and ginst7358 (P1_U3845, P1_U5063, P1_U5064, P1_U5065);
  and ginst7359 (P1_U3846, P1_U5070, P1_U5071, P1_U5072);
  and ginst7360 (P1_U3847, P1_U5073, P1_U5074, P1_U5075);
  and ginst7361 (P1_U3848, P1_U5080, P1_U5081, P1_U5082);
  and ginst7362 (P1_U3849, P1_U5083, P1_U5084, P1_U5085);
  and ginst7363 (P1_U3850, P1_STATE_REG_SCAN_IN, P1_U3428);
  and ginst7364 (P1_U3851, P1_U3424, P1_U3850);
  and ginst7365 (P1_U3852, P1_U6111, P1_U6114, P1_U6117);
  and ginst7366 (P1_U3853, P1_U3852, P1_U3854, P1_U6129);
  and ginst7367 (P1_U3854, P1_U6120, P1_U6123, P1_U6126);
  and ginst7368 (P1_U3855, P1_U6135, P1_U6138, P1_U6141);
  and ginst7369 (P1_U3856, P1_U6144, P1_U6147, P1_U6150);
  and ginst7370 (P1_U3857, P1_U3855, P1_U3856, P1_U6132);
  and ginst7371 (P1_U3858, P1_U3862, P1_U3863, P1_U6075, P1_U6078, P1_U6081);
  and ginst7372 (P1_U3859, P1_U6156, P1_U6159, P1_U6162, P1_U6165, P1_U6168);
  and ginst7373 (P1_U3860, P1_U3853, P1_U3857, P1_U3859, P1_U6108, P1_U6153);
  and ginst7374 (P1_U3861, P1_U3858, P1_U6102);
  and ginst7375 (P1_U3862, P1_U6084, P1_U6087, P1_U6090, P1_U6093);
  and ginst7376 (P1_U3863, P1_U6096, P1_U6099);
  and ginst7377 (P1_U3864, P1_U5087, P1_U5090, P1_U5091);
  and ginst7378 (P1_U3865, P1_U3052, P1_U5690);
  and ginst7379 (P1_U3866, P1_U5651, P1_U5652);
  and ginst7380 (P1_U3867, P1_U3451, P1_U3452);
  and ginst7381 (P1_U3868, P1_U3369, P1_U3371, P1_U3420);
  and ginst7382 (P1_U3869, P1_U3969, P1_U5677);
  and ginst7383 (P1_U3870, P1_U3424, P1_U3869);
  and ginst7384 (P1_U3871, P1_U3022, P1_U5100);
  and ginst7385 (P1_U3872, P1_U5146, P1_U5147);
  and ginst7386 (P1_U3873, P1_U3078, P1_U3994);
  and ginst7387 (P1_U3874, P1_U5187, P1_U5188);
  and ginst7388 (P1_U3875, P1_U5190, P1_U5191);
  and ginst7389 (P1_U3876, P1_U5280, P1_U5281);
  and ginst7390 (P1_U3877, P1_U3433, P1_U5366);
  and ginst7391 (P1_U3878, P1_U5431, P1_U5432);
  and ginst7392 (P1_U3879, P1_U3438, P1_U5514);
  and ginst7393 (P1_U3880, P1_U3438, P1_U5516);
  and ginst7394 (P1_U3881, P1_U3438, P1_U5518);
  and ginst7395 (P1_U3882, P1_U3438, P1_U5520);
  and ginst7396 (P1_U3883, P1_U3438, P1_U5522);
  and ginst7397 (P1_U3884, P1_U3438, P1_U5524);
  and ginst7398 (P1_U3885, P1_U3438, P1_U5526);
  and ginst7399 (P1_U3886, P1_U3438, P1_U5528);
  and ginst7400 (P1_U3887, P1_U3438, P1_U5530);
  and ginst7401 (P1_U3888, P1_U3438, P1_U5533);
  and ginst7402 (P1_U3889, P1_U3438, P1_U5535);
  and ginst7403 (P1_U3890, P1_U3438, P1_U5537);
  and ginst7404 (P1_U3891, P1_U3438, P1_U5539);
  and ginst7405 (P1_U3892, P1_U3438, P1_U5541);
  and ginst7406 (P1_U3893, P1_U3438, P1_U5543);
  and ginst7407 (P1_U3894, P1_U3438, P1_U5555);
  and ginst7408 (P1_U3895, P1_U5585, P1_U5587);
  and ginst7409 (P1_U3896, P1_U5588, P1_U5590);
  and ginst7410 (P1_U3897, P1_U5591, P1_U5593);
  and ginst7411 (P1_U3898, P1_U5594, P1_U5596);
  and ginst7412 (P1_U3899, P1_U5597, P1_U5599);
  and ginst7413 (P1_U3900, P1_U5600, P1_U5602);
  and ginst7414 (P1_U3901, P1_U5603, P1_U5605);
  and ginst7415 (P1_U3902, P1_U5606, P1_U5608);
  and ginst7416 (P1_U3903, P1_U5609, P1_U5611);
  and ginst7417 (P1_U3904, P1_U5615, P1_U5617);
  and ginst7418 (P1_U3905, P1_U5618, P1_U5620);
  and ginst7419 (P1_U3906, P1_U5621, P1_U5623);
  and ginst7420 (P1_U3907, P1_U5624, P1_U5626);
  and ginst7421 (P1_U3908, P1_U5627, P1_U5629);
  and ginst7422 (P1_U3909, P1_U5630, P1_U5632);
  not ginst7423 (P1_U3910, P1_IR_REG_31__SCAN_IN);
  nand ginst7424 (P1_U3911, P1_U3022, P1_U3360);
  nand ginst7425 (P1_U3912, P1_U5699, P1_U5702);
  nand ginst7426 (P1_U3913, P1_U3047, P1_U3632);
  nand ginst7427 (P1_U3914, P1_U3047, P1_U3748);
  and ginst7428 (P1_U3915, P1_U5941, P1_U5942);
  and ginst7429 (P1_U3916, P1_U5943, P1_U5944);
  and ginst7430 (P1_U3917, P1_U5945, P1_U5946);
  and ginst7431 (P1_U3918, P1_U5947, P1_U5948);
  and ginst7432 (P1_U3919, P1_U5949, P1_U5950);
  and ginst7433 (P1_U3920, P1_U5951, P1_U5952);
  and ginst7434 (P1_U3921, P1_U5953, P1_U5954);
  and ginst7435 (P1_U3922, P1_U5955, P1_U5956);
  and ginst7436 (P1_U3923, P1_U5957, P1_U5958);
  and ginst7437 (P1_U3924, P1_U5959, P1_U5960);
  and ginst7438 (P1_U3925, P1_U5961, P1_U5962);
  and ginst7439 (P1_U3926, P1_U5963, P1_U5964);
  and ginst7440 (P1_U3927, P1_U5965, P1_U5966);
  and ginst7441 (P1_U3928, P1_U5967, P1_U5968);
  and ginst7442 (P1_U3929, P1_U5969, P1_U5970);
  and ginst7443 (P1_U3930, P1_U5971, P1_U5972);
  and ginst7444 (P1_U3931, P1_U5973, P1_U5974);
  and ginst7445 (P1_U3932, P1_U5975, P1_U5976);
  and ginst7446 (P1_U3933, P1_U5977, P1_U5978);
  and ginst7447 (P1_U3934, P1_U5979, P1_U5980);
  and ginst7448 (P1_U3935, P1_U5981, P1_U5982);
  and ginst7449 (P1_U3936, P1_U5983, P1_U5984);
  and ginst7450 (P1_U3937, P1_U5985, P1_U5986);
  and ginst7451 (P1_U3938, P1_U5987, P1_U5988);
  and ginst7452 (P1_U3939, P1_U5989, P1_U5990);
  and ginst7453 (P1_U3940, P1_U5991, P1_U5992);
  and ginst7454 (P1_U3941, P1_U5993, P1_U5994);
  and ginst7455 (P1_U3942, P1_U5995, P1_U5996);
  and ginst7456 (P1_U3943, P1_U5997, P1_U5998);
  and ginst7457 (P1_U3944, P1_U5999, P1_U6000);
  nand ginst7458 (P1_U3945, P1_U3056, P1_U3747);
  and ginst7459 (P1_U3946, P1_U6001, P1_U6002);
  and ginst7460 (P1_U3947, P1_U6003, P1_U6004);
  not ginst7461 (P1_U3948, P1_R1375_U14);
  not ginst7462 (P1_U3949, P1_R1360_U14);
  and ginst7463 (P1_U3950, P1_U6071, P1_U6072);
  nand ginst7464 (P1_U3951, P1_U3860, P1_U3861, P1_U6105);
  not ginst7465 (P1_U3952, P1_R1352_U6);
  not ginst7466 (P1_U3953, P1_U3372);
  not ginst7467 (P1_U3954, P1_U3426);
  not ginst7468 (P1_U3955, P1_U3428);
  not ginst7469 (P1_U3956, P1_U3370);
  not ginst7470 (P1_U3957, P1_U3419);
  not ginst7471 (P1_U3958, P1_U3366);
  not ginst7472 (P1_U3959, P1_U3365);
  not ginst7473 (P1_U3960, P1_U3368);
  not ginst7474 (P1_U3961, P1_U3361);
  not ginst7475 (P1_U3962, P1_U3364);
  not ginst7476 (P1_U3963, P1_U3362);
  not ginst7477 (P1_U3964, P1_U3420);
  not ginst7478 (P1_U3965, P1_U3418);
  nand ginst7479 (P1_U3966, P1_U3049, P1_U4001);
  not ginst7480 (P1_U3967, P1_U3371);
  not ginst7481 (P1_U3968, P1_U3369);
  nand ginst7482 (P1_U3969, P1_U3367, P1_U3987);
  nand ginst7483 (P1_U3970, P1_U3049, P1_U3421);
  not ginst7484 (P1_U3971, P1_U3912);
  not ginst7485 (P1_U3972, P1_U3430);
  not ginst7486 (P1_U3973, P1_U3425);
  not ginst7487 (P1_U3974, P1_U3411);
  not ginst7488 (P1_U3975, P1_U3409);
  not ginst7489 (P1_U3976, P1_U3407);
  not ginst7490 (P1_U3977, P1_U3405);
  not ginst7491 (P1_U3978, P1_U3403);
  not ginst7492 (P1_U3979, P1_U3401);
  not ginst7493 (P1_U3980, P1_U3399);
  not ginst7494 (P1_U3981, P1_U3397);
  not ginst7495 (P1_U3982, P1_U3395);
  not ginst7496 (P1_U3983, P1_U3415);
  not ginst7497 (P1_U3984, P1_U3414);
  not ginst7498 (P1_U3985, P1_U3413);
  not ginst7499 (P1_U3986, P1_U3427);
  not ginst7500 (P1_U3987, P1_U3373);
  not ginst7501 (P1_U3988, P1_U3416);
  not ginst7502 (P1_U3989, P1_U3417);
  not ginst7503 (P1_U3990, P1_U3914);
  not ginst7504 (P1_U3991, P1_U3913);
  not ginst7505 (P1_U3992, P1_U3911);
  not ginst7506 (P1_U3993, P1_U3945);
  not ginst7507 (P1_U3994, P1_U3431);
  nand ginst7508 (P1_U3995, P1_STATE_REG_SCAN_IN, P1_U3432);
  nand ginst7509 (P1_U3996, P1_U3022, P1_U3965);
  not ginst7510 (P1_U3997, P1_U3429);
  nand ginst7511 (P1_U3998, P1_U3212, P1_U3973);
  not ginst7512 (P1_U3999, P1_U3424);
  not ginst7513 (P1_U4000, P1_U3433);
  not ginst7514 (P1_U4001, P1_U3363);
  not ginst7515 (P1_U4002, P1_U3367);
  not ginst7516 (P1_U4003, P1_U3358);
  not ginst7517 (P1_U4004, P1_U3357);
  nand ginst7518 (P1_U4005, P1_U3086, U88);
  nand ginst7519 (P1_U4006, P1_IR_REG_0__SCAN_IN, P1_U3028);
  nand ginst7520 (P1_U4007, P1_IR_REG_0__SCAN_IN, P1_U4004);
  nand ginst7521 (P1_U4008, P1_U3086, U77);
  nand ginst7522 (P1_U4009, P1_SUB_84_U40, P1_U3028);
  nand ginst7523 (P1_U4010, P1_IR_REG_1__SCAN_IN, P1_U4004);
  nand ginst7524 (P1_U4011, P1_U3086, U66);
  nand ginst7525 (P1_U4012, P1_SUB_84_U21, P1_U3028);
  nand ginst7526 (P1_U4013, P1_IR_REG_2__SCAN_IN, P1_U4004);
  nand ginst7527 (P1_U4014, P1_U3086, U63);
  nand ginst7528 (P1_U4015, P1_SUB_84_U22, P1_U3028);
  nand ginst7529 (P1_U4016, P1_IR_REG_3__SCAN_IN, P1_U4004);
  nand ginst7530 (P1_U4017, P1_U3086, U62);
  nand ginst7531 (P1_U4018, P1_SUB_84_U23, P1_U3028);
  nand ginst7532 (P1_U4019, P1_IR_REG_4__SCAN_IN, P1_U4004);
  nand ginst7533 (P1_U4020, P1_U3086, U61);
  nand ginst7534 (P1_U4021, P1_SUB_84_U162, P1_U3028);
  nand ginst7535 (P1_U4022, P1_IR_REG_5__SCAN_IN, P1_U4004);
  nand ginst7536 (P1_U4023, P1_U3086, U60);
  nand ginst7537 (P1_U4024, P1_SUB_84_U24, P1_U3028);
  nand ginst7538 (P1_U4025, P1_IR_REG_6__SCAN_IN, P1_U4004);
  nand ginst7539 (P1_U4026, P1_U3086, U59);
  nand ginst7540 (P1_U4027, P1_SUB_84_U25, P1_U3028);
  nand ginst7541 (P1_U4028, P1_IR_REG_7__SCAN_IN, P1_U4004);
  nand ginst7542 (P1_U4029, P1_U3086, U58);
  nand ginst7543 (P1_U4030, P1_SUB_84_U26, P1_U3028);
  nand ginst7544 (P1_U4031, P1_IR_REG_8__SCAN_IN, P1_U4004);
  nand ginst7545 (P1_U4032, P1_U3086, U57);
  nand ginst7546 (P1_U4033, P1_SUB_84_U160, P1_U3028);
  nand ginst7547 (P1_U4034, P1_IR_REG_9__SCAN_IN, P1_U4004);
  nand ginst7548 (P1_U4035, P1_U3086, U87);
  nand ginst7549 (P1_U4036, P1_SUB_84_U6, P1_U3028);
  nand ginst7550 (P1_U4037, P1_IR_REG_10__SCAN_IN, P1_U4004);
  nand ginst7551 (P1_U4038, P1_U3086, U86);
  nand ginst7552 (P1_U4039, P1_SUB_84_U7, P1_U3028);
  nand ginst7553 (P1_U4040, P1_IR_REG_11__SCAN_IN, P1_U4004);
  nand ginst7554 (P1_U4041, P1_U3086, U85);
  nand ginst7555 (P1_U4042, P1_SUB_84_U8, P1_U3028);
  nand ginst7556 (P1_U4043, P1_IR_REG_12__SCAN_IN, P1_U4004);
  nand ginst7557 (P1_U4044, P1_U3086, U84);
  nand ginst7558 (P1_U4045, P1_SUB_84_U179, P1_U3028);
  nand ginst7559 (P1_U4046, P1_IR_REG_13__SCAN_IN, P1_U4004);
  nand ginst7560 (P1_U4047, P1_U3086, U83);
  nand ginst7561 (P1_U4048, P1_SUB_84_U9, P1_U3028);
  nand ginst7562 (P1_U4049, P1_IR_REG_14__SCAN_IN, P1_U4004);
  nand ginst7563 (P1_U4050, P1_U3086, U82);
  nand ginst7564 (P1_U4051, P1_SUB_84_U10, P1_U3028);
  nand ginst7565 (P1_U4052, P1_IR_REG_15__SCAN_IN, P1_U4004);
  nand ginst7566 (P1_U4053, P1_U3086, U81);
  nand ginst7567 (P1_U4054, P1_SUB_84_U11, P1_U3028);
  nand ginst7568 (P1_U4055, P1_IR_REG_16__SCAN_IN, P1_U4004);
  nand ginst7569 (P1_U4056, P1_U3086, U80);
  nand ginst7570 (P1_U4057, P1_SUB_84_U177, P1_U3028);
  nand ginst7571 (P1_U4058, P1_IR_REG_17__SCAN_IN, P1_U4004);
  nand ginst7572 (P1_U4059, P1_U3086, U79);
  nand ginst7573 (P1_U4060, P1_SUB_84_U12, P1_U3028);
  nand ginst7574 (P1_U4061, P1_IR_REG_18__SCAN_IN, P1_U4004);
  nand ginst7575 (P1_U4062, P1_U3086, U78);
  nand ginst7576 (P1_U4063, P1_SUB_84_U13, P1_U3028);
  nand ginst7577 (P1_U4064, P1_IR_REG_19__SCAN_IN, P1_U4004);
  nand ginst7578 (P1_U4065, P1_U3086, U76);
  nand ginst7579 (P1_U4066, P1_SUB_84_U14, P1_U3028);
  nand ginst7580 (P1_U4067, P1_IR_REG_20__SCAN_IN, P1_U4004);
  nand ginst7581 (P1_U4068, P1_U3086, U75);
  nand ginst7582 (P1_U4069, P1_SUB_84_U173, P1_U3028);
  nand ginst7583 (P1_U4070, P1_IR_REG_21__SCAN_IN, P1_U4004);
  nand ginst7584 (P1_U4071, P1_U3086, U74);
  nand ginst7585 (P1_U4072, P1_SUB_84_U15, P1_U3028);
  nand ginst7586 (P1_U4073, P1_IR_REG_22__SCAN_IN, P1_U4004);
  nand ginst7587 (P1_U4074, P1_U3086, U73);
  nand ginst7588 (P1_U4075, P1_SUB_84_U16, P1_U3028);
  nand ginst7589 (P1_U4076, P1_IR_REG_23__SCAN_IN, P1_U4004);
  nand ginst7590 (P1_U4077, P1_U3086, U72);
  nand ginst7591 (P1_U4078, P1_SUB_84_U17, P1_U3028);
  nand ginst7592 (P1_U4079, P1_IR_REG_24__SCAN_IN, P1_U4004);
  nand ginst7593 (P1_U4080, P1_U3086, U71);
  nand ginst7594 (P1_U4081, P1_SUB_84_U170, P1_U3028);
  nand ginst7595 (P1_U4082, P1_IR_REG_25__SCAN_IN, P1_U4004);
  nand ginst7596 (P1_U4083, P1_U3086, U70);
  nand ginst7597 (P1_U4084, P1_SUB_84_U18, P1_U3028);
  nand ginst7598 (P1_U4085, P1_IR_REG_26__SCAN_IN, P1_U4004);
  nand ginst7599 (P1_U4086, P1_U3086, U69);
  nand ginst7600 (P1_U4087, P1_SUB_84_U42, P1_U3028);
  nand ginst7601 (P1_U4088, P1_IR_REG_27__SCAN_IN, P1_U4004);
  nand ginst7602 (P1_U4089, P1_U3086, U68);
  nand ginst7603 (P1_U4090, P1_SUB_84_U19, P1_U3028);
  nand ginst7604 (P1_U4091, P1_IR_REG_28__SCAN_IN, P1_U4004);
  nand ginst7605 (P1_U4092, P1_U3086, U67);
  nand ginst7606 (P1_U4093, P1_SUB_84_U20, P1_U3028);
  nand ginst7607 (P1_U4094, P1_IR_REG_29__SCAN_IN, P1_U4004);
  nand ginst7608 (P1_U4095, P1_U3086, U65);
  nand ginst7609 (P1_U4096, P1_SUB_84_U165, P1_U3028);
  nand ginst7610 (P1_U4097, P1_IR_REG_30__SCAN_IN, P1_U4004);
  nand ginst7611 (P1_U4098, P1_U3086, U64);
  nand ginst7612 (P1_U4099, P1_SUB_84_U41, P1_U3028);
  nand ginst7613 (P1_U4100, P1_IR_REG_31__SCAN_IN, P1_U4004);
  not ginst7614 (P1_U4101, P1_U3360);
  not ginst7615 (P1_U4102, P1_U3421);
  nand ginst7616 (P1_U4103, P1_U3358, P1_U5666);
  nand ginst7617 (P1_U4104, P1_U3358, P1_U5669);
  nand ginst7618 (P1_U4105, P1_D_REG_10__SCAN_IN, P1_U4101);
  nand ginst7619 (P1_U4106, P1_D_REG_11__SCAN_IN, P1_U4101);
  nand ginst7620 (P1_U4107, P1_D_REG_12__SCAN_IN, P1_U4101);
  nand ginst7621 (P1_U4108, P1_D_REG_13__SCAN_IN, P1_U4101);
  nand ginst7622 (P1_U4109, P1_D_REG_14__SCAN_IN, P1_U4101);
  nand ginst7623 (P1_U4110, P1_D_REG_15__SCAN_IN, P1_U4101);
  nand ginst7624 (P1_U4111, P1_D_REG_16__SCAN_IN, P1_U4101);
  nand ginst7625 (P1_U4112, P1_D_REG_17__SCAN_IN, P1_U4101);
  nand ginst7626 (P1_U4113, P1_D_REG_18__SCAN_IN, P1_U4101);
  nand ginst7627 (P1_U4114, P1_D_REG_19__SCAN_IN, P1_U4101);
  nand ginst7628 (P1_U4115, P1_D_REG_20__SCAN_IN, P1_U4101);
  nand ginst7629 (P1_U4116, P1_D_REG_21__SCAN_IN, P1_U4101);
  nand ginst7630 (P1_U4117, P1_D_REG_22__SCAN_IN, P1_U4101);
  nand ginst7631 (P1_U4118, P1_D_REG_23__SCAN_IN, P1_U4101);
  nand ginst7632 (P1_U4119, P1_D_REG_24__SCAN_IN, P1_U4101);
  nand ginst7633 (P1_U4120, P1_D_REG_25__SCAN_IN, P1_U4101);
  nand ginst7634 (P1_U4121, P1_D_REG_26__SCAN_IN, P1_U4101);
  nand ginst7635 (P1_U4122, P1_D_REG_27__SCAN_IN, P1_U4101);
  nand ginst7636 (P1_U4123, P1_D_REG_28__SCAN_IN, P1_U4101);
  nand ginst7637 (P1_U4124, P1_D_REG_29__SCAN_IN, P1_U4101);
  nand ginst7638 (P1_U4125, P1_D_REG_2__SCAN_IN, P1_U4101);
  nand ginst7639 (P1_U4126, P1_D_REG_30__SCAN_IN, P1_U4101);
  nand ginst7640 (P1_U4127, P1_D_REG_31__SCAN_IN, P1_U4101);
  nand ginst7641 (P1_U4128, P1_D_REG_3__SCAN_IN, P1_U4101);
  nand ginst7642 (P1_U4129, P1_D_REG_4__SCAN_IN, P1_U4101);
  nand ginst7643 (P1_U4130, P1_D_REG_5__SCAN_IN, P1_U4101);
  nand ginst7644 (P1_U4131, P1_D_REG_6__SCAN_IN, P1_U4101);
  nand ginst7645 (P1_U4132, P1_D_REG_7__SCAN_IN, P1_U4101);
  nand ginst7646 (P1_U4133, P1_D_REG_8__SCAN_IN, P1_U4101);
  nand ginst7647 (P1_U4134, P1_D_REG_9__SCAN_IN, P1_U4101);
  nand ginst7648 (P1_U4135, P1_U5690, P1_U5693);
  nand ginst7649 (P1_U4136, P1_U3367, P1_U5712, P1_U5713);
  nand ginst7650 (P1_U4137, P1_REG2_REG_1__SCAN_IN, P1_U3018);
  nand ginst7651 (P1_U4138, P1_REG1_REG_1__SCAN_IN, P1_U3019);
  nand ginst7652 (P1_U4139, P1_REG0_REG_1__SCAN_IN, P1_U3020);
  nand ginst7653 (P1_U4140, P1_REG3_REG_1__SCAN_IN, P1_U3017);
  not ginst7654 (P1_U4141, P1_U3078);
  nand ginst7655 (P1_U4142, P1_U3416, P1_U3966);
  nand ginst7656 (P1_U4143, P1_R1150_U18, P1_U3961);
  nand ginst7657 (P1_U4144, P1_R1117_U18, P1_U3963);
  nand ginst7658 (P1_U4145, P1_R1138_U96, P1_U3962);
  nand ginst7659 (P1_U4146, P1_R1192_U18, P1_U3959);
  nand ginst7660 (P1_U4147, P1_R1207_U18, P1_U3958);
  nand ginst7661 (P1_U4148, P1_R1171_U96, P1_U3968);
  nand ginst7662 (P1_U4149, P1_R1240_U96, P1_U3967);
  not ginst7663 (P1_U4150, P1_U3374);
  nand ginst7664 (P1_U4151, P1_R1222_U96, P1_U3026);
  nand ginst7665 (P1_U4152, P1_U3025, P1_U3078);
  nand ginst7666 (P1_U4153, P1_U3023, P1_U3450);
  nand ginst7667 (P1_U4154, P1_U3450, P1_U4142);
  nand ginst7668 (P1_U4155, P1_U3620, P1_U4150);
  nand ginst7669 (P1_U4156, P1_REG2_REG_2__SCAN_IN, P1_U3018);
  nand ginst7670 (P1_U4157, P1_REG1_REG_2__SCAN_IN, P1_U3019);
  nand ginst7671 (P1_U4158, P1_REG0_REG_2__SCAN_IN, P1_U3020);
  nand ginst7672 (P1_U4159, P1_REG3_REG_2__SCAN_IN, P1_U3017);
  not ginst7673 (P1_U4160, P1_U3068);
  nand ginst7674 (P1_U4161, P1_REG0_REG_0__SCAN_IN, P1_U3020);
  nand ginst7675 (P1_U4162, P1_REG1_REG_0__SCAN_IN, P1_U3019);
  nand ginst7676 (P1_U4163, P1_REG2_REG_0__SCAN_IN, P1_U3018);
  nand ginst7677 (P1_U4164, P1_REG3_REG_0__SCAN_IN, P1_U3017);
  not ginst7678 (P1_U4165, P1_U3077);
  nand ginst7679 (P1_U4166, P1_U3033, P1_U3077);
  nand ginst7680 (P1_U4167, P1_R1150_U96, P1_U3961);
  nand ginst7681 (P1_U4168, P1_R1117_U96, P1_U3963);
  nand ginst7682 (P1_U4169, P1_R1138_U95, P1_U3962);
  nand ginst7683 (P1_U4170, P1_R1192_U96, P1_U3959);
  nand ginst7684 (P1_U4171, P1_R1207_U96, P1_U3958);
  nand ginst7685 (P1_U4172, P1_R1171_U95, P1_U3968);
  nand ginst7686 (P1_U4173, P1_R1240_U95, P1_U3967);
  not ginst7687 (P1_U4174, P1_U3376);
  nand ginst7688 (P1_U4175, P1_R1222_U95, P1_U3026);
  nand ginst7689 (P1_U4176, P1_U3025, P1_U3068);
  nand ginst7690 (P1_U4177, P1_R1282_U57, P1_U3023);
  nand ginst7691 (P1_U4178, P1_U3455, P1_U4142);
  nand ginst7692 (P1_U4179, P1_U3636, P1_U4174);
  nand ginst7693 (P1_U4180, P1_REG2_REG_3__SCAN_IN, P1_U3018);
  nand ginst7694 (P1_U4181, P1_REG1_REG_3__SCAN_IN, P1_U3019);
  nand ginst7695 (P1_U4182, P1_REG0_REG_3__SCAN_IN, P1_U3020);
  nand ginst7696 (P1_U4183, P1_ADD_95_U4, P1_U3017);
  not ginst7697 (P1_U4184, P1_U3064);
  nand ginst7698 (P1_U4185, P1_U3033, P1_U3078);
  nand ginst7699 (P1_U4186, P1_R1150_U106, P1_U3961);
  nand ginst7700 (P1_U4187, P1_R1117_U106, P1_U3963);
  nand ginst7701 (P1_U4188, P1_R1138_U17, P1_U3962);
  nand ginst7702 (P1_U4189, P1_R1192_U106, P1_U3959);
  nand ginst7703 (P1_U4190, P1_R1207_U106, P1_U3958);
  nand ginst7704 (P1_U4191, P1_R1171_U17, P1_U3968);
  nand ginst7705 (P1_U4192, P1_R1240_U17, P1_U3967);
  not ginst7706 (P1_U4193, P1_U3377);
  nand ginst7707 (P1_U4194, P1_R1222_U17, P1_U3026);
  nand ginst7708 (P1_U4195, P1_U3025, P1_U3064);
  nand ginst7709 (P1_U4196, P1_R1282_U18, P1_U3023);
  nand ginst7710 (P1_U4197, P1_U3458, P1_U4142);
  nand ginst7711 (P1_U4198, P1_U3640, P1_U4193);
  nand ginst7712 (P1_U4199, P1_REG2_REG_4__SCAN_IN, P1_U3018);
  nand ginst7713 (P1_U4200, P1_REG1_REG_4__SCAN_IN, P1_U3019);
  nand ginst7714 (P1_U4201, P1_REG0_REG_4__SCAN_IN, P1_U3020);
  nand ginst7715 (P1_U4202, P1_ADD_95_U59, P1_U3017);
  not ginst7716 (P1_U4203, P1_U3060);
  nand ginst7717 (P1_U4204, P1_U3033, P1_U3068);
  nand ginst7718 (P1_U4205, P1_R1150_U15, P1_U3961);
  nand ginst7719 (P1_U4206, P1_R1117_U15, P1_U3963);
  nand ginst7720 (P1_U4207, P1_R1138_U101, P1_U3962);
  nand ginst7721 (P1_U4208, P1_R1192_U15, P1_U3959);
  nand ginst7722 (P1_U4209, P1_R1207_U15, P1_U3958);
  nand ginst7723 (P1_U4210, P1_R1171_U101, P1_U3968);
  nand ginst7724 (P1_U4211, P1_R1240_U101, P1_U3967);
  not ginst7725 (P1_U4212, P1_U3378);
  nand ginst7726 (P1_U4213, P1_R1222_U101, P1_U3026);
  nand ginst7727 (P1_U4214, P1_U3025, P1_U3060);
  nand ginst7728 (P1_U4215, P1_R1282_U20, P1_U3023);
  nand ginst7729 (P1_U4216, P1_U3461, P1_U4142);
  nand ginst7730 (P1_U4217, P1_U3643, P1_U4212);
  nand ginst7731 (P1_U4218, P1_REG2_REG_5__SCAN_IN, P1_U3018);
  nand ginst7732 (P1_U4219, P1_REG1_REG_5__SCAN_IN, P1_U3019);
  nand ginst7733 (P1_U4220, P1_REG0_REG_5__SCAN_IN, P1_U3020);
  nand ginst7734 (P1_U4221, P1_ADD_95_U58, P1_U3017);
  not ginst7735 (P1_U4222, P1_U3067);
  nand ginst7736 (P1_U4223, P1_U3033, P1_U3064);
  nand ginst7737 (P1_U4224, P1_R1150_U105, P1_U3961);
  nand ginst7738 (P1_U4225, P1_R1117_U105, P1_U3963);
  nand ginst7739 (P1_U4226, P1_R1138_U100, P1_U3962);
  nand ginst7740 (P1_U4227, P1_R1192_U105, P1_U3959);
  nand ginst7741 (P1_U4228, P1_R1207_U105, P1_U3958);
  nand ginst7742 (P1_U4229, P1_R1171_U100, P1_U3968);
  nand ginst7743 (P1_U4230, P1_R1240_U100, P1_U3967);
  not ginst7744 (P1_U4231, P1_U3379);
  nand ginst7745 (P1_U4232, P1_R1222_U100, P1_U3026);
  nand ginst7746 (P1_U4233, P1_U3025, P1_U3067);
  nand ginst7747 (P1_U4234, P1_R1282_U21, P1_U3023);
  nand ginst7748 (P1_U4235, P1_U3464, P1_U4142);
  nand ginst7749 (P1_U4236, P1_U3646, P1_U4231);
  nand ginst7750 (P1_U4237, P1_REG2_REG_6__SCAN_IN, P1_U3018);
  nand ginst7751 (P1_U4238, P1_REG1_REG_6__SCAN_IN, P1_U3019);
  nand ginst7752 (P1_U4239, P1_REG0_REG_6__SCAN_IN, P1_U3020);
  nand ginst7753 (P1_U4240, P1_ADD_95_U57, P1_U3017);
  not ginst7754 (P1_U4241, P1_U3071);
  nand ginst7755 (P1_U4242, P1_U3033, P1_U3060);
  nand ginst7756 (P1_U4243, P1_R1150_U104, P1_U3961);
  nand ginst7757 (P1_U4244, P1_R1117_U104, P1_U3963);
  nand ginst7758 (P1_U4245, P1_R1138_U18, P1_U3962);
  nand ginst7759 (P1_U4246, P1_R1192_U104, P1_U3959);
  nand ginst7760 (P1_U4247, P1_R1207_U104, P1_U3958);
  nand ginst7761 (P1_U4248, P1_R1171_U18, P1_U3968);
  nand ginst7762 (P1_U4249, P1_R1240_U18, P1_U3967);
  not ginst7763 (P1_U4250, P1_U3380);
  nand ginst7764 (P1_U4251, P1_R1222_U18, P1_U3026);
  nand ginst7765 (P1_U4252, P1_U3025, P1_U3071);
  nand ginst7766 (P1_U4253, P1_R1282_U65, P1_U3023);
  nand ginst7767 (P1_U4254, P1_U3467, P1_U4142);
  nand ginst7768 (P1_U4255, P1_U3650, P1_U4250);
  nand ginst7769 (P1_U4256, P1_REG2_REG_7__SCAN_IN, P1_U3018);
  nand ginst7770 (P1_U4257, P1_REG1_REG_7__SCAN_IN, P1_U3019);
  nand ginst7771 (P1_U4258, P1_REG0_REG_7__SCAN_IN, P1_U3020);
  nand ginst7772 (P1_U4259, P1_ADD_95_U56, P1_U3017);
  not ginst7773 (P1_U4260, P1_U3070);
  nand ginst7774 (P1_U4261, P1_U3033, P1_U3067);
  nand ginst7775 (P1_U4262, P1_R1150_U16, P1_U3961);
  nand ginst7776 (P1_U4263, P1_R1117_U16, P1_U3963);
  nand ginst7777 (P1_U4264, P1_R1138_U99, P1_U3962);
  nand ginst7778 (P1_U4265, P1_R1192_U16, P1_U3959);
  nand ginst7779 (P1_U4266, P1_R1207_U16, P1_U3958);
  nand ginst7780 (P1_U4267, P1_R1171_U99, P1_U3968);
  nand ginst7781 (P1_U4268, P1_R1240_U99, P1_U3967);
  not ginst7782 (P1_U4269, P1_U3381);
  nand ginst7783 (P1_U4270, P1_R1222_U99, P1_U3026);
  nand ginst7784 (P1_U4271, P1_U3025, P1_U3070);
  nand ginst7785 (P1_U4272, P1_R1282_U22, P1_U3023);
  nand ginst7786 (P1_U4273, P1_U3470, P1_U4142);
  nand ginst7787 (P1_U4274, P1_U3654, P1_U4269);
  nand ginst7788 (P1_U4275, P1_REG2_REG_8__SCAN_IN, P1_U3018);
  nand ginst7789 (P1_U4276, P1_REG1_REG_8__SCAN_IN, P1_U3019);
  nand ginst7790 (P1_U4277, P1_REG0_REG_8__SCAN_IN, P1_U3020);
  nand ginst7791 (P1_U4278, P1_ADD_95_U55, P1_U3017);
  not ginst7792 (P1_U4279, P1_U3084);
  nand ginst7793 (P1_U4280, P1_U3033, P1_U3071);
  nand ginst7794 (P1_U4281, P1_R1150_U103, P1_U3961);
  nand ginst7795 (P1_U4282, P1_R1117_U103, P1_U3963);
  nand ginst7796 (P1_U4283, P1_R1138_U19, P1_U3962);
  nand ginst7797 (P1_U4284, P1_R1192_U103, P1_U3959);
  nand ginst7798 (P1_U4285, P1_R1207_U103, P1_U3958);
  nand ginst7799 (P1_U4286, P1_R1171_U19, P1_U3968);
  nand ginst7800 (P1_U4287, P1_R1240_U19, P1_U3967);
  not ginst7801 (P1_U4288, P1_U3382);
  nand ginst7802 (P1_U4289, P1_R1222_U19, P1_U3026);
  nand ginst7803 (P1_U4290, P1_U3025, P1_U3084);
  nand ginst7804 (P1_U4291, P1_R1282_U23, P1_U3023);
  nand ginst7805 (P1_U4292, P1_U3473, P1_U4142);
  nand ginst7806 (P1_U4293, P1_U3658, P1_U4288);
  nand ginst7807 (P1_U4294, P1_REG2_REG_9__SCAN_IN, P1_U3018);
  nand ginst7808 (P1_U4295, P1_REG1_REG_9__SCAN_IN, P1_U3019);
  nand ginst7809 (P1_U4296, P1_REG0_REG_9__SCAN_IN, P1_U3020);
  nand ginst7810 (P1_U4297, P1_ADD_95_U54, P1_U3017);
  not ginst7811 (P1_U4298, P1_U3083);
  nand ginst7812 (P1_U4299, P1_U3033, P1_U3070);
  nand ginst7813 (P1_U4300, P1_R1150_U17, P1_U3961);
  nand ginst7814 (P1_U4301, P1_R1117_U17, P1_U3963);
  nand ginst7815 (P1_U4302, P1_R1138_U98, P1_U3962);
  nand ginst7816 (P1_U4303, P1_R1192_U17, P1_U3959);
  nand ginst7817 (P1_U4304, P1_R1207_U17, P1_U3958);
  nand ginst7818 (P1_U4305, P1_R1171_U98, P1_U3968);
  nand ginst7819 (P1_U4306, P1_R1240_U98, P1_U3967);
  not ginst7820 (P1_U4307, P1_U3383);
  nand ginst7821 (P1_U4308, P1_R1222_U98, P1_U3026);
  nand ginst7822 (P1_U4309, P1_U3025, P1_U3083);
  nand ginst7823 (P1_U4310, P1_R1282_U24, P1_U3023);
  nand ginst7824 (P1_U4311, P1_U3476, P1_U4142);
  nand ginst7825 (P1_U4312, P1_U3662, P1_U4307);
  nand ginst7826 (P1_U4313, P1_REG2_REG_10__SCAN_IN, P1_U3018);
  nand ginst7827 (P1_U4314, P1_REG1_REG_10__SCAN_IN, P1_U3019);
  nand ginst7828 (P1_U4315, P1_REG0_REG_10__SCAN_IN, P1_U3020);
  nand ginst7829 (P1_U4316, P1_ADD_95_U78, P1_U3017);
  not ginst7830 (P1_U4317, P1_U3062);
  nand ginst7831 (P1_U4318, P1_U3033, P1_U3084);
  nand ginst7832 (P1_U4319, P1_R1150_U102, P1_U3961);
  nand ginst7833 (P1_U4320, P1_R1117_U102, P1_U3963);
  nand ginst7834 (P1_U4321, P1_R1138_U97, P1_U3962);
  nand ginst7835 (P1_U4322, P1_R1192_U102, P1_U3959);
  nand ginst7836 (P1_U4323, P1_R1207_U102, P1_U3958);
  nand ginst7837 (P1_U4324, P1_R1171_U97, P1_U3968);
  nand ginst7838 (P1_U4325, P1_R1240_U97, P1_U3967);
  not ginst7839 (P1_U4326, P1_U3384);
  nand ginst7840 (P1_U4327, P1_R1222_U97, P1_U3026);
  nand ginst7841 (P1_U4328, P1_U3025, P1_U3062);
  nand ginst7842 (P1_U4329, P1_R1282_U63, P1_U3023);
  nand ginst7843 (P1_U4330, P1_U3479, P1_U4142);
  nand ginst7844 (P1_U4331, P1_U3666, P1_U4326);
  nand ginst7845 (P1_U4332, P1_REG2_REG_11__SCAN_IN, P1_U3018);
  nand ginst7846 (P1_U4333, P1_REG1_REG_11__SCAN_IN, P1_U3019);
  nand ginst7847 (P1_U4334, P1_REG0_REG_11__SCAN_IN, P1_U3020);
  nand ginst7848 (P1_U4335, P1_ADD_95_U77, P1_U3017);
  not ginst7849 (P1_U4336, P1_U3063);
  nand ginst7850 (P1_U4337, P1_U3033, P1_U3083);
  nand ginst7851 (P1_U4338, P1_R1150_U112, P1_U3961);
  nand ginst7852 (P1_U4339, P1_R1117_U112, P1_U3963);
  nand ginst7853 (P1_U4340, P1_R1138_U11, P1_U3962);
  nand ginst7854 (P1_U4341, P1_R1192_U112, P1_U3959);
  nand ginst7855 (P1_U4342, P1_R1207_U112, P1_U3958);
  nand ginst7856 (P1_U4343, P1_R1171_U11, P1_U3968);
  nand ginst7857 (P1_U4344, P1_R1240_U11, P1_U3967);
  not ginst7858 (P1_U4345, P1_U3385);
  nand ginst7859 (P1_U4346, P1_R1222_U11, P1_U3026);
  nand ginst7860 (P1_U4347, P1_U3025, P1_U3063);
  nand ginst7861 (P1_U4348, P1_R1282_U6, P1_U3023);
  nand ginst7862 (P1_U4349, P1_U3482, P1_U4142);
  nand ginst7863 (P1_U4350, P1_U3670, P1_U4345);
  nand ginst7864 (P1_U4351, P1_REG2_REG_12__SCAN_IN, P1_U3018);
  nand ginst7865 (P1_U4352, P1_REG1_REG_12__SCAN_IN, P1_U3019);
  nand ginst7866 (P1_U4353, P1_REG0_REG_12__SCAN_IN, P1_U3020);
  nand ginst7867 (P1_U4354, P1_ADD_95_U76, P1_U3017);
  not ginst7868 (P1_U4355, P1_U3072);
  nand ginst7869 (P1_U4356, P1_U3033, P1_U3062);
  nand ginst7870 (P1_U4357, P1_R1150_U10, P1_U3961);
  nand ginst7871 (P1_U4358, P1_R1117_U10, P1_U3963);
  nand ginst7872 (P1_U4359, P1_R1138_U115, P1_U3962);
  nand ginst7873 (P1_U4360, P1_R1192_U10, P1_U3959);
  nand ginst7874 (P1_U4361, P1_R1207_U10, P1_U3958);
  nand ginst7875 (P1_U4362, P1_R1171_U115, P1_U3968);
  nand ginst7876 (P1_U4363, P1_R1240_U115, P1_U3967);
  not ginst7877 (P1_U4364, P1_U3386);
  nand ginst7878 (P1_U4365, P1_R1222_U115, P1_U3026);
  nand ginst7879 (P1_U4366, P1_U3025, P1_U3072);
  nand ginst7880 (P1_U4367, P1_R1282_U7, P1_U3023);
  nand ginst7881 (P1_U4368, P1_U3485, P1_U4142);
  nand ginst7882 (P1_U4369, P1_U3674, P1_U4364);
  nand ginst7883 (P1_U4370, P1_REG2_REG_13__SCAN_IN, P1_U3018);
  nand ginst7884 (P1_U4371, P1_REG1_REG_13__SCAN_IN, P1_U3019);
  nand ginst7885 (P1_U4372, P1_REG0_REG_13__SCAN_IN, P1_U3020);
  nand ginst7886 (P1_U4373, P1_ADD_95_U75, P1_U3017);
  not ginst7887 (P1_U4374, P1_U3080);
  nand ginst7888 (P1_U4375, P1_U3033, P1_U3063);
  nand ginst7889 (P1_U4376, P1_R1150_U101, P1_U3961);
  nand ginst7890 (P1_U4377, P1_R1117_U101, P1_U3963);
  nand ginst7891 (P1_U4378, P1_R1138_U114, P1_U3962);
  nand ginst7892 (P1_U4379, P1_R1192_U101, P1_U3959);
  nand ginst7893 (P1_U4380, P1_R1207_U101, P1_U3958);
  nand ginst7894 (P1_U4381, P1_R1171_U114, P1_U3968);
  nand ginst7895 (P1_U4382, P1_R1240_U114, P1_U3967);
  not ginst7896 (P1_U4383, P1_U3387);
  nand ginst7897 (P1_U4384, P1_R1222_U114, P1_U3026);
  nand ginst7898 (P1_U4385, P1_U3025, P1_U3080);
  nand ginst7899 (P1_U4386, P1_R1282_U8, P1_U3023);
  nand ginst7900 (P1_U4387, P1_U3488, P1_U4142);
  nand ginst7901 (P1_U4388, P1_U3678, P1_U4383);
  nand ginst7902 (P1_U4389, P1_REG2_REG_14__SCAN_IN, P1_U3018);
  nand ginst7903 (P1_U4390, P1_REG1_REG_14__SCAN_IN, P1_U3019);
  nand ginst7904 (P1_U4391, P1_REG0_REG_14__SCAN_IN, P1_U3020);
  nand ginst7905 (P1_U4392, P1_ADD_95_U74, P1_U3017);
  not ginst7906 (P1_U4393, P1_U3079);
  nand ginst7907 (P1_U4394, P1_U3033, P1_U3072);
  nand ginst7908 (P1_U4395, P1_R1150_U100, P1_U3961);
  nand ginst7909 (P1_U4396, P1_R1117_U100, P1_U3963);
  nand ginst7910 (P1_U4397, P1_R1138_U12, P1_U3962);
  nand ginst7911 (P1_U4398, P1_R1192_U100, P1_U3959);
  nand ginst7912 (P1_U4399, P1_R1207_U100, P1_U3958);
  nand ginst7913 (P1_U4400, P1_R1171_U12, P1_U3968);
  nand ginst7914 (P1_U4401, P1_R1240_U12, P1_U3967);
  not ginst7915 (P1_U4402, P1_U3388);
  nand ginst7916 (P1_U4403, P1_R1222_U12, P1_U3026);
  nand ginst7917 (P1_U4404, P1_U3025, P1_U3079);
  nand ginst7918 (P1_U4405, P1_R1282_U86, P1_U3023);
  nand ginst7919 (P1_U4406, P1_U3491, P1_U4142);
  nand ginst7920 (P1_U4407, P1_U3682, P1_U4402);
  nand ginst7921 (P1_U4408, P1_REG2_REG_15__SCAN_IN, P1_U3018);
  nand ginst7922 (P1_U4409, P1_REG1_REG_15__SCAN_IN, P1_U3019);
  nand ginst7923 (P1_U4410, P1_REG0_REG_15__SCAN_IN, P1_U3020);
  nand ginst7924 (P1_U4411, P1_ADD_95_U73, P1_U3017);
  not ginst7925 (P1_U4412, P1_U3074);
  nand ginst7926 (P1_U4413, P1_U3033, P1_U3080);
  nand ginst7927 (P1_U4414, P1_R1150_U111, P1_U3961);
  nand ginst7928 (P1_U4415, P1_R1117_U111, P1_U3963);
  nand ginst7929 (P1_U4416, P1_R1138_U113, P1_U3962);
  nand ginst7930 (P1_U4417, P1_R1192_U111, P1_U3959);
  nand ginst7931 (P1_U4418, P1_R1207_U111, P1_U3958);
  nand ginst7932 (P1_U4419, P1_R1171_U113, P1_U3968);
  nand ginst7933 (P1_U4420, P1_R1240_U113, P1_U3967);
  not ginst7934 (P1_U4421, P1_U3389);
  nand ginst7935 (P1_U4422, P1_R1222_U113, P1_U3026);
  nand ginst7936 (P1_U4423, P1_U3025, P1_U3074);
  nand ginst7937 (P1_U4424, P1_R1282_U9, P1_U3023);
  nand ginst7938 (P1_U4425, P1_U3494, P1_U4142);
  nand ginst7939 (P1_U4426, P1_U3686, P1_U4421);
  nand ginst7940 (P1_U4427, P1_REG2_REG_16__SCAN_IN, P1_U3018);
  nand ginst7941 (P1_U4428, P1_REG1_REG_16__SCAN_IN, P1_U3019);
  nand ginst7942 (P1_U4429, P1_REG0_REG_16__SCAN_IN, P1_U3020);
  nand ginst7943 (P1_U4430, P1_ADD_95_U72, P1_U3017);
  not ginst7944 (P1_U4431, P1_U3073);
  nand ginst7945 (P1_U4432, P1_U3033, P1_U3079);
  nand ginst7946 (P1_U4433, P1_R1150_U110, P1_U3961);
  nand ginst7947 (P1_U4434, P1_R1117_U110, P1_U3963);
  nand ginst7948 (P1_U4435, P1_R1138_U112, P1_U3962);
  nand ginst7949 (P1_U4436, P1_R1192_U110, P1_U3959);
  nand ginst7950 (P1_U4437, P1_R1207_U110, P1_U3958);
  nand ginst7951 (P1_U4438, P1_R1171_U112, P1_U3968);
  nand ginst7952 (P1_U4439, P1_R1240_U112, P1_U3967);
  not ginst7953 (P1_U4440, P1_U3390);
  nand ginst7954 (P1_U4441, P1_R1222_U112, P1_U3026);
  nand ginst7955 (P1_U4442, P1_U3025, P1_U3073);
  nand ginst7956 (P1_U4443, P1_R1282_U10, P1_U3023);
  nand ginst7957 (P1_U4444, P1_U3497, P1_U4142);
  nand ginst7958 (P1_U4445, P1_U3690, P1_U4440);
  nand ginst7959 (P1_U4446, P1_REG2_REG_17__SCAN_IN, P1_U3018);
  nand ginst7960 (P1_U4447, P1_REG1_REG_17__SCAN_IN, P1_U3019);
  nand ginst7961 (P1_U4448, P1_REG0_REG_17__SCAN_IN, P1_U3020);
  nand ginst7962 (P1_U4449, P1_ADD_95_U71, P1_U3017);
  not ginst7963 (P1_U4450, P1_U3069);
  nand ginst7964 (P1_U4451, P1_U3033, P1_U3074);
  nand ginst7965 (P1_U4452, P1_R1150_U11, P1_U3961);
  nand ginst7966 (P1_U4453, P1_R1117_U11, P1_U3963);
  nand ginst7967 (P1_U4454, P1_R1138_U111, P1_U3962);
  nand ginst7968 (P1_U4455, P1_R1192_U11, P1_U3959);
  nand ginst7969 (P1_U4456, P1_R1207_U11, P1_U3958);
  nand ginst7970 (P1_U4457, P1_R1171_U111, P1_U3968);
  nand ginst7971 (P1_U4458, P1_R1240_U111, P1_U3967);
  not ginst7972 (P1_U4459, P1_U3391);
  nand ginst7973 (P1_U4460, P1_R1222_U111, P1_U3026);
  nand ginst7974 (P1_U4461, P1_U3025, P1_U3069);
  nand ginst7975 (P1_U4462, P1_R1282_U11, P1_U3023);
  nand ginst7976 (P1_U4463, P1_U3500, P1_U4142);
  nand ginst7977 (P1_U4464, P1_U3694, P1_U4459);
  nand ginst7978 (P1_U4465, P1_REG2_REG_18__SCAN_IN, P1_U3018);
  nand ginst7979 (P1_U4466, P1_REG1_REG_18__SCAN_IN, P1_U3019);
  nand ginst7980 (P1_U4467, P1_REG0_REG_18__SCAN_IN, P1_U3020);
  nand ginst7981 (P1_U4468, P1_ADD_95_U70, P1_U3017);
  not ginst7982 (P1_U4469, P1_U3082);
  nand ginst7983 (P1_U4470, P1_U3033, P1_U3073);
  nand ginst7984 (P1_U4471, P1_R1150_U99, P1_U3961);
  nand ginst7985 (P1_U4472, P1_R1117_U99, P1_U3963);
  nand ginst7986 (P1_U4473, P1_R1138_U13, P1_U3962);
  nand ginst7987 (P1_U4474, P1_R1192_U99, P1_U3959);
  nand ginst7988 (P1_U4475, P1_R1207_U99, P1_U3958);
  nand ginst7989 (P1_U4476, P1_R1171_U13, P1_U3968);
  nand ginst7990 (P1_U4477, P1_R1240_U13, P1_U3967);
  not ginst7991 (P1_U4478, P1_U3392);
  nand ginst7992 (P1_U4479, P1_R1222_U13, P1_U3026);
  nand ginst7993 (P1_U4480, P1_U3025, P1_U3082);
  nand ginst7994 (P1_U4481, P1_R1282_U84, P1_U3023);
  nand ginst7995 (P1_U4482, P1_U3503, P1_U4142);
  nand ginst7996 (P1_U4483, P1_U3698, P1_U4478);
  nand ginst7997 (P1_U4484, P1_REG2_REG_19__SCAN_IN, P1_U3018);
  nand ginst7998 (P1_U4485, P1_REG1_REG_19__SCAN_IN, P1_U3019);
  nand ginst7999 (P1_U4486, P1_REG0_REG_19__SCAN_IN, P1_U3020);
  nand ginst8000 (P1_U4487, P1_ADD_95_U69, P1_U3017);
  not ginst8001 (P1_U4488, P1_U3081);
  nand ginst8002 (P1_U4489, P1_U3033, P1_U3069);
  nand ginst8003 (P1_U4490, P1_R1150_U98, P1_U3961);
  nand ginst8004 (P1_U4491, P1_R1117_U98, P1_U3963);
  nand ginst8005 (P1_U4492, P1_R1138_U110, P1_U3962);
  nand ginst8006 (P1_U4493, P1_R1192_U98, P1_U3959);
  nand ginst8007 (P1_U4494, P1_R1207_U98, P1_U3958);
  nand ginst8008 (P1_U4495, P1_R1171_U110, P1_U3968);
  nand ginst8009 (P1_U4496, P1_R1240_U110, P1_U3967);
  not ginst8010 (P1_U4497, P1_U3393);
  nand ginst8011 (P1_U4498, P1_R1222_U110, P1_U3026);
  nand ginst8012 (P1_U4499, P1_U3025, P1_U3081);
  nand ginst8013 (P1_U4500, P1_R1282_U12, P1_U3023);
  nand ginst8014 (P1_U4501, P1_U3506, P1_U4142);
  nand ginst8015 (P1_U4502, P1_U3702, P1_U4497);
  nand ginst8016 (P1_U4503, P1_REG2_REG_20__SCAN_IN, P1_U3018);
  nand ginst8017 (P1_U4504, P1_REG1_REG_20__SCAN_IN, P1_U3019);
  nand ginst8018 (P1_U4505, P1_REG0_REG_20__SCAN_IN, P1_U3020);
  nand ginst8019 (P1_U4506, P1_ADD_95_U68, P1_U3017);
  not ginst8020 (P1_U4507, P1_U3076);
  nand ginst8021 (P1_U4508, P1_U3033, P1_U3082);
  nand ginst8022 (P1_U4509, P1_R1150_U97, P1_U3961);
  nand ginst8023 (P1_U4510, P1_R1117_U97, P1_U3963);
  nand ginst8024 (P1_U4511, P1_R1138_U109, P1_U3962);
  nand ginst8025 (P1_U4512, P1_R1192_U97, P1_U3959);
  nand ginst8026 (P1_U4513, P1_R1207_U97, P1_U3958);
  nand ginst8027 (P1_U4514, P1_R1171_U109, P1_U3968);
  nand ginst8028 (P1_U4515, P1_R1240_U109, P1_U3967);
  not ginst8029 (P1_U4516, P1_U3394);
  nand ginst8030 (P1_U4517, P1_R1222_U109, P1_U3026);
  nand ginst8031 (P1_U4518, P1_U3025, P1_U3076);
  nand ginst8032 (P1_U4519, P1_R1282_U82, P1_U3023);
  nand ginst8033 (P1_U4520, P1_U3508, P1_U4142);
  nand ginst8034 (P1_U4521, P1_U3706, P1_U4516);
  nand ginst8035 (P1_U4522, P1_REG2_REG_21__SCAN_IN, P1_U3018);
  nand ginst8036 (P1_U4523, P1_REG1_REG_21__SCAN_IN, P1_U3019);
  nand ginst8037 (P1_U4524, P1_REG0_REG_21__SCAN_IN, P1_U3020);
  nand ginst8038 (P1_U4525, P1_ADD_95_U67, P1_U3017);
  not ginst8039 (P1_U4526, P1_U3075);
  nand ginst8040 (P1_U4527, P1_U3033, P1_U3081);
  nand ginst8041 (P1_U4528, P1_R1150_U95, P1_U3961);
  nand ginst8042 (P1_U4529, P1_R1117_U95, P1_U3963);
  nand ginst8043 (P1_U4530, P1_R1138_U14, P1_U3962);
  nand ginst8044 (P1_U4531, P1_R1192_U95, P1_U3959);
  nand ginst8045 (P1_U4532, P1_R1207_U95, P1_U3958);
  nand ginst8046 (P1_U4533, P1_R1171_U14, P1_U3968);
  nand ginst8047 (P1_U4534, P1_R1240_U14, P1_U3967);
  not ginst8048 (P1_U4535, P1_U3396);
  nand ginst8049 (P1_U4536, P1_R1222_U14, P1_U3026);
  nand ginst8050 (P1_U4537, P1_U3025, P1_U3075);
  nand ginst8051 (P1_U4538, P1_R1282_U13, P1_U3023);
  nand ginst8052 (P1_U4539, P1_U3982, P1_U4142);
  nand ginst8053 (P1_U4540, P1_U3710, P1_U4535);
  nand ginst8054 (P1_U4541, P1_REG2_REG_22__SCAN_IN, P1_U3018);
  nand ginst8055 (P1_U4542, P1_REG1_REG_22__SCAN_IN, P1_U3019);
  nand ginst8056 (P1_U4543, P1_REG0_REG_22__SCAN_IN, P1_U3020);
  nand ginst8057 (P1_U4544, P1_ADD_95_U66, P1_U3017);
  not ginst8058 (P1_U4545, P1_U3061);
  nand ginst8059 (P1_U4546, P1_U3033, P1_U3076);
  nand ginst8060 (P1_U4547, P1_R1150_U109, P1_U3961);
  nand ginst8061 (P1_U4548, P1_R1117_U109, P1_U3963);
  nand ginst8062 (P1_U4549, P1_R1138_U15, P1_U3962);
  nand ginst8063 (P1_U4550, P1_R1192_U109, P1_U3959);
  nand ginst8064 (P1_U4551, P1_R1207_U109, P1_U3958);
  nand ginst8065 (P1_U4552, P1_R1171_U15, P1_U3968);
  nand ginst8066 (P1_U4553, P1_R1240_U15, P1_U3967);
  not ginst8067 (P1_U4554, P1_U3398);
  nand ginst8068 (P1_U4555, P1_R1222_U15, P1_U3026);
  nand ginst8069 (P1_U4556, P1_U3025, P1_U3061);
  nand ginst8070 (P1_U4557, P1_R1282_U78, P1_U3023);
  nand ginst8071 (P1_U4558, P1_U3981, P1_U4142);
  nand ginst8072 (P1_U4559, P1_U3714, P1_U4554);
  nand ginst8073 (P1_U4560, P1_REG2_REG_23__SCAN_IN, P1_U3018);
  nand ginst8074 (P1_U4561, P1_REG1_REG_23__SCAN_IN, P1_U3019);
  nand ginst8075 (P1_U4562, P1_REG0_REG_23__SCAN_IN, P1_U3020);
  nand ginst8076 (P1_U4563, P1_ADD_95_U65, P1_U3017);
  not ginst8077 (P1_U4564, P1_U3066);
  nand ginst8078 (P1_U4565, P1_U3033, P1_U3075);
  nand ginst8079 (P1_U4566, P1_R1150_U108, P1_U3961);
  nand ginst8080 (P1_U4567, P1_R1117_U108, P1_U3963);
  nand ginst8081 (P1_U4568, P1_R1138_U108, P1_U3962);
  nand ginst8082 (P1_U4569, P1_R1192_U108, P1_U3959);
  nand ginst8083 (P1_U4570, P1_R1207_U108, P1_U3958);
  nand ginst8084 (P1_U4571, P1_R1171_U108, P1_U3968);
  nand ginst8085 (P1_U4572, P1_R1240_U108, P1_U3967);
  not ginst8086 (P1_U4573, P1_U3400);
  nand ginst8087 (P1_U4574, P1_R1222_U108, P1_U3026);
  nand ginst8088 (P1_U4575, P1_U3025, P1_U3066);
  nand ginst8089 (P1_U4576, P1_R1282_U14, P1_U3023);
  nand ginst8090 (P1_U4577, P1_U3980, P1_U4142);
  nand ginst8091 (P1_U4578, P1_U3718, P1_U4573);
  nand ginst8092 (P1_U4579, P1_REG2_REG_24__SCAN_IN, P1_U3018);
  nand ginst8093 (P1_U4580, P1_REG1_REG_24__SCAN_IN, P1_U3019);
  nand ginst8094 (P1_U4581, P1_REG0_REG_24__SCAN_IN, P1_U3020);
  nand ginst8095 (P1_U4582, P1_ADD_95_U64, P1_U3017);
  not ginst8096 (P1_U4583, P1_U3065);
  nand ginst8097 (P1_U4584, P1_U3033, P1_U3061);
  nand ginst8098 (P1_U4585, P1_R1150_U12, P1_U3961);
  nand ginst8099 (P1_U4586, P1_R1117_U12, P1_U3963);
  nand ginst8100 (P1_U4587, P1_R1138_U107, P1_U3962);
  nand ginst8101 (P1_U4588, P1_R1192_U12, P1_U3959);
  nand ginst8102 (P1_U4589, P1_R1207_U12, P1_U3958);
  nand ginst8103 (P1_U4590, P1_R1171_U107, P1_U3968);
  nand ginst8104 (P1_U4591, P1_R1240_U107, P1_U3967);
  not ginst8105 (P1_U4592, P1_U3402);
  nand ginst8106 (P1_U4593, P1_R1222_U107, P1_U3026);
  nand ginst8107 (P1_U4594, P1_U3025, P1_U3065);
  nand ginst8108 (P1_U4595, P1_R1282_U76, P1_U3023);
  nand ginst8109 (P1_U4596, P1_U3979, P1_U4142);
  nand ginst8110 (P1_U4597, P1_U3722, P1_U4592);
  nand ginst8111 (P1_U4598, P1_REG2_REG_25__SCAN_IN, P1_U3018);
  nand ginst8112 (P1_U4599, P1_REG1_REG_25__SCAN_IN, P1_U3019);
  nand ginst8113 (P1_U4600, P1_REG0_REG_25__SCAN_IN, P1_U3020);
  nand ginst8114 (P1_U4601, P1_ADD_95_U63, P1_U3017);
  not ginst8115 (P1_U4602, P1_U3058);
  nand ginst8116 (P1_U4603, P1_U3033, P1_U3066);
  nand ginst8117 (P1_U4604, P1_R1150_U94, P1_U3961);
  nand ginst8118 (P1_U4605, P1_R1117_U94, P1_U3963);
  nand ginst8119 (P1_U4606, P1_R1138_U106, P1_U3962);
  nand ginst8120 (P1_U4607, P1_R1192_U94, P1_U3959);
  nand ginst8121 (P1_U4608, P1_R1207_U94, P1_U3958);
  nand ginst8122 (P1_U4609, P1_R1171_U106, P1_U3968);
  nand ginst8123 (P1_U4610, P1_R1240_U106, P1_U3967);
  not ginst8124 (P1_U4611, P1_U3404);
  nand ginst8125 (P1_U4612, P1_R1222_U106, P1_U3026);
  nand ginst8126 (P1_U4613, P1_U3025, P1_U3058);
  nand ginst8127 (P1_U4614, P1_R1282_U15, P1_U3023);
  nand ginst8128 (P1_U4615, P1_U3978, P1_U4142);
  nand ginst8129 (P1_U4616, P1_U3726, P1_U4611);
  nand ginst8130 (P1_U4617, P1_REG2_REG_26__SCAN_IN, P1_U3018);
  nand ginst8131 (P1_U4618, P1_REG1_REG_26__SCAN_IN, P1_U3019);
  nand ginst8132 (P1_U4619, P1_REG0_REG_26__SCAN_IN, P1_U3020);
  nand ginst8133 (P1_U4620, P1_ADD_95_U62, P1_U3017);
  not ginst8134 (P1_U4621, P1_U3057);
  nand ginst8135 (P1_U4622, P1_U3033, P1_U3065);
  nand ginst8136 (P1_U4623, P1_R1150_U93, P1_U3961);
  nand ginst8137 (P1_U4624, P1_R1117_U93, P1_U3963);
  nand ginst8138 (P1_U4625, P1_R1138_U105, P1_U3962);
  nand ginst8139 (P1_U4626, P1_R1192_U93, P1_U3959);
  nand ginst8140 (P1_U4627, P1_R1207_U93, P1_U3958);
  nand ginst8141 (P1_U4628, P1_R1171_U105, P1_U3968);
  nand ginst8142 (P1_U4629, P1_R1240_U105, P1_U3967);
  not ginst8143 (P1_U4630, P1_U3406);
  nand ginst8144 (P1_U4631, P1_R1222_U105, P1_U3026);
  nand ginst8145 (P1_U4632, P1_U3025, P1_U3057);
  nand ginst8146 (P1_U4633, P1_R1282_U74, P1_U3023);
  nand ginst8147 (P1_U4634, P1_U3977, P1_U4142);
  nand ginst8148 (P1_U4635, P1_U3730, P1_U4630);
  nand ginst8149 (P1_U4636, P1_REG2_REG_27__SCAN_IN, P1_U3018);
  nand ginst8150 (P1_U4637, P1_REG1_REG_27__SCAN_IN, P1_U3019);
  nand ginst8151 (P1_U4638, P1_REG0_REG_27__SCAN_IN, P1_U3020);
  nand ginst8152 (P1_U4639, P1_ADD_95_U61, P1_U3017);
  not ginst8153 (P1_U4640, P1_U3053);
  nand ginst8154 (P1_U4641, P1_U3033, P1_U3058);
  nand ginst8155 (P1_U4642, P1_R1150_U107, P1_U3961);
  nand ginst8156 (P1_U4643, P1_R1117_U107, P1_U3963);
  nand ginst8157 (P1_U4644, P1_R1138_U16, P1_U3962);
  nand ginst8158 (P1_U4645, P1_R1192_U107, P1_U3959);
  nand ginst8159 (P1_U4646, P1_R1207_U107, P1_U3958);
  nand ginst8160 (P1_U4647, P1_R1171_U16, P1_U3968);
  nand ginst8161 (P1_U4648, P1_R1240_U16, P1_U3967);
  not ginst8162 (P1_U4649, P1_U3408);
  nand ginst8163 (P1_U4650, P1_R1222_U16, P1_U3026);
  nand ginst8164 (P1_U4651, P1_U3025, P1_U3053);
  nand ginst8165 (P1_U4652, P1_R1282_U16, P1_U3023);
  nand ginst8166 (P1_U4653, P1_U3976, P1_U4142);
  nand ginst8167 (P1_U4654, P1_U3734, P1_U4649);
  nand ginst8168 (P1_U4655, P1_REG2_REG_28__SCAN_IN, P1_U3018);
  nand ginst8169 (P1_U4656, P1_REG1_REG_28__SCAN_IN, P1_U3019);
  nand ginst8170 (P1_U4657, P1_REG0_REG_28__SCAN_IN, P1_U3020);
  nand ginst8171 (P1_U4658, P1_ADD_95_U60, P1_U3017);
  not ginst8172 (P1_U4659, P1_U3054);
  nand ginst8173 (P1_U4660, P1_U3033, P1_U3057);
  nand ginst8174 (P1_U4661, P1_R1150_U13, P1_U3961);
  nand ginst8175 (P1_U4662, P1_R1117_U13, P1_U3963);
  nand ginst8176 (P1_U4663, P1_R1138_U104, P1_U3962);
  nand ginst8177 (P1_U4664, P1_R1192_U13, P1_U3959);
  nand ginst8178 (P1_U4665, P1_R1207_U13, P1_U3958);
  nand ginst8179 (P1_U4666, P1_R1171_U104, P1_U3968);
  nand ginst8180 (P1_U4667, P1_R1240_U104, P1_U3967);
  not ginst8181 (P1_U4668, P1_U3410);
  nand ginst8182 (P1_U4669, P1_R1222_U104, P1_U3026);
  nand ginst8183 (P1_U4670, P1_U3025, P1_U3054);
  nand ginst8184 (P1_U4671, P1_R1282_U72, P1_U3023);
  nand ginst8185 (P1_U4672, P1_U3975, P1_U4142);
  nand ginst8186 (P1_U4673, P1_U3738, P1_U4668);
  nand ginst8187 (P1_U4674, P1_ADD_95_U5, P1_U3017);
  nand ginst8188 (P1_U4675, P1_REG2_REG_29__SCAN_IN, P1_U3018);
  nand ginst8189 (P1_U4676, P1_REG1_REG_29__SCAN_IN, P1_U3019);
  nand ginst8190 (P1_U4677, P1_REG0_REG_29__SCAN_IN, P1_U3020);
  not ginst8191 (P1_U4678, P1_U3055);
  nand ginst8192 (P1_U4679, P1_U3033, P1_U3053);
  nand ginst8193 (P1_U4680, P1_R1150_U92, P1_U3961);
  nand ginst8194 (P1_U4681, P1_R1117_U92, P1_U3963);
  nand ginst8195 (P1_U4682, P1_R1138_U103, P1_U3962);
  nand ginst8196 (P1_U4683, P1_R1192_U92, P1_U3959);
  nand ginst8197 (P1_U4684, P1_R1207_U92, P1_U3958);
  nand ginst8198 (P1_U4685, P1_R1171_U103, P1_U3968);
  nand ginst8199 (P1_U4686, P1_R1240_U103, P1_U3967);
  not ginst8200 (P1_U4687, P1_U3412);
  nand ginst8201 (P1_U4688, P1_R1222_U103, P1_U3026);
  nand ginst8202 (P1_U4689, P1_U3025, P1_U3055);
  nand ginst8203 (P1_U4690, P1_R1282_U17, P1_U3023);
  nand ginst8204 (P1_U4691, P1_U3974, P1_U4142);
  nand ginst8205 (P1_U4692, P1_U3742, P1_U4687);
  nand ginst8206 (P1_U4693, P1_REG2_REG_30__SCAN_IN, P1_U3018);
  nand ginst8207 (P1_U4694, P1_REG1_REG_30__SCAN_IN, P1_U3019);
  nand ginst8208 (P1_U4695, P1_REG0_REG_30__SCAN_IN, P1_U3020);
  not ginst8209 (P1_U4696, P1_U3059);
  nand ginst8210 (P1_U4697, P1_U3359, P1_U5699);
  nand ginst8211 (P1_U4698, P1_U3912, P1_U4697);
  nand ginst8212 (P1_U4699, P1_U3059, P1_U3743);
  nand ginst8213 (P1_U4700, P1_U3033, P1_U3054);
  nand ginst8214 (P1_U4701, P1_R1150_U14, P1_U3961);
  nand ginst8215 (P1_U4702, P1_R1117_U14, P1_U3963);
  nand ginst8216 (P1_U4703, P1_R1138_U102, P1_U3962);
  nand ginst8217 (P1_U4704, P1_R1192_U14, P1_U3959);
  nand ginst8218 (P1_U4705, P1_R1207_U14, P1_U3958);
  nand ginst8219 (P1_U4706, P1_R1171_U102, P1_U3968);
  nand ginst8220 (P1_U4707, P1_R1240_U102, P1_U3967);
  nand ginst8221 (P1_U4708, P1_U3051, P1_U3801, P1_U3802);
  nand ginst8222 (P1_U4709, P1_R1222_U102, P1_U3026);
  nand ginst8223 (P1_U4710, P1_R1282_U70, P1_U3023);
  nand ginst8224 (P1_U4711, P1_U3985, P1_U4142);
  nand ginst8225 (P1_U4712, P1_U3051, P1_U3744, P1_U3745, P1_U3746);
  nand ginst8226 (P1_U4713, P1_REG2_REG_31__SCAN_IN, P1_U3018);
  nand ginst8227 (P1_U4714, P1_REG1_REG_31__SCAN_IN, P1_U3019);
  nand ginst8228 (P1_U4715, P1_REG0_REG_31__SCAN_IN, P1_U3020);
  not ginst8229 (P1_U4716, P1_U3056);
  nand ginst8230 (P1_U4717, P1_R1282_U19, P1_U3023);
  nand ginst8231 (P1_U4718, P1_U3984, P1_U4142);
  nand ginst8232 (P1_U4719, P1_U3945, P1_U4717, P1_U4718);
  nand ginst8233 (P1_U4720, P1_R1282_U68, P1_U3023);
  nand ginst8234 (P1_U4721, P1_U3983, P1_U4142);
  nand ginst8235 (P1_U4722, P1_U3945, P1_U4720, P1_U4721);
  nand ginst8236 (P1_U4723, P1_U3016, P1_U3749);
  nand ginst8237 (P1_U4724, P1_U3418, P1_U4723);
  nand ginst8238 (P1_U4725, P1_U3441, P1_U3988);
  not ginst8239 (P1_U4726, P1_U3422);
  nand ginst8240 (P1_U4727, P1_U3035, P1_U3078);
  nand ginst8241 (P1_U4728, P1_REG3_REG_0__SCAN_IN, P1_U3032);
  nand ginst8242 (P1_U4729, P1_R1222_U96, P1_U3031);
  nand ginst8243 (P1_U4730, P1_U3030, P1_U3450);
  nand ginst8244 (P1_U4731, P1_U3029, P1_U3450);
  nand ginst8245 (P1_U4732, P1_U3035, P1_U3068);
  nand ginst8246 (P1_U4733, P1_REG3_REG_1__SCAN_IN, P1_U3032);
  nand ginst8247 (P1_U4734, P1_R1222_U95, P1_U3031);
  nand ginst8248 (P1_U4735, P1_U3030, P1_U3455);
  nand ginst8249 (P1_U4736, P1_R1282_U57, P1_U3029);
  nand ginst8250 (P1_U4737, P1_U3035, P1_U3064);
  nand ginst8251 (P1_U4738, P1_REG3_REG_2__SCAN_IN, P1_U3032);
  nand ginst8252 (P1_U4739, P1_R1222_U17, P1_U3031);
  nand ginst8253 (P1_U4740, P1_U3030, P1_U3458);
  nand ginst8254 (P1_U4741, P1_R1282_U18, P1_U3029);
  nand ginst8255 (P1_U4742, P1_U3035, P1_U3060);
  nand ginst8256 (P1_U4743, P1_ADD_95_U4, P1_U3032);
  nand ginst8257 (P1_U4744, P1_R1222_U101, P1_U3031);
  nand ginst8258 (P1_U4745, P1_U3030, P1_U3461);
  nand ginst8259 (P1_U4746, P1_R1282_U20, P1_U3029);
  nand ginst8260 (P1_U4747, P1_U3035, P1_U3067);
  nand ginst8261 (P1_U4748, P1_ADD_95_U59, P1_U3032);
  nand ginst8262 (P1_U4749, P1_R1222_U100, P1_U3031);
  nand ginst8263 (P1_U4750, P1_U3030, P1_U3464);
  nand ginst8264 (P1_U4751, P1_R1282_U21, P1_U3029);
  nand ginst8265 (P1_U4752, P1_U3035, P1_U3071);
  nand ginst8266 (P1_U4753, P1_ADD_95_U58, P1_U3032);
  nand ginst8267 (P1_U4754, P1_R1222_U18, P1_U3031);
  nand ginst8268 (P1_U4755, P1_U3030, P1_U3467);
  nand ginst8269 (P1_U4756, P1_R1282_U65, P1_U3029);
  nand ginst8270 (P1_U4757, P1_U3035, P1_U3070);
  nand ginst8271 (P1_U4758, P1_ADD_95_U57, P1_U3032);
  nand ginst8272 (P1_U4759, P1_R1222_U99, P1_U3031);
  nand ginst8273 (P1_U4760, P1_U3030, P1_U3470);
  nand ginst8274 (P1_U4761, P1_R1282_U22, P1_U3029);
  nand ginst8275 (P1_U4762, P1_U3035, P1_U3084);
  nand ginst8276 (P1_U4763, P1_ADD_95_U56, P1_U3032);
  nand ginst8277 (P1_U4764, P1_R1222_U19, P1_U3031);
  nand ginst8278 (P1_U4765, P1_U3030, P1_U3473);
  nand ginst8279 (P1_U4766, P1_R1282_U23, P1_U3029);
  nand ginst8280 (P1_U4767, P1_U3035, P1_U3083);
  nand ginst8281 (P1_U4768, P1_ADD_95_U55, P1_U3032);
  nand ginst8282 (P1_U4769, P1_R1222_U98, P1_U3031);
  nand ginst8283 (P1_U4770, P1_U3030, P1_U3476);
  nand ginst8284 (P1_U4771, P1_R1282_U24, P1_U3029);
  nand ginst8285 (P1_U4772, P1_U3035, P1_U3062);
  nand ginst8286 (P1_U4773, P1_ADD_95_U54, P1_U3032);
  nand ginst8287 (P1_U4774, P1_R1222_U97, P1_U3031);
  nand ginst8288 (P1_U4775, P1_U3030, P1_U3479);
  nand ginst8289 (P1_U4776, P1_R1282_U63, P1_U3029);
  nand ginst8290 (P1_U4777, P1_U3035, P1_U3063);
  nand ginst8291 (P1_U4778, P1_ADD_95_U78, P1_U3032);
  nand ginst8292 (P1_U4779, P1_R1222_U11, P1_U3031);
  nand ginst8293 (P1_U4780, P1_U3030, P1_U3482);
  nand ginst8294 (P1_U4781, P1_R1282_U6, P1_U3029);
  nand ginst8295 (P1_U4782, P1_U3035, P1_U3072);
  nand ginst8296 (P1_U4783, P1_ADD_95_U77, P1_U3032);
  nand ginst8297 (P1_U4784, P1_R1222_U115, P1_U3031);
  nand ginst8298 (P1_U4785, P1_U3030, P1_U3485);
  nand ginst8299 (P1_U4786, P1_R1282_U7, P1_U3029);
  nand ginst8300 (P1_U4787, P1_U3035, P1_U3080);
  nand ginst8301 (P1_U4788, P1_ADD_95_U76, P1_U3032);
  nand ginst8302 (P1_U4789, P1_R1222_U114, P1_U3031);
  nand ginst8303 (P1_U4790, P1_U3030, P1_U3488);
  nand ginst8304 (P1_U4791, P1_R1282_U8, P1_U3029);
  nand ginst8305 (P1_U4792, P1_U3035, P1_U3079);
  nand ginst8306 (P1_U4793, P1_ADD_95_U75, P1_U3032);
  nand ginst8307 (P1_U4794, P1_R1222_U12, P1_U3031);
  nand ginst8308 (P1_U4795, P1_U3030, P1_U3491);
  nand ginst8309 (P1_U4796, P1_R1282_U86, P1_U3029);
  nand ginst8310 (P1_U4797, P1_U3035, P1_U3074);
  nand ginst8311 (P1_U4798, P1_ADD_95_U74, P1_U3032);
  nand ginst8312 (P1_U4799, P1_R1222_U113, P1_U3031);
  nand ginst8313 (P1_U4800, P1_U3030, P1_U3494);
  nand ginst8314 (P1_U4801, P1_R1282_U9, P1_U3029);
  nand ginst8315 (P1_U4802, P1_U3035, P1_U3073);
  nand ginst8316 (P1_U4803, P1_ADD_95_U73, P1_U3032);
  nand ginst8317 (P1_U4804, P1_R1222_U112, P1_U3031);
  nand ginst8318 (P1_U4805, P1_U3030, P1_U3497);
  nand ginst8319 (P1_U4806, P1_R1282_U10, P1_U3029);
  nand ginst8320 (P1_U4807, P1_U3035, P1_U3069);
  nand ginst8321 (P1_U4808, P1_ADD_95_U72, P1_U3032);
  nand ginst8322 (P1_U4809, P1_R1222_U111, P1_U3031);
  nand ginst8323 (P1_U4810, P1_U3030, P1_U3500);
  nand ginst8324 (P1_U4811, P1_R1282_U11, P1_U3029);
  nand ginst8325 (P1_U4812, P1_U3035, P1_U3082);
  nand ginst8326 (P1_U4813, P1_ADD_95_U71, P1_U3032);
  nand ginst8327 (P1_U4814, P1_R1222_U13, P1_U3031);
  nand ginst8328 (P1_U4815, P1_U3030, P1_U3503);
  nand ginst8329 (P1_U4816, P1_R1282_U84, P1_U3029);
  nand ginst8330 (P1_U4817, P1_U3035, P1_U3081);
  nand ginst8331 (P1_U4818, P1_ADD_95_U70, P1_U3032);
  nand ginst8332 (P1_U4819, P1_R1222_U110, P1_U3031);
  nand ginst8333 (P1_U4820, P1_U3030, P1_U3506);
  nand ginst8334 (P1_U4821, P1_R1282_U12, P1_U3029);
  nand ginst8335 (P1_U4822, P1_U3035, P1_U3076);
  nand ginst8336 (P1_U4823, P1_ADD_95_U69, P1_U3032);
  nand ginst8337 (P1_U4824, P1_R1222_U109, P1_U3031);
  nand ginst8338 (P1_U4825, P1_U3030, P1_U3508);
  nand ginst8339 (P1_U4826, P1_R1282_U82, P1_U3029);
  nand ginst8340 (P1_U4827, P1_U3035, P1_U3075);
  nand ginst8341 (P1_U4828, P1_ADD_95_U68, P1_U3032);
  nand ginst8342 (P1_U4829, P1_R1222_U14, P1_U3031);
  nand ginst8343 (P1_U4830, P1_U3030, P1_U3982);
  nand ginst8344 (P1_U4831, P1_R1282_U13, P1_U3029);
  nand ginst8345 (P1_U4832, P1_U3035, P1_U3061);
  nand ginst8346 (P1_U4833, P1_ADD_95_U67, P1_U3032);
  nand ginst8347 (P1_U4834, P1_R1222_U15, P1_U3031);
  nand ginst8348 (P1_U4835, P1_U3030, P1_U3981);
  nand ginst8349 (P1_U4836, P1_R1282_U78, P1_U3029);
  nand ginst8350 (P1_U4837, P1_U3035, P1_U3066);
  nand ginst8351 (P1_U4838, P1_ADD_95_U66, P1_U3032);
  nand ginst8352 (P1_U4839, P1_R1222_U108, P1_U3031);
  nand ginst8353 (P1_U4840, P1_U3030, P1_U3980);
  nand ginst8354 (P1_U4841, P1_R1282_U14, P1_U3029);
  nand ginst8355 (P1_U4842, P1_U3035, P1_U3065);
  nand ginst8356 (P1_U4843, P1_ADD_95_U65, P1_U3032);
  nand ginst8357 (P1_U4844, P1_R1222_U107, P1_U3031);
  nand ginst8358 (P1_U4845, P1_U3030, P1_U3979);
  nand ginst8359 (P1_U4846, P1_R1282_U76, P1_U3029);
  nand ginst8360 (P1_U4847, P1_U3035, P1_U3058);
  nand ginst8361 (P1_U4848, P1_ADD_95_U64, P1_U3032);
  nand ginst8362 (P1_U4849, P1_R1222_U106, P1_U3031);
  nand ginst8363 (P1_U4850, P1_U3030, P1_U3978);
  nand ginst8364 (P1_U4851, P1_R1282_U15, P1_U3029);
  nand ginst8365 (P1_U4852, P1_U3035, P1_U3057);
  nand ginst8366 (P1_U4853, P1_ADD_95_U63, P1_U3032);
  nand ginst8367 (P1_U4854, P1_R1222_U105, P1_U3031);
  nand ginst8368 (P1_U4855, P1_U3030, P1_U3977);
  nand ginst8369 (P1_U4856, P1_R1282_U74, P1_U3029);
  nand ginst8370 (P1_U4857, P1_U3035, P1_U3053);
  nand ginst8371 (P1_U4858, P1_ADD_95_U62, P1_U3032);
  nand ginst8372 (P1_U4859, P1_R1222_U16, P1_U3031);
  nand ginst8373 (P1_U4860, P1_U3030, P1_U3976);
  nand ginst8374 (P1_U4861, P1_R1282_U16, P1_U3029);
  nand ginst8375 (P1_U4862, P1_U3035, P1_U3054);
  nand ginst8376 (P1_U4863, P1_ADD_95_U61, P1_U3032);
  nand ginst8377 (P1_U4864, P1_R1222_U104, P1_U3031);
  nand ginst8378 (P1_U4865, P1_U3030, P1_U3975);
  nand ginst8379 (P1_U4866, P1_R1282_U72, P1_U3029);
  nand ginst8380 (P1_U4867, P1_U3035, P1_U3055);
  nand ginst8381 (P1_U4868, P1_ADD_95_U60, P1_U3032);
  nand ginst8382 (P1_U4869, P1_R1222_U103, P1_U3031);
  nand ginst8383 (P1_U4870, P1_U3030, P1_U3974);
  nand ginst8384 (P1_U4871, P1_R1282_U17, P1_U3029);
  nand ginst8385 (P1_U4872, P1_ADD_95_U5, P1_U3032);
  nand ginst8386 (P1_U4873, P1_R1222_U102, P1_U3031);
  nand ginst8387 (P1_U4874, P1_U3030, P1_U3985);
  nand ginst8388 (P1_U4875, P1_R1282_U70, P1_U3029);
  nand ginst8389 (P1_U4876, P1_U3030, P1_U3984);
  nand ginst8390 (P1_U4877, P1_R1282_U19, P1_U3029);
  nand ginst8391 (P1_U4878, P1_U3030, P1_U3983);
  nand ginst8392 (P1_U4879, P1_R1282_U68, P1_U3029);
  nand ginst8393 (P1_U4880, P1_U3418, P1_U3803, P1_U3804, P1_U3806, P1_U4726);
  nand ginst8394 (P1_U4881, P1_R1105_U13, P1_U3041);
  nand ginst8395 (P1_U4882, P1_U3039, P1_U3442);
  nand ginst8396 (P1_U4883, P1_R1162_U13, P1_U3037);
  nand ginst8397 (P1_U4884, P1_U4881, P1_U4882, P1_U4883);
  nand ginst8398 (P1_U4885, P1_U3046, P1_U3373);
  nand ginst8399 (P1_U4886, P1_U4885, P1_U5677);
  nand ginst8400 (P1_U4887, P1_U3912, P1_U4886);
  not ginst8401 (P1_U4888, P1_U3085);
  not ginst8402 (P1_U4889, P1_U3423);
  nand ginst8403 (P1_U4890, P1_U3043, P1_U4884);
  nand ginst8404 (P1_U4891, P1_R1105_U13, P1_U3042);
  nand ginst8405 (P1_U4892, P1_REG3_REG_19__SCAN_IN, P1_U3086);
  nand ginst8406 (P1_U4893, P1_U3040, P1_U3442);
  nand ginst8407 (P1_U4894, P1_R1162_U13, P1_U3038);
  nand ginst8408 (P1_U4895, P1_ADDR_REG_19__SCAN_IN, P1_U4889);
  nand ginst8409 (P1_U4896, P1_R1105_U75, P1_U3041);
  nand ginst8410 (P1_U4897, P1_U3039, P1_U3505);
  nand ginst8411 (P1_U4898, P1_R1162_U75, P1_U3037);
  nand ginst8412 (P1_U4899, P1_U4896, P1_U4897, P1_U4898);
  nand ginst8413 (P1_U4900, P1_U3043, P1_U4899);
  nand ginst8414 (P1_U4901, P1_R1105_U75, P1_U3042);
  nand ginst8415 (P1_U4902, P1_REG3_REG_18__SCAN_IN, P1_U3086);
  nand ginst8416 (P1_U4903, P1_U3040, P1_U3505);
  nand ginst8417 (P1_U4904, P1_R1162_U75, P1_U3038);
  nand ginst8418 (P1_U4905, P1_ADDR_REG_18__SCAN_IN, P1_U4889);
  nand ginst8419 (P1_U4906, P1_R1105_U12, P1_U3041);
  nand ginst8420 (P1_U4907, P1_U3039, P1_U3502);
  nand ginst8421 (P1_U4908, P1_R1162_U12, P1_U3037);
  nand ginst8422 (P1_U4909, P1_U4906, P1_U4907, P1_U4908);
  nand ginst8423 (P1_U4910, P1_U3043, P1_U4909);
  nand ginst8424 (P1_U4911, P1_R1105_U12, P1_U3042);
  nand ginst8425 (P1_U4912, P1_REG3_REG_17__SCAN_IN, P1_U3086);
  nand ginst8426 (P1_U4913, P1_U3040, P1_U3502);
  nand ginst8427 (P1_U4914, P1_R1162_U12, P1_U3038);
  nand ginst8428 (P1_U4915, P1_ADDR_REG_17__SCAN_IN, P1_U4889);
  nand ginst8429 (P1_U4916, P1_R1105_U76, P1_U3041);
  nand ginst8430 (P1_U4917, P1_U3039, P1_U3499);
  nand ginst8431 (P1_U4918, P1_R1162_U76, P1_U3037);
  nand ginst8432 (P1_U4919, P1_U4916, P1_U4917, P1_U4918);
  nand ginst8433 (P1_U4920, P1_U3043, P1_U4919);
  nand ginst8434 (P1_U4921, P1_R1105_U76, P1_U3042);
  nand ginst8435 (P1_U4922, P1_REG3_REG_16__SCAN_IN, P1_U3086);
  nand ginst8436 (P1_U4923, P1_U3040, P1_U3499);
  nand ginst8437 (P1_U4924, P1_R1162_U76, P1_U3038);
  nand ginst8438 (P1_U4925, P1_ADDR_REG_16__SCAN_IN, P1_U4889);
  nand ginst8439 (P1_U4926, P1_R1105_U77, P1_U3041);
  nand ginst8440 (P1_U4927, P1_U3039, P1_U3496);
  nand ginst8441 (P1_U4928, P1_R1162_U77, P1_U3037);
  nand ginst8442 (P1_U4929, P1_U4926, P1_U4927, P1_U4928);
  nand ginst8443 (P1_U4930, P1_U3043, P1_U4929);
  nand ginst8444 (P1_U4931, P1_R1105_U77, P1_U3042);
  nand ginst8445 (P1_U4932, P1_REG3_REG_15__SCAN_IN, P1_U3086);
  nand ginst8446 (P1_U4933, P1_U3040, P1_U3496);
  nand ginst8447 (P1_U4934, P1_R1162_U77, P1_U3038);
  nand ginst8448 (P1_U4935, P1_ADDR_REG_15__SCAN_IN, P1_U4889);
  nand ginst8449 (P1_U4936, P1_R1105_U78, P1_U3041);
  nand ginst8450 (P1_U4937, P1_U3039, P1_U3493);
  nand ginst8451 (P1_U4938, P1_R1162_U78, P1_U3037);
  nand ginst8452 (P1_U4939, P1_U4936, P1_U4937, P1_U4938);
  nand ginst8453 (P1_U4940, P1_U3043, P1_U4939);
  nand ginst8454 (P1_U4941, P1_R1105_U78, P1_U3042);
  nand ginst8455 (P1_U4942, P1_REG3_REG_14__SCAN_IN, P1_U3086);
  nand ginst8456 (P1_U4943, P1_U3040, P1_U3493);
  nand ginst8457 (P1_U4944, P1_R1162_U78, P1_U3038);
  nand ginst8458 (P1_U4945, P1_ADDR_REG_14__SCAN_IN, P1_U4889);
  nand ginst8459 (P1_U4946, P1_R1105_U11, P1_U3041);
  nand ginst8460 (P1_U4947, P1_U3039, P1_U3490);
  nand ginst8461 (P1_U4948, P1_R1162_U11, P1_U3037);
  nand ginst8462 (P1_U4949, P1_U4946, P1_U4947, P1_U4948);
  nand ginst8463 (P1_U4950, P1_U3043, P1_U4949);
  nand ginst8464 (P1_U4951, P1_R1105_U11, P1_U3042);
  nand ginst8465 (P1_U4952, P1_REG3_REG_13__SCAN_IN, P1_U3086);
  nand ginst8466 (P1_U4953, P1_U3040, P1_U3490);
  nand ginst8467 (P1_U4954, P1_R1162_U11, P1_U3038);
  nand ginst8468 (P1_U4955, P1_ADDR_REG_13__SCAN_IN, P1_U4889);
  nand ginst8469 (P1_U4956, P1_R1105_U79, P1_U3041);
  nand ginst8470 (P1_U4957, P1_U3039, P1_U3487);
  nand ginst8471 (P1_U4958, P1_R1162_U79, P1_U3037);
  nand ginst8472 (P1_U4959, P1_U4956, P1_U4957, P1_U4958);
  nand ginst8473 (P1_U4960, P1_U3043, P1_U4959);
  nand ginst8474 (P1_U4961, P1_R1105_U79, P1_U3042);
  nand ginst8475 (P1_U4962, P1_REG3_REG_12__SCAN_IN, P1_U3086);
  nand ginst8476 (P1_U4963, P1_U3040, P1_U3487);
  nand ginst8477 (P1_U4964, P1_R1162_U79, P1_U3038);
  nand ginst8478 (P1_U4965, P1_ADDR_REG_12__SCAN_IN, P1_U4889);
  nand ginst8479 (P1_U4966, P1_R1105_U80, P1_U3041);
  nand ginst8480 (P1_U4967, P1_U3039, P1_U3484);
  nand ginst8481 (P1_U4968, P1_R1162_U80, P1_U3037);
  nand ginst8482 (P1_U4969, P1_U4966, P1_U4967, P1_U4968);
  nand ginst8483 (P1_U4970, P1_U3043, P1_U4969);
  nand ginst8484 (P1_U4971, P1_R1105_U80, P1_U3042);
  nand ginst8485 (P1_U4972, P1_REG3_REG_11__SCAN_IN, P1_U3086);
  nand ginst8486 (P1_U4973, P1_U3040, P1_U3484);
  nand ginst8487 (P1_U4974, P1_R1162_U80, P1_U3038);
  nand ginst8488 (P1_U4975, P1_ADDR_REG_11__SCAN_IN, P1_U4889);
  nand ginst8489 (P1_U4976, P1_R1105_U10, P1_U3041);
  nand ginst8490 (P1_U4977, P1_U3039, P1_U3481);
  nand ginst8491 (P1_U4978, P1_R1162_U10, P1_U3037);
  nand ginst8492 (P1_U4979, P1_U4976, P1_U4977, P1_U4978);
  nand ginst8493 (P1_U4980, P1_U3043, P1_U4979);
  nand ginst8494 (P1_U4981, P1_R1105_U10, P1_U3042);
  nand ginst8495 (P1_U4982, P1_REG3_REG_10__SCAN_IN, P1_U3086);
  nand ginst8496 (P1_U4983, P1_U3040, P1_U3481);
  nand ginst8497 (P1_U4984, P1_R1162_U10, P1_U3038);
  nand ginst8498 (P1_U4985, P1_ADDR_REG_10__SCAN_IN, P1_U4889);
  nand ginst8499 (P1_U4986, P1_R1105_U70, P1_U3041);
  nand ginst8500 (P1_U4987, P1_U3039, P1_U3478);
  nand ginst8501 (P1_U4988, P1_R1162_U70, P1_U3037);
  nand ginst8502 (P1_U4989, P1_U4986, P1_U4987, P1_U4988);
  nand ginst8503 (P1_U4990, P1_U3043, P1_U4989);
  nand ginst8504 (P1_U4991, P1_R1105_U70, P1_U3042);
  nand ginst8505 (P1_U4992, P1_REG3_REG_9__SCAN_IN, P1_U3086);
  nand ginst8506 (P1_U4993, P1_U3040, P1_U3478);
  nand ginst8507 (P1_U4994, P1_R1162_U70, P1_U3038);
  nand ginst8508 (P1_U4995, P1_ADDR_REG_9__SCAN_IN, P1_U4889);
  nand ginst8509 (P1_U4996, P1_R1105_U71, P1_U3041);
  nand ginst8510 (P1_U4997, P1_U3039, P1_U3475);
  nand ginst8511 (P1_U4998, P1_R1162_U71, P1_U3037);
  nand ginst8512 (P1_U4999, P1_U4996, P1_U4997, P1_U4998);
  nand ginst8513 (P1_U5000, P1_U3043, P1_U4999);
  nand ginst8514 (P1_U5001, P1_R1105_U71, P1_U3042);
  nand ginst8515 (P1_U5002, P1_REG3_REG_8__SCAN_IN, P1_U3086);
  nand ginst8516 (P1_U5003, P1_U3040, P1_U3475);
  nand ginst8517 (P1_U5004, P1_R1162_U71, P1_U3038);
  nand ginst8518 (P1_U5005, P1_ADDR_REG_8__SCAN_IN, P1_U4889);
  nand ginst8519 (P1_U5006, P1_R1105_U16, P1_U3041);
  nand ginst8520 (P1_U5007, P1_U3039, P1_U3472);
  nand ginst8521 (P1_U5008, P1_R1162_U16, P1_U3037);
  nand ginst8522 (P1_U5009, P1_U5006, P1_U5007, P1_U5008);
  nand ginst8523 (P1_U5010, P1_U3043, P1_U5009);
  nand ginst8524 (P1_U5011, P1_R1105_U16, P1_U3042);
  nand ginst8525 (P1_U5012, P1_REG3_REG_7__SCAN_IN, P1_U3086);
  nand ginst8526 (P1_U5013, P1_U3040, P1_U3472);
  nand ginst8527 (P1_U5014, P1_R1162_U16, P1_U3038);
  nand ginst8528 (P1_U5015, P1_ADDR_REG_7__SCAN_IN, P1_U4889);
  nand ginst8529 (P1_U5016, P1_R1105_U72, P1_U3041);
  nand ginst8530 (P1_U5017, P1_U3039, P1_U3469);
  nand ginst8531 (P1_U5018, P1_R1162_U72, P1_U3037);
  nand ginst8532 (P1_U5019, P1_U5016, P1_U5017, P1_U5018);
  nand ginst8533 (P1_U5020, P1_U3043, P1_U5019);
  nand ginst8534 (P1_U5021, P1_R1105_U72, P1_U3042);
  nand ginst8535 (P1_U5022, P1_REG3_REG_6__SCAN_IN, P1_U3086);
  nand ginst8536 (P1_U5023, P1_U3040, P1_U3469);
  nand ginst8537 (P1_U5024, P1_R1162_U72, P1_U3038);
  nand ginst8538 (P1_U5025, P1_ADDR_REG_6__SCAN_IN, P1_U4889);
  nand ginst8539 (P1_U5026, P1_R1105_U15, P1_U3041);
  nand ginst8540 (P1_U5027, P1_U3039, P1_U3466);
  nand ginst8541 (P1_U5028, P1_R1162_U15, P1_U3037);
  nand ginst8542 (P1_U5029, P1_U5026, P1_U5027, P1_U5028);
  nand ginst8543 (P1_U5030, P1_U3043, P1_U5029);
  nand ginst8544 (P1_U5031, P1_R1105_U15, P1_U3042);
  nand ginst8545 (P1_U5032, P1_REG3_REG_5__SCAN_IN, P1_U3086);
  nand ginst8546 (P1_U5033, P1_U3040, P1_U3466);
  nand ginst8547 (P1_U5034, P1_R1162_U15, P1_U3038);
  nand ginst8548 (P1_U5035, P1_ADDR_REG_5__SCAN_IN, P1_U4889);
  nand ginst8549 (P1_U5036, P1_R1105_U73, P1_U3041);
  nand ginst8550 (P1_U5037, P1_U3039, P1_U3463);
  nand ginst8551 (P1_U5038, P1_R1162_U73, P1_U3037);
  nand ginst8552 (P1_U5039, P1_U5036, P1_U5037, P1_U5038);
  nand ginst8553 (P1_U5040, P1_U3043, P1_U5039);
  nand ginst8554 (P1_U5041, P1_R1105_U73, P1_U3042);
  nand ginst8555 (P1_U5042, P1_REG3_REG_4__SCAN_IN, P1_U3086);
  nand ginst8556 (P1_U5043, P1_U3040, P1_U3463);
  nand ginst8557 (P1_U5044, P1_R1162_U73, P1_U3038);
  nand ginst8558 (P1_U5045, P1_ADDR_REG_4__SCAN_IN, P1_U4889);
  nand ginst8559 (P1_U5046, P1_R1105_U74, P1_U3041);
  nand ginst8560 (P1_U5047, P1_U3039, P1_U3460);
  nand ginst8561 (P1_U5048, P1_R1162_U74, P1_U3037);
  nand ginst8562 (P1_U5049, P1_U5046, P1_U5047, P1_U5048);
  nand ginst8563 (P1_U5050, P1_U3043, P1_U5049);
  nand ginst8564 (P1_U5051, P1_R1105_U74, P1_U3042);
  nand ginst8565 (P1_U5052, P1_REG3_REG_3__SCAN_IN, P1_U3086);
  nand ginst8566 (P1_U5053, P1_U3040, P1_U3460);
  nand ginst8567 (P1_U5054, P1_R1162_U74, P1_U3038);
  nand ginst8568 (P1_U5055, P1_ADDR_REG_3__SCAN_IN, P1_U4889);
  nand ginst8569 (P1_U5056, P1_R1105_U14, P1_U3041);
  nand ginst8570 (P1_U5057, P1_U3039, P1_U3457);
  nand ginst8571 (P1_U5058, P1_R1162_U14, P1_U3037);
  nand ginst8572 (P1_U5059, P1_U5056, P1_U5057, P1_U5058);
  nand ginst8573 (P1_U5060, P1_U3043, P1_U5059);
  nand ginst8574 (P1_U5061, P1_R1105_U14, P1_U3042);
  nand ginst8575 (P1_U5062, P1_REG3_REG_2__SCAN_IN, P1_U3086);
  nand ginst8576 (P1_U5063, P1_U3040, P1_U3457);
  nand ginst8577 (P1_U5064, P1_R1162_U14, P1_U3038);
  nand ginst8578 (P1_U5065, P1_ADDR_REG_2__SCAN_IN, P1_U4889);
  nand ginst8579 (P1_U5066, P1_R1105_U68, P1_U3041);
  nand ginst8580 (P1_U5067, P1_U3039, P1_U3454);
  nand ginst8581 (P1_U5068, P1_R1162_U68, P1_U3037);
  nand ginst8582 (P1_U5069, P1_U5066, P1_U5067, P1_U5068);
  nand ginst8583 (P1_U5070, P1_U3043, P1_U5069);
  nand ginst8584 (P1_U5071, P1_R1105_U68, P1_U3042);
  nand ginst8585 (P1_U5072, P1_REG3_REG_1__SCAN_IN, P1_U3086);
  nand ginst8586 (P1_U5073, P1_U3040, P1_U3454);
  nand ginst8587 (P1_U5074, P1_R1162_U68, P1_U3038);
  nand ginst8588 (P1_U5075, P1_ADDR_REG_1__SCAN_IN, P1_U4889);
  nand ginst8589 (P1_U5076, P1_R1105_U69, P1_U3041);
  nand ginst8590 (P1_U5077, P1_U3039, P1_U3448);
  nand ginst8591 (P1_U5078, P1_R1162_U69, P1_U3037);
  nand ginst8592 (P1_U5079, P1_U5076, P1_U5077, P1_U5078);
  nand ginst8593 (P1_U5080, P1_U3043, P1_U5079);
  nand ginst8594 (P1_U5081, P1_R1105_U69, P1_U3042);
  nand ginst8595 (P1_U5082, P1_REG3_REG_0__SCAN_IN, P1_U3086);
  nand ginst8596 (P1_U5083, P1_U3040, P1_U3448);
  nand ginst8597 (P1_U5084, P1_R1162_U69, P1_U3038);
  nand ginst8598 (P1_U5085, P1_ADDR_REG_0__SCAN_IN, P1_U4889);
  not ginst8599 (P1_U5086, P1_U3951);
  nand ginst8600 (P1_U5087, P1_LT_197_U13, P1_U3954, P1_U3987);
  nand ginst8601 (P1_U5088, P1_U3427, P1_U5677);
  nand ginst8602 (P1_U5089, P1_U3851, P1_U5088);
  nand ginst8603 (P1_U5090, P1_U3022, P1_U3949, P1_U3986);
  nand ginst8604 (P1_U5091, P1_B_REG_SCAN_IN, P1_U5089);
  nand ginst8605 (P1_U5092, P1_U3036, P1_U3079);
  nand ginst8606 (P1_U5093, P1_U3034, P1_U3073);
  nand ginst8607 (P1_U5094, P1_ADD_95_U73, P1_U3430);
  nand ginst8608 (P1_U5095, P1_U5092, P1_U5093, P1_U5094);
  nand ginst8609 (P1_U5096, P1_U3361, P1_U3362, P1_U3364);
  nand ginst8610 (P1_U5097, P1_U3365, P1_U3366, P1_U3419);
  nand ginst8611 (P1_U5098, P1_U5097, P1_U5684);
  nand ginst8612 (P1_U5099, P1_U5096, P1_U5693);
  nand ginst8613 (P1_U5100, P1_U3868, P1_U5098, P1_U5099);
  nand ginst8614 (P1_U5101, P1_U3430, P1_U5100);
  not ginst8615 (P1_U5102, P1_U3432);
  nand ginst8616 (P1_U5103, P1_U3497, P1_U5656);
  nand ginst8617 (P1_U5104, P1_ADD_95_U73, P1_U5655);
  nand ginst8618 (P1_U5105, P1_U3994, P1_U5095);
  nand ginst8619 (P1_U5106, P1_R1165_U104, P1_U3027);
  nand ginst8620 (P1_U5107, P1_REG3_REG_15__SCAN_IN, P1_U3086);
  nand ginst8621 (P1_U5108, P1_U3036, P1_U3058);
  nand ginst8622 (P1_U5109, P1_U3034, P1_U3053);
  nand ginst8623 (P1_U5110, P1_ADD_95_U62, P1_U3430);
  nand ginst8624 (P1_U5111, P1_U5108, P1_U5109, P1_U5110);
  nand ginst8625 (P1_U5112, P1_U3422, P1_U3430);
  nand ginst8626 (P1_U5113, P1_U5102, P1_U5112);
  nand ginst8627 (P1_U5114, P1_U3422, P1_U3972);
  nand ginst8628 (P1_U5115, P1_U3418, P1_U5114);
  nand ginst8629 (P1_U5116, P1_U3045, P1_U3976);
  nand ginst8630 (P1_U5117, P1_ADD_95_U62, P1_U3044);
  nand ginst8631 (P1_U5118, P1_U3994, P1_U5111);
  nand ginst8632 (P1_U5119, P1_R1165_U13, P1_U3027);
  nand ginst8633 (P1_U5120, P1_REG3_REG_26__SCAN_IN, P1_U3086);
  nand ginst8634 (P1_U5121, P1_U3036, P1_U3067);
  nand ginst8635 (P1_U5122, P1_U3034, P1_U3070);
  nand ginst8636 (P1_U5123, P1_ADD_95_U57, P1_U3430);
  nand ginst8637 (P1_U5124, P1_U5121, P1_U5122, P1_U5123);
  nand ginst8638 (P1_U5125, P1_U3470, P1_U5656);
  nand ginst8639 (P1_U5126, P1_ADD_95_U57, P1_U5655);
  nand ginst8640 (P1_U5127, P1_U3994, P1_U5124);
  nand ginst8641 (P1_U5128, P1_R1165_U89, P1_U3027);
  nand ginst8642 (P1_U5129, P1_REG3_REG_6__SCAN_IN, P1_U3086);
  nand ginst8643 (P1_U5130, P1_U3036, P1_U3069);
  nand ginst8644 (P1_U5131, P1_U3034, P1_U3081);
  nand ginst8645 (P1_U5132, P1_ADD_95_U70, P1_U3430);
  nand ginst8646 (P1_U5133, P1_U5130, P1_U5131, P1_U5132);
  nand ginst8647 (P1_U5134, P1_U3506, P1_U5656);
  nand ginst8648 (P1_U5135, P1_ADD_95_U70, P1_U5655);
  nand ginst8649 (P1_U5136, P1_U3994, P1_U5133);
  nand ginst8650 (P1_U5137, P1_R1165_U102, P1_U3027);
  nand ginst8651 (P1_U5138, P1_REG3_REG_18__SCAN_IN, P1_U3086);
  nand ginst8652 (P1_U5139, P1_U3036, P1_U3078);
  nand ginst8653 (P1_U5140, P1_U3034, P1_U3064);
  nand ginst8654 (P1_U5141, P1_REG3_REG_2__SCAN_IN, P1_U3430);
  nand ginst8655 (P1_U5142, P1_U5139, P1_U5140, P1_U5141);
  nand ginst8656 (P1_U5143, P1_U3458, P1_U5656);
  nand ginst8657 (P1_U5144, P1_REG3_REG_2__SCAN_IN, P1_U5655);
  nand ginst8658 (P1_U5145, P1_U3994, P1_U5142);
  nand ginst8659 (P1_U5146, P1_R1165_U92, P1_U3027);
  nand ginst8660 (P1_U5147, P1_REG3_REG_2__SCAN_IN, P1_U3086);
  nand ginst8661 (P1_U5148, P1_U3036, P1_U3062);
  nand ginst8662 (P1_U5149, P1_U3034, P1_U3072);
  nand ginst8663 (P1_U5150, P1_ADD_95_U77, P1_U3430);
  nand ginst8664 (P1_U5151, P1_U5148, P1_U5149, P1_U5150);
  nand ginst8665 (P1_U5152, P1_U3485, P1_U5656);
  nand ginst8666 (P1_U5153, P1_ADD_95_U77, P1_U5655);
  nand ginst8667 (P1_U5154, P1_U3994, P1_U5151);
  nand ginst8668 (P1_U5155, P1_R1165_U107, P1_U3027);
  nand ginst8669 (P1_U5156, P1_REG3_REG_11__SCAN_IN, P1_U3086);
  nand ginst8670 (P1_U5157, P1_U3036, P1_U3075);
  nand ginst8671 (P1_U5158, P1_U3034, P1_U3066);
  nand ginst8672 (P1_U5159, P1_ADD_95_U66, P1_U3430);
  nand ginst8673 (P1_U5160, P1_U5157, P1_U5158, P1_U5159);
  nand ginst8674 (P1_U5161, P1_U3045, P1_U3980);
  nand ginst8675 (P1_U5162, P1_ADD_95_U66, P1_U3044);
  nand ginst8676 (P1_U5163, P1_U3994, P1_U5160);
  nand ginst8677 (P1_U5164, P1_R1165_U98, P1_U3027);
  nand ginst8678 (P1_U5165, P1_REG3_REG_22__SCAN_IN, P1_U3086);
  nand ginst8679 (P1_U5166, P1_U3036, P1_U3072);
  nand ginst8680 (P1_U5167, P1_U3034, P1_U3079);
  nand ginst8681 (P1_U5168, P1_ADD_95_U75, P1_U3430);
  nand ginst8682 (P1_U5169, P1_U5166, P1_U5167, P1_U5168);
  nand ginst8683 (P1_U5170, P1_U3491, P1_U5656);
  nand ginst8684 (P1_U5171, P1_ADD_95_U75, P1_U5655);
  nand ginst8685 (P1_U5172, P1_U3994, P1_U5169);
  nand ginst8686 (P1_U5173, P1_R1165_U10, P1_U3027);
  nand ginst8687 (P1_U5174, P1_REG3_REG_13__SCAN_IN, P1_U3086);
  nand ginst8688 (P1_U5175, P1_U3036, P1_U3081);
  nand ginst8689 (P1_U5176, P1_U3034, P1_U3075);
  nand ginst8690 (P1_U5177, P1_ADD_95_U68, P1_U3430);
  nand ginst8691 (P1_U5178, P1_U5175, P1_U5176, P1_U5177);
  nand ginst8692 (P1_U5179, P1_U3045, P1_U3982);
  nand ginst8693 (P1_U5180, P1_ADD_95_U68, P1_U3044);
  nand ginst8694 (P1_U5181, P1_U3994, P1_U5178);
  nand ginst8695 (P1_U5182, P1_R1165_U99, P1_U3027);
  nand ginst8696 (P1_U5183, P1_REG3_REG_20__SCAN_IN, P1_U3086);
  nand ginst8697 (P1_U5184, P1_U3429, P1_U3431);
  nand ginst8698 (P1_U5185, P1_U3430, P1_U5184);
  nand ginst8699 (P1_U5186, P1_U3995, P1_U5185);
  nand ginst8700 (P1_U5187, P1_U3034, P1_U3873);
  nand ginst8701 (P1_U5188, P1_U3450, P1_U5656);
  nand ginst8702 (P1_U5189, P1_REG3_REG_0__SCAN_IN, P1_U5186);
  nand ginst8703 (P1_U5190, P1_R1165_U86, P1_U3027);
  nand ginst8704 (P1_U5191, P1_REG3_REG_0__SCAN_IN, P1_U3086);
  nand ginst8705 (P1_U5192, P1_U3036, P1_U3084);
  nand ginst8706 (P1_U5193, P1_U3034, P1_U3062);
  nand ginst8707 (P1_U5194, P1_ADD_95_U54, P1_U3430);
  nand ginst8708 (P1_U5195, P1_U5192, P1_U5193, P1_U5194);
  nand ginst8709 (P1_U5196, P1_U3479, P1_U5656);
  nand ginst8710 (P1_U5197, P1_ADD_95_U54, P1_U5655);
  nand ginst8711 (P1_U5198, P1_U3994, P1_U5195);
  nand ginst8712 (P1_U5199, P1_R1165_U87, P1_U3027);
  nand ginst8713 (P1_U5200, P1_REG3_REG_9__SCAN_IN, P1_U3086);
  nand ginst8714 (P1_U5201, P1_U3036, P1_U3064);
  nand ginst8715 (P1_U5202, P1_U3034, P1_U3067);
  nand ginst8716 (P1_U5203, P1_ADD_95_U59, P1_U3430);
  nand ginst8717 (P1_U5204, P1_U5201, P1_U5202, P1_U5203);
  nand ginst8718 (P1_U5205, P1_U3464, P1_U5656);
  nand ginst8719 (P1_U5206, P1_ADD_95_U59, P1_U5655);
  nand ginst8720 (P1_U5207, P1_U3994, P1_U5204);
  nand ginst8721 (P1_U5208, P1_R1165_U91, P1_U3027);
  nand ginst8722 (P1_U5209, P1_REG3_REG_4__SCAN_IN, P1_U3086);
  nand ginst8723 (P1_U5210, P1_U3036, P1_U3066);
  nand ginst8724 (P1_U5211, P1_U3034, P1_U3058);
  nand ginst8725 (P1_U5212, P1_ADD_95_U64, P1_U3430);
  nand ginst8726 (P1_U5213, P1_U5210, P1_U5211, P1_U5212);
  nand ginst8727 (P1_U5214, P1_U3045, P1_U3978);
  nand ginst8728 (P1_U5215, P1_ADD_95_U64, P1_U3044);
  nand ginst8729 (P1_U5216, P1_U3994, P1_U5213);
  nand ginst8730 (P1_U5217, P1_R1165_U96, P1_U3027);
  nand ginst8731 (P1_U5218, P1_REG3_REG_24__SCAN_IN, P1_U3086);
  nand ginst8732 (P1_U5219, P1_U3036, P1_U3073);
  nand ginst8733 (P1_U5220, P1_U3034, P1_U3082);
  nand ginst8734 (P1_U5221, P1_ADD_95_U71, P1_U3430);
  nand ginst8735 (P1_U5222, P1_U5219, P1_U5220, P1_U5221);
  nand ginst8736 (P1_U5223, P1_U3503, P1_U5656);
  nand ginst8737 (P1_U5224, P1_ADD_95_U71, P1_U5655);
  nand ginst8738 (P1_U5225, P1_U3994, P1_U5222);
  nand ginst8739 (P1_U5226, P1_R1165_U11, P1_U3027);
  nand ginst8740 (P1_U5227, P1_REG3_REG_17__SCAN_IN, P1_U3086);
  nand ginst8741 (P1_U5228, P1_U3036, P1_U3060);
  nand ginst8742 (P1_U5229, P1_U3034, P1_U3071);
  nand ginst8743 (P1_U5230, P1_ADD_95_U58, P1_U3430);
  nand ginst8744 (P1_U5231, P1_U5228, P1_U5229, P1_U5230);
  nand ginst8745 (P1_U5232, P1_U3467, P1_U5656);
  nand ginst8746 (P1_U5233, P1_ADD_95_U58, P1_U5655);
  nand ginst8747 (P1_U5234, P1_U3994, P1_U5231);
  nand ginst8748 (P1_U5235, P1_R1165_U90, P1_U3027);
  nand ginst8749 (P1_U5236, P1_REG3_REG_5__SCAN_IN, P1_U3086);
  nand ginst8750 (P1_U5237, P1_U3036, P1_U3074);
  nand ginst8751 (P1_U5238, P1_U3034, P1_U3069);
  nand ginst8752 (P1_U5239, P1_ADD_95_U72, P1_U3430);
  nand ginst8753 (P1_U5240, P1_U5237, P1_U5238, P1_U5239);
  nand ginst8754 (P1_U5241, P1_U3500, P1_U5656);
  nand ginst8755 (P1_U5242, P1_ADD_95_U72, P1_U5655);
  nand ginst8756 (P1_U5243, P1_U3994, P1_U5240);
  nand ginst8757 (P1_U5244, P1_R1165_U103, P1_U3027);
  nand ginst8758 (P1_U5245, P1_REG3_REG_16__SCAN_IN, P1_U3086);
  nand ginst8759 (P1_U5246, P1_U3036, P1_U3065);
  nand ginst8760 (P1_U5247, P1_U3034, P1_U3057);
  nand ginst8761 (P1_U5248, P1_ADD_95_U63, P1_U3430);
  nand ginst8762 (P1_U5249, P1_U5246, P1_U5247, P1_U5248);
  nand ginst8763 (P1_U5250, P1_U3045, P1_U3977);
  nand ginst8764 (P1_U5251, P1_ADD_95_U63, P1_U3044);
  nand ginst8765 (P1_U5252, P1_U3994, P1_U5249);
  nand ginst8766 (P1_U5253, P1_R1165_U95, P1_U3027);
  nand ginst8767 (P1_U5254, P1_REG3_REG_25__SCAN_IN, P1_U3086);
  nand ginst8768 (P1_U5255, P1_U3036, P1_U3063);
  nand ginst8769 (P1_U5256, P1_U3034, P1_U3080);
  nand ginst8770 (P1_U5257, P1_ADD_95_U76, P1_U3430);
  nand ginst8771 (P1_U5258, P1_U5255, P1_U5256, P1_U5257);
  nand ginst8772 (P1_U5259, P1_U3488, P1_U5656);
  nand ginst8773 (P1_U5260, P1_ADD_95_U76, P1_U5655);
  nand ginst8774 (P1_U5261, P1_U3994, P1_U5258);
  nand ginst8775 (P1_U5262, P1_R1165_U106, P1_U3027);
  nand ginst8776 (P1_U5263, P1_REG3_REG_12__SCAN_IN, P1_U3086);
  nand ginst8777 (P1_U5264, P1_U3036, P1_U3076);
  nand ginst8778 (P1_U5265, P1_U3034, P1_U3061);
  nand ginst8779 (P1_U5266, P1_ADD_95_U67, P1_U3430);
  nand ginst8780 (P1_U5267, P1_U5264, P1_U5265, P1_U5266);
  nand ginst8781 (P1_U5268, P1_U3045, P1_U3981);
  nand ginst8782 (P1_U5269, P1_ADD_95_U67, P1_U3044);
  nand ginst8783 (P1_U5270, P1_U3994, P1_U5267);
  nand ginst8784 (P1_U5271, P1_R1165_U12, P1_U3027);
  nand ginst8785 (P1_U5272, P1_REG3_REG_21__SCAN_IN, P1_U3086);
  nand ginst8786 (P1_U5273, P1_U3036, P1_U3077);
  nand ginst8787 (P1_U5274, P1_U3034, P1_U3068);
  nand ginst8788 (P1_U5275, P1_REG3_REG_1__SCAN_IN, P1_U3430);
  nand ginst8789 (P1_U5276, P1_U5273, P1_U5274, P1_U5275);
  nand ginst8790 (P1_U5277, P1_U3455, P1_U5656);
  nand ginst8791 (P1_U5278, P1_REG3_REG_1__SCAN_IN, P1_U5655);
  nand ginst8792 (P1_U5279, P1_U3994, P1_U5276);
  nand ginst8793 (P1_U5280, P1_R1165_U100, P1_U3027);
  nand ginst8794 (P1_U5281, P1_REG3_REG_1__SCAN_IN, P1_U3086);
  nand ginst8795 (P1_U5282, P1_U3036, P1_U3070);
  nand ginst8796 (P1_U5283, P1_U3034, P1_U3083);
  nand ginst8797 (P1_U5284, P1_ADD_95_U55, P1_U3430);
  nand ginst8798 (P1_U5285, P1_U5282, P1_U5283, P1_U5284);
  nand ginst8799 (P1_U5286, P1_U3476, P1_U5656);
  nand ginst8800 (P1_U5287, P1_ADD_95_U55, P1_U5655);
  nand ginst8801 (P1_U5288, P1_U3994, P1_U5285);
  nand ginst8802 (P1_U5289, P1_R1165_U88, P1_U3027);
  nand ginst8803 (P1_U5290, P1_REG3_REG_8__SCAN_IN, P1_U3086);
  nand ginst8804 (P1_U5291, P1_U3036, P1_U3053);
  nand ginst8805 (P1_U5292, P1_U3034, P1_U3055);
  nand ginst8806 (P1_U5293, P1_ADD_95_U60, P1_U3430);
  nand ginst8807 (P1_U5294, P1_U5291, P1_U5292, P1_U5293);
  nand ginst8808 (P1_U5295, P1_U3045, P1_U3974);
  nand ginst8809 (P1_U5296, P1_ADD_95_U60, P1_U3044);
  nand ginst8810 (P1_U5297, P1_U3994, P1_U5294);
  nand ginst8811 (P1_U5298, P1_R1165_U93, P1_U3027);
  nand ginst8812 (P1_U5299, P1_REG3_REG_28__SCAN_IN, P1_U3086);
  nand ginst8813 (P1_U5300, P1_U3036, P1_U3082);
  nand ginst8814 (P1_U5301, P1_U3034, P1_U3076);
  nand ginst8815 (P1_U5302, P1_ADD_95_U69, P1_U3430);
  nand ginst8816 (P1_U5303, P1_U5300, P1_U5301, P1_U5302);
  nand ginst8817 (P1_U5304, P1_U3508, P1_U5656);
  nand ginst8818 (P1_U5305, P1_ADD_95_U69, P1_U5655);
  nand ginst8819 (P1_U5306, P1_U3994, P1_U5303);
  nand ginst8820 (P1_U5307, P1_R1165_U101, P1_U3027);
  nand ginst8821 (P1_U5308, P1_REG3_REG_19__SCAN_IN, P1_U3086);
  nand ginst8822 (P1_U5309, P1_U3036, P1_U3068);
  nand ginst8823 (P1_U5310, P1_U3034, P1_U3060);
  nand ginst8824 (P1_U5311, P1_ADD_95_U4, P1_U3430);
  nand ginst8825 (P1_U5312, P1_U5309, P1_U5310, P1_U5311);
  nand ginst8826 (P1_U5313, P1_U3461, P1_U5656);
  nand ginst8827 (P1_U5314, P1_ADD_95_U4, P1_U5655);
  nand ginst8828 (P1_U5315, P1_U3994, P1_U5312);
  nand ginst8829 (P1_U5316, P1_R1165_U14, P1_U3027);
  nand ginst8830 (P1_U5317, P1_REG3_REG_3__SCAN_IN, P1_U3086);
  nand ginst8831 (P1_U5318, P1_U3036, P1_U3083);
  nand ginst8832 (P1_U5319, P1_U3034, P1_U3063);
  nand ginst8833 (P1_U5320, P1_ADD_95_U78, P1_U3430);
  nand ginst8834 (P1_U5321, P1_U5318, P1_U5319, P1_U5320);
  nand ginst8835 (P1_U5322, P1_U3482, P1_U5656);
  nand ginst8836 (P1_U5323, P1_ADD_95_U78, P1_U5655);
  nand ginst8837 (P1_U5324, P1_U3994, P1_U5321);
  nand ginst8838 (P1_U5325, P1_R1165_U108, P1_U3027);
  nand ginst8839 (P1_U5326, P1_REG3_REG_10__SCAN_IN, P1_U3086);
  nand ginst8840 (P1_U5327, P1_U3036, P1_U3061);
  nand ginst8841 (P1_U5328, P1_U3034, P1_U3065);
  nand ginst8842 (P1_U5329, P1_ADD_95_U65, P1_U3430);
  nand ginst8843 (P1_U5330, P1_U5327, P1_U5328, P1_U5329);
  nand ginst8844 (P1_U5331, P1_U3045, P1_U3979);
  nand ginst8845 (P1_U5332, P1_ADD_95_U65, P1_U3044);
  nand ginst8846 (P1_U5333, P1_U3994, P1_U5330);
  nand ginst8847 (P1_U5334, P1_R1165_U97, P1_U3027);
  nand ginst8848 (P1_U5335, P1_REG3_REG_23__SCAN_IN, P1_U3086);
  nand ginst8849 (P1_U5336, P1_U3036, P1_U3080);
  nand ginst8850 (P1_U5337, P1_U3034, P1_U3074);
  nand ginst8851 (P1_U5338, P1_ADD_95_U74, P1_U3430);
  nand ginst8852 (P1_U5339, P1_U5336, P1_U5337, P1_U5338);
  nand ginst8853 (P1_U5340, P1_U3494, P1_U5656);
  nand ginst8854 (P1_U5341, P1_ADD_95_U74, P1_U5655);
  nand ginst8855 (P1_U5342, P1_U3994, P1_U5339);
  nand ginst8856 (P1_U5343, P1_R1165_U105, P1_U3027);
  nand ginst8857 (P1_U5344, P1_REG3_REG_14__SCAN_IN, P1_U3086);
  nand ginst8858 (P1_U5345, P1_U3036, P1_U3057);
  nand ginst8859 (P1_U5346, P1_U3034, P1_U3054);
  nand ginst8860 (P1_U5347, P1_ADD_95_U61, P1_U3430);
  nand ginst8861 (P1_U5348, P1_U5345, P1_U5346, P1_U5347);
  nand ginst8862 (P1_U5349, P1_U3045, P1_U3975);
  nand ginst8863 (P1_U5350, P1_ADD_95_U61, P1_U3044);
  nand ginst8864 (P1_U5351, P1_U3994, P1_U5348);
  nand ginst8865 (P1_U5352, P1_R1165_U94, P1_U3027);
  nand ginst8866 (P1_U5353, P1_REG3_REG_27__SCAN_IN, P1_U3086);
  nand ginst8867 (P1_U5354, P1_U3036, P1_U3071);
  nand ginst8868 (P1_U5355, P1_U3034, P1_U3084);
  nand ginst8869 (P1_U5356, P1_ADD_95_U56, P1_U3430);
  nand ginst8870 (P1_U5357, P1_U5354, P1_U5355, P1_U5356);
  nand ginst8871 (P1_U5358, P1_U3473, P1_U5656);
  nand ginst8872 (P1_U5359, P1_ADD_95_U56, P1_U5655);
  nand ginst8873 (P1_U5360, P1_U3994, P1_U5357);
  nand ginst8874 (P1_U5361, P1_R1165_U15, P1_U3027);
  nand ginst8875 (P1_U5362, P1_REG3_REG_7__SCAN_IN, P1_U3086);
  nand ginst8876 (P1_U5363, P1_U3375, P1_U3449);
  nand ginst8877 (P1_U5364, P1_U3446, P1_U5363);
  nand ginst8878 (P1_U5365, P1_R1165_U86, P1_U3446, P1_U5702);
  nand ginst8879 (P1_U5366, P1_U3441, P1_U3447);
  nand ginst8880 (P1_U5367, P1_U3877, P1_U3970);
  nand ginst8881 (P1_U5368, P1_U3370, P1_U3419);
  nand ginst8882 (P1_U5369, P1_U3363, P1_U3365, P1_U3368);
  nand ginst8883 (P1_U5370, P1_U3421, P1_U4000);
  nand ginst8884 (P1_U5371, P1_U3421, P1_U5369);
  not ginst8885 (P1_U5372, P1_U3434);
  nand ginst8886 (P1_U5373, P1_U3970, P1_U5372);
  nand ginst8887 (P1_U5374, P1_U3479, P1_U5373);
  nand ginst8888 (P1_U5375, P1_U3021, P1_U3083);
  nand ginst8889 (P1_U5376, P1_U3476, P1_U5373);
  nand ginst8890 (P1_U5377, P1_U3021, P1_U3084);
  nand ginst8891 (P1_U5378, P1_U3473, P1_U5373);
  nand ginst8892 (P1_U5379, P1_U3021, P1_U3070);
  nand ginst8893 (P1_U5380, P1_U3470, P1_U5373);
  nand ginst8894 (P1_U5381, P1_U3021, P1_U3071);
  nand ginst8895 (P1_U5382, P1_U3467, P1_U5373);
  nand ginst8896 (P1_U5383, P1_U3021, P1_U3067);
  nand ginst8897 (P1_U5384, P1_U3464, P1_U5373);
  nand ginst8898 (P1_U5385, P1_U3021, P1_U3060);
  nand ginst8899 (P1_U5386, P1_U3461, P1_U5373);
  nand ginst8900 (P1_U5387, P1_U3021, P1_U3064);
  nand ginst8901 (P1_U5388, P1_U3974, P1_U5373);
  nand ginst8902 (P1_U5389, P1_U3021, P1_U3054);
  nand ginst8903 (P1_U5390, P1_U3975, P1_U5373);
  nand ginst8904 (P1_U5391, P1_U3021, P1_U3053);
  nand ginst8905 (P1_U5392, P1_U3976, P1_U5373);
  nand ginst8906 (P1_U5393, P1_U3021, P1_U3057);
  nand ginst8907 (P1_U5394, P1_U3977, P1_U5373);
  nand ginst8908 (P1_U5395, P1_U3021, P1_U3058);
  nand ginst8909 (P1_U5396, P1_U3978, P1_U5373);
  nand ginst8910 (P1_U5397, P1_U3021, P1_U3065);
  nand ginst8911 (P1_U5398, P1_U3979, P1_U5373);
  nand ginst8912 (P1_U5399, P1_U3021, P1_U3066);
  nand ginst8913 (P1_U5400, P1_U3980, P1_U5373);
  nand ginst8914 (P1_U5401, P1_U3021, P1_U3061);
  nand ginst8915 (P1_U5402, P1_U3981, P1_U5373);
  nand ginst8916 (P1_U5403, P1_U3021, P1_U3075);
  nand ginst8917 (P1_U5404, P1_U3982, P1_U5373);
  nand ginst8918 (P1_U5405, P1_U3021, P1_U3076);
  nand ginst8919 (P1_U5406, P1_U3458, P1_U5373);
  nand ginst8920 (P1_U5407, P1_U3021, P1_U3068);
  nand ginst8921 (P1_U5408, P1_U3508, P1_U5373);
  nand ginst8922 (P1_U5409, P1_U3021, P1_U3081);
  nand ginst8923 (P1_U5410, P1_U3506, P1_U5373);
  nand ginst8924 (P1_U5411, P1_U3021, P1_U3082);
  nand ginst8925 (P1_U5412, P1_U3503, P1_U5373);
  nand ginst8926 (P1_U5413, P1_U3021, P1_U3069);
  nand ginst8927 (P1_U5414, P1_U3500, P1_U5373);
  nand ginst8928 (P1_U5415, P1_U3021, P1_U3073);
  nand ginst8929 (P1_U5416, P1_U3497, P1_U5373);
  nand ginst8930 (P1_U5417, P1_U3021, P1_U3074);
  nand ginst8931 (P1_U5418, P1_U3494, P1_U5373);
  nand ginst8932 (P1_U5419, P1_U3021, P1_U3079);
  nand ginst8933 (P1_U5420, P1_U3491, P1_U5373);
  nand ginst8934 (P1_U5421, P1_U3021, P1_U3080);
  nand ginst8935 (P1_U5422, P1_U3488, P1_U5373);
  nand ginst8936 (P1_U5423, P1_U3021, P1_U3072);
  nand ginst8937 (P1_U5424, P1_U3485, P1_U5373);
  nand ginst8938 (P1_U5425, P1_U3021, P1_U3063);
  nand ginst8939 (P1_U5426, P1_U3482, P1_U5373);
  nand ginst8940 (P1_U5427, P1_U3021, P1_U3062);
  nand ginst8941 (P1_U5428, P1_U3455, P1_U5373);
  nand ginst8942 (P1_U5429, P1_U3021, P1_U3078);
  nand ginst8943 (P1_U5430, P1_U3450, P1_U5373);
  nand ginst8944 (P1_U5431, P1_U3021, P1_U3077);
  nand ginst8945 (P1_U5432, P1_REG1_REG_0__SCAN_IN, P1_U4102);
  nand ginst8946 (P1_U5433, P1_U3021, P1_U3479);
  nand ginst8947 (P1_U5434, P1_U3083, P1_U3434);
  nand ginst8948 (P1_U5435, P1_U3021, P1_U3476);
  nand ginst8949 (P1_U5436, P1_U3084, P1_U3434);
  nand ginst8950 (P1_U5437, P1_U3021, P1_U3473);
  nand ginst8951 (P1_U5438, P1_U3070, P1_U3434);
  nand ginst8952 (P1_U5439, P1_U3021, P1_U3470);
  nand ginst8953 (P1_U5440, P1_U3071, P1_U3434);
  nand ginst8954 (P1_U5441, P1_U3021, P1_U3467);
  nand ginst8955 (P1_U5442, P1_U3067, P1_U3434);
  nand ginst8956 (P1_U5443, P1_U3021, P1_U3464);
  nand ginst8957 (P1_U5444, P1_U3060, P1_U3434);
  nand ginst8958 (P1_U5445, P1_U3021, P1_U3461);
  nand ginst8959 (P1_U5446, P1_U3064, P1_U3434);
  nand ginst8960 (P1_U5447, P1_U3021, P1_U3974);
  nand ginst8961 (P1_U5448, P1_U3054, P1_U3434);
  nand ginst8962 (P1_U5449, P1_U3021, P1_U3975);
  nand ginst8963 (P1_U5450, P1_U3053, P1_U3434);
  nand ginst8964 (P1_U5451, P1_U3021, P1_U3976);
  nand ginst8965 (P1_U5452, P1_U3057, P1_U3434);
  nand ginst8966 (P1_U5453, P1_U3021, P1_U3977);
  nand ginst8967 (P1_U5454, P1_U3058, P1_U3434);
  nand ginst8968 (P1_U5455, P1_U3021, P1_U3978);
  nand ginst8969 (P1_U5456, P1_U3065, P1_U3434);
  nand ginst8970 (P1_U5457, P1_U3021, P1_U3979);
  nand ginst8971 (P1_U5458, P1_U3066, P1_U3434);
  nand ginst8972 (P1_U5459, P1_U3021, P1_U3980);
  nand ginst8973 (P1_U5460, P1_U3061, P1_U3434);
  nand ginst8974 (P1_U5461, P1_U3021, P1_U3981);
  nand ginst8975 (P1_U5462, P1_U3075, P1_U3434);
  nand ginst8976 (P1_U5463, P1_U3021, P1_U3982);
  nand ginst8977 (P1_U5464, P1_U3076, P1_U3434);
  nand ginst8978 (P1_U5465, P1_U3021, P1_U3458);
  nand ginst8979 (P1_U5466, P1_U3068, P1_U3434);
  nand ginst8980 (P1_U5467, P1_U3021, P1_U3508);
  nand ginst8981 (P1_U5468, P1_U3081, P1_U3434);
  nand ginst8982 (P1_U5469, P1_U3021, P1_U3506);
  nand ginst8983 (P1_U5470, P1_U3082, P1_U3434);
  nand ginst8984 (P1_U5471, P1_U3021, P1_U3503);
  nand ginst8985 (P1_U5472, P1_U3069, P1_U3434);
  nand ginst8986 (P1_U5473, P1_U3021, P1_U3500);
  nand ginst8987 (P1_U5474, P1_U3073, P1_U3434);
  nand ginst8988 (P1_U5475, P1_U3021, P1_U3497);
  nand ginst8989 (P1_U5476, P1_U3074, P1_U3434);
  nand ginst8990 (P1_U5477, P1_U3021, P1_U3494);
  nand ginst8991 (P1_U5478, P1_U3079, P1_U3434);
  nand ginst8992 (P1_U5479, P1_U3021, P1_U3491);
  nand ginst8993 (P1_U5480, P1_U3080, P1_U3434);
  nand ginst8994 (P1_U5481, P1_U3021, P1_U3488);
  nand ginst8995 (P1_U5482, P1_U3072, P1_U3434);
  nand ginst8996 (P1_U5483, P1_U3021, P1_U3485);
  nand ginst8997 (P1_U5484, P1_U3063, P1_U3434);
  nand ginst8998 (P1_U5485, P1_U3021, P1_U3482);
  nand ginst8999 (P1_U5486, P1_U3062, P1_U3434);
  nand ginst9000 (P1_U5487, P1_U3021, P1_U3455);
  nand ginst9001 (P1_U5488, P1_U3078, P1_U3434);
  nand ginst9002 (P1_U5489, P1_U3021, P1_U3450);
  nand ginst9003 (P1_U5490, P1_U3077, P1_U3434);
  nand ginst9004 (P1_U5491, P1_U3448, P1_U4102);
  nand ginst9005 (P1_U5492, P1_U3426, P1_U3428);
  nand ginst9006 (P1_U5493, P1_U3479, P1_U3953);
  nand ginst9007 (P1_U5494, P1_U3586, P1_U5492);
  nand ginst9008 (P1_U5495, P1_U3476, P1_U3953);
  nand ginst9009 (P1_U5496, P1_U3587, P1_U5492);
  nand ginst9010 (P1_U5497, P1_U3473, P1_U3953);
  nand ginst9011 (P1_U5498, P1_U3588, P1_U5492);
  nand ginst9012 (P1_U5499, P1_U3470, P1_U3953);
  nand ginst9013 (P1_U5500, P1_U3589, P1_U5492);
  nand ginst9014 (P1_U5501, P1_U3467, P1_U3953);
  nand ginst9015 (P1_U5502, P1_U3590, P1_U5492);
  nand ginst9016 (P1_U5503, P1_U3464, P1_U3953);
  nand ginst9017 (P1_U5504, P1_U3591, P1_U5492);
  nand ginst9018 (P1_U5505, P1_U3593, P1_U5492);
  nand ginst9019 (P1_U5506, P1_U3953, P1_U3983);
  nand ginst9020 (P1_U5507, P1_U3594, P1_U5492);
  nand ginst9021 (P1_U5508, P1_U3953, P1_U3984);
  nand ginst9022 (P1_U5509, P1_U3461, P1_U3953);
  nand ginst9023 (P1_U5510, P1_U3592, P1_U5492);
  nand ginst9024 (P1_U5511, P1_U3596, P1_U5492);
  nand ginst9025 (P1_U5512, P1_U3953, P1_U3985);
  nand ginst9026 (P1_U5513, P1_U3597, P1_U5492);
  nand ginst9027 (P1_U5514, P1_U3953, P1_U3974);
  nand ginst9028 (P1_U5515, P1_U3598, P1_U5492);
  nand ginst9029 (P1_U5516, P1_U3953, P1_U3975);
  nand ginst9030 (P1_U5517, P1_U3599, P1_U5492);
  nand ginst9031 (P1_U5518, P1_U3953, P1_U3976);
  nand ginst9032 (P1_U5519, P1_U3600, P1_U5492);
  nand ginst9033 (P1_U5520, P1_U3953, P1_U3977);
  nand ginst9034 (P1_U5521, P1_U3601, P1_U5492);
  nand ginst9035 (P1_U5522, P1_U3953, P1_U3978);
  nand ginst9036 (P1_U5523, P1_U3602, P1_U5492);
  nand ginst9037 (P1_U5524, P1_U3953, P1_U3979);
  nand ginst9038 (P1_U5525, P1_U3603, P1_U5492);
  nand ginst9039 (P1_U5526, P1_U3953, P1_U3980);
  nand ginst9040 (P1_U5527, P1_U3604, P1_U5492);
  nand ginst9041 (P1_U5528, P1_U3953, P1_U3981);
  nand ginst9042 (P1_U5529, P1_U3605, P1_U5492);
  nand ginst9043 (P1_U5530, P1_U3953, P1_U3982);
  nand ginst9044 (P1_U5531, P1_U3458, P1_U3953);
  nand ginst9045 (P1_U5532, P1_U3595, P1_U5492);
  nand ginst9046 (P1_U5533, P1_U3508, P1_U3953);
  nand ginst9047 (P1_U5534, P1_U3607, P1_U5492);
  nand ginst9048 (P1_U5535, P1_U3506, P1_U3953);
  nand ginst9049 (P1_U5536, P1_U3608, P1_U5492);
  nand ginst9050 (P1_U5537, P1_U3503, P1_U3953);
  nand ginst9051 (P1_U5538, P1_U3609, P1_U5492);
  nand ginst9052 (P1_U5539, P1_U3500, P1_U3953);
  nand ginst9053 (P1_U5540, P1_U3610, P1_U5492);
  nand ginst9054 (P1_U5541, P1_U3497, P1_U3953);
  nand ginst9055 (P1_U5542, P1_U3611, P1_U5492);
  nand ginst9056 (P1_U5543, P1_U3494, P1_U3953);
  nand ginst9057 (P1_U5544, P1_U3612, P1_U5492);
  nand ginst9058 (P1_U5545, P1_U3491, P1_U3953);
  nand ginst9059 (P1_U5546, P1_U3613, P1_U5492);
  nand ginst9060 (P1_U5547, P1_U3488, P1_U3953);
  nand ginst9061 (P1_U5548, P1_U3614, P1_U5492);
  nand ginst9062 (P1_U5549, P1_U3485, P1_U3953);
  nand ginst9063 (P1_U5550, P1_U3615, P1_U5492);
  nand ginst9064 (P1_U5551, P1_U3482, P1_U3953);
  nand ginst9065 (P1_U5552, P1_U3616, P1_U5492);
  nand ginst9066 (P1_U5553, P1_U3455, P1_U3953);
  nand ginst9067 (P1_U5554, P1_U3606, P1_U5492);
  nand ginst9068 (P1_U5555, P1_U3450, P1_U3953);
  nand ginst9069 (P1_U5556, P1_U3617, P1_U5492);
  nand ginst9070 (P1_U5557, P1_U3479, P1_U5492);
  nand ginst9071 (P1_U5558, P1_U3586, P1_U3953);
  nand ginst9072 (P1_U5559, P1_U3084, P1_U5677);
  nand ginst9073 (P1_U5560, P1_U3476, P1_U5492);
  nand ginst9074 (P1_U5561, P1_U3587, P1_U3953);
  nand ginst9075 (P1_U5562, P1_U3070, P1_U5677);
  nand ginst9076 (P1_U5563, P1_U3473, P1_U5492);
  nand ginst9077 (P1_U5564, P1_U3588, P1_U3953);
  nand ginst9078 (P1_U5565, P1_U3071, P1_U5677);
  nand ginst9079 (P1_U5566, P1_U3470, P1_U5492);
  nand ginst9080 (P1_U5567, P1_U3589, P1_U3953);
  nand ginst9081 (P1_U5568, P1_U3067, P1_U5677);
  nand ginst9082 (P1_U5569, P1_U3467, P1_U5492);
  nand ginst9083 (P1_U5570, P1_U3590, P1_U3953);
  nand ginst9084 (P1_U5571, P1_U3060, P1_U5677);
  nand ginst9085 (P1_U5572, P1_U3464, P1_U5492);
  nand ginst9086 (P1_U5573, P1_U3591, P1_U3953);
  nand ginst9087 (P1_U5574, P1_U3064, P1_U5677);
  nand ginst9088 (P1_U5575, P1_U3983, P1_U5492);
  nand ginst9089 (P1_U5576, P1_U3593, P1_U3953);
  nand ginst9090 (P1_U5577, P1_U3984, P1_U5492);
  nand ginst9091 (P1_U5578, P1_U3594, P1_U3953);
  nand ginst9092 (P1_U5579, P1_U3461, P1_U5492);
  nand ginst9093 (P1_U5580, P1_U3592, P1_U3953);
  nand ginst9094 (P1_U5581, P1_U3068, P1_U5677);
  nand ginst9095 (P1_U5582, P1_U3985, P1_U5492);
  nand ginst9096 (P1_U5583, P1_U3596, P1_U3953);
  nand ginst9097 (P1_U5584, P1_U3054, P1_U5677);
  nand ginst9098 (P1_U5585, P1_U3974, P1_U5492);
  nand ginst9099 (P1_U5586, P1_U3597, P1_U3953);
  nand ginst9100 (P1_U5587, P1_U3053, P1_U5677);
  nand ginst9101 (P1_U5588, P1_U3975, P1_U5492);
  nand ginst9102 (P1_U5589, P1_U3598, P1_U3953);
  nand ginst9103 (P1_U5590, P1_U3057, P1_U5677);
  nand ginst9104 (P1_U5591, P1_U3976, P1_U5492);
  nand ginst9105 (P1_U5592, P1_U3599, P1_U3953);
  nand ginst9106 (P1_U5593, P1_U3058, P1_U5677);
  nand ginst9107 (P1_U5594, P1_U3977, P1_U5492);
  nand ginst9108 (P1_U5595, P1_U3600, P1_U3953);
  nand ginst9109 (P1_U5596, P1_U3065, P1_U5677);
  nand ginst9110 (P1_U5597, P1_U3978, P1_U5492);
  nand ginst9111 (P1_U5598, P1_U3601, P1_U3953);
  nand ginst9112 (P1_U5599, P1_U3066, P1_U5677);
  nand ginst9113 (P1_U5600, P1_U3979, P1_U5492);
  nand ginst9114 (P1_U5601, P1_U3602, P1_U3953);
  nand ginst9115 (P1_U5602, P1_U3061, P1_U5677);
  nand ginst9116 (P1_U5603, P1_U3980, P1_U5492);
  nand ginst9117 (P1_U5604, P1_U3603, P1_U3953);
  nand ginst9118 (P1_U5605, P1_U3075, P1_U5677);
  nand ginst9119 (P1_U5606, P1_U3981, P1_U5492);
  nand ginst9120 (P1_U5607, P1_U3604, P1_U3953);
  nand ginst9121 (P1_U5608, P1_U3076, P1_U5677);
  nand ginst9122 (P1_U5609, P1_U3982, P1_U5492);
  nand ginst9123 (P1_U5610, P1_U3605, P1_U3953);
  nand ginst9124 (P1_U5611, P1_U3081, P1_U5677);
  nand ginst9125 (P1_U5612, P1_U3458, P1_U5492);
  nand ginst9126 (P1_U5613, P1_U3595, P1_U3953);
  nand ginst9127 (P1_U5614, P1_U3078, P1_U5677);
  nand ginst9128 (P1_U5615, P1_U3508, P1_U5492);
  nand ginst9129 (P1_U5616, P1_U3607, P1_U3953);
  nand ginst9130 (P1_U5617, P1_U3082, P1_U5677);
  nand ginst9131 (P1_U5618, P1_U3506, P1_U5492);
  nand ginst9132 (P1_U5619, P1_U3608, P1_U3953);
  nand ginst9133 (P1_U5620, P1_U3069, P1_U5677);
  nand ginst9134 (P1_U5621, P1_U3503, P1_U5492);
  nand ginst9135 (P1_U5622, P1_U3609, P1_U3953);
  nand ginst9136 (P1_U5623, P1_U3073, P1_U5677);
  nand ginst9137 (P1_U5624, P1_U3500, P1_U5492);
  nand ginst9138 (P1_U5625, P1_U3610, P1_U3953);
  nand ginst9139 (P1_U5626, P1_U3074, P1_U5677);
  nand ginst9140 (P1_U5627, P1_U3497, P1_U5492);
  nand ginst9141 (P1_U5628, P1_U3611, P1_U3953);
  nand ginst9142 (P1_U5629, P1_U3079, P1_U5677);
  nand ginst9143 (P1_U5630, P1_U3494, P1_U5492);
  nand ginst9144 (P1_U5631, P1_U3612, P1_U3953);
  nand ginst9145 (P1_U5632, P1_U3080, P1_U5677);
  nand ginst9146 (P1_U5633, P1_U3491, P1_U5492);
  nand ginst9147 (P1_U5634, P1_U3613, P1_U3953);
  nand ginst9148 (P1_U5635, P1_U3072, P1_U5677);
  nand ginst9149 (P1_U5636, P1_U3488, P1_U5492);
  nand ginst9150 (P1_U5637, P1_U3614, P1_U3953);
  nand ginst9151 (P1_U5638, P1_U3063, P1_U5677);
  nand ginst9152 (P1_U5639, P1_U3485, P1_U5492);
  nand ginst9153 (P1_U5640, P1_U3615, P1_U3953);
  nand ginst9154 (P1_U5641, P1_U3062, P1_U5677);
  nand ginst9155 (P1_U5642, P1_U3482, P1_U5492);
  nand ginst9156 (P1_U5643, P1_U3616, P1_U3953);
  nand ginst9157 (P1_U5644, P1_U3083, P1_U5677);
  nand ginst9158 (P1_U5645, P1_U3455, P1_U5492);
  nand ginst9159 (P1_U5646, P1_U3606, P1_U3953);
  nand ginst9160 (P1_U5647, P1_U3077, P1_U5677);
  nand ginst9161 (P1_U5648, P1_U3450, P1_U5492);
  nand ginst9162 (P1_U5649, P1_U3617, P1_U3953);
  nand ginst9163 (P1_U5650, P1_U3052, P1_U3864, P1_U3950, P1_U5662);
  nand ginst9164 (P1_U5651, P1_U3086, P1_U5091);
  nand ginst9165 (P1_U5652, P1_U3865, P1_U5090, P1_U5091);
  nand ginst9166 (P1_U5653, P1_U3430, P1_U3997);
  nand ginst9167 (P1_U5654, P1_U3972, P1_U3997);
  nand ginst9168 (P1_U5655, P1_U3995, P1_U5653);
  nand ginst9169 (P1_U5656, P1_U3996, P1_U5654);
  nand ginst9170 (P1_U5657, P1_R1207_U14, P1_U3958);
  nand ginst9171 (P1_U5658, P1_R1192_U14, P1_U3959);
  nand ginst9172 (P1_U5659, P1_R1150_U14, P1_U3961);
  nand ginst9173 (P1_U5660, P1_R1117_U14, P1_U3963);
  nand ginst9174 (P1_U5661, P1_U5666, P1_U5672);
  nand ginst9175 (P1_U5662, P1_U5693, P1_U6169, P1_U6170);
  nand ginst9176 (P1_U5663, P1_U3438, P1_U3442);
  nand ginst9177 (P1_U5664, P1_IR_REG_24__SCAN_IN, P1_U3910);
  nand ginst9178 (P1_U5665, P1_IR_REG_31__SCAN_IN, P1_SUB_84_U17);
  not ginst9179 (P1_U5666, P1_U3435);
  nand ginst9180 (P1_U5667, P1_IR_REG_25__SCAN_IN, P1_U3910);
  nand ginst9181 (P1_U5668, P1_IR_REG_31__SCAN_IN, P1_SUB_84_U170);
  not ginst9182 (P1_U5669, P1_U3436);
  nand ginst9183 (P1_U5670, P1_IR_REG_26__SCAN_IN, P1_U3910);
  nand ginst9184 (P1_U5671, P1_IR_REG_31__SCAN_IN, P1_SUB_84_U18);
  not ginst9185 (P1_U5672, P1_U3437);
  nand ginst9186 (P1_U5673, P1_U3050, P1_U3359);
  nand ginst9187 (P1_U5674, P1_B_REG_SCAN_IN, P1_U4003, P1_U5666);
  nand ginst9188 (P1_U5675, P1_IR_REG_23__SCAN_IN, P1_U3910);
  nand ginst9189 (P1_U5676, P1_IR_REG_31__SCAN_IN, P1_SUB_84_U16);
  not ginst9190 (P1_U5677, P1_U3438);
  nand ginst9191 (P1_U5678, P1_D_REG_0__SCAN_IN, P1_U3911);
  nand ginst9192 (P1_U5679, P1_U3992, P1_U4103);
  nand ginst9193 (P1_U5680, P1_D_REG_1__SCAN_IN, P1_U3911);
  nand ginst9194 (P1_U5681, P1_U3992, P1_U4104);
  nand ginst9195 (P1_U5682, P1_IR_REG_22__SCAN_IN, P1_U3910);
  nand ginst9196 (P1_U5683, P1_IR_REG_31__SCAN_IN, P1_SUB_84_U15);
  not ginst9197 (P1_U5684, P1_U3443);
  nand ginst9198 (P1_U5685, P1_IR_REG_19__SCAN_IN, P1_U3910);
  nand ginst9199 (P1_U5686, P1_IR_REG_31__SCAN_IN, P1_SUB_84_U13);
  not ginst9200 (P1_U5687, P1_U3442);
  nand ginst9201 (P1_U5688, P1_IR_REG_20__SCAN_IN, P1_U3910);
  nand ginst9202 (P1_U5689, P1_IR_REG_31__SCAN_IN, P1_SUB_84_U14);
  not ginst9203 (P1_U5690, P1_U3441);
  nand ginst9204 (P1_U5691, P1_IR_REG_21__SCAN_IN, P1_U3910);
  nand ginst9205 (P1_U5692, P1_IR_REG_31__SCAN_IN, P1_SUB_84_U173);
  not ginst9206 (P1_U5693, P1_U3447);
  nand ginst9207 (P1_U5694, P1_IR_REG_0__SCAN_IN, P1_U3910);
  nand ginst9208 (P1_U5695, P1_IR_REG_0__SCAN_IN, P1_IR_REG_31__SCAN_IN);
  not ginst9209 (P1_U5696, P1_U3448);
  nand ginst9210 (P1_U5697, P1_IR_REG_28__SCAN_IN, P1_U3910);
  nand ginst9211 (P1_U5698, P1_IR_REG_31__SCAN_IN, P1_SUB_84_U19);
  not ginst9212 (P1_U5699, P1_U3446);
  nand ginst9213 (P1_U5700, P1_IR_REG_27__SCAN_IN, P1_U3910);
  nand ginst9214 (P1_U5701, P1_IR_REG_31__SCAN_IN, P1_SUB_84_U42);
  not ginst9215 (P1_U5702, P1_U3449);
  nand ginst9216 (P1_U5703, P1_U3912, U88);
  nand ginst9217 (P1_U5704, P1_U3448, P1_U3971);
  not ginst9218 (P1_U5705, P1_U3450);
  nand ginst9219 (P1_U5706, P1_IR_REG_30__SCAN_IN, P1_U3910);
  nand ginst9220 (P1_U5707, P1_IR_REG_31__SCAN_IN, P1_SUB_84_U165);
  not ginst9221 (P1_U5708, P1_U3444);
  nand ginst9222 (P1_U5709, P1_IR_REG_29__SCAN_IN, P1_U3910);
  nand ginst9223 (P1_U5710, P1_IR_REG_31__SCAN_IN, P1_SUB_84_U20);
  not ginst9224 (P1_U5711, P1_U3445);
  nand ginst9225 (P1_U5712, P1_U3443, P1_U5693);
  nand ginst9226 (P1_U5713, P1_U4135, P1_U5684);
  nand ginst9227 (P1_U5714, P1_D_REG_1__SCAN_IN, P1_U4101);
  nand ginst9228 (P1_U5715, P1_U3360, P1_U4104);
  not ginst9229 (P1_U5716, P1_U3452);
  nand ginst9230 (P1_U5717, P1_U3360, P1_U5661);
  nand ginst9231 (P1_U5718, P1_D_REG_0__SCAN_IN, P1_U4101);
  not ginst9232 (P1_U5719, P1_U3451);
  nand ginst9233 (P1_U5720, P1_REG0_REG_0__SCAN_IN, P1_U3913);
  nand ginst9234 (P1_U5721, P1_U3991, P1_U4155);
  nand ginst9235 (P1_U5722, P1_IR_REG_1__SCAN_IN, P1_U3910);
  nand ginst9236 (P1_U5723, P1_IR_REG_31__SCAN_IN, P1_SUB_84_U40);
  nand ginst9237 (P1_U5724, P1_U3912, U77);
  nand ginst9238 (P1_U5725, P1_U3454, P1_U3971);
  not ginst9239 (P1_U5726, P1_U3455);
  nand ginst9240 (P1_U5727, P1_REG0_REG_1__SCAN_IN, P1_U3913);
  nand ginst9241 (P1_U5728, P1_U3991, P1_U4179);
  nand ginst9242 (P1_U5729, P1_IR_REG_2__SCAN_IN, P1_U3910);
  nand ginst9243 (P1_U5730, P1_IR_REG_31__SCAN_IN, P1_SUB_84_U21);
  nand ginst9244 (P1_U5731, P1_U3912, U66);
  nand ginst9245 (P1_U5732, P1_U3457, P1_U3971);
  not ginst9246 (P1_U5733, P1_U3458);
  nand ginst9247 (P1_U5734, P1_REG0_REG_2__SCAN_IN, P1_U3913);
  nand ginst9248 (P1_U5735, P1_U3991, P1_U4198);
  nand ginst9249 (P1_U5736, P1_IR_REG_3__SCAN_IN, P1_U3910);
  nand ginst9250 (P1_U5737, P1_IR_REG_31__SCAN_IN, P1_SUB_84_U22);
  nand ginst9251 (P1_U5738, P1_U3912, U63);
  nand ginst9252 (P1_U5739, P1_U3460, P1_U3971);
  not ginst9253 (P1_U5740, P1_U3461);
  nand ginst9254 (P1_U5741, P1_REG0_REG_3__SCAN_IN, P1_U3913);
  nand ginst9255 (P1_U5742, P1_U3991, P1_U4217);
  nand ginst9256 (P1_U5743, P1_IR_REG_4__SCAN_IN, P1_U3910);
  nand ginst9257 (P1_U5744, P1_IR_REG_31__SCAN_IN, P1_SUB_84_U23);
  nand ginst9258 (P1_U5745, P1_U3912, U62);
  nand ginst9259 (P1_U5746, P1_U3463, P1_U3971);
  not ginst9260 (P1_U5747, P1_U3464);
  nand ginst9261 (P1_U5748, P1_REG0_REG_4__SCAN_IN, P1_U3913);
  nand ginst9262 (P1_U5749, P1_U3991, P1_U4236);
  nand ginst9263 (P1_U5750, P1_IR_REG_5__SCAN_IN, P1_U3910);
  nand ginst9264 (P1_U5751, P1_IR_REG_31__SCAN_IN, P1_SUB_84_U162);
  nand ginst9265 (P1_U5752, P1_U3912, U61);
  nand ginst9266 (P1_U5753, P1_U3466, P1_U3971);
  not ginst9267 (P1_U5754, P1_U3467);
  nand ginst9268 (P1_U5755, P1_REG0_REG_5__SCAN_IN, P1_U3913);
  nand ginst9269 (P1_U5756, P1_U3991, P1_U4255);
  nand ginst9270 (P1_U5757, P1_IR_REG_6__SCAN_IN, P1_U3910);
  nand ginst9271 (P1_U5758, P1_IR_REG_31__SCAN_IN, P1_SUB_84_U24);
  nand ginst9272 (P1_U5759, P1_U3912, U60);
  nand ginst9273 (P1_U5760, P1_U3469, P1_U3971);
  not ginst9274 (P1_U5761, P1_U3470);
  nand ginst9275 (P1_U5762, P1_REG0_REG_6__SCAN_IN, P1_U3913);
  nand ginst9276 (P1_U5763, P1_U3991, P1_U4274);
  nand ginst9277 (P1_U5764, P1_IR_REG_7__SCAN_IN, P1_U3910);
  nand ginst9278 (P1_U5765, P1_IR_REG_31__SCAN_IN, P1_SUB_84_U25);
  nand ginst9279 (P1_U5766, P1_U3912, U59);
  nand ginst9280 (P1_U5767, P1_U3472, P1_U3971);
  not ginst9281 (P1_U5768, P1_U3473);
  nand ginst9282 (P1_U5769, P1_REG0_REG_7__SCAN_IN, P1_U3913);
  nand ginst9283 (P1_U5770, P1_U3991, P1_U4293);
  nand ginst9284 (P1_U5771, P1_IR_REG_8__SCAN_IN, P1_U3910);
  nand ginst9285 (P1_U5772, P1_IR_REG_31__SCAN_IN, P1_SUB_84_U26);
  nand ginst9286 (P1_U5773, P1_U3912, U58);
  nand ginst9287 (P1_U5774, P1_U3475, P1_U3971);
  not ginst9288 (P1_U5775, P1_U3476);
  nand ginst9289 (P1_U5776, P1_REG0_REG_8__SCAN_IN, P1_U3913);
  nand ginst9290 (P1_U5777, P1_U3991, P1_U4312);
  nand ginst9291 (P1_U5778, P1_IR_REG_9__SCAN_IN, P1_U3910);
  nand ginst9292 (P1_U5779, P1_IR_REG_31__SCAN_IN, P1_SUB_84_U160);
  nand ginst9293 (P1_U5780, P1_U3912, U57);
  nand ginst9294 (P1_U5781, P1_U3478, P1_U3971);
  not ginst9295 (P1_U5782, P1_U3479);
  nand ginst9296 (P1_U5783, P1_REG0_REG_9__SCAN_IN, P1_U3913);
  nand ginst9297 (P1_U5784, P1_U3991, P1_U4331);
  nand ginst9298 (P1_U5785, P1_IR_REG_10__SCAN_IN, P1_U3910);
  nand ginst9299 (P1_U5786, P1_IR_REG_31__SCAN_IN, P1_SUB_84_U6);
  nand ginst9300 (P1_U5787, P1_U3912, U87);
  nand ginst9301 (P1_U5788, P1_U3481, P1_U3971);
  not ginst9302 (P1_U5789, P1_U3482);
  nand ginst9303 (P1_U5790, P1_REG0_REG_10__SCAN_IN, P1_U3913);
  nand ginst9304 (P1_U5791, P1_U3991, P1_U4350);
  nand ginst9305 (P1_U5792, P1_IR_REG_11__SCAN_IN, P1_U3910);
  nand ginst9306 (P1_U5793, P1_IR_REG_31__SCAN_IN, P1_SUB_84_U7);
  nand ginst9307 (P1_U5794, P1_U3912, U86);
  nand ginst9308 (P1_U5795, P1_U3484, P1_U3971);
  not ginst9309 (P1_U5796, P1_U3485);
  nand ginst9310 (P1_U5797, P1_REG0_REG_11__SCAN_IN, P1_U3913);
  nand ginst9311 (P1_U5798, P1_U3991, P1_U4369);
  nand ginst9312 (P1_U5799, P1_IR_REG_12__SCAN_IN, P1_U3910);
  nand ginst9313 (P1_U5800, P1_IR_REG_31__SCAN_IN, P1_SUB_84_U8);
  nand ginst9314 (P1_U5801, P1_U3912, U85);
  nand ginst9315 (P1_U5802, P1_U3487, P1_U3971);
  not ginst9316 (P1_U5803, P1_U3488);
  nand ginst9317 (P1_U5804, P1_REG0_REG_12__SCAN_IN, P1_U3913);
  nand ginst9318 (P1_U5805, P1_U3991, P1_U4388);
  nand ginst9319 (P1_U5806, P1_IR_REG_13__SCAN_IN, P1_U3910);
  nand ginst9320 (P1_U5807, P1_IR_REG_31__SCAN_IN, P1_SUB_84_U179);
  nand ginst9321 (P1_U5808, P1_U3912, U84);
  nand ginst9322 (P1_U5809, P1_U3490, P1_U3971);
  not ginst9323 (P1_U5810, P1_U3491);
  nand ginst9324 (P1_U5811, P1_REG0_REG_13__SCAN_IN, P1_U3913);
  nand ginst9325 (P1_U5812, P1_U3991, P1_U4407);
  nand ginst9326 (P1_U5813, P1_IR_REG_14__SCAN_IN, P1_U3910);
  nand ginst9327 (P1_U5814, P1_IR_REG_31__SCAN_IN, P1_SUB_84_U9);
  nand ginst9328 (P1_U5815, P1_U3912, U83);
  nand ginst9329 (P1_U5816, P1_U3493, P1_U3971);
  not ginst9330 (P1_U5817, P1_U3494);
  nand ginst9331 (P1_U5818, P1_REG0_REG_14__SCAN_IN, P1_U3913);
  nand ginst9332 (P1_U5819, P1_U3991, P1_U4426);
  nand ginst9333 (P1_U5820, P1_IR_REG_15__SCAN_IN, P1_U3910);
  nand ginst9334 (P1_U5821, P1_IR_REG_31__SCAN_IN, P1_SUB_84_U10);
  nand ginst9335 (P1_U5822, P1_U3912, U82);
  nand ginst9336 (P1_U5823, P1_U3496, P1_U3971);
  not ginst9337 (P1_U5824, P1_U3497);
  nand ginst9338 (P1_U5825, P1_REG0_REG_15__SCAN_IN, P1_U3913);
  nand ginst9339 (P1_U5826, P1_U3991, P1_U4445);
  nand ginst9340 (P1_U5827, P1_IR_REG_16__SCAN_IN, P1_U3910);
  nand ginst9341 (P1_U5828, P1_IR_REG_31__SCAN_IN, P1_SUB_84_U11);
  nand ginst9342 (P1_U5829, P1_U3912, U81);
  nand ginst9343 (P1_U5830, P1_U3499, P1_U3971);
  not ginst9344 (P1_U5831, P1_U3500);
  nand ginst9345 (P1_U5832, P1_REG0_REG_16__SCAN_IN, P1_U3913);
  nand ginst9346 (P1_U5833, P1_U3991, P1_U4464);
  nand ginst9347 (P1_U5834, P1_IR_REG_17__SCAN_IN, P1_U3910);
  nand ginst9348 (P1_U5835, P1_IR_REG_31__SCAN_IN, P1_SUB_84_U177);
  nand ginst9349 (P1_U5836, P1_U3912, U80);
  nand ginst9350 (P1_U5837, P1_U3502, P1_U3971);
  not ginst9351 (P1_U5838, P1_U3503);
  nand ginst9352 (P1_U5839, P1_REG0_REG_17__SCAN_IN, P1_U3913);
  nand ginst9353 (P1_U5840, P1_U3991, P1_U4483);
  nand ginst9354 (P1_U5841, P1_IR_REG_18__SCAN_IN, P1_U3910);
  nand ginst9355 (P1_U5842, P1_IR_REG_31__SCAN_IN, P1_SUB_84_U12);
  nand ginst9356 (P1_U5843, P1_U3912, U79);
  nand ginst9357 (P1_U5844, P1_U3505, P1_U3971);
  not ginst9358 (P1_U5845, P1_U3506);
  nand ginst9359 (P1_U5846, P1_REG0_REG_18__SCAN_IN, P1_U3913);
  nand ginst9360 (P1_U5847, P1_U3991, P1_U4502);
  nand ginst9361 (P1_U5848, P1_U3912, U78);
  nand ginst9362 (P1_U5849, P1_U3442, P1_U3971);
  not ginst9363 (P1_U5850, P1_U3508);
  nand ginst9364 (P1_U5851, P1_REG0_REG_19__SCAN_IN, P1_U3913);
  nand ginst9365 (P1_U5852, P1_U3991, P1_U4521);
  nand ginst9366 (P1_U5853, P1_REG0_REG_20__SCAN_IN, P1_U3913);
  nand ginst9367 (P1_U5854, P1_U3991, P1_U4540);
  nand ginst9368 (P1_U5855, P1_REG0_REG_21__SCAN_IN, P1_U3913);
  nand ginst9369 (P1_U5856, P1_U3991, P1_U4559);
  nand ginst9370 (P1_U5857, P1_REG0_REG_22__SCAN_IN, P1_U3913);
  nand ginst9371 (P1_U5858, P1_U3991, P1_U4578);
  nand ginst9372 (P1_U5859, P1_REG0_REG_23__SCAN_IN, P1_U3913);
  nand ginst9373 (P1_U5860, P1_U3991, P1_U4597);
  nand ginst9374 (P1_U5861, P1_REG0_REG_24__SCAN_IN, P1_U3913);
  nand ginst9375 (P1_U5862, P1_U3991, P1_U4616);
  nand ginst9376 (P1_U5863, P1_REG0_REG_25__SCAN_IN, P1_U3913);
  nand ginst9377 (P1_U5864, P1_U3991, P1_U4635);
  nand ginst9378 (P1_U5865, P1_REG0_REG_26__SCAN_IN, P1_U3913);
  nand ginst9379 (P1_U5866, P1_U3991, P1_U4654);
  nand ginst9380 (P1_U5867, P1_REG0_REG_27__SCAN_IN, P1_U3913);
  nand ginst9381 (P1_U5868, P1_U3991, P1_U4673);
  nand ginst9382 (P1_U5869, P1_REG0_REG_28__SCAN_IN, P1_U3913);
  nand ginst9383 (P1_U5870, P1_U3991, P1_U4692);
  nand ginst9384 (P1_U5871, P1_REG0_REG_29__SCAN_IN, P1_U3913);
  nand ginst9385 (P1_U5872, P1_U3991, P1_U4712);
  nand ginst9386 (P1_U5873, P1_REG0_REG_30__SCAN_IN, P1_U3913);
  nand ginst9387 (P1_U5874, P1_U3991, P1_U4719);
  nand ginst9388 (P1_U5875, P1_REG0_REG_31__SCAN_IN, P1_U3913);
  nand ginst9389 (P1_U5876, P1_U3991, P1_U4722);
  nand ginst9390 (P1_U5877, P1_REG1_REG_0__SCAN_IN, P1_U3914);
  nand ginst9391 (P1_U5878, P1_U3990, P1_U4155);
  nand ginst9392 (P1_U5879, P1_REG1_REG_1__SCAN_IN, P1_U3914);
  nand ginst9393 (P1_U5880, P1_U3990, P1_U4179);
  nand ginst9394 (P1_U5881, P1_REG1_REG_2__SCAN_IN, P1_U3914);
  nand ginst9395 (P1_U5882, P1_U3990, P1_U4198);
  nand ginst9396 (P1_U5883, P1_REG1_REG_3__SCAN_IN, P1_U3914);
  nand ginst9397 (P1_U5884, P1_U3990, P1_U4217);
  nand ginst9398 (P1_U5885, P1_REG1_REG_4__SCAN_IN, P1_U3914);
  nand ginst9399 (P1_U5886, P1_U3990, P1_U4236);
  nand ginst9400 (P1_U5887, P1_REG1_REG_5__SCAN_IN, P1_U3914);
  nand ginst9401 (P1_U5888, P1_U3990, P1_U4255);
  nand ginst9402 (P1_U5889, P1_REG1_REG_6__SCAN_IN, P1_U3914);
  nand ginst9403 (P1_U5890, P1_U3990, P1_U4274);
  nand ginst9404 (P1_U5891, P1_REG1_REG_7__SCAN_IN, P1_U3914);
  nand ginst9405 (P1_U5892, P1_U3990, P1_U4293);
  nand ginst9406 (P1_U5893, P1_REG1_REG_8__SCAN_IN, P1_U3914);
  nand ginst9407 (P1_U5894, P1_U3990, P1_U4312);
  nand ginst9408 (P1_U5895, P1_REG1_REG_9__SCAN_IN, P1_U3914);
  nand ginst9409 (P1_U5896, P1_U3990, P1_U4331);
  nand ginst9410 (P1_U5897, P1_REG1_REG_10__SCAN_IN, P1_U3914);
  nand ginst9411 (P1_U5898, P1_U3990, P1_U4350);
  nand ginst9412 (P1_U5899, P1_REG1_REG_11__SCAN_IN, P1_U3914);
  nand ginst9413 (P1_U5900, P1_U3990, P1_U4369);
  nand ginst9414 (P1_U5901, P1_REG1_REG_12__SCAN_IN, P1_U3914);
  nand ginst9415 (P1_U5902, P1_U3990, P1_U4388);
  nand ginst9416 (P1_U5903, P1_REG1_REG_13__SCAN_IN, P1_U3914);
  nand ginst9417 (P1_U5904, P1_U3990, P1_U4407);
  nand ginst9418 (P1_U5905, P1_REG1_REG_14__SCAN_IN, P1_U3914);
  nand ginst9419 (P1_U5906, P1_U3990, P1_U4426);
  nand ginst9420 (P1_U5907, P1_REG1_REG_15__SCAN_IN, P1_U3914);
  nand ginst9421 (P1_U5908, P1_U3990, P1_U4445);
  nand ginst9422 (P1_U5909, P1_REG1_REG_16__SCAN_IN, P1_U3914);
  nand ginst9423 (P1_U5910, P1_U3990, P1_U4464);
  nand ginst9424 (P1_U5911, P1_REG1_REG_17__SCAN_IN, P1_U3914);
  nand ginst9425 (P1_U5912, P1_U3990, P1_U4483);
  nand ginst9426 (P1_U5913, P1_REG1_REG_18__SCAN_IN, P1_U3914);
  nand ginst9427 (P1_U5914, P1_U3990, P1_U4502);
  nand ginst9428 (P1_U5915, P1_REG1_REG_19__SCAN_IN, P1_U3914);
  nand ginst9429 (P1_U5916, P1_U3990, P1_U4521);
  nand ginst9430 (P1_U5917, P1_REG1_REG_20__SCAN_IN, P1_U3914);
  nand ginst9431 (P1_U5918, P1_U3990, P1_U4540);
  nand ginst9432 (P1_U5919, P1_REG1_REG_21__SCAN_IN, P1_U3914);
  nand ginst9433 (P1_U5920, P1_U3990, P1_U4559);
  nand ginst9434 (P1_U5921, P1_REG1_REG_22__SCAN_IN, P1_U3914);
  nand ginst9435 (P1_U5922, P1_U3990, P1_U4578);
  nand ginst9436 (P1_U5923, P1_REG1_REG_23__SCAN_IN, P1_U3914);
  nand ginst9437 (P1_U5924, P1_U3990, P1_U4597);
  nand ginst9438 (P1_U5925, P1_REG1_REG_24__SCAN_IN, P1_U3914);
  nand ginst9439 (P1_U5926, P1_U3990, P1_U4616);
  nand ginst9440 (P1_U5927, P1_REG1_REG_25__SCAN_IN, P1_U3914);
  nand ginst9441 (P1_U5928, P1_U3990, P1_U4635);
  nand ginst9442 (P1_U5929, P1_REG1_REG_26__SCAN_IN, P1_U3914);
  nand ginst9443 (P1_U5930, P1_U3990, P1_U4654);
  nand ginst9444 (P1_U5931, P1_REG1_REG_27__SCAN_IN, P1_U3914);
  nand ginst9445 (P1_U5932, P1_U3990, P1_U4673);
  nand ginst9446 (P1_U5933, P1_REG1_REG_28__SCAN_IN, P1_U3914);
  nand ginst9447 (P1_U5934, P1_U3990, P1_U4692);
  nand ginst9448 (P1_U5935, P1_REG1_REG_29__SCAN_IN, P1_U3914);
  nand ginst9449 (P1_U5936, P1_U3990, P1_U4712);
  nand ginst9450 (P1_U5937, P1_REG1_REG_30__SCAN_IN, P1_U3914);
  nand ginst9451 (P1_U5938, P1_U3990, P1_U4719);
  nand ginst9452 (P1_U5939, P1_REG1_REG_31__SCAN_IN, P1_U3914);
  nand ginst9453 (P1_U5940, P1_U3990, P1_U4722);
  nand ginst9454 (P1_U5941, P1_REG2_REG_0__SCAN_IN, P1_U3417);
  nand ginst9455 (P1_U5942, P1_U3374, P1_U3989);
  nand ginst9456 (P1_U5943, P1_REG2_REG_1__SCAN_IN, P1_U3417);
  nand ginst9457 (P1_U5944, P1_U3376, P1_U3989);
  nand ginst9458 (P1_U5945, P1_REG2_REG_2__SCAN_IN, P1_U3417);
  nand ginst9459 (P1_U5946, P1_U3377, P1_U3989);
  nand ginst9460 (P1_U5947, P1_REG2_REG_3__SCAN_IN, P1_U3417);
  nand ginst9461 (P1_U5948, P1_U3378, P1_U3989);
  nand ginst9462 (P1_U5949, P1_REG2_REG_4__SCAN_IN, P1_U3417);
  nand ginst9463 (P1_U5950, P1_U3379, P1_U3989);
  nand ginst9464 (P1_U5951, P1_REG2_REG_5__SCAN_IN, P1_U3417);
  nand ginst9465 (P1_U5952, P1_U3380, P1_U3989);
  nand ginst9466 (P1_U5953, P1_REG2_REG_6__SCAN_IN, P1_U3417);
  nand ginst9467 (P1_U5954, P1_U3381, P1_U3989);
  nand ginst9468 (P1_U5955, P1_REG2_REG_7__SCAN_IN, P1_U3417);
  nand ginst9469 (P1_U5956, P1_U3382, P1_U3989);
  nand ginst9470 (P1_U5957, P1_REG2_REG_8__SCAN_IN, P1_U3417);
  nand ginst9471 (P1_U5958, P1_U3383, P1_U3989);
  nand ginst9472 (P1_U5959, P1_REG2_REG_9__SCAN_IN, P1_U3417);
  nand ginst9473 (P1_U5960, P1_U3384, P1_U3989);
  nand ginst9474 (P1_U5961, P1_REG2_REG_10__SCAN_IN, P1_U3417);
  nand ginst9475 (P1_U5962, P1_U3385, P1_U3989);
  nand ginst9476 (P1_U5963, P1_REG2_REG_11__SCAN_IN, P1_U3417);
  nand ginst9477 (P1_U5964, P1_U3386, P1_U3989);
  nand ginst9478 (P1_U5965, P1_REG2_REG_12__SCAN_IN, P1_U3417);
  nand ginst9479 (P1_U5966, P1_U3387, P1_U3989);
  nand ginst9480 (P1_U5967, P1_REG2_REG_13__SCAN_IN, P1_U3417);
  nand ginst9481 (P1_U5968, P1_U3388, P1_U3989);
  nand ginst9482 (P1_U5969, P1_REG2_REG_14__SCAN_IN, P1_U3417);
  nand ginst9483 (P1_U5970, P1_U3389, P1_U3989);
  nand ginst9484 (P1_U5971, P1_REG2_REG_15__SCAN_IN, P1_U3417);
  nand ginst9485 (P1_U5972, P1_U3390, P1_U3989);
  nand ginst9486 (P1_U5973, P1_REG2_REG_16__SCAN_IN, P1_U3417);
  nand ginst9487 (P1_U5974, P1_U3391, P1_U3989);
  nand ginst9488 (P1_U5975, P1_REG2_REG_17__SCAN_IN, P1_U3417);
  nand ginst9489 (P1_U5976, P1_U3392, P1_U3989);
  nand ginst9490 (P1_U5977, P1_REG2_REG_18__SCAN_IN, P1_U3417);
  nand ginst9491 (P1_U5978, P1_U3393, P1_U3989);
  nand ginst9492 (P1_U5979, P1_REG2_REG_19__SCAN_IN, P1_U3417);
  nand ginst9493 (P1_U5980, P1_U3394, P1_U3989);
  nand ginst9494 (P1_U5981, P1_REG2_REG_20__SCAN_IN, P1_U3417);
  nand ginst9495 (P1_U5982, P1_U3396, P1_U3989);
  nand ginst9496 (P1_U5983, P1_REG2_REG_21__SCAN_IN, P1_U3417);
  nand ginst9497 (P1_U5984, P1_U3398, P1_U3989);
  nand ginst9498 (P1_U5985, P1_REG2_REG_22__SCAN_IN, P1_U3417);
  nand ginst9499 (P1_U5986, P1_U3400, P1_U3989);
  nand ginst9500 (P1_U5987, P1_REG2_REG_23__SCAN_IN, P1_U3417);
  nand ginst9501 (P1_U5988, P1_U3402, P1_U3989);
  nand ginst9502 (P1_U5989, P1_REG2_REG_24__SCAN_IN, P1_U3417);
  nand ginst9503 (P1_U5990, P1_U3404, P1_U3989);
  nand ginst9504 (P1_U5991, P1_REG2_REG_25__SCAN_IN, P1_U3417);
  nand ginst9505 (P1_U5992, P1_U3406, P1_U3989);
  nand ginst9506 (P1_U5993, P1_REG2_REG_26__SCAN_IN, P1_U3417);
  nand ginst9507 (P1_U5994, P1_U3408, P1_U3989);
  nand ginst9508 (P1_U5995, P1_REG2_REG_27__SCAN_IN, P1_U3417);
  nand ginst9509 (P1_U5996, P1_U3410, P1_U3989);
  nand ginst9510 (P1_U5997, P1_REG2_REG_28__SCAN_IN, P1_U3417);
  nand ginst9511 (P1_U5998, P1_U3412, P1_U3989);
  nand ginst9512 (P1_U5999, P1_REG2_REG_29__SCAN_IN, P1_U3417);
  nand ginst9513 (P1_U6000, P1_U3989, P1_U4708);
  nand ginst9514 (P1_U6001, P1_REG2_REG_30__SCAN_IN, P1_U3417);
  nand ginst9515 (P1_U6002, P1_U3989, P1_U3993);
  nand ginst9516 (P1_U6003, P1_REG2_REG_31__SCAN_IN, P1_U3417);
  nand ginst9517 (P1_U6004, P1_U3989, P1_U3993);
  nand ginst9518 (P1_U6005, P1_DATAO_REG_0__SCAN_IN, P1_U3425);
  nand ginst9519 (P1_U6006, P1_U3077, P1_U3973);
  nand ginst9520 (P1_U6007, P1_DATAO_REG_1__SCAN_IN, P1_U3425);
  nand ginst9521 (P1_U6008, P1_U3078, P1_U3973);
  nand ginst9522 (P1_U6009, P1_DATAO_REG_2__SCAN_IN, P1_U3425);
  nand ginst9523 (P1_U6010, P1_U3068, P1_U3973);
  nand ginst9524 (P1_U6011, P1_DATAO_REG_3__SCAN_IN, P1_U3425);
  nand ginst9525 (P1_U6012, P1_U3064, P1_U3973);
  nand ginst9526 (P1_U6013, P1_DATAO_REG_4__SCAN_IN, P1_U3425);
  nand ginst9527 (P1_U6014, P1_U3060, P1_U3973);
  nand ginst9528 (P1_U6015, P1_DATAO_REG_5__SCAN_IN, P1_U3425);
  nand ginst9529 (P1_U6016, P1_U3067, P1_U3973);
  nand ginst9530 (P1_U6017, P1_DATAO_REG_6__SCAN_IN, P1_U3425);
  nand ginst9531 (P1_U6018, P1_U3071, P1_U3973);
  nand ginst9532 (P1_U6019, P1_DATAO_REG_7__SCAN_IN, P1_U3425);
  nand ginst9533 (P1_U6020, P1_U3070, P1_U3973);
  nand ginst9534 (P1_U6021, P1_DATAO_REG_8__SCAN_IN, P1_U3425);
  nand ginst9535 (P1_U6022, P1_U3084, P1_U3973);
  nand ginst9536 (P1_U6023, P1_DATAO_REG_9__SCAN_IN, P1_U3425);
  nand ginst9537 (P1_U6024, P1_U3083, P1_U3973);
  nand ginst9538 (P1_U6025, P1_DATAO_REG_10__SCAN_IN, P1_U3425);
  nand ginst9539 (P1_U6026, P1_U3062, P1_U3973);
  nand ginst9540 (P1_U6027, P1_DATAO_REG_11__SCAN_IN, P1_U3425);
  nand ginst9541 (P1_U6028, P1_U3063, P1_U3973);
  nand ginst9542 (P1_U6029, P1_DATAO_REG_12__SCAN_IN, P1_U3425);
  nand ginst9543 (P1_U6030, P1_U3072, P1_U3973);
  nand ginst9544 (P1_U6031, P1_DATAO_REG_13__SCAN_IN, P1_U3425);
  nand ginst9545 (P1_U6032, P1_U3080, P1_U3973);
  nand ginst9546 (P1_U6033, P1_DATAO_REG_14__SCAN_IN, P1_U3425);
  nand ginst9547 (P1_U6034, P1_U3079, P1_U3973);
  nand ginst9548 (P1_U6035, P1_DATAO_REG_15__SCAN_IN, P1_U3425);
  nand ginst9549 (P1_U6036, P1_U3074, P1_U3973);
  nand ginst9550 (P1_U6037, P1_DATAO_REG_16__SCAN_IN, P1_U3425);
  nand ginst9551 (P1_U6038, P1_U3073, P1_U3973);
  nand ginst9552 (P1_U6039, P1_DATAO_REG_17__SCAN_IN, P1_U3425);
  nand ginst9553 (P1_U6040, P1_U3069, P1_U3973);
  nand ginst9554 (P1_U6041, P1_DATAO_REG_18__SCAN_IN, P1_U3425);
  nand ginst9555 (P1_U6042, P1_U3082, P1_U3973);
  nand ginst9556 (P1_U6043, P1_DATAO_REG_19__SCAN_IN, P1_U3425);
  nand ginst9557 (P1_U6044, P1_U3081, P1_U3973);
  nand ginst9558 (P1_U6045, P1_DATAO_REG_20__SCAN_IN, P1_U3425);
  nand ginst9559 (P1_U6046, P1_U3076, P1_U3973);
  nand ginst9560 (P1_U6047, P1_DATAO_REG_21__SCAN_IN, P1_U3425);
  nand ginst9561 (P1_U6048, P1_U3075, P1_U3973);
  nand ginst9562 (P1_U6049, P1_DATAO_REG_22__SCAN_IN, P1_U3425);
  nand ginst9563 (P1_U6050, P1_U3061, P1_U3973);
  nand ginst9564 (P1_U6051, P1_DATAO_REG_23__SCAN_IN, P1_U3425);
  nand ginst9565 (P1_U6052, P1_U3066, P1_U3973);
  nand ginst9566 (P1_U6053, P1_DATAO_REG_24__SCAN_IN, P1_U3425);
  nand ginst9567 (P1_U6054, P1_U3065, P1_U3973);
  nand ginst9568 (P1_U6055, P1_DATAO_REG_25__SCAN_IN, P1_U3425);
  nand ginst9569 (P1_U6056, P1_U3058, P1_U3973);
  nand ginst9570 (P1_U6057, P1_DATAO_REG_26__SCAN_IN, P1_U3425);
  nand ginst9571 (P1_U6058, P1_U3057, P1_U3973);
  nand ginst9572 (P1_U6059, P1_DATAO_REG_27__SCAN_IN, P1_U3425);
  nand ginst9573 (P1_U6060, P1_U3053, P1_U3973);
  nand ginst9574 (P1_U6061, P1_DATAO_REG_28__SCAN_IN, P1_U3425);
  nand ginst9575 (P1_U6062, P1_U3054, P1_U3973);
  nand ginst9576 (P1_U6063, P1_DATAO_REG_29__SCAN_IN, P1_U3425);
  nand ginst9577 (P1_U6064, P1_U3055, P1_U3973);
  nand ginst9578 (P1_U6065, P1_DATAO_REG_30__SCAN_IN, P1_U3425);
  nand ginst9579 (P1_U6066, P1_U3059, P1_U3973);
  nand ginst9580 (P1_U6067, P1_DATAO_REG_31__SCAN_IN, P1_U3425);
  nand ginst9581 (P1_U6068, P1_U3056, P1_U3973);
  nand ginst9582 (P1_U6069, P1_U3048, P1_U3438, P1_U3948);
  nand ginst9583 (P1_U6070, P1_R1375_U14, P1_U3954, P1_U5690);
  nand ginst9584 (P1_U6071, P1_U3438, P1_U3447, P1_U3949, P1_U5684);
  nand ginst9585 (P1_U6072, P1_R1360_U14, P1_U3955, P1_U3959);
  nand ginst9586 (P1_U6073, P1_U3055, P1_U3985);
  nand ginst9587 (P1_U6074, P1_U3413, P1_U4678);
  nand ginst9588 (P1_U6075, P1_U6073, P1_U6074);
  nand ginst9589 (P1_U6076, P1_U3054, P1_U3974);
  nand ginst9590 (P1_U6077, P1_U3411, P1_U4659);
  nand ginst9591 (P1_U6078, P1_U6076, P1_U6077);
  nand ginst9592 (P1_U6079, P1_U3053, P1_U3975);
  nand ginst9593 (P1_U6080, P1_U3409, P1_U4640);
  nand ginst9594 (P1_U6081, P1_U6079, P1_U6080);
  nand ginst9595 (P1_U6082, P1_U3065, P1_U3978);
  nand ginst9596 (P1_U6083, P1_U3403, P1_U4583);
  nand ginst9597 (P1_U6084, P1_U6082, P1_U6083);
  nand ginst9598 (P1_U6085, P1_U3066, P1_U3979);
  nand ginst9599 (P1_U6086, P1_U3401, P1_U4564);
  nand ginst9600 (P1_U6087, P1_U6085, P1_U6086);
  nand ginst9601 (P1_U6088, P1_U3075, P1_U3981);
  nand ginst9602 (P1_U6089, P1_U3397, P1_U4526);
  nand ginst9603 (P1_U6090, P1_U6088, P1_U6089);
  nand ginst9604 (P1_U6091, P1_U3061, P1_U3980);
  nand ginst9605 (P1_U6092, P1_U3399, P1_U4545);
  nand ginst9606 (P1_U6093, P1_U6091, P1_U6092);
  nand ginst9607 (P1_U6094, P1_U3058, P1_U3977);
  nand ginst9608 (P1_U6095, P1_U3405, P1_U4602);
  nand ginst9609 (P1_U6096, P1_U6094, P1_U6095);
  nand ginst9610 (P1_U6097, P1_U3057, P1_U3976);
  nand ginst9611 (P1_U6098, P1_U3407, P1_U4621);
  nand ginst9612 (P1_U6099, P1_U6097, P1_U6098);
  nand ginst9613 (P1_U6100, P1_U3059, P1_U3984);
  nand ginst9614 (P1_U6101, P1_U3414, P1_U4696);
  nand ginst9615 (P1_U6102, P1_U6100, P1_U6101);
  nand ginst9616 (P1_U6103, P1_U3056, P1_U3983);
  nand ginst9617 (P1_U6104, P1_U3415, P1_U4716);
  nand ginst9618 (P1_U6105, P1_U6103, P1_U6104);
  nand ginst9619 (P1_U6106, P1_U4450, P1_U5838);
  nand ginst9620 (P1_U6107, P1_U3069, P1_U3503);
  nand ginst9621 (P1_U6108, P1_U6106, P1_U6107);
  nand ginst9622 (P1_U6109, P1_U4279, P1_U5775);
  nand ginst9623 (P1_U6110, P1_U3084, P1_U3476);
  nand ginst9624 (P1_U6111, P1_U6109, P1_U6110);
  nand ginst9625 (P1_U6112, P1_U4298, P1_U5782);
  nand ginst9626 (P1_U6113, P1_U3083, P1_U3479);
  nand ginst9627 (P1_U6114, P1_U6112, P1_U6113);
  nand ginst9628 (P1_U6115, P1_U4374, P1_U5810);
  nand ginst9629 (P1_U6116, P1_U3080, P1_U3491);
  nand ginst9630 (P1_U6117, P1_U6115, P1_U6116);
  nand ginst9631 (P1_U6118, P1_U4393, P1_U5817);
  nand ginst9632 (P1_U6119, P1_U3079, P1_U3494);
  nand ginst9633 (P1_U6120, P1_U6118, P1_U6119);
  nand ginst9634 (P1_U6121, P1_U4165, P1_U5705);
  nand ginst9635 (P1_U6122, P1_U3077, P1_U3450);
  nand ginst9636 (P1_U6123, P1_U6121, P1_U6122);
  nand ginst9637 (P1_U6124, P1_U4141, P1_U5726);
  nand ginst9638 (P1_U6125, P1_U3078, P1_U3455);
  nand ginst9639 (P1_U6126, P1_U6124, P1_U6125);
  nand ginst9640 (P1_U6127, P1_U4412, P1_U5824);
  nand ginst9641 (P1_U6128, P1_U3074, P1_U3497);
  nand ginst9642 (P1_U6129, P1_U6127, P1_U6128);
  nand ginst9643 (P1_U6130, P1_U4431, P1_U5831);
  nand ginst9644 (P1_U6131, P1_U3073, P1_U3500);
  nand ginst9645 (P1_U6132, P1_U6130, P1_U6131);
  nand ginst9646 (P1_U6133, P1_U4241, P1_U5761);
  nand ginst9647 (P1_U6134, P1_U3071, P1_U3470);
  nand ginst9648 (P1_U6135, P1_U6133, P1_U6134);
  nand ginst9649 (P1_U6136, P1_U4260, P1_U5768);
  nand ginst9650 (P1_U6137, P1_U3070, P1_U3473);
  nand ginst9651 (P1_U6138, P1_U6136, P1_U6137);
  nand ginst9652 (P1_U6139, P1_U4355, P1_U5803);
  nand ginst9653 (P1_U6140, P1_U3072, P1_U3488);
  nand ginst9654 (P1_U6141, P1_U6139, P1_U6140);
  nand ginst9655 (P1_U6142, P1_U4160, P1_U5733);
  nand ginst9656 (P1_U6143, P1_U3068, P1_U3458);
  nand ginst9657 (P1_U6144, P1_U6142, P1_U6143);
  nand ginst9658 (P1_U6145, P1_U4184, P1_U5740);
  nand ginst9659 (P1_U6146, P1_U3064, P1_U3461);
  nand ginst9660 (P1_U6147, P1_U6145, P1_U6146);
  nand ginst9661 (P1_U6148, P1_U4222, P1_U5754);
  nand ginst9662 (P1_U6149, P1_U3067, P1_U3467);
  nand ginst9663 (P1_U6150, P1_U6148, P1_U6149);
  nand ginst9664 (P1_U6151, P1_U4469, P1_U5845);
  nand ginst9665 (P1_U6152, P1_U3082, P1_U3506);
  nand ginst9666 (P1_U6153, P1_U6151, P1_U6152);
  nand ginst9667 (P1_U6154, P1_U4488, P1_U5850);
  nand ginst9668 (P1_U6155, P1_U3081, P1_U3508);
  nand ginst9669 (P1_U6156, P1_U6154, P1_U6155);
  nand ginst9670 (P1_U6157, P1_U4203, P1_U5747);
  nand ginst9671 (P1_U6158, P1_U3060, P1_U3464);
  nand ginst9672 (P1_U6159, P1_U6157, P1_U6158);
  nand ginst9673 (P1_U6160, P1_U4336, P1_U5796);
  nand ginst9674 (P1_U6161, P1_U3063, P1_U3485);
  nand ginst9675 (P1_U6162, P1_U6160, P1_U6161);
  nand ginst9676 (P1_U6163, P1_U4317, P1_U5789);
  nand ginst9677 (P1_U6164, P1_U3062, P1_U3482);
  nand ginst9678 (P1_U6165, P1_U6163, P1_U6164);
  nand ginst9679 (P1_U6166, P1_U3076, P1_U3982);
  nand ginst9680 (P1_U6167, P1_U3395, P1_U4507);
  nand ginst9681 (P1_U6168, P1_U6166, P1_U6167);
  nand ginst9682 (P1_U6169, P1_U3951, P1_U5663);
  nand ginst9683 (P1_U6170, P1_U3426, P1_U5086);
  nand ginst9684 (P1_U6171, P1_R1352_U6, P1_U3083);
  nand ginst9685 (P1_U6172, P1_U3083, P1_U3952);
  nand ginst9686 (P1_U6173, P1_R1352_U6, P1_U3084);
  nand ginst9687 (P1_U6174, P1_U3084, P1_U3952);
  nand ginst9688 (P1_U6175, P1_R1352_U6, P1_U3070);
  nand ginst9689 (P1_U6176, P1_U3070, P1_U3952);
  nand ginst9690 (P1_U6177, P1_R1352_U6, P1_U3071);
  nand ginst9691 (P1_U6178, P1_U3071, P1_U3952);
  nand ginst9692 (P1_U6179, P1_R1352_U6, P1_U3067);
  nand ginst9693 (P1_U6180, P1_U3067, P1_U3952);
  nand ginst9694 (P1_U6181, P1_R1352_U6, P1_U3060);
  nand ginst9695 (P1_U6182, P1_U3060, P1_U3952);
  nand ginst9696 (P1_U6183, P1_R1352_U6, P1_U3064);
  nand ginst9697 (P1_U6184, P1_U3064, P1_U3952);
  nand ginst9698 (P1_U6185, P1_R1309_U8, P1_R1352_U6);
  nand ginst9699 (P1_U6186, P1_U3056, P1_U3952);
  nand ginst9700 (P1_U6187, P1_R1309_U6, P1_R1352_U6);
  nand ginst9701 (P1_U6188, P1_U3059, P1_U3952);
  nand ginst9702 (P1_U6189, P1_R1352_U6, P1_U3068);
  nand ginst9703 (P1_U6190, P1_U3068, P1_U3952);
  nand ginst9704 (P1_U6191, P1_R1352_U6, P1_U3055);
  nand ginst9705 (P1_U6192, P1_U3055, P1_U3952);
  nand ginst9706 (P1_U6193, P1_R1352_U6, P1_U3054);
  nand ginst9707 (P1_U6194, P1_U3054, P1_U3952);
  nand ginst9708 (P1_U6195, P1_R1352_U6, P1_U3053);
  nand ginst9709 (P1_U6196, P1_U3053, P1_U3952);
  nand ginst9710 (P1_U6197, P1_R1352_U6, P1_U3057);
  nand ginst9711 (P1_U6198, P1_U3057, P1_U3952);
  nand ginst9712 (P1_U6199, P1_R1352_U6, P1_U3058);
  nand ginst9713 (P1_U6200, P1_U3058, P1_U3952);
  nand ginst9714 (P1_U6201, P1_R1352_U6, P1_U3065);
  nand ginst9715 (P1_U6202, P1_U3065, P1_U3952);
  nand ginst9716 (P1_U6203, P1_R1352_U6, P1_U3066);
  nand ginst9717 (P1_U6204, P1_U3066, P1_U3952);
  nand ginst9718 (P1_U6205, P1_R1352_U6, P1_U3061);
  nand ginst9719 (P1_U6206, P1_U3061, P1_U3952);
  nand ginst9720 (P1_U6207, P1_R1352_U6, P1_U3075);
  nand ginst9721 (P1_U6208, P1_U3075, P1_U3952);
  nand ginst9722 (P1_U6209, P1_R1352_U6, P1_U3076);
  nand ginst9723 (P1_U6210, P1_U3076, P1_U3952);
  nand ginst9724 (P1_U6211, P1_R1352_U6, P1_U3078);
  nand ginst9725 (P1_U6212, P1_U3078, P1_U3952);
  nand ginst9726 (P1_U6213, P1_R1352_U6, P1_U3081);
  nand ginst9727 (P1_U6214, P1_U3081, P1_U3952);
  nand ginst9728 (P1_U6215, P1_R1352_U6, P1_U3082);
  nand ginst9729 (P1_U6216, P1_U3082, P1_U3952);
  nand ginst9730 (P1_U6217, P1_R1352_U6, P1_U3069);
  nand ginst9731 (P1_U6218, P1_U3069, P1_U3952);
  nand ginst9732 (P1_U6219, P1_R1352_U6, P1_U3073);
  nand ginst9733 (P1_U6220, P1_U3073, P1_U3952);
  nand ginst9734 (P1_U6221, P1_R1352_U6, P1_U3074);
  nand ginst9735 (P1_U6222, P1_U3074, P1_U3952);
  nand ginst9736 (P1_U6223, P1_R1352_U6, P1_U3079);
  nand ginst9737 (P1_U6224, P1_U3079, P1_U3952);
  nand ginst9738 (P1_U6225, P1_R1352_U6, P1_U3080);
  nand ginst9739 (P1_U6226, P1_U3080, P1_U3952);
  nand ginst9740 (P1_U6227, P1_R1352_U6, P1_U3072);
  nand ginst9741 (P1_U6228, P1_U3072, P1_U3952);
  nand ginst9742 (P1_U6229, P1_R1352_U6, P1_U3063);
  nand ginst9743 (P1_U6230, P1_U3063, P1_U3952);
  nand ginst9744 (P1_U6231, P1_R1352_U6, P1_U3062);
  nand ginst9745 (P1_U6232, P1_U3062, P1_U3952);
  nand ginst9746 (P1_U6233, P1_R1352_U6, P1_U3077);
  nand ginst9747 (P1_U6234, P1_U3077, P1_U3952);
  nand ginst9748 (P1_U6235, P1_U3448, P1_U5364);
  nand ginst9749 (P1_U6236, P1_REG2_REG_0__SCAN_IN, P1_U3015, P1_U5696);
  and ginst9750 (P2_R1054_U10, P2_R1054_U100, P2_R1054_U174);
  nand ginst9751 (P2_R1054_U100, P2_R1054_U56, P2_U3433);
  nand ginst9752 (P2_R1054_U101, P2_R1054_U24, P2_U3394);
  nand ginst9753 (P2_R1054_U102, P2_R1054_U31, P2_U3403);
  nand ginst9754 (P2_R1054_U103, P2_R1054_U35, P2_U3409);
  not ginst9755 (P2_R1054_U104, P2_R1054_U58);
  not ginst9756 (P2_R1054_U105, P2_R1054_U33);
  not ginst9757 (P2_R1054_U106, P2_R1054_U47);
  not ginst9758 (P2_R1054_U107, P2_R1054_U21);
  nand ginst9759 (P2_R1054_U108, P2_R1054_U107, P2_R1054_U22);
  nand ginst9760 (P2_R1054_U109, P2_R1054_U108, P2_R1054_U88);
  and ginst9761 (P2_R1054_U11, P2_R1054_U175, P2_R1054_U176);
  nand ginst9762 (P2_R1054_U110, P2_R1054_U21, P2_U3573);
  not ginst9763 (P2_R1054_U111, P2_R1054_U42);
  nand ginst9764 (P2_R1054_U112, P2_R1054_U26, P2_U3397);
  nand ginst9765 (P2_R1054_U113, P2_R1054_U101, P2_R1054_U112, P2_R1054_U42);
  nand ginst9766 (P2_R1054_U114, P2_R1054_U25, P2_R1054_U26);
  nand ginst9767 (P2_R1054_U115, P2_R1054_U114, P2_R1054_U23);
  nand ginst9768 (P2_R1054_U116, P2_R1054_U97, P2_U3561);
  not ginst9769 (P2_R1054_U117, P2_R1054_U87);
  nand ginst9770 (P2_R1054_U118, P2_R1054_U30, P2_U3406);
  nand ginst9771 (P2_R1054_U119, P2_R1054_U27, P2_U3558);
  nand ginst9772 (P2_R1054_U12, P2_R1054_U207, P2_R1054_U210);
  nand ginst9773 (P2_R1054_U120, P2_R1054_U28, P2_U3559);
  nand ginst9774 (P2_R1054_U121, P2_R1054_U105, P2_R1054_U6);
  nand ginst9775 (P2_R1054_U122, P2_R1054_U121, P2_R1054_U7);
  nand ginst9776 (P2_R1054_U123, P2_R1054_U32, P2_U3400);
  nand ginst9777 (P2_R1054_U124, P2_R1054_U30, P2_U3406);
  nand ginst9778 (P2_R1054_U125, P2_R1054_U123, P2_R1054_U6, P2_R1054_U87);
  nand ginst9779 (P2_R1054_U126, P2_R1054_U122, P2_R1054_U124);
  not ginst9780 (P2_R1054_U127, P2_R1054_U40);
  nand ginst9781 (P2_R1054_U128, P2_R1054_U37, P2_U3412);
  nand ginst9782 (P2_R1054_U129, P2_R1054_U103, P2_R1054_U128, P2_R1054_U40);
  nand ginst9783 (P2_R1054_U13, P2_R1054_U196, P2_R1054_U199);
  nand ginst9784 (P2_R1054_U130, P2_R1054_U36, P2_R1054_U37);
  nand ginst9785 (P2_R1054_U131, P2_R1054_U130, P2_R1054_U34);
  nand ginst9786 (P2_R1054_U132, P2_R1054_U98, P2_U3556);
  not ginst9787 (P2_R1054_U133, P2_R1054_U86);
  nand ginst9788 (P2_R1054_U134, P2_R1054_U39, P2_U3415);
  nand ginst9789 (P2_R1054_U135, P2_R1054_U134, P2_R1054_U47);
  nand ginst9790 (P2_R1054_U136, P2_R1054_U127, P2_R1054_U36);
  nand ginst9791 (P2_R1054_U137, P2_R1054_U103, P2_R1054_U136, P2_R1054_U222);
  nand ginst9792 (P2_R1054_U138, P2_R1054_U103, P2_R1054_U40);
  nand ginst9793 (P2_R1054_U139, P2_R1054_U138, P2_R1054_U218, P2_R1054_U219, P2_R1054_U36);
  nand ginst9794 (P2_R1054_U14, P2_R1054_U153, P2_R1054_U155);
  nand ginst9795 (P2_R1054_U140, P2_R1054_U103, P2_R1054_U36);
  nand ginst9796 (P2_R1054_U141, P2_R1054_U123, P2_R1054_U87);
  not ginst9797 (P2_R1054_U142, P2_R1054_U41);
  nand ginst9798 (P2_R1054_U143, P2_R1054_U28, P2_U3559);
  nand ginst9799 (P2_R1054_U144, P2_R1054_U142, P2_R1054_U143);
  nand ginst9800 (P2_R1054_U145, P2_R1054_U102, P2_R1054_U144, P2_R1054_U229);
  nand ginst9801 (P2_R1054_U146, P2_R1054_U102, P2_R1054_U41);
  nand ginst9802 (P2_R1054_U147, P2_R1054_U30, P2_U3406);
  nand ginst9803 (P2_R1054_U148, P2_R1054_U146, P2_R1054_U147, P2_R1054_U7);
  nand ginst9804 (P2_R1054_U149, P2_R1054_U28, P2_U3559);
  nand ginst9805 (P2_R1054_U15, P2_R1054_U145, P2_R1054_U148);
  nand ginst9806 (P2_R1054_U150, P2_R1054_U102, P2_R1054_U149);
  nand ginst9807 (P2_R1054_U151, P2_R1054_U123, P2_R1054_U33);
  nand ginst9808 (P2_R1054_U152, P2_R1054_U111, P2_R1054_U25);
  nand ginst9809 (P2_R1054_U153, P2_R1054_U101, P2_R1054_U152, P2_R1054_U242);
  nand ginst9810 (P2_R1054_U154, P2_R1054_U101, P2_R1054_U42);
  nand ginst9811 (P2_R1054_U155, P2_R1054_U154, P2_R1054_U238, P2_R1054_U239, P2_R1054_U25);
  nand ginst9812 (P2_R1054_U156, P2_R1054_U101, P2_R1054_U25);
  nand ginst9813 (P2_R1054_U157, P2_R1054_U45, P2_U3421);
  nand ginst9814 (P2_R1054_U158, P2_R1054_U43, P2_U3571);
  nand ginst9815 (P2_R1054_U159, P2_R1054_U44, P2_U3572);
  nand ginst9816 (P2_R1054_U16, P2_R1054_U137, P2_R1054_U139);
  nand ginst9817 (P2_R1054_U160, P2_R1054_U106, P2_R1054_U8);
  nand ginst9818 (P2_R1054_U161, P2_R1054_U160, P2_R1054_U9);
  nand ginst9819 (P2_R1054_U162, P2_R1054_U45, P2_U3421);
  nand ginst9820 (P2_R1054_U163, P2_R1054_U134, P2_R1054_U8, P2_R1054_U86);
  nand ginst9821 (P2_R1054_U164, P2_R1054_U161, P2_R1054_U162);
  not ginst9822 (P2_R1054_U165, P2_R1054_U96);
  nand ginst9823 (P2_R1054_U166, P2_R1054_U49, P2_U3424);
  nand ginst9824 (P2_R1054_U167, P2_R1054_U166, P2_R1054_U96);
  nand ginst9825 (P2_R1054_U168, P2_R1054_U48, P2_U3570);
  not ginst9826 (P2_R1054_U169, P2_R1054_U95);
  nand ginst9827 (P2_R1054_U17, P2_R1054_U21, P2_R1054_U213);
  nand ginst9828 (P2_R1054_U170, P2_R1054_U51, P2_U3427);
  nand ginst9829 (P2_R1054_U171, P2_R1054_U170, P2_R1054_U95);
  nand ginst9830 (P2_R1054_U172, P2_R1054_U50, P2_U3569);
  not ginst9831 (P2_R1054_U173, P2_R1054_U94);
  nand ginst9832 (P2_R1054_U174, P2_R1054_U55, P2_U3436);
  nand ginst9833 (P2_R1054_U175, P2_R1054_U52, P2_U3566);
  nand ginst9834 (P2_R1054_U176, P2_R1054_U53, P2_U3567);
  nand ginst9835 (P2_R1054_U177, P2_R1054_U10, P2_R1054_U104);
  nand ginst9836 (P2_R1054_U178, P2_R1054_U11, P2_R1054_U177);
  nand ginst9837 (P2_R1054_U179, P2_R1054_U57, P2_U3430);
  not ginst9838 (P2_R1054_U18, P2_U3409);
  nand ginst9839 (P2_R1054_U180, P2_R1054_U55, P2_U3436);
  nand ginst9840 (P2_R1054_U181, P2_R1054_U10, P2_R1054_U179, P2_R1054_U94);
  nand ginst9841 (P2_R1054_U182, P2_R1054_U178, P2_R1054_U180);
  not ginst9842 (P2_R1054_U183, P2_R1054_U93);
  nand ginst9843 (P2_R1054_U184, P2_R1054_U60, P2_U3439);
  nand ginst9844 (P2_R1054_U185, P2_R1054_U184, P2_R1054_U93);
  nand ginst9845 (P2_R1054_U186, P2_R1054_U59, P2_U3565);
  not ginst9846 (P2_R1054_U187, P2_R1054_U61);
  nand ginst9847 (P2_R1054_U188, P2_R1054_U187, P2_R1054_U62);
  nand ginst9848 (P2_R1054_U189, P2_R1054_U188, P2_R1054_U92);
  not ginst9849 (P2_R1054_U19, P2_U3394);
  nand ginst9850 (P2_R1054_U190, P2_R1054_U61, P2_U3564);
  not ginst9851 (P2_R1054_U191, P2_R1054_U91);
  nand ginst9852 (P2_R1054_U192, P2_R1054_U179, P2_R1054_U94);
  not ginst9853 (P2_R1054_U193, P2_R1054_U63);
  nand ginst9854 (P2_R1054_U194, P2_R1054_U53, P2_U3567);
  nand ginst9855 (P2_R1054_U195, P2_R1054_U193, P2_R1054_U194);
  nand ginst9856 (P2_R1054_U196, P2_R1054_U100, P2_R1054_U195, P2_R1054_U269);
  nand ginst9857 (P2_R1054_U197, P2_R1054_U100, P2_R1054_U63);
  nand ginst9858 (P2_R1054_U198, P2_R1054_U55, P2_U3436);
  nand ginst9859 (P2_R1054_U199, P2_R1054_U11, P2_R1054_U197, P2_R1054_U198);
  not ginst9860 (P2_R1054_U20, P2_U3386);
  nand ginst9861 (P2_R1054_U200, P2_R1054_U53, P2_U3567);
  nand ginst9862 (P2_R1054_U201, P2_R1054_U100, P2_R1054_U200);
  nand ginst9863 (P2_R1054_U202, P2_R1054_U179, P2_R1054_U58);
  nand ginst9864 (P2_R1054_U203, P2_R1054_U134, P2_R1054_U86);
  not ginst9865 (P2_R1054_U204, P2_R1054_U64);
  nand ginst9866 (P2_R1054_U205, P2_R1054_U44, P2_U3572);
  nand ginst9867 (P2_R1054_U206, P2_R1054_U204, P2_R1054_U205);
  nand ginst9868 (P2_R1054_U207, P2_R1054_U206, P2_R1054_U290, P2_R1054_U99);
  nand ginst9869 (P2_R1054_U208, P2_R1054_U64, P2_R1054_U99);
  nand ginst9870 (P2_R1054_U209, P2_R1054_U45, P2_U3421);
  nand ginst9871 (P2_R1054_U21, P2_R1054_U65, P2_U3386);
  nand ginst9872 (P2_R1054_U210, P2_R1054_U208, P2_R1054_U209, P2_R1054_U9);
  nand ginst9873 (P2_R1054_U211, P2_R1054_U44, P2_U3572);
  nand ginst9874 (P2_R1054_U212, P2_R1054_U211, P2_R1054_U99);
  nand ginst9875 (P2_R1054_U213, P2_R1054_U20, P2_U3574);
  nand ginst9876 (P2_R1054_U214, P2_R1054_U39, P2_U3415);
  nand ginst9877 (P2_R1054_U215, P2_R1054_U38, P2_U3555);
  nand ginst9878 (P2_R1054_U216, P2_R1054_U135, P2_R1054_U86);
  nand ginst9879 (P2_R1054_U217, P2_R1054_U133, P2_R1054_U214, P2_R1054_U215);
  nand ginst9880 (P2_R1054_U218, P2_R1054_U37, P2_U3412);
  nand ginst9881 (P2_R1054_U219, P2_R1054_U34, P2_U3556);
  not ginst9882 (P2_R1054_U22, P2_U3573);
  nand ginst9883 (P2_R1054_U220, P2_R1054_U37, P2_U3412);
  nand ginst9884 (P2_R1054_U221, P2_R1054_U34, P2_U3556);
  nand ginst9885 (P2_R1054_U222, P2_R1054_U220, P2_R1054_U221);
  nand ginst9886 (P2_R1054_U223, P2_R1054_U35, P2_U3409);
  nand ginst9887 (P2_R1054_U224, P2_R1054_U18, P2_U3557);
  nand ginst9888 (P2_R1054_U225, P2_R1054_U140, P2_R1054_U40);
  nand ginst9889 (P2_R1054_U226, P2_R1054_U127, P2_R1054_U223, P2_R1054_U224);
  nand ginst9890 (P2_R1054_U227, P2_R1054_U30, P2_U3406);
  nand ginst9891 (P2_R1054_U228, P2_R1054_U27, P2_U3558);
  nand ginst9892 (P2_R1054_U229, P2_R1054_U227, P2_R1054_U228);
  not ginst9893 (P2_R1054_U23, P2_U3397);
  nand ginst9894 (P2_R1054_U230, P2_R1054_U31, P2_U3403);
  nand ginst9895 (P2_R1054_U231, P2_R1054_U28, P2_U3559);
  nand ginst9896 (P2_R1054_U232, P2_R1054_U150, P2_R1054_U41);
  nand ginst9897 (P2_R1054_U233, P2_R1054_U142, P2_R1054_U230, P2_R1054_U231);
  nand ginst9898 (P2_R1054_U234, P2_R1054_U32, P2_U3400);
  nand ginst9899 (P2_R1054_U235, P2_R1054_U29, P2_U3560);
  nand ginst9900 (P2_R1054_U236, P2_R1054_U151, P2_R1054_U87);
  nand ginst9901 (P2_R1054_U237, P2_R1054_U117, P2_R1054_U234, P2_R1054_U235);
  nand ginst9902 (P2_R1054_U238, P2_R1054_U26, P2_U3397);
  nand ginst9903 (P2_R1054_U239, P2_R1054_U23, P2_U3561);
  not ginst9904 (P2_R1054_U24, P2_U3562);
  nand ginst9905 (P2_R1054_U240, P2_R1054_U26, P2_U3397);
  nand ginst9906 (P2_R1054_U241, P2_R1054_U23, P2_U3561);
  nand ginst9907 (P2_R1054_U242, P2_R1054_U240, P2_R1054_U241);
  nand ginst9908 (P2_R1054_U243, P2_R1054_U24, P2_U3394);
  nand ginst9909 (P2_R1054_U244, P2_R1054_U19, P2_U3562);
  nand ginst9910 (P2_R1054_U245, P2_R1054_U156, P2_R1054_U42);
  nand ginst9911 (P2_R1054_U246, P2_R1054_U111, P2_R1054_U243, P2_R1054_U244);
  nand ginst9912 (P2_R1054_U247, P2_R1054_U22, P2_U3391);
  nand ginst9913 (P2_R1054_U248, P2_R1054_U88, P2_U3573);
  not ginst9914 (P2_R1054_U249, P2_R1054_U80);
  nand ginst9915 (P2_R1054_U25, P2_R1054_U19, P2_U3562);
  nand ginst9916 (P2_R1054_U250, P2_R1054_U107, P2_R1054_U249);
  nand ginst9917 (P2_R1054_U251, P2_R1054_U21, P2_R1054_U80);
  nand ginst9918 (P2_R1054_U252, P2_R1054_U90, P2_U3379);
  nand ginst9919 (P2_R1054_U253, P2_R1054_U89, P2_U3563);
  not ginst9920 (P2_R1054_U254, P2_R1054_U81);
  nand ginst9921 (P2_R1054_U255, P2_R1054_U191, P2_R1054_U254);
  nand ginst9922 (P2_R1054_U256, P2_R1054_U81, P2_R1054_U91);
  nand ginst9923 (P2_R1054_U257, P2_R1054_U62, P2_U3442);
  nand ginst9924 (P2_R1054_U258, P2_R1054_U92, P2_U3564);
  not ginst9925 (P2_R1054_U259, P2_R1054_U82);
  not ginst9926 (P2_R1054_U26, P2_U3561);
  nand ginst9927 (P2_R1054_U260, P2_R1054_U187, P2_R1054_U259);
  nand ginst9928 (P2_R1054_U261, P2_R1054_U61, P2_R1054_U82);
  nand ginst9929 (P2_R1054_U262, P2_R1054_U60, P2_U3439);
  nand ginst9930 (P2_R1054_U263, P2_R1054_U59, P2_U3565);
  not ginst9931 (P2_R1054_U264, P2_R1054_U83);
  nand ginst9932 (P2_R1054_U265, P2_R1054_U183, P2_R1054_U264);
  nand ginst9933 (P2_R1054_U266, P2_R1054_U83, P2_R1054_U93);
  nand ginst9934 (P2_R1054_U267, P2_R1054_U55, P2_U3436);
  nand ginst9935 (P2_R1054_U268, P2_R1054_U52, P2_U3566);
  nand ginst9936 (P2_R1054_U269, P2_R1054_U267, P2_R1054_U268);
  not ginst9937 (P2_R1054_U27, P2_U3406);
  nand ginst9938 (P2_R1054_U270, P2_R1054_U56, P2_U3433);
  nand ginst9939 (P2_R1054_U271, P2_R1054_U53, P2_U3567);
  nand ginst9940 (P2_R1054_U272, P2_R1054_U201, P2_R1054_U63);
  nand ginst9941 (P2_R1054_U273, P2_R1054_U193, P2_R1054_U270, P2_R1054_U271);
  nand ginst9942 (P2_R1054_U274, P2_R1054_U57, P2_U3430);
  nand ginst9943 (P2_R1054_U275, P2_R1054_U54, P2_U3568);
  nand ginst9944 (P2_R1054_U276, P2_R1054_U202, P2_R1054_U94);
  nand ginst9945 (P2_R1054_U277, P2_R1054_U173, P2_R1054_U274, P2_R1054_U275);
  nand ginst9946 (P2_R1054_U278, P2_R1054_U51, P2_U3427);
  nand ginst9947 (P2_R1054_U279, P2_R1054_U50, P2_U3569);
  not ginst9948 (P2_R1054_U28, P2_U3403);
  not ginst9949 (P2_R1054_U280, P2_R1054_U84);
  nand ginst9950 (P2_R1054_U281, P2_R1054_U169, P2_R1054_U280);
  nand ginst9951 (P2_R1054_U282, P2_R1054_U84, P2_R1054_U95);
  nand ginst9952 (P2_R1054_U283, P2_R1054_U49, P2_U3424);
  nand ginst9953 (P2_R1054_U284, P2_R1054_U48, P2_U3570);
  not ginst9954 (P2_R1054_U285, P2_R1054_U85);
  nand ginst9955 (P2_R1054_U286, P2_R1054_U165, P2_R1054_U285);
  nand ginst9956 (P2_R1054_U287, P2_R1054_U85, P2_R1054_U96);
  nand ginst9957 (P2_R1054_U288, P2_R1054_U45, P2_U3421);
  nand ginst9958 (P2_R1054_U289, P2_R1054_U43, P2_U3571);
  not ginst9959 (P2_R1054_U29, P2_U3400);
  nand ginst9960 (P2_R1054_U290, P2_R1054_U288, P2_R1054_U289);
  nand ginst9961 (P2_R1054_U291, P2_R1054_U46, P2_U3418);
  nand ginst9962 (P2_R1054_U292, P2_R1054_U44, P2_U3572);
  nand ginst9963 (P2_R1054_U293, P2_R1054_U212, P2_R1054_U64);
  nand ginst9964 (P2_R1054_U294, P2_R1054_U204, P2_R1054_U291, P2_R1054_U292);
  not ginst9965 (P2_R1054_U30, P2_U3558);
  not ginst9966 (P2_R1054_U31, P2_U3559);
  not ginst9967 (P2_R1054_U32, P2_U3560);
  nand ginst9968 (P2_R1054_U33, P2_R1054_U29, P2_U3560);
  not ginst9969 (P2_R1054_U34, P2_U3412);
  not ginst9970 (P2_R1054_U35, P2_U3557);
  nand ginst9971 (P2_R1054_U36, P2_R1054_U18, P2_U3557);
  not ginst9972 (P2_R1054_U37, P2_U3556);
  not ginst9973 (P2_R1054_U38, P2_U3415);
  not ginst9974 (P2_R1054_U39, P2_U3555);
  nand ginst9975 (P2_R1054_U40, P2_R1054_U125, P2_R1054_U126);
  nand ginst9976 (P2_R1054_U41, P2_R1054_U141, P2_R1054_U33);
  nand ginst9977 (P2_R1054_U42, P2_R1054_U109, P2_R1054_U110);
  not ginst9978 (P2_R1054_U43, P2_U3421);
  not ginst9979 (P2_R1054_U44, P2_U3418);
  not ginst9980 (P2_R1054_U45, P2_U3571);
  not ginst9981 (P2_R1054_U46, P2_U3572);
  nand ginst9982 (P2_R1054_U47, P2_R1054_U38, P2_U3555);
  not ginst9983 (P2_R1054_U48, P2_U3424);
  not ginst9984 (P2_R1054_U49, P2_U3570);
  not ginst9985 (P2_R1054_U50, P2_U3427);
  not ginst9986 (P2_R1054_U51, P2_U3569);
  not ginst9987 (P2_R1054_U52, P2_U3436);
  not ginst9988 (P2_R1054_U53, P2_U3433);
  not ginst9989 (P2_R1054_U54, P2_U3430);
  not ginst9990 (P2_R1054_U55, P2_U3566);
  not ginst9991 (P2_R1054_U56, P2_U3567);
  not ginst9992 (P2_R1054_U57, P2_U3568);
  nand ginst9993 (P2_R1054_U58, P2_R1054_U54, P2_U3568);
  not ginst9994 (P2_R1054_U59, P2_U3439);
  and ginst9995 (P2_R1054_U6, P2_R1054_U102, P2_R1054_U118);
  not ginst9996 (P2_R1054_U60, P2_U3565);
  nand ginst9997 (P2_R1054_U61, P2_R1054_U185, P2_R1054_U186);
  not ginst9998 (P2_R1054_U62, P2_U3564);
  nand ginst9999 (P2_R1054_U63, P2_R1054_U192, P2_R1054_U58);
  nand ginst10000 (P2_R1054_U64, P2_R1054_U203, P2_R1054_U47);
  not ginst10001 (P2_R1054_U65, P2_U3574);
  nand ginst10002 (P2_R1054_U66, P2_R1054_U250, P2_R1054_U251);
  nand ginst10003 (P2_R1054_U67, P2_R1054_U255, P2_R1054_U256);
  nand ginst10004 (P2_R1054_U68, P2_R1054_U260, P2_R1054_U261);
  nand ginst10005 (P2_R1054_U69, P2_R1054_U265, P2_R1054_U266);
  and ginst10006 (P2_R1054_U7, P2_R1054_U119, P2_R1054_U120);
  nand ginst10007 (P2_R1054_U70, P2_R1054_U281, P2_R1054_U282);
  nand ginst10008 (P2_R1054_U71, P2_R1054_U286, P2_R1054_U287);
  nand ginst10009 (P2_R1054_U72, P2_R1054_U216, P2_R1054_U217);
  nand ginst10010 (P2_R1054_U73, P2_R1054_U225, P2_R1054_U226);
  nand ginst10011 (P2_R1054_U74, P2_R1054_U232, P2_R1054_U233);
  nand ginst10012 (P2_R1054_U75, P2_R1054_U236, P2_R1054_U237);
  nand ginst10013 (P2_R1054_U76, P2_R1054_U245, P2_R1054_U246);
  nand ginst10014 (P2_R1054_U77, P2_R1054_U272, P2_R1054_U273);
  nand ginst10015 (P2_R1054_U78, P2_R1054_U276, P2_R1054_U277);
  nand ginst10016 (P2_R1054_U79, P2_R1054_U293, P2_R1054_U294);
  and ginst10017 (P2_R1054_U8, P2_R1054_U157, P2_R1054_U99);
  nand ginst10018 (P2_R1054_U80, P2_R1054_U247, P2_R1054_U248);
  nand ginst10019 (P2_R1054_U81, P2_R1054_U252, P2_R1054_U253);
  nand ginst10020 (P2_R1054_U82, P2_R1054_U257, P2_R1054_U258);
  nand ginst10021 (P2_R1054_U83, P2_R1054_U262, P2_R1054_U263);
  nand ginst10022 (P2_R1054_U84, P2_R1054_U278, P2_R1054_U279);
  nand ginst10023 (P2_R1054_U85, P2_R1054_U283, P2_R1054_U284);
  nand ginst10024 (P2_R1054_U86, P2_R1054_U129, P2_R1054_U131, P2_R1054_U132);
  nand ginst10025 (P2_R1054_U87, P2_R1054_U113, P2_R1054_U115, P2_R1054_U116);
  not ginst10026 (P2_R1054_U88, P2_U3391);
  not ginst10027 (P2_R1054_U89, P2_U3379);
  and ginst10028 (P2_R1054_U9, P2_R1054_U158, P2_R1054_U159);
  not ginst10029 (P2_R1054_U90, P2_U3563);
  nand ginst10030 (P2_R1054_U91, P2_R1054_U189, P2_R1054_U190);
  not ginst10031 (P2_R1054_U92, P2_U3442);
  nand ginst10032 (P2_R1054_U93, P2_R1054_U181, P2_R1054_U182);
  nand ginst10033 (P2_R1054_U94, P2_R1054_U171, P2_R1054_U172);
  nand ginst10034 (P2_R1054_U95, P2_R1054_U167, P2_R1054_U168);
  nand ginst10035 (P2_R1054_U96, P2_R1054_U163, P2_R1054_U164);
  not ginst10036 (P2_R1054_U97, P2_R1054_U25);
  not ginst10037 (P2_R1054_U98, P2_R1054_U36);
  nand ginst10038 (P2_R1054_U99, P2_R1054_U46, P2_U3418);
  and ginst10039 (P2_R1077_U10, P2_R1077_U348, P2_R1077_U351);
  nand ginst10040 (P2_R1077_U100, P2_R1077_U398, P2_R1077_U399);
  nand ginst10041 (P2_R1077_U101, P2_R1077_U407, P2_R1077_U408);
  nand ginst10042 (P2_R1077_U102, P2_R1077_U414, P2_R1077_U415);
  nand ginst10043 (P2_R1077_U103, P2_R1077_U421, P2_R1077_U422);
  nand ginst10044 (P2_R1077_U104, P2_R1077_U428, P2_R1077_U429);
  nand ginst10045 (P2_R1077_U105, P2_R1077_U433, P2_R1077_U434);
  nand ginst10046 (P2_R1077_U106, P2_R1077_U440, P2_R1077_U441);
  nand ginst10047 (P2_R1077_U107, P2_R1077_U447, P2_R1077_U448);
  nand ginst10048 (P2_R1077_U108, P2_R1077_U461, P2_R1077_U462);
  nand ginst10049 (P2_R1077_U109, P2_R1077_U466, P2_R1077_U467);
  and ginst10050 (P2_R1077_U11, P2_R1077_U341, P2_R1077_U344);
  nand ginst10051 (P2_R1077_U110, P2_R1077_U473, P2_R1077_U474);
  nand ginst10052 (P2_R1077_U111, P2_R1077_U480, P2_R1077_U481);
  nand ginst10053 (P2_R1077_U112, P2_R1077_U487, P2_R1077_U488);
  nand ginst10054 (P2_R1077_U113, P2_R1077_U494, P2_R1077_U495);
  nand ginst10055 (P2_R1077_U114, P2_R1077_U499, P2_R1077_U500);
  and ginst10056 (P2_R1077_U115, P2_R1077_U187, P2_R1077_U189);
  and ginst10057 (P2_R1077_U116, P2_R1077_U180, P2_R1077_U4);
  and ginst10058 (P2_R1077_U117, P2_R1077_U192, P2_R1077_U194);
  and ginst10059 (P2_R1077_U118, P2_R1077_U200, P2_R1077_U201);
  and ginst10060 (P2_R1077_U119, P2_R1077_U22, P2_R1077_U381, P2_R1077_U382);
  and ginst10061 (P2_R1077_U12, P2_R1077_U332, P2_R1077_U335);
  and ginst10062 (P2_R1077_U120, P2_R1077_U212, P2_R1077_U5);
  and ginst10063 (P2_R1077_U121, P2_R1077_U180, P2_R1077_U181);
  and ginst10064 (P2_R1077_U122, P2_R1077_U218, P2_R1077_U220);
  and ginst10065 (P2_R1077_U123, P2_R1077_U34, P2_R1077_U388, P2_R1077_U389);
  and ginst10066 (P2_R1077_U124, P2_R1077_U226, P2_R1077_U4);
  and ginst10067 (P2_R1077_U125, P2_R1077_U181, P2_R1077_U234);
  and ginst10068 (P2_R1077_U126, P2_R1077_U204, P2_R1077_U6);
  and ginst10069 (P2_R1077_U127, P2_R1077_U239, P2_R1077_U243);
  and ginst10070 (P2_R1077_U128, P2_R1077_U250, P2_R1077_U7);
  and ginst10071 (P2_R1077_U129, P2_R1077_U248, P2_R1077_U253);
  and ginst10072 (P2_R1077_U13, P2_R1077_U323, P2_R1077_U326);
  and ginst10073 (P2_R1077_U130, P2_R1077_U267, P2_R1077_U268);
  and ginst10074 (P2_R1077_U131, P2_R1077_U282, P2_R1077_U9);
  and ginst10075 (P2_R1077_U132, P2_R1077_U280, P2_R1077_U285);
  and ginst10076 (P2_R1077_U133, P2_R1077_U298, P2_R1077_U301);
  and ginst10077 (P2_R1077_U134, P2_R1077_U302, P2_R1077_U368);
  and ginst10078 (P2_R1077_U135, P2_R1077_U160, P2_R1077_U278);
  and ginst10079 (P2_R1077_U136, P2_R1077_U454, P2_R1077_U455, P2_R1077_U80);
  and ginst10080 (P2_R1077_U137, P2_R1077_U325, P2_R1077_U9);
  and ginst10081 (P2_R1077_U138, P2_R1077_U468, P2_R1077_U469, P2_R1077_U59);
  and ginst10082 (P2_R1077_U139, P2_R1077_U334, P2_R1077_U8);
  and ginst10083 (P2_R1077_U14, P2_R1077_U318, P2_R1077_U320);
  and ginst10084 (P2_R1077_U140, P2_R1077_U172, P2_R1077_U489, P2_R1077_U490);
  and ginst10085 (P2_R1077_U141, P2_R1077_U343, P2_R1077_U7);
  and ginst10086 (P2_R1077_U142, P2_R1077_U171, P2_R1077_U501, P2_R1077_U502);
  and ginst10087 (P2_R1077_U143, P2_R1077_U350, P2_R1077_U6);
  nand ginst10088 (P2_R1077_U144, P2_R1077_U118, P2_R1077_U202);
  nand ginst10089 (P2_R1077_U145, P2_R1077_U217, P2_R1077_U229);
  not ginst10090 (P2_R1077_U146, P2_U3054);
  not ginst10091 (P2_R1077_U147, P2_U3904);
  and ginst10092 (P2_R1077_U148, P2_R1077_U402, P2_R1077_U403);
  nand ginst10093 (P2_R1077_U149, P2_R1077_U169, P2_R1077_U304, P2_R1077_U364);
  and ginst10094 (P2_R1077_U15, P2_R1077_U310, P2_R1077_U313);
  and ginst10095 (P2_R1077_U150, P2_R1077_U409, P2_R1077_U410);
  nand ginst10096 (P2_R1077_U151, P2_R1077_U134, P2_R1077_U369, P2_R1077_U370);
  and ginst10097 (P2_R1077_U152, P2_R1077_U416, P2_R1077_U417);
  nand ginst10098 (P2_R1077_U153, P2_R1077_U299, P2_R1077_U365, P2_R1077_U86);
  and ginst10099 (P2_R1077_U154, P2_R1077_U423, P2_R1077_U424);
  nand ginst10100 (P2_R1077_U155, P2_R1077_U292, P2_R1077_U293);
  and ginst10101 (P2_R1077_U156, P2_R1077_U435, P2_R1077_U436);
  nand ginst10102 (P2_R1077_U157, P2_R1077_U288, P2_R1077_U289);
  and ginst10103 (P2_R1077_U158, P2_R1077_U442, P2_R1077_U443);
  nand ginst10104 (P2_R1077_U159, P2_R1077_U132, P2_R1077_U284);
  and ginst10105 (P2_R1077_U16, P2_R1077_U232, P2_R1077_U235);
  and ginst10106 (P2_R1077_U160, P2_R1077_U449, P2_R1077_U450);
  nand ginst10107 (P2_R1077_U161, P2_R1077_U327, P2_R1077_U43);
  nand ginst10108 (P2_R1077_U162, P2_R1077_U130, P2_R1077_U269);
  and ginst10109 (P2_R1077_U163, P2_R1077_U475, P2_R1077_U476);
  nand ginst10110 (P2_R1077_U164, P2_R1077_U256, P2_R1077_U257);
  and ginst10111 (P2_R1077_U165, P2_R1077_U482, P2_R1077_U483);
  nand ginst10112 (P2_R1077_U166, P2_R1077_U129, P2_R1077_U252);
  nand ginst10113 (P2_R1077_U167, P2_R1077_U127, P2_R1077_U242);
  nand ginst10114 (P2_R1077_U168, P2_R1077_U366, P2_R1077_U367);
  nand ginst10115 (P2_R1077_U169, P2_R1077_U151, P2_U3053);
  and ginst10116 (P2_R1077_U17, P2_R1077_U224, P2_R1077_U227);
  not ginst10117 (P2_R1077_U170, P2_R1077_U34);
  nand ginst10118 (P2_R1077_U171, P2_U3082, P2_U3416);
  nand ginst10119 (P2_R1077_U172, P2_U3071, P2_U3425);
  nand ginst10120 (P2_R1077_U173, P2_U3057, P2_U3898);
  not ginst10121 (P2_R1077_U174, P2_R1077_U68);
  not ginst10122 (P2_R1077_U175, P2_R1077_U77);
  nand ginst10123 (P2_R1077_U176, P2_U3064, P2_U3899);
  not ginst10124 (P2_R1077_U177, P2_R1077_U65);
  or ginst10125 (P2_R1077_U178, P2_U3066, P2_U3404);
  or ginst10126 (P2_R1077_U179, P2_U3059, P2_U3401);
  and ginst10127 (P2_R1077_U18, P2_R1077_U210, P2_R1077_U213);
  or ginst10128 (P2_R1077_U180, P2_U3063, P2_U3398);
  or ginst10129 (P2_R1077_U181, P2_U3067, P2_U3395);
  not ginst10130 (P2_R1077_U182, P2_R1077_U31);
  or ginst10131 (P2_R1077_U183, P2_U3077, P2_U3392);
  not ginst10132 (P2_R1077_U184, P2_R1077_U42);
  not ginst10133 (P2_R1077_U185, P2_R1077_U43);
  nand ginst10134 (P2_R1077_U186, P2_R1077_U42, P2_R1077_U43);
  nand ginst10135 (P2_R1077_U187, P2_U3067, P2_U3395);
  nand ginst10136 (P2_R1077_U188, P2_R1077_U181, P2_R1077_U186);
  nand ginst10137 (P2_R1077_U189, P2_U3063, P2_U3398);
  not ginst10138 (P2_R1077_U19, P2_U3407);
  nand ginst10139 (P2_R1077_U190, P2_R1077_U115, P2_R1077_U188);
  nand ginst10140 (P2_R1077_U191, P2_R1077_U34, P2_R1077_U35);
  nand ginst10141 (P2_R1077_U192, P2_R1077_U191, P2_U3066);
  nand ginst10142 (P2_R1077_U193, P2_R1077_U116, P2_R1077_U190);
  nand ginst10143 (P2_R1077_U194, P2_R1077_U170, P2_U3404);
  not ginst10144 (P2_R1077_U195, P2_R1077_U41);
  or ginst10145 (P2_R1077_U196, P2_U3069, P2_U3410);
  or ginst10146 (P2_R1077_U197, P2_U3070, P2_U3407);
  not ginst10147 (P2_R1077_U198, P2_R1077_U22);
  nand ginst10148 (P2_R1077_U199, P2_R1077_U22, P2_R1077_U23);
  not ginst10149 (P2_R1077_U20, P2_U3070);
  nand ginst10150 (P2_R1077_U200, P2_R1077_U199, P2_U3069);
  nand ginst10151 (P2_R1077_U201, P2_R1077_U198, P2_U3410);
  nand ginst10152 (P2_R1077_U202, P2_R1077_U41, P2_R1077_U5);
  not ginst10153 (P2_R1077_U203, P2_R1077_U144);
  or ginst10154 (P2_R1077_U204, P2_U3083, P2_U3413);
  nand ginst10155 (P2_R1077_U205, P2_R1077_U144, P2_R1077_U204);
  not ginst10156 (P2_R1077_U206, P2_R1077_U40);
  or ginst10157 (P2_R1077_U207, P2_U3082, P2_U3416);
  or ginst10158 (P2_R1077_U208, P2_U3070, P2_U3407);
  nand ginst10159 (P2_R1077_U209, P2_R1077_U208, P2_R1077_U41);
  not ginst10160 (P2_R1077_U21, P2_U3069);
  nand ginst10161 (P2_R1077_U210, P2_R1077_U119, P2_R1077_U209);
  nand ginst10162 (P2_R1077_U211, P2_R1077_U195, P2_R1077_U22);
  nand ginst10163 (P2_R1077_U212, P2_U3069, P2_U3410);
  nand ginst10164 (P2_R1077_U213, P2_R1077_U120, P2_R1077_U211);
  or ginst10165 (P2_R1077_U214, P2_U3070, P2_U3407);
  nand ginst10166 (P2_R1077_U215, P2_R1077_U181, P2_R1077_U185);
  nand ginst10167 (P2_R1077_U216, P2_U3067, P2_U3395);
  not ginst10168 (P2_R1077_U217, P2_R1077_U45);
  nand ginst10169 (P2_R1077_U218, P2_R1077_U121, P2_R1077_U184);
  nand ginst10170 (P2_R1077_U219, P2_R1077_U180, P2_R1077_U45);
  nand ginst10171 (P2_R1077_U22, P2_U3070, P2_U3407);
  nand ginst10172 (P2_R1077_U220, P2_U3063, P2_U3398);
  not ginst10173 (P2_R1077_U221, P2_R1077_U44);
  or ginst10174 (P2_R1077_U222, P2_U3059, P2_U3401);
  nand ginst10175 (P2_R1077_U223, P2_R1077_U222, P2_R1077_U44);
  nand ginst10176 (P2_R1077_U224, P2_R1077_U123, P2_R1077_U223);
  nand ginst10177 (P2_R1077_U225, P2_R1077_U221, P2_R1077_U34);
  nand ginst10178 (P2_R1077_U226, P2_U3066, P2_U3404);
  nand ginst10179 (P2_R1077_U227, P2_R1077_U124, P2_R1077_U225);
  or ginst10180 (P2_R1077_U228, P2_U3059, P2_U3401);
  nand ginst10181 (P2_R1077_U229, P2_R1077_U181, P2_R1077_U184);
  not ginst10182 (P2_R1077_U23, P2_U3410);
  not ginst10183 (P2_R1077_U230, P2_R1077_U145);
  nand ginst10184 (P2_R1077_U231, P2_U3063, P2_U3398);
  nand ginst10185 (P2_R1077_U232, P2_R1077_U400, P2_R1077_U401, P2_R1077_U42, P2_R1077_U43);
  nand ginst10186 (P2_R1077_U233, P2_R1077_U42, P2_R1077_U43);
  nand ginst10187 (P2_R1077_U234, P2_U3067, P2_U3395);
  nand ginst10188 (P2_R1077_U235, P2_R1077_U125, P2_R1077_U233);
  or ginst10189 (P2_R1077_U236, P2_U3082, P2_U3416);
  or ginst10190 (P2_R1077_U237, P2_U3061, P2_U3419);
  nand ginst10191 (P2_R1077_U238, P2_R1077_U177, P2_R1077_U6);
  nand ginst10192 (P2_R1077_U239, P2_U3061, P2_U3419);
  not ginst10193 (P2_R1077_U24, P2_U3401);
  nand ginst10194 (P2_R1077_U240, P2_R1077_U171, P2_R1077_U238);
  or ginst10195 (P2_R1077_U241, P2_U3061, P2_U3419);
  nand ginst10196 (P2_R1077_U242, P2_R1077_U126, P2_R1077_U144);
  nand ginst10197 (P2_R1077_U243, P2_R1077_U240, P2_R1077_U241);
  not ginst10198 (P2_R1077_U244, P2_R1077_U167);
  or ginst10199 (P2_R1077_U245, P2_U3079, P2_U3428);
  or ginst10200 (P2_R1077_U246, P2_U3071, P2_U3425);
  nand ginst10201 (P2_R1077_U247, P2_R1077_U174, P2_R1077_U7);
  nand ginst10202 (P2_R1077_U248, P2_U3079, P2_U3428);
  nand ginst10203 (P2_R1077_U249, P2_R1077_U172, P2_R1077_U247);
  not ginst10204 (P2_R1077_U25, P2_U3059);
  or ginst10205 (P2_R1077_U250, P2_U3062, P2_U3422);
  or ginst10206 (P2_R1077_U251, P2_U3079, P2_U3428);
  nand ginst10207 (P2_R1077_U252, P2_R1077_U128, P2_R1077_U167);
  nand ginst10208 (P2_R1077_U253, P2_R1077_U249, P2_R1077_U251);
  not ginst10209 (P2_R1077_U254, P2_R1077_U166);
  or ginst10210 (P2_R1077_U255, P2_U3078, P2_U3431);
  nand ginst10211 (P2_R1077_U256, P2_R1077_U166, P2_R1077_U255);
  nand ginst10212 (P2_R1077_U257, P2_U3078, P2_U3431);
  not ginst10213 (P2_R1077_U258, P2_R1077_U164);
  or ginst10214 (P2_R1077_U259, P2_U3073, P2_U3434);
  not ginst10215 (P2_R1077_U26, P2_U3066);
  nand ginst10216 (P2_R1077_U260, P2_R1077_U164, P2_R1077_U259);
  nand ginst10217 (P2_R1077_U261, P2_U3073, P2_U3434);
  not ginst10218 (P2_R1077_U262, P2_R1077_U92);
  or ginst10219 (P2_R1077_U263, P2_U3068, P2_U3440);
  or ginst10220 (P2_R1077_U264, P2_U3072, P2_U3437);
  not ginst10221 (P2_R1077_U265, P2_R1077_U59);
  nand ginst10222 (P2_R1077_U266, P2_R1077_U59, P2_R1077_U60);
  nand ginst10223 (P2_R1077_U267, P2_R1077_U266, P2_U3068);
  nand ginst10224 (P2_R1077_U268, P2_R1077_U265, P2_U3440);
  nand ginst10225 (P2_R1077_U269, P2_R1077_U8, P2_R1077_U92);
  not ginst10226 (P2_R1077_U27, P2_U3395);
  not ginst10227 (P2_R1077_U270, P2_R1077_U162);
  or ginst10228 (P2_R1077_U271, P2_U3075, P2_U3903);
  or ginst10229 (P2_R1077_U272, P2_U3080, P2_U3445);
  or ginst10230 (P2_R1077_U273, P2_U3074, P2_U3902);
  not ginst10231 (P2_R1077_U274, P2_R1077_U80);
  nand ginst10232 (P2_R1077_U275, P2_R1077_U274, P2_U3903);
  nand ginst10233 (P2_R1077_U276, P2_R1077_U275, P2_R1077_U90);
  nand ginst10234 (P2_R1077_U277, P2_R1077_U80, P2_R1077_U81);
  nand ginst10235 (P2_R1077_U278, P2_R1077_U276, P2_R1077_U277);
  nand ginst10236 (P2_R1077_U279, P2_R1077_U175, P2_R1077_U9);
  not ginst10237 (P2_R1077_U28, P2_U3067);
  nand ginst10238 (P2_R1077_U280, P2_U3074, P2_U3902);
  nand ginst10239 (P2_R1077_U281, P2_R1077_U278, P2_R1077_U279);
  or ginst10240 (P2_R1077_U282, P2_U3081, P2_U3443);
  or ginst10241 (P2_R1077_U283, P2_U3074, P2_U3902);
  nand ginst10242 (P2_R1077_U284, P2_R1077_U131, P2_R1077_U162, P2_R1077_U273);
  nand ginst10243 (P2_R1077_U285, P2_R1077_U281, P2_R1077_U283);
  not ginst10244 (P2_R1077_U286, P2_R1077_U159);
  or ginst10245 (P2_R1077_U287, P2_U3060, P2_U3901);
  nand ginst10246 (P2_R1077_U288, P2_R1077_U159, P2_R1077_U287);
  nand ginst10247 (P2_R1077_U289, P2_U3060, P2_U3901);
  not ginst10248 (P2_R1077_U29, P2_U3387);
  not ginst10249 (P2_R1077_U290, P2_R1077_U157);
  or ginst10250 (P2_R1077_U291, P2_U3065, P2_U3900);
  nand ginst10251 (P2_R1077_U292, P2_R1077_U157, P2_R1077_U291);
  nand ginst10252 (P2_R1077_U293, P2_U3065, P2_U3900);
  not ginst10253 (P2_R1077_U294, P2_R1077_U155);
  or ginst10254 (P2_R1077_U295, P2_U3057, P2_U3898);
  nand ginst10255 (P2_R1077_U296, P2_R1077_U173, P2_R1077_U176);
  not ginst10256 (P2_R1077_U297, P2_R1077_U86);
  or ginst10257 (P2_R1077_U298, P2_U3064, P2_U3899);
  nand ginst10258 (P2_R1077_U299, P2_R1077_U155, P2_R1077_U168, P2_R1077_U298);
  not ginst10259 (P2_R1077_U30, P2_U3076);
  not ginst10260 (P2_R1077_U300, P2_R1077_U153);
  or ginst10261 (P2_R1077_U301, P2_U3052, P2_U3896);
  nand ginst10262 (P2_R1077_U302, P2_U3052, P2_U3896);
  not ginst10263 (P2_R1077_U303, P2_R1077_U151);
  nand ginst10264 (P2_R1077_U304, P2_R1077_U151, P2_U3895);
  not ginst10265 (P2_R1077_U305, P2_R1077_U149);
  nand ginst10266 (P2_R1077_U306, P2_R1077_U155, P2_R1077_U298);
  not ginst10267 (P2_R1077_U307, P2_R1077_U89);
  or ginst10268 (P2_R1077_U308, P2_U3057, P2_U3898);
  nand ginst10269 (P2_R1077_U309, P2_R1077_U308, P2_R1077_U89);
  nand ginst10270 (P2_R1077_U31, P2_U3076, P2_U3387);
  nand ginst10271 (P2_R1077_U310, P2_R1077_U154, P2_R1077_U173, P2_R1077_U309);
  nand ginst10272 (P2_R1077_U311, P2_R1077_U173, P2_R1077_U307);
  nand ginst10273 (P2_R1077_U312, P2_U3056, P2_U3897);
  nand ginst10274 (P2_R1077_U313, P2_R1077_U168, P2_R1077_U311, P2_R1077_U312);
  or ginst10275 (P2_R1077_U314, P2_U3057, P2_U3898);
  nand ginst10276 (P2_R1077_U315, P2_R1077_U162, P2_R1077_U282);
  not ginst10277 (P2_R1077_U316, P2_R1077_U91);
  nand ginst10278 (P2_R1077_U317, P2_R1077_U9, P2_R1077_U91);
  nand ginst10279 (P2_R1077_U318, P2_R1077_U135, P2_R1077_U317);
  nand ginst10280 (P2_R1077_U319, P2_R1077_U278, P2_R1077_U317);
  not ginst10281 (P2_R1077_U32, P2_U3398);
  nand ginst10282 (P2_R1077_U320, P2_R1077_U319, P2_R1077_U453);
  or ginst10283 (P2_R1077_U321, P2_U3080, P2_U3445);
  nand ginst10284 (P2_R1077_U322, P2_R1077_U321, P2_R1077_U91);
  nand ginst10285 (P2_R1077_U323, P2_R1077_U136, P2_R1077_U322);
  nand ginst10286 (P2_R1077_U324, P2_R1077_U316, P2_R1077_U80);
  nand ginst10287 (P2_R1077_U325, P2_U3075, P2_U3903);
  nand ginst10288 (P2_R1077_U326, P2_R1077_U137, P2_R1077_U324);
  or ginst10289 (P2_R1077_U327, P2_U3077, P2_U3392);
  not ginst10290 (P2_R1077_U328, P2_R1077_U161);
  or ginst10291 (P2_R1077_U329, P2_U3080, P2_U3445);
  not ginst10292 (P2_R1077_U33, P2_U3063);
  or ginst10293 (P2_R1077_U330, P2_U3072, P2_U3437);
  nand ginst10294 (P2_R1077_U331, P2_R1077_U330, P2_R1077_U92);
  nand ginst10295 (P2_R1077_U332, P2_R1077_U138, P2_R1077_U331);
  nand ginst10296 (P2_R1077_U333, P2_R1077_U262, P2_R1077_U59);
  nand ginst10297 (P2_R1077_U334, P2_U3068, P2_U3440);
  nand ginst10298 (P2_R1077_U335, P2_R1077_U139, P2_R1077_U333);
  or ginst10299 (P2_R1077_U336, P2_U3072, P2_U3437);
  nand ginst10300 (P2_R1077_U337, P2_R1077_U167, P2_R1077_U250);
  not ginst10301 (P2_R1077_U338, P2_R1077_U93);
  or ginst10302 (P2_R1077_U339, P2_U3071, P2_U3425);
  nand ginst10303 (P2_R1077_U34, P2_U3059, P2_U3401);
  nand ginst10304 (P2_R1077_U340, P2_R1077_U339, P2_R1077_U93);
  nand ginst10305 (P2_R1077_U341, P2_R1077_U140, P2_R1077_U340);
  nand ginst10306 (P2_R1077_U342, P2_R1077_U172, P2_R1077_U338);
  nand ginst10307 (P2_R1077_U343, P2_U3079, P2_U3428);
  nand ginst10308 (P2_R1077_U344, P2_R1077_U141, P2_R1077_U342);
  or ginst10309 (P2_R1077_U345, P2_U3071, P2_U3425);
  or ginst10310 (P2_R1077_U346, P2_U3082, P2_U3416);
  nand ginst10311 (P2_R1077_U347, P2_R1077_U346, P2_R1077_U40);
  nand ginst10312 (P2_R1077_U348, P2_R1077_U142, P2_R1077_U347);
  nand ginst10313 (P2_R1077_U349, P2_R1077_U171, P2_R1077_U206);
  not ginst10314 (P2_R1077_U35, P2_U3404);
  nand ginst10315 (P2_R1077_U350, P2_U3061, P2_U3419);
  nand ginst10316 (P2_R1077_U351, P2_R1077_U143, P2_R1077_U349);
  nand ginst10317 (P2_R1077_U352, P2_R1077_U171, P2_R1077_U207);
  nand ginst10318 (P2_R1077_U353, P2_R1077_U204, P2_R1077_U65);
  nand ginst10319 (P2_R1077_U354, P2_R1077_U214, P2_R1077_U22);
  nand ginst10320 (P2_R1077_U355, P2_R1077_U228, P2_R1077_U34);
  nand ginst10321 (P2_R1077_U356, P2_R1077_U180, P2_R1077_U231);
  nand ginst10322 (P2_R1077_U357, P2_R1077_U173, P2_R1077_U314);
  nand ginst10323 (P2_R1077_U358, P2_R1077_U176, P2_R1077_U298);
  nand ginst10324 (P2_R1077_U359, P2_R1077_U329, P2_R1077_U80);
  not ginst10325 (P2_R1077_U36, P2_U3413);
  nand ginst10326 (P2_R1077_U360, P2_R1077_U282, P2_R1077_U77);
  nand ginst10327 (P2_R1077_U361, P2_R1077_U336, P2_R1077_U59);
  nand ginst10328 (P2_R1077_U362, P2_R1077_U172, P2_R1077_U345);
  nand ginst10329 (P2_R1077_U363, P2_R1077_U250, P2_R1077_U68);
  nand ginst10330 (P2_R1077_U364, P2_U3053, P2_U3895);
  nand ginst10331 (P2_R1077_U365, P2_R1077_U168, P2_R1077_U296);
  nand ginst10332 (P2_R1077_U366, P2_R1077_U295, P2_U3056);
  nand ginst10333 (P2_R1077_U367, P2_R1077_U295, P2_U3897);
  nand ginst10334 (P2_R1077_U368, P2_R1077_U168, P2_R1077_U296, P2_R1077_U301);
  nand ginst10335 (P2_R1077_U369, P2_R1077_U133, P2_R1077_U155, P2_R1077_U168);
  not ginst10336 (P2_R1077_U37, P2_U3083);
  nand ginst10337 (P2_R1077_U370, P2_R1077_U297, P2_R1077_U301);
  nand ginst10338 (P2_R1077_U371, P2_R1077_U39, P2_U3082);
  nand ginst10339 (P2_R1077_U372, P2_R1077_U38, P2_U3416);
  nand ginst10340 (P2_R1077_U373, P2_R1077_U371, P2_R1077_U372);
  nand ginst10341 (P2_R1077_U374, P2_R1077_U352, P2_R1077_U40);
  nand ginst10342 (P2_R1077_U375, P2_R1077_U206, P2_R1077_U373);
  nand ginst10343 (P2_R1077_U376, P2_R1077_U36, P2_U3083);
  nand ginst10344 (P2_R1077_U377, P2_R1077_U37, P2_U3413);
  nand ginst10345 (P2_R1077_U378, P2_R1077_U376, P2_R1077_U377);
  nand ginst10346 (P2_R1077_U379, P2_R1077_U144, P2_R1077_U353);
  not ginst10347 (P2_R1077_U38, P2_U3082);
  nand ginst10348 (P2_R1077_U380, P2_R1077_U203, P2_R1077_U378);
  nand ginst10349 (P2_R1077_U381, P2_R1077_U23, P2_U3069);
  nand ginst10350 (P2_R1077_U382, P2_R1077_U21, P2_U3410);
  nand ginst10351 (P2_R1077_U383, P2_R1077_U19, P2_U3070);
  nand ginst10352 (P2_R1077_U384, P2_R1077_U20, P2_U3407);
  nand ginst10353 (P2_R1077_U385, P2_R1077_U383, P2_R1077_U384);
  nand ginst10354 (P2_R1077_U386, P2_R1077_U354, P2_R1077_U41);
  nand ginst10355 (P2_R1077_U387, P2_R1077_U195, P2_R1077_U385);
  nand ginst10356 (P2_R1077_U388, P2_R1077_U35, P2_U3066);
  nand ginst10357 (P2_R1077_U389, P2_R1077_U26, P2_U3404);
  not ginst10358 (P2_R1077_U39, P2_U3416);
  nand ginst10359 (P2_R1077_U390, P2_R1077_U24, P2_U3059);
  nand ginst10360 (P2_R1077_U391, P2_R1077_U25, P2_U3401);
  nand ginst10361 (P2_R1077_U392, P2_R1077_U390, P2_R1077_U391);
  nand ginst10362 (P2_R1077_U393, P2_R1077_U355, P2_R1077_U44);
  nand ginst10363 (P2_R1077_U394, P2_R1077_U221, P2_R1077_U392);
  nand ginst10364 (P2_R1077_U395, P2_R1077_U32, P2_U3063);
  nand ginst10365 (P2_R1077_U396, P2_R1077_U33, P2_U3398);
  nand ginst10366 (P2_R1077_U397, P2_R1077_U395, P2_R1077_U396);
  nand ginst10367 (P2_R1077_U398, P2_R1077_U145, P2_R1077_U356);
  nand ginst10368 (P2_R1077_U399, P2_R1077_U230, P2_R1077_U397);
  and ginst10369 (P2_R1077_U4, P2_R1077_U178, P2_R1077_U179);
  nand ginst10370 (P2_R1077_U40, P2_R1077_U205, P2_R1077_U65);
  nand ginst10371 (P2_R1077_U400, P2_R1077_U27, P2_U3067);
  nand ginst10372 (P2_R1077_U401, P2_R1077_U28, P2_U3395);
  nand ginst10373 (P2_R1077_U402, P2_R1077_U147, P2_U3054);
  nand ginst10374 (P2_R1077_U403, P2_R1077_U146, P2_U3904);
  nand ginst10375 (P2_R1077_U404, P2_R1077_U147, P2_U3054);
  nand ginst10376 (P2_R1077_U405, P2_R1077_U146, P2_U3904);
  nand ginst10377 (P2_R1077_U406, P2_R1077_U404, P2_R1077_U405);
  nand ginst10378 (P2_R1077_U407, P2_R1077_U148, P2_R1077_U149);
  nand ginst10379 (P2_R1077_U408, P2_R1077_U305, P2_R1077_U406);
  nand ginst10380 (P2_R1077_U409, P2_R1077_U88, P2_U3053);
  nand ginst10381 (P2_R1077_U41, P2_R1077_U117, P2_R1077_U193);
  nand ginst10382 (P2_R1077_U410, P2_R1077_U87, P2_U3895);
  nand ginst10383 (P2_R1077_U411, P2_R1077_U88, P2_U3053);
  nand ginst10384 (P2_R1077_U412, P2_R1077_U87, P2_U3895);
  nand ginst10385 (P2_R1077_U413, P2_R1077_U411, P2_R1077_U412);
  nand ginst10386 (P2_R1077_U414, P2_R1077_U150, P2_R1077_U151);
  nand ginst10387 (P2_R1077_U415, P2_R1077_U303, P2_R1077_U413);
  nand ginst10388 (P2_R1077_U416, P2_R1077_U46, P2_U3052);
  nand ginst10389 (P2_R1077_U417, P2_R1077_U47, P2_U3896);
  nand ginst10390 (P2_R1077_U418, P2_R1077_U46, P2_U3052);
  nand ginst10391 (P2_R1077_U419, P2_R1077_U47, P2_U3896);
  nand ginst10392 (P2_R1077_U42, P2_R1077_U182, P2_R1077_U183);
  nand ginst10393 (P2_R1077_U420, P2_R1077_U418, P2_R1077_U419);
  nand ginst10394 (P2_R1077_U421, P2_R1077_U152, P2_R1077_U153);
  nand ginst10395 (P2_R1077_U422, P2_R1077_U300, P2_R1077_U420);
  nand ginst10396 (P2_R1077_U423, P2_R1077_U49, P2_U3056);
  nand ginst10397 (P2_R1077_U424, P2_R1077_U48, P2_U3897);
  nand ginst10398 (P2_R1077_U425, P2_R1077_U50, P2_U3057);
  nand ginst10399 (P2_R1077_U426, P2_R1077_U51, P2_U3898);
  nand ginst10400 (P2_R1077_U427, P2_R1077_U425, P2_R1077_U426);
  nand ginst10401 (P2_R1077_U428, P2_R1077_U357, P2_R1077_U89);
  nand ginst10402 (P2_R1077_U429, P2_R1077_U307, P2_R1077_U427);
  nand ginst10403 (P2_R1077_U43, P2_U3077, P2_U3392);
  nand ginst10404 (P2_R1077_U430, P2_R1077_U52, P2_U3064);
  nand ginst10405 (P2_R1077_U431, P2_R1077_U53, P2_U3899);
  nand ginst10406 (P2_R1077_U432, P2_R1077_U430, P2_R1077_U431);
  nand ginst10407 (P2_R1077_U433, P2_R1077_U155, P2_R1077_U358);
  nand ginst10408 (P2_R1077_U434, P2_R1077_U294, P2_R1077_U432);
  nand ginst10409 (P2_R1077_U435, P2_R1077_U84, P2_U3065);
  nand ginst10410 (P2_R1077_U436, P2_R1077_U85, P2_U3900);
  nand ginst10411 (P2_R1077_U437, P2_R1077_U84, P2_U3065);
  nand ginst10412 (P2_R1077_U438, P2_R1077_U85, P2_U3900);
  nand ginst10413 (P2_R1077_U439, P2_R1077_U437, P2_R1077_U438);
  nand ginst10414 (P2_R1077_U44, P2_R1077_U122, P2_R1077_U219);
  nand ginst10415 (P2_R1077_U440, P2_R1077_U156, P2_R1077_U157);
  nand ginst10416 (P2_R1077_U441, P2_R1077_U290, P2_R1077_U439);
  nand ginst10417 (P2_R1077_U442, P2_R1077_U82, P2_U3060);
  nand ginst10418 (P2_R1077_U443, P2_R1077_U83, P2_U3901);
  nand ginst10419 (P2_R1077_U444, P2_R1077_U82, P2_U3060);
  nand ginst10420 (P2_R1077_U445, P2_R1077_U83, P2_U3901);
  nand ginst10421 (P2_R1077_U446, P2_R1077_U444, P2_R1077_U445);
  nand ginst10422 (P2_R1077_U447, P2_R1077_U158, P2_R1077_U159);
  nand ginst10423 (P2_R1077_U448, P2_R1077_U286, P2_R1077_U446);
  nand ginst10424 (P2_R1077_U449, P2_R1077_U54, P2_U3074);
  nand ginst10425 (P2_R1077_U45, P2_R1077_U215, P2_R1077_U216);
  nand ginst10426 (P2_R1077_U450, P2_R1077_U55, P2_U3902);
  nand ginst10427 (P2_R1077_U451, P2_R1077_U54, P2_U3074);
  nand ginst10428 (P2_R1077_U452, P2_R1077_U55, P2_U3902);
  nand ginst10429 (P2_R1077_U453, P2_R1077_U451, P2_R1077_U452);
  nand ginst10430 (P2_R1077_U454, P2_R1077_U81, P2_U3075);
  nand ginst10431 (P2_R1077_U455, P2_R1077_U90, P2_U3903);
  nand ginst10432 (P2_R1077_U456, P2_R1077_U161, P2_R1077_U182);
  nand ginst10433 (P2_R1077_U457, P2_R1077_U31, P2_R1077_U328);
  nand ginst10434 (P2_R1077_U458, P2_R1077_U78, P2_U3080);
  nand ginst10435 (P2_R1077_U459, P2_R1077_U79, P2_U3445);
  not ginst10436 (P2_R1077_U46, P2_U3896);
  nand ginst10437 (P2_R1077_U460, P2_R1077_U458, P2_R1077_U459);
  nand ginst10438 (P2_R1077_U461, P2_R1077_U359, P2_R1077_U91);
  nand ginst10439 (P2_R1077_U462, P2_R1077_U316, P2_R1077_U460);
  nand ginst10440 (P2_R1077_U463, P2_R1077_U75, P2_U3081);
  nand ginst10441 (P2_R1077_U464, P2_R1077_U76, P2_U3443);
  nand ginst10442 (P2_R1077_U465, P2_R1077_U463, P2_R1077_U464);
  nand ginst10443 (P2_R1077_U466, P2_R1077_U162, P2_R1077_U360);
  nand ginst10444 (P2_R1077_U467, P2_R1077_U270, P2_R1077_U465);
  nand ginst10445 (P2_R1077_U468, P2_R1077_U60, P2_U3068);
  nand ginst10446 (P2_R1077_U469, P2_R1077_U58, P2_U3440);
  not ginst10447 (P2_R1077_U47, P2_U3052);
  nand ginst10448 (P2_R1077_U470, P2_R1077_U56, P2_U3072);
  nand ginst10449 (P2_R1077_U471, P2_R1077_U57, P2_U3437);
  nand ginst10450 (P2_R1077_U472, P2_R1077_U470, P2_R1077_U471);
  nand ginst10451 (P2_R1077_U473, P2_R1077_U361, P2_R1077_U92);
  nand ginst10452 (P2_R1077_U474, P2_R1077_U262, P2_R1077_U472);
  nand ginst10453 (P2_R1077_U475, P2_R1077_U73, P2_U3073);
  nand ginst10454 (P2_R1077_U476, P2_R1077_U74, P2_U3434);
  nand ginst10455 (P2_R1077_U477, P2_R1077_U73, P2_U3073);
  nand ginst10456 (P2_R1077_U478, P2_R1077_U74, P2_U3434);
  nand ginst10457 (P2_R1077_U479, P2_R1077_U477, P2_R1077_U478);
  not ginst10458 (P2_R1077_U48, P2_U3056);
  nand ginst10459 (P2_R1077_U480, P2_R1077_U163, P2_R1077_U164);
  nand ginst10460 (P2_R1077_U481, P2_R1077_U258, P2_R1077_U479);
  nand ginst10461 (P2_R1077_U482, P2_R1077_U71, P2_U3078);
  nand ginst10462 (P2_R1077_U483, P2_R1077_U72, P2_U3431);
  nand ginst10463 (P2_R1077_U484, P2_R1077_U71, P2_U3078);
  nand ginst10464 (P2_R1077_U485, P2_R1077_U72, P2_U3431);
  nand ginst10465 (P2_R1077_U486, P2_R1077_U484, P2_R1077_U485);
  nand ginst10466 (P2_R1077_U487, P2_R1077_U165, P2_R1077_U166);
  nand ginst10467 (P2_R1077_U488, P2_R1077_U254, P2_R1077_U486);
  nand ginst10468 (P2_R1077_U489, P2_R1077_U61, P2_U3079);
  not ginst10469 (P2_R1077_U49, P2_U3897);
  nand ginst10470 (P2_R1077_U490, P2_R1077_U62, P2_U3428);
  nand ginst10471 (P2_R1077_U491, P2_R1077_U69, P2_U3071);
  nand ginst10472 (P2_R1077_U492, P2_R1077_U70, P2_U3425);
  nand ginst10473 (P2_R1077_U493, P2_R1077_U491, P2_R1077_U492);
  nand ginst10474 (P2_R1077_U494, P2_R1077_U362, P2_R1077_U93);
  nand ginst10475 (P2_R1077_U495, P2_R1077_U338, P2_R1077_U493);
  nand ginst10476 (P2_R1077_U496, P2_R1077_U66, P2_U3062);
  nand ginst10477 (P2_R1077_U497, P2_R1077_U67, P2_U3422);
  nand ginst10478 (P2_R1077_U498, P2_R1077_U496, P2_R1077_U497);
  nand ginst10479 (P2_R1077_U499, P2_R1077_U167, P2_R1077_U363);
  and ginst10480 (P2_R1077_U5, P2_R1077_U196, P2_R1077_U197);
  not ginst10481 (P2_R1077_U50, P2_U3898);
  nand ginst10482 (P2_R1077_U500, P2_R1077_U244, P2_R1077_U498);
  nand ginst10483 (P2_R1077_U501, P2_R1077_U63, P2_U3061);
  nand ginst10484 (P2_R1077_U502, P2_R1077_U64, P2_U3419);
  nand ginst10485 (P2_R1077_U503, P2_R1077_U29, P2_U3076);
  nand ginst10486 (P2_R1077_U504, P2_R1077_U30, P2_U3387);
  not ginst10487 (P2_R1077_U51, P2_U3057);
  not ginst10488 (P2_R1077_U52, P2_U3899);
  not ginst10489 (P2_R1077_U53, P2_U3064);
  not ginst10490 (P2_R1077_U54, P2_U3902);
  not ginst10491 (P2_R1077_U55, P2_U3074);
  not ginst10492 (P2_R1077_U56, P2_U3437);
  not ginst10493 (P2_R1077_U57, P2_U3072);
  not ginst10494 (P2_R1077_U58, P2_U3068);
  nand ginst10495 (P2_R1077_U59, P2_U3072, P2_U3437);
  and ginst10496 (P2_R1077_U6, P2_R1077_U236, P2_R1077_U237);
  not ginst10497 (P2_R1077_U60, P2_U3440);
  not ginst10498 (P2_R1077_U61, P2_U3428);
  not ginst10499 (P2_R1077_U62, P2_U3079);
  not ginst10500 (P2_R1077_U63, P2_U3419);
  not ginst10501 (P2_R1077_U64, P2_U3061);
  nand ginst10502 (P2_R1077_U65, P2_U3083, P2_U3413);
  not ginst10503 (P2_R1077_U66, P2_U3422);
  not ginst10504 (P2_R1077_U67, P2_U3062);
  nand ginst10505 (P2_R1077_U68, P2_U3062, P2_U3422);
  not ginst10506 (P2_R1077_U69, P2_U3425);
  and ginst10507 (P2_R1077_U7, P2_R1077_U245, P2_R1077_U246);
  not ginst10508 (P2_R1077_U70, P2_U3071);
  not ginst10509 (P2_R1077_U71, P2_U3431);
  not ginst10510 (P2_R1077_U72, P2_U3078);
  not ginst10511 (P2_R1077_U73, P2_U3434);
  not ginst10512 (P2_R1077_U74, P2_U3073);
  not ginst10513 (P2_R1077_U75, P2_U3443);
  not ginst10514 (P2_R1077_U76, P2_U3081);
  nand ginst10515 (P2_R1077_U77, P2_U3081, P2_U3443);
  not ginst10516 (P2_R1077_U78, P2_U3445);
  not ginst10517 (P2_R1077_U79, P2_U3080);
  and ginst10518 (P2_R1077_U8, P2_R1077_U263, P2_R1077_U264);
  nand ginst10519 (P2_R1077_U80, P2_U3080, P2_U3445);
  not ginst10520 (P2_R1077_U81, P2_U3903);
  not ginst10521 (P2_R1077_U82, P2_U3901);
  not ginst10522 (P2_R1077_U83, P2_U3060);
  not ginst10523 (P2_R1077_U84, P2_U3900);
  not ginst10524 (P2_R1077_U85, P2_U3065);
  nand ginst10525 (P2_R1077_U86, P2_U3056, P2_U3897);
  not ginst10526 (P2_R1077_U87, P2_U3053);
  not ginst10527 (P2_R1077_U88, P2_U3895);
  nand ginst10528 (P2_R1077_U89, P2_R1077_U176, P2_R1077_U306);
  and ginst10529 (P2_R1077_U9, P2_R1077_U271, P2_R1077_U272);
  not ginst10530 (P2_R1077_U90, P2_U3075);
  nand ginst10531 (P2_R1077_U91, P2_R1077_U315, P2_R1077_U77);
  nand ginst10532 (P2_R1077_U92, P2_R1077_U260, P2_R1077_U261);
  nand ginst10533 (P2_R1077_U93, P2_R1077_U337, P2_R1077_U68);
  nand ginst10534 (P2_R1077_U94, P2_R1077_U456, P2_R1077_U457);
  nand ginst10535 (P2_R1077_U95, P2_R1077_U503, P2_R1077_U504);
  nand ginst10536 (P2_R1077_U96, P2_R1077_U374, P2_R1077_U375);
  nand ginst10537 (P2_R1077_U97, P2_R1077_U379, P2_R1077_U380);
  nand ginst10538 (P2_R1077_U98, P2_R1077_U386, P2_R1077_U387);
  nand ginst10539 (P2_R1077_U99, P2_R1077_U393, P2_R1077_U394);
  and ginst10540 (P2_R1095_U10, P2_R1095_U194, P2_R1095_U281);
  nand ginst10541 (P2_R1095_U100, P2_R1095_U424, P2_R1095_U425);
  nand ginst10542 (P2_R1095_U101, P2_R1095_U440, P2_R1095_U441);
  nand ginst10543 (P2_R1095_U102, P2_R1095_U445, P2_R1095_U446);
  nand ginst10544 (P2_R1095_U103, P2_R1095_U450, P2_R1095_U451);
  nand ginst10545 (P2_R1095_U104, P2_R1095_U455, P2_R1095_U456);
  nand ginst10546 (P2_R1095_U105, P2_R1095_U460, P2_R1095_U461);
  nand ginst10547 (P2_R1095_U106, P2_R1095_U476, P2_R1095_U477);
  nand ginst10548 (P2_R1095_U107, P2_R1095_U481, P2_R1095_U482);
  nand ginst10549 (P2_R1095_U108, P2_R1095_U364, P2_R1095_U365);
  nand ginst10550 (P2_R1095_U109, P2_R1095_U373, P2_R1095_U374);
  and ginst10551 (P2_R1095_U11, P2_R1095_U282, P2_R1095_U283);
  nand ginst10552 (P2_R1095_U110, P2_R1095_U380, P2_R1095_U381);
  nand ginst10553 (P2_R1095_U111, P2_R1095_U384, P2_R1095_U385);
  nand ginst10554 (P2_R1095_U112, P2_R1095_U393, P2_R1095_U394);
  nand ginst10555 (P2_R1095_U113, P2_R1095_U414, P2_R1095_U415);
  nand ginst10556 (P2_R1095_U114, P2_R1095_U431, P2_R1095_U432);
  nand ginst10557 (P2_R1095_U115, P2_R1095_U435, P2_R1095_U436);
  nand ginst10558 (P2_R1095_U116, P2_R1095_U467, P2_R1095_U468);
  nand ginst10559 (P2_R1095_U117, P2_R1095_U471, P2_R1095_U472);
  nand ginst10560 (P2_R1095_U118, P2_R1095_U488, P2_R1095_U489);
  and ginst10561 (P2_R1095_U119, P2_R1095_U196, P2_R1095_U206);
  and ginst10562 (P2_R1095_U12, P2_R1095_U195, P2_R1095_U299);
  and ginst10563 (P2_R1095_U120, P2_R1095_U208, P2_R1095_U209);
  and ginst10564 (P2_R1095_U121, P2_R1095_U13, P2_R1095_U14);
  and ginst10565 (P2_R1095_U122, P2_R1095_U222, P2_R1095_U340);
  and ginst10566 (P2_R1095_U123, P2_R1095_U122, P2_R1095_U342);
  and ginst10567 (P2_R1095_U124, P2_R1095_U27, P2_R1095_U366, P2_R1095_U367);
  and ginst10568 (P2_R1095_U125, P2_R1095_U198, P2_R1095_U370);
  and ginst10569 (P2_R1095_U126, P2_R1095_U237, P2_R1095_U6);
  and ginst10570 (P2_R1095_U127, P2_R1095_U197, P2_R1095_U377);
  and ginst10571 (P2_R1095_U128, P2_R1095_U35, P2_R1095_U386, P2_R1095_U387);
  and ginst10572 (P2_R1095_U129, P2_R1095_U196, P2_R1095_U390);
  and ginst10573 (P2_R1095_U13, P2_R1095_U197, P2_R1095_U210, P2_R1095_U215);
  and ginst10574 (P2_R1095_U130, P2_R1095_U15, P2_R1095_U251);
  and ginst10575 (P2_R1095_U131, P2_R1095_U252, P2_R1095_U343);
  and ginst10576 (P2_R1095_U132, P2_R1095_U262, P2_R1095_U8);
  and ginst10577 (P2_R1095_U133, P2_R1095_U10, P2_R1095_U286);
  and ginst10578 (P2_R1095_U134, P2_R1095_U301, P2_R1095_U302);
  and ginst10579 (P2_R1095_U135, P2_R1095_U303, P2_R1095_U397);
  and ginst10580 (P2_R1095_U136, P2_R1095_U16, P2_R1095_U301, P2_R1095_U302, P2_R1095_U304);
  and ginst10581 (P2_R1095_U137, P2_R1095_U165, P2_R1095_U359);
  nand ginst10582 (P2_R1095_U138, P2_R1095_U402, P2_R1095_U403);
  and ginst10583 (P2_R1095_U139, P2_R1095_U407, P2_R1095_U408, P2_R1095_U53);
  and ginst10584 (P2_R1095_U14, P2_R1095_U198, P2_R1095_U220);
  and ginst10585 (P2_R1095_U140, P2_R1095_U195, P2_R1095_U411);
  nand ginst10586 (P2_R1095_U141, P2_R1095_U416, P2_R1095_U417);
  nand ginst10587 (P2_R1095_U142, P2_R1095_U421, P2_R1095_U422);
  and ginst10588 (P2_R1095_U143, P2_R1095_U11, P2_R1095_U313);
  and ginst10589 (P2_R1095_U144, P2_R1095_U194, P2_R1095_U428);
  nand ginst10590 (P2_R1095_U145, P2_R1095_U437, P2_R1095_U438);
  nand ginst10591 (P2_R1095_U146, P2_R1095_U442, P2_R1095_U443);
  nand ginst10592 (P2_R1095_U147, P2_R1095_U447, P2_R1095_U448);
  nand ginst10593 (P2_R1095_U148, P2_R1095_U452, P2_R1095_U453);
  nand ginst10594 (P2_R1095_U149, P2_R1095_U457, P2_R1095_U458);
  and ginst10595 (P2_R1095_U15, P2_R1095_U192, P2_R1095_U224, P2_R1095_U244);
  and ginst10596 (P2_R1095_U150, P2_R1095_U324, P2_R1095_U9);
  and ginst10597 (P2_R1095_U151, P2_R1095_U193, P2_R1095_U464);
  nand ginst10598 (P2_R1095_U152, P2_R1095_U473, P2_R1095_U474);
  nand ginst10599 (P2_R1095_U153, P2_R1095_U478, P2_R1095_U479);
  and ginst10600 (P2_R1095_U154, P2_R1095_U333, P2_R1095_U7);
  and ginst10601 (P2_R1095_U155, P2_R1095_U192, P2_R1095_U485);
  and ginst10602 (P2_R1095_U156, P2_R1095_U362, P2_R1095_U363);
  nand ginst10603 (P2_R1095_U157, P2_R1095_U123, P2_R1095_U341);
  and ginst10604 (P2_R1095_U158, P2_R1095_U371, P2_R1095_U372);
  and ginst10605 (P2_R1095_U159, P2_R1095_U378, P2_R1095_U379);
  and ginst10606 (P2_R1095_U16, P2_R1095_U398, P2_R1095_U399);
  and ginst10607 (P2_R1095_U160, P2_R1095_U382, P2_R1095_U383);
  nand ginst10608 (P2_R1095_U161, P2_R1095_U120, P2_R1095_U344);
  and ginst10609 (P2_R1095_U162, P2_R1095_U391, P2_R1095_U392);
  not ginst10610 (P2_R1095_U163, P2_U3904);
  not ginst10611 (P2_R1095_U164, P2_U3054);
  and ginst10612 (P2_R1095_U165, P2_R1095_U400, P2_R1095_U401);
  nand ginst10613 (P2_R1095_U166, P2_R1095_U134, P2_R1095_U360);
  and ginst10614 (P2_R1095_U167, P2_R1095_U412, P2_R1095_U413);
  nand ginst10615 (P2_R1095_U168, P2_R1095_U292, P2_R1095_U293);
  nand ginst10616 (P2_R1095_U169, P2_R1095_U288, P2_R1095_U289);
  nand ginst10617 (P2_R1095_U17, P2_R1095_U331, P2_R1095_U334);
  and ginst10618 (P2_R1095_U170, P2_R1095_U429, P2_R1095_U430);
  and ginst10619 (P2_R1095_U171, P2_R1095_U433, P2_R1095_U434);
  nand ginst10620 (P2_R1095_U172, P2_R1095_U278, P2_R1095_U279);
  nand ginst10621 (P2_R1095_U173, P2_R1095_U274, P2_R1095_U275);
  not ginst10622 (P2_R1095_U174, P2_U3392);
  nand ginst10623 (P2_R1095_U175, P2_R1095_U97, P2_U3387);
  nand ginst10624 (P2_R1095_U176, P2_R1095_U187, P2_R1095_U271, P2_R1095_U339);
  not ginst10625 (P2_R1095_U177, P2_U3443);
  nand ginst10626 (P2_R1095_U178, P2_R1095_U268, P2_R1095_U269);
  nand ginst10627 (P2_R1095_U179, P2_R1095_U264, P2_R1095_U265);
  nand ginst10628 (P2_R1095_U18, P2_R1095_U322, P2_R1095_U325);
  and ginst10629 (P2_R1095_U180, P2_R1095_U465, P2_R1095_U466);
  and ginst10630 (P2_R1095_U181, P2_R1095_U469, P2_R1095_U470);
  nand ginst10631 (P2_R1095_U182, P2_R1095_U254, P2_R1095_U255);
  nand ginst10632 (P2_R1095_U183, P2_R1095_U131, P2_R1095_U353);
  nand ginst10633 (P2_R1095_U184, P2_R1095_U351, P2_R1095_U62);
  and ginst10634 (P2_R1095_U185, P2_R1095_U486, P2_R1095_U487);
  nand ginst10635 (P2_R1095_U186, P2_R1095_U135, P2_R1095_U166);
  nand ginst10636 (P2_R1095_U187, P2_R1095_U177, P2_R1095_U178);
  nand ginst10637 (P2_R1095_U188, P2_R1095_U174, P2_R1095_U175);
  not ginst10638 (P2_R1095_U189, P2_R1095_U53);
  nand ginst10639 (P2_R1095_U19, P2_R1095_U311, P2_R1095_U314);
  not ginst10640 (P2_R1095_U190, P2_R1095_U35);
  not ginst10641 (P2_R1095_U191, P2_R1095_U27);
  nand ginst10642 (P2_R1095_U192, P2_R1095_U57, P2_U3419);
  nand ginst10643 (P2_R1095_U193, P2_R1095_U69, P2_U3434);
  nand ginst10644 (P2_R1095_U194, P2_R1095_U83, P2_U3901);
  nand ginst10645 (P2_R1095_U195, P2_R1095_U52, P2_U3897);
  nand ginst10646 (P2_R1095_U196, P2_R1095_U34, P2_U3395);
  nand ginst10647 (P2_R1095_U197, P2_R1095_U42, P2_U3404);
  nand ginst10648 (P2_R1095_U198, P2_R1095_U26, P2_U3410);
  not ginst10649 (P2_R1095_U199, P2_R1095_U71);
  nand ginst10650 (P2_R1095_U20, P2_R1095_U305, P2_R1095_U357);
  not ginst10651 (P2_R1095_U200, P2_R1095_U85);
  not ginst10652 (P2_R1095_U201, P2_R1095_U44);
  not ginst10653 (P2_R1095_U202, P2_R1095_U59);
  not ginst10654 (P2_R1095_U203, P2_R1095_U175);
  nand ginst10655 (P2_R1095_U204, P2_R1095_U175, P2_U3077);
  not ginst10656 (P2_R1095_U205, P2_R1095_U50);
  nand ginst10657 (P2_R1095_U206, P2_R1095_U36, P2_U3398);
  nand ginst10658 (P2_R1095_U207, P2_R1095_U35, P2_R1095_U36);
  nand ginst10659 (P2_R1095_U208, P2_R1095_U207, P2_R1095_U40);
  nand ginst10660 (P2_R1095_U209, P2_R1095_U190, P2_U3063);
  nand ginst10661 (P2_R1095_U21, P2_R1095_U137, P2_R1095_U186);
  nand ginst10662 (P2_R1095_U210, P2_R1095_U41, P2_U3407);
  nand ginst10663 (P2_R1095_U211, P2_R1095_U30, P2_U3070);
  nand ginst10664 (P2_R1095_U212, P2_R1095_U29, P2_U3066);
  nand ginst10665 (P2_R1095_U213, P2_R1095_U197, P2_R1095_U201);
  nand ginst10666 (P2_R1095_U214, P2_R1095_U213, P2_R1095_U6);
  nand ginst10667 (P2_R1095_U215, P2_R1095_U43, P2_U3401);
  nand ginst10668 (P2_R1095_U216, P2_R1095_U41, P2_U3407);
  nand ginst10669 (P2_R1095_U217, P2_R1095_U13, P2_R1095_U161);
  not ginst10670 (P2_R1095_U218, P2_R1095_U45);
  not ginst10671 (P2_R1095_U219, P2_R1095_U48);
  nand ginst10672 (P2_R1095_U22, P2_R1095_U242, P2_R1095_U347);
  nand ginst10673 (P2_R1095_U220, P2_R1095_U28, P2_U3413);
  nand ginst10674 (P2_R1095_U221, P2_R1095_U27, P2_R1095_U28);
  nand ginst10675 (P2_R1095_U222, P2_R1095_U191, P2_U3083);
  not ginst10676 (P2_R1095_U223, P2_R1095_U157);
  nand ginst10677 (P2_R1095_U224, P2_R1095_U47, P2_U3416);
  nand ginst10678 (P2_R1095_U225, P2_R1095_U224, P2_R1095_U59);
  nand ginst10679 (P2_R1095_U226, P2_R1095_U219, P2_R1095_U27);
  nand ginst10680 (P2_R1095_U227, P2_R1095_U125, P2_R1095_U226);
  nand ginst10681 (P2_R1095_U228, P2_R1095_U198, P2_R1095_U48);
  nand ginst10682 (P2_R1095_U229, P2_R1095_U124, P2_R1095_U228);
  nand ginst10683 (P2_R1095_U23, P2_R1095_U235, P2_R1095_U238);
  nand ginst10684 (P2_R1095_U230, P2_R1095_U198, P2_R1095_U27);
  nand ginst10685 (P2_R1095_U231, P2_R1095_U161, P2_R1095_U215);
  not ginst10686 (P2_R1095_U232, P2_R1095_U49);
  nand ginst10687 (P2_R1095_U233, P2_R1095_U29, P2_U3066);
  nand ginst10688 (P2_R1095_U234, P2_R1095_U232, P2_R1095_U233);
  nand ginst10689 (P2_R1095_U235, P2_R1095_U127, P2_R1095_U234);
  nand ginst10690 (P2_R1095_U236, P2_R1095_U197, P2_R1095_U49);
  nand ginst10691 (P2_R1095_U237, P2_R1095_U41, P2_U3407);
  nand ginst10692 (P2_R1095_U238, P2_R1095_U126, P2_R1095_U236);
  nand ginst10693 (P2_R1095_U239, P2_R1095_U29, P2_U3066);
  nand ginst10694 (P2_R1095_U24, P2_R1095_U227, P2_R1095_U229);
  nand ginst10695 (P2_R1095_U240, P2_R1095_U197, P2_R1095_U239);
  nand ginst10696 (P2_R1095_U241, P2_R1095_U215, P2_R1095_U44);
  nand ginst10697 (P2_R1095_U242, P2_R1095_U129, P2_R1095_U348);
  nand ginst10698 (P2_R1095_U243, P2_R1095_U196, P2_R1095_U35);
  nand ginst10699 (P2_R1095_U244, P2_R1095_U56, P2_U3422);
  nand ginst10700 (P2_R1095_U245, P2_R1095_U60, P2_U3062);
  nand ginst10701 (P2_R1095_U246, P2_R1095_U58, P2_U3061);
  nand ginst10702 (P2_R1095_U247, P2_R1095_U192, P2_R1095_U202);
  nand ginst10703 (P2_R1095_U248, P2_R1095_U247, P2_R1095_U7);
  nand ginst10704 (P2_R1095_U249, P2_R1095_U56, P2_U3422);
  nand ginst10705 (P2_R1095_U25, P2_R1095_U175, P2_R1095_U337);
  not ginst10706 (P2_R1095_U250, P2_R1095_U62);
  nand ginst10707 (P2_R1095_U251, P2_R1095_U55, P2_U3425);
  nand ginst10708 (P2_R1095_U252, P2_R1095_U61, P2_U3071);
  nand ginst10709 (P2_R1095_U253, P2_R1095_U64, P2_U3428);
  nand ginst10710 (P2_R1095_U254, P2_R1095_U183, P2_R1095_U253);
  nand ginst10711 (P2_R1095_U255, P2_R1095_U63, P2_U3079);
  not ginst10712 (P2_R1095_U256, P2_R1095_U182);
  nand ginst10713 (P2_R1095_U257, P2_R1095_U68, P2_U3437);
  nand ginst10714 (P2_R1095_U258, P2_R1095_U65, P2_U3072);
  nand ginst10715 (P2_R1095_U259, P2_R1095_U66, P2_U3073);
  not ginst10716 (P2_R1095_U26, P2_U3069);
  nand ginst10717 (P2_R1095_U260, P2_R1095_U199, P2_R1095_U8);
  nand ginst10718 (P2_R1095_U261, P2_R1095_U260, P2_R1095_U9);
  nand ginst10719 (P2_R1095_U262, P2_R1095_U70, P2_U3431);
  nand ginst10720 (P2_R1095_U263, P2_R1095_U68, P2_U3437);
  nand ginst10721 (P2_R1095_U264, P2_R1095_U132, P2_R1095_U182);
  nand ginst10722 (P2_R1095_U265, P2_R1095_U261, P2_R1095_U263);
  not ginst10723 (P2_R1095_U266, P2_R1095_U179);
  nand ginst10724 (P2_R1095_U267, P2_R1095_U73, P2_U3440);
  nand ginst10725 (P2_R1095_U268, P2_R1095_U179, P2_R1095_U267);
  nand ginst10726 (P2_R1095_U269, P2_R1095_U72, P2_U3068);
  nand ginst10727 (P2_R1095_U27, P2_R1095_U32, P2_U3069);
  not ginst10728 (P2_R1095_U270, P2_R1095_U178);
  nand ginst10729 (P2_R1095_U271, P2_R1095_U178, P2_U3081);
  not ginst10730 (P2_R1095_U272, P2_R1095_U176);
  nand ginst10731 (P2_R1095_U273, P2_R1095_U76, P2_U3445);
  nand ginst10732 (P2_R1095_U274, P2_R1095_U176, P2_R1095_U273);
  nand ginst10733 (P2_R1095_U275, P2_R1095_U75, P2_U3080);
  not ginst10734 (P2_R1095_U276, P2_R1095_U173);
  nand ginst10735 (P2_R1095_U277, P2_R1095_U78, P2_U3903);
  nand ginst10736 (P2_R1095_U278, P2_R1095_U173, P2_R1095_U277);
  nand ginst10737 (P2_R1095_U279, P2_R1095_U77, P2_U3075);
  not ginst10738 (P2_R1095_U28, P2_U3083);
  not ginst10739 (P2_R1095_U280, P2_R1095_U172);
  nand ginst10740 (P2_R1095_U281, P2_R1095_U82, P2_U3900);
  nand ginst10741 (P2_R1095_U282, P2_R1095_U79, P2_U3065);
  nand ginst10742 (P2_R1095_U283, P2_R1095_U80, P2_U3060);
  nand ginst10743 (P2_R1095_U284, P2_R1095_U10, P2_R1095_U200);
  nand ginst10744 (P2_R1095_U285, P2_R1095_U11, P2_R1095_U284);
  nand ginst10745 (P2_R1095_U286, P2_R1095_U84, P2_U3902);
  nand ginst10746 (P2_R1095_U287, P2_R1095_U82, P2_U3900);
  nand ginst10747 (P2_R1095_U288, P2_R1095_U133, P2_R1095_U172);
  nand ginst10748 (P2_R1095_U289, P2_R1095_U285, P2_R1095_U287);
  not ginst10749 (P2_R1095_U29, P2_U3404);
  not ginst10750 (P2_R1095_U290, P2_R1095_U169);
  nand ginst10751 (P2_R1095_U291, P2_R1095_U87, P2_U3899);
  nand ginst10752 (P2_R1095_U292, P2_R1095_U169, P2_R1095_U291);
  nand ginst10753 (P2_R1095_U293, P2_R1095_U86, P2_U3064);
  not ginst10754 (P2_R1095_U294, P2_R1095_U168);
  nand ginst10755 (P2_R1095_U295, P2_R1095_U89, P2_U3898);
  nand ginst10756 (P2_R1095_U296, P2_R1095_U168, P2_R1095_U295);
  nand ginst10757 (P2_R1095_U297, P2_R1095_U88, P2_U3057);
  not ginst10758 (P2_R1095_U298, P2_R1095_U93);
  nand ginst10759 (P2_R1095_U299, P2_R1095_U54, P2_U3896);
  not ginst10760 (P2_R1095_U30, P2_U3407);
  nand ginst10761 (P2_R1095_U300, P2_R1095_U53, P2_R1095_U54);
  nand ginst10762 (P2_R1095_U301, P2_R1095_U300, P2_R1095_U91);
  nand ginst10763 (P2_R1095_U302, P2_R1095_U189, P2_U3052);
  nand ginst10764 (P2_R1095_U303, P2_R1095_U92, P2_U3895);
  nand ginst10765 (P2_R1095_U304, P2_R1095_U51, P2_U3053);
  nand ginst10766 (P2_R1095_U305, P2_R1095_U140, P2_R1095_U355);
  nand ginst10767 (P2_R1095_U306, P2_R1095_U195, P2_R1095_U53);
  nand ginst10768 (P2_R1095_U307, P2_R1095_U172, P2_R1095_U286);
  not ginst10769 (P2_R1095_U308, P2_R1095_U94);
  nand ginst10770 (P2_R1095_U309, P2_R1095_U80, P2_U3060);
  not ginst10771 (P2_R1095_U31, P2_U3401);
  nand ginst10772 (P2_R1095_U310, P2_R1095_U308, P2_R1095_U309);
  nand ginst10773 (P2_R1095_U311, P2_R1095_U144, P2_R1095_U310);
  nand ginst10774 (P2_R1095_U312, P2_R1095_U194, P2_R1095_U94);
  nand ginst10775 (P2_R1095_U313, P2_R1095_U82, P2_U3900);
  nand ginst10776 (P2_R1095_U314, P2_R1095_U143, P2_R1095_U312);
  nand ginst10777 (P2_R1095_U315, P2_R1095_U80, P2_U3060);
  nand ginst10778 (P2_R1095_U316, P2_R1095_U194, P2_R1095_U315);
  nand ginst10779 (P2_R1095_U317, P2_R1095_U286, P2_R1095_U85);
  nand ginst10780 (P2_R1095_U318, P2_R1095_U182, P2_R1095_U262);
  not ginst10781 (P2_R1095_U319, P2_R1095_U95);
  not ginst10782 (P2_R1095_U32, P2_U3410);
  nand ginst10783 (P2_R1095_U320, P2_R1095_U66, P2_U3073);
  nand ginst10784 (P2_R1095_U321, P2_R1095_U319, P2_R1095_U320);
  nand ginst10785 (P2_R1095_U322, P2_R1095_U151, P2_R1095_U321);
  nand ginst10786 (P2_R1095_U323, P2_R1095_U193, P2_R1095_U95);
  nand ginst10787 (P2_R1095_U324, P2_R1095_U68, P2_U3437);
  nand ginst10788 (P2_R1095_U325, P2_R1095_U150, P2_R1095_U323);
  nand ginst10789 (P2_R1095_U326, P2_R1095_U66, P2_U3073);
  nand ginst10790 (P2_R1095_U327, P2_R1095_U193, P2_R1095_U326);
  nand ginst10791 (P2_R1095_U328, P2_R1095_U262, P2_R1095_U71);
  nand ginst10792 (P2_R1095_U329, P2_R1095_U58, P2_U3061);
  not ginst10793 (P2_R1095_U33, P2_U3413);
  nand ginst10794 (P2_R1095_U330, P2_R1095_U329, P2_R1095_U350);
  nand ginst10795 (P2_R1095_U331, P2_R1095_U155, P2_R1095_U330);
  nand ginst10796 (P2_R1095_U332, P2_R1095_U192, P2_R1095_U96);
  nand ginst10797 (P2_R1095_U333, P2_R1095_U56, P2_U3422);
  nand ginst10798 (P2_R1095_U334, P2_R1095_U154, P2_R1095_U332);
  nand ginst10799 (P2_R1095_U335, P2_R1095_U58, P2_U3061);
  nand ginst10800 (P2_R1095_U336, P2_R1095_U192, P2_R1095_U335);
  nand ginst10801 (P2_R1095_U337, P2_R1095_U38, P2_U3076);
  nand ginst10802 (P2_R1095_U338, P2_R1095_U174, P2_U3077);
  nand ginst10803 (P2_R1095_U339, P2_R1095_U177, P2_U3081);
  not ginst10804 (P2_R1095_U34, P2_U3067);
  nand ginst10805 (P2_R1095_U340, P2_R1095_U221, P2_R1095_U33);
  nand ginst10806 (P2_R1095_U341, P2_R1095_U121, P2_R1095_U161);
  nand ginst10807 (P2_R1095_U342, P2_R1095_U14, P2_R1095_U218);
  nand ginst10808 (P2_R1095_U343, P2_R1095_U250, P2_R1095_U251);
  nand ginst10809 (P2_R1095_U344, P2_R1095_U119, P2_R1095_U50);
  not ginst10810 (P2_R1095_U345, P2_R1095_U161);
  nand ginst10811 (P2_R1095_U346, P2_R1095_U196, P2_R1095_U50);
  nand ginst10812 (P2_R1095_U347, P2_R1095_U128, P2_R1095_U346);
  nand ginst10813 (P2_R1095_U348, P2_R1095_U205, P2_R1095_U35);
  nand ginst10814 (P2_R1095_U349, P2_R1095_U157, P2_R1095_U224);
  nand ginst10815 (P2_R1095_U35, P2_R1095_U37, P2_U3067);
  not ginst10816 (P2_R1095_U350, P2_R1095_U96);
  nand ginst10817 (P2_R1095_U351, P2_R1095_U15, P2_R1095_U157);
  not ginst10818 (P2_R1095_U352, P2_R1095_U184);
  nand ginst10819 (P2_R1095_U353, P2_R1095_U130, P2_R1095_U157);
  not ginst10820 (P2_R1095_U354, P2_R1095_U183);
  nand ginst10821 (P2_R1095_U355, P2_R1095_U298, P2_R1095_U53);
  nand ginst10822 (P2_R1095_U356, P2_R1095_U195, P2_R1095_U93);
  nand ginst10823 (P2_R1095_U357, P2_R1095_U139, P2_R1095_U356);
  nand ginst10824 (P2_R1095_U358, P2_R1095_U12, P2_R1095_U93);
  nand ginst10825 (P2_R1095_U359, P2_R1095_U136, P2_R1095_U358);
  not ginst10826 (P2_R1095_U36, P2_U3063);
  nand ginst10827 (P2_R1095_U360, P2_R1095_U12, P2_R1095_U93);
  not ginst10828 (P2_R1095_U361, P2_R1095_U166);
  nand ginst10829 (P2_R1095_U362, P2_R1095_U47, P2_U3416);
  nand ginst10830 (P2_R1095_U363, P2_R1095_U46, P2_U3082);
  nand ginst10831 (P2_R1095_U364, P2_R1095_U157, P2_R1095_U225);
  nand ginst10832 (P2_R1095_U365, P2_R1095_U156, P2_R1095_U223);
  nand ginst10833 (P2_R1095_U366, P2_R1095_U28, P2_U3413);
  nand ginst10834 (P2_R1095_U367, P2_R1095_U33, P2_U3083);
  nand ginst10835 (P2_R1095_U368, P2_R1095_U28, P2_U3413);
  nand ginst10836 (P2_R1095_U369, P2_R1095_U33, P2_U3083);
  not ginst10837 (P2_R1095_U37, P2_U3395);
  nand ginst10838 (P2_R1095_U370, P2_R1095_U368, P2_R1095_U369);
  nand ginst10839 (P2_R1095_U371, P2_R1095_U26, P2_U3410);
  nand ginst10840 (P2_R1095_U372, P2_R1095_U32, P2_U3069);
  nand ginst10841 (P2_R1095_U373, P2_R1095_U230, P2_R1095_U48);
  nand ginst10842 (P2_R1095_U374, P2_R1095_U158, P2_R1095_U219);
  nand ginst10843 (P2_R1095_U375, P2_R1095_U41, P2_U3407);
  nand ginst10844 (P2_R1095_U376, P2_R1095_U30, P2_U3070);
  nand ginst10845 (P2_R1095_U377, P2_R1095_U375, P2_R1095_U376);
  nand ginst10846 (P2_R1095_U378, P2_R1095_U42, P2_U3404);
  nand ginst10847 (P2_R1095_U379, P2_R1095_U29, P2_U3066);
  not ginst10848 (P2_R1095_U38, P2_U3387);
  nand ginst10849 (P2_R1095_U380, P2_R1095_U240, P2_R1095_U49);
  nand ginst10850 (P2_R1095_U381, P2_R1095_U159, P2_R1095_U232);
  nand ginst10851 (P2_R1095_U382, P2_R1095_U43, P2_U3401);
  nand ginst10852 (P2_R1095_U383, P2_R1095_U31, P2_U3059);
  nand ginst10853 (P2_R1095_U384, P2_R1095_U161, P2_R1095_U241);
  nand ginst10854 (P2_R1095_U385, P2_R1095_U160, P2_R1095_U345);
  nand ginst10855 (P2_R1095_U386, P2_R1095_U36, P2_U3398);
  nand ginst10856 (P2_R1095_U387, P2_R1095_U40, P2_U3063);
  nand ginst10857 (P2_R1095_U388, P2_R1095_U36, P2_U3398);
  nand ginst10858 (P2_R1095_U389, P2_R1095_U40, P2_U3063);
  not ginst10859 (P2_R1095_U39, P2_U3077);
  nand ginst10860 (P2_R1095_U390, P2_R1095_U388, P2_R1095_U389);
  nand ginst10861 (P2_R1095_U391, P2_R1095_U34, P2_U3395);
  nand ginst10862 (P2_R1095_U392, P2_R1095_U37, P2_U3067);
  nand ginst10863 (P2_R1095_U393, P2_R1095_U243, P2_R1095_U50);
  nand ginst10864 (P2_R1095_U394, P2_R1095_U162, P2_R1095_U205);
  nand ginst10865 (P2_R1095_U395, P2_R1095_U164, P2_U3904);
  nand ginst10866 (P2_R1095_U396, P2_R1095_U163, P2_U3054);
  nand ginst10867 (P2_R1095_U397, P2_R1095_U395, P2_R1095_U396);
  nand ginst10868 (P2_R1095_U398, P2_R1095_U164, P2_U3904);
  nand ginst10869 (P2_R1095_U399, P2_R1095_U163, P2_U3054);
  not ginst10870 (P2_R1095_U40, P2_U3398);
  nand ginst10871 (P2_R1095_U400, P2_R1095_U397, P2_R1095_U51, P2_U3053);
  nand ginst10872 (P2_R1095_U401, P2_R1095_U16, P2_R1095_U92, P2_U3895);
  nand ginst10873 (P2_R1095_U402, P2_R1095_U92, P2_U3895);
  nand ginst10874 (P2_R1095_U403, P2_R1095_U51, P2_U3053);
  not ginst10875 (P2_R1095_U404, P2_R1095_U138);
  nand ginst10876 (P2_R1095_U405, P2_R1095_U361, P2_R1095_U404);
  nand ginst10877 (P2_R1095_U406, P2_R1095_U138, P2_R1095_U166);
  nand ginst10878 (P2_R1095_U407, P2_R1095_U54, P2_U3896);
  nand ginst10879 (P2_R1095_U408, P2_R1095_U91, P2_U3052);
  nand ginst10880 (P2_R1095_U409, P2_R1095_U54, P2_U3896);
  not ginst10881 (P2_R1095_U41, P2_U3070);
  nand ginst10882 (P2_R1095_U410, P2_R1095_U91, P2_U3052);
  nand ginst10883 (P2_R1095_U411, P2_R1095_U409, P2_R1095_U410);
  nand ginst10884 (P2_R1095_U412, P2_R1095_U52, P2_U3897);
  nand ginst10885 (P2_R1095_U413, P2_R1095_U90, P2_U3056);
  nand ginst10886 (P2_R1095_U414, P2_R1095_U306, P2_R1095_U93);
  nand ginst10887 (P2_R1095_U415, P2_R1095_U167, P2_R1095_U298);
  nand ginst10888 (P2_R1095_U416, P2_R1095_U89, P2_U3898);
  nand ginst10889 (P2_R1095_U417, P2_R1095_U88, P2_U3057);
  not ginst10890 (P2_R1095_U418, P2_R1095_U141);
  nand ginst10891 (P2_R1095_U419, P2_R1095_U294, P2_R1095_U418);
  not ginst10892 (P2_R1095_U42, P2_U3066);
  nand ginst10893 (P2_R1095_U420, P2_R1095_U141, P2_R1095_U168);
  nand ginst10894 (P2_R1095_U421, P2_R1095_U87, P2_U3899);
  nand ginst10895 (P2_R1095_U422, P2_R1095_U86, P2_U3064);
  not ginst10896 (P2_R1095_U423, P2_R1095_U142);
  nand ginst10897 (P2_R1095_U424, P2_R1095_U290, P2_R1095_U423);
  nand ginst10898 (P2_R1095_U425, P2_R1095_U142, P2_R1095_U169);
  nand ginst10899 (P2_R1095_U426, P2_R1095_U82, P2_U3900);
  nand ginst10900 (P2_R1095_U427, P2_R1095_U79, P2_U3065);
  nand ginst10901 (P2_R1095_U428, P2_R1095_U426, P2_R1095_U427);
  nand ginst10902 (P2_R1095_U429, P2_R1095_U83, P2_U3901);
  not ginst10903 (P2_R1095_U43, P2_U3059);
  nand ginst10904 (P2_R1095_U430, P2_R1095_U80, P2_U3060);
  nand ginst10905 (P2_R1095_U431, P2_R1095_U316, P2_R1095_U94);
  nand ginst10906 (P2_R1095_U432, P2_R1095_U170, P2_R1095_U308);
  nand ginst10907 (P2_R1095_U433, P2_R1095_U84, P2_U3902);
  nand ginst10908 (P2_R1095_U434, P2_R1095_U81, P2_U3074);
  nand ginst10909 (P2_R1095_U435, P2_R1095_U172, P2_R1095_U317);
  nand ginst10910 (P2_R1095_U436, P2_R1095_U171, P2_R1095_U280);
  nand ginst10911 (P2_R1095_U437, P2_R1095_U78, P2_U3903);
  nand ginst10912 (P2_R1095_U438, P2_R1095_U77, P2_U3075);
  not ginst10913 (P2_R1095_U439, P2_R1095_U145);
  nand ginst10914 (P2_R1095_U44, P2_R1095_U31, P2_U3059);
  nand ginst10915 (P2_R1095_U440, P2_R1095_U276, P2_R1095_U439);
  nand ginst10916 (P2_R1095_U441, P2_R1095_U145, P2_R1095_U173);
  nand ginst10917 (P2_R1095_U442, P2_R1095_U39, P2_U3392);
  nand ginst10918 (P2_R1095_U443, P2_R1095_U174, P2_U3077);
  not ginst10919 (P2_R1095_U444, P2_R1095_U146);
  nand ginst10920 (P2_R1095_U445, P2_R1095_U203, P2_R1095_U444);
  nand ginst10921 (P2_R1095_U446, P2_R1095_U146, P2_R1095_U175);
  nand ginst10922 (P2_R1095_U447, P2_R1095_U76, P2_U3445);
  nand ginst10923 (P2_R1095_U448, P2_R1095_U75, P2_U3080);
  not ginst10924 (P2_R1095_U449, P2_R1095_U147);
  nand ginst10925 (P2_R1095_U45, P2_R1095_U214, P2_R1095_U216);
  nand ginst10926 (P2_R1095_U450, P2_R1095_U272, P2_R1095_U449);
  nand ginst10927 (P2_R1095_U451, P2_R1095_U147, P2_R1095_U176);
  nand ginst10928 (P2_R1095_U452, P2_R1095_U74, P2_U3443);
  nand ginst10929 (P2_R1095_U453, P2_R1095_U177, P2_U3081);
  not ginst10930 (P2_R1095_U454, P2_R1095_U148);
  nand ginst10931 (P2_R1095_U455, P2_R1095_U270, P2_R1095_U454);
  nand ginst10932 (P2_R1095_U456, P2_R1095_U148, P2_R1095_U178);
  nand ginst10933 (P2_R1095_U457, P2_R1095_U73, P2_U3440);
  nand ginst10934 (P2_R1095_U458, P2_R1095_U72, P2_U3068);
  not ginst10935 (P2_R1095_U459, P2_R1095_U149);
  not ginst10936 (P2_R1095_U46, P2_U3416);
  nand ginst10937 (P2_R1095_U460, P2_R1095_U266, P2_R1095_U459);
  nand ginst10938 (P2_R1095_U461, P2_R1095_U149, P2_R1095_U179);
  nand ginst10939 (P2_R1095_U462, P2_R1095_U68, P2_U3437);
  nand ginst10940 (P2_R1095_U463, P2_R1095_U65, P2_U3072);
  nand ginst10941 (P2_R1095_U464, P2_R1095_U462, P2_R1095_U463);
  nand ginst10942 (P2_R1095_U465, P2_R1095_U69, P2_U3434);
  nand ginst10943 (P2_R1095_U466, P2_R1095_U66, P2_U3073);
  nand ginst10944 (P2_R1095_U467, P2_R1095_U327, P2_R1095_U95);
  nand ginst10945 (P2_R1095_U468, P2_R1095_U180, P2_R1095_U319);
  nand ginst10946 (P2_R1095_U469, P2_R1095_U70, P2_U3431);
  not ginst10947 (P2_R1095_U47, P2_U3082);
  nand ginst10948 (P2_R1095_U470, P2_R1095_U67, P2_U3078);
  nand ginst10949 (P2_R1095_U471, P2_R1095_U182, P2_R1095_U328);
  nand ginst10950 (P2_R1095_U472, P2_R1095_U181, P2_R1095_U256);
  nand ginst10951 (P2_R1095_U473, P2_R1095_U64, P2_U3428);
  nand ginst10952 (P2_R1095_U474, P2_R1095_U63, P2_U3079);
  not ginst10953 (P2_R1095_U475, P2_R1095_U152);
  nand ginst10954 (P2_R1095_U476, P2_R1095_U354, P2_R1095_U475);
  nand ginst10955 (P2_R1095_U477, P2_R1095_U152, P2_R1095_U183);
  nand ginst10956 (P2_R1095_U478, P2_R1095_U55, P2_U3425);
  nand ginst10957 (P2_R1095_U479, P2_R1095_U61, P2_U3071);
  nand ginst10958 (P2_R1095_U48, P2_R1095_U217, P2_R1095_U45);
  not ginst10959 (P2_R1095_U480, P2_R1095_U153);
  nand ginst10960 (P2_R1095_U481, P2_R1095_U352, P2_R1095_U480);
  nand ginst10961 (P2_R1095_U482, P2_R1095_U153, P2_R1095_U184);
  nand ginst10962 (P2_R1095_U483, P2_R1095_U56, P2_U3422);
  nand ginst10963 (P2_R1095_U484, P2_R1095_U60, P2_U3062);
  nand ginst10964 (P2_R1095_U485, P2_R1095_U483, P2_R1095_U484);
  nand ginst10965 (P2_R1095_U486, P2_R1095_U57, P2_U3419);
  nand ginst10966 (P2_R1095_U487, P2_R1095_U58, P2_U3061);
  nand ginst10967 (P2_R1095_U488, P2_R1095_U336, P2_R1095_U96);
  nand ginst10968 (P2_R1095_U489, P2_R1095_U185, P2_R1095_U350);
  nand ginst10969 (P2_R1095_U49, P2_R1095_U231, P2_R1095_U44);
  nand ginst10970 (P2_R1095_U50, P2_R1095_U188, P2_R1095_U204, P2_R1095_U338);
  not ginst10971 (P2_R1095_U51, P2_U3895);
  not ginst10972 (P2_R1095_U52, P2_U3056);
  nand ginst10973 (P2_R1095_U53, P2_R1095_U90, P2_U3056);
  not ginst10974 (P2_R1095_U54, P2_U3052);
  not ginst10975 (P2_R1095_U55, P2_U3071);
  not ginst10976 (P2_R1095_U56, P2_U3062);
  not ginst10977 (P2_R1095_U57, P2_U3061);
  not ginst10978 (P2_R1095_U58, P2_U3419);
  nand ginst10979 (P2_R1095_U59, P2_R1095_U46, P2_U3082);
  and ginst10980 (P2_R1095_U6, P2_R1095_U211, P2_R1095_U212);
  not ginst10981 (P2_R1095_U60, P2_U3422);
  not ginst10982 (P2_R1095_U61, P2_U3425);
  nand ginst10983 (P2_R1095_U62, P2_R1095_U248, P2_R1095_U249);
  not ginst10984 (P2_R1095_U63, P2_U3428);
  not ginst10985 (P2_R1095_U64, P2_U3079);
  not ginst10986 (P2_R1095_U65, P2_U3437);
  not ginst10987 (P2_R1095_U66, P2_U3434);
  not ginst10988 (P2_R1095_U67, P2_U3431);
  not ginst10989 (P2_R1095_U68, P2_U3072);
  not ginst10990 (P2_R1095_U69, P2_U3073);
  and ginst10991 (P2_R1095_U7, P2_R1095_U245, P2_R1095_U246);
  not ginst10992 (P2_R1095_U70, P2_U3078);
  nand ginst10993 (P2_R1095_U71, P2_R1095_U67, P2_U3078);
  not ginst10994 (P2_R1095_U72, P2_U3440);
  not ginst10995 (P2_R1095_U73, P2_U3068);
  not ginst10996 (P2_R1095_U74, P2_U3081);
  not ginst10997 (P2_R1095_U75, P2_U3445);
  not ginst10998 (P2_R1095_U76, P2_U3080);
  not ginst10999 (P2_R1095_U77, P2_U3903);
  not ginst11000 (P2_R1095_U78, P2_U3075);
  not ginst11001 (P2_R1095_U79, P2_U3900);
  and ginst11002 (P2_R1095_U8, P2_R1095_U193, P2_R1095_U257);
  not ginst11003 (P2_R1095_U80, P2_U3901);
  not ginst11004 (P2_R1095_U81, P2_U3902);
  not ginst11005 (P2_R1095_U82, P2_U3065);
  not ginst11006 (P2_R1095_U83, P2_U3060);
  not ginst11007 (P2_R1095_U84, P2_U3074);
  nand ginst11008 (P2_R1095_U85, P2_R1095_U81, P2_U3074);
  not ginst11009 (P2_R1095_U86, P2_U3899);
  not ginst11010 (P2_R1095_U87, P2_U3064);
  not ginst11011 (P2_R1095_U88, P2_U3898);
  not ginst11012 (P2_R1095_U89, P2_U3057);
  and ginst11013 (P2_R1095_U9, P2_R1095_U258, P2_R1095_U259);
  not ginst11014 (P2_R1095_U90, P2_U3897);
  not ginst11015 (P2_R1095_U91, P2_U3896);
  not ginst11016 (P2_R1095_U92, P2_U3053);
  nand ginst11017 (P2_R1095_U93, P2_R1095_U296, P2_R1095_U297);
  nand ginst11018 (P2_R1095_U94, P2_R1095_U307, P2_R1095_U85);
  nand ginst11019 (P2_R1095_U95, P2_R1095_U318, P2_R1095_U71);
  nand ginst11020 (P2_R1095_U96, P2_R1095_U349, P2_R1095_U59);
  not ginst11021 (P2_R1095_U97, P2_U3076);
  nand ginst11022 (P2_R1095_U98, P2_R1095_U405, P2_R1095_U406);
  nand ginst11023 (P2_R1095_U99, P2_R1095_U419, P2_R1095_U420);
  and ginst11024 (P2_R1110_U10, P2_R1110_U348, P2_R1110_U351);
  nand ginst11025 (P2_R1110_U100, P2_R1110_U398, P2_R1110_U399);
  nand ginst11026 (P2_R1110_U101, P2_R1110_U407, P2_R1110_U408);
  nand ginst11027 (P2_R1110_U102, P2_R1110_U414, P2_R1110_U415);
  nand ginst11028 (P2_R1110_U103, P2_R1110_U421, P2_R1110_U422);
  nand ginst11029 (P2_R1110_U104, P2_R1110_U428, P2_R1110_U429);
  nand ginst11030 (P2_R1110_U105, P2_R1110_U433, P2_R1110_U434);
  nand ginst11031 (P2_R1110_U106, P2_R1110_U440, P2_R1110_U441);
  nand ginst11032 (P2_R1110_U107, P2_R1110_U447, P2_R1110_U448);
  nand ginst11033 (P2_R1110_U108, P2_R1110_U461, P2_R1110_U462);
  nand ginst11034 (P2_R1110_U109, P2_R1110_U466, P2_R1110_U467);
  and ginst11035 (P2_R1110_U11, P2_R1110_U341, P2_R1110_U344);
  nand ginst11036 (P2_R1110_U110, P2_R1110_U473, P2_R1110_U474);
  nand ginst11037 (P2_R1110_U111, P2_R1110_U480, P2_R1110_U481);
  nand ginst11038 (P2_R1110_U112, P2_R1110_U487, P2_R1110_U488);
  nand ginst11039 (P2_R1110_U113, P2_R1110_U494, P2_R1110_U495);
  nand ginst11040 (P2_R1110_U114, P2_R1110_U499, P2_R1110_U500);
  and ginst11041 (P2_R1110_U115, P2_R1110_U187, P2_R1110_U189);
  and ginst11042 (P2_R1110_U116, P2_R1110_U180, P2_R1110_U4);
  and ginst11043 (P2_R1110_U117, P2_R1110_U192, P2_R1110_U194);
  and ginst11044 (P2_R1110_U118, P2_R1110_U200, P2_R1110_U201);
  and ginst11045 (P2_R1110_U119, P2_R1110_U22, P2_R1110_U381, P2_R1110_U382);
  and ginst11046 (P2_R1110_U12, P2_R1110_U332, P2_R1110_U335);
  and ginst11047 (P2_R1110_U120, P2_R1110_U212, P2_R1110_U5);
  and ginst11048 (P2_R1110_U121, P2_R1110_U180, P2_R1110_U181);
  and ginst11049 (P2_R1110_U122, P2_R1110_U218, P2_R1110_U220);
  and ginst11050 (P2_R1110_U123, P2_R1110_U34, P2_R1110_U388, P2_R1110_U389);
  and ginst11051 (P2_R1110_U124, P2_R1110_U226, P2_R1110_U4);
  and ginst11052 (P2_R1110_U125, P2_R1110_U181, P2_R1110_U234);
  and ginst11053 (P2_R1110_U126, P2_R1110_U204, P2_R1110_U6);
  and ginst11054 (P2_R1110_U127, P2_R1110_U239, P2_R1110_U243);
  and ginst11055 (P2_R1110_U128, P2_R1110_U250, P2_R1110_U7);
  and ginst11056 (P2_R1110_U129, P2_R1110_U248, P2_R1110_U253);
  and ginst11057 (P2_R1110_U13, P2_R1110_U323, P2_R1110_U326);
  and ginst11058 (P2_R1110_U130, P2_R1110_U267, P2_R1110_U268);
  and ginst11059 (P2_R1110_U131, P2_R1110_U282, P2_R1110_U9);
  and ginst11060 (P2_R1110_U132, P2_R1110_U280, P2_R1110_U285);
  and ginst11061 (P2_R1110_U133, P2_R1110_U298, P2_R1110_U301);
  and ginst11062 (P2_R1110_U134, P2_R1110_U302, P2_R1110_U368);
  and ginst11063 (P2_R1110_U135, P2_R1110_U160, P2_R1110_U278);
  and ginst11064 (P2_R1110_U136, P2_R1110_U454, P2_R1110_U455, P2_R1110_U80);
  and ginst11065 (P2_R1110_U137, P2_R1110_U325, P2_R1110_U9);
  and ginst11066 (P2_R1110_U138, P2_R1110_U468, P2_R1110_U469, P2_R1110_U59);
  and ginst11067 (P2_R1110_U139, P2_R1110_U334, P2_R1110_U8);
  and ginst11068 (P2_R1110_U14, P2_R1110_U318, P2_R1110_U320);
  and ginst11069 (P2_R1110_U140, P2_R1110_U172, P2_R1110_U489, P2_R1110_U490);
  and ginst11070 (P2_R1110_U141, P2_R1110_U343, P2_R1110_U7);
  and ginst11071 (P2_R1110_U142, P2_R1110_U171, P2_R1110_U501, P2_R1110_U502);
  and ginst11072 (P2_R1110_U143, P2_R1110_U350, P2_R1110_U6);
  nand ginst11073 (P2_R1110_U144, P2_R1110_U118, P2_R1110_U202);
  nand ginst11074 (P2_R1110_U145, P2_R1110_U217, P2_R1110_U229);
  not ginst11075 (P2_R1110_U146, P2_U3054);
  not ginst11076 (P2_R1110_U147, P2_U3904);
  and ginst11077 (P2_R1110_U148, P2_R1110_U402, P2_R1110_U403);
  nand ginst11078 (P2_R1110_U149, P2_R1110_U169, P2_R1110_U304, P2_R1110_U364);
  and ginst11079 (P2_R1110_U15, P2_R1110_U310, P2_R1110_U313);
  and ginst11080 (P2_R1110_U150, P2_R1110_U409, P2_R1110_U410);
  nand ginst11081 (P2_R1110_U151, P2_R1110_U134, P2_R1110_U369, P2_R1110_U370);
  and ginst11082 (P2_R1110_U152, P2_R1110_U416, P2_R1110_U417);
  nand ginst11083 (P2_R1110_U153, P2_R1110_U299, P2_R1110_U365, P2_R1110_U86);
  and ginst11084 (P2_R1110_U154, P2_R1110_U423, P2_R1110_U424);
  nand ginst11085 (P2_R1110_U155, P2_R1110_U292, P2_R1110_U293);
  and ginst11086 (P2_R1110_U156, P2_R1110_U435, P2_R1110_U436);
  nand ginst11087 (P2_R1110_U157, P2_R1110_U288, P2_R1110_U289);
  and ginst11088 (P2_R1110_U158, P2_R1110_U442, P2_R1110_U443);
  nand ginst11089 (P2_R1110_U159, P2_R1110_U132, P2_R1110_U284);
  and ginst11090 (P2_R1110_U16, P2_R1110_U232, P2_R1110_U235);
  and ginst11091 (P2_R1110_U160, P2_R1110_U449, P2_R1110_U450);
  nand ginst11092 (P2_R1110_U161, P2_R1110_U327, P2_R1110_U43);
  nand ginst11093 (P2_R1110_U162, P2_R1110_U130, P2_R1110_U269);
  and ginst11094 (P2_R1110_U163, P2_R1110_U475, P2_R1110_U476);
  nand ginst11095 (P2_R1110_U164, P2_R1110_U256, P2_R1110_U257);
  and ginst11096 (P2_R1110_U165, P2_R1110_U482, P2_R1110_U483);
  nand ginst11097 (P2_R1110_U166, P2_R1110_U129, P2_R1110_U252);
  nand ginst11098 (P2_R1110_U167, P2_R1110_U127, P2_R1110_U242);
  nand ginst11099 (P2_R1110_U168, P2_R1110_U366, P2_R1110_U367);
  nand ginst11100 (P2_R1110_U169, P2_R1110_U151, P2_U3053);
  and ginst11101 (P2_R1110_U17, P2_R1110_U224, P2_R1110_U227);
  not ginst11102 (P2_R1110_U170, P2_R1110_U34);
  nand ginst11103 (P2_R1110_U171, P2_U3082, P2_U3416);
  nand ginst11104 (P2_R1110_U172, P2_U3071, P2_U3425);
  nand ginst11105 (P2_R1110_U173, P2_U3057, P2_U3898);
  not ginst11106 (P2_R1110_U174, P2_R1110_U68);
  not ginst11107 (P2_R1110_U175, P2_R1110_U77);
  nand ginst11108 (P2_R1110_U176, P2_U3064, P2_U3899);
  not ginst11109 (P2_R1110_U177, P2_R1110_U65);
  or ginst11110 (P2_R1110_U178, P2_U3066, P2_U3404);
  or ginst11111 (P2_R1110_U179, P2_U3059, P2_U3401);
  and ginst11112 (P2_R1110_U18, P2_R1110_U210, P2_R1110_U213);
  or ginst11113 (P2_R1110_U180, P2_U3063, P2_U3398);
  or ginst11114 (P2_R1110_U181, P2_U3067, P2_U3395);
  not ginst11115 (P2_R1110_U182, P2_R1110_U31);
  or ginst11116 (P2_R1110_U183, P2_U3077, P2_U3392);
  not ginst11117 (P2_R1110_U184, P2_R1110_U42);
  not ginst11118 (P2_R1110_U185, P2_R1110_U43);
  nand ginst11119 (P2_R1110_U186, P2_R1110_U42, P2_R1110_U43);
  nand ginst11120 (P2_R1110_U187, P2_U3067, P2_U3395);
  nand ginst11121 (P2_R1110_U188, P2_R1110_U181, P2_R1110_U186);
  nand ginst11122 (P2_R1110_U189, P2_U3063, P2_U3398);
  not ginst11123 (P2_R1110_U19, P2_U3407);
  nand ginst11124 (P2_R1110_U190, P2_R1110_U115, P2_R1110_U188);
  nand ginst11125 (P2_R1110_U191, P2_R1110_U34, P2_R1110_U35);
  nand ginst11126 (P2_R1110_U192, P2_R1110_U191, P2_U3066);
  nand ginst11127 (P2_R1110_U193, P2_R1110_U116, P2_R1110_U190);
  nand ginst11128 (P2_R1110_U194, P2_R1110_U170, P2_U3404);
  not ginst11129 (P2_R1110_U195, P2_R1110_U41);
  or ginst11130 (P2_R1110_U196, P2_U3069, P2_U3410);
  or ginst11131 (P2_R1110_U197, P2_U3070, P2_U3407);
  not ginst11132 (P2_R1110_U198, P2_R1110_U22);
  nand ginst11133 (P2_R1110_U199, P2_R1110_U22, P2_R1110_U23);
  not ginst11134 (P2_R1110_U20, P2_U3070);
  nand ginst11135 (P2_R1110_U200, P2_R1110_U199, P2_U3069);
  nand ginst11136 (P2_R1110_U201, P2_R1110_U198, P2_U3410);
  nand ginst11137 (P2_R1110_U202, P2_R1110_U41, P2_R1110_U5);
  not ginst11138 (P2_R1110_U203, P2_R1110_U144);
  or ginst11139 (P2_R1110_U204, P2_U3083, P2_U3413);
  nand ginst11140 (P2_R1110_U205, P2_R1110_U144, P2_R1110_U204);
  not ginst11141 (P2_R1110_U206, P2_R1110_U40);
  or ginst11142 (P2_R1110_U207, P2_U3082, P2_U3416);
  or ginst11143 (P2_R1110_U208, P2_U3070, P2_U3407);
  nand ginst11144 (P2_R1110_U209, P2_R1110_U208, P2_R1110_U41);
  not ginst11145 (P2_R1110_U21, P2_U3069);
  nand ginst11146 (P2_R1110_U210, P2_R1110_U119, P2_R1110_U209);
  nand ginst11147 (P2_R1110_U211, P2_R1110_U195, P2_R1110_U22);
  nand ginst11148 (P2_R1110_U212, P2_U3069, P2_U3410);
  nand ginst11149 (P2_R1110_U213, P2_R1110_U120, P2_R1110_U211);
  or ginst11150 (P2_R1110_U214, P2_U3070, P2_U3407);
  nand ginst11151 (P2_R1110_U215, P2_R1110_U181, P2_R1110_U185);
  nand ginst11152 (P2_R1110_U216, P2_U3067, P2_U3395);
  not ginst11153 (P2_R1110_U217, P2_R1110_U45);
  nand ginst11154 (P2_R1110_U218, P2_R1110_U121, P2_R1110_U184);
  nand ginst11155 (P2_R1110_U219, P2_R1110_U180, P2_R1110_U45);
  nand ginst11156 (P2_R1110_U22, P2_U3070, P2_U3407);
  nand ginst11157 (P2_R1110_U220, P2_U3063, P2_U3398);
  not ginst11158 (P2_R1110_U221, P2_R1110_U44);
  or ginst11159 (P2_R1110_U222, P2_U3059, P2_U3401);
  nand ginst11160 (P2_R1110_U223, P2_R1110_U222, P2_R1110_U44);
  nand ginst11161 (P2_R1110_U224, P2_R1110_U123, P2_R1110_U223);
  nand ginst11162 (P2_R1110_U225, P2_R1110_U221, P2_R1110_U34);
  nand ginst11163 (P2_R1110_U226, P2_U3066, P2_U3404);
  nand ginst11164 (P2_R1110_U227, P2_R1110_U124, P2_R1110_U225);
  or ginst11165 (P2_R1110_U228, P2_U3059, P2_U3401);
  nand ginst11166 (P2_R1110_U229, P2_R1110_U181, P2_R1110_U184);
  not ginst11167 (P2_R1110_U23, P2_U3410);
  not ginst11168 (P2_R1110_U230, P2_R1110_U145);
  nand ginst11169 (P2_R1110_U231, P2_U3063, P2_U3398);
  nand ginst11170 (P2_R1110_U232, P2_R1110_U400, P2_R1110_U401, P2_R1110_U42, P2_R1110_U43);
  nand ginst11171 (P2_R1110_U233, P2_R1110_U42, P2_R1110_U43);
  nand ginst11172 (P2_R1110_U234, P2_U3067, P2_U3395);
  nand ginst11173 (P2_R1110_U235, P2_R1110_U125, P2_R1110_U233);
  or ginst11174 (P2_R1110_U236, P2_U3082, P2_U3416);
  or ginst11175 (P2_R1110_U237, P2_U3061, P2_U3419);
  nand ginst11176 (P2_R1110_U238, P2_R1110_U177, P2_R1110_U6);
  nand ginst11177 (P2_R1110_U239, P2_U3061, P2_U3419);
  not ginst11178 (P2_R1110_U24, P2_U3401);
  nand ginst11179 (P2_R1110_U240, P2_R1110_U171, P2_R1110_U238);
  or ginst11180 (P2_R1110_U241, P2_U3061, P2_U3419);
  nand ginst11181 (P2_R1110_U242, P2_R1110_U126, P2_R1110_U144);
  nand ginst11182 (P2_R1110_U243, P2_R1110_U240, P2_R1110_U241);
  not ginst11183 (P2_R1110_U244, P2_R1110_U167);
  or ginst11184 (P2_R1110_U245, P2_U3079, P2_U3428);
  or ginst11185 (P2_R1110_U246, P2_U3071, P2_U3425);
  nand ginst11186 (P2_R1110_U247, P2_R1110_U174, P2_R1110_U7);
  nand ginst11187 (P2_R1110_U248, P2_U3079, P2_U3428);
  nand ginst11188 (P2_R1110_U249, P2_R1110_U172, P2_R1110_U247);
  not ginst11189 (P2_R1110_U25, P2_U3059);
  or ginst11190 (P2_R1110_U250, P2_U3062, P2_U3422);
  or ginst11191 (P2_R1110_U251, P2_U3079, P2_U3428);
  nand ginst11192 (P2_R1110_U252, P2_R1110_U128, P2_R1110_U167);
  nand ginst11193 (P2_R1110_U253, P2_R1110_U249, P2_R1110_U251);
  not ginst11194 (P2_R1110_U254, P2_R1110_U166);
  or ginst11195 (P2_R1110_U255, P2_U3078, P2_U3431);
  nand ginst11196 (P2_R1110_U256, P2_R1110_U166, P2_R1110_U255);
  nand ginst11197 (P2_R1110_U257, P2_U3078, P2_U3431);
  not ginst11198 (P2_R1110_U258, P2_R1110_U164);
  or ginst11199 (P2_R1110_U259, P2_U3073, P2_U3434);
  not ginst11200 (P2_R1110_U26, P2_U3066);
  nand ginst11201 (P2_R1110_U260, P2_R1110_U164, P2_R1110_U259);
  nand ginst11202 (P2_R1110_U261, P2_U3073, P2_U3434);
  not ginst11203 (P2_R1110_U262, P2_R1110_U92);
  or ginst11204 (P2_R1110_U263, P2_U3068, P2_U3440);
  or ginst11205 (P2_R1110_U264, P2_U3072, P2_U3437);
  not ginst11206 (P2_R1110_U265, P2_R1110_U59);
  nand ginst11207 (P2_R1110_U266, P2_R1110_U59, P2_R1110_U60);
  nand ginst11208 (P2_R1110_U267, P2_R1110_U266, P2_U3068);
  nand ginst11209 (P2_R1110_U268, P2_R1110_U265, P2_U3440);
  nand ginst11210 (P2_R1110_U269, P2_R1110_U8, P2_R1110_U92);
  not ginst11211 (P2_R1110_U27, P2_U3395);
  not ginst11212 (P2_R1110_U270, P2_R1110_U162);
  or ginst11213 (P2_R1110_U271, P2_U3075, P2_U3903);
  or ginst11214 (P2_R1110_U272, P2_U3080, P2_U3445);
  or ginst11215 (P2_R1110_U273, P2_U3074, P2_U3902);
  not ginst11216 (P2_R1110_U274, P2_R1110_U80);
  nand ginst11217 (P2_R1110_U275, P2_R1110_U274, P2_U3903);
  nand ginst11218 (P2_R1110_U276, P2_R1110_U275, P2_R1110_U90);
  nand ginst11219 (P2_R1110_U277, P2_R1110_U80, P2_R1110_U81);
  nand ginst11220 (P2_R1110_U278, P2_R1110_U276, P2_R1110_U277);
  nand ginst11221 (P2_R1110_U279, P2_R1110_U175, P2_R1110_U9);
  not ginst11222 (P2_R1110_U28, P2_U3067);
  nand ginst11223 (P2_R1110_U280, P2_U3074, P2_U3902);
  nand ginst11224 (P2_R1110_U281, P2_R1110_U278, P2_R1110_U279);
  or ginst11225 (P2_R1110_U282, P2_U3081, P2_U3443);
  or ginst11226 (P2_R1110_U283, P2_U3074, P2_U3902);
  nand ginst11227 (P2_R1110_U284, P2_R1110_U131, P2_R1110_U162, P2_R1110_U273);
  nand ginst11228 (P2_R1110_U285, P2_R1110_U281, P2_R1110_U283);
  not ginst11229 (P2_R1110_U286, P2_R1110_U159);
  or ginst11230 (P2_R1110_U287, P2_U3060, P2_U3901);
  nand ginst11231 (P2_R1110_U288, P2_R1110_U159, P2_R1110_U287);
  nand ginst11232 (P2_R1110_U289, P2_U3060, P2_U3901);
  not ginst11233 (P2_R1110_U29, P2_U3387);
  not ginst11234 (P2_R1110_U290, P2_R1110_U157);
  or ginst11235 (P2_R1110_U291, P2_U3065, P2_U3900);
  nand ginst11236 (P2_R1110_U292, P2_R1110_U157, P2_R1110_U291);
  nand ginst11237 (P2_R1110_U293, P2_U3065, P2_U3900);
  not ginst11238 (P2_R1110_U294, P2_R1110_U155);
  or ginst11239 (P2_R1110_U295, P2_U3057, P2_U3898);
  nand ginst11240 (P2_R1110_U296, P2_R1110_U173, P2_R1110_U176);
  not ginst11241 (P2_R1110_U297, P2_R1110_U86);
  or ginst11242 (P2_R1110_U298, P2_U3064, P2_U3899);
  nand ginst11243 (P2_R1110_U299, P2_R1110_U155, P2_R1110_U168, P2_R1110_U298);
  not ginst11244 (P2_R1110_U30, P2_U3076);
  not ginst11245 (P2_R1110_U300, P2_R1110_U153);
  or ginst11246 (P2_R1110_U301, P2_U3052, P2_U3896);
  nand ginst11247 (P2_R1110_U302, P2_U3052, P2_U3896);
  not ginst11248 (P2_R1110_U303, P2_R1110_U151);
  nand ginst11249 (P2_R1110_U304, P2_R1110_U151, P2_U3895);
  not ginst11250 (P2_R1110_U305, P2_R1110_U149);
  nand ginst11251 (P2_R1110_U306, P2_R1110_U155, P2_R1110_U298);
  not ginst11252 (P2_R1110_U307, P2_R1110_U89);
  or ginst11253 (P2_R1110_U308, P2_U3057, P2_U3898);
  nand ginst11254 (P2_R1110_U309, P2_R1110_U308, P2_R1110_U89);
  nand ginst11255 (P2_R1110_U31, P2_U3076, P2_U3387);
  nand ginst11256 (P2_R1110_U310, P2_R1110_U154, P2_R1110_U173, P2_R1110_U309);
  nand ginst11257 (P2_R1110_U311, P2_R1110_U173, P2_R1110_U307);
  nand ginst11258 (P2_R1110_U312, P2_U3056, P2_U3897);
  nand ginst11259 (P2_R1110_U313, P2_R1110_U168, P2_R1110_U311, P2_R1110_U312);
  or ginst11260 (P2_R1110_U314, P2_U3057, P2_U3898);
  nand ginst11261 (P2_R1110_U315, P2_R1110_U162, P2_R1110_U282);
  not ginst11262 (P2_R1110_U316, P2_R1110_U91);
  nand ginst11263 (P2_R1110_U317, P2_R1110_U9, P2_R1110_U91);
  nand ginst11264 (P2_R1110_U318, P2_R1110_U135, P2_R1110_U317);
  nand ginst11265 (P2_R1110_U319, P2_R1110_U278, P2_R1110_U317);
  not ginst11266 (P2_R1110_U32, P2_U3398);
  nand ginst11267 (P2_R1110_U320, P2_R1110_U319, P2_R1110_U453);
  or ginst11268 (P2_R1110_U321, P2_U3080, P2_U3445);
  nand ginst11269 (P2_R1110_U322, P2_R1110_U321, P2_R1110_U91);
  nand ginst11270 (P2_R1110_U323, P2_R1110_U136, P2_R1110_U322);
  nand ginst11271 (P2_R1110_U324, P2_R1110_U316, P2_R1110_U80);
  nand ginst11272 (P2_R1110_U325, P2_U3075, P2_U3903);
  nand ginst11273 (P2_R1110_U326, P2_R1110_U137, P2_R1110_U324);
  or ginst11274 (P2_R1110_U327, P2_U3077, P2_U3392);
  not ginst11275 (P2_R1110_U328, P2_R1110_U161);
  or ginst11276 (P2_R1110_U329, P2_U3080, P2_U3445);
  not ginst11277 (P2_R1110_U33, P2_U3063);
  or ginst11278 (P2_R1110_U330, P2_U3072, P2_U3437);
  nand ginst11279 (P2_R1110_U331, P2_R1110_U330, P2_R1110_U92);
  nand ginst11280 (P2_R1110_U332, P2_R1110_U138, P2_R1110_U331);
  nand ginst11281 (P2_R1110_U333, P2_R1110_U262, P2_R1110_U59);
  nand ginst11282 (P2_R1110_U334, P2_U3068, P2_U3440);
  nand ginst11283 (P2_R1110_U335, P2_R1110_U139, P2_R1110_U333);
  or ginst11284 (P2_R1110_U336, P2_U3072, P2_U3437);
  nand ginst11285 (P2_R1110_U337, P2_R1110_U167, P2_R1110_U250);
  not ginst11286 (P2_R1110_U338, P2_R1110_U93);
  or ginst11287 (P2_R1110_U339, P2_U3071, P2_U3425);
  nand ginst11288 (P2_R1110_U34, P2_U3059, P2_U3401);
  nand ginst11289 (P2_R1110_U340, P2_R1110_U339, P2_R1110_U93);
  nand ginst11290 (P2_R1110_U341, P2_R1110_U140, P2_R1110_U340);
  nand ginst11291 (P2_R1110_U342, P2_R1110_U172, P2_R1110_U338);
  nand ginst11292 (P2_R1110_U343, P2_U3079, P2_U3428);
  nand ginst11293 (P2_R1110_U344, P2_R1110_U141, P2_R1110_U342);
  or ginst11294 (P2_R1110_U345, P2_U3071, P2_U3425);
  or ginst11295 (P2_R1110_U346, P2_U3082, P2_U3416);
  nand ginst11296 (P2_R1110_U347, P2_R1110_U346, P2_R1110_U40);
  nand ginst11297 (P2_R1110_U348, P2_R1110_U142, P2_R1110_U347);
  nand ginst11298 (P2_R1110_U349, P2_R1110_U171, P2_R1110_U206);
  not ginst11299 (P2_R1110_U35, P2_U3404);
  nand ginst11300 (P2_R1110_U350, P2_U3061, P2_U3419);
  nand ginst11301 (P2_R1110_U351, P2_R1110_U143, P2_R1110_U349);
  nand ginst11302 (P2_R1110_U352, P2_R1110_U171, P2_R1110_U207);
  nand ginst11303 (P2_R1110_U353, P2_R1110_U204, P2_R1110_U65);
  nand ginst11304 (P2_R1110_U354, P2_R1110_U214, P2_R1110_U22);
  nand ginst11305 (P2_R1110_U355, P2_R1110_U228, P2_R1110_U34);
  nand ginst11306 (P2_R1110_U356, P2_R1110_U180, P2_R1110_U231);
  nand ginst11307 (P2_R1110_U357, P2_R1110_U173, P2_R1110_U314);
  nand ginst11308 (P2_R1110_U358, P2_R1110_U176, P2_R1110_U298);
  nand ginst11309 (P2_R1110_U359, P2_R1110_U329, P2_R1110_U80);
  not ginst11310 (P2_R1110_U36, P2_U3413);
  nand ginst11311 (P2_R1110_U360, P2_R1110_U282, P2_R1110_U77);
  nand ginst11312 (P2_R1110_U361, P2_R1110_U336, P2_R1110_U59);
  nand ginst11313 (P2_R1110_U362, P2_R1110_U172, P2_R1110_U345);
  nand ginst11314 (P2_R1110_U363, P2_R1110_U250, P2_R1110_U68);
  nand ginst11315 (P2_R1110_U364, P2_U3053, P2_U3895);
  nand ginst11316 (P2_R1110_U365, P2_R1110_U168, P2_R1110_U296);
  nand ginst11317 (P2_R1110_U366, P2_R1110_U295, P2_U3056);
  nand ginst11318 (P2_R1110_U367, P2_R1110_U295, P2_U3897);
  nand ginst11319 (P2_R1110_U368, P2_R1110_U168, P2_R1110_U296, P2_R1110_U301);
  nand ginst11320 (P2_R1110_U369, P2_R1110_U133, P2_R1110_U155, P2_R1110_U168);
  not ginst11321 (P2_R1110_U37, P2_U3083);
  nand ginst11322 (P2_R1110_U370, P2_R1110_U297, P2_R1110_U301);
  nand ginst11323 (P2_R1110_U371, P2_R1110_U39, P2_U3082);
  nand ginst11324 (P2_R1110_U372, P2_R1110_U38, P2_U3416);
  nand ginst11325 (P2_R1110_U373, P2_R1110_U371, P2_R1110_U372);
  nand ginst11326 (P2_R1110_U374, P2_R1110_U352, P2_R1110_U40);
  nand ginst11327 (P2_R1110_U375, P2_R1110_U206, P2_R1110_U373);
  nand ginst11328 (P2_R1110_U376, P2_R1110_U36, P2_U3083);
  nand ginst11329 (P2_R1110_U377, P2_R1110_U37, P2_U3413);
  nand ginst11330 (P2_R1110_U378, P2_R1110_U376, P2_R1110_U377);
  nand ginst11331 (P2_R1110_U379, P2_R1110_U144, P2_R1110_U353);
  not ginst11332 (P2_R1110_U38, P2_U3082);
  nand ginst11333 (P2_R1110_U380, P2_R1110_U203, P2_R1110_U378);
  nand ginst11334 (P2_R1110_U381, P2_R1110_U23, P2_U3069);
  nand ginst11335 (P2_R1110_U382, P2_R1110_U21, P2_U3410);
  nand ginst11336 (P2_R1110_U383, P2_R1110_U19, P2_U3070);
  nand ginst11337 (P2_R1110_U384, P2_R1110_U20, P2_U3407);
  nand ginst11338 (P2_R1110_U385, P2_R1110_U383, P2_R1110_U384);
  nand ginst11339 (P2_R1110_U386, P2_R1110_U354, P2_R1110_U41);
  nand ginst11340 (P2_R1110_U387, P2_R1110_U195, P2_R1110_U385);
  nand ginst11341 (P2_R1110_U388, P2_R1110_U35, P2_U3066);
  nand ginst11342 (P2_R1110_U389, P2_R1110_U26, P2_U3404);
  not ginst11343 (P2_R1110_U39, P2_U3416);
  nand ginst11344 (P2_R1110_U390, P2_R1110_U24, P2_U3059);
  nand ginst11345 (P2_R1110_U391, P2_R1110_U25, P2_U3401);
  nand ginst11346 (P2_R1110_U392, P2_R1110_U390, P2_R1110_U391);
  nand ginst11347 (P2_R1110_U393, P2_R1110_U355, P2_R1110_U44);
  nand ginst11348 (P2_R1110_U394, P2_R1110_U221, P2_R1110_U392);
  nand ginst11349 (P2_R1110_U395, P2_R1110_U32, P2_U3063);
  nand ginst11350 (P2_R1110_U396, P2_R1110_U33, P2_U3398);
  nand ginst11351 (P2_R1110_U397, P2_R1110_U395, P2_R1110_U396);
  nand ginst11352 (P2_R1110_U398, P2_R1110_U145, P2_R1110_U356);
  nand ginst11353 (P2_R1110_U399, P2_R1110_U230, P2_R1110_U397);
  and ginst11354 (P2_R1110_U4, P2_R1110_U178, P2_R1110_U179);
  nand ginst11355 (P2_R1110_U40, P2_R1110_U205, P2_R1110_U65);
  nand ginst11356 (P2_R1110_U400, P2_R1110_U27, P2_U3067);
  nand ginst11357 (P2_R1110_U401, P2_R1110_U28, P2_U3395);
  nand ginst11358 (P2_R1110_U402, P2_R1110_U147, P2_U3054);
  nand ginst11359 (P2_R1110_U403, P2_R1110_U146, P2_U3904);
  nand ginst11360 (P2_R1110_U404, P2_R1110_U147, P2_U3054);
  nand ginst11361 (P2_R1110_U405, P2_R1110_U146, P2_U3904);
  nand ginst11362 (P2_R1110_U406, P2_R1110_U404, P2_R1110_U405);
  nand ginst11363 (P2_R1110_U407, P2_R1110_U148, P2_R1110_U149);
  nand ginst11364 (P2_R1110_U408, P2_R1110_U305, P2_R1110_U406);
  nand ginst11365 (P2_R1110_U409, P2_R1110_U88, P2_U3053);
  nand ginst11366 (P2_R1110_U41, P2_R1110_U117, P2_R1110_U193);
  nand ginst11367 (P2_R1110_U410, P2_R1110_U87, P2_U3895);
  nand ginst11368 (P2_R1110_U411, P2_R1110_U88, P2_U3053);
  nand ginst11369 (P2_R1110_U412, P2_R1110_U87, P2_U3895);
  nand ginst11370 (P2_R1110_U413, P2_R1110_U411, P2_R1110_U412);
  nand ginst11371 (P2_R1110_U414, P2_R1110_U150, P2_R1110_U151);
  nand ginst11372 (P2_R1110_U415, P2_R1110_U303, P2_R1110_U413);
  nand ginst11373 (P2_R1110_U416, P2_R1110_U46, P2_U3052);
  nand ginst11374 (P2_R1110_U417, P2_R1110_U47, P2_U3896);
  nand ginst11375 (P2_R1110_U418, P2_R1110_U46, P2_U3052);
  nand ginst11376 (P2_R1110_U419, P2_R1110_U47, P2_U3896);
  nand ginst11377 (P2_R1110_U42, P2_R1110_U182, P2_R1110_U183);
  nand ginst11378 (P2_R1110_U420, P2_R1110_U418, P2_R1110_U419);
  nand ginst11379 (P2_R1110_U421, P2_R1110_U152, P2_R1110_U153);
  nand ginst11380 (P2_R1110_U422, P2_R1110_U300, P2_R1110_U420);
  nand ginst11381 (P2_R1110_U423, P2_R1110_U49, P2_U3056);
  nand ginst11382 (P2_R1110_U424, P2_R1110_U48, P2_U3897);
  nand ginst11383 (P2_R1110_U425, P2_R1110_U50, P2_U3057);
  nand ginst11384 (P2_R1110_U426, P2_R1110_U51, P2_U3898);
  nand ginst11385 (P2_R1110_U427, P2_R1110_U425, P2_R1110_U426);
  nand ginst11386 (P2_R1110_U428, P2_R1110_U357, P2_R1110_U89);
  nand ginst11387 (P2_R1110_U429, P2_R1110_U307, P2_R1110_U427);
  nand ginst11388 (P2_R1110_U43, P2_U3077, P2_U3392);
  nand ginst11389 (P2_R1110_U430, P2_R1110_U52, P2_U3064);
  nand ginst11390 (P2_R1110_U431, P2_R1110_U53, P2_U3899);
  nand ginst11391 (P2_R1110_U432, P2_R1110_U430, P2_R1110_U431);
  nand ginst11392 (P2_R1110_U433, P2_R1110_U155, P2_R1110_U358);
  nand ginst11393 (P2_R1110_U434, P2_R1110_U294, P2_R1110_U432);
  nand ginst11394 (P2_R1110_U435, P2_R1110_U84, P2_U3065);
  nand ginst11395 (P2_R1110_U436, P2_R1110_U85, P2_U3900);
  nand ginst11396 (P2_R1110_U437, P2_R1110_U84, P2_U3065);
  nand ginst11397 (P2_R1110_U438, P2_R1110_U85, P2_U3900);
  nand ginst11398 (P2_R1110_U439, P2_R1110_U437, P2_R1110_U438);
  nand ginst11399 (P2_R1110_U44, P2_R1110_U122, P2_R1110_U219);
  nand ginst11400 (P2_R1110_U440, P2_R1110_U156, P2_R1110_U157);
  nand ginst11401 (P2_R1110_U441, P2_R1110_U290, P2_R1110_U439);
  nand ginst11402 (P2_R1110_U442, P2_R1110_U82, P2_U3060);
  nand ginst11403 (P2_R1110_U443, P2_R1110_U83, P2_U3901);
  nand ginst11404 (P2_R1110_U444, P2_R1110_U82, P2_U3060);
  nand ginst11405 (P2_R1110_U445, P2_R1110_U83, P2_U3901);
  nand ginst11406 (P2_R1110_U446, P2_R1110_U444, P2_R1110_U445);
  nand ginst11407 (P2_R1110_U447, P2_R1110_U158, P2_R1110_U159);
  nand ginst11408 (P2_R1110_U448, P2_R1110_U286, P2_R1110_U446);
  nand ginst11409 (P2_R1110_U449, P2_R1110_U54, P2_U3074);
  nand ginst11410 (P2_R1110_U45, P2_R1110_U215, P2_R1110_U216);
  nand ginst11411 (P2_R1110_U450, P2_R1110_U55, P2_U3902);
  nand ginst11412 (P2_R1110_U451, P2_R1110_U54, P2_U3074);
  nand ginst11413 (P2_R1110_U452, P2_R1110_U55, P2_U3902);
  nand ginst11414 (P2_R1110_U453, P2_R1110_U451, P2_R1110_U452);
  nand ginst11415 (P2_R1110_U454, P2_R1110_U81, P2_U3075);
  nand ginst11416 (P2_R1110_U455, P2_R1110_U90, P2_U3903);
  nand ginst11417 (P2_R1110_U456, P2_R1110_U161, P2_R1110_U182);
  nand ginst11418 (P2_R1110_U457, P2_R1110_U31, P2_R1110_U328);
  nand ginst11419 (P2_R1110_U458, P2_R1110_U78, P2_U3080);
  nand ginst11420 (P2_R1110_U459, P2_R1110_U79, P2_U3445);
  not ginst11421 (P2_R1110_U46, P2_U3896);
  nand ginst11422 (P2_R1110_U460, P2_R1110_U458, P2_R1110_U459);
  nand ginst11423 (P2_R1110_U461, P2_R1110_U359, P2_R1110_U91);
  nand ginst11424 (P2_R1110_U462, P2_R1110_U316, P2_R1110_U460);
  nand ginst11425 (P2_R1110_U463, P2_R1110_U75, P2_U3081);
  nand ginst11426 (P2_R1110_U464, P2_R1110_U76, P2_U3443);
  nand ginst11427 (P2_R1110_U465, P2_R1110_U463, P2_R1110_U464);
  nand ginst11428 (P2_R1110_U466, P2_R1110_U162, P2_R1110_U360);
  nand ginst11429 (P2_R1110_U467, P2_R1110_U270, P2_R1110_U465);
  nand ginst11430 (P2_R1110_U468, P2_R1110_U60, P2_U3068);
  nand ginst11431 (P2_R1110_U469, P2_R1110_U58, P2_U3440);
  not ginst11432 (P2_R1110_U47, P2_U3052);
  nand ginst11433 (P2_R1110_U470, P2_R1110_U56, P2_U3072);
  nand ginst11434 (P2_R1110_U471, P2_R1110_U57, P2_U3437);
  nand ginst11435 (P2_R1110_U472, P2_R1110_U470, P2_R1110_U471);
  nand ginst11436 (P2_R1110_U473, P2_R1110_U361, P2_R1110_U92);
  nand ginst11437 (P2_R1110_U474, P2_R1110_U262, P2_R1110_U472);
  nand ginst11438 (P2_R1110_U475, P2_R1110_U73, P2_U3073);
  nand ginst11439 (P2_R1110_U476, P2_R1110_U74, P2_U3434);
  nand ginst11440 (P2_R1110_U477, P2_R1110_U73, P2_U3073);
  nand ginst11441 (P2_R1110_U478, P2_R1110_U74, P2_U3434);
  nand ginst11442 (P2_R1110_U479, P2_R1110_U477, P2_R1110_U478);
  not ginst11443 (P2_R1110_U48, P2_U3056);
  nand ginst11444 (P2_R1110_U480, P2_R1110_U163, P2_R1110_U164);
  nand ginst11445 (P2_R1110_U481, P2_R1110_U258, P2_R1110_U479);
  nand ginst11446 (P2_R1110_U482, P2_R1110_U71, P2_U3078);
  nand ginst11447 (P2_R1110_U483, P2_R1110_U72, P2_U3431);
  nand ginst11448 (P2_R1110_U484, P2_R1110_U71, P2_U3078);
  nand ginst11449 (P2_R1110_U485, P2_R1110_U72, P2_U3431);
  nand ginst11450 (P2_R1110_U486, P2_R1110_U484, P2_R1110_U485);
  nand ginst11451 (P2_R1110_U487, P2_R1110_U165, P2_R1110_U166);
  nand ginst11452 (P2_R1110_U488, P2_R1110_U254, P2_R1110_U486);
  nand ginst11453 (P2_R1110_U489, P2_R1110_U61, P2_U3079);
  not ginst11454 (P2_R1110_U49, P2_U3897);
  nand ginst11455 (P2_R1110_U490, P2_R1110_U62, P2_U3428);
  nand ginst11456 (P2_R1110_U491, P2_R1110_U69, P2_U3071);
  nand ginst11457 (P2_R1110_U492, P2_R1110_U70, P2_U3425);
  nand ginst11458 (P2_R1110_U493, P2_R1110_U491, P2_R1110_U492);
  nand ginst11459 (P2_R1110_U494, P2_R1110_U362, P2_R1110_U93);
  nand ginst11460 (P2_R1110_U495, P2_R1110_U338, P2_R1110_U493);
  nand ginst11461 (P2_R1110_U496, P2_R1110_U66, P2_U3062);
  nand ginst11462 (P2_R1110_U497, P2_R1110_U67, P2_U3422);
  nand ginst11463 (P2_R1110_U498, P2_R1110_U496, P2_R1110_U497);
  nand ginst11464 (P2_R1110_U499, P2_R1110_U167, P2_R1110_U363);
  and ginst11465 (P2_R1110_U5, P2_R1110_U196, P2_R1110_U197);
  not ginst11466 (P2_R1110_U50, P2_U3898);
  nand ginst11467 (P2_R1110_U500, P2_R1110_U244, P2_R1110_U498);
  nand ginst11468 (P2_R1110_U501, P2_R1110_U63, P2_U3061);
  nand ginst11469 (P2_R1110_U502, P2_R1110_U64, P2_U3419);
  nand ginst11470 (P2_R1110_U503, P2_R1110_U29, P2_U3076);
  nand ginst11471 (P2_R1110_U504, P2_R1110_U30, P2_U3387);
  not ginst11472 (P2_R1110_U51, P2_U3057);
  not ginst11473 (P2_R1110_U52, P2_U3899);
  not ginst11474 (P2_R1110_U53, P2_U3064);
  not ginst11475 (P2_R1110_U54, P2_U3902);
  not ginst11476 (P2_R1110_U55, P2_U3074);
  not ginst11477 (P2_R1110_U56, P2_U3437);
  not ginst11478 (P2_R1110_U57, P2_U3072);
  not ginst11479 (P2_R1110_U58, P2_U3068);
  nand ginst11480 (P2_R1110_U59, P2_U3072, P2_U3437);
  and ginst11481 (P2_R1110_U6, P2_R1110_U236, P2_R1110_U237);
  not ginst11482 (P2_R1110_U60, P2_U3440);
  not ginst11483 (P2_R1110_U61, P2_U3428);
  not ginst11484 (P2_R1110_U62, P2_U3079);
  not ginst11485 (P2_R1110_U63, P2_U3419);
  not ginst11486 (P2_R1110_U64, P2_U3061);
  nand ginst11487 (P2_R1110_U65, P2_U3083, P2_U3413);
  not ginst11488 (P2_R1110_U66, P2_U3422);
  not ginst11489 (P2_R1110_U67, P2_U3062);
  nand ginst11490 (P2_R1110_U68, P2_U3062, P2_U3422);
  not ginst11491 (P2_R1110_U69, P2_U3425);
  and ginst11492 (P2_R1110_U7, P2_R1110_U245, P2_R1110_U246);
  not ginst11493 (P2_R1110_U70, P2_U3071);
  not ginst11494 (P2_R1110_U71, P2_U3431);
  not ginst11495 (P2_R1110_U72, P2_U3078);
  not ginst11496 (P2_R1110_U73, P2_U3434);
  not ginst11497 (P2_R1110_U74, P2_U3073);
  not ginst11498 (P2_R1110_U75, P2_U3443);
  not ginst11499 (P2_R1110_U76, P2_U3081);
  nand ginst11500 (P2_R1110_U77, P2_U3081, P2_U3443);
  not ginst11501 (P2_R1110_U78, P2_U3445);
  not ginst11502 (P2_R1110_U79, P2_U3080);
  and ginst11503 (P2_R1110_U8, P2_R1110_U263, P2_R1110_U264);
  nand ginst11504 (P2_R1110_U80, P2_U3080, P2_U3445);
  not ginst11505 (P2_R1110_U81, P2_U3903);
  not ginst11506 (P2_R1110_U82, P2_U3901);
  not ginst11507 (P2_R1110_U83, P2_U3060);
  not ginst11508 (P2_R1110_U84, P2_U3900);
  not ginst11509 (P2_R1110_U85, P2_U3065);
  nand ginst11510 (P2_R1110_U86, P2_U3056, P2_U3897);
  not ginst11511 (P2_R1110_U87, P2_U3053);
  not ginst11512 (P2_R1110_U88, P2_U3895);
  nand ginst11513 (P2_R1110_U89, P2_R1110_U176, P2_R1110_U306);
  and ginst11514 (P2_R1110_U9, P2_R1110_U271, P2_R1110_U272);
  not ginst11515 (P2_R1110_U90, P2_U3075);
  nand ginst11516 (P2_R1110_U91, P2_R1110_U315, P2_R1110_U77);
  nand ginst11517 (P2_R1110_U92, P2_R1110_U260, P2_R1110_U261);
  nand ginst11518 (P2_R1110_U93, P2_R1110_U337, P2_R1110_U68);
  nand ginst11519 (P2_R1110_U94, P2_R1110_U456, P2_R1110_U457);
  nand ginst11520 (P2_R1110_U95, P2_R1110_U503, P2_R1110_U504);
  nand ginst11521 (P2_R1110_U96, P2_R1110_U374, P2_R1110_U375);
  nand ginst11522 (P2_R1110_U97, P2_R1110_U379, P2_R1110_U380);
  nand ginst11523 (P2_R1110_U98, P2_R1110_U386, P2_R1110_U387);
  nand ginst11524 (P2_R1110_U99, P2_R1110_U393, P2_R1110_U394);
  and ginst11525 (P2_R1131_U10, P2_R1131_U194, P2_R1131_U281);
  nand ginst11526 (P2_R1131_U100, P2_R1131_U424, P2_R1131_U425);
  nand ginst11527 (P2_R1131_U101, P2_R1131_U440, P2_R1131_U441);
  nand ginst11528 (P2_R1131_U102, P2_R1131_U445, P2_R1131_U446);
  nand ginst11529 (P2_R1131_U103, P2_R1131_U450, P2_R1131_U451);
  nand ginst11530 (P2_R1131_U104, P2_R1131_U455, P2_R1131_U456);
  nand ginst11531 (P2_R1131_U105, P2_R1131_U460, P2_R1131_U461);
  nand ginst11532 (P2_R1131_U106, P2_R1131_U476, P2_R1131_U477);
  nand ginst11533 (P2_R1131_U107, P2_R1131_U481, P2_R1131_U482);
  nand ginst11534 (P2_R1131_U108, P2_R1131_U364, P2_R1131_U365);
  nand ginst11535 (P2_R1131_U109, P2_R1131_U373, P2_R1131_U374);
  and ginst11536 (P2_R1131_U11, P2_R1131_U282, P2_R1131_U283);
  nand ginst11537 (P2_R1131_U110, P2_R1131_U380, P2_R1131_U381);
  nand ginst11538 (P2_R1131_U111, P2_R1131_U384, P2_R1131_U385);
  nand ginst11539 (P2_R1131_U112, P2_R1131_U393, P2_R1131_U394);
  nand ginst11540 (P2_R1131_U113, P2_R1131_U414, P2_R1131_U415);
  nand ginst11541 (P2_R1131_U114, P2_R1131_U431, P2_R1131_U432);
  nand ginst11542 (P2_R1131_U115, P2_R1131_U435, P2_R1131_U436);
  nand ginst11543 (P2_R1131_U116, P2_R1131_U467, P2_R1131_U468);
  nand ginst11544 (P2_R1131_U117, P2_R1131_U471, P2_R1131_U472);
  nand ginst11545 (P2_R1131_U118, P2_R1131_U488, P2_R1131_U489);
  and ginst11546 (P2_R1131_U119, P2_R1131_U196, P2_R1131_U206);
  and ginst11547 (P2_R1131_U12, P2_R1131_U195, P2_R1131_U299);
  and ginst11548 (P2_R1131_U120, P2_R1131_U208, P2_R1131_U209);
  and ginst11549 (P2_R1131_U121, P2_R1131_U13, P2_R1131_U14);
  and ginst11550 (P2_R1131_U122, P2_R1131_U222, P2_R1131_U340);
  and ginst11551 (P2_R1131_U123, P2_R1131_U122, P2_R1131_U342);
  and ginst11552 (P2_R1131_U124, P2_R1131_U27, P2_R1131_U366, P2_R1131_U367);
  and ginst11553 (P2_R1131_U125, P2_R1131_U198, P2_R1131_U370);
  and ginst11554 (P2_R1131_U126, P2_R1131_U237, P2_R1131_U6);
  and ginst11555 (P2_R1131_U127, P2_R1131_U197, P2_R1131_U377);
  and ginst11556 (P2_R1131_U128, P2_R1131_U35, P2_R1131_U386, P2_R1131_U387);
  and ginst11557 (P2_R1131_U129, P2_R1131_U196, P2_R1131_U390);
  and ginst11558 (P2_R1131_U13, P2_R1131_U197, P2_R1131_U210, P2_R1131_U215);
  and ginst11559 (P2_R1131_U130, P2_R1131_U15, P2_R1131_U251);
  and ginst11560 (P2_R1131_U131, P2_R1131_U252, P2_R1131_U343);
  and ginst11561 (P2_R1131_U132, P2_R1131_U262, P2_R1131_U8);
  and ginst11562 (P2_R1131_U133, P2_R1131_U10, P2_R1131_U286);
  and ginst11563 (P2_R1131_U134, P2_R1131_U301, P2_R1131_U302);
  and ginst11564 (P2_R1131_U135, P2_R1131_U303, P2_R1131_U397);
  and ginst11565 (P2_R1131_U136, P2_R1131_U16, P2_R1131_U301, P2_R1131_U302, P2_R1131_U304);
  and ginst11566 (P2_R1131_U137, P2_R1131_U165, P2_R1131_U359);
  nand ginst11567 (P2_R1131_U138, P2_R1131_U402, P2_R1131_U403);
  and ginst11568 (P2_R1131_U139, P2_R1131_U407, P2_R1131_U408, P2_R1131_U53);
  and ginst11569 (P2_R1131_U14, P2_R1131_U198, P2_R1131_U220);
  and ginst11570 (P2_R1131_U140, P2_R1131_U195, P2_R1131_U411);
  nand ginst11571 (P2_R1131_U141, P2_R1131_U416, P2_R1131_U417);
  nand ginst11572 (P2_R1131_U142, P2_R1131_U421, P2_R1131_U422);
  and ginst11573 (P2_R1131_U143, P2_R1131_U11, P2_R1131_U313);
  and ginst11574 (P2_R1131_U144, P2_R1131_U194, P2_R1131_U428);
  nand ginst11575 (P2_R1131_U145, P2_R1131_U437, P2_R1131_U438);
  nand ginst11576 (P2_R1131_U146, P2_R1131_U442, P2_R1131_U443);
  nand ginst11577 (P2_R1131_U147, P2_R1131_U447, P2_R1131_U448);
  nand ginst11578 (P2_R1131_U148, P2_R1131_U452, P2_R1131_U453);
  nand ginst11579 (P2_R1131_U149, P2_R1131_U457, P2_R1131_U458);
  and ginst11580 (P2_R1131_U15, P2_R1131_U192, P2_R1131_U224, P2_R1131_U244);
  and ginst11581 (P2_R1131_U150, P2_R1131_U324, P2_R1131_U9);
  and ginst11582 (P2_R1131_U151, P2_R1131_U193, P2_R1131_U464);
  nand ginst11583 (P2_R1131_U152, P2_R1131_U473, P2_R1131_U474);
  nand ginst11584 (P2_R1131_U153, P2_R1131_U478, P2_R1131_U479);
  and ginst11585 (P2_R1131_U154, P2_R1131_U333, P2_R1131_U7);
  and ginst11586 (P2_R1131_U155, P2_R1131_U192, P2_R1131_U485);
  and ginst11587 (P2_R1131_U156, P2_R1131_U362, P2_R1131_U363);
  nand ginst11588 (P2_R1131_U157, P2_R1131_U123, P2_R1131_U341);
  and ginst11589 (P2_R1131_U158, P2_R1131_U371, P2_R1131_U372);
  and ginst11590 (P2_R1131_U159, P2_R1131_U378, P2_R1131_U379);
  and ginst11591 (P2_R1131_U16, P2_R1131_U398, P2_R1131_U399);
  and ginst11592 (P2_R1131_U160, P2_R1131_U382, P2_R1131_U383);
  nand ginst11593 (P2_R1131_U161, P2_R1131_U120, P2_R1131_U344);
  and ginst11594 (P2_R1131_U162, P2_R1131_U391, P2_R1131_U392);
  not ginst11595 (P2_R1131_U163, P2_U3904);
  not ginst11596 (P2_R1131_U164, P2_U3054);
  and ginst11597 (P2_R1131_U165, P2_R1131_U400, P2_R1131_U401);
  nand ginst11598 (P2_R1131_U166, P2_R1131_U134, P2_R1131_U360);
  and ginst11599 (P2_R1131_U167, P2_R1131_U412, P2_R1131_U413);
  nand ginst11600 (P2_R1131_U168, P2_R1131_U292, P2_R1131_U293);
  nand ginst11601 (P2_R1131_U169, P2_R1131_U288, P2_R1131_U289);
  nand ginst11602 (P2_R1131_U17, P2_R1131_U331, P2_R1131_U334);
  and ginst11603 (P2_R1131_U170, P2_R1131_U429, P2_R1131_U430);
  and ginst11604 (P2_R1131_U171, P2_R1131_U433, P2_R1131_U434);
  nand ginst11605 (P2_R1131_U172, P2_R1131_U278, P2_R1131_U279);
  nand ginst11606 (P2_R1131_U173, P2_R1131_U274, P2_R1131_U275);
  not ginst11607 (P2_R1131_U174, P2_U3392);
  nand ginst11608 (P2_R1131_U175, P2_R1131_U97, P2_U3387);
  nand ginst11609 (P2_R1131_U176, P2_R1131_U187, P2_R1131_U271, P2_R1131_U339);
  not ginst11610 (P2_R1131_U177, P2_U3443);
  nand ginst11611 (P2_R1131_U178, P2_R1131_U268, P2_R1131_U269);
  nand ginst11612 (P2_R1131_U179, P2_R1131_U264, P2_R1131_U265);
  nand ginst11613 (P2_R1131_U18, P2_R1131_U322, P2_R1131_U325);
  and ginst11614 (P2_R1131_U180, P2_R1131_U465, P2_R1131_U466);
  and ginst11615 (P2_R1131_U181, P2_R1131_U469, P2_R1131_U470);
  nand ginst11616 (P2_R1131_U182, P2_R1131_U254, P2_R1131_U255);
  nand ginst11617 (P2_R1131_U183, P2_R1131_U131, P2_R1131_U353);
  nand ginst11618 (P2_R1131_U184, P2_R1131_U351, P2_R1131_U62);
  and ginst11619 (P2_R1131_U185, P2_R1131_U486, P2_R1131_U487);
  nand ginst11620 (P2_R1131_U186, P2_R1131_U135, P2_R1131_U166);
  nand ginst11621 (P2_R1131_U187, P2_R1131_U177, P2_R1131_U178);
  nand ginst11622 (P2_R1131_U188, P2_R1131_U174, P2_R1131_U175);
  not ginst11623 (P2_R1131_U189, P2_R1131_U53);
  nand ginst11624 (P2_R1131_U19, P2_R1131_U311, P2_R1131_U314);
  not ginst11625 (P2_R1131_U190, P2_R1131_U35);
  not ginst11626 (P2_R1131_U191, P2_R1131_U27);
  nand ginst11627 (P2_R1131_U192, P2_R1131_U57, P2_U3419);
  nand ginst11628 (P2_R1131_U193, P2_R1131_U69, P2_U3434);
  nand ginst11629 (P2_R1131_U194, P2_R1131_U83, P2_U3901);
  nand ginst11630 (P2_R1131_U195, P2_R1131_U52, P2_U3897);
  nand ginst11631 (P2_R1131_U196, P2_R1131_U34, P2_U3395);
  nand ginst11632 (P2_R1131_U197, P2_R1131_U42, P2_U3404);
  nand ginst11633 (P2_R1131_U198, P2_R1131_U26, P2_U3410);
  not ginst11634 (P2_R1131_U199, P2_R1131_U71);
  nand ginst11635 (P2_R1131_U20, P2_R1131_U305, P2_R1131_U357);
  not ginst11636 (P2_R1131_U200, P2_R1131_U85);
  not ginst11637 (P2_R1131_U201, P2_R1131_U44);
  not ginst11638 (P2_R1131_U202, P2_R1131_U59);
  not ginst11639 (P2_R1131_U203, P2_R1131_U175);
  nand ginst11640 (P2_R1131_U204, P2_R1131_U175, P2_U3077);
  not ginst11641 (P2_R1131_U205, P2_R1131_U50);
  nand ginst11642 (P2_R1131_U206, P2_R1131_U36, P2_U3398);
  nand ginst11643 (P2_R1131_U207, P2_R1131_U35, P2_R1131_U36);
  nand ginst11644 (P2_R1131_U208, P2_R1131_U207, P2_R1131_U40);
  nand ginst11645 (P2_R1131_U209, P2_R1131_U190, P2_U3063);
  nand ginst11646 (P2_R1131_U21, P2_R1131_U137, P2_R1131_U186);
  nand ginst11647 (P2_R1131_U210, P2_R1131_U41, P2_U3407);
  nand ginst11648 (P2_R1131_U211, P2_R1131_U30, P2_U3070);
  nand ginst11649 (P2_R1131_U212, P2_R1131_U29, P2_U3066);
  nand ginst11650 (P2_R1131_U213, P2_R1131_U197, P2_R1131_U201);
  nand ginst11651 (P2_R1131_U214, P2_R1131_U213, P2_R1131_U6);
  nand ginst11652 (P2_R1131_U215, P2_R1131_U43, P2_U3401);
  nand ginst11653 (P2_R1131_U216, P2_R1131_U41, P2_U3407);
  nand ginst11654 (P2_R1131_U217, P2_R1131_U13, P2_R1131_U161);
  not ginst11655 (P2_R1131_U218, P2_R1131_U45);
  not ginst11656 (P2_R1131_U219, P2_R1131_U48);
  nand ginst11657 (P2_R1131_U22, P2_R1131_U242, P2_R1131_U347);
  nand ginst11658 (P2_R1131_U220, P2_R1131_U28, P2_U3413);
  nand ginst11659 (P2_R1131_U221, P2_R1131_U27, P2_R1131_U28);
  nand ginst11660 (P2_R1131_U222, P2_R1131_U191, P2_U3083);
  not ginst11661 (P2_R1131_U223, P2_R1131_U157);
  nand ginst11662 (P2_R1131_U224, P2_R1131_U47, P2_U3416);
  nand ginst11663 (P2_R1131_U225, P2_R1131_U224, P2_R1131_U59);
  nand ginst11664 (P2_R1131_U226, P2_R1131_U219, P2_R1131_U27);
  nand ginst11665 (P2_R1131_U227, P2_R1131_U125, P2_R1131_U226);
  nand ginst11666 (P2_R1131_U228, P2_R1131_U198, P2_R1131_U48);
  nand ginst11667 (P2_R1131_U229, P2_R1131_U124, P2_R1131_U228);
  nand ginst11668 (P2_R1131_U23, P2_R1131_U235, P2_R1131_U238);
  nand ginst11669 (P2_R1131_U230, P2_R1131_U198, P2_R1131_U27);
  nand ginst11670 (P2_R1131_U231, P2_R1131_U161, P2_R1131_U215);
  not ginst11671 (P2_R1131_U232, P2_R1131_U49);
  nand ginst11672 (P2_R1131_U233, P2_R1131_U29, P2_U3066);
  nand ginst11673 (P2_R1131_U234, P2_R1131_U232, P2_R1131_U233);
  nand ginst11674 (P2_R1131_U235, P2_R1131_U127, P2_R1131_U234);
  nand ginst11675 (P2_R1131_U236, P2_R1131_U197, P2_R1131_U49);
  nand ginst11676 (P2_R1131_U237, P2_R1131_U41, P2_U3407);
  nand ginst11677 (P2_R1131_U238, P2_R1131_U126, P2_R1131_U236);
  nand ginst11678 (P2_R1131_U239, P2_R1131_U29, P2_U3066);
  nand ginst11679 (P2_R1131_U24, P2_R1131_U227, P2_R1131_U229);
  nand ginst11680 (P2_R1131_U240, P2_R1131_U197, P2_R1131_U239);
  nand ginst11681 (P2_R1131_U241, P2_R1131_U215, P2_R1131_U44);
  nand ginst11682 (P2_R1131_U242, P2_R1131_U129, P2_R1131_U348);
  nand ginst11683 (P2_R1131_U243, P2_R1131_U196, P2_R1131_U35);
  nand ginst11684 (P2_R1131_U244, P2_R1131_U56, P2_U3422);
  nand ginst11685 (P2_R1131_U245, P2_R1131_U60, P2_U3062);
  nand ginst11686 (P2_R1131_U246, P2_R1131_U58, P2_U3061);
  nand ginst11687 (P2_R1131_U247, P2_R1131_U192, P2_R1131_U202);
  nand ginst11688 (P2_R1131_U248, P2_R1131_U247, P2_R1131_U7);
  nand ginst11689 (P2_R1131_U249, P2_R1131_U56, P2_U3422);
  nand ginst11690 (P2_R1131_U25, P2_R1131_U175, P2_R1131_U337);
  not ginst11691 (P2_R1131_U250, P2_R1131_U62);
  nand ginst11692 (P2_R1131_U251, P2_R1131_U55, P2_U3425);
  nand ginst11693 (P2_R1131_U252, P2_R1131_U61, P2_U3071);
  nand ginst11694 (P2_R1131_U253, P2_R1131_U64, P2_U3428);
  nand ginst11695 (P2_R1131_U254, P2_R1131_U183, P2_R1131_U253);
  nand ginst11696 (P2_R1131_U255, P2_R1131_U63, P2_U3079);
  not ginst11697 (P2_R1131_U256, P2_R1131_U182);
  nand ginst11698 (P2_R1131_U257, P2_R1131_U68, P2_U3437);
  nand ginst11699 (P2_R1131_U258, P2_R1131_U65, P2_U3072);
  nand ginst11700 (P2_R1131_U259, P2_R1131_U66, P2_U3073);
  not ginst11701 (P2_R1131_U26, P2_U3069);
  nand ginst11702 (P2_R1131_U260, P2_R1131_U199, P2_R1131_U8);
  nand ginst11703 (P2_R1131_U261, P2_R1131_U260, P2_R1131_U9);
  nand ginst11704 (P2_R1131_U262, P2_R1131_U70, P2_U3431);
  nand ginst11705 (P2_R1131_U263, P2_R1131_U68, P2_U3437);
  nand ginst11706 (P2_R1131_U264, P2_R1131_U132, P2_R1131_U182);
  nand ginst11707 (P2_R1131_U265, P2_R1131_U261, P2_R1131_U263);
  not ginst11708 (P2_R1131_U266, P2_R1131_U179);
  nand ginst11709 (P2_R1131_U267, P2_R1131_U73, P2_U3440);
  nand ginst11710 (P2_R1131_U268, P2_R1131_U179, P2_R1131_U267);
  nand ginst11711 (P2_R1131_U269, P2_R1131_U72, P2_U3068);
  nand ginst11712 (P2_R1131_U27, P2_R1131_U32, P2_U3069);
  not ginst11713 (P2_R1131_U270, P2_R1131_U178);
  nand ginst11714 (P2_R1131_U271, P2_R1131_U178, P2_U3081);
  not ginst11715 (P2_R1131_U272, P2_R1131_U176);
  nand ginst11716 (P2_R1131_U273, P2_R1131_U76, P2_U3445);
  nand ginst11717 (P2_R1131_U274, P2_R1131_U176, P2_R1131_U273);
  nand ginst11718 (P2_R1131_U275, P2_R1131_U75, P2_U3080);
  not ginst11719 (P2_R1131_U276, P2_R1131_U173);
  nand ginst11720 (P2_R1131_U277, P2_R1131_U78, P2_U3903);
  nand ginst11721 (P2_R1131_U278, P2_R1131_U173, P2_R1131_U277);
  nand ginst11722 (P2_R1131_U279, P2_R1131_U77, P2_U3075);
  not ginst11723 (P2_R1131_U28, P2_U3083);
  not ginst11724 (P2_R1131_U280, P2_R1131_U172);
  nand ginst11725 (P2_R1131_U281, P2_R1131_U82, P2_U3900);
  nand ginst11726 (P2_R1131_U282, P2_R1131_U79, P2_U3065);
  nand ginst11727 (P2_R1131_U283, P2_R1131_U80, P2_U3060);
  nand ginst11728 (P2_R1131_U284, P2_R1131_U10, P2_R1131_U200);
  nand ginst11729 (P2_R1131_U285, P2_R1131_U11, P2_R1131_U284);
  nand ginst11730 (P2_R1131_U286, P2_R1131_U84, P2_U3902);
  nand ginst11731 (P2_R1131_U287, P2_R1131_U82, P2_U3900);
  nand ginst11732 (P2_R1131_U288, P2_R1131_U133, P2_R1131_U172);
  nand ginst11733 (P2_R1131_U289, P2_R1131_U285, P2_R1131_U287);
  not ginst11734 (P2_R1131_U29, P2_U3404);
  not ginst11735 (P2_R1131_U290, P2_R1131_U169);
  nand ginst11736 (P2_R1131_U291, P2_R1131_U87, P2_U3899);
  nand ginst11737 (P2_R1131_U292, P2_R1131_U169, P2_R1131_U291);
  nand ginst11738 (P2_R1131_U293, P2_R1131_U86, P2_U3064);
  not ginst11739 (P2_R1131_U294, P2_R1131_U168);
  nand ginst11740 (P2_R1131_U295, P2_R1131_U89, P2_U3898);
  nand ginst11741 (P2_R1131_U296, P2_R1131_U168, P2_R1131_U295);
  nand ginst11742 (P2_R1131_U297, P2_R1131_U88, P2_U3057);
  not ginst11743 (P2_R1131_U298, P2_R1131_U93);
  nand ginst11744 (P2_R1131_U299, P2_R1131_U54, P2_U3896);
  not ginst11745 (P2_R1131_U30, P2_U3407);
  nand ginst11746 (P2_R1131_U300, P2_R1131_U53, P2_R1131_U54);
  nand ginst11747 (P2_R1131_U301, P2_R1131_U300, P2_R1131_U91);
  nand ginst11748 (P2_R1131_U302, P2_R1131_U189, P2_U3052);
  nand ginst11749 (P2_R1131_U303, P2_R1131_U92, P2_U3895);
  nand ginst11750 (P2_R1131_U304, P2_R1131_U51, P2_U3053);
  nand ginst11751 (P2_R1131_U305, P2_R1131_U140, P2_R1131_U355);
  nand ginst11752 (P2_R1131_U306, P2_R1131_U195, P2_R1131_U53);
  nand ginst11753 (P2_R1131_U307, P2_R1131_U172, P2_R1131_U286);
  not ginst11754 (P2_R1131_U308, P2_R1131_U94);
  nand ginst11755 (P2_R1131_U309, P2_R1131_U80, P2_U3060);
  not ginst11756 (P2_R1131_U31, P2_U3401);
  nand ginst11757 (P2_R1131_U310, P2_R1131_U308, P2_R1131_U309);
  nand ginst11758 (P2_R1131_U311, P2_R1131_U144, P2_R1131_U310);
  nand ginst11759 (P2_R1131_U312, P2_R1131_U194, P2_R1131_U94);
  nand ginst11760 (P2_R1131_U313, P2_R1131_U82, P2_U3900);
  nand ginst11761 (P2_R1131_U314, P2_R1131_U143, P2_R1131_U312);
  nand ginst11762 (P2_R1131_U315, P2_R1131_U80, P2_U3060);
  nand ginst11763 (P2_R1131_U316, P2_R1131_U194, P2_R1131_U315);
  nand ginst11764 (P2_R1131_U317, P2_R1131_U286, P2_R1131_U85);
  nand ginst11765 (P2_R1131_U318, P2_R1131_U182, P2_R1131_U262);
  not ginst11766 (P2_R1131_U319, P2_R1131_U95);
  not ginst11767 (P2_R1131_U32, P2_U3410);
  nand ginst11768 (P2_R1131_U320, P2_R1131_U66, P2_U3073);
  nand ginst11769 (P2_R1131_U321, P2_R1131_U319, P2_R1131_U320);
  nand ginst11770 (P2_R1131_U322, P2_R1131_U151, P2_R1131_U321);
  nand ginst11771 (P2_R1131_U323, P2_R1131_U193, P2_R1131_U95);
  nand ginst11772 (P2_R1131_U324, P2_R1131_U68, P2_U3437);
  nand ginst11773 (P2_R1131_U325, P2_R1131_U150, P2_R1131_U323);
  nand ginst11774 (P2_R1131_U326, P2_R1131_U66, P2_U3073);
  nand ginst11775 (P2_R1131_U327, P2_R1131_U193, P2_R1131_U326);
  nand ginst11776 (P2_R1131_U328, P2_R1131_U262, P2_R1131_U71);
  nand ginst11777 (P2_R1131_U329, P2_R1131_U58, P2_U3061);
  not ginst11778 (P2_R1131_U33, P2_U3413);
  nand ginst11779 (P2_R1131_U330, P2_R1131_U329, P2_R1131_U350);
  nand ginst11780 (P2_R1131_U331, P2_R1131_U155, P2_R1131_U330);
  nand ginst11781 (P2_R1131_U332, P2_R1131_U192, P2_R1131_U96);
  nand ginst11782 (P2_R1131_U333, P2_R1131_U56, P2_U3422);
  nand ginst11783 (P2_R1131_U334, P2_R1131_U154, P2_R1131_U332);
  nand ginst11784 (P2_R1131_U335, P2_R1131_U58, P2_U3061);
  nand ginst11785 (P2_R1131_U336, P2_R1131_U192, P2_R1131_U335);
  nand ginst11786 (P2_R1131_U337, P2_R1131_U38, P2_U3076);
  nand ginst11787 (P2_R1131_U338, P2_R1131_U174, P2_U3077);
  nand ginst11788 (P2_R1131_U339, P2_R1131_U177, P2_U3081);
  not ginst11789 (P2_R1131_U34, P2_U3067);
  nand ginst11790 (P2_R1131_U340, P2_R1131_U221, P2_R1131_U33);
  nand ginst11791 (P2_R1131_U341, P2_R1131_U121, P2_R1131_U161);
  nand ginst11792 (P2_R1131_U342, P2_R1131_U14, P2_R1131_U218);
  nand ginst11793 (P2_R1131_U343, P2_R1131_U250, P2_R1131_U251);
  nand ginst11794 (P2_R1131_U344, P2_R1131_U119, P2_R1131_U50);
  not ginst11795 (P2_R1131_U345, P2_R1131_U161);
  nand ginst11796 (P2_R1131_U346, P2_R1131_U196, P2_R1131_U50);
  nand ginst11797 (P2_R1131_U347, P2_R1131_U128, P2_R1131_U346);
  nand ginst11798 (P2_R1131_U348, P2_R1131_U205, P2_R1131_U35);
  nand ginst11799 (P2_R1131_U349, P2_R1131_U157, P2_R1131_U224);
  nand ginst11800 (P2_R1131_U35, P2_R1131_U37, P2_U3067);
  not ginst11801 (P2_R1131_U350, P2_R1131_U96);
  nand ginst11802 (P2_R1131_U351, P2_R1131_U15, P2_R1131_U157);
  not ginst11803 (P2_R1131_U352, P2_R1131_U184);
  nand ginst11804 (P2_R1131_U353, P2_R1131_U130, P2_R1131_U157);
  not ginst11805 (P2_R1131_U354, P2_R1131_U183);
  nand ginst11806 (P2_R1131_U355, P2_R1131_U298, P2_R1131_U53);
  nand ginst11807 (P2_R1131_U356, P2_R1131_U195, P2_R1131_U93);
  nand ginst11808 (P2_R1131_U357, P2_R1131_U139, P2_R1131_U356);
  nand ginst11809 (P2_R1131_U358, P2_R1131_U12, P2_R1131_U93);
  nand ginst11810 (P2_R1131_U359, P2_R1131_U136, P2_R1131_U358);
  not ginst11811 (P2_R1131_U36, P2_U3063);
  nand ginst11812 (P2_R1131_U360, P2_R1131_U12, P2_R1131_U93);
  not ginst11813 (P2_R1131_U361, P2_R1131_U166);
  nand ginst11814 (P2_R1131_U362, P2_R1131_U47, P2_U3416);
  nand ginst11815 (P2_R1131_U363, P2_R1131_U46, P2_U3082);
  nand ginst11816 (P2_R1131_U364, P2_R1131_U157, P2_R1131_U225);
  nand ginst11817 (P2_R1131_U365, P2_R1131_U156, P2_R1131_U223);
  nand ginst11818 (P2_R1131_U366, P2_R1131_U28, P2_U3413);
  nand ginst11819 (P2_R1131_U367, P2_R1131_U33, P2_U3083);
  nand ginst11820 (P2_R1131_U368, P2_R1131_U28, P2_U3413);
  nand ginst11821 (P2_R1131_U369, P2_R1131_U33, P2_U3083);
  not ginst11822 (P2_R1131_U37, P2_U3395);
  nand ginst11823 (P2_R1131_U370, P2_R1131_U368, P2_R1131_U369);
  nand ginst11824 (P2_R1131_U371, P2_R1131_U26, P2_U3410);
  nand ginst11825 (P2_R1131_U372, P2_R1131_U32, P2_U3069);
  nand ginst11826 (P2_R1131_U373, P2_R1131_U230, P2_R1131_U48);
  nand ginst11827 (P2_R1131_U374, P2_R1131_U158, P2_R1131_U219);
  nand ginst11828 (P2_R1131_U375, P2_R1131_U41, P2_U3407);
  nand ginst11829 (P2_R1131_U376, P2_R1131_U30, P2_U3070);
  nand ginst11830 (P2_R1131_U377, P2_R1131_U375, P2_R1131_U376);
  nand ginst11831 (P2_R1131_U378, P2_R1131_U42, P2_U3404);
  nand ginst11832 (P2_R1131_U379, P2_R1131_U29, P2_U3066);
  not ginst11833 (P2_R1131_U38, P2_U3387);
  nand ginst11834 (P2_R1131_U380, P2_R1131_U240, P2_R1131_U49);
  nand ginst11835 (P2_R1131_U381, P2_R1131_U159, P2_R1131_U232);
  nand ginst11836 (P2_R1131_U382, P2_R1131_U43, P2_U3401);
  nand ginst11837 (P2_R1131_U383, P2_R1131_U31, P2_U3059);
  nand ginst11838 (P2_R1131_U384, P2_R1131_U161, P2_R1131_U241);
  nand ginst11839 (P2_R1131_U385, P2_R1131_U160, P2_R1131_U345);
  nand ginst11840 (P2_R1131_U386, P2_R1131_U36, P2_U3398);
  nand ginst11841 (P2_R1131_U387, P2_R1131_U40, P2_U3063);
  nand ginst11842 (P2_R1131_U388, P2_R1131_U36, P2_U3398);
  nand ginst11843 (P2_R1131_U389, P2_R1131_U40, P2_U3063);
  not ginst11844 (P2_R1131_U39, P2_U3077);
  nand ginst11845 (P2_R1131_U390, P2_R1131_U388, P2_R1131_U389);
  nand ginst11846 (P2_R1131_U391, P2_R1131_U34, P2_U3395);
  nand ginst11847 (P2_R1131_U392, P2_R1131_U37, P2_U3067);
  nand ginst11848 (P2_R1131_U393, P2_R1131_U243, P2_R1131_U50);
  nand ginst11849 (P2_R1131_U394, P2_R1131_U162, P2_R1131_U205);
  nand ginst11850 (P2_R1131_U395, P2_R1131_U164, P2_U3904);
  nand ginst11851 (P2_R1131_U396, P2_R1131_U163, P2_U3054);
  nand ginst11852 (P2_R1131_U397, P2_R1131_U395, P2_R1131_U396);
  nand ginst11853 (P2_R1131_U398, P2_R1131_U164, P2_U3904);
  nand ginst11854 (P2_R1131_U399, P2_R1131_U163, P2_U3054);
  not ginst11855 (P2_R1131_U40, P2_U3398);
  nand ginst11856 (P2_R1131_U400, P2_R1131_U397, P2_R1131_U51, P2_U3053);
  nand ginst11857 (P2_R1131_U401, P2_R1131_U16, P2_R1131_U92, P2_U3895);
  nand ginst11858 (P2_R1131_U402, P2_R1131_U92, P2_U3895);
  nand ginst11859 (P2_R1131_U403, P2_R1131_U51, P2_U3053);
  not ginst11860 (P2_R1131_U404, P2_R1131_U138);
  nand ginst11861 (P2_R1131_U405, P2_R1131_U361, P2_R1131_U404);
  nand ginst11862 (P2_R1131_U406, P2_R1131_U138, P2_R1131_U166);
  nand ginst11863 (P2_R1131_U407, P2_R1131_U54, P2_U3896);
  nand ginst11864 (P2_R1131_U408, P2_R1131_U91, P2_U3052);
  nand ginst11865 (P2_R1131_U409, P2_R1131_U54, P2_U3896);
  not ginst11866 (P2_R1131_U41, P2_U3070);
  nand ginst11867 (P2_R1131_U410, P2_R1131_U91, P2_U3052);
  nand ginst11868 (P2_R1131_U411, P2_R1131_U409, P2_R1131_U410);
  nand ginst11869 (P2_R1131_U412, P2_R1131_U52, P2_U3897);
  nand ginst11870 (P2_R1131_U413, P2_R1131_U90, P2_U3056);
  nand ginst11871 (P2_R1131_U414, P2_R1131_U306, P2_R1131_U93);
  nand ginst11872 (P2_R1131_U415, P2_R1131_U167, P2_R1131_U298);
  nand ginst11873 (P2_R1131_U416, P2_R1131_U89, P2_U3898);
  nand ginst11874 (P2_R1131_U417, P2_R1131_U88, P2_U3057);
  not ginst11875 (P2_R1131_U418, P2_R1131_U141);
  nand ginst11876 (P2_R1131_U419, P2_R1131_U294, P2_R1131_U418);
  not ginst11877 (P2_R1131_U42, P2_U3066);
  nand ginst11878 (P2_R1131_U420, P2_R1131_U141, P2_R1131_U168);
  nand ginst11879 (P2_R1131_U421, P2_R1131_U87, P2_U3899);
  nand ginst11880 (P2_R1131_U422, P2_R1131_U86, P2_U3064);
  not ginst11881 (P2_R1131_U423, P2_R1131_U142);
  nand ginst11882 (P2_R1131_U424, P2_R1131_U290, P2_R1131_U423);
  nand ginst11883 (P2_R1131_U425, P2_R1131_U142, P2_R1131_U169);
  nand ginst11884 (P2_R1131_U426, P2_R1131_U82, P2_U3900);
  nand ginst11885 (P2_R1131_U427, P2_R1131_U79, P2_U3065);
  nand ginst11886 (P2_R1131_U428, P2_R1131_U426, P2_R1131_U427);
  nand ginst11887 (P2_R1131_U429, P2_R1131_U83, P2_U3901);
  not ginst11888 (P2_R1131_U43, P2_U3059);
  nand ginst11889 (P2_R1131_U430, P2_R1131_U80, P2_U3060);
  nand ginst11890 (P2_R1131_U431, P2_R1131_U316, P2_R1131_U94);
  nand ginst11891 (P2_R1131_U432, P2_R1131_U170, P2_R1131_U308);
  nand ginst11892 (P2_R1131_U433, P2_R1131_U84, P2_U3902);
  nand ginst11893 (P2_R1131_U434, P2_R1131_U81, P2_U3074);
  nand ginst11894 (P2_R1131_U435, P2_R1131_U172, P2_R1131_U317);
  nand ginst11895 (P2_R1131_U436, P2_R1131_U171, P2_R1131_U280);
  nand ginst11896 (P2_R1131_U437, P2_R1131_U78, P2_U3903);
  nand ginst11897 (P2_R1131_U438, P2_R1131_U77, P2_U3075);
  not ginst11898 (P2_R1131_U439, P2_R1131_U145);
  nand ginst11899 (P2_R1131_U44, P2_R1131_U31, P2_U3059);
  nand ginst11900 (P2_R1131_U440, P2_R1131_U276, P2_R1131_U439);
  nand ginst11901 (P2_R1131_U441, P2_R1131_U145, P2_R1131_U173);
  nand ginst11902 (P2_R1131_U442, P2_R1131_U39, P2_U3392);
  nand ginst11903 (P2_R1131_U443, P2_R1131_U174, P2_U3077);
  not ginst11904 (P2_R1131_U444, P2_R1131_U146);
  nand ginst11905 (P2_R1131_U445, P2_R1131_U203, P2_R1131_U444);
  nand ginst11906 (P2_R1131_U446, P2_R1131_U146, P2_R1131_U175);
  nand ginst11907 (P2_R1131_U447, P2_R1131_U76, P2_U3445);
  nand ginst11908 (P2_R1131_U448, P2_R1131_U75, P2_U3080);
  not ginst11909 (P2_R1131_U449, P2_R1131_U147);
  nand ginst11910 (P2_R1131_U45, P2_R1131_U214, P2_R1131_U216);
  nand ginst11911 (P2_R1131_U450, P2_R1131_U272, P2_R1131_U449);
  nand ginst11912 (P2_R1131_U451, P2_R1131_U147, P2_R1131_U176);
  nand ginst11913 (P2_R1131_U452, P2_R1131_U74, P2_U3443);
  nand ginst11914 (P2_R1131_U453, P2_R1131_U177, P2_U3081);
  not ginst11915 (P2_R1131_U454, P2_R1131_U148);
  nand ginst11916 (P2_R1131_U455, P2_R1131_U270, P2_R1131_U454);
  nand ginst11917 (P2_R1131_U456, P2_R1131_U148, P2_R1131_U178);
  nand ginst11918 (P2_R1131_U457, P2_R1131_U73, P2_U3440);
  nand ginst11919 (P2_R1131_U458, P2_R1131_U72, P2_U3068);
  not ginst11920 (P2_R1131_U459, P2_R1131_U149);
  not ginst11921 (P2_R1131_U46, P2_U3416);
  nand ginst11922 (P2_R1131_U460, P2_R1131_U266, P2_R1131_U459);
  nand ginst11923 (P2_R1131_U461, P2_R1131_U149, P2_R1131_U179);
  nand ginst11924 (P2_R1131_U462, P2_R1131_U68, P2_U3437);
  nand ginst11925 (P2_R1131_U463, P2_R1131_U65, P2_U3072);
  nand ginst11926 (P2_R1131_U464, P2_R1131_U462, P2_R1131_U463);
  nand ginst11927 (P2_R1131_U465, P2_R1131_U69, P2_U3434);
  nand ginst11928 (P2_R1131_U466, P2_R1131_U66, P2_U3073);
  nand ginst11929 (P2_R1131_U467, P2_R1131_U327, P2_R1131_U95);
  nand ginst11930 (P2_R1131_U468, P2_R1131_U180, P2_R1131_U319);
  nand ginst11931 (P2_R1131_U469, P2_R1131_U70, P2_U3431);
  not ginst11932 (P2_R1131_U47, P2_U3082);
  nand ginst11933 (P2_R1131_U470, P2_R1131_U67, P2_U3078);
  nand ginst11934 (P2_R1131_U471, P2_R1131_U182, P2_R1131_U328);
  nand ginst11935 (P2_R1131_U472, P2_R1131_U181, P2_R1131_U256);
  nand ginst11936 (P2_R1131_U473, P2_R1131_U64, P2_U3428);
  nand ginst11937 (P2_R1131_U474, P2_R1131_U63, P2_U3079);
  not ginst11938 (P2_R1131_U475, P2_R1131_U152);
  nand ginst11939 (P2_R1131_U476, P2_R1131_U354, P2_R1131_U475);
  nand ginst11940 (P2_R1131_U477, P2_R1131_U152, P2_R1131_U183);
  nand ginst11941 (P2_R1131_U478, P2_R1131_U55, P2_U3425);
  nand ginst11942 (P2_R1131_U479, P2_R1131_U61, P2_U3071);
  nand ginst11943 (P2_R1131_U48, P2_R1131_U217, P2_R1131_U45);
  not ginst11944 (P2_R1131_U480, P2_R1131_U153);
  nand ginst11945 (P2_R1131_U481, P2_R1131_U352, P2_R1131_U480);
  nand ginst11946 (P2_R1131_U482, P2_R1131_U153, P2_R1131_U184);
  nand ginst11947 (P2_R1131_U483, P2_R1131_U56, P2_U3422);
  nand ginst11948 (P2_R1131_U484, P2_R1131_U60, P2_U3062);
  nand ginst11949 (P2_R1131_U485, P2_R1131_U483, P2_R1131_U484);
  nand ginst11950 (P2_R1131_U486, P2_R1131_U57, P2_U3419);
  nand ginst11951 (P2_R1131_U487, P2_R1131_U58, P2_U3061);
  nand ginst11952 (P2_R1131_U488, P2_R1131_U336, P2_R1131_U96);
  nand ginst11953 (P2_R1131_U489, P2_R1131_U185, P2_R1131_U350);
  nand ginst11954 (P2_R1131_U49, P2_R1131_U231, P2_R1131_U44);
  nand ginst11955 (P2_R1131_U50, P2_R1131_U188, P2_R1131_U204, P2_R1131_U338);
  not ginst11956 (P2_R1131_U51, P2_U3895);
  not ginst11957 (P2_R1131_U52, P2_U3056);
  nand ginst11958 (P2_R1131_U53, P2_R1131_U90, P2_U3056);
  not ginst11959 (P2_R1131_U54, P2_U3052);
  not ginst11960 (P2_R1131_U55, P2_U3071);
  not ginst11961 (P2_R1131_U56, P2_U3062);
  not ginst11962 (P2_R1131_U57, P2_U3061);
  not ginst11963 (P2_R1131_U58, P2_U3419);
  nand ginst11964 (P2_R1131_U59, P2_R1131_U46, P2_U3082);
  and ginst11965 (P2_R1131_U6, P2_R1131_U211, P2_R1131_U212);
  not ginst11966 (P2_R1131_U60, P2_U3422);
  not ginst11967 (P2_R1131_U61, P2_U3425);
  nand ginst11968 (P2_R1131_U62, P2_R1131_U248, P2_R1131_U249);
  not ginst11969 (P2_R1131_U63, P2_U3428);
  not ginst11970 (P2_R1131_U64, P2_U3079);
  not ginst11971 (P2_R1131_U65, P2_U3437);
  not ginst11972 (P2_R1131_U66, P2_U3434);
  not ginst11973 (P2_R1131_U67, P2_U3431);
  not ginst11974 (P2_R1131_U68, P2_U3072);
  not ginst11975 (P2_R1131_U69, P2_U3073);
  and ginst11976 (P2_R1131_U7, P2_R1131_U245, P2_R1131_U246);
  not ginst11977 (P2_R1131_U70, P2_U3078);
  nand ginst11978 (P2_R1131_U71, P2_R1131_U67, P2_U3078);
  not ginst11979 (P2_R1131_U72, P2_U3440);
  not ginst11980 (P2_R1131_U73, P2_U3068);
  not ginst11981 (P2_R1131_U74, P2_U3081);
  not ginst11982 (P2_R1131_U75, P2_U3445);
  not ginst11983 (P2_R1131_U76, P2_U3080);
  not ginst11984 (P2_R1131_U77, P2_U3903);
  not ginst11985 (P2_R1131_U78, P2_U3075);
  not ginst11986 (P2_R1131_U79, P2_U3900);
  and ginst11987 (P2_R1131_U8, P2_R1131_U193, P2_R1131_U257);
  not ginst11988 (P2_R1131_U80, P2_U3901);
  not ginst11989 (P2_R1131_U81, P2_U3902);
  not ginst11990 (P2_R1131_U82, P2_U3065);
  not ginst11991 (P2_R1131_U83, P2_U3060);
  not ginst11992 (P2_R1131_U84, P2_U3074);
  nand ginst11993 (P2_R1131_U85, P2_R1131_U81, P2_U3074);
  not ginst11994 (P2_R1131_U86, P2_U3899);
  not ginst11995 (P2_R1131_U87, P2_U3064);
  not ginst11996 (P2_R1131_U88, P2_U3898);
  not ginst11997 (P2_R1131_U89, P2_U3057);
  and ginst11998 (P2_R1131_U9, P2_R1131_U258, P2_R1131_U259);
  not ginst11999 (P2_R1131_U90, P2_U3897);
  not ginst12000 (P2_R1131_U91, P2_U3896);
  not ginst12001 (P2_R1131_U92, P2_U3053);
  nand ginst12002 (P2_R1131_U93, P2_R1131_U296, P2_R1131_U297);
  nand ginst12003 (P2_R1131_U94, P2_R1131_U307, P2_R1131_U85);
  nand ginst12004 (P2_R1131_U95, P2_R1131_U318, P2_R1131_U71);
  nand ginst12005 (P2_R1131_U96, P2_R1131_U349, P2_R1131_U59);
  not ginst12006 (P2_R1131_U97, P2_U3076);
  nand ginst12007 (P2_R1131_U98, P2_R1131_U405, P2_R1131_U406);
  nand ginst12008 (P2_R1131_U99, P2_R1131_U419, P2_R1131_U420);
  and ginst12009 (P2_R1143_U10, P2_R1143_U348, P2_R1143_U351);
  nand ginst12010 (P2_R1143_U100, P2_R1143_U398, P2_R1143_U399);
  nand ginst12011 (P2_R1143_U101, P2_R1143_U407, P2_R1143_U408);
  nand ginst12012 (P2_R1143_U102, P2_R1143_U414, P2_R1143_U415);
  nand ginst12013 (P2_R1143_U103, P2_R1143_U421, P2_R1143_U422);
  nand ginst12014 (P2_R1143_U104, P2_R1143_U428, P2_R1143_U429);
  nand ginst12015 (P2_R1143_U105, P2_R1143_U433, P2_R1143_U434);
  nand ginst12016 (P2_R1143_U106, P2_R1143_U440, P2_R1143_U441);
  nand ginst12017 (P2_R1143_U107, P2_R1143_U447, P2_R1143_U448);
  nand ginst12018 (P2_R1143_U108, P2_R1143_U461, P2_R1143_U462);
  nand ginst12019 (P2_R1143_U109, P2_R1143_U466, P2_R1143_U467);
  and ginst12020 (P2_R1143_U11, P2_R1143_U341, P2_R1143_U344);
  nand ginst12021 (P2_R1143_U110, P2_R1143_U473, P2_R1143_U474);
  nand ginst12022 (P2_R1143_U111, P2_R1143_U480, P2_R1143_U481);
  nand ginst12023 (P2_R1143_U112, P2_R1143_U487, P2_R1143_U488);
  nand ginst12024 (P2_R1143_U113, P2_R1143_U494, P2_R1143_U495);
  nand ginst12025 (P2_R1143_U114, P2_R1143_U499, P2_R1143_U500);
  and ginst12026 (P2_R1143_U115, P2_R1143_U187, P2_R1143_U189);
  and ginst12027 (P2_R1143_U116, P2_R1143_U180, P2_R1143_U4);
  and ginst12028 (P2_R1143_U117, P2_R1143_U192, P2_R1143_U194);
  and ginst12029 (P2_R1143_U118, P2_R1143_U200, P2_R1143_U201);
  and ginst12030 (P2_R1143_U119, P2_R1143_U22, P2_R1143_U381, P2_R1143_U382);
  and ginst12031 (P2_R1143_U12, P2_R1143_U332, P2_R1143_U335);
  and ginst12032 (P2_R1143_U120, P2_R1143_U212, P2_R1143_U5);
  and ginst12033 (P2_R1143_U121, P2_R1143_U180, P2_R1143_U181);
  and ginst12034 (P2_R1143_U122, P2_R1143_U218, P2_R1143_U220);
  and ginst12035 (P2_R1143_U123, P2_R1143_U34, P2_R1143_U388, P2_R1143_U389);
  and ginst12036 (P2_R1143_U124, P2_R1143_U226, P2_R1143_U4);
  and ginst12037 (P2_R1143_U125, P2_R1143_U181, P2_R1143_U234);
  and ginst12038 (P2_R1143_U126, P2_R1143_U204, P2_R1143_U6);
  and ginst12039 (P2_R1143_U127, P2_R1143_U239, P2_R1143_U243);
  and ginst12040 (P2_R1143_U128, P2_R1143_U250, P2_R1143_U7);
  and ginst12041 (P2_R1143_U129, P2_R1143_U248, P2_R1143_U253);
  and ginst12042 (P2_R1143_U13, P2_R1143_U323, P2_R1143_U326);
  and ginst12043 (P2_R1143_U130, P2_R1143_U267, P2_R1143_U268);
  and ginst12044 (P2_R1143_U131, P2_R1143_U282, P2_R1143_U9);
  and ginst12045 (P2_R1143_U132, P2_R1143_U280, P2_R1143_U285);
  and ginst12046 (P2_R1143_U133, P2_R1143_U298, P2_R1143_U301);
  and ginst12047 (P2_R1143_U134, P2_R1143_U302, P2_R1143_U368);
  and ginst12048 (P2_R1143_U135, P2_R1143_U160, P2_R1143_U278);
  and ginst12049 (P2_R1143_U136, P2_R1143_U454, P2_R1143_U455, P2_R1143_U80);
  and ginst12050 (P2_R1143_U137, P2_R1143_U325, P2_R1143_U9);
  and ginst12051 (P2_R1143_U138, P2_R1143_U468, P2_R1143_U469, P2_R1143_U59);
  and ginst12052 (P2_R1143_U139, P2_R1143_U334, P2_R1143_U8);
  and ginst12053 (P2_R1143_U14, P2_R1143_U318, P2_R1143_U320);
  and ginst12054 (P2_R1143_U140, P2_R1143_U172, P2_R1143_U489, P2_R1143_U490);
  and ginst12055 (P2_R1143_U141, P2_R1143_U343, P2_R1143_U7);
  and ginst12056 (P2_R1143_U142, P2_R1143_U171, P2_R1143_U501, P2_R1143_U502);
  and ginst12057 (P2_R1143_U143, P2_R1143_U350, P2_R1143_U6);
  nand ginst12058 (P2_R1143_U144, P2_R1143_U118, P2_R1143_U202);
  nand ginst12059 (P2_R1143_U145, P2_R1143_U217, P2_R1143_U229);
  not ginst12060 (P2_R1143_U146, P2_U3054);
  not ginst12061 (P2_R1143_U147, P2_U3904);
  and ginst12062 (P2_R1143_U148, P2_R1143_U402, P2_R1143_U403);
  nand ginst12063 (P2_R1143_U149, P2_R1143_U169, P2_R1143_U304, P2_R1143_U364);
  and ginst12064 (P2_R1143_U15, P2_R1143_U310, P2_R1143_U313);
  and ginst12065 (P2_R1143_U150, P2_R1143_U409, P2_R1143_U410);
  nand ginst12066 (P2_R1143_U151, P2_R1143_U134, P2_R1143_U369, P2_R1143_U370);
  and ginst12067 (P2_R1143_U152, P2_R1143_U416, P2_R1143_U417);
  nand ginst12068 (P2_R1143_U153, P2_R1143_U299, P2_R1143_U365, P2_R1143_U86);
  and ginst12069 (P2_R1143_U154, P2_R1143_U423, P2_R1143_U424);
  nand ginst12070 (P2_R1143_U155, P2_R1143_U292, P2_R1143_U293);
  and ginst12071 (P2_R1143_U156, P2_R1143_U435, P2_R1143_U436);
  nand ginst12072 (P2_R1143_U157, P2_R1143_U288, P2_R1143_U289);
  and ginst12073 (P2_R1143_U158, P2_R1143_U442, P2_R1143_U443);
  nand ginst12074 (P2_R1143_U159, P2_R1143_U132, P2_R1143_U284);
  and ginst12075 (P2_R1143_U16, P2_R1143_U232, P2_R1143_U235);
  and ginst12076 (P2_R1143_U160, P2_R1143_U449, P2_R1143_U450);
  nand ginst12077 (P2_R1143_U161, P2_R1143_U327, P2_R1143_U43);
  nand ginst12078 (P2_R1143_U162, P2_R1143_U130, P2_R1143_U269);
  and ginst12079 (P2_R1143_U163, P2_R1143_U475, P2_R1143_U476);
  nand ginst12080 (P2_R1143_U164, P2_R1143_U256, P2_R1143_U257);
  and ginst12081 (P2_R1143_U165, P2_R1143_U482, P2_R1143_U483);
  nand ginst12082 (P2_R1143_U166, P2_R1143_U129, P2_R1143_U252);
  nand ginst12083 (P2_R1143_U167, P2_R1143_U127, P2_R1143_U242);
  nand ginst12084 (P2_R1143_U168, P2_R1143_U366, P2_R1143_U367);
  nand ginst12085 (P2_R1143_U169, P2_R1143_U151, P2_U3053);
  and ginst12086 (P2_R1143_U17, P2_R1143_U224, P2_R1143_U227);
  not ginst12087 (P2_R1143_U170, P2_R1143_U34);
  nand ginst12088 (P2_R1143_U171, P2_U3082, P2_U3416);
  nand ginst12089 (P2_R1143_U172, P2_U3071, P2_U3425);
  nand ginst12090 (P2_R1143_U173, P2_U3057, P2_U3898);
  not ginst12091 (P2_R1143_U174, P2_R1143_U68);
  not ginst12092 (P2_R1143_U175, P2_R1143_U77);
  nand ginst12093 (P2_R1143_U176, P2_U3064, P2_U3899);
  not ginst12094 (P2_R1143_U177, P2_R1143_U65);
  or ginst12095 (P2_R1143_U178, P2_U3066, P2_U3404);
  or ginst12096 (P2_R1143_U179, P2_U3059, P2_U3401);
  and ginst12097 (P2_R1143_U18, P2_R1143_U210, P2_R1143_U213);
  or ginst12098 (P2_R1143_U180, P2_U3063, P2_U3398);
  or ginst12099 (P2_R1143_U181, P2_U3067, P2_U3395);
  not ginst12100 (P2_R1143_U182, P2_R1143_U31);
  or ginst12101 (P2_R1143_U183, P2_U3077, P2_U3392);
  not ginst12102 (P2_R1143_U184, P2_R1143_U42);
  not ginst12103 (P2_R1143_U185, P2_R1143_U43);
  nand ginst12104 (P2_R1143_U186, P2_R1143_U42, P2_R1143_U43);
  nand ginst12105 (P2_R1143_U187, P2_U3067, P2_U3395);
  nand ginst12106 (P2_R1143_U188, P2_R1143_U181, P2_R1143_U186);
  nand ginst12107 (P2_R1143_U189, P2_U3063, P2_U3398);
  not ginst12108 (P2_R1143_U19, P2_U3407);
  nand ginst12109 (P2_R1143_U190, P2_R1143_U115, P2_R1143_U188);
  nand ginst12110 (P2_R1143_U191, P2_R1143_U34, P2_R1143_U35);
  nand ginst12111 (P2_R1143_U192, P2_R1143_U191, P2_U3066);
  nand ginst12112 (P2_R1143_U193, P2_R1143_U116, P2_R1143_U190);
  nand ginst12113 (P2_R1143_U194, P2_R1143_U170, P2_U3404);
  not ginst12114 (P2_R1143_U195, P2_R1143_U41);
  or ginst12115 (P2_R1143_U196, P2_U3069, P2_U3410);
  or ginst12116 (P2_R1143_U197, P2_U3070, P2_U3407);
  not ginst12117 (P2_R1143_U198, P2_R1143_U22);
  nand ginst12118 (P2_R1143_U199, P2_R1143_U22, P2_R1143_U23);
  not ginst12119 (P2_R1143_U20, P2_U3070);
  nand ginst12120 (P2_R1143_U200, P2_R1143_U199, P2_U3069);
  nand ginst12121 (P2_R1143_U201, P2_R1143_U198, P2_U3410);
  nand ginst12122 (P2_R1143_U202, P2_R1143_U41, P2_R1143_U5);
  not ginst12123 (P2_R1143_U203, P2_R1143_U144);
  or ginst12124 (P2_R1143_U204, P2_U3083, P2_U3413);
  nand ginst12125 (P2_R1143_U205, P2_R1143_U144, P2_R1143_U204);
  not ginst12126 (P2_R1143_U206, P2_R1143_U40);
  or ginst12127 (P2_R1143_U207, P2_U3082, P2_U3416);
  or ginst12128 (P2_R1143_U208, P2_U3070, P2_U3407);
  nand ginst12129 (P2_R1143_U209, P2_R1143_U208, P2_R1143_U41);
  not ginst12130 (P2_R1143_U21, P2_U3069);
  nand ginst12131 (P2_R1143_U210, P2_R1143_U119, P2_R1143_U209);
  nand ginst12132 (P2_R1143_U211, P2_R1143_U195, P2_R1143_U22);
  nand ginst12133 (P2_R1143_U212, P2_U3069, P2_U3410);
  nand ginst12134 (P2_R1143_U213, P2_R1143_U120, P2_R1143_U211);
  or ginst12135 (P2_R1143_U214, P2_U3070, P2_U3407);
  nand ginst12136 (P2_R1143_U215, P2_R1143_U181, P2_R1143_U185);
  nand ginst12137 (P2_R1143_U216, P2_U3067, P2_U3395);
  not ginst12138 (P2_R1143_U217, P2_R1143_U45);
  nand ginst12139 (P2_R1143_U218, P2_R1143_U121, P2_R1143_U184);
  nand ginst12140 (P2_R1143_U219, P2_R1143_U180, P2_R1143_U45);
  nand ginst12141 (P2_R1143_U22, P2_U3070, P2_U3407);
  nand ginst12142 (P2_R1143_U220, P2_U3063, P2_U3398);
  not ginst12143 (P2_R1143_U221, P2_R1143_U44);
  or ginst12144 (P2_R1143_U222, P2_U3059, P2_U3401);
  nand ginst12145 (P2_R1143_U223, P2_R1143_U222, P2_R1143_U44);
  nand ginst12146 (P2_R1143_U224, P2_R1143_U123, P2_R1143_U223);
  nand ginst12147 (P2_R1143_U225, P2_R1143_U221, P2_R1143_U34);
  nand ginst12148 (P2_R1143_U226, P2_U3066, P2_U3404);
  nand ginst12149 (P2_R1143_U227, P2_R1143_U124, P2_R1143_U225);
  or ginst12150 (P2_R1143_U228, P2_U3059, P2_U3401);
  nand ginst12151 (P2_R1143_U229, P2_R1143_U181, P2_R1143_U184);
  not ginst12152 (P2_R1143_U23, P2_U3410);
  not ginst12153 (P2_R1143_U230, P2_R1143_U145);
  nand ginst12154 (P2_R1143_U231, P2_U3063, P2_U3398);
  nand ginst12155 (P2_R1143_U232, P2_R1143_U400, P2_R1143_U401, P2_R1143_U42, P2_R1143_U43);
  nand ginst12156 (P2_R1143_U233, P2_R1143_U42, P2_R1143_U43);
  nand ginst12157 (P2_R1143_U234, P2_U3067, P2_U3395);
  nand ginst12158 (P2_R1143_U235, P2_R1143_U125, P2_R1143_U233);
  or ginst12159 (P2_R1143_U236, P2_U3082, P2_U3416);
  or ginst12160 (P2_R1143_U237, P2_U3061, P2_U3419);
  nand ginst12161 (P2_R1143_U238, P2_R1143_U177, P2_R1143_U6);
  nand ginst12162 (P2_R1143_U239, P2_U3061, P2_U3419);
  not ginst12163 (P2_R1143_U24, P2_U3401);
  nand ginst12164 (P2_R1143_U240, P2_R1143_U171, P2_R1143_U238);
  or ginst12165 (P2_R1143_U241, P2_U3061, P2_U3419);
  nand ginst12166 (P2_R1143_U242, P2_R1143_U126, P2_R1143_U144);
  nand ginst12167 (P2_R1143_U243, P2_R1143_U240, P2_R1143_U241);
  not ginst12168 (P2_R1143_U244, P2_R1143_U167);
  or ginst12169 (P2_R1143_U245, P2_U3079, P2_U3428);
  or ginst12170 (P2_R1143_U246, P2_U3071, P2_U3425);
  nand ginst12171 (P2_R1143_U247, P2_R1143_U174, P2_R1143_U7);
  nand ginst12172 (P2_R1143_U248, P2_U3079, P2_U3428);
  nand ginst12173 (P2_R1143_U249, P2_R1143_U172, P2_R1143_U247);
  not ginst12174 (P2_R1143_U25, P2_U3059);
  or ginst12175 (P2_R1143_U250, P2_U3062, P2_U3422);
  or ginst12176 (P2_R1143_U251, P2_U3079, P2_U3428);
  nand ginst12177 (P2_R1143_U252, P2_R1143_U128, P2_R1143_U167);
  nand ginst12178 (P2_R1143_U253, P2_R1143_U249, P2_R1143_U251);
  not ginst12179 (P2_R1143_U254, P2_R1143_U166);
  or ginst12180 (P2_R1143_U255, P2_U3078, P2_U3431);
  nand ginst12181 (P2_R1143_U256, P2_R1143_U166, P2_R1143_U255);
  nand ginst12182 (P2_R1143_U257, P2_U3078, P2_U3431);
  not ginst12183 (P2_R1143_U258, P2_R1143_U164);
  or ginst12184 (P2_R1143_U259, P2_U3073, P2_U3434);
  not ginst12185 (P2_R1143_U26, P2_U3066);
  nand ginst12186 (P2_R1143_U260, P2_R1143_U164, P2_R1143_U259);
  nand ginst12187 (P2_R1143_U261, P2_U3073, P2_U3434);
  not ginst12188 (P2_R1143_U262, P2_R1143_U92);
  or ginst12189 (P2_R1143_U263, P2_U3068, P2_U3440);
  or ginst12190 (P2_R1143_U264, P2_U3072, P2_U3437);
  not ginst12191 (P2_R1143_U265, P2_R1143_U59);
  nand ginst12192 (P2_R1143_U266, P2_R1143_U59, P2_R1143_U60);
  nand ginst12193 (P2_R1143_U267, P2_R1143_U266, P2_U3068);
  nand ginst12194 (P2_R1143_U268, P2_R1143_U265, P2_U3440);
  nand ginst12195 (P2_R1143_U269, P2_R1143_U8, P2_R1143_U92);
  not ginst12196 (P2_R1143_U27, P2_U3395);
  not ginst12197 (P2_R1143_U270, P2_R1143_U162);
  or ginst12198 (P2_R1143_U271, P2_U3075, P2_U3903);
  or ginst12199 (P2_R1143_U272, P2_U3080, P2_U3445);
  or ginst12200 (P2_R1143_U273, P2_U3074, P2_U3902);
  not ginst12201 (P2_R1143_U274, P2_R1143_U80);
  nand ginst12202 (P2_R1143_U275, P2_R1143_U274, P2_U3903);
  nand ginst12203 (P2_R1143_U276, P2_R1143_U275, P2_R1143_U90);
  nand ginst12204 (P2_R1143_U277, P2_R1143_U80, P2_R1143_U81);
  nand ginst12205 (P2_R1143_U278, P2_R1143_U276, P2_R1143_U277);
  nand ginst12206 (P2_R1143_U279, P2_R1143_U175, P2_R1143_U9);
  not ginst12207 (P2_R1143_U28, P2_U3067);
  nand ginst12208 (P2_R1143_U280, P2_U3074, P2_U3902);
  nand ginst12209 (P2_R1143_U281, P2_R1143_U278, P2_R1143_U279);
  or ginst12210 (P2_R1143_U282, P2_U3081, P2_U3443);
  or ginst12211 (P2_R1143_U283, P2_U3074, P2_U3902);
  nand ginst12212 (P2_R1143_U284, P2_R1143_U131, P2_R1143_U162, P2_R1143_U273);
  nand ginst12213 (P2_R1143_U285, P2_R1143_U281, P2_R1143_U283);
  not ginst12214 (P2_R1143_U286, P2_R1143_U159);
  or ginst12215 (P2_R1143_U287, P2_U3060, P2_U3901);
  nand ginst12216 (P2_R1143_U288, P2_R1143_U159, P2_R1143_U287);
  nand ginst12217 (P2_R1143_U289, P2_U3060, P2_U3901);
  not ginst12218 (P2_R1143_U29, P2_U3387);
  not ginst12219 (P2_R1143_U290, P2_R1143_U157);
  or ginst12220 (P2_R1143_U291, P2_U3065, P2_U3900);
  nand ginst12221 (P2_R1143_U292, P2_R1143_U157, P2_R1143_U291);
  nand ginst12222 (P2_R1143_U293, P2_U3065, P2_U3900);
  not ginst12223 (P2_R1143_U294, P2_R1143_U155);
  or ginst12224 (P2_R1143_U295, P2_U3057, P2_U3898);
  nand ginst12225 (P2_R1143_U296, P2_R1143_U173, P2_R1143_U176);
  not ginst12226 (P2_R1143_U297, P2_R1143_U86);
  or ginst12227 (P2_R1143_U298, P2_U3064, P2_U3899);
  nand ginst12228 (P2_R1143_U299, P2_R1143_U155, P2_R1143_U168, P2_R1143_U298);
  not ginst12229 (P2_R1143_U30, P2_U3076);
  not ginst12230 (P2_R1143_U300, P2_R1143_U153);
  or ginst12231 (P2_R1143_U301, P2_U3052, P2_U3896);
  nand ginst12232 (P2_R1143_U302, P2_U3052, P2_U3896);
  not ginst12233 (P2_R1143_U303, P2_R1143_U151);
  nand ginst12234 (P2_R1143_U304, P2_R1143_U151, P2_U3895);
  not ginst12235 (P2_R1143_U305, P2_R1143_U149);
  nand ginst12236 (P2_R1143_U306, P2_R1143_U155, P2_R1143_U298);
  not ginst12237 (P2_R1143_U307, P2_R1143_U89);
  or ginst12238 (P2_R1143_U308, P2_U3057, P2_U3898);
  nand ginst12239 (P2_R1143_U309, P2_R1143_U308, P2_R1143_U89);
  nand ginst12240 (P2_R1143_U31, P2_U3076, P2_U3387);
  nand ginst12241 (P2_R1143_U310, P2_R1143_U154, P2_R1143_U173, P2_R1143_U309);
  nand ginst12242 (P2_R1143_U311, P2_R1143_U173, P2_R1143_U307);
  nand ginst12243 (P2_R1143_U312, P2_U3056, P2_U3897);
  nand ginst12244 (P2_R1143_U313, P2_R1143_U168, P2_R1143_U311, P2_R1143_U312);
  or ginst12245 (P2_R1143_U314, P2_U3057, P2_U3898);
  nand ginst12246 (P2_R1143_U315, P2_R1143_U162, P2_R1143_U282);
  not ginst12247 (P2_R1143_U316, P2_R1143_U91);
  nand ginst12248 (P2_R1143_U317, P2_R1143_U9, P2_R1143_U91);
  nand ginst12249 (P2_R1143_U318, P2_R1143_U135, P2_R1143_U317);
  nand ginst12250 (P2_R1143_U319, P2_R1143_U278, P2_R1143_U317);
  not ginst12251 (P2_R1143_U32, P2_U3398);
  nand ginst12252 (P2_R1143_U320, P2_R1143_U319, P2_R1143_U453);
  or ginst12253 (P2_R1143_U321, P2_U3080, P2_U3445);
  nand ginst12254 (P2_R1143_U322, P2_R1143_U321, P2_R1143_U91);
  nand ginst12255 (P2_R1143_U323, P2_R1143_U136, P2_R1143_U322);
  nand ginst12256 (P2_R1143_U324, P2_R1143_U316, P2_R1143_U80);
  nand ginst12257 (P2_R1143_U325, P2_U3075, P2_U3903);
  nand ginst12258 (P2_R1143_U326, P2_R1143_U137, P2_R1143_U324);
  or ginst12259 (P2_R1143_U327, P2_U3077, P2_U3392);
  not ginst12260 (P2_R1143_U328, P2_R1143_U161);
  or ginst12261 (P2_R1143_U329, P2_U3080, P2_U3445);
  not ginst12262 (P2_R1143_U33, P2_U3063);
  or ginst12263 (P2_R1143_U330, P2_U3072, P2_U3437);
  nand ginst12264 (P2_R1143_U331, P2_R1143_U330, P2_R1143_U92);
  nand ginst12265 (P2_R1143_U332, P2_R1143_U138, P2_R1143_U331);
  nand ginst12266 (P2_R1143_U333, P2_R1143_U262, P2_R1143_U59);
  nand ginst12267 (P2_R1143_U334, P2_U3068, P2_U3440);
  nand ginst12268 (P2_R1143_U335, P2_R1143_U139, P2_R1143_U333);
  or ginst12269 (P2_R1143_U336, P2_U3072, P2_U3437);
  nand ginst12270 (P2_R1143_U337, P2_R1143_U167, P2_R1143_U250);
  not ginst12271 (P2_R1143_U338, P2_R1143_U93);
  or ginst12272 (P2_R1143_U339, P2_U3071, P2_U3425);
  nand ginst12273 (P2_R1143_U34, P2_U3059, P2_U3401);
  nand ginst12274 (P2_R1143_U340, P2_R1143_U339, P2_R1143_U93);
  nand ginst12275 (P2_R1143_U341, P2_R1143_U140, P2_R1143_U340);
  nand ginst12276 (P2_R1143_U342, P2_R1143_U172, P2_R1143_U338);
  nand ginst12277 (P2_R1143_U343, P2_U3079, P2_U3428);
  nand ginst12278 (P2_R1143_U344, P2_R1143_U141, P2_R1143_U342);
  or ginst12279 (P2_R1143_U345, P2_U3071, P2_U3425);
  or ginst12280 (P2_R1143_U346, P2_U3082, P2_U3416);
  nand ginst12281 (P2_R1143_U347, P2_R1143_U346, P2_R1143_U40);
  nand ginst12282 (P2_R1143_U348, P2_R1143_U142, P2_R1143_U347);
  nand ginst12283 (P2_R1143_U349, P2_R1143_U171, P2_R1143_U206);
  not ginst12284 (P2_R1143_U35, P2_U3404);
  nand ginst12285 (P2_R1143_U350, P2_U3061, P2_U3419);
  nand ginst12286 (P2_R1143_U351, P2_R1143_U143, P2_R1143_U349);
  nand ginst12287 (P2_R1143_U352, P2_R1143_U171, P2_R1143_U207);
  nand ginst12288 (P2_R1143_U353, P2_R1143_U204, P2_R1143_U65);
  nand ginst12289 (P2_R1143_U354, P2_R1143_U214, P2_R1143_U22);
  nand ginst12290 (P2_R1143_U355, P2_R1143_U228, P2_R1143_U34);
  nand ginst12291 (P2_R1143_U356, P2_R1143_U180, P2_R1143_U231);
  nand ginst12292 (P2_R1143_U357, P2_R1143_U173, P2_R1143_U314);
  nand ginst12293 (P2_R1143_U358, P2_R1143_U176, P2_R1143_U298);
  nand ginst12294 (P2_R1143_U359, P2_R1143_U329, P2_R1143_U80);
  not ginst12295 (P2_R1143_U36, P2_U3413);
  nand ginst12296 (P2_R1143_U360, P2_R1143_U282, P2_R1143_U77);
  nand ginst12297 (P2_R1143_U361, P2_R1143_U336, P2_R1143_U59);
  nand ginst12298 (P2_R1143_U362, P2_R1143_U172, P2_R1143_U345);
  nand ginst12299 (P2_R1143_U363, P2_R1143_U250, P2_R1143_U68);
  nand ginst12300 (P2_R1143_U364, P2_U3053, P2_U3895);
  nand ginst12301 (P2_R1143_U365, P2_R1143_U168, P2_R1143_U296);
  nand ginst12302 (P2_R1143_U366, P2_R1143_U295, P2_U3056);
  nand ginst12303 (P2_R1143_U367, P2_R1143_U295, P2_U3897);
  nand ginst12304 (P2_R1143_U368, P2_R1143_U168, P2_R1143_U296, P2_R1143_U301);
  nand ginst12305 (P2_R1143_U369, P2_R1143_U133, P2_R1143_U155, P2_R1143_U168);
  not ginst12306 (P2_R1143_U37, P2_U3083);
  nand ginst12307 (P2_R1143_U370, P2_R1143_U297, P2_R1143_U301);
  nand ginst12308 (P2_R1143_U371, P2_R1143_U39, P2_U3082);
  nand ginst12309 (P2_R1143_U372, P2_R1143_U38, P2_U3416);
  nand ginst12310 (P2_R1143_U373, P2_R1143_U371, P2_R1143_U372);
  nand ginst12311 (P2_R1143_U374, P2_R1143_U352, P2_R1143_U40);
  nand ginst12312 (P2_R1143_U375, P2_R1143_U206, P2_R1143_U373);
  nand ginst12313 (P2_R1143_U376, P2_R1143_U36, P2_U3083);
  nand ginst12314 (P2_R1143_U377, P2_R1143_U37, P2_U3413);
  nand ginst12315 (P2_R1143_U378, P2_R1143_U376, P2_R1143_U377);
  nand ginst12316 (P2_R1143_U379, P2_R1143_U144, P2_R1143_U353);
  not ginst12317 (P2_R1143_U38, P2_U3082);
  nand ginst12318 (P2_R1143_U380, P2_R1143_U203, P2_R1143_U378);
  nand ginst12319 (P2_R1143_U381, P2_R1143_U23, P2_U3069);
  nand ginst12320 (P2_R1143_U382, P2_R1143_U21, P2_U3410);
  nand ginst12321 (P2_R1143_U383, P2_R1143_U19, P2_U3070);
  nand ginst12322 (P2_R1143_U384, P2_R1143_U20, P2_U3407);
  nand ginst12323 (P2_R1143_U385, P2_R1143_U383, P2_R1143_U384);
  nand ginst12324 (P2_R1143_U386, P2_R1143_U354, P2_R1143_U41);
  nand ginst12325 (P2_R1143_U387, P2_R1143_U195, P2_R1143_U385);
  nand ginst12326 (P2_R1143_U388, P2_R1143_U35, P2_U3066);
  nand ginst12327 (P2_R1143_U389, P2_R1143_U26, P2_U3404);
  not ginst12328 (P2_R1143_U39, P2_U3416);
  nand ginst12329 (P2_R1143_U390, P2_R1143_U24, P2_U3059);
  nand ginst12330 (P2_R1143_U391, P2_R1143_U25, P2_U3401);
  nand ginst12331 (P2_R1143_U392, P2_R1143_U390, P2_R1143_U391);
  nand ginst12332 (P2_R1143_U393, P2_R1143_U355, P2_R1143_U44);
  nand ginst12333 (P2_R1143_U394, P2_R1143_U221, P2_R1143_U392);
  nand ginst12334 (P2_R1143_U395, P2_R1143_U32, P2_U3063);
  nand ginst12335 (P2_R1143_U396, P2_R1143_U33, P2_U3398);
  nand ginst12336 (P2_R1143_U397, P2_R1143_U395, P2_R1143_U396);
  nand ginst12337 (P2_R1143_U398, P2_R1143_U145, P2_R1143_U356);
  nand ginst12338 (P2_R1143_U399, P2_R1143_U230, P2_R1143_U397);
  and ginst12339 (P2_R1143_U4, P2_R1143_U178, P2_R1143_U179);
  nand ginst12340 (P2_R1143_U40, P2_R1143_U205, P2_R1143_U65);
  nand ginst12341 (P2_R1143_U400, P2_R1143_U27, P2_U3067);
  nand ginst12342 (P2_R1143_U401, P2_R1143_U28, P2_U3395);
  nand ginst12343 (P2_R1143_U402, P2_R1143_U147, P2_U3054);
  nand ginst12344 (P2_R1143_U403, P2_R1143_U146, P2_U3904);
  nand ginst12345 (P2_R1143_U404, P2_R1143_U147, P2_U3054);
  nand ginst12346 (P2_R1143_U405, P2_R1143_U146, P2_U3904);
  nand ginst12347 (P2_R1143_U406, P2_R1143_U404, P2_R1143_U405);
  nand ginst12348 (P2_R1143_U407, P2_R1143_U148, P2_R1143_U149);
  nand ginst12349 (P2_R1143_U408, P2_R1143_U305, P2_R1143_U406);
  nand ginst12350 (P2_R1143_U409, P2_R1143_U88, P2_U3053);
  nand ginst12351 (P2_R1143_U41, P2_R1143_U117, P2_R1143_U193);
  nand ginst12352 (P2_R1143_U410, P2_R1143_U87, P2_U3895);
  nand ginst12353 (P2_R1143_U411, P2_R1143_U88, P2_U3053);
  nand ginst12354 (P2_R1143_U412, P2_R1143_U87, P2_U3895);
  nand ginst12355 (P2_R1143_U413, P2_R1143_U411, P2_R1143_U412);
  nand ginst12356 (P2_R1143_U414, P2_R1143_U150, P2_R1143_U151);
  nand ginst12357 (P2_R1143_U415, P2_R1143_U303, P2_R1143_U413);
  nand ginst12358 (P2_R1143_U416, P2_R1143_U46, P2_U3052);
  nand ginst12359 (P2_R1143_U417, P2_R1143_U47, P2_U3896);
  nand ginst12360 (P2_R1143_U418, P2_R1143_U46, P2_U3052);
  nand ginst12361 (P2_R1143_U419, P2_R1143_U47, P2_U3896);
  nand ginst12362 (P2_R1143_U42, P2_R1143_U182, P2_R1143_U183);
  nand ginst12363 (P2_R1143_U420, P2_R1143_U418, P2_R1143_U419);
  nand ginst12364 (P2_R1143_U421, P2_R1143_U152, P2_R1143_U153);
  nand ginst12365 (P2_R1143_U422, P2_R1143_U300, P2_R1143_U420);
  nand ginst12366 (P2_R1143_U423, P2_R1143_U49, P2_U3056);
  nand ginst12367 (P2_R1143_U424, P2_R1143_U48, P2_U3897);
  nand ginst12368 (P2_R1143_U425, P2_R1143_U50, P2_U3057);
  nand ginst12369 (P2_R1143_U426, P2_R1143_U51, P2_U3898);
  nand ginst12370 (P2_R1143_U427, P2_R1143_U425, P2_R1143_U426);
  nand ginst12371 (P2_R1143_U428, P2_R1143_U357, P2_R1143_U89);
  nand ginst12372 (P2_R1143_U429, P2_R1143_U307, P2_R1143_U427);
  nand ginst12373 (P2_R1143_U43, P2_U3077, P2_U3392);
  nand ginst12374 (P2_R1143_U430, P2_R1143_U52, P2_U3064);
  nand ginst12375 (P2_R1143_U431, P2_R1143_U53, P2_U3899);
  nand ginst12376 (P2_R1143_U432, P2_R1143_U430, P2_R1143_U431);
  nand ginst12377 (P2_R1143_U433, P2_R1143_U155, P2_R1143_U358);
  nand ginst12378 (P2_R1143_U434, P2_R1143_U294, P2_R1143_U432);
  nand ginst12379 (P2_R1143_U435, P2_R1143_U84, P2_U3065);
  nand ginst12380 (P2_R1143_U436, P2_R1143_U85, P2_U3900);
  nand ginst12381 (P2_R1143_U437, P2_R1143_U84, P2_U3065);
  nand ginst12382 (P2_R1143_U438, P2_R1143_U85, P2_U3900);
  nand ginst12383 (P2_R1143_U439, P2_R1143_U437, P2_R1143_U438);
  nand ginst12384 (P2_R1143_U44, P2_R1143_U122, P2_R1143_U219);
  nand ginst12385 (P2_R1143_U440, P2_R1143_U156, P2_R1143_U157);
  nand ginst12386 (P2_R1143_U441, P2_R1143_U290, P2_R1143_U439);
  nand ginst12387 (P2_R1143_U442, P2_R1143_U82, P2_U3060);
  nand ginst12388 (P2_R1143_U443, P2_R1143_U83, P2_U3901);
  nand ginst12389 (P2_R1143_U444, P2_R1143_U82, P2_U3060);
  nand ginst12390 (P2_R1143_U445, P2_R1143_U83, P2_U3901);
  nand ginst12391 (P2_R1143_U446, P2_R1143_U444, P2_R1143_U445);
  nand ginst12392 (P2_R1143_U447, P2_R1143_U158, P2_R1143_U159);
  nand ginst12393 (P2_R1143_U448, P2_R1143_U286, P2_R1143_U446);
  nand ginst12394 (P2_R1143_U449, P2_R1143_U54, P2_U3074);
  nand ginst12395 (P2_R1143_U45, P2_R1143_U215, P2_R1143_U216);
  nand ginst12396 (P2_R1143_U450, P2_R1143_U55, P2_U3902);
  nand ginst12397 (P2_R1143_U451, P2_R1143_U54, P2_U3074);
  nand ginst12398 (P2_R1143_U452, P2_R1143_U55, P2_U3902);
  nand ginst12399 (P2_R1143_U453, P2_R1143_U451, P2_R1143_U452);
  nand ginst12400 (P2_R1143_U454, P2_R1143_U81, P2_U3075);
  nand ginst12401 (P2_R1143_U455, P2_R1143_U90, P2_U3903);
  nand ginst12402 (P2_R1143_U456, P2_R1143_U161, P2_R1143_U182);
  nand ginst12403 (P2_R1143_U457, P2_R1143_U31, P2_R1143_U328);
  nand ginst12404 (P2_R1143_U458, P2_R1143_U78, P2_U3080);
  nand ginst12405 (P2_R1143_U459, P2_R1143_U79, P2_U3445);
  not ginst12406 (P2_R1143_U46, P2_U3896);
  nand ginst12407 (P2_R1143_U460, P2_R1143_U458, P2_R1143_U459);
  nand ginst12408 (P2_R1143_U461, P2_R1143_U359, P2_R1143_U91);
  nand ginst12409 (P2_R1143_U462, P2_R1143_U316, P2_R1143_U460);
  nand ginst12410 (P2_R1143_U463, P2_R1143_U75, P2_U3081);
  nand ginst12411 (P2_R1143_U464, P2_R1143_U76, P2_U3443);
  nand ginst12412 (P2_R1143_U465, P2_R1143_U463, P2_R1143_U464);
  nand ginst12413 (P2_R1143_U466, P2_R1143_U162, P2_R1143_U360);
  nand ginst12414 (P2_R1143_U467, P2_R1143_U270, P2_R1143_U465);
  nand ginst12415 (P2_R1143_U468, P2_R1143_U60, P2_U3068);
  nand ginst12416 (P2_R1143_U469, P2_R1143_U58, P2_U3440);
  not ginst12417 (P2_R1143_U47, P2_U3052);
  nand ginst12418 (P2_R1143_U470, P2_R1143_U56, P2_U3072);
  nand ginst12419 (P2_R1143_U471, P2_R1143_U57, P2_U3437);
  nand ginst12420 (P2_R1143_U472, P2_R1143_U470, P2_R1143_U471);
  nand ginst12421 (P2_R1143_U473, P2_R1143_U361, P2_R1143_U92);
  nand ginst12422 (P2_R1143_U474, P2_R1143_U262, P2_R1143_U472);
  nand ginst12423 (P2_R1143_U475, P2_R1143_U73, P2_U3073);
  nand ginst12424 (P2_R1143_U476, P2_R1143_U74, P2_U3434);
  nand ginst12425 (P2_R1143_U477, P2_R1143_U73, P2_U3073);
  nand ginst12426 (P2_R1143_U478, P2_R1143_U74, P2_U3434);
  nand ginst12427 (P2_R1143_U479, P2_R1143_U477, P2_R1143_U478);
  not ginst12428 (P2_R1143_U48, P2_U3056);
  nand ginst12429 (P2_R1143_U480, P2_R1143_U163, P2_R1143_U164);
  nand ginst12430 (P2_R1143_U481, P2_R1143_U258, P2_R1143_U479);
  nand ginst12431 (P2_R1143_U482, P2_R1143_U71, P2_U3078);
  nand ginst12432 (P2_R1143_U483, P2_R1143_U72, P2_U3431);
  nand ginst12433 (P2_R1143_U484, P2_R1143_U71, P2_U3078);
  nand ginst12434 (P2_R1143_U485, P2_R1143_U72, P2_U3431);
  nand ginst12435 (P2_R1143_U486, P2_R1143_U484, P2_R1143_U485);
  nand ginst12436 (P2_R1143_U487, P2_R1143_U165, P2_R1143_U166);
  nand ginst12437 (P2_R1143_U488, P2_R1143_U254, P2_R1143_U486);
  nand ginst12438 (P2_R1143_U489, P2_R1143_U61, P2_U3079);
  not ginst12439 (P2_R1143_U49, P2_U3897);
  nand ginst12440 (P2_R1143_U490, P2_R1143_U62, P2_U3428);
  nand ginst12441 (P2_R1143_U491, P2_R1143_U69, P2_U3071);
  nand ginst12442 (P2_R1143_U492, P2_R1143_U70, P2_U3425);
  nand ginst12443 (P2_R1143_U493, P2_R1143_U491, P2_R1143_U492);
  nand ginst12444 (P2_R1143_U494, P2_R1143_U362, P2_R1143_U93);
  nand ginst12445 (P2_R1143_U495, P2_R1143_U338, P2_R1143_U493);
  nand ginst12446 (P2_R1143_U496, P2_R1143_U66, P2_U3062);
  nand ginst12447 (P2_R1143_U497, P2_R1143_U67, P2_U3422);
  nand ginst12448 (P2_R1143_U498, P2_R1143_U496, P2_R1143_U497);
  nand ginst12449 (P2_R1143_U499, P2_R1143_U167, P2_R1143_U363);
  and ginst12450 (P2_R1143_U5, P2_R1143_U196, P2_R1143_U197);
  not ginst12451 (P2_R1143_U50, P2_U3898);
  nand ginst12452 (P2_R1143_U500, P2_R1143_U244, P2_R1143_U498);
  nand ginst12453 (P2_R1143_U501, P2_R1143_U63, P2_U3061);
  nand ginst12454 (P2_R1143_U502, P2_R1143_U64, P2_U3419);
  nand ginst12455 (P2_R1143_U503, P2_R1143_U29, P2_U3076);
  nand ginst12456 (P2_R1143_U504, P2_R1143_U30, P2_U3387);
  not ginst12457 (P2_R1143_U51, P2_U3057);
  not ginst12458 (P2_R1143_U52, P2_U3899);
  not ginst12459 (P2_R1143_U53, P2_U3064);
  not ginst12460 (P2_R1143_U54, P2_U3902);
  not ginst12461 (P2_R1143_U55, P2_U3074);
  not ginst12462 (P2_R1143_U56, P2_U3437);
  not ginst12463 (P2_R1143_U57, P2_U3072);
  not ginst12464 (P2_R1143_U58, P2_U3068);
  nand ginst12465 (P2_R1143_U59, P2_U3072, P2_U3437);
  and ginst12466 (P2_R1143_U6, P2_R1143_U236, P2_R1143_U237);
  not ginst12467 (P2_R1143_U60, P2_U3440);
  not ginst12468 (P2_R1143_U61, P2_U3428);
  not ginst12469 (P2_R1143_U62, P2_U3079);
  not ginst12470 (P2_R1143_U63, P2_U3419);
  not ginst12471 (P2_R1143_U64, P2_U3061);
  nand ginst12472 (P2_R1143_U65, P2_U3083, P2_U3413);
  not ginst12473 (P2_R1143_U66, P2_U3422);
  not ginst12474 (P2_R1143_U67, P2_U3062);
  nand ginst12475 (P2_R1143_U68, P2_U3062, P2_U3422);
  not ginst12476 (P2_R1143_U69, P2_U3425);
  and ginst12477 (P2_R1143_U7, P2_R1143_U245, P2_R1143_U246);
  not ginst12478 (P2_R1143_U70, P2_U3071);
  not ginst12479 (P2_R1143_U71, P2_U3431);
  not ginst12480 (P2_R1143_U72, P2_U3078);
  not ginst12481 (P2_R1143_U73, P2_U3434);
  not ginst12482 (P2_R1143_U74, P2_U3073);
  not ginst12483 (P2_R1143_U75, P2_U3443);
  not ginst12484 (P2_R1143_U76, P2_U3081);
  nand ginst12485 (P2_R1143_U77, P2_U3081, P2_U3443);
  not ginst12486 (P2_R1143_U78, P2_U3445);
  not ginst12487 (P2_R1143_U79, P2_U3080);
  and ginst12488 (P2_R1143_U8, P2_R1143_U263, P2_R1143_U264);
  nand ginst12489 (P2_R1143_U80, P2_U3080, P2_U3445);
  not ginst12490 (P2_R1143_U81, P2_U3903);
  not ginst12491 (P2_R1143_U82, P2_U3901);
  not ginst12492 (P2_R1143_U83, P2_U3060);
  not ginst12493 (P2_R1143_U84, P2_U3900);
  not ginst12494 (P2_R1143_U85, P2_U3065);
  nand ginst12495 (P2_R1143_U86, P2_U3056, P2_U3897);
  not ginst12496 (P2_R1143_U87, P2_U3053);
  not ginst12497 (P2_R1143_U88, P2_U3895);
  nand ginst12498 (P2_R1143_U89, P2_R1143_U176, P2_R1143_U306);
  and ginst12499 (P2_R1143_U9, P2_R1143_U271, P2_R1143_U272);
  not ginst12500 (P2_R1143_U90, P2_U3075);
  nand ginst12501 (P2_R1143_U91, P2_R1143_U315, P2_R1143_U77);
  nand ginst12502 (P2_R1143_U92, P2_R1143_U260, P2_R1143_U261);
  nand ginst12503 (P2_R1143_U93, P2_R1143_U337, P2_R1143_U68);
  nand ginst12504 (P2_R1143_U94, P2_R1143_U456, P2_R1143_U457);
  nand ginst12505 (P2_R1143_U95, P2_R1143_U503, P2_R1143_U504);
  nand ginst12506 (P2_R1143_U96, P2_R1143_U374, P2_R1143_U375);
  nand ginst12507 (P2_R1143_U97, P2_R1143_U379, P2_R1143_U380);
  nand ginst12508 (P2_R1143_U98, P2_R1143_U386, P2_R1143_U387);
  nand ginst12509 (P2_R1143_U99, P2_R1143_U393, P2_R1143_U394);
  and ginst12510 (P2_R1158_U10, P2_R1158_U235, P2_R1158_U5);
  nand ginst12511 (P2_R1158_U100, P2_R1158_U451, P2_R1158_U452);
  nand ginst12512 (P2_R1158_U101, P2_R1158_U458, P2_R1158_U459);
  nand ginst12513 (P2_R1158_U102, P2_R1158_U465, P2_R1158_U466);
  nand ginst12514 (P2_R1158_U103, P2_R1158_U527, P2_R1158_U528);
  nand ginst12515 (P2_R1158_U104, P2_R1158_U534, P2_R1158_U535);
  nand ginst12516 (P2_R1158_U105, P2_R1158_U543, P2_R1158_U544);
  nand ginst12517 (P2_R1158_U106, P2_R1158_U548, P2_R1158_U549);
  nand ginst12518 (P2_R1158_U107, P2_R1158_U555, P2_R1158_U556);
  nand ginst12519 (P2_R1158_U108, P2_R1158_U562, P2_R1158_U563);
  nand ginst12520 (P2_R1158_U109, P2_R1158_U569, P2_R1158_U570);
  and ginst12521 (P2_R1158_U11, P2_R1158_U261, P2_R1158_U9);
  nand ginst12522 (P2_R1158_U110, P2_R1158_U576, P2_R1158_U577);
  nand ginst12523 (P2_R1158_U111, P2_R1158_U581, P2_R1158_U582);
  nand ginst12524 (P2_R1158_U112, P2_R1158_U588, P2_R1158_U589);
  nand ginst12525 (P2_R1158_U113, P2_R1158_U595, P2_R1158_U596);
  nand ginst12526 (P2_R1158_U114, P2_R1158_U602, P2_R1158_U603);
  nand ginst12527 (P2_R1158_U115, P2_R1158_U609, P2_R1158_U610);
  nand ginst12528 (P2_R1158_U116, P2_R1158_U616, P2_R1158_U617);
  nand ginst12529 (P2_R1158_U117, P2_R1158_U621, P2_R1158_U622);
  nand ginst12530 (P2_R1158_U118, P2_R1158_U628, P2_R1158_U629);
  and ginst12531 (P2_R1158_U119, P2_R1158_U75, P2_U3152);
  and ginst12532 (P2_R1158_U12, P2_R1158_U11, P2_R1158_U271);
  and ginst12533 (P2_R1158_U120, P2_R1158_U229, P2_R1158_U230);
  and ginst12534 (P2_R1158_U121, P2_R1158_U10, P2_R1158_U243);
  and ginst12535 (P2_R1158_U122, P2_R1158_U244, P2_R1158_U361);
  and ginst12536 (P2_R1158_U123, P2_R1158_U24, P2_R1158_U439, P2_R1158_U440);
  and ginst12537 (P2_R1158_U124, P2_R1158_U249, P2_R1158_U5);
  and ginst12538 (P2_R1158_U125, P2_R1158_U29, P2_R1158_U460, P2_R1158_U461);
  and ginst12539 (P2_R1158_U126, P2_R1158_U256, P2_R1158_U4);
  and ginst12540 (P2_R1158_U127, P2_R1158_U213, P2_R1158_U266);
  and ginst12541 (P2_R1158_U128, P2_R1158_U12, P2_R1158_U273);
  and ginst12542 (P2_R1158_U129, P2_R1158_U274, P2_R1158_U372);
  and ginst12543 (P2_R1158_U13, P2_R1158_U536, P2_R1158_U537);
  and ginst12544 (P2_R1158_U130, P2_R1158_U279, P2_R1158_U280);
  and ginst12545 (P2_R1158_U131, P2_R1158_U292, P2_R1158_U8);
  and ginst12546 (P2_R1158_U132, P2_R1158_U214, P2_R1158_U290);
  and ginst12547 (P2_R1158_U133, P2_R1158_U313, P2_R1158_U375);
  and ginst12548 (P2_R1158_U134, P2_R1158_U306, P2_R1158_U315);
  and ginst12549 (P2_R1158_U135, P2_R1158_U315, P2_R1158_U369);
  and ginst12550 (P2_R1158_U136, P2_R1158_U314, P2_R1158_U373);
  nand ginst12551 (P2_R1158_U137, P2_R1158_U521, P2_R1158_U522);
  and ginst12552 (P2_R1158_U138, P2_R1158_U215, P2_R1158_U318);
  and ginst12553 (P2_R1158_U139, P2_R1158_U39, P2_R1158_U517);
  and ginst12554 (P2_R1158_U14, P2_R1158_U340, P2_R1158_U343);
  and ginst12555 (P2_R1158_U140, P2_R1158_U209, P2_R1158_U318);
  and ginst12556 (P2_R1158_U141, P2_R1158_U13, P2_R1158_U60);
  and ginst12557 (P2_R1158_U142, P2_R1158_U392, P2_R1158_U393);
  and ginst12558 (P2_R1158_U143, P2_R1158_U214, P2_R1158_U564, P2_R1158_U565);
  and ginst12559 (P2_R1158_U144, P2_R1158_U326, P2_R1158_U8);
  and ginst12560 (P2_R1158_U145, P2_R1158_U43, P2_R1158_U590, P2_R1158_U591);
  and ginst12561 (P2_R1158_U146, P2_R1158_U333, P2_R1158_U7);
  and ginst12562 (P2_R1158_U147, P2_R1158_U213, P2_R1158_U611, P2_R1158_U612);
  and ginst12563 (P2_R1158_U148, P2_R1158_U342, P2_R1158_U6);
  nand ginst12564 (P2_R1158_U149, P2_R1158_U630, P2_R1158_U631);
  and ginst12565 (P2_R1158_U15, P2_R1158_U331, P2_R1158_U334);
  not ginst12566 (P2_R1158_U150, P2_U3416);
  and ginst12567 (P2_R1158_U151, P2_R1158_U398, P2_R1158_U399);
  not ginst12568 (P2_R1158_U152, P2_U3401);
  not ginst12569 (P2_R1158_U153, P2_U3392);
  not ginst12570 (P2_R1158_U154, P2_U3387);
  not ginst12571 (P2_R1158_U155, P2_U3398);
  not ginst12572 (P2_R1158_U156, P2_U3395);
  not ginst12573 (P2_R1158_U157, P2_U3404);
  not ginst12574 (P2_R1158_U158, P2_U3410);
  not ginst12575 (P2_R1158_U159, P2_U3407);
  and ginst12576 (P2_R1158_U16, P2_R1158_U324, P2_R1158_U327);
  not ginst12577 (P2_R1158_U160, P2_U3413);
  nand ginst12578 (P2_R1158_U161, P2_R1158_U122, P2_R1158_U390);
  and ginst12579 (P2_R1158_U162, P2_R1158_U432, P2_R1158_U433);
  nand ginst12580 (P2_R1158_U163, P2_R1158_U360, P2_R1158_U388);
  and ginst12581 (P2_R1158_U164, P2_R1158_U446, P2_R1158_U447);
  nand ginst12582 (P2_R1158_U165, P2_R1158_U211, P2_R1158_U233, P2_R1158_U354);
  and ginst12583 (P2_R1158_U166, P2_R1158_U453, P2_R1158_U454);
  nand ginst12584 (P2_R1158_U167, P2_R1158_U120, P2_R1158_U231);
  not ginst12585 (P2_R1158_U168, P2_U3896);
  not ginst12586 (P2_R1158_U169, P2_U3431);
  and ginst12587 (P2_R1158_U17, P2_R1158_U142, P2_R1158_U394, P2_R1158_U538, P2_R1158_U539);
  not ginst12588 (P2_R1158_U170, P2_U3419);
  not ginst12589 (P2_R1158_U171, P2_U3422);
  not ginst12590 (P2_R1158_U172, P2_U3428);
  not ginst12591 (P2_R1158_U173, P2_U3425);
  not ginst12592 (P2_R1158_U174, P2_U3434);
  not ginst12593 (P2_R1158_U175, P2_U3440);
  not ginst12594 (P2_R1158_U176, P2_U3437);
  not ginst12595 (P2_R1158_U177, P2_U3443);
  not ginst12596 (P2_R1158_U178, P2_U3902);
  not ginst12597 (P2_R1158_U179, P2_U3903);
  and ginst12598 (P2_R1158_U18, P2_R1158_U254, P2_R1158_U257);
  not ginst12599 (P2_R1158_U180, P2_U3445);
  not ginst12600 (P2_R1158_U181, P2_U3901);
  not ginst12601 (P2_R1158_U182, P2_U3900);
  not ginst12602 (P2_R1158_U183, P2_U3897);
  not ginst12603 (P2_R1158_U184, P2_U3898);
  not ginst12604 (P2_R1158_U185, P2_U3899);
  not ginst12605 (P2_R1158_U186, P2_U3053);
  not ginst12606 (P2_R1158_U187, P2_U3895);
  and ginst12607 (P2_R1158_U188, P2_R1158_U529, P2_R1158_U530);
  nand ginst12608 (P2_R1158_U189, P2_R1158_U309, P2_R1158_U310);
  and ginst12609 (P2_R1158_U19, P2_R1158_U247, P2_R1158_U250);
  nand ginst12610 (P2_R1158_U190, P2_R1158_U79, P2_U3064);
  nand ginst12611 (P2_R1158_U191, P2_R1158_U190, P2_R1158_U61);
  nand ginst12612 (P2_R1158_U192, P2_R1158_U302, P2_R1158_U303);
  and ginst12613 (P2_R1158_U193, P2_R1158_U550, P2_R1158_U551);
  nand ginst12614 (P2_R1158_U194, P2_R1158_U298, P2_R1158_U299);
  and ginst12615 (P2_R1158_U195, P2_R1158_U557, P2_R1158_U558);
  nand ginst12616 (P2_R1158_U196, P2_R1158_U294, P2_R1158_U295);
  and ginst12617 (P2_R1158_U197, P2_R1158_U571, P2_R1158_U572);
  nand ginst12618 (P2_R1158_U198, P2_R1158_U220, P2_R1158_U221);
  nand ginst12619 (P2_R1158_U199, P2_R1158_U284, P2_R1158_U285);
  nand ginst12620 (P2_R1158_U20, P2_R1158_U305, P2_U3056);
  and ginst12621 (P2_R1158_U200, P2_R1158_U583, P2_R1158_U584);
  nand ginst12622 (P2_R1158_U201, P2_R1158_U130, P2_R1158_U281);
  and ginst12623 (P2_R1158_U202, P2_R1158_U597, P2_R1158_U598);
  nand ginst12624 (P2_R1158_U203, P2_R1158_U368, P2_R1158_U382);
  and ginst12625 (P2_R1158_U204, P2_R1158_U604, P2_R1158_U605);
  nand ginst12626 (P2_R1158_U205, P2_R1158_U363, P2_R1158_U380);
  nand ginst12627 (P2_R1158_U206, P2_R1158_U378, P2_R1158_U52);
  and ginst12628 (P2_R1158_U207, P2_R1158_U623, P2_R1158_U624);
  nand ginst12629 (P2_R1158_U208, P2_R1158_U210, P2_R1158_U259, P2_R1158_U355);
  nand ginst12630 (P2_R1158_U209, P2_R1158_U20, P2_R1158_U366);
  not ginst12631 (P2_R1158_U21, P2_U3152);
  nand ginst12632 (P2_R1158_U210, P2_R1158_U161, P2_R1158_U67);
  nand ginst12633 (P2_R1158_U211, P2_R1158_U167, P2_R1158_U76);
  not ginst12634 (P2_R1158_U212, P2_R1158_U29);
  nand ginst12635 (P2_R1158_U213, P2_R1158_U85, P2_U3071);
  nand ginst12636 (P2_R1158_U214, P2_R1158_U92, P2_U3075);
  not ginst12637 (P2_R1158_U215, P2_R1158_U60);
  not ginst12638 (P2_R1158_U216, P2_R1158_U49);
  not ginst12639 (P2_R1158_U217, P2_R1158_U56);
  not ginst12640 (P2_R1158_U218, P2_R1158_U190);
  nand ginst12641 (P2_R1158_U219, P2_R1158_U21, P2_R1158_U411);
  not ginst12642 (P2_R1158_U22, P2_U3083);
  nand ginst12643 (P2_R1158_U220, P2_R1158_U219, P2_U3076);
  nand ginst12644 (P2_R1158_U221, P2_R1158_U75, P2_U3152);
  not ginst12645 (P2_R1158_U222, P2_R1158_U198);
  nand ginst12646 (P2_R1158_U223, P2_R1158_U31, P2_R1158_U408);
  nand ginst12647 (P2_R1158_U224, P2_R1158_U74, P2_U3077);
  not ginst12648 (P2_R1158_U225, P2_R1158_U37);
  nand ginst12649 (P2_R1158_U226, P2_R1158_U30, P2_R1158_U414);
  nand ginst12650 (P2_R1158_U227, P2_R1158_U28, P2_R1158_U417);
  nand ginst12651 (P2_R1158_U228, P2_R1158_U29, P2_R1158_U30);
  nand ginst12652 (P2_R1158_U229, P2_R1158_U228, P2_R1158_U73);
  not ginst12653 (P2_R1158_U23, P2_U3070);
  nand ginst12654 (P2_R1158_U230, P2_R1158_U212, P2_U3063);
  nand ginst12655 (P2_R1158_U231, P2_R1158_U37, P2_R1158_U4);
  not ginst12656 (P2_R1158_U232, P2_R1158_U167);
  nand ginst12657 (P2_R1158_U233, P2_R1158_U167, P2_U3059);
  not ginst12658 (P2_R1158_U234, P2_R1158_U165);
  nand ginst12659 (P2_R1158_U235, P2_R1158_U26, P2_R1158_U420);
  not ginst12660 (P2_R1158_U236, P2_R1158_U27);
  nand ginst12661 (P2_R1158_U237, P2_R1158_U25, P2_R1158_U423);
  nand ginst12662 (P2_R1158_U238, P2_R1158_U23, P2_R1158_U426);
  not ginst12663 (P2_R1158_U239, P2_R1158_U24);
  nand ginst12664 (P2_R1158_U24, P2_R1158_U69, P2_U3070);
  nand ginst12665 (P2_R1158_U240, P2_R1158_U24, P2_R1158_U25);
  nand ginst12666 (P2_R1158_U241, P2_R1158_U240, P2_R1158_U70);
  nand ginst12667 (P2_R1158_U242, P2_R1158_U239, P2_U3069);
  nand ginst12668 (P2_R1158_U243, P2_R1158_U22, P2_R1158_U429);
  nand ginst12669 (P2_R1158_U244, P2_R1158_U68, P2_U3083);
  nand ginst12670 (P2_R1158_U245, P2_R1158_U23, P2_R1158_U426);
  nand ginst12671 (P2_R1158_U246, P2_R1158_U245, P2_R1158_U36);
  nand ginst12672 (P2_R1158_U247, P2_R1158_U123, P2_R1158_U246);
  nand ginst12673 (P2_R1158_U248, P2_R1158_U24, P2_R1158_U387);
  nand ginst12674 (P2_R1158_U249, P2_R1158_U70, P2_U3069);
  not ginst12675 (P2_R1158_U25, P2_U3069);
  nand ginst12676 (P2_R1158_U250, P2_R1158_U124, P2_R1158_U248);
  nand ginst12677 (P2_R1158_U251, P2_R1158_U23, P2_R1158_U426);
  nand ginst12678 (P2_R1158_U252, P2_R1158_U28, P2_R1158_U417);
  nand ginst12679 (P2_R1158_U253, P2_R1158_U252, P2_R1158_U37);
  nand ginst12680 (P2_R1158_U254, P2_R1158_U125, P2_R1158_U253);
  nand ginst12681 (P2_R1158_U255, P2_R1158_U225, P2_R1158_U29);
  nand ginst12682 (P2_R1158_U256, P2_R1158_U73, P2_U3063);
  nand ginst12683 (P2_R1158_U257, P2_R1158_U126, P2_R1158_U255);
  nand ginst12684 (P2_R1158_U258, P2_R1158_U28, P2_R1158_U417);
  nand ginst12685 (P2_R1158_U259, P2_R1158_U161, P2_U3082);
  not ginst12686 (P2_R1158_U26, P2_U3066);
  not ginst12687 (P2_R1158_U260, P2_R1158_U208);
  nand ginst12688 (P2_R1158_U261, P2_R1158_U475, P2_R1158_U51);
  not ginst12689 (P2_R1158_U262, P2_R1158_U52);
  nand ginst12690 (P2_R1158_U263, P2_R1158_U481, P2_R1158_U50);
  nand ginst12691 (P2_R1158_U264, P2_R1158_U47, P2_R1158_U484);
  nand ginst12692 (P2_R1158_U265, P2_R1158_U216, P2_R1158_U6);
  nand ginst12693 (P2_R1158_U266, P2_R1158_U86, P2_U3079);
  nand ginst12694 (P2_R1158_U267, P2_R1158_U127, P2_R1158_U265);
  nand ginst12695 (P2_R1158_U268, P2_R1158_U478, P2_R1158_U48);
  nand ginst12696 (P2_R1158_U269, P2_R1158_U481, P2_R1158_U50);
  nand ginst12697 (P2_R1158_U27, P2_R1158_U71, P2_U3066);
  nand ginst12698 (P2_R1158_U270, P2_R1158_U267, P2_R1158_U269);
  nand ginst12699 (P2_R1158_U271, P2_R1158_U46, P2_R1158_U472);
  nand ginst12700 (P2_R1158_U272, P2_R1158_U84, P2_U3078);
  nand ginst12701 (P2_R1158_U273, P2_R1158_U45, P2_R1158_U487);
  nand ginst12702 (P2_R1158_U274, P2_R1158_U83, P2_U3073);
  nand ginst12703 (P2_R1158_U275, P2_R1158_U44, P2_R1158_U490);
  nand ginst12704 (P2_R1158_U276, P2_R1158_U42, P2_R1158_U493);
  not ginst12705 (P2_R1158_U277, P2_R1158_U43);
  nand ginst12706 (P2_R1158_U278, P2_R1158_U43, P2_R1158_U44);
  nand ginst12707 (P2_R1158_U279, P2_R1158_U278, P2_R1158_U82);
  not ginst12708 (P2_R1158_U28, P2_U3067);
  nand ginst12709 (P2_R1158_U280, P2_R1158_U277, P2_U3068);
  nand ginst12710 (P2_R1158_U281, P2_R1158_U63, P2_R1158_U7);
  not ginst12711 (P2_R1158_U282, P2_R1158_U201);
  nand ginst12712 (P2_R1158_U283, P2_R1158_U496, P2_R1158_U53);
  nand ginst12713 (P2_R1158_U284, P2_R1158_U201, P2_R1158_U283);
  nand ginst12714 (P2_R1158_U285, P2_R1158_U89, P2_U3081);
  not ginst12715 (P2_R1158_U286, P2_R1158_U199);
  nand ginst12716 (P2_R1158_U287, P2_R1158_U499, P2_R1158_U57);
  nand ginst12717 (P2_R1158_U288, P2_R1158_U502, P2_R1158_U54);
  nand ginst12718 (P2_R1158_U289, P2_R1158_U217, P2_R1158_U8);
  nand ginst12719 (P2_R1158_U29, P2_R1158_U72, P2_U3067);
  nand ginst12720 (P2_R1158_U290, P2_R1158_U91, P2_U3074);
  nand ginst12721 (P2_R1158_U291, P2_R1158_U132, P2_R1158_U289);
  nand ginst12722 (P2_R1158_U292, P2_R1158_U505, P2_R1158_U55);
  nand ginst12723 (P2_R1158_U293, P2_R1158_U499, P2_R1158_U57);
  nand ginst12724 (P2_R1158_U294, P2_R1158_U131, P2_R1158_U199);
  nand ginst12725 (P2_R1158_U295, P2_R1158_U291, P2_R1158_U293);
  not ginst12726 (P2_R1158_U296, P2_R1158_U196);
  nand ginst12727 (P2_R1158_U297, P2_R1158_U508, P2_R1158_U58);
  nand ginst12728 (P2_R1158_U298, P2_R1158_U196, P2_R1158_U297);
  nand ginst12729 (P2_R1158_U299, P2_R1158_U93, P2_U3060);
  not ginst12730 (P2_R1158_U30, P2_U3063);
  not ginst12731 (P2_R1158_U300, P2_R1158_U194);
  nand ginst12732 (P2_R1158_U301, P2_R1158_U511, P2_R1158_U59);
  nand ginst12733 (P2_R1158_U302, P2_R1158_U194, P2_R1158_U301);
  nand ginst12734 (P2_R1158_U303, P2_R1158_U94, P2_U3065);
  not ginst12735 (P2_R1158_U304, P2_R1158_U192);
  nand ginst12736 (P2_R1158_U305, P2_R1158_U39, P2_R1158_U517);
  nand ginst12737 (P2_R1158_U306, P2_R1158_U190, P2_R1158_U307, P2_R1158_U60);
  nand ginst12738 (P2_R1158_U307, P2_R1158_U80, P2_U3056);
  nand ginst12739 (P2_R1158_U308, P2_R1158_U40, P2_R1158_U520);
  nand ginst12740 (P2_R1158_U309, P2_R1158_U192, P2_R1158_U369);
  not ginst12741 (P2_R1158_U31, P2_U3077);
  nand ginst12742 (P2_R1158_U310, P2_R1158_U306, P2_R1158_U365);
  not ginst12743 (P2_R1158_U311, P2_R1158_U189);
  nand ginst12744 (P2_R1158_U312, P2_R1158_U38, P2_R1158_U469);
  nand ginst12745 (P2_R1158_U313, P2_R1158_U77, P2_U3052);
  nand ginst12746 (P2_R1158_U314, P2_R1158_U77, P2_U3052);
  nand ginst12747 (P2_R1158_U315, P2_R1158_U38, P2_R1158_U469);
  not ginst12748 (P2_R1158_U316, P2_R1158_U61);
  not ginst12749 (P2_R1158_U317, P2_R1158_U191);
  nand ginst12750 (P2_R1158_U318, P2_R1158_U80, P2_U3056);
  nand ginst12751 (P2_R1158_U319, P2_R1158_U39, P2_R1158_U517);
  not ginst12752 (P2_R1158_U32, P2_U3076);
  nand ginst12753 (P2_R1158_U320, P2_R1158_U199, P2_R1158_U292);
  not ginst12754 (P2_R1158_U321, P2_R1158_U62);
  nand ginst12755 (P2_R1158_U322, P2_R1158_U502, P2_R1158_U54);
  nand ginst12756 (P2_R1158_U323, P2_R1158_U322, P2_R1158_U62);
  nand ginst12757 (P2_R1158_U324, P2_R1158_U143, P2_R1158_U323);
  nand ginst12758 (P2_R1158_U325, P2_R1158_U214, P2_R1158_U321);
  nand ginst12759 (P2_R1158_U326, P2_R1158_U91, P2_U3074);
  nand ginst12760 (P2_R1158_U327, P2_R1158_U144, P2_R1158_U325);
  nand ginst12761 (P2_R1158_U328, P2_R1158_U502, P2_R1158_U54);
  nand ginst12762 (P2_R1158_U329, P2_R1158_U42, P2_R1158_U493);
  not ginst12763 (P2_R1158_U33, P2_U3059);
  nand ginst12764 (P2_R1158_U330, P2_R1158_U329, P2_R1158_U63);
  nand ginst12765 (P2_R1158_U331, P2_R1158_U145, P2_R1158_U330);
  nand ginst12766 (P2_R1158_U332, P2_R1158_U385, P2_R1158_U43);
  nand ginst12767 (P2_R1158_U333, P2_R1158_U82, P2_U3068);
  nand ginst12768 (P2_R1158_U334, P2_R1158_U146, P2_R1158_U332);
  nand ginst12769 (P2_R1158_U335, P2_R1158_U42, P2_R1158_U493);
  nand ginst12770 (P2_R1158_U336, P2_R1158_U206, P2_R1158_U268);
  not ginst12771 (P2_R1158_U337, P2_R1158_U66);
  nand ginst12772 (P2_R1158_U338, P2_R1158_U47, P2_R1158_U484);
  nand ginst12773 (P2_R1158_U339, P2_R1158_U338, P2_R1158_U66);
  not ginst12774 (P2_R1158_U34, P2_U3082);
  nand ginst12775 (P2_R1158_U340, P2_R1158_U147, P2_R1158_U339);
  nand ginst12776 (P2_R1158_U341, P2_R1158_U213, P2_R1158_U337);
  nand ginst12777 (P2_R1158_U342, P2_R1158_U86, P2_U3079);
  nand ginst12778 (P2_R1158_U343, P2_R1158_U148, P2_R1158_U341);
  nand ginst12779 (P2_R1158_U344, P2_R1158_U47, P2_R1158_U484);
  nand ginst12780 (P2_R1158_U345, P2_R1158_U24, P2_R1158_U251);
  nand ginst12781 (P2_R1158_U346, P2_R1158_U258, P2_R1158_U29);
  nand ginst12782 (P2_R1158_U347, P2_R1158_U319, P2_R1158_U60);
  nand ginst12783 (P2_R1158_U348, P2_R1158_U190, P2_R1158_U308);
  nand ginst12784 (P2_R1158_U349, P2_R1158_U214, P2_R1158_U328);
  nand ginst12785 (P2_R1158_U35, P2_R1158_U241, P2_R1158_U242, P2_R1158_U359);
  nand ginst12786 (P2_R1158_U350, P2_R1158_U292, P2_R1158_U56);
  nand ginst12787 (P2_R1158_U351, P2_R1158_U335, P2_R1158_U43);
  nand ginst12788 (P2_R1158_U352, P2_R1158_U213, P2_R1158_U344);
  nand ginst12789 (P2_R1158_U353, P2_R1158_U268, P2_R1158_U49);
  nand ginst12790 (P2_R1158_U354, P2_R1158_U76, P2_U3059);
  nand ginst12791 (P2_R1158_U355, P2_R1158_U67, P2_U3082);
  nand ginst12792 (P2_R1158_U356, P2_R1158_U133, P2_R1158_U309);
  nand ginst12793 (P2_R1158_U357, P2_R1158_U219, P2_R1158_U223, P2_U3076);
  nand ginst12794 (P2_R1158_U358, P2_R1158_U119, P2_R1158_U223);
  nand ginst12795 (P2_R1158_U359, P2_R1158_U236, P2_R1158_U5);
  nand ginst12796 (P2_R1158_U36, P2_R1158_U27, P2_R1158_U386);
  not ginst12797 (P2_R1158_U360, P2_R1158_U35);
  nand ginst12798 (P2_R1158_U361, P2_R1158_U243, P2_R1158_U35);
  nand ginst12799 (P2_R1158_U362, P2_R1158_U262, P2_R1158_U9);
  not ginst12800 (P2_R1158_U363, P2_R1158_U65);
  nand ginst12801 (P2_R1158_U364, P2_R1158_U271, P2_R1158_U65);
  nand ginst12802 (P2_R1158_U365, P2_R1158_U20, P2_R1158_U307, P2_R1158_U366);
  nand ginst12803 (P2_R1158_U366, P2_R1158_U305, P2_R1158_U80);
  not ginst12804 (P2_R1158_U367, P2_R1158_U20);
  not ginst12805 (P2_R1158_U368, P2_R1158_U64);
  nand ginst12806 (P2_R1158_U369, P2_R1158_U370, P2_R1158_U371);
  nand ginst12807 (P2_R1158_U37, P2_R1158_U224, P2_R1158_U357, P2_R1158_U358);
  nand ginst12808 (P2_R1158_U370, P2_R1158_U305, P2_R1158_U308, P2_R1158_U80);
  nand ginst12809 (P2_R1158_U371, P2_R1158_U308, P2_R1158_U367);
  nand ginst12810 (P2_R1158_U372, P2_R1158_U273, P2_R1158_U64);
  nand ginst12811 (P2_R1158_U373, P2_R1158_U134, P2_R1158_U365);
  nand ginst12812 (P2_R1158_U374, P2_R1158_U135, P2_R1158_U192);
  nand ginst12813 (P2_R1158_U375, P2_R1158_U376, P2_R1158_U377);
  nand ginst12814 (P2_R1158_U376, P2_R1158_U190, P2_R1158_U307, P2_R1158_U60);
  nand ginst12815 (P2_R1158_U377, P2_R1158_U20, P2_R1158_U307, P2_R1158_U366);
  nand ginst12816 (P2_R1158_U378, P2_R1158_U208, P2_R1158_U261);
  not ginst12817 (P2_R1158_U379, P2_R1158_U206);
  not ginst12818 (P2_R1158_U38, P2_U3052);
  nand ginst12819 (P2_R1158_U380, P2_R1158_U11, P2_R1158_U208);
  not ginst12820 (P2_R1158_U381, P2_R1158_U205);
  nand ginst12821 (P2_R1158_U382, P2_R1158_U12, P2_R1158_U208);
  not ginst12822 (P2_R1158_U383, P2_R1158_U203);
  nand ginst12823 (P2_R1158_U384, P2_R1158_U128, P2_R1158_U208);
  not ginst12824 (P2_R1158_U385, P2_R1158_U63);
  nand ginst12825 (P2_R1158_U386, P2_R1158_U165, P2_R1158_U235);
  not ginst12826 (P2_R1158_U387, P2_R1158_U36);
  nand ginst12827 (P2_R1158_U388, P2_R1158_U10, P2_R1158_U165);
  not ginst12828 (P2_R1158_U389, P2_R1158_U163);
  not ginst12829 (P2_R1158_U39, P2_U3057);
  nand ginst12830 (P2_R1158_U390, P2_R1158_U121, P2_R1158_U165);
  not ginst12831 (P2_R1158_U391, P2_R1158_U161);
  nand ginst12832 (P2_R1158_U392, P2_R1158_U138, P2_R1158_U209);
  nand ginst12833 (P2_R1158_U393, P2_R1158_U13, P2_R1158_U139);
  nand ginst12834 (P2_R1158_U394, P2_R1158_U140, P2_R1158_U316);
  nand ginst12835 (P2_R1158_U395, P2_R1158_U150, P2_U3152);
  nand ginst12836 (P2_R1158_U396, P2_R1158_U21, P2_U3416);
  not ginst12837 (P2_R1158_U397, P2_R1158_U67);
  nand ginst12838 (P2_R1158_U398, P2_R1158_U397, P2_U3082);
  nand ginst12839 (P2_R1158_U399, P2_R1158_U34, P2_R1158_U67);
  and ginst12840 (P2_R1158_U4, P2_R1158_U226, P2_R1158_U227);
  not ginst12841 (P2_R1158_U40, P2_U3064);
  nand ginst12842 (P2_R1158_U400, P2_R1158_U397, P2_U3082);
  nand ginst12843 (P2_R1158_U401, P2_R1158_U34, P2_R1158_U67);
  nand ginst12844 (P2_R1158_U402, P2_R1158_U400, P2_R1158_U401);
  nand ginst12845 (P2_R1158_U403, P2_R1158_U152, P2_U3152);
  nand ginst12846 (P2_R1158_U404, P2_R1158_U21, P2_U3401);
  not ginst12847 (P2_R1158_U405, P2_R1158_U76);
  nand ginst12848 (P2_R1158_U406, P2_R1158_U153, P2_U3152);
  nand ginst12849 (P2_R1158_U407, P2_R1158_U21, P2_U3392);
  not ginst12850 (P2_R1158_U408, P2_R1158_U74);
  nand ginst12851 (P2_R1158_U409, P2_R1158_U154, P2_U3152);
  not ginst12852 (P2_R1158_U41, P2_U3056);
  nand ginst12853 (P2_R1158_U410, P2_R1158_U21, P2_U3387);
  not ginst12854 (P2_R1158_U411, P2_R1158_U75);
  nand ginst12855 (P2_R1158_U412, P2_R1158_U155, P2_U3152);
  nand ginst12856 (P2_R1158_U413, P2_R1158_U21, P2_U3398);
  not ginst12857 (P2_R1158_U414, P2_R1158_U73);
  nand ginst12858 (P2_R1158_U415, P2_R1158_U156, P2_U3152);
  nand ginst12859 (P2_R1158_U416, P2_R1158_U21, P2_U3395);
  not ginst12860 (P2_R1158_U417, P2_R1158_U72);
  nand ginst12861 (P2_R1158_U418, P2_R1158_U157, P2_U3152);
  nand ginst12862 (P2_R1158_U419, P2_R1158_U21, P2_U3404);
  not ginst12863 (P2_R1158_U42, P2_U3072);
  not ginst12864 (P2_R1158_U420, P2_R1158_U71);
  nand ginst12865 (P2_R1158_U421, P2_R1158_U158, P2_U3152);
  nand ginst12866 (P2_R1158_U422, P2_R1158_U21, P2_U3410);
  not ginst12867 (P2_R1158_U423, P2_R1158_U70);
  nand ginst12868 (P2_R1158_U424, P2_R1158_U159, P2_U3152);
  nand ginst12869 (P2_R1158_U425, P2_R1158_U21, P2_U3407);
  not ginst12870 (P2_R1158_U426, P2_R1158_U69);
  nand ginst12871 (P2_R1158_U427, P2_R1158_U160, P2_U3152);
  nand ginst12872 (P2_R1158_U428, P2_R1158_U21, P2_U3413);
  not ginst12873 (P2_R1158_U429, P2_R1158_U68);
  nand ginst12874 (P2_R1158_U43, P2_R1158_U81, P2_U3072);
  nand ginst12875 (P2_R1158_U430, P2_R1158_U151, P2_R1158_U161);
  nand ginst12876 (P2_R1158_U431, P2_R1158_U391, P2_R1158_U402);
  nand ginst12877 (P2_R1158_U432, P2_R1158_U429, P2_U3083);
  nand ginst12878 (P2_R1158_U433, P2_R1158_U22, P2_R1158_U68);
  nand ginst12879 (P2_R1158_U434, P2_R1158_U429, P2_U3083);
  nand ginst12880 (P2_R1158_U435, P2_R1158_U22, P2_R1158_U68);
  nand ginst12881 (P2_R1158_U436, P2_R1158_U434, P2_R1158_U435);
  nand ginst12882 (P2_R1158_U437, P2_R1158_U162, P2_R1158_U163);
  nand ginst12883 (P2_R1158_U438, P2_R1158_U389, P2_R1158_U436);
  nand ginst12884 (P2_R1158_U439, P2_R1158_U423, P2_U3069);
  not ginst12885 (P2_R1158_U44, P2_U3068);
  nand ginst12886 (P2_R1158_U440, P2_R1158_U25, P2_R1158_U70);
  nand ginst12887 (P2_R1158_U441, P2_R1158_U426, P2_U3070);
  nand ginst12888 (P2_R1158_U442, P2_R1158_U23, P2_R1158_U69);
  nand ginst12889 (P2_R1158_U443, P2_R1158_U441, P2_R1158_U442);
  nand ginst12890 (P2_R1158_U444, P2_R1158_U345, P2_R1158_U36);
  nand ginst12891 (P2_R1158_U445, P2_R1158_U387, P2_R1158_U443);
  nand ginst12892 (P2_R1158_U446, P2_R1158_U420, P2_U3066);
  nand ginst12893 (P2_R1158_U447, P2_R1158_U26, P2_R1158_U71);
  nand ginst12894 (P2_R1158_U448, P2_R1158_U420, P2_U3066);
  nand ginst12895 (P2_R1158_U449, P2_R1158_U26, P2_R1158_U71);
  not ginst12896 (P2_R1158_U45, P2_U3073);
  nand ginst12897 (P2_R1158_U450, P2_R1158_U448, P2_R1158_U449);
  nand ginst12898 (P2_R1158_U451, P2_R1158_U164, P2_R1158_U165);
  nand ginst12899 (P2_R1158_U452, P2_R1158_U234, P2_R1158_U450);
  nand ginst12900 (P2_R1158_U453, P2_R1158_U405, P2_U3059);
  nand ginst12901 (P2_R1158_U454, P2_R1158_U33, P2_R1158_U76);
  nand ginst12902 (P2_R1158_U455, P2_R1158_U405, P2_U3059);
  nand ginst12903 (P2_R1158_U456, P2_R1158_U33, P2_R1158_U76);
  nand ginst12904 (P2_R1158_U457, P2_R1158_U455, P2_R1158_U456);
  nand ginst12905 (P2_R1158_U458, P2_R1158_U166, P2_R1158_U167);
  nand ginst12906 (P2_R1158_U459, P2_R1158_U232, P2_R1158_U457);
  not ginst12907 (P2_R1158_U46, P2_U3078);
  nand ginst12908 (P2_R1158_U460, P2_R1158_U414, P2_U3063);
  nand ginst12909 (P2_R1158_U461, P2_R1158_U30, P2_R1158_U73);
  nand ginst12910 (P2_R1158_U462, P2_R1158_U417, P2_U3067);
  nand ginst12911 (P2_R1158_U463, P2_R1158_U28, P2_R1158_U72);
  nand ginst12912 (P2_R1158_U464, P2_R1158_U462, P2_R1158_U463);
  nand ginst12913 (P2_R1158_U465, P2_R1158_U346, P2_R1158_U37);
  nand ginst12914 (P2_R1158_U466, P2_R1158_U225, P2_R1158_U464);
  nand ginst12915 (P2_R1158_U467, P2_R1158_U168, P2_U3152);
  nand ginst12916 (P2_R1158_U468, P2_R1158_U21, P2_U3896);
  not ginst12917 (P2_R1158_U469, P2_R1158_U77);
  not ginst12918 (P2_R1158_U47, P2_U3071);
  nand ginst12919 (P2_R1158_U470, P2_R1158_U169, P2_U3152);
  nand ginst12920 (P2_R1158_U471, P2_R1158_U21, P2_U3431);
  not ginst12921 (P2_R1158_U472, P2_R1158_U84);
  nand ginst12922 (P2_R1158_U473, P2_R1158_U170, P2_U3152);
  nand ginst12923 (P2_R1158_U474, P2_R1158_U21, P2_U3419);
  not ginst12924 (P2_R1158_U475, P2_R1158_U88);
  nand ginst12925 (P2_R1158_U476, P2_R1158_U171, P2_U3152);
  nand ginst12926 (P2_R1158_U477, P2_R1158_U21, P2_U3422);
  not ginst12927 (P2_R1158_U478, P2_R1158_U87);
  nand ginst12928 (P2_R1158_U479, P2_R1158_U172, P2_U3152);
  not ginst12929 (P2_R1158_U48, P2_U3062);
  nand ginst12930 (P2_R1158_U480, P2_R1158_U21, P2_U3428);
  not ginst12931 (P2_R1158_U481, P2_R1158_U86);
  nand ginst12932 (P2_R1158_U482, P2_R1158_U173, P2_U3152);
  nand ginst12933 (P2_R1158_U483, P2_R1158_U21, P2_U3425);
  not ginst12934 (P2_R1158_U484, P2_R1158_U85);
  nand ginst12935 (P2_R1158_U485, P2_R1158_U174, P2_U3152);
  nand ginst12936 (P2_R1158_U486, P2_R1158_U21, P2_U3434);
  not ginst12937 (P2_R1158_U487, P2_R1158_U83);
  nand ginst12938 (P2_R1158_U488, P2_R1158_U175, P2_U3152);
  nand ginst12939 (P2_R1158_U489, P2_R1158_U21, P2_U3440);
  nand ginst12940 (P2_R1158_U49, P2_R1158_U87, P2_U3062);
  not ginst12941 (P2_R1158_U490, P2_R1158_U82);
  nand ginst12942 (P2_R1158_U491, P2_R1158_U176, P2_U3152);
  nand ginst12943 (P2_R1158_U492, P2_R1158_U21, P2_U3437);
  not ginst12944 (P2_R1158_U493, P2_R1158_U81);
  nand ginst12945 (P2_R1158_U494, P2_R1158_U177, P2_U3152);
  nand ginst12946 (P2_R1158_U495, P2_R1158_U21, P2_U3443);
  not ginst12947 (P2_R1158_U496, P2_R1158_U89);
  nand ginst12948 (P2_R1158_U497, P2_R1158_U178, P2_U3152);
  nand ginst12949 (P2_R1158_U498, P2_R1158_U21, P2_U3902);
  not ginst12950 (P2_R1158_U499, P2_R1158_U91);
  and ginst12951 (P2_R1158_U5, P2_R1158_U237, P2_R1158_U238);
  not ginst12952 (P2_R1158_U50, P2_U3079);
  nand ginst12953 (P2_R1158_U500, P2_R1158_U179, P2_U3152);
  nand ginst12954 (P2_R1158_U501, P2_R1158_U21, P2_U3903);
  not ginst12955 (P2_R1158_U502, P2_R1158_U92);
  nand ginst12956 (P2_R1158_U503, P2_R1158_U180, P2_U3152);
  nand ginst12957 (P2_R1158_U504, P2_R1158_U21, P2_U3445);
  not ginst12958 (P2_R1158_U505, P2_R1158_U90);
  nand ginst12959 (P2_R1158_U506, P2_R1158_U181, P2_U3152);
  nand ginst12960 (P2_R1158_U507, P2_R1158_U21, P2_U3901);
  not ginst12961 (P2_R1158_U508, P2_R1158_U93);
  nand ginst12962 (P2_R1158_U509, P2_R1158_U182, P2_U3152);
  not ginst12963 (P2_R1158_U51, P2_U3061);
  nand ginst12964 (P2_R1158_U510, P2_R1158_U21, P2_U3900);
  not ginst12965 (P2_R1158_U511, P2_R1158_U94);
  nand ginst12966 (P2_R1158_U512, P2_R1158_U183, P2_U3152);
  nand ginst12967 (P2_R1158_U513, P2_R1158_U21, P2_U3897);
  not ginst12968 (P2_R1158_U514, P2_R1158_U80);
  nand ginst12969 (P2_R1158_U515, P2_R1158_U184, P2_U3152);
  nand ginst12970 (P2_R1158_U516, P2_R1158_U21, P2_U3898);
  not ginst12971 (P2_R1158_U517, P2_R1158_U78);
  nand ginst12972 (P2_R1158_U518, P2_R1158_U185, P2_U3152);
  nand ginst12973 (P2_R1158_U519, P2_R1158_U21, P2_U3899);
  nand ginst12974 (P2_R1158_U52, P2_R1158_U88, P2_U3061);
  not ginst12975 (P2_R1158_U520, P2_R1158_U79);
  nand ginst12976 (P2_R1158_U521, P2_R1158_U186, P2_U3152);
  nand ginst12977 (P2_R1158_U522, P2_R1158_U21, P2_U3053);
  not ginst12978 (P2_R1158_U523, P2_R1158_U137);
  nand ginst12979 (P2_R1158_U524, P2_R1158_U523, P2_U3895);
  nand ginst12980 (P2_R1158_U525, P2_R1158_U137, P2_R1158_U187);
  not ginst12981 (P2_R1158_U526, P2_R1158_U95);
  nand ginst12982 (P2_R1158_U527, P2_R1158_U312, P2_R1158_U356, P2_R1158_U526);
  nand ginst12983 (P2_R1158_U528, P2_R1158_U136, P2_R1158_U374, P2_R1158_U95);
  nand ginst12984 (P2_R1158_U529, P2_R1158_U469, P2_U3052);
  not ginst12985 (P2_R1158_U53, P2_U3081);
  nand ginst12986 (P2_R1158_U530, P2_R1158_U38, P2_R1158_U77);
  nand ginst12987 (P2_R1158_U531, P2_R1158_U469, P2_U3052);
  nand ginst12988 (P2_R1158_U532, P2_R1158_U38, P2_R1158_U77);
  nand ginst12989 (P2_R1158_U533, P2_R1158_U531, P2_R1158_U532);
  nand ginst12990 (P2_R1158_U534, P2_R1158_U188, P2_R1158_U189);
  nand ginst12991 (P2_R1158_U535, P2_R1158_U311, P2_R1158_U533);
  nand ginst12992 (P2_R1158_U536, P2_R1158_U514, P2_U3056);
  nand ginst12993 (P2_R1158_U537, P2_R1158_U41, P2_R1158_U80);
  nand ginst12994 (P2_R1158_U538, P2_R1158_U141, P2_R1158_U190, P2_R1158_U61);
  nand ginst12995 (P2_R1158_U539, P2_R1158_U209, P2_R1158_U218, P2_R1158_U318);
  not ginst12996 (P2_R1158_U54, P2_U3075);
  nand ginst12997 (P2_R1158_U540, P2_R1158_U517, P2_U3057);
  nand ginst12998 (P2_R1158_U541, P2_R1158_U39, P2_R1158_U78);
  nand ginst12999 (P2_R1158_U542, P2_R1158_U540, P2_R1158_U541);
  nand ginst13000 (P2_R1158_U543, P2_R1158_U191, P2_R1158_U347);
  nand ginst13001 (P2_R1158_U544, P2_R1158_U317, P2_R1158_U542);
  nand ginst13002 (P2_R1158_U545, P2_R1158_U520, P2_U3064);
  nand ginst13003 (P2_R1158_U546, P2_R1158_U40, P2_R1158_U79);
  nand ginst13004 (P2_R1158_U547, P2_R1158_U545, P2_R1158_U546);
  nand ginst13005 (P2_R1158_U548, P2_R1158_U192, P2_R1158_U348);
  nand ginst13006 (P2_R1158_U549, P2_R1158_U304, P2_R1158_U547);
  not ginst13007 (P2_R1158_U55, P2_U3080);
  nand ginst13008 (P2_R1158_U550, P2_R1158_U511, P2_U3065);
  nand ginst13009 (P2_R1158_U551, P2_R1158_U59, P2_R1158_U94);
  nand ginst13010 (P2_R1158_U552, P2_R1158_U511, P2_U3065);
  nand ginst13011 (P2_R1158_U553, P2_R1158_U59, P2_R1158_U94);
  nand ginst13012 (P2_R1158_U554, P2_R1158_U552, P2_R1158_U553);
  nand ginst13013 (P2_R1158_U555, P2_R1158_U193, P2_R1158_U194);
  nand ginst13014 (P2_R1158_U556, P2_R1158_U300, P2_R1158_U554);
  nand ginst13015 (P2_R1158_U557, P2_R1158_U508, P2_U3060);
  nand ginst13016 (P2_R1158_U558, P2_R1158_U58, P2_R1158_U93);
  nand ginst13017 (P2_R1158_U559, P2_R1158_U508, P2_U3060);
  nand ginst13018 (P2_R1158_U56, P2_R1158_U90, P2_U3080);
  nand ginst13019 (P2_R1158_U560, P2_R1158_U58, P2_R1158_U93);
  nand ginst13020 (P2_R1158_U561, P2_R1158_U559, P2_R1158_U560);
  nand ginst13021 (P2_R1158_U562, P2_R1158_U195, P2_R1158_U196);
  nand ginst13022 (P2_R1158_U563, P2_R1158_U296, P2_R1158_U561);
  nand ginst13023 (P2_R1158_U564, P2_R1158_U499, P2_U3074);
  nand ginst13024 (P2_R1158_U565, P2_R1158_U57, P2_R1158_U91);
  nand ginst13025 (P2_R1158_U566, P2_R1158_U502, P2_U3075);
  nand ginst13026 (P2_R1158_U567, P2_R1158_U54, P2_R1158_U92);
  nand ginst13027 (P2_R1158_U568, P2_R1158_U566, P2_R1158_U567);
  nand ginst13028 (P2_R1158_U569, P2_R1158_U349, P2_R1158_U62);
  not ginst13029 (P2_R1158_U57, P2_U3074);
  nand ginst13030 (P2_R1158_U570, P2_R1158_U321, P2_R1158_U568);
  nand ginst13031 (P2_R1158_U571, P2_R1158_U408, P2_U3077);
  nand ginst13032 (P2_R1158_U572, P2_R1158_U31, P2_R1158_U74);
  nand ginst13033 (P2_R1158_U573, P2_R1158_U408, P2_U3077);
  nand ginst13034 (P2_R1158_U574, P2_R1158_U31, P2_R1158_U74);
  nand ginst13035 (P2_R1158_U575, P2_R1158_U573, P2_R1158_U574);
  nand ginst13036 (P2_R1158_U576, P2_R1158_U197, P2_R1158_U198);
  nand ginst13037 (P2_R1158_U577, P2_R1158_U222, P2_R1158_U575);
  nand ginst13038 (P2_R1158_U578, P2_R1158_U505, P2_U3080);
  nand ginst13039 (P2_R1158_U579, P2_R1158_U55, P2_R1158_U90);
  not ginst13040 (P2_R1158_U58, P2_U3060);
  nand ginst13041 (P2_R1158_U580, P2_R1158_U578, P2_R1158_U579);
  nand ginst13042 (P2_R1158_U581, P2_R1158_U199, P2_R1158_U350);
  nand ginst13043 (P2_R1158_U582, P2_R1158_U286, P2_R1158_U580);
  nand ginst13044 (P2_R1158_U583, P2_R1158_U496, P2_U3081);
  nand ginst13045 (P2_R1158_U584, P2_R1158_U53, P2_R1158_U89);
  nand ginst13046 (P2_R1158_U585, P2_R1158_U496, P2_U3081);
  nand ginst13047 (P2_R1158_U586, P2_R1158_U53, P2_R1158_U89);
  nand ginst13048 (P2_R1158_U587, P2_R1158_U585, P2_R1158_U586);
  nand ginst13049 (P2_R1158_U588, P2_R1158_U200, P2_R1158_U201);
  nand ginst13050 (P2_R1158_U589, P2_R1158_U282, P2_R1158_U587);
  not ginst13051 (P2_R1158_U59, P2_U3065);
  nand ginst13052 (P2_R1158_U590, P2_R1158_U490, P2_U3068);
  nand ginst13053 (P2_R1158_U591, P2_R1158_U44, P2_R1158_U82);
  nand ginst13054 (P2_R1158_U592, P2_R1158_U493, P2_U3072);
  nand ginst13055 (P2_R1158_U593, P2_R1158_U42, P2_R1158_U81);
  nand ginst13056 (P2_R1158_U594, P2_R1158_U592, P2_R1158_U593);
  nand ginst13057 (P2_R1158_U595, P2_R1158_U351, P2_R1158_U63);
  nand ginst13058 (P2_R1158_U596, P2_R1158_U385, P2_R1158_U594);
  nand ginst13059 (P2_R1158_U597, P2_R1158_U487, P2_U3073);
  nand ginst13060 (P2_R1158_U598, P2_R1158_U45, P2_R1158_U83);
  nand ginst13061 (P2_R1158_U599, P2_R1158_U487, P2_U3073);
  and ginst13062 (P2_R1158_U6, P2_R1158_U263, P2_R1158_U264);
  nand ginst13063 (P2_R1158_U60, P2_R1158_U78, P2_U3057);
  nand ginst13064 (P2_R1158_U600, P2_R1158_U45, P2_R1158_U83);
  nand ginst13065 (P2_R1158_U601, P2_R1158_U599, P2_R1158_U600);
  nand ginst13066 (P2_R1158_U602, P2_R1158_U202, P2_R1158_U203);
  nand ginst13067 (P2_R1158_U603, P2_R1158_U383, P2_R1158_U601);
  nand ginst13068 (P2_R1158_U604, P2_R1158_U472, P2_U3078);
  nand ginst13069 (P2_R1158_U605, P2_R1158_U46, P2_R1158_U84);
  nand ginst13070 (P2_R1158_U606, P2_R1158_U472, P2_U3078);
  nand ginst13071 (P2_R1158_U607, P2_R1158_U46, P2_R1158_U84);
  nand ginst13072 (P2_R1158_U608, P2_R1158_U606, P2_R1158_U607);
  nand ginst13073 (P2_R1158_U609, P2_R1158_U204, P2_R1158_U205);
  nand ginst13074 (P2_R1158_U61, P2_R1158_U192, P2_R1158_U308);
  nand ginst13075 (P2_R1158_U610, P2_R1158_U381, P2_R1158_U608);
  nand ginst13076 (P2_R1158_U611, P2_R1158_U481, P2_U3079);
  nand ginst13077 (P2_R1158_U612, P2_R1158_U50, P2_R1158_U86);
  nand ginst13078 (P2_R1158_U613, P2_R1158_U484, P2_U3071);
  nand ginst13079 (P2_R1158_U614, P2_R1158_U47, P2_R1158_U85);
  nand ginst13080 (P2_R1158_U615, P2_R1158_U613, P2_R1158_U614);
  nand ginst13081 (P2_R1158_U616, P2_R1158_U352, P2_R1158_U66);
  nand ginst13082 (P2_R1158_U617, P2_R1158_U337, P2_R1158_U615);
  nand ginst13083 (P2_R1158_U618, P2_R1158_U478, P2_U3062);
  nand ginst13084 (P2_R1158_U619, P2_R1158_U48, P2_R1158_U87);
  nand ginst13085 (P2_R1158_U62, P2_R1158_U320, P2_R1158_U56);
  nand ginst13086 (P2_R1158_U620, P2_R1158_U618, P2_R1158_U619);
  nand ginst13087 (P2_R1158_U621, P2_R1158_U206, P2_R1158_U353);
  nand ginst13088 (P2_R1158_U622, P2_R1158_U379, P2_R1158_U620);
  nand ginst13089 (P2_R1158_U623, P2_R1158_U475, P2_U3061);
  nand ginst13090 (P2_R1158_U624, P2_R1158_U51, P2_R1158_U88);
  nand ginst13091 (P2_R1158_U625, P2_R1158_U475, P2_U3061);
  nand ginst13092 (P2_R1158_U626, P2_R1158_U51, P2_R1158_U88);
  nand ginst13093 (P2_R1158_U627, P2_R1158_U625, P2_R1158_U626);
  nand ginst13094 (P2_R1158_U628, P2_R1158_U207, P2_R1158_U208);
  nand ginst13095 (P2_R1158_U629, P2_R1158_U260, P2_R1158_U627);
  nand ginst13096 (P2_R1158_U63, P2_R1158_U129, P2_R1158_U384);
  nand ginst13097 (P2_R1158_U630, P2_R1158_U21, P2_R1158_U75);
  nand ginst13098 (P2_R1158_U631, P2_R1158_U411, P2_U3152);
  not ginst13099 (P2_R1158_U632, P2_R1158_U149);
  nand ginst13100 (P2_R1158_U633, P2_R1158_U632, P2_U3076);
  nand ginst13101 (P2_R1158_U634, P2_R1158_U149, P2_R1158_U32);
  nand ginst13102 (P2_R1158_U64, P2_R1158_U272, P2_R1158_U364);
  nand ginst13103 (P2_R1158_U65, P2_R1158_U270, P2_R1158_U362);
  nand ginst13104 (P2_R1158_U66, P2_R1158_U336, P2_R1158_U49);
  nand ginst13105 (P2_R1158_U67, P2_R1158_U395, P2_R1158_U396);
  nand ginst13106 (P2_R1158_U68, P2_R1158_U427, P2_R1158_U428);
  nand ginst13107 (P2_R1158_U69, P2_R1158_U424, P2_R1158_U425);
  and ginst13108 (P2_R1158_U7, P2_R1158_U275, P2_R1158_U276);
  nand ginst13109 (P2_R1158_U70, P2_R1158_U421, P2_R1158_U422);
  nand ginst13110 (P2_R1158_U71, P2_R1158_U418, P2_R1158_U419);
  nand ginst13111 (P2_R1158_U72, P2_R1158_U415, P2_R1158_U416);
  nand ginst13112 (P2_R1158_U73, P2_R1158_U412, P2_R1158_U413);
  nand ginst13113 (P2_R1158_U74, P2_R1158_U406, P2_R1158_U407);
  nand ginst13114 (P2_R1158_U75, P2_R1158_U409, P2_R1158_U410);
  nand ginst13115 (P2_R1158_U76, P2_R1158_U403, P2_R1158_U404);
  nand ginst13116 (P2_R1158_U77, P2_R1158_U467, P2_R1158_U468);
  nand ginst13117 (P2_R1158_U78, P2_R1158_U515, P2_R1158_U516);
  nand ginst13118 (P2_R1158_U79, P2_R1158_U518, P2_R1158_U519);
  and ginst13119 (P2_R1158_U8, P2_R1158_U287, P2_R1158_U288);
  nand ginst13120 (P2_R1158_U80, P2_R1158_U512, P2_R1158_U513);
  nand ginst13121 (P2_R1158_U81, P2_R1158_U491, P2_R1158_U492);
  nand ginst13122 (P2_R1158_U82, P2_R1158_U488, P2_R1158_U489);
  nand ginst13123 (P2_R1158_U83, P2_R1158_U485, P2_R1158_U486);
  nand ginst13124 (P2_R1158_U84, P2_R1158_U470, P2_R1158_U471);
  nand ginst13125 (P2_R1158_U85, P2_R1158_U482, P2_R1158_U483);
  nand ginst13126 (P2_R1158_U86, P2_R1158_U479, P2_R1158_U480);
  nand ginst13127 (P2_R1158_U87, P2_R1158_U476, P2_R1158_U477);
  nand ginst13128 (P2_R1158_U88, P2_R1158_U473, P2_R1158_U474);
  nand ginst13129 (P2_R1158_U89, P2_R1158_U494, P2_R1158_U495);
  and ginst13130 (P2_R1158_U9, P2_R1158_U268, P2_R1158_U6);
  nand ginst13131 (P2_R1158_U90, P2_R1158_U503, P2_R1158_U504);
  nand ginst13132 (P2_R1158_U91, P2_R1158_U497, P2_R1158_U498);
  nand ginst13133 (P2_R1158_U92, P2_R1158_U500, P2_R1158_U501);
  nand ginst13134 (P2_R1158_U93, P2_R1158_U506, P2_R1158_U507);
  nand ginst13135 (P2_R1158_U94, P2_R1158_U509, P2_R1158_U510);
  nand ginst13136 (P2_R1158_U95, P2_R1158_U524, P2_R1158_U525);
  nand ginst13137 (P2_R1158_U96, P2_R1158_U633, P2_R1158_U634);
  nand ginst13138 (P2_R1158_U97, P2_R1158_U430, P2_R1158_U431);
  nand ginst13139 (P2_R1158_U98, P2_R1158_U437, P2_R1158_U438);
  nand ginst13140 (P2_R1158_U99, P2_R1158_U444, P2_R1158_U445);
  and ginst13141 (P2_R1161_U10, P2_R1161_U348, P2_R1161_U351);
  nand ginst13142 (P2_R1161_U100, P2_R1161_U398, P2_R1161_U399);
  nand ginst13143 (P2_R1161_U101, P2_R1161_U407, P2_R1161_U408);
  nand ginst13144 (P2_R1161_U102, P2_R1161_U414, P2_R1161_U415);
  nand ginst13145 (P2_R1161_U103, P2_R1161_U421, P2_R1161_U422);
  nand ginst13146 (P2_R1161_U104, P2_R1161_U428, P2_R1161_U429);
  nand ginst13147 (P2_R1161_U105, P2_R1161_U433, P2_R1161_U434);
  nand ginst13148 (P2_R1161_U106, P2_R1161_U440, P2_R1161_U441);
  nand ginst13149 (P2_R1161_U107, P2_R1161_U447, P2_R1161_U448);
  nand ginst13150 (P2_R1161_U108, P2_R1161_U461, P2_R1161_U462);
  nand ginst13151 (P2_R1161_U109, P2_R1161_U466, P2_R1161_U467);
  and ginst13152 (P2_R1161_U11, P2_R1161_U341, P2_R1161_U344);
  nand ginst13153 (P2_R1161_U110, P2_R1161_U473, P2_R1161_U474);
  nand ginst13154 (P2_R1161_U111, P2_R1161_U480, P2_R1161_U481);
  nand ginst13155 (P2_R1161_U112, P2_R1161_U487, P2_R1161_U488);
  nand ginst13156 (P2_R1161_U113, P2_R1161_U494, P2_R1161_U495);
  nand ginst13157 (P2_R1161_U114, P2_R1161_U499, P2_R1161_U500);
  and ginst13158 (P2_R1161_U115, P2_R1161_U187, P2_R1161_U189);
  and ginst13159 (P2_R1161_U116, P2_R1161_U180, P2_R1161_U4);
  and ginst13160 (P2_R1161_U117, P2_R1161_U192, P2_R1161_U194);
  and ginst13161 (P2_R1161_U118, P2_R1161_U200, P2_R1161_U201);
  and ginst13162 (P2_R1161_U119, P2_R1161_U22, P2_R1161_U381, P2_R1161_U382);
  and ginst13163 (P2_R1161_U12, P2_R1161_U332, P2_R1161_U335);
  and ginst13164 (P2_R1161_U120, P2_R1161_U212, P2_R1161_U5);
  and ginst13165 (P2_R1161_U121, P2_R1161_U180, P2_R1161_U181);
  and ginst13166 (P2_R1161_U122, P2_R1161_U218, P2_R1161_U220);
  and ginst13167 (P2_R1161_U123, P2_R1161_U34, P2_R1161_U388, P2_R1161_U389);
  and ginst13168 (P2_R1161_U124, P2_R1161_U226, P2_R1161_U4);
  and ginst13169 (P2_R1161_U125, P2_R1161_U181, P2_R1161_U234);
  and ginst13170 (P2_R1161_U126, P2_R1161_U204, P2_R1161_U6);
  and ginst13171 (P2_R1161_U127, P2_R1161_U239, P2_R1161_U243);
  and ginst13172 (P2_R1161_U128, P2_R1161_U250, P2_R1161_U7);
  and ginst13173 (P2_R1161_U129, P2_R1161_U248, P2_R1161_U253);
  and ginst13174 (P2_R1161_U13, P2_R1161_U323, P2_R1161_U326);
  and ginst13175 (P2_R1161_U130, P2_R1161_U267, P2_R1161_U268);
  and ginst13176 (P2_R1161_U131, P2_R1161_U282, P2_R1161_U9);
  and ginst13177 (P2_R1161_U132, P2_R1161_U280, P2_R1161_U285);
  and ginst13178 (P2_R1161_U133, P2_R1161_U298, P2_R1161_U301);
  and ginst13179 (P2_R1161_U134, P2_R1161_U302, P2_R1161_U368);
  and ginst13180 (P2_R1161_U135, P2_R1161_U160, P2_R1161_U278);
  and ginst13181 (P2_R1161_U136, P2_R1161_U454, P2_R1161_U455, P2_R1161_U80);
  and ginst13182 (P2_R1161_U137, P2_R1161_U325, P2_R1161_U9);
  and ginst13183 (P2_R1161_U138, P2_R1161_U468, P2_R1161_U469, P2_R1161_U59);
  and ginst13184 (P2_R1161_U139, P2_R1161_U334, P2_R1161_U8);
  and ginst13185 (P2_R1161_U14, P2_R1161_U318, P2_R1161_U320);
  and ginst13186 (P2_R1161_U140, P2_R1161_U172, P2_R1161_U489, P2_R1161_U490);
  and ginst13187 (P2_R1161_U141, P2_R1161_U343, P2_R1161_U7);
  and ginst13188 (P2_R1161_U142, P2_R1161_U171, P2_R1161_U501, P2_R1161_U502);
  and ginst13189 (P2_R1161_U143, P2_R1161_U350, P2_R1161_U6);
  nand ginst13190 (P2_R1161_U144, P2_R1161_U118, P2_R1161_U202);
  nand ginst13191 (P2_R1161_U145, P2_R1161_U217, P2_R1161_U229);
  not ginst13192 (P2_R1161_U146, P2_U3054);
  not ginst13193 (P2_R1161_U147, P2_U3904);
  and ginst13194 (P2_R1161_U148, P2_R1161_U402, P2_R1161_U403);
  nand ginst13195 (P2_R1161_U149, P2_R1161_U169, P2_R1161_U304, P2_R1161_U364);
  and ginst13196 (P2_R1161_U15, P2_R1161_U310, P2_R1161_U313);
  and ginst13197 (P2_R1161_U150, P2_R1161_U409, P2_R1161_U410);
  nand ginst13198 (P2_R1161_U151, P2_R1161_U134, P2_R1161_U369, P2_R1161_U370);
  and ginst13199 (P2_R1161_U152, P2_R1161_U416, P2_R1161_U417);
  nand ginst13200 (P2_R1161_U153, P2_R1161_U299, P2_R1161_U365, P2_R1161_U86);
  and ginst13201 (P2_R1161_U154, P2_R1161_U423, P2_R1161_U424);
  nand ginst13202 (P2_R1161_U155, P2_R1161_U292, P2_R1161_U293);
  and ginst13203 (P2_R1161_U156, P2_R1161_U435, P2_R1161_U436);
  nand ginst13204 (P2_R1161_U157, P2_R1161_U288, P2_R1161_U289);
  and ginst13205 (P2_R1161_U158, P2_R1161_U442, P2_R1161_U443);
  nand ginst13206 (P2_R1161_U159, P2_R1161_U132, P2_R1161_U284);
  and ginst13207 (P2_R1161_U16, P2_R1161_U232, P2_R1161_U235);
  and ginst13208 (P2_R1161_U160, P2_R1161_U449, P2_R1161_U450);
  nand ginst13209 (P2_R1161_U161, P2_R1161_U327, P2_R1161_U43);
  nand ginst13210 (P2_R1161_U162, P2_R1161_U130, P2_R1161_U269);
  and ginst13211 (P2_R1161_U163, P2_R1161_U475, P2_R1161_U476);
  nand ginst13212 (P2_R1161_U164, P2_R1161_U256, P2_R1161_U257);
  and ginst13213 (P2_R1161_U165, P2_R1161_U482, P2_R1161_U483);
  nand ginst13214 (P2_R1161_U166, P2_R1161_U129, P2_R1161_U252);
  nand ginst13215 (P2_R1161_U167, P2_R1161_U127, P2_R1161_U242);
  nand ginst13216 (P2_R1161_U168, P2_R1161_U366, P2_R1161_U367);
  nand ginst13217 (P2_R1161_U169, P2_R1161_U151, P2_U3053);
  and ginst13218 (P2_R1161_U17, P2_R1161_U224, P2_R1161_U227);
  not ginst13219 (P2_R1161_U170, P2_R1161_U34);
  nand ginst13220 (P2_R1161_U171, P2_U3082, P2_U3416);
  nand ginst13221 (P2_R1161_U172, P2_U3071, P2_U3425);
  nand ginst13222 (P2_R1161_U173, P2_U3057, P2_U3898);
  not ginst13223 (P2_R1161_U174, P2_R1161_U68);
  not ginst13224 (P2_R1161_U175, P2_R1161_U77);
  nand ginst13225 (P2_R1161_U176, P2_U3064, P2_U3899);
  not ginst13226 (P2_R1161_U177, P2_R1161_U65);
  or ginst13227 (P2_R1161_U178, P2_U3066, P2_U3404);
  or ginst13228 (P2_R1161_U179, P2_U3059, P2_U3401);
  and ginst13229 (P2_R1161_U18, P2_R1161_U210, P2_R1161_U213);
  or ginst13230 (P2_R1161_U180, P2_U3063, P2_U3398);
  or ginst13231 (P2_R1161_U181, P2_U3067, P2_U3395);
  not ginst13232 (P2_R1161_U182, P2_R1161_U31);
  or ginst13233 (P2_R1161_U183, P2_U3077, P2_U3392);
  not ginst13234 (P2_R1161_U184, P2_R1161_U42);
  not ginst13235 (P2_R1161_U185, P2_R1161_U43);
  nand ginst13236 (P2_R1161_U186, P2_R1161_U42, P2_R1161_U43);
  nand ginst13237 (P2_R1161_U187, P2_U3067, P2_U3395);
  nand ginst13238 (P2_R1161_U188, P2_R1161_U181, P2_R1161_U186);
  nand ginst13239 (P2_R1161_U189, P2_U3063, P2_U3398);
  not ginst13240 (P2_R1161_U19, P2_U3407);
  nand ginst13241 (P2_R1161_U190, P2_R1161_U115, P2_R1161_U188);
  nand ginst13242 (P2_R1161_U191, P2_R1161_U34, P2_R1161_U35);
  nand ginst13243 (P2_R1161_U192, P2_R1161_U191, P2_U3066);
  nand ginst13244 (P2_R1161_U193, P2_R1161_U116, P2_R1161_U190);
  nand ginst13245 (P2_R1161_U194, P2_R1161_U170, P2_U3404);
  not ginst13246 (P2_R1161_U195, P2_R1161_U41);
  or ginst13247 (P2_R1161_U196, P2_U3069, P2_U3410);
  or ginst13248 (P2_R1161_U197, P2_U3070, P2_U3407);
  not ginst13249 (P2_R1161_U198, P2_R1161_U22);
  nand ginst13250 (P2_R1161_U199, P2_R1161_U22, P2_R1161_U23);
  not ginst13251 (P2_R1161_U20, P2_U3070);
  nand ginst13252 (P2_R1161_U200, P2_R1161_U199, P2_U3069);
  nand ginst13253 (P2_R1161_U201, P2_R1161_U198, P2_U3410);
  nand ginst13254 (P2_R1161_U202, P2_R1161_U41, P2_R1161_U5);
  not ginst13255 (P2_R1161_U203, P2_R1161_U144);
  or ginst13256 (P2_R1161_U204, P2_U3083, P2_U3413);
  nand ginst13257 (P2_R1161_U205, P2_R1161_U144, P2_R1161_U204);
  not ginst13258 (P2_R1161_U206, P2_R1161_U40);
  or ginst13259 (P2_R1161_U207, P2_U3082, P2_U3416);
  or ginst13260 (P2_R1161_U208, P2_U3070, P2_U3407);
  nand ginst13261 (P2_R1161_U209, P2_R1161_U208, P2_R1161_U41);
  not ginst13262 (P2_R1161_U21, P2_U3069);
  nand ginst13263 (P2_R1161_U210, P2_R1161_U119, P2_R1161_U209);
  nand ginst13264 (P2_R1161_U211, P2_R1161_U195, P2_R1161_U22);
  nand ginst13265 (P2_R1161_U212, P2_U3069, P2_U3410);
  nand ginst13266 (P2_R1161_U213, P2_R1161_U120, P2_R1161_U211);
  or ginst13267 (P2_R1161_U214, P2_U3070, P2_U3407);
  nand ginst13268 (P2_R1161_U215, P2_R1161_U181, P2_R1161_U185);
  nand ginst13269 (P2_R1161_U216, P2_U3067, P2_U3395);
  not ginst13270 (P2_R1161_U217, P2_R1161_U45);
  nand ginst13271 (P2_R1161_U218, P2_R1161_U121, P2_R1161_U184);
  nand ginst13272 (P2_R1161_U219, P2_R1161_U180, P2_R1161_U45);
  nand ginst13273 (P2_R1161_U22, P2_U3070, P2_U3407);
  nand ginst13274 (P2_R1161_U220, P2_U3063, P2_U3398);
  not ginst13275 (P2_R1161_U221, P2_R1161_U44);
  or ginst13276 (P2_R1161_U222, P2_U3059, P2_U3401);
  nand ginst13277 (P2_R1161_U223, P2_R1161_U222, P2_R1161_U44);
  nand ginst13278 (P2_R1161_U224, P2_R1161_U123, P2_R1161_U223);
  nand ginst13279 (P2_R1161_U225, P2_R1161_U221, P2_R1161_U34);
  nand ginst13280 (P2_R1161_U226, P2_U3066, P2_U3404);
  nand ginst13281 (P2_R1161_U227, P2_R1161_U124, P2_R1161_U225);
  or ginst13282 (P2_R1161_U228, P2_U3059, P2_U3401);
  nand ginst13283 (P2_R1161_U229, P2_R1161_U181, P2_R1161_U184);
  not ginst13284 (P2_R1161_U23, P2_U3410);
  not ginst13285 (P2_R1161_U230, P2_R1161_U145);
  nand ginst13286 (P2_R1161_U231, P2_U3063, P2_U3398);
  nand ginst13287 (P2_R1161_U232, P2_R1161_U400, P2_R1161_U401, P2_R1161_U42, P2_R1161_U43);
  nand ginst13288 (P2_R1161_U233, P2_R1161_U42, P2_R1161_U43);
  nand ginst13289 (P2_R1161_U234, P2_U3067, P2_U3395);
  nand ginst13290 (P2_R1161_U235, P2_R1161_U125, P2_R1161_U233);
  or ginst13291 (P2_R1161_U236, P2_U3082, P2_U3416);
  or ginst13292 (P2_R1161_U237, P2_U3061, P2_U3419);
  nand ginst13293 (P2_R1161_U238, P2_R1161_U177, P2_R1161_U6);
  nand ginst13294 (P2_R1161_U239, P2_U3061, P2_U3419);
  not ginst13295 (P2_R1161_U24, P2_U3401);
  nand ginst13296 (P2_R1161_U240, P2_R1161_U171, P2_R1161_U238);
  or ginst13297 (P2_R1161_U241, P2_U3061, P2_U3419);
  nand ginst13298 (P2_R1161_U242, P2_R1161_U126, P2_R1161_U144);
  nand ginst13299 (P2_R1161_U243, P2_R1161_U240, P2_R1161_U241);
  not ginst13300 (P2_R1161_U244, P2_R1161_U167);
  or ginst13301 (P2_R1161_U245, P2_U3079, P2_U3428);
  or ginst13302 (P2_R1161_U246, P2_U3071, P2_U3425);
  nand ginst13303 (P2_R1161_U247, P2_R1161_U174, P2_R1161_U7);
  nand ginst13304 (P2_R1161_U248, P2_U3079, P2_U3428);
  nand ginst13305 (P2_R1161_U249, P2_R1161_U172, P2_R1161_U247);
  not ginst13306 (P2_R1161_U25, P2_U3059);
  or ginst13307 (P2_R1161_U250, P2_U3062, P2_U3422);
  or ginst13308 (P2_R1161_U251, P2_U3079, P2_U3428);
  nand ginst13309 (P2_R1161_U252, P2_R1161_U128, P2_R1161_U167);
  nand ginst13310 (P2_R1161_U253, P2_R1161_U249, P2_R1161_U251);
  not ginst13311 (P2_R1161_U254, P2_R1161_U166);
  or ginst13312 (P2_R1161_U255, P2_U3078, P2_U3431);
  nand ginst13313 (P2_R1161_U256, P2_R1161_U166, P2_R1161_U255);
  nand ginst13314 (P2_R1161_U257, P2_U3078, P2_U3431);
  not ginst13315 (P2_R1161_U258, P2_R1161_U164);
  or ginst13316 (P2_R1161_U259, P2_U3073, P2_U3434);
  not ginst13317 (P2_R1161_U26, P2_U3066);
  nand ginst13318 (P2_R1161_U260, P2_R1161_U164, P2_R1161_U259);
  nand ginst13319 (P2_R1161_U261, P2_U3073, P2_U3434);
  not ginst13320 (P2_R1161_U262, P2_R1161_U92);
  or ginst13321 (P2_R1161_U263, P2_U3068, P2_U3440);
  or ginst13322 (P2_R1161_U264, P2_U3072, P2_U3437);
  not ginst13323 (P2_R1161_U265, P2_R1161_U59);
  nand ginst13324 (P2_R1161_U266, P2_R1161_U59, P2_R1161_U60);
  nand ginst13325 (P2_R1161_U267, P2_R1161_U266, P2_U3068);
  nand ginst13326 (P2_R1161_U268, P2_R1161_U265, P2_U3440);
  nand ginst13327 (P2_R1161_U269, P2_R1161_U8, P2_R1161_U92);
  not ginst13328 (P2_R1161_U27, P2_U3395);
  not ginst13329 (P2_R1161_U270, P2_R1161_U162);
  or ginst13330 (P2_R1161_U271, P2_U3075, P2_U3903);
  or ginst13331 (P2_R1161_U272, P2_U3080, P2_U3445);
  or ginst13332 (P2_R1161_U273, P2_U3074, P2_U3902);
  not ginst13333 (P2_R1161_U274, P2_R1161_U80);
  nand ginst13334 (P2_R1161_U275, P2_R1161_U274, P2_U3903);
  nand ginst13335 (P2_R1161_U276, P2_R1161_U275, P2_R1161_U90);
  nand ginst13336 (P2_R1161_U277, P2_R1161_U80, P2_R1161_U81);
  nand ginst13337 (P2_R1161_U278, P2_R1161_U276, P2_R1161_U277);
  nand ginst13338 (P2_R1161_U279, P2_R1161_U175, P2_R1161_U9);
  not ginst13339 (P2_R1161_U28, P2_U3067);
  nand ginst13340 (P2_R1161_U280, P2_U3074, P2_U3902);
  nand ginst13341 (P2_R1161_U281, P2_R1161_U278, P2_R1161_U279);
  or ginst13342 (P2_R1161_U282, P2_U3081, P2_U3443);
  or ginst13343 (P2_R1161_U283, P2_U3074, P2_U3902);
  nand ginst13344 (P2_R1161_U284, P2_R1161_U131, P2_R1161_U162, P2_R1161_U273);
  nand ginst13345 (P2_R1161_U285, P2_R1161_U281, P2_R1161_U283);
  not ginst13346 (P2_R1161_U286, P2_R1161_U159);
  or ginst13347 (P2_R1161_U287, P2_U3060, P2_U3901);
  nand ginst13348 (P2_R1161_U288, P2_R1161_U159, P2_R1161_U287);
  nand ginst13349 (P2_R1161_U289, P2_U3060, P2_U3901);
  not ginst13350 (P2_R1161_U29, P2_U3387);
  not ginst13351 (P2_R1161_U290, P2_R1161_U157);
  or ginst13352 (P2_R1161_U291, P2_U3065, P2_U3900);
  nand ginst13353 (P2_R1161_U292, P2_R1161_U157, P2_R1161_U291);
  nand ginst13354 (P2_R1161_U293, P2_U3065, P2_U3900);
  not ginst13355 (P2_R1161_U294, P2_R1161_U155);
  or ginst13356 (P2_R1161_U295, P2_U3057, P2_U3898);
  nand ginst13357 (P2_R1161_U296, P2_R1161_U173, P2_R1161_U176);
  not ginst13358 (P2_R1161_U297, P2_R1161_U86);
  or ginst13359 (P2_R1161_U298, P2_U3064, P2_U3899);
  nand ginst13360 (P2_R1161_U299, P2_R1161_U155, P2_R1161_U168, P2_R1161_U298);
  not ginst13361 (P2_R1161_U30, P2_U3076);
  not ginst13362 (P2_R1161_U300, P2_R1161_U153);
  or ginst13363 (P2_R1161_U301, P2_U3052, P2_U3896);
  nand ginst13364 (P2_R1161_U302, P2_U3052, P2_U3896);
  not ginst13365 (P2_R1161_U303, P2_R1161_U151);
  nand ginst13366 (P2_R1161_U304, P2_R1161_U151, P2_U3895);
  not ginst13367 (P2_R1161_U305, P2_R1161_U149);
  nand ginst13368 (P2_R1161_U306, P2_R1161_U155, P2_R1161_U298);
  not ginst13369 (P2_R1161_U307, P2_R1161_U89);
  or ginst13370 (P2_R1161_U308, P2_U3057, P2_U3898);
  nand ginst13371 (P2_R1161_U309, P2_R1161_U308, P2_R1161_U89);
  nand ginst13372 (P2_R1161_U31, P2_U3076, P2_U3387);
  nand ginst13373 (P2_R1161_U310, P2_R1161_U154, P2_R1161_U173, P2_R1161_U309);
  nand ginst13374 (P2_R1161_U311, P2_R1161_U173, P2_R1161_U307);
  nand ginst13375 (P2_R1161_U312, P2_U3056, P2_U3897);
  nand ginst13376 (P2_R1161_U313, P2_R1161_U168, P2_R1161_U311, P2_R1161_U312);
  or ginst13377 (P2_R1161_U314, P2_U3057, P2_U3898);
  nand ginst13378 (P2_R1161_U315, P2_R1161_U162, P2_R1161_U282);
  not ginst13379 (P2_R1161_U316, P2_R1161_U91);
  nand ginst13380 (P2_R1161_U317, P2_R1161_U9, P2_R1161_U91);
  nand ginst13381 (P2_R1161_U318, P2_R1161_U135, P2_R1161_U317);
  nand ginst13382 (P2_R1161_U319, P2_R1161_U278, P2_R1161_U317);
  not ginst13383 (P2_R1161_U32, P2_U3398);
  nand ginst13384 (P2_R1161_U320, P2_R1161_U319, P2_R1161_U453);
  or ginst13385 (P2_R1161_U321, P2_U3080, P2_U3445);
  nand ginst13386 (P2_R1161_U322, P2_R1161_U321, P2_R1161_U91);
  nand ginst13387 (P2_R1161_U323, P2_R1161_U136, P2_R1161_U322);
  nand ginst13388 (P2_R1161_U324, P2_R1161_U316, P2_R1161_U80);
  nand ginst13389 (P2_R1161_U325, P2_U3075, P2_U3903);
  nand ginst13390 (P2_R1161_U326, P2_R1161_U137, P2_R1161_U324);
  or ginst13391 (P2_R1161_U327, P2_U3077, P2_U3392);
  not ginst13392 (P2_R1161_U328, P2_R1161_U161);
  or ginst13393 (P2_R1161_U329, P2_U3080, P2_U3445);
  not ginst13394 (P2_R1161_U33, P2_U3063);
  or ginst13395 (P2_R1161_U330, P2_U3072, P2_U3437);
  nand ginst13396 (P2_R1161_U331, P2_R1161_U330, P2_R1161_U92);
  nand ginst13397 (P2_R1161_U332, P2_R1161_U138, P2_R1161_U331);
  nand ginst13398 (P2_R1161_U333, P2_R1161_U262, P2_R1161_U59);
  nand ginst13399 (P2_R1161_U334, P2_U3068, P2_U3440);
  nand ginst13400 (P2_R1161_U335, P2_R1161_U139, P2_R1161_U333);
  or ginst13401 (P2_R1161_U336, P2_U3072, P2_U3437);
  nand ginst13402 (P2_R1161_U337, P2_R1161_U167, P2_R1161_U250);
  not ginst13403 (P2_R1161_U338, P2_R1161_U93);
  or ginst13404 (P2_R1161_U339, P2_U3071, P2_U3425);
  nand ginst13405 (P2_R1161_U34, P2_U3059, P2_U3401);
  nand ginst13406 (P2_R1161_U340, P2_R1161_U339, P2_R1161_U93);
  nand ginst13407 (P2_R1161_U341, P2_R1161_U140, P2_R1161_U340);
  nand ginst13408 (P2_R1161_U342, P2_R1161_U172, P2_R1161_U338);
  nand ginst13409 (P2_R1161_U343, P2_U3079, P2_U3428);
  nand ginst13410 (P2_R1161_U344, P2_R1161_U141, P2_R1161_U342);
  or ginst13411 (P2_R1161_U345, P2_U3071, P2_U3425);
  or ginst13412 (P2_R1161_U346, P2_U3082, P2_U3416);
  nand ginst13413 (P2_R1161_U347, P2_R1161_U346, P2_R1161_U40);
  nand ginst13414 (P2_R1161_U348, P2_R1161_U142, P2_R1161_U347);
  nand ginst13415 (P2_R1161_U349, P2_R1161_U171, P2_R1161_U206);
  not ginst13416 (P2_R1161_U35, P2_U3404);
  nand ginst13417 (P2_R1161_U350, P2_U3061, P2_U3419);
  nand ginst13418 (P2_R1161_U351, P2_R1161_U143, P2_R1161_U349);
  nand ginst13419 (P2_R1161_U352, P2_R1161_U171, P2_R1161_U207);
  nand ginst13420 (P2_R1161_U353, P2_R1161_U204, P2_R1161_U65);
  nand ginst13421 (P2_R1161_U354, P2_R1161_U214, P2_R1161_U22);
  nand ginst13422 (P2_R1161_U355, P2_R1161_U228, P2_R1161_U34);
  nand ginst13423 (P2_R1161_U356, P2_R1161_U180, P2_R1161_U231);
  nand ginst13424 (P2_R1161_U357, P2_R1161_U173, P2_R1161_U314);
  nand ginst13425 (P2_R1161_U358, P2_R1161_U176, P2_R1161_U298);
  nand ginst13426 (P2_R1161_U359, P2_R1161_U329, P2_R1161_U80);
  not ginst13427 (P2_R1161_U36, P2_U3413);
  nand ginst13428 (P2_R1161_U360, P2_R1161_U282, P2_R1161_U77);
  nand ginst13429 (P2_R1161_U361, P2_R1161_U336, P2_R1161_U59);
  nand ginst13430 (P2_R1161_U362, P2_R1161_U172, P2_R1161_U345);
  nand ginst13431 (P2_R1161_U363, P2_R1161_U250, P2_R1161_U68);
  nand ginst13432 (P2_R1161_U364, P2_U3053, P2_U3895);
  nand ginst13433 (P2_R1161_U365, P2_R1161_U168, P2_R1161_U296);
  nand ginst13434 (P2_R1161_U366, P2_R1161_U295, P2_U3056);
  nand ginst13435 (P2_R1161_U367, P2_R1161_U295, P2_U3897);
  nand ginst13436 (P2_R1161_U368, P2_R1161_U168, P2_R1161_U296, P2_R1161_U301);
  nand ginst13437 (P2_R1161_U369, P2_R1161_U133, P2_R1161_U155, P2_R1161_U168);
  not ginst13438 (P2_R1161_U37, P2_U3083);
  nand ginst13439 (P2_R1161_U370, P2_R1161_U297, P2_R1161_U301);
  nand ginst13440 (P2_R1161_U371, P2_R1161_U39, P2_U3082);
  nand ginst13441 (P2_R1161_U372, P2_R1161_U38, P2_U3416);
  nand ginst13442 (P2_R1161_U373, P2_R1161_U371, P2_R1161_U372);
  nand ginst13443 (P2_R1161_U374, P2_R1161_U352, P2_R1161_U40);
  nand ginst13444 (P2_R1161_U375, P2_R1161_U206, P2_R1161_U373);
  nand ginst13445 (P2_R1161_U376, P2_R1161_U36, P2_U3083);
  nand ginst13446 (P2_R1161_U377, P2_R1161_U37, P2_U3413);
  nand ginst13447 (P2_R1161_U378, P2_R1161_U376, P2_R1161_U377);
  nand ginst13448 (P2_R1161_U379, P2_R1161_U144, P2_R1161_U353);
  not ginst13449 (P2_R1161_U38, P2_U3082);
  nand ginst13450 (P2_R1161_U380, P2_R1161_U203, P2_R1161_U378);
  nand ginst13451 (P2_R1161_U381, P2_R1161_U23, P2_U3069);
  nand ginst13452 (P2_R1161_U382, P2_R1161_U21, P2_U3410);
  nand ginst13453 (P2_R1161_U383, P2_R1161_U19, P2_U3070);
  nand ginst13454 (P2_R1161_U384, P2_R1161_U20, P2_U3407);
  nand ginst13455 (P2_R1161_U385, P2_R1161_U383, P2_R1161_U384);
  nand ginst13456 (P2_R1161_U386, P2_R1161_U354, P2_R1161_U41);
  nand ginst13457 (P2_R1161_U387, P2_R1161_U195, P2_R1161_U385);
  nand ginst13458 (P2_R1161_U388, P2_R1161_U35, P2_U3066);
  nand ginst13459 (P2_R1161_U389, P2_R1161_U26, P2_U3404);
  not ginst13460 (P2_R1161_U39, P2_U3416);
  nand ginst13461 (P2_R1161_U390, P2_R1161_U24, P2_U3059);
  nand ginst13462 (P2_R1161_U391, P2_R1161_U25, P2_U3401);
  nand ginst13463 (P2_R1161_U392, P2_R1161_U390, P2_R1161_U391);
  nand ginst13464 (P2_R1161_U393, P2_R1161_U355, P2_R1161_U44);
  nand ginst13465 (P2_R1161_U394, P2_R1161_U221, P2_R1161_U392);
  nand ginst13466 (P2_R1161_U395, P2_R1161_U32, P2_U3063);
  nand ginst13467 (P2_R1161_U396, P2_R1161_U33, P2_U3398);
  nand ginst13468 (P2_R1161_U397, P2_R1161_U395, P2_R1161_U396);
  nand ginst13469 (P2_R1161_U398, P2_R1161_U145, P2_R1161_U356);
  nand ginst13470 (P2_R1161_U399, P2_R1161_U230, P2_R1161_U397);
  and ginst13471 (P2_R1161_U4, P2_R1161_U178, P2_R1161_U179);
  nand ginst13472 (P2_R1161_U40, P2_R1161_U205, P2_R1161_U65);
  nand ginst13473 (P2_R1161_U400, P2_R1161_U27, P2_U3067);
  nand ginst13474 (P2_R1161_U401, P2_R1161_U28, P2_U3395);
  nand ginst13475 (P2_R1161_U402, P2_R1161_U147, P2_U3054);
  nand ginst13476 (P2_R1161_U403, P2_R1161_U146, P2_U3904);
  nand ginst13477 (P2_R1161_U404, P2_R1161_U147, P2_U3054);
  nand ginst13478 (P2_R1161_U405, P2_R1161_U146, P2_U3904);
  nand ginst13479 (P2_R1161_U406, P2_R1161_U404, P2_R1161_U405);
  nand ginst13480 (P2_R1161_U407, P2_R1161_U148, P2_R1161_U149);
  nand ginst13481 (P2_R1161_U408, P2_R1161_U305, P2_R1161_U406);
  nand ginst13482 (P2_R1161_U409, P2_R1161_U88, P2_U3053);
  nand ginst13483 (P2_R1161_U41, P2_R1161_U117, P2_R1161_U193);
  nand ginst13484 (P2_R1161_U410, P2_R1161_U87, P2_U3895);
  nand ginst13485 (P2_R1161_U411, P2_R1161_U88, P2_U3053);
  nand ginst13486 (P2_R1161_U412, P2_R1161_U87, P2_U3895);
  nand ginst13487 (P2_R1161_U413, P2_R1161_U411, P2_R1161_U412);
  nand ginst13488 (P2_R1161_U414, P2_R1161_U150, P2_R1161_U151);
  nand ginst13489 (P2_R1161_U415, P2_R1161_U303, P2_R1161_U413);
  nand ginst13490 (P2_R1161_U416, P2_R1161_U46, P2_U3052);
  nand ginst13491 (P2_R1161_U417, P2_R1161_U47, P2_U3896);
  nand ginst13492 (P2_R1161_U418, P2_R1161_U46, P2_U3052);
  nand ginst13493 (P2_R1161_U419, P2_R1161_U47, P2_U3896);
  nand ginst13494 (P2_R1161_U42, P2_R1161_U182, P2_R1161_U183);
  nand ginst13495 (P2_R1161_U420, P2_R1161_U418, P2_R1161_U419);
  nand ginst13496 (P2_R1161_U421, P2_R1161_U152, P2_R1161_U153);
  nand ginst13497 (P2_R1161_U422, P2_R1161_U300, P2_R1161_U420);
  nand ginst13498 (P2_R1161_U423, P2_R1161_U49, P2_U3056);
  nand ginst13499 (P2_R1161_U424, P2_R1161_U48, P2_U3897);
  nand ginst13500 (P2_R1161_U425, P2_R1161_U50, P2_U3057);
  nand ginst13501 (P2_R1161_U426, P2_R1161_U51, P2_U3898);
  nand ginst13502 (P2_R1161_U427, P2_R1161_U425, P2_R1161_U426);
  nand ginst13503 (P2_R1161_U428, P2_R1161_U357, P2_R1161_U89);
  nand ginst13504 (P2_R1161_U429, P2_R1161_U307, P2_R1161_U427);
  nand ginst13505 (P2_R1161_U43, P2_U3077, P2_U3392);
  nand ginst13506 (P2_R1161_U430, P2_R1161_U52, P2_U3064);
  nand ginst13507 (P2_R1161_U431, P2_R1161_U53, P2_U3899);
  nand ginst13508 (P2_R1161_U432, P2_R1161_U430, P2_R1161_U431);
  nand ginst13509 (P2_R1161_U433, P2_R1161_U155, P2_R1161_U358);
  nand ginst13510 (P2_R1161_U434, P2_R1161_U294, P2_R1161_U432);
  nand ginst13511 (P2_R1161_U435, P2_R1161_U84, P2_U3065);
  nand ginst13512 (P2_R1161_U436, P2_R1161_U85, P2_U3900);
  nand ginst13513 (P2_R1161_U437, P2_R1161_U84, P2_U3065);
  nand ginst13514 (P2_R1161_U438, P2_R1161_U85, P2_U3900);
  nand ginst13515 (P2_R1161_U439, P2_R1161_U437, P2_R1161_U438);
  nand ginst13516 (P2_R1161_U44, P2_R1161_U122, P2_R1161_U219);
  nand ginst13517 (P2_R1161_U440, P2_R1161_U156, P2_R1161_U157);
  nand ginst13518 (P2_R1161_U441, P2_R1161_U290, P2_R1161_U439);
  nand ginst13519 (P2_R1161_U442, P2_R1161_U82, P2_U3060);
  nand ginst13520 (P2_R1161_U443, P2_R1161_U83, P2_U3901);
  nand ginst13521 (P2_R1161_U444, P2_R1161_U82, P2_U3060);
  nand ginst13522 (P2_R1161_U445, P2_R1161_U83, P2_U3901);
  nand ginst13523 (P2_R1161_U446, P2_R1161_U444, P2_R1161_U445);
  nand ginst13524 (P2_R1161_U447, P2_R1161_U158, P2_R1161_U159);
  nand ginst13525 (P2_R1161_U448, P2_R1161_U286, P2_R1161_U446);
  nand ginst13526 (P2_R1161_U449, P2_R1161_U54, P2_U3074);
  nand ginst13527 (P2_R1161_U45, P2_R1161_U215, P2_R1161_U216);
  nand ginst13528 (P2_R1161_U450, P2_R1161_U55, P2_U3902);
  nand ginst13529 (P2_R1161_U451, P2_R1161_U54, P2_U3074);
  nand ginst13530 (P2_R1161_U452, P2_R1161_U55, P2_U3902);
  nand ginst13531 (P2_R1161_U453, P2_R1161_U451, P2_R1161_U452);
  nand ginst13532 (P2_R1161_U454, P2_R1161_U81, P2_U3075);
  nand ginst13533 (P2_R1161_U455, P2_R1161_U90, P2_U3903);
  nand ginst13534 (P2_R1161_U456, P2_R1161_U161, P2_R1161_U182);
  nand ginst13535 (P2_R1161_U457, P2_R1161_U31, P2_R1161_U328);
  nand ginst13536 (P2_R1161_U458, P2_R1161_U78, P2_U3080);
  nand ginst13537 (P2_R1161_U459, P2_R1161_U79, P2_U3445);
  not ginst13538 (P2_R1161_U46, P2_U3896);
  nand ginst13539 (P2_R1161_U460, P2_R1161_U458, P2_R1161_U459);
  nand ginst13540 (P2_R1161_U461, P2_R1161_U359, P2_R1161_U91);
  nand ginst13541 (P2_R1161_U462, P2_R1161_U316, P2_R1161_U460);
  nand ginst13542 (P2_R1161_U463, P2_R1161_U75, P2_U3081);
  nand ginst13543 (P2_R1161_U464, P2_R1161_U76, P2_U3443);
  nand ginst13544 (P2_R1161_U465, P2_R1161_U463, P2_R1161_U464);
  nand ginst13545 (P2_R1161_U466, P2_R1161_U162, P2_R1161_U360);
  nand ginst13546 (P2_R1161_U467, P2_R1161_U270, P2_R1161_U465);
  nand ginst13547 (P2_R1161_U468, P2_R1161_U60, P2_U3068);
  nand ginst13548 (P2_R1161_U469, P2_R1161_U58, P2_U3440);
  not ginst13549 (P2_R1161_U47, P2_U3052);
  nand ginst13550 (P2_R1161_U470, P2_R1161_U56, P2_U3072);
  nand ginst13551 (P2_R1161_U471, P2_R1161_U57, P2_U3437);
  nand ginst13552 (P2_R1161_U472, P2_R1161_U470, P2_R1161_U471);
  nand ginst13553 (P2_R1161_U473, P2_R1161_U361, P2_R1161_U92);
  nand ginst13554 (P2_R1161_U474, P2_R1161_U262, P2_R1161_U472);
  nand ginst13555 (P2_R1161_U475, P2_R1161_U73, P2_U3073);
  nand ginst13556 (P2_R1161_U476, P2_R1161_U74, P2_U3434);
  nand ginst13557 (P2_R1161_U477, P2_R1161_U73, P2_U3073);
  nand ginst13558 (P2_R1161_U478, P2_R1161_U74, P2_U3434);
  nand ginst13559 (P2_R1161_U479, P2_R1161_U477, P2_R1161_U478);
  not ginst13560 (P2_R1161_U48, P2_U3056);
  nand ginst13561 (P2_R1161_U480, P2_R1161_U163, P2_R1161_U164);
  nand ginst13562 (P2_R1161_U481, P2_R1161_U258, P2_R1161_U479);
  nand ginst13563 (P2_R1161_U482, P2_R1161_U71, P2_U3078);
  nand ginst13564 (P2_R1161_U483, P2_R1161_U72, P2_U3431);
  nand ginst13565 (P2_R1161_U484, P2_R1161_U71, P2_U3078);
  nand ginst13566 (P2_R1161_U485, P2_R1161_U72, P2_U3431);
  nand ginst13567 (P2_R1161_U486, P2_R1161_U484, P2_R1161_U485);
  nand ginst13568 (P2_R1161_U487, P2_R1161_U165, P2_R1161_U166);
  nand ginst13569 (P2_R1161_U488, P2_R1161_U254, P2_R1161_U486);
  nand ginst13570 (P2_R1161_U489, P2_R1161_U61, P2_U3079);
  not ginst13571 (P2_R1161_U49, P2_U3897);
  nand ginst13572 (P2_R1161_U490, P2_R1161_U62, P2_U3428);
  nand ginst13573 (P2_R1161_U491, P2_R1161_U69, P2_U3071);
  nand ginst13574 (P2_R1161_U492, P2_R1161_U70, P2_U3425);
  nand ginst13575 (P2_R1161_U493, P2_R1161_U491, P2_R1161_U492);
  nand ginst13576 (P2_R1161_U494, P2_R1161_U362, P2_R1161_U93);
  nand ginst13577 (P2_R1161_U495, P2_R1161_U338, P2_R1161_U493);
  nand ginst13578 (P2_R1161_U496, P2_R1161_U66, P2_U3062);
  nand ginst13579 (P2_R1161_U497, P2_R1161_U67, P2_U3422);
  nand ginst13580 (P2_R1161_U498, P2_R1161_U496, P2_R1161_U497);
  nand ginst13581 (P2_R1161_U499, P2_R1161_U167, P2_R1161_U363);
  and ginst13582 (P2_R1161_U5, P2_R1161_U196, P2_R1161_U197);
  not ginst13583 (P2_R1161_U50, P2_U3898);
  nand ginst13584 (P2_R1161_U500, P2_R1161_U244, P2_R1161_U498);
  nand ginst13585 (P2_R1161_U501, P2_R1161_U63, P2_U3061);
  nand ginst13586 (P2_R1161_U502, P2_R1161_U64, P2_U3419);
  nand ginst13587 (P2_R1161_U503, P2_R1161_U29, P2_U3076);
  nand ginst13588 (P2_R1161_U504, P2_R1161_U30, P2_U3387);
  not ginst13589 (P2_R1161_U51, P2_U3057);
  not ginst13590 (P2_R1161_U52, P2_U3899);
  not ginst13591 (P2_R1161_U53, P2_U3064);
  not ginst13592 (P2_R1161_U54, P2_U3902);
  not ginst13593 (P2_R1161_U55, P2_U3074);
  not ginst13594 (P2_R1161_U56, P2_U3437);
  not ginst13595 (P2_R1161_U57, P2_U3072);
  not ginst13596 (P2_R1161_U58, P2_U3068);
  nand ginst13597 (P2_R1161_U59, P2_U3072, P2_U3437);
  and ginst13598 (P2_R1161_U6, P2_R1161_U236, P2_R1161_U237);
  not ginst13599 (P2_R1161_U60, P2_U3440);
  not ginst13600 (P2_R1161_U61, P2_U3428);
  not ginst13601 (P2_R1161_U62, P2_U3079);
  not ginst13602 (P2_R1161_U63, P2_U3419);
  not ginst13603 (P2_R1161_U64, P2_U3061);
  nand ginst13604 (P2_R1161_U65, P2_U3083, P2_U3413);
  not ginst13605 (P2_R1161_U66, P2_U3422);
  not ginst13606 (P2_R1161_U67, P2_U3062);
  nand ginst13607 (P2_R1161_U68, P2_U3062, P2_U3422);
  not ginst13608 (P2_R1161_U69, P2_U3425);
  and ginst13609 (P2_R1161_U7, P2_R1161_U245, P2_R1161_U246);
  not ginst13610 (P2_R1161_U70, P2_U3071);
  not ginst13611 (P2_R1161_U71, P2_U3431);
  not ginst13612 (P2_R1161_U72, P2_U3078);
  not ginst13613 (P2_R1161_U73, P2_U3434);
  not ginst13614 (P2_R1161_U74, P2_U3073);
  not ginst13615 (P2_R1161_U75, P2_U3443);
  not ginst13616 (P2_R1161_U76, P2_U3081);
  nand ginst13617 (P2_R1161_U77, P2_U3081, P2_U3443);
  not ginst13618 (P2_R1161_U78, P2_U3445);
  not ginst13619 (P2_R1161_U79, P2_U3080);
  and ginst13620 (P2_R1161_U8, P2_R1161_U263, P2_R1161_U264);
  nand ginst13621 (P2_R1161_U80, P2_U3080, P2_U3445);
  not ginst13622 (P2_R1161_U81, P2_U3903);
  not ginst13623 (P2_R1161_U82, P2_U3901);
  not ginst13624 (P2_R1161_U83, P2_U3060);
  not ginst13625 (P2_R1161_U84, P2_U3900);
  not ginst13626 (P2_R1161_U85, P2_U3065);
  nand ginst13627 (P2_R1161_U86, P2_U3056, P2_U3897);
  not ginst13628 (P2_R1161_U87, P2_U3053);
  not ginst13629 (P2_R1161_U88, P2_U3895);
  nand ginst13630 (P2_R1161_U89, P2_R1161_U176, P2_R1161_U306);
  and ginst13631 (P2_R1161_U9, P2_R1161_U271, P2_R1161_U272);
  not ginst13632 (P2_R1161_U90, P2_U3075);
  nand ginst13633 (P2_R1161_U91, P2_R1161_U315, P2_R1161_U77);
  nand ginst13634 (P2_R1161_U92, P2_R1161_U260, P2_R1161_U261);
  nand ginst13635 (P2_R1161_U93, P2_R1161_U337, P2_R1161_U68);
  nand ginst13636 (P2_R1161_U94, P2_R1161_U456, P2_R1161_U457);
  nand ginst13637 (P2_R1161_U95, P2_R1161_U503, P2_R1161_U504);
  nand ginst13638 (P2_R1161_U96, P2_R1161_U374, P2_R1161_U375);
  nand ginst13639 (P2_R1161_U97, P2_R1161_U379, P2_R1161_U380);
  nand ginst13640 (P2_R1161_U98, P2_R1161_U386, P2_R1161_U387);
  nand ginst13641 (P2_R1161_U99, P2_R1161_U393, P2_R1161_U394);
  and ginst13642 (P2_R1179_U10, P2_R1179_U194, P2_R1179_U281);
  nand ginst13643 (P2_R1179_U100, P2_R1179_U424, P2_R1179_U425);
  nand ginst13644 (P2_R1179_U101, P2_R1179_U440, P2_R1179_U441);
  nand ginst13645 (P2_R1179_U102, P2_R1179_U445, P2_R1179_U446);
  nand ginst13646 (P2_R1179_U103, P2_R1179_U450, P2_R1179_U451);
  nand ginst13647 (P2_R1179_U104, P2_R1179_U455, P2_R1179_U456);
  nand ginst13648 (P2_R1179_U105, P2_R1179_U460, P2_R1179_U461);
  nand ginst13649 (P2_R1179_U106, P2_R1179_U476, P2_R1179_U477);
  nand ginst13650 (P2_R1179_U107, P2_R1179_U481, P2_R1179_U482);
  nand ginst13651 (P2_R1179_U108, P2_R1179_U364, P2_R1179_U365);
  nand ginst13652 (P2_R1179_U109, P2_R1179_U373, P2_R1179_U374);
  and ginst13653 (P2_R1179_U11, P2_R1179_U282, P2_R1179_U283);
  nand ginst13654 (P2_R1179_U110, P2_R1179_U380, P2_R1179_U381);
  nand ginst13655 (P2_R1179_U111, P2_R1179_U384, P2_R1179_U385);
  nand ginst13656 (P2_R1179_U112, P2_R1179_U393, P2_R1179_U394);
  nand ginst13657 (P2_R1179_U113, P2_R1179_U414, P2_R1179_U415);
  nand ginst13658 (P2_R1179_U114, P2_R1179_U431, P2_R1179_U432);
  nand ginst13659 (P2_R1179_U115, P2_R1179_U435, P2_R1179_U436);
  nand ginst13660 (P2_R1179_U116, P2_R1179_U467, P2_R1179_U468);
  nand ginst13661 (P2_R1179_U117, P2_R1179_U471, P2_R1179_U472);
  nand ginst13662 (P2_R1179_U118, P2_R1179_U488, P2_R1179_U489);
  and ginst13663 (P2_R1179_U119, P2_R1179_U196, P2_R1179_U206);
  and ginst13664 (P2_R1179_U12, P2_R1179_U195, P2_R1179_U299);
  and ginst13665 (P2_R1179_U120, P2_R1179_U208, P2_R1179_U209);
  and ginst13666 (P2_R1179_U121, P2_R1179_U13, P2_R1179_U14);
  and ginst13667 (P2_R1179_U122, P2_R1179_U222, P2_R1179_U340);
  and ginst13668 (P2_R1179_U123, P2_R1179_U122, P2_R1179_U342);
  and ginst13669 (P2_R1179_U124, P2_R1179_U27, P2_R1179_U366, P2_R1179_U367);
  and ginst13670 (P2_R1179_U125, P2_R1179_U198, P2_R1179_U370);
  and ginst13671 (P2_R1179_U126, P2_R1179_U237, P2_R1179_U6);
  and ginst13672 (P2_R1179_U127, P2_R1179_U197, P2_R1179_U377);
  and ginst13673 (P2_R1179_U128, P2_R1179_U35, P2_R1179_U386, P2_R1179_U387);
  and ginst13674 (P2_R1179_U129, P2_R1179_U196, P2_R1179_U390);
  and ginst13675 (P2_R1179_U13, P2_R1179_U197, P2_R1179_U210, P2_R1179_U215);
  and ginst13676 (P2_R1179_U130, P2_R1179_U15, P2_R1179_U251);
  and ginst13677 (P2_R1179_U131, P2_R1179_U252, P2_R1179_U343);
  and ginst13678 (P2_R1179_U132, P2_R1179_U262, P2_R1179_U8);
  and ginst13679 (P2_R1179_U133, P2_R1179_U10, P2_R1179_U286);
  and ginst13680 (P2_R1179_U134, P2_R1179_U301, P2_R1179_U302);
  and ginst13681 (P2_R1179_U135, P2_R1179_U303, P2_R1179_U397);
  and ginst13682 (P2_R1179_U136, P2_R1179_U16, P2_R1179_U301, P2_R1179_U302, P2_R1179_U304);
  and ginst13683 (P2_R1179_U137, P2_R1179_U165, P2_R1179_U359);
  nand ginst13684 (P2_R1179_U138, P2_R1179_U402, P2_R1179_U403);
  and ginst13685 (P2_R1179_U139, P2_R1179_U407, P2_R1179_U408, P2_R1179_U53);
  and ginst13686 (P2_R1179_U14, P2_R1179_U198, P2_R1179_U220);
  and ginst13687 (P2_R1179_U140, P2_R1179_U195, P2_R1179_U411);
  nand ginst13688 (P2_R1179_U141, P2_R1179_U416, P2_R1179_U417);
  nand ginst13689 (P2_R1179_U142, P2_R1179_U421, P2_R1179_U422);
  and ginst13690 (P2_R1179_U143, P2_R1179_U11, P2_R1179_U313);
  and ginst13691 (P2_R1179_U144, P2_R1179_U194, P2_R1179_U428);
  nand ginst13692 (P2_R1179_U145, P2_R1179_U437, P2_R1179_U438);
  nand ginst13693 (P2_R1179_U146, P2_R1179_U442, P2_R1179_U443);
  nand ginst13694 (P2_R1179_U147, P2_R1179_U447, P2_R1179_U448);
  nand ginst13695 (P2_R1179_U148, P2_R1179_U452, P2_R1179_U453);
  nand ginst13696 (P2_R1179_U149, P2_R1179_U457, P2_R1179_U458);
  and ginst13697 (P2_R1179_U15, P2_R1179_U192, P2_R1179_U224, P2_R1179_U244);
  and ginst13698 (P2_R1179_U150, P2_R1179_U324, P2_R1179_U9);
  and ginst13699 (P2_R1179_U151, P2_R1179_U193, P2_R1179_U464);
  nand ginst13700 (P2_R1179_U152, P2_R1179_U473, P2_R1179_U474);
  nand ginst13701 (P2_R1179_U153, P2_R1179_U478, P2_R1179_U479);
  and ginst13702 (P2_R1179_U154, P2_R1179_U333, P2_R1179_U7);
  and ginst13703 (P2_R1179_U155, P2_R1179_U192, P2_R1179_U485);
  and ginst13704 (P2_R1179_U156, P2_R1179_U362, P2_R1179_U363);
  nand ginst13705 (P2_R1179_U157, P2_R1179_U123, P2_R1179_U341);
  and ginst13706 (P2_R1179_U158, P2_R1179_U371, P2_R1179_U372);
  and ginst13707 (P2_R1179_U159, P2_R1179_U378, P2_R1179_U379);
  and ginst13708 (P2_R1179_U16, P2_R1179_U398, P2_R1179_U399);
  and ginst13709 (P2_R1179_U160, P2_R1179_U382, P2_R1179_U383);
  nand ginst13710 (P2_R1179_U161, P2_R1179_U120, P2_R1179_U344);
  and ginst13711 (P2_R1179_U162, P2_R1179_U391, P2_R1179_U392);
  not ginst13712 (P2_R1179_U163, P2_U3904);
  not ginst13713 (P2_R1179_U164, P2_U3054);
  and ginst13714 (P2_R1179_U165, P2_R1179_U400, P2_R1179_U401);
  nand ginst13715 (P2_R1179_U166, P2_R1179_U134, P2_R1179_U360);
  and ginst13716 (P2_R1179_U167, P2_R1179_U412, P2_R1179_U413);
  nand ginst13717 (P2_R1179_U168, P2_R1179_U292, P2_R1179_U293);
  nand ginst13718 (P2_R1179_U169, P2_R1179_U288, P2_R1179_U289);
  nand ginst13719 (P2_R1179_U17, P2_R1179_U331, P2_R1179_U334);
  and ginst13720 (P2_R1179_U170, P2_R1179_U429, P2_R1179_U430);
  and ginst13721 (P2_R1179_U171, P2_R1179_U433, P2_R1179_U434);
  nand ginst13722 (P2_R1179_U172, P2_R1179_U278, P2_R1179_U279);
  nand ginst13723 (P2_R1179_U173, P2_R1179_U274, P2_R1179_U275);
  not ginst13724 (P2_R1179_U174, P2_U3392);
  nand ginst13725 (P2_R1179_U175, P2_R1179_U97, P2_U3387);
  nand ginst13726 (P2_R1179_U176, P2_R1179_U187, P2_R1179_U271, P2_R1179_U339);
  not ginst13727 (P2_R1179_U177, P2_U3443);
  nand ginst13728 (P2_R1179_U178, P2_R1179_U268, P2_R1179_U269);
  nand ginst13729 (P2_R1179_U179, P2_R1179_U264, P2_R1179_U265);
  nand ginst13730 (P2_R1179_U18, P2_R1179_U322, P2_R1179_U325);
  and ginst13731 (P2_R1179_U180, P2_R1179_U465, P2_R1179_U466);
  and ginst13732 (P2_R1179_U181, P2_R1179_U469, P2_R1179_U470);
  nand ginst13733 (P2_R1179_U182, P2_R1179_U254, P2_R1179_U255);
  nand ginst13734 (P2_R1179_U183, P2_R1179_U131, P2_R1179_U353);
  nand ginst13735 (P2_R1179_U184, P2_R1179_U351, P2_R1179_U62);
  and ginst13736 (P2_R1179_U185, P2_R1179_U486, P2_R1179_U487);
  nand ginst13737 (P2_R1179_U186, P2_R1179_U135, P2_R1179_U166);
  nand ginst13738 (P2_R1179_U187, P2_R1179_U177, P2_R1179_U178);
  nand ginst13739 (P2_R1179_U188, P2_R1179_U174, P2_R1179_U175);
  not ginst13740 (P2_R1179_U189, P2_R1179_U53);
  nand ginst13741 (P2_R1179_U19, P2_R1179_U311, P2_R1179_U314);
  not ginst13742 (P2_R1179_U190, P2_R1179_U35);
  not ginst13743 (P2_R1179_U191, P2_R1179_U27);
  nand ginst13744 (P2_R1179_U192, P2_R1179_U57, P2_U3419);
  nand ginst13745 (P2_R1179_U193, P2_R1179_U69, P2_U3434);
  nand ginst13746 (P2_R1179_U194, P2_R1179_U83, P2_U3901);
  nand ginst13747 (P2_R1179_U195, P2_R1179_U52, P2_U3897);
  nand ginst13748 (P2_R1179_U196, P2_R1179_U34, P2_U3395);
  nand ginst13749 (P2_R1179_U197, P2_R1179_U42, P2_U3404);
  nand ginst13750 (P2_R1179_U198, P2_R1179_U26, P2_U3410);
  not ginst13751 (P2_R1179_U199, P2_R1179_U71);
  nand ginst13752 (P2_R1179_U20, P2_R1179_U305, P2_R1179_U357);
  not ginst13753 (P2_R1179_U200, P2_R1179_U85);
  not ginst13754 (P2_R1179_U201, P2_R1179_U44);
  not ginst13755 (P2_R1179_U202, P2_R1179_U59);
  not ginst13756 (P2_R1179_U203, P2_R1179_U175);
  nand ginst13757 (P2_R1179_U204, P2_R1179_U175, P2_U3077);
  not ginst13758 (P2_R1179_U205, P2_R1179_U50);
  nand ginst13759 (P2_R1179_U206, P2_R1179_U36, P2_U3398);
  nand ginst13760 (P2_R1179_U207, P2_R1179_U35, P2_R1179_U36);
  nand ginst13761 (P2_R1179_U208, P2_R1179_U207, P2_R1179_U40);
  nand ginst13762 (P2_R1179_U209, P2_R1179_U190, P2_U3063);
  nand ginst13763 (P2_R1179_U21, P2_R1179_U137, P2_R1179_U186);
  nand ginst13764 (P2_R1179_U210, P2_R1179_U41, P2_U3407);
  nand ginst13765 (P2_R1179_U211, P2_R1179_U30, P2_U3070);
  nand ginst13766 (P2_R1179_U212, P2_R1179_U29, P2_U3066);
  nand ginst13767 (P2_R1179_U213, P2_R1179_U197, P2_R1179_U201);
  nand ginst13768 (P2_R1179_U214, P2_R1179_U213, P2_R1179_U6);
  nand ginst13769 (P2_R1179_U215, P2_R1179_U43, P2_U3401);
  nand ginst13770 (P2_R1179_U216, P2_R1179_U41, P2_U3407);
  nand ginst13771 (P2_R1179_U217, P2_R1179_U13, P2_R1179_U161);
  not ginst13772 (P2_R1179_U218, P2_R1179_U45);
  not ginst13773 (P2_R1179_U219, P2_R1179_U48);
  nand ginst13774 (P2_R1179_U22, P2_R1179_U242, P2_R1179_U347);
  nand ginst13775 (P2_R1179_U220, P2_R1179_U28, P2_U3413);
  nand ginst13776 (P2_R1179_U221, P2_R1179_U27, P2_R1179_U28);
  nand ginst13777 (P2_R1179_U222, P2_R1179_U191, P2_U3083);
  not ginst13778 (P2_R1179_U223, P2_R1179_U157);
  nand ginst13779 (P2_R1179_U224, P2_R1179_U47, P2_U3416);
  nand ginst13780 (P2_R1179_U225, P2_R1179_U224, P2_R1179_U59);
  nand ginst13781 (P2_R1179_U226, P2_R1179_U219, P2_R1179_U27);
  nand ginst13782 (P2_R1179_U227, P2_R1179_U125, P2_R1179_U226);
  nand ginst13783 (P2_R1179_U228, P2_R1179_U198, P2_R1179_U48);
  nand ginst13784 (P2_R1179_U229, P2_R1179_U124, P2_R1179_U228);
  nand ginst13785 (P2_R1179_U23, P2_R1179_U235, P2_R1179_U238);
  nand ginst13786 (P2_R1179_U230, P2_R1179_U198, P2_R1179_U27);
  nand ginst13787 (P2_R1179_U231, P2_R1179_U161, P2_R1179_U215);
  not ginst13788 (P2_R1179_U232, P2_R1179_U49);
  nand ginst13789 (P2_R1179_U233, P2_R1179_U29, P2_U3066);
  nand ginst13790 (P2_R1179_U234, P2_R1179_U232, P2_R1179_U233);
  nand ginst13791 (P2_R1179_U235, P2_R1179_U127, P2_R1179_U234);
  nand ginst13792 (P2_R1179_U236, P2_R1179_U197, P2_R1179_U49);
  nand ginst13793 (P2_R1179_U237, P2_R1179_U41, P2_U3407);
  nand ginst13794 (P2_R1179_U238, P2_R1179_U126, P2_R1179_U236);
  nand ginst13795 (P2_R1179_U239, P2_R1179_U29, P2_U3066);
  nand ginst13796 (P2_R1179_U24, P2_R1179_U227, P2_R1179_U229);
  nand ginst13797 (P2_R1179_U240, P2_R1179_U197, P2_R1179_U239);
  nand ginst13798 (P2_R1179_U241, P2_R1179_U215, P2_R1179_U44);
  nand ginst13799 (P2_R1179_U242, P2_R1179_U129, P2_R1179_U348);
  nand ginst13800 (P2_R1179_U243, P2_R1179_U196, P2_R1179_U35);
  nand ginst13801 (P2_R1179_U244, P2_R1179_U56, P2_U3422);
  nand ginst13802 (P2_R1179_U245, P2_R1179_U60, P2_U3062);
  nand ginst13803 (P2_R1179_U246, P2_R1179_U58, P2_U3061);
  nand ginst13804 (P2_R1179_U247, P2_R1179_U192, P2_R1179_U202);
  nand ginst13805 (P2_R1179_U248, P2_R1179_U247, P2_R1179_U7);
  nand ginst13806 (P2_R1179_U249, P2_R1179_U56, P2_U3422);
  nand ginst13807 (P2_R1179_U25, P2_R1179_U175, P2_R1179_U337);
  not ginst13808 (P2_R1179_U250, P2_R1179_U62);
  nand ginst13809 (P2_R1179_U251, P2_R1179_U55, P2_U3425);
  nand ginst13810 (P2_R1179_U252, P2_R1179_U61, P2_U3071);
  nand ginst13811 (P2_R1179_U253, P2_R1179_U64, P2_U3428);
  nand ginst13812 (P2_R1179_U254, P2_R1179_U183, P2_R1179_U253);
  nand ginst13813 (P2_R1179_U255, P2_R1179_U63, P2_U3079);
  not ginst13814 (P2_R1179_U256, P2_R1179_U182);
  nand ginst13815 (P2_R1179_U257, P2_R1179_U68, P2_U3437);
  nand ginst13816 (P2_R1179_U258, P2_R1179_U65, P2_U3072);
  nand ginst13817 (P2_R1179_U259, P2_R1179_U66, P2_U3073);
  not ginst13818 (P2_R1179_U26, P2_U3069);
  nand ginst13819 (P2_R1179_U260, P2_R1179_U199, P2_R1179_U8);
  nand ginst13820 (P2_R1179_U261, P2_R1179_U260, P2_R1179_U9);
  nand ginst13821 (P2_R1179_U262, P2_R1179_U70, P2_U3431);
  nand ginst13822 (P2_R1179_U263, P2_R1179_U68, P2_U3437);
  nand ginst13823 (P2_R1179_U264, P2_R1179_U132, P2_R1179_U182);
  nand ginst13824 (P2_R1179_U265, P2_R1179_U261, P2_R1179_U263);
  not ginst13825 (P2_R1179_U266, P2_R1179_U179);
  nand ginst13826 (P2_R1179_U267, P2_R1179_U73, P2_U3440);
  nand ginst13827 (P2_R1179_U268, P2_R1179_U179, P2_R1179_U267);
  nand ginst13828 (P2_R1179_U269, P2_R1179_U72, P2_U3068);
  nand ginst13829 (P2_R1179_U27, P2_R1179_U32, P2_U3069);
  not ginst13830 (P2_R1179_U270, P2_R1179_U178);
  nand ginst13831 (P2_R1179_U271, P2_R1179_U178, P2_U3081);
  not ginst13832 (P2_R1179_U272, P2_R1179_U176);
  nand ginst13833 (P2_R1179_U273, P2_R1179_U76, P2_U3445);
  nand ginst13834 (P2_R1179_U274, P2_R1179_U176, P2_R1179_U273);
  nand ginst13835 (P2_R1179_U275, P2_R1179_U75, P2_U3080);
  not ginst13836 (P2_R1179_U276, P2_R1179_U173);
  nand ginst13837 (P2_R1179_U277, P2_R1179_U78, P2_U3903);
  nand ginst13838 (P2_R1179_U278, P2_R1179_U173, P2_R1179_U277);
  nand ginst13839 (P2_R1179_U279, P2_R1179_U77, P2_U3075);
  not ginst13840 (P2_R1179_U28, P2_U3083);
  not ginst13841 (P2_R1179_U280, P2_R1179_U172);
  nand ginst13842 (P2_R1179_U281, P2_R1179_U82, P2_U3900);
  nand ginst13843 (P2_R1179_U282, P2_R1179_U79, P2_U3065);
  nand ginst13844 (P2_R1179_U283, P2_R1179_U80, P2_U3060);
  nand ginst13845 (P2_R1179_U284, P2_R1179_U10, P2_R1179_U200);
  nand ginst13846 (P2_R1179_U285, P2_R1179_U11, P2_R1179_U284);
  nand ginst13847 (P2_R1179_U286, P2_R1179_U84, P2_U3902);
  nand ginst13848 (P2_R1179_U287, P2_R1179_U82, P2_U3900);
  nand ginst13849 (P2_R1179_U288, P2_R1179_U133, P2_R1179_U172);
  nand ginst13850 (P2_R1179_U289, P2_R1179_U285, P2_R1179_U287);
  not ginst13851 (P2_R1179_U29, P2_U3404);
  not ginst13852 (P2_R1179_U290, P2_R1179_U169);
  nand ginst13853 (P2_R1179_U291, P2_R1179_U87, P2_U3899);
  nand ginst13854 (P2_R1179_U292, P2_R1179_U169, P2_R1179_U291);
  nand ginst13855 (P2_R1179_U293, P2_R1179_U86, P2_U3064);
  not ginst13856 (P2_R1179_U294, P2_R1179_U168);
  nand ginst13857 (P2_R1179_U295, P2_R1179_U89, P2_U3898);
  nand ginst13858 (P2_R1179_U296, P2_R1179_U168, P2_R1179_U295);
  nand ginst13859 (P2_R1179_U297, P2_R1179_U88, P2_U3057);
  not ginst13860 (P2_R1179_U298, P2_R1179_U93);
  nand ginst13861 (P2_R1179_U299, P2_R1179_U54, P2_U3896);
  not ginst13862 (P2_R1179_U30, P2_U3407);
  nand ginst13863 (P2_R1179_U300, P2_R1179_U53, P2_R1179_U54);
  nand ginst13864 (P2_R1179_U301, P2_R1179_U300, P2_R1179_U91);
  nand ginst13865 (P2_R1179_U302, P2_R1179_U189, P2_U3052);
  nand ginst13866 (P2_R1179_U303, P2_R1179_U92, P2_U3895);
  nand ginst13867 (P2_R1179_U304, P2_R1179_U51, P2_U3053);
  nand ginst13868 (P2_R1179_U305, P2_R1179_U140, P2_R1179_U355);
  nand ginst13869 (P2_R1179_U306, P2_R1179_U195, P2_R1179_U53);
  nand ginst13870 (P2_R1179_U307, P2_R1179_U172, P2_R1179_U286);
  not ginst13871 (P2_R1179_U308, P2_R1179_U94);
  nand ginst13872 (P2_R1179_U309, P2_R1179_U80, P2_U3060);
  not ginst13873 (P2_R1179_U31, P2_U3401);
  nand ginst13874 (P2_R1179_U310, P2_R1179_U308, P2_R1179_U309);
  nand ginst13875 (P2_R1179_U311, P2_R1179_U144, P2_R1179_U310);
  nand ginst13876 (P2_R1179_U312, P2_R1179_U194, P2_R1179_U94);
  nand ginst13877 (P2_R1179_U313, P2_R1179_U82, P2_U3900);
  nand ginst13878 (P2_R1179_U314, P2_R1179_U143, P2_R1179_U312);
  nand ginst13879 (P2_R1179_U315, P2_R1179_U80, P2_U3060);
  nand ginst13880 (P2_R1179_U316, P2_R1179_U194, P2_R1179_U315);
  nand ginst13881 (P2_R1179_U317, P2_R1179_U286, P2_R1179_U85);
  nand ginst13882 (P2_R1179_U318, P2_R1179_U182, P2_R1179_U262);
  not ginst13883 (P2_R1179_U319, P2_R1179_U95);
  not ginst13884 (P2_R1179_U32, P2_U3410);
  nand ginst13885 (P2_R1179_U320, P2_R1179_U66, P2_U3073);
  nand ginst13886 (P2_R1179_U321, P2_R1179_U319, P2_R1179_U320);
  nand ginst13887 (P2_R1179_U322, P2_R1179_U151, P2_R1179_U321);
  nand ginst13888 (P2_R1179_U323, P2_R1179_U193, P2_R1179_U95);
  nand ginst13889 (P2_R1179_U324, P2_R1179_U68, P2_U3437);
  nand ginst13890 (P2_R1179_U325, P2_R1179_U150, P2_R1179_U323);
  nand ginst13891 (P2_R1179_U326, P2_R1179_U66, P2_U3073);
  nand ginst13892 (P2_R1179_U327, P2_R1179_U193, P2_R1179_U326);
  nand ginst13893 (P2_R1179_U328, P2_R1179_U262, P2_R1179_U71);
  nand ginst13894 (P2_R1179_U329, P2_R1179_U58, P2_U3061);
  not ginst13895 (P2_R1179_U33, P2_U3413);
  nand ginst13896 (P2_R1179_U330, P2_R1179_U329, P2_R1179_U350);
  nand ginst13897 (P2_R1179_U331, P2_R1179_U155, P2_R1179_U330);
  nand ginst13898 (P2_R1179_U332, P2_R1179_U192, P2_R1179_U96);
  nand ginst13899 (P2_R1179_U333, P2_R1179_U56, P2_U3422);
  nand ginst13900 (P2_R1179_U334, P2_R1179_U154, P2_R1179_U332);
  nand ginst13901 (P2_R1179_U335, P2_R1179_U58, P2_U3061);
  nand ginst13902 (P2_R1179_U336, P2_R1179_U192, P2_R1179_U335);
  nand ginst13903 (P2_R1179_U337, P2_R1179_U38, P2_U3076);
  nand ginst13904 (P2_R1179_U338, P2_R1179_U174, P2_U3077);
  nand ginst13905 (P2_R1179_U339, P2_R1179_U177, P2_U3081);
  not ginst13906 (P2_R1179_U34, P2_U3067);
  nand ginst13907 (P2_R1179_U340, P2_R1179_U221, P2_R1179_U33);
  nand ginst13908 (P2_R1179_U341, P2_R1179_U121, P2_R1179_U161);
  nand ginst13909 (P2_R1179_U342, P2_R1179_U14, P2_R1179_U218);
  nand ginst13910 (P2_R1179_U343, P2_R1179_U250, P2_R1179_U251);
  nand ginst13911 (P2_R1179_U344, P2_R1179_U119, P2_R1179_U50);
  not ginst13912 (P2_R1179_U345, P2_R1179_U161);
  nand ginst13913 (P2_R1179_U346, P2_R1179_U196, P2_R1179_U50);
  nand ginst13914 (P2_R1179_U347, P2_R1179_U128, P2_R1179_U346);
  nand ginst13915 (P2_R1179_U348, P2_R1179_U205, P2_R1179_U35);
  nand ginst13916 (P2_R1179_U349, P2_R1179_U157, P2_R1179_U224);
  nand ginst13917 (P2_R1179_U35, P2_R1179_U37, P2_U3067);
  not ginst13918 (P2_R1179_U350, P2_R1179_U96);
  nand ginst13919 (P2_R1179_U351, P2_R1179_U15, P2_R1179_U157);
  not ginst13920 (P2_R1179_U352, P2_R1179_U184);
  nand ginst13921 (P2_R1179_U353, P2_R1179_U130, P2_R1179_U157);
  not ginst13922 (P2_R1179_U354, P2_R1179_U183);
  nand ginst13923 (P2_R1179_U355, P2_R1179_U298, P2_R1179_U53);
  nand ginst13924 (P2_R1179_U356, P2_R1179_U195, P2_R1179_U93);
  nand ginst13925 (P2_R1179_U357, P2_R1179_U139, P2_R1179_U356);
  nand ginst13926 (P2_R1179_U358, P2_R1179_U12, P2_R1179_U93);
  nand ginst13927 (P2_R1179_U359, P2_R1179_U136, P2_R1179_U358);
  not ginst13928 (P2_R1179_U36, P2_U3063);
  nand ginst13929 (P2_R1179_U360, P2_R1179_U12, P2_R1179_U93);
  not ginst13930 (P2_R1179_U361, P2_R1179_U166);
  nand ginst13931 (P2_R1179_U362, P2_R1179_U47, P2_U3416);
  nand ginst13932 (P2_R1179_U363, P2_R1179_U46, P2_U3082);
  nand ginst13933 (P2_R1179_U364, P2_R1179_U157, P2_R1179_U225);
  nand ginst13934 (P2_R1179_U365, P2_R1179_U156, P2_R1179_U223);
  nand ginst13935 (P2_R1179_U366, P2_R1179_U28, P2_U3413);
  nand ginst13936 (P2_R1179_U367, P2_R1179_U33, P2_U3083);
  nand ginst13937 (P2_R1179_U368, P2_R1179_U28, P2_U3413);
  nand ginst13938 (P2_R1179_U369, P2_R1179_U33, P2_U3083);
  not ginst13939 (P2_R1179_U37, P2_U3395);
  nand ginst13940 (P2_R1179_U370, P2_R1179_U368, P2_R1179_U369);
  nand ginst13941 (P2_R1179_U371, P2_R1179_U26, P2_U3410);
  nand ginst13942 (P2_R1179_U372, P2_R1179_U32, P2_U3069);
  nand ginst13943 (P2_R1179_U373, P2_R1179_U230, P2_R1179_U48);
  nand ginst13944 (P2_R1179_U374, P2_R1179_U158, P2_R1179_U219);
  nand ginst13945 (P2_R1179_U375, P2_R1179_U41, P2_U3407);
  nand ginst13946 (P2_R1179_U376, P2_R1179_U30, P2_U3070);
  nand ginst13947 (P2_R1179_U377, P2_R1179_U375, P2_R1179_U376);
  nand ginst13948 (P2_R1179_U378, P2_R1179_U42, P2_U3404);
  nand ginst13949 (P2_R1179_U379, P2_R1179_U29, P2_U3066);
  not ginst13950 (P2_R1179_U38, P2_U3387);
  nand ginst13951 (P2_R1179_U380, P2_R1179_U240, P2_R1179_U49);
  nand ginst13952 (P2_R1179_U381, P2_R1179_U159, P2_R1179_U232);
  nand ginst13953 (P2_R1179_U382, P2_R1179_U43, P2_U3401);
  nand ginst13954 (P2_R1179_U383, P2_R1179_U31, P2_U3059);
  nand ginst13955 (P2_R1179_U384, P2_R1179_U161, P2_R1179_U241);
  nand ginst13956 (P2_R1179_U385, P2_R1179_U160, P2_R1179_U345);
  nand ginst13957 (P2_R1179_U386, P2_R1179_U36, P2_U3398);
  nand ginst13958 (P2_R1179_U387, P2_R1179_U40, P2_U3063);
  nand ginst13959 (P2_R1179_U388, P2_R1179_U36, P2_U3398);
  nand ginst13960 (P2_R1179_U389, P2_R1179_U40, P2_U3063);
  not ginst13961 (P2_R1179_U39, P2_U3077);
  nand ginst13962 (P2_R1179_U390, P2_R1179_U388, P2_R1179_U389);
  nand ginst13963 (P2_R1179_U391, P2_R1179_U34, P2_U3395);
  nand ginst13964 (P2_R1179_U392, P2_R1179_U37, P2_U3067);
  nand ginst13965 (P2_R1179_U393, P2_R1179_U243, P2_R1179_U50);
  nand ginst13966 (P2_R1179_U394, P2_R1179_U162, P2_R1179_U205);
  nand ginst13967 (P2_R1179_U395, P2_R1179_U164, P2_U3904);
  nand ginst13968 (P2_R1179_U396, P2_R1179_U163, P2_U3054);
  nand ginst13969 (P2_R1179_U397, P2_R1179_U395, P2_R1179_U396);
  nand ginst13970 (P2_R1179_U398, P2_R1179_U164, P2_U3904);
  nand ginst13971 (P2_R1179_U399, P2_R1179_U163, P2_U3054);
  not ginst13972 (P2_R1179_U40, P2_U3398);
  nand ginst13973 (P2_R1179_U400, P2_R1179_U397, P2_R1179_U51, P2_U3053);
  nand ginst13974 (P2_R1179_U401, P2_R1179_U16, P2_R1179_U92, P2_U3895);
  nand ginst13975 (P2_R1179_U402, P2_R1179_U92, P2_U3895);
  nand ginst13976 (P2_R1179_U403, P2_R1179_U51, P2_U3053);
  not ginst13977 (P2_R1179_U404, P2_R1179_U138);
  nand ginst13978 (P2_R1179_U405, P2_R1179_U361, P2_R1179_U404);
  nand ginst13979 (P2_R1179_U406, P2_R1179_U138, P2_R1179_U166);
  nand ginst13980 (P2_R1179_U407, P2_R1179_U54, P2_U3896);
  nand ginst13981 (P2_R1179_U408, P2_R1179_U91, P2_U3052);
  nand ginst13982 (P2_R1179_U409, P2_R1179_U54, P2_U3896);
  not ginst13983 (P2_R1179_U41, P2_U3070);
  nand ginst13984 (P2_R1179_U410, P2_R1179_U91, P2_U3052);
  nand ginst13985 (P2_R1179_U411, P2_R1179_U409, P2_R1179_U410);
  nand ginst13986 (P2_R1179_U412, P2_R1179_U52, P2_U3897);
  nand ginst13987 (P2_R1179_U413, P2_R1179_U90, P2_U3056);
  nand ginst13988 (P2_R1179_U414, P2_R1179_U306, P2_R1179_U93);
  nand ginst13989 (P2_R1179_U415, P2_R1179_U167, P2_R1179_U298);
  nand ginst13990 (P2_R1179_U416, P2_R1179_U89, P2_U3898);
  nand ginst13991 (P2_R1179_U417, P2_R1179_U88, P2_U3057);
  not ginst13992 (P2_R1179_U418, P2_R1179_U141);
  nand ginst13993 (P2_R1179_U419, P2_R1179_U294, P2_R1179_U418);
  not ginst13994 (P2_R1179_U42, P2_U3066);
  nand ginst13995 (P2_R1179_U420, P2_R1179_U141, P2_R1179_U168);
  nand ginst13996 (P2_R1179_U421, P2_R1179_U87, P2_U3899);
  nand ginst13997 (P2_R1179_U422, P2_R1179_U86, P2_U3064);
  not ginst13998 (P2_R1179_U423, P2_R1179_U142);
  nand ginst13999 (P2_R1179_U424, P2_R1179_U290, P2_R1179_U423);
  nand ginst14000 (P2_R1179_U425, P2_R1179_U142, P2_R1179_U169);
  nand ginst14001 (P2_R1179_U426, P2_R1179_U82, P2_U3900);
  nand ginst14002 (P2_R1179_U427, P2_R1179_U79, P2_U3065);
  nand ginst14003 (P2_R1179_U428, P2_R1179_U426, P2_R1179_U427);
  nand ginst14004 (P2_R1179_U429, P2_R1179_U83, P2_U3901);
  not ginst14005 (P2_R1179_U43, P2_U3059);
  nand ginst14006 (P2_R1179_U430, P2_R1179_U80, P2_U3060);
  nand ginst14007 (P2_R1179_U431, P2_R1179_U316, P2_R1179_U94);
  nand ginst14008 (P2_R1179_U432, P2_R1179_U170, P2_R1179_U308);
  nand ginst14009 (P2_R1179_U433, P2_R1179_U84, P2_U3902);
  nand ginst14010 (P2_R1179_U434, P2_R1179_U81, P2_U3074);
  nand ginst14011 (P2_R1179_U435, P2_R1179_U172, P2_R1179_U317);
  nand ginst14012 (P2_R1179_U436, P2_R1179_U171, P2_R1179_U280);
  nand ginst14013 (P2_R1179_U437, P2_R1179_U78, P2_U3903);
  nand ginst14014 (P2_R1179_U438, P2_R1179_U77, P2_U3075);
  not ginst14015 (P2_R1179_U439, P2_R1179_U145);
  nand ginst14016 (P2_R1179_U44, P2_R1179_U31, P2_U3059);
  nand ginst14017 (P2_R1179_U440, P2_R1179_U276, P2_R1179_U439);
  nand ginst14018 (P2_R1179_U441, P2_R1179_U145, P2_R1179_U173);
  nand ginst14019 (P2_R1179_U442, P2_R1179_U39, P2_U3392);
  nand ginst14020 (P2_R1179_U443, P2_R1179_U174, P2_U3077);
  not ginst14021 (P2_R1179_U444, P2_R1179_U146);
  nand ginst14022 (P2_R1179_U445, P2_R1179_U203, P2_R1179_U444);
  nand ginst14023 (P2_R1179_U446, P2_R1179_U146, P2_R1179_U175);
  nand ginst14024 (P2_R1179_U447, P2_R1179_U76, P2_U3445);
  nand ginst14025 (P2_R1179_U448, P2_R1179_U75, P2_U3080);
  not ginst14026 (P2_R1179_U449, P2_R1179_U147);
  nand ginst14027 (P2_R1179_U45, P2_R1179_U214, P2_R1179_U216);
  nand ginst14028 (P2_R1179_U450, P2_R1179_U272, P2_R1179_U449);
  nand ginst14029 (P2_R1179_U451, P2_R1179_U147, P2_R1179_U176);
  nand ginst14030 (P2_R1179_U452, P2_R1179_U74, P2_U3443);
  nand ginst14031 (P2_R1179_U453, P2_R1179_U177, P2_U3081);
  not ginst14032 (P2_R1179_U454, P2_R1179_U148);
  nand ginst14033 (P2_R1179_U455, P2_R1179_U270, P2_R1179_U454);
  nand ginst14034 (P2_R1179_U456, P2_R1179_U148, P2_R1179_U178);
  nand ginst14035 (P2_R1179_U457, P2_R1179_U73, P2_U3440);
  nand ginst14036 (P2_R1179_U458, P2_R1179_U72, P2_U3068);
  not ginst14037 (P2_R1179_U459, P2_R1179_U149);
  not ginst14038 (P2_R1179_U46, P2_U3416);
  nand ginst14039 (P2_R1179_U460, P2_R1179_U266, P2_R1179_U459);
  nand ginst14040 (P2_R1179_U461, P2_R1179_U149, P2_R1179_U179);
  nand ginst14041 (P2_R1179_U462, P2_R1179_U68, P2_U3437);
  nand ginst14042 (P2_R1179_U463, P2_R1179_U65, P2_U3072);
  nand ginst14043 (P2_R1179_U464, P2_R1179_U462, P2_R1179_U463);
  nand ginst14044 (P2_R1179_U465, P2_R1179_U69, P2_U3434);
  nand ginst14045 (P2_R1179_U466, P2_R1179_U66, P2_U3073);
  nand ginst14046 (P2_R1179_U467, P2_R1179_U327, P2_R1179_U95);
  nand ginst14047 (P2_R1179_U468, P2_R1179_U180, P2_R1179_U319);
  nand ginst14048 (P2_R1179_U469, P2_R1179_U70, P2_U3431);
  not ginst14049 (P2_R1179_U47, P2_U3082);
  nand ginst14050 (P2_R1179_U470, P2_R1179_U67, P2_U3078);
  nand ginst14051 (P2_R1179_U471, P2_R1179_U182, P2_R1179_U328);
  nand ginst14052 (P2_R1179_U472, P2_R1179_U181, P2_R1179_U256);
  nand ginst14053 (P2_R1179_U473, P2_R1179_U64, P2_U3428);
  nand ginst14054 (P2_R1179_U474, P2_R1179_U63, P2_U3079);
  not ginst14055 (P2_R1179_U475, P2_R1179_U152);
  nand ginst14056 (P2_R1179_U476, P2_R1179_U354, P2_R1179_U475);
  nand ginst14057 (P2_R1179_U477, P2_R1179_U152, P2_R1179_U183);
  nand ginst14058 (P2_R1179_U478, P2_R1179_U55, P2_U3425);
  nand ginst14059 (P2_R1179_U479, P2_R1179_U61, P2_U3071);
  nand ginst14060 (P2_R1179_U48, P2_R1179_U217, P2_R1179_U45);
  not ginst14061 (P2_R1179_U480, P2_R1179_U153);
  nand ginst14062 (P2_R1179_U481, P2_R1179_U352, P2_R1179_U480);
  nand ginst14063 (P2_R1179_U482, P2_R1179_U153, P2_R1179_U184);
  nand ginst14064 (P2_R1179_U483, P2_R1179_U56, P2_U3422);
  nand ginst14065 (P2_R1179_U484, P2_R1179_U60, P2_U3062);
  nand ginst14066 (P2_R1179_U485, P2_R1179_U483, P2_R1179_U484);
  nand ginst14067 (P2_R1179_U486, P2_R1179_U57, P2_U3419);
  nand ginst14068 (P2_R1179_U487, P2_R1179_U58, P2_U3061);
  nand ginst14069 (P2_R1179_U488, P2_R1179_U336, P2_R1179_U96);
  nand ginst14070 (P2_R1179_U489, P2_R1179_U185, P2_R1179_U350);
  nand ginst14071 (P2_R1179_U49, P2_R1179_U231, P2_R1179_U44);
  nand ginst14072 (P2_R1179_U50, P2_R1179_U188, P2_R1179_U204, P2_R1179_U338);
  not ginst14073 (P2_R1179_U51, P2_U3895);
  not ginst14074 (P2_R1179_U52, P2_U3056);
  nand ginst14075 (P2_R1179_U53, P2_R1179_U90, P2_U3056);
  not ginst14076 (P2_R1179_U54, P2_U3052);
  not ginst14077 (P2_R1179_U55, P2_U3071);
  not ginst14078 (P2_R1179_U56, P2_U3062);
  not ginst14079 (P2_R1179_U57, P2_U3061);
  not ginst14080 (P2_R1179_U58, P2_U3419);
  nand ginst14081 (P2_R1179_U59, P2_R1179_U46, P2_U3082);
  and ginst14082 (P2_R1179_U6, P2_R1179_U211, P2_R1179_U212);
  not ginst14083 (P2_R1179_U60, P2_U3422);
  not ginst14084 (P2_R1179_U61, P2_U3425);
  nand ginst14085 (P2_R1179_U62, P2_R1179_U248, P2_R1179_U249);
  not ginst14086 (P2_R1179_U63, P2_U3428);
  not ginst14087 (P2_R1179_U64, P2_U3079);
  not ginst14088 (P2_R1179_U65, P2_U3437);
  not ginst14089 (P2_R1179_U66, P2_U3434);
  not ginst14090 (P2_R1179_U67, P2_U3431);
  not ginst14091 (P2_R1179_U68, P2_U3072);
  not ginst14092 (P2_R1179_U69, P2_U3073);
  and ginst14093 (P2_R1179_U7, P2_R1179_U245, P2_R1179_U246);
  not ginst14094 (P2_R1179_U70, P2_U3078);
  nand ginst14095 (P2_R1179_U71, P2_R1179_U67, P2_U3078);
  not ginst14096 (P2_R1179_U72, P2_U3440);
  not ginst14097 (P2_R1179_U73, P2_U3068);
  not ginst14098 (P2_R1179_U74, P2_U3081);
  not ginst14099 (P2_R1179_U75, P2_U3445);
  not ginst14100 (P2_R1179_U76, P2_U3080);
  not ginst14101 (P2_R1179_U77, P2_U3903);
  not ginst14102 (P2_R1179_U78, P2_U3075);
  not ginst14103 (P2_R1179_U79, P2_U3900);
  and ginst14104 (P2_R1179_U8, P2_R1179_U193, P2_R1179_U257);
  not ginst14105 (P2_R1179_U80, P2_U3901);
  not ginst14106 (P2_R1179_U81, P2_U3902);
  not ginst14107 (P2_R1179_U82, P2_U3065);
  not ginst14108 (P2_R1179_U83, P2_U3060);
  not ginst14109 (P2_R1179_U84, P2_U3074);
  nand ginst14110 (P2_R1179_U85, P2_R1179_U81, P2_U3074);
  not ginst14111 (P2_R1179_U86, P2_U3899);
  not ginst14112 (P2_R1179_U87, P2_U3064);
  not ginst14113 (P2_R1179_U88, P2_U3898);
  not ginst14114 (P2_R1179_U89, P2_U3057);
  and ginst14115 (P2_R1179_U9, P2_R1179_U258, P2_R1179_U259);
  not ginst14116 (P2_R1179_U90, P2_U3897);
  not ginst14117 (P2_R1179_U91, P2_U3896);
  not ginst14118 (P2_R1179_U92, P2_U3053);
  nand ginst14119 (P2_R1179_U93, P2_R1179_U296, P2_R1179_U297);
  nand ginst14120 (P2_R1179_U94, P2_R1179_U307, P2_R1179_U85);
  nand ginst14121 (P2_R1179_U95, P2_R1179_U318, P2_R1179_U71);
  nand ginst14122 (P2_R1179_U96, P2_R1179_U349, P2_R1179_U59);
  not ginst14123 (P2_R1179_U97, P2_U3076);
  nand ginst14124 (P2_R1179_U98, P2_R1179_U405, P2_R1179_U406);
  nand ginst14125 (P2_R1179_U99, P2_R1179_U419, P2_R1179_U420);
  and ginst14126 (P2_R1200_U10, P2_R1200_U194, P2_R1200_U281);
  nand ginst14127 (P2_R1200_U100, P2_R1200_U424, P2_R1200_U425);
  nand ginst14128 (P2_R1200_U101, P2_R1200_U440, P2_R1200_U441);
  nand ginst14129 (P2_R1200_U102, P2_R1200_U445, P2_R1200_U446);
  nand ginst14130 (P2_R1200_U103, P2_R1200_U450, P2_R1200_U451);
  nand ginst14131 (P2_R1200_U104, P2_R1200_U455, P2_R1200_U456);
  nand ginst14132 (P2_R1200_U105, P2_R1200_U460, P2_R1200_U461);
  nand ginst14133 (P2_R1200_U106, P2_R1200_U476, P2_R1200_U477);
  nand ginst14134 (P2_R1200_U107, P2_R1200_U481, P2_R1200_U482);
  nand ginst14135 (P2_R1200_U108, P2_R1200_U364, P2_R1200_U365);
  nand ginst14136 (P2_R1200_U109, P2_R1200_U373, P2_R1200_U374);
  and ginst14137 (P2_R1200_U11, P2_R1200_U282, P2_R1200_U283);
  nand ginst14138 (P2_R1200_U110, P2_R1200_U380, P2_R1200_U381);
  nand ginst14139 (P2_R1200_U111, P2_R1200_U384, P2_R1200_U385);
  nand ginst14140 (P2_R1200_U112, P2_R1200_U393, P2_R1200_U394);
  nand ginst14141 (P2_R1200_U113, P2_R1200_U414, P2_R1200_U415);
  nand ginst14142 (P2_R1200_U114, P2_R1200_U431, P2_R1200_U432);
  nand ginst14143 (P2_R1200_U115, P2_R1200_U435, P2_R1200_U436);
  nand ginst14144 (P2_R1200_U116, P2_R1200_U467, P2_R1200_U468);
  nand ginst14145 (P2_R1200_U117, P2_R1200_U471, P2_R1200_U472);
  nand ginst14146 (P2_R1200_U118, P2_R1200_U488, P2_R1200_U489);
  and ginst14147 (P2_R1200_U119, P2_R1200_U196, P2_R1200_U206);
  and ginst14148 (P2_R1200_U12, P2_R1200_U195, P2_R1200_U299);
  and ginst14149 (P2_R1200_U120, P2_R1200_U208, P2_R1200_U209);
  and ginst14150 (P2_R1200_U121, P2_R1200_U13, P2_R1200_U14);
  and ginst14151 (P2_R1200_U122, P2_R1200_U222, P2_R1200_U340);
  and ginst14152 (P2_R1200_U123, P2_R1200_U122, P2_R1200_U342);
  and ginst14153 (P2_R1200_U124, P2_R1200_U27, P2_R1200_U366, P2_R1200_U367);
  and ginst14154 (P2_R1200_U125, P2_R1200_U198, P2_R1200_U370);
  and ginst14155 (P2_R1200_U126, P2_R1200_U237, P2_R1200_U6);
  and ginst14156 (P2_R1200_U127, P2_R1200_U197, P2_R1200_U377);
  and ginst14157 (P2_R1200_U128, P2_R1200_U35, P2_R1200_U386, P2_R1200_U387);
  and ginst14158 (P2_R1200_U129, P2_R1200_U196, P2_R1200_U390);
  and ginst14159 (P2_R1200_U13, P2_R1200_U197, P2_R1200_U210, P2_R1200_U215);
  and ginst14160 (P2_R1200_U130, P2_R1200_U15, P2_R1200_U251);
  and ginst14161 (P2_R1200_U131, P2_R1200_U252, P2_R1200_U343);
  and ginst14162 (P2_R1200_U132, P2_R1200_U262, P2_R1200_U8);
  and ginst14163 (P2_R1200_U133, P2_R1200_U10, P2_R1200_U286);
  and ginst14164 (P2_R1200_U134, P2_R1200_U301, P2_R1200_U302);
  and ginst14165 (P2_R1200_U135, P2_R1200_U303, P2_R1200_U397);
  and ginst14166 (P2_R1200_U136, P2_R1200_U16, P2_R1200_U301, P2_R1200_U302, P2_R1200_U304);
  and ginst14167 (P2_R1200_U137, P2_R1200_U165, P2_R1200_U359);
  nand ginst14168 (P2_R1200_U138, P2_R1200_U402, P2_R1200_U403);
  and ginst14169 (P2_R1200_U139, P2_R1200_U407, P2_R1200_U408, P2_R1200_U53);
  and ginst14170 (P2_R1200_U14, P2_R1200_U198, P2_R1200_U220);
  and ginst14171 (P2_R1200_U140, P2_R1200_U195, P2_R1200_U411);
  nand ginst14172 (P2_R1200_U141, P2_R1200_U416, P2_R1200_U417);
  nand ginst14173 (P2_R1200_U142, P2_R1200_U421, P2_R1200_U422);
  and ginst14174 (P2_R1200_U143, P2_R1200_U11, P2_R1200_U313);
  and ginst14175 (P2_R1200_U144, P2_R1200_U194, P2_R1200_U428);
  nand ginst14176 (P2_R1200_U145, P2_R1200_U437, P2_R1200_U438);
  nand ginst14177 (P2_R1200_U146, P2_R1200_U442, P2_R1200_U443);
  nand ginst14178 (P2_R1200_U147, P2_R1200_U447, P2_R1200_U448);
  nand ginst14179 (P2_R1200_U148, P2_R1200_U452, P2_R1200_U453);
  nand ginst14180 (P2_R1200_U149, P2_R1200_U457, P2_R1200_U458);
  and ginst14181 (P2_R1200_U15, P2_R1200_U192, P2_R1200_U224, P2_R1200_U244);
  and ginst14182 (P2_R1200_U150, P2_R1200_U324, P2_R1200_U9);
  and ginst14183 (P2_R1200_U151, P2_R1200_U193, P2_R1200_U464);
  nand ginst14184 (P2_R1200_U152, P2_R1200_U473, P2_R1200_U474);
  nand ginst14185 (P2_R1200_U153, P2_R1200_U478, P2_R1200_U479);
  and ginst14186 (P2_R1200_U154, P2_R1200_U333, P2_R1200_U7);
  and ginst14187 (P2_R1200_U155, P2_R1200_U192, P2_R1200_U485);
  and ginst14188 (P2_R1200_U156, P2_R1200_U362, P2_R1200_U363);
  nand ginst14189 (P2_R1200_U157, P2_R1200_U123, P2_R1200_U341);
  and ginst14190 (P2_R1200_U158, P2_R1200_U371, P2_R1200_U372);
  and ginst14191 (P2_R1200_U159, P2_R1200_U378, P2_R1200_U379);
  and ginst14192 (P2_R1200_U16, P2_R1200_U398, P2_R1200_U399);
  and ginst14193 (P2_R1200_U160, P2_R1200_U382, P2_R1200_U383);
  nand ginst14194 (P2_R1200_U161, P2_R1200_U120, P2_R1200_U344);
  and ginst14195 (P2_R1200_U162, P2_R1200_U391, P2_R1200_U392);
  not ginst14196 (P2_R1200_U163, P2_U3904);
  not ginst14197 (P2_R1200_U164, P2_U3054);
  and ginst14198 (P2_R1200_U165, P2_R1200_U400, P2_R1200_U401);
  nand ginst14199 (P2_R1200_U166, P2_R1200_U134, P2_R1200_U360);
  and ginst14200 (P2_R1200_U167, P2_R1200_U412, P2_R1200_U413);
  nand ginst14201 (P2_R1200_U168, P2_R1200_U292, P2_R1200_U293);
  nand ginst14202 (P2_R1200_U169, P2_R1200_U288, P2_R1200_U289);
  nand ginst14203 (P2_R1200_U17, P2_R1200_U331, P2_R1200_U334);
  and ginst14204 (P2_R1200_U170, P2_R1200_U429, P2_R1200_U430);
  and ginst14205 (P2_R1200_U171, P2_R1200_U433, P2_R1200_U434);
  nand ginst14206 (P2_R1200_U172, P2_R1200_U278, P2_R1200_U279);
  nand ginst14207 (P2_R1200_U173, P2_R1200_U274, P2_R1200_U275);
  not ginst14208 (P2_R1200_U174, P2_U3392);
  nand ginst14209 (P2_R1200_U175, P2_R1200_U97, P2_U3387);
  nand ginst14210 (P2_R1200_U176, P2_R1200_U187, P2_R1200_U271, P2_R1200_U339);
  not ginst14211 (P2_R1200_U177, P2_U3443);
  nand ginst14212 (P2_R1200_U178, P2_R1200_U268, P2_R1200_U269);
  nand ginst14213 (P2_R1200_U179, P2_R1200_U264, P2_R1200_U265);
  nand ginst14214 (P2_R1200_U18, P2_R1200_U322, P2_R1200_U325);
  and ginst14215 (P2_R1200_U180, P2_R1200_U465, P2_R1200_U466);
  and ginst14216 (P2_R1200_U181, P2_R1200_U469, P2_R1200_U470);
  nand ginst14217 (P2_R1200_U182, P2_R1200_U254, P2_R1200_U255);
  nand ginst14218 (P2_R1200_U183, P2_R1200_U131, P2_R1200_U353);
  nand ginst14219 (P2_R1200_U184, P2_R1200_U351, P2_R1200_U62);
  and ginst14220 (P2_R1200_U185, P2_R1200_U486, P2_R1200_U487);
  nand ginst14221 (P2_R1200_U186, P2_R1200_U135, P2_R1200_U166);
  nand ginst14222 (P2_R1200_U187, P2_R1200_U177, P2_R1200_U178);
  nand ginst14223 (P2_R1200_U188, P2_R1200_U174, P2_R1200_U175);
  not ginst14224 (P2_R1200_U189, P2_R1200_U53);
  nand ginst14225 (P2_R1200_U19, P2_R1200_U311, P2_R1200_U314);
  not ginst14226 (P2_R1200_U190, P2_R1200_U35);
  not ginst14227 (P2_R1200_U191, P2_R1200_U27);
  nand ginst14228 (P2_R1200_U192, P2_R1200_U57, P2_U3419);
  nand ginst14229 (P2_R1200_U193, P2_R1200_U69, P2_U3434);
  nand ginst14230 (P2_R1200_U194, P2_R1200_U83, P2_U3901);
  nand ginst14231 (P2_R1200_U195, P2_R1200_U52, P2_U3897);
  nand ginst14232 (P2_R1200_U196, P2_R1200_U34, P2_U3395);
  nand ginst14233 (P2_R1200_U197, P2_R1200_U42, P2_U3404);
  nand ginst14234 (P2_R1200_U198, P2_R1200_U26, P2_U3410);
  not ginst14235 (P2_R1200_U199, P2_R1200_U71);
  nand ginst14236 (P2_R1200_U20, P2_R1200_U305, P2_R1200_U357);
  not ginst14237 (P2_R1200_U200, P2_R1200_U85);
  not ginst14238 (P2_R1200_U201, P2_R1200_U44);
  not ginst14239 (P2_R1200_U202, P2_R1200_U59);
  not ginst14240 (P2_R1200_U203, P2_R1200_U175);
  nand ginst14241 (P2_R1200_U204, P2_R1200_U175, P2_U3077);
  not ginst14242 (P2_R1200_U205, P2_R1200_U50);
  nand ginst14243 (P2_R1200_U206, P2_R1200_U36, P2_U3398);
  nand ginst14244 (P2_R1200_U207, P2_R1200_U35, P2_R1200_U36);
  nand ginst14245 (P2_R1200_U208, P2_R1200_U207, P2_R1200_U40);
  nand ginst14246 (P2_R1200_U209, P2_R1200_U190, P2_U3063);
  nand ginst14247 (P2_R1200_U21, P2_R1200_U137, P2_R1200_U186);
  nand ginst14248 (P2_R1200_U210, P2_R1200_U41, P2_U3407);
  nand ginst14249 (P2_R1200_U211, P2_R1200_U30, P2_U3070);
  nand ginst14250 (P2_R1200_U212, P2_R1200_U29, P2_U3066);
  nand ginst14251 (P2_R1200_U213, P2_R1200_U197, P2_R1200_U201);
  nand ginst14252 (P2_R1200_U214, P2_R1200_U213, P2_R1200_U6);
  nand ginst14253 (P2_R1200_U215, P2_R1200_U43, P2_U3401);
  nand ginst14254 (P2_R1200_U216, P2_R1200_U41, P2_U3407);
  nand ginst14255 (P2_R1200_U217, P2_R1200_U13, P2_R1200_U161);
  not ginst14256 (P2_R1200_U218, P2_R1200_U45);
  not ginst14257 (P2_R1200_U219, P2_R1200_U48);
  nand ginst14258 (P2_R1200_U22, P2_R1200_U242, P2_R1200_U347);
  nand ginst14259 (P2_R1200_U220, P2_R1200_U28, P2_U3413);
  nand ginst14260 (P2_R1200_U221, P2_R1200_U27, P2_R1200_U28);
  nand ginst14261 (P2_R1200_U222, P2_R1200_U191, P2_U3083);
  not ginst14262 (P2_R1200_U223, P2_R1200_U157);
  nand ginst14263 (P2_R1200_U224, P2_R1200_U47, P2_U3416);
  nand ginst14264 (P2_R1200_U225, P2_R1200_U224, P2_R1200_U59);
  nand ginst14265 (P2_R1200_U226, P2_R1200_U219, P2_R1200_U27);
  nand ginst14266 (P2_R1200_U227, P2_R1200_U125, P2_R1200_U226);
  nand ginst14267 (P2_R1200_U228, P2_R1200_U198, P2_R1200_U48);
  nand ginst14268 (P2_R1200_U229, P2_R1200_U124, P2_R1200_U228);
  nand ginst14269 (P2_R1200_U23, P2_R1200_U235, P2_R1200_U238);
  nand ginst14270 (P2_R1200_U230, P2_R1200_U198, P2_R1200_U27);
  nand ginst14271 (P2_R1200_U231, P2_R1200_U161, P2_R1200_U215);
  not ginst14272 (P2_R1200_U232, P2_R1200_U49);
  nand ginst14273 (P2_R1200_U233, P2_R1200_U29, P2_U3066);
  nand ginst14274 (P2_R1200_U234, P2_R1200_U232, P2_R1200_U233);
  nand ginst14275 (P2_R1200_U235, P2_R1200_U127, P2_R1200_U234);
  nand ginst14276 (P2_R1200_U236, P2_R1200_U197, P2_R1200_U49);
  nand ginst14277 (P2_R1200_U237, P2_R1200_U41, P2_U3407);
  nand ginst14278 (P2_R1200_U238, P2_R1200_U126, P2_R1200_U236);
  nand ginst14279 (P2_R1200_U239, P2_R1200_U29, P2_U3066);
  nand ginst14280 (P2_R1200_U24, P2_R1200_U227, P2_R1200_U229);
  nand ginst14281 (P2_R1200_U240, P2_R1200_U197, P2_R1200_U239);
  nand ginst14282 (P2_R1200_U241, P2_R1200_U215, P2_R1200_U44);
  nand ginst14283 (P2_R1200_U242, P2_R1200_U129, P2_R1200_U348);
  nand ginst14284 (P2_R1200_U243, P2_R1200_U196, P2_R1200_U35);
  nand ginst14285 (P2_R1200_U244, P2_R1200_U56, P2_U3422);
  nand ginst14286 (P2_R1200_U245, P2_R1200_U60, P2_U3062);
  nand ginst14287 (P2_R1200_U246, P2_R1200_U58, P2_U3061);
  nand ginst14288 (P2_R1200_U247, P2_R1200_U192, P2_R1200_U202);
  nand ginst14289 (P2_R1200_U248, P2_R1200_U247, P2_R1200_U7);
  nand ginst14290 (P2_R1200_U249, P2_R1200_U56, P2_U3422);
  nand ginst14291 (P2_R1200_U25, P2_R1200_U175, P2_R1200_U337);
  not ginst14292 (P2_R1200_U250, P2_R1200_U62);
  nand ginst14293 (P2_R1200_U251, P2_R1200_U55, P2_U3425);
  nand ginst14294 (P2_R1200_U252, P2_R1200_U61, P2_U3071);
  nand ginst14295 (P2_R1200_U253, P2_R1200_U64, P2_U3428);
  nand ginst14296 (P2_R1200_U254, P2_R1200_U183, P2_R1200_U253);
  nand ginst14297 (P2_R1200_U255, P2_R1200_U63, P2_U3079);
  not ginst14298 (P2_R1200_U256, P2_R1200_U182);
  nand ginst14299 (P2_R1200_U257, P2_R1200_U68, P2_U3437);
  nand ginst14300 (P2_R1200_U258, P2_R1200_U65, P2_U3072);
  nand ginst14301 (P2_R1200_U259, P2_R1200_U66, P2_U3073);
  not ginst14302 (P2_R1200_U26, P2_U3069);
  nand ginst14303 (P2_R1200_U260, P2_R1200_U199, P2_R1200_U8);
  nand ginst14304 (P2_R1200_U261, P2_R1200_U260, P2_R1200_U9);
  nand ginst14305 (P2_R1200_U262, P2_R1200_U70, P2_U3431);
  nand ginst14306 (P2_R1200_U263, P2_R1200_U68, P2_U3437);
  nand ginst14307 (P2_R1200_U264, P2_R1200_U132, P2_R1200_U182);
  nand ginst14308 (P2_R1200_U265, P2_R1200_U261, P2_R1200_U263);
  not ginst14309 (P2_R1200_U266, P2_R1200_U179);
  nand ginst14310 (P2_R1200_U267, P2_R1200_U73, P2_U3440);
  nand ginst14311 (P2_R1200_U268, P2_R1200_U179, P2_R1200_U267);
  nand ginst14312 (P2_R1200_U269, P2_R1200_U72, P2_U3068);
  nand ginst14313 (P2_R1200_U27, P2_R1200_U32, P2_U3069);
  not ginst14314 (P2_R1200_U270, P2_R1200_U178);
  nand ginst14315 (P2_R1200_U271, P2_R1200_U178, P2_U3081);
  not ginst14316 (P2_R1200_U272, P2_R1200_U176);
  nand ginst14317 (P2_R1200_U273, P2_R1200_U76, P2_U3445);
  nand ginst14318 (P2_R1200_U274, P2_R1200_U176, P2_R1200_U273);
  nand ginst14319 (P2_R1200_U275, P2_R1200_U75, P2_U3080);
  not ginst14320 (P2_R1200_U276, P2_R1200_U173);
  nand ginst14321 (P2_R1200_U277, P2_R1200_U78, P2_U3903);
  nand ginst14322 (P2_R1200_U278, P2_R1200_U173, P2_R1200_U277);
  nand ginst14323 (P2_R1200_U279, P2_R1200_U77, P2_U3075);
  not ginst14324 (P2_R1200_U28, P2_U3083);
  not ginst14325 (P2_R1200_U280, P2_R1200_U172);
  nand ginst14326 (P2_R1200_U281, P2_R1200_U82, P2_U3900);
  nand ginst14327 (P2_R1200_U282, P2_R1200_U79, P2_U3065);
  nand ginst14328 (P2_R1200_U283, P2_R1200_U80, P2_U3060);
  nand ginst14329 (P2_R1200_U284, P2_R1200_U10, P2_R1200_U200);
  nand ginst14330 (P2_R1200_U285, P2_R1200_U11, P2_R1200_U284);
  nand ginst14331 (P2_R1200_U286, P2_R1200_U84, P2_U3902);
  nand ginst14332 (P2_R1200_U287, P2_R1200_U82, P2_U3900);
  nand ginst14333 (P2_R1200_U288, P2_R1200_U133, P2_R1200_U172);
  nand ginst14334 (P2_R1200_U289, P2_R1200_U285, P2_R1200_U287);
  not ginst14335 (P2_R1200_U29, P2_U3404);
  not ginst14336 (P2_R1200_U290, P2_R1200_U169);
  nand ginst14337 (P2_R1200_U291, P2_R1200_U87, P2_U3899);
  nand ginst14338 (P2_R1200_U292, P2_R1200_U169, P2_R1200_U291);
  nand ginst14339 (P2_R1200_U293, P2_R1200_U86, P2_U3064);
  not ginst14340 (P2_R1200_U294, P2_R1200_U168);
  nand ginst14341 (P2_R1200_U295, P2_R1200_U89, P2_U3898);
  nand ginst14342 (P2_R1200_U296, P2_R1200_U168, P2_R1200_U295);
  nand ginst14343 (P2_R1200_U297, P2_R1200_U88, P2_U3057);
  not ginst14344 (P2_R1200_U298, P2_R1200_U93);
  nand ginst14345 (P2_R1200_U299, P2_R1200_U54, P2_U3896);
  not ginst14346 (P2_R1200_U30, P2_U3407);
  nand ginst14347 (P2_R1200_U300, P2_R1200_U53, P2_R1200_U54);
  nand ginst14348 (P2_R1200_U301, P2_R1200_U300, P2_R1200_U91);
  nand ginst14349 (P2_R1200_U302, P2_R1200_U189, P2_U3052);
  nand ginst14350 (P2_R1200_U303, P2_R1200_U92, P2_U3895);
  nand ginst14351 (P2_R1200_U304, P2_R1200_U51, P2_U3053);
  nand ginst14352 (P2_R1200_U305, P2_R1200_U140, P2_R1200_U355);
  nand ginst14353 (P2_R1200_U306, P2_R1200_U195, P2_R1200_U53);
  nand ginst14354 (P2_R1200_U307, P2_R1200_U172, P2_R1200_U286);
  not ginst14355 (P2_R1200_U308, P2_R1200_U94);
  nand ginst14356 (P2_R1200_U309, P2_R1200_U80, P2_U3060);
  not ginst14357 (P2_R1200_U31, P2_U3401);
  nand ginst14358 (P2_R1200_U310, P2_R1200_U308, P2_R1200_U309);
  nand ginst14359 (P2_R1200_U311, P2_R1200_U144, P2_R1200_U310);
  nand ginst14360 (P2_R1200_U312, P2_R1200_U194, P2_R1200_U94);
  nand ginst14361 (P2_R1200_U313, P2_R1200_U82, P2_U3900);
  nand ginst14362 (P2_R1200_U314, P2_R1200_U143, P2_R1200_U312);
  nand ginst14363 (P2_R1200_U315, P2_R1200_U80, P2_U3060);
  nand ginst14364 (P2_R1200_U316, P2_R1200_U194, P2_R1200_U315);
  nand ginst14365 (P2_R1200_U317, P2_R1200_U286, P2_R1200_U85);
  nand ginst14366 (P2_R1200_U318, P2_R1200_U182, P2_R1200_U262);
  not ginst14367 (P2_R1200_U319, P2_R1200_U95);
  not ginst14368 (P2_R1200_U32, P2_U3410);
  nand ginst14369 (P2_R1200_U320, P2_R1200_U66, P2_U3073);
  nand ginst14370 (P2_R1200_U321, P2_R1200_U319, P2_R1200_U320);
  nand ginst14371 (P2_R1200_U322, P2_R1200_U151, P2_R1200_U321);
  nand ginst14372 (P2_R1200_U323, P2_R1200_U193, P2_R1200_U95);
  nand ginst14373 (P2_R1200_U324, P2_R1200_U68, P2_U3437);
  nand ginst14374 (P2_R1200_U325, P2_R1200_U150, P2_R1200_U323);
  nand ginst14375 (P2_R1200_U326, P2_R1200_U66, P2_U3073);
  nand ginst14376 (P2_R1200_U327, P2_R1200_U193, P2_R1200_U326);
  nand ginst14377 (P2_R1200_U328, P2_R1200_U262, P2_R1200_U71);
  nand ginst14378 (P2_R1200_U329, P2_R1200_U58, P2_U3061);
  not ginst14379 (P2_R1200_U33, P2_U3413);
  nand ginst14380 (P2_R1200_U330, P2_R1200_U329, P2_R1200_U350);
  nand ginst14381 (P2_R1200_U331, P2_R1200_U155, P2_R1200_U330);
  nand ginst14382 (P2_R1200_U332, P2_R1200_U192, P2_R1200_U96);
  nand ginst14383 (P2_R1200_U333, P2_R1200_U56, P2_U3422);
  nand ginst14384 (P2_R1200_U334, P2_R1200_U154, P2_R1200_U332);
  nand ginst14385 (P2_R1200_U335, P2_R1200_U58, P2_U3061);
  nand ginst14386 (P2_R1200_U336, P2_R1200_U192, P2_R1200_U335);
  nand ginst14387 (P2_R1200_U337, P2_R1200_U38, P2_U3076);
  nand ginst14388 (P2_R1200_U338, P2_R1200_U174, P2_U3077);
  nand ginst14389 (P2_R1200_U339, P2_R1200_U177, P2_U3081);
  not ginst14390 (P2_R1200_U34, P2_U3067);
  nand ginst14391 (P2_R1200_U340, P2_R1200_U221, P2_R1200_U33);
  nand ginst14392 (P2_R1200_U341, P2_R1200_U121, P2_R1200_U161);
  nand ginst14393 (P2_R1200_U342, P2_R1200_U14, P2_R1200_U218);
  nand ginst14394 (P2_R1200_U343, P2_R1200_U250, P2_R1200_U251);
  nand ginst14395 (P2_R1200_U344, P2_R1200_U119, P2_R1200_U50);
  not ginst14396 (P2_R1200_U345, P2_R1200_U161);
  nand ginst14397 (P2_R1200_U346, P2_R1200_U196, P2_R1200_U50);
  nand ginst14398 (P2_R1200_U347, P2_R1200_U128, P2_R1200_U346);
  nand ginst14399 (P2_R1200_U348, P2_R1200_U205, P2_R1200_U35);
  nand ginst14400 (P2_R1200_U349, P2_R1200_U157, P2_R1200_U224);
  nand ginst14401 (P2_R1200_U35, P2_R1200_U37, P2_U3067);
  not ginst14402 (P2_R1200_U350, P2_R1200_U96);
  nand ginst14403 (P2_R1200_U351, P2_R1200_U15, P2_R1200_U157);
  not ginst14404 (P2_R1200_U352, P2_R1200_U184);
  nand ginst14405 (P2_R1200_U353, P2_R1200_U130, P2_R1200_U157);
  not ginst14406 (P2_R1200_U354, P2_R1200_U183);
  nand ginst14407 (P2_R1200_U355, P2_R1200_U298, P2_R1200_U53);
  nand ginst14408 (P2_R1200_U356, P2_R1200_U195, P2_R1200_U93);
  nand ginst14409 (P2_R1200_U357, P2_R1200_U139, P2_R1200_U356);
  nand ginst14410 (P2_R1200_U358, P2_R1200_U12, P2_R1200_U93);
  nand ginst14411 (P2_R1200_U359, P2_R1200_U136, P2_R1200_U358);
  not ginst14412 (P2_R1200_U36, P2_U3063);
  nand ginst14413 (P2_R1200_U360, P2_R1200_U12, P2_R1200_U93);
  not ginst14414 (P2_R1200_U361, P2_R1200_U166);
  nand ginst14415 (P2_R1200_U362, P2_R1200_U47, P2_U3416);
  nand ginst14416 (P2_R1200_U363, P2_R1200_U46, P2_U3082);
  nand ginst14417 (P2_R1200_U364, P2_R1200_U157, P2_R1200_U225);
  nand ginst14418 (P2_R1200_U365, P2_R1200_U156, P2_R1200_U223);
  nand ginst14419 (P2_R1200_U366, P2_R1200_U28, P2_U3413);
  nand ginst14420 (P2_R1200_U367, P2_R1200_U33, P2_U3083);
  nand ginst14421 (P2_R1200_U368, P2_R1200_U28, P2_U3413);
  nand ginst14422 (P2_R1200_U369, P2_R1200_U33, P2_U3083);
  not ginst14423 (P2_R1200_U37, P2_U3395);
  nand ginst14424 (P2_R1200_U370, P2_R1200_U368, P2_R1200_U369);
  nand ginst14425 (P2_R1200_U371, P2_R1200_U26, P2_U3410);
  nand ginst14426 (P2_R1200_U372, P2_R1200_U32, P2_U3069);
  nand ginst14427 (P2_R1200_U373, P2_R1200_U230, P2_R1200_U48);
  nand ginst14428 (P2_R1200_U374, P2_R1200_U158, P2_R1200_U219);
  nand ginst14429 (P2_R1200_U375, P2_R1200_U41, P2_U3407);
  nand ginst14430 (P2_R1200_U376, P2_R1200_U30, P2_U3070);
  nand ginst14431 (P2_R1200_U377, P2_R1200_U375, P2_R1200_U376);
  nand ginst14432 (P2_R1200_U378, P2_R1200_U42, P2_U3404);
  nand ginst14433 (P2_R1200_U379, P2_R1200_U29, P2_U3066);
  not ginst14434 (P2_R1200_U38, P2_U3387);
  nand ginst14435 (P2_R1200_U380, P2_R1200_U240, P2_R1200_U49);
  nand ginst14436 (P2_R1200_U381, P2_R1200_U159, P2_R1200_U232);
  nand ginst14437 (P2_R1200_U382, P2_R1200_U43, P2_U3401);
  nand ginst14438 (P2_R1200_U383, P2_R1200_U31, P2_U3059);
  nand ginst14439 (P2_R1200_U384, P2_R1200_U161, P2_R1200_U241);
  nand ginst14440 (P2_R1200_U385, P2_R1200_U160, P2_R1200_U345);
  nand ginst14441 (P2_R1200_U386, P2_R1200_U36, P2_U3398);
  nand ginst14442 (P2_R1200_U387, P2_R1200_U40, P2_U3063);
  nand ginst14443 (P2_R1200_U388, P2_R1200_U36, P2_U3398);
  nand ginst14444 (P2_R1200_U389, P2_R1200_U40, P2_U3063);
  not ginst14445 (P2_R1200_U39, P2_U3077);
  nand ginst14446 (P2_R1200_U390, P2_R1200_U388, P2_R1200_U389);
  nand ginst14447 (P2_R1200_U391, P2_R1200_U34, P2_U3395);
  nand ginst14448 (P2_R1200_U392, P2_R1200_U37, P2_U3067);
  nand ginst14449 (P2_R1200_U393, P2_R1200_U243, P2_R1200_U50);
  nand ginst14450 (P2_R1200_U394, P2_R1200_U162, P2_R1200_U205);
  nand ginst14451 (P2_R1200_U395, P2_R1200_U164, P2_U3904);
  nand ginst14452 (P2_R1200_U396, P2_R1200_U163, P2_U3054);
  nand ginst14453 (P2_R1200_U397, P2_R1200_U395, P2_R1200_U396);
  nand ginst14454 (P2_R1200_U398, P2_R1200_U164, P2_U3904);
  nand ginst14455 (P2_R1200_U399, P2_R1200_U163, P2_U3054);
  not ginst14456 (P2_R1200_U40, P2_U3398);
  nand ginst14457 (P2_R1200_U400, P2_R1200_U397, P2_R1200_U51, P2_U3053);
  nand ginst14458 (P2_R1200_U401, P2_R1200_U16, P2_R1200_U92, P2_U3895);
  nand ginst14459 (P2_R1200_U402, P2_R1200_U92, P2_U3895);
  nand ginst14460 (P2_R1200_U403, P2_R1200_U51, P2_U3053);
  not ginst14461 (P2_R1200_U404, P2_R1200_U138);
  nand ginst14462 (P2_R1200_U405, P2_R1200_U361, P2_R1200_U404);
  nand ginst14463 (P2_R1200_U406, P2_R1200_U138, P2_R1200_U166);
  nand ginst14464 (P2_R1200_U407, P2_R1200_U54, P2_U3896);
  nand ginst14465 (P2_R1200_U408, P2_R1200_U91, P2_U3052);
  nand ginst14466 (P2_R1200_U409, P2_R1200_U54, P2_U3896);
  not ginst14467 (P2_R1200_U41, P2_U3070);
  nand ginst14468 (P2_R1200_U410, P2_R1200_U91, P2_U3052);
  nand ginst14469 (P2_R1200_U411, P2_R1200_U409, P2_R1200_U410);
  nand ginst14470 (P2_R1200_U412, P2_R1200_U52, P2_U3897);
  nand ginst14471 (P2_R1200_U413, P2_R1200_U90, P2_U3056);
  nand ginst14472 (P2_R1200_U414, P2_R1200_U306, P2_R1200_U93);
  nand ginst14473 (P2_R1200_U415, P2_R1200_U167, P2_R1200_U298);
  nand ginst14474 (P2_R1200_U416, P2_R1200_U89, P2_U3898);
  nand ginst14475 (P2_R1200_U417, P2_R1200_U88, P2_U3057);
  not ginst14476 (P2_R1200_U418, P2_R1200_U141);
  nand ginst14477 (P2_R1200_U419, P2_R1200_U294, P2_R1200_U418);
  not ginst14478 (P2_R1200_U42, P2_U3066);
  nand ginst14479 (P2_R1200_U420, P2_R1200_U141, P2_R1200_U168);
  nand ginst14480 (P2_R1200_U421, P2_R1200_U87, P2_U3899);
  nand ginst14481 (P2_R1200_U422, P2_R1200_U86, P2_U3064);
  not ginst14482 (P2_R1200_U423, P2_R1200_U142);
  nand ginst14483 (P2_R1200_U424, P2_R1200_U290, P2_R1200_U423);
  nand ginst14484 (P2_R1200_U425, P2_R1200_U142, P2_R1200_U169);
  nand ginst14485 (P2_R1200_U426, P2_R1200_U82, P2_U3900);
  nand ginst14486 (P2_R1200_U427, P2_R1200_U79, P2_U3065);
  nand ginst14487 (P2_R1200_U428, P2_R1200_U426, P2_R1200_U427);
  nand ginst14488 (P2_R1200_U429, P2_R1200_U83, P2_U3901);
  not ginst14489 (P2_R1200_U43, P2_U3059);
  nand ginst14490 (P2_R1200_U430, P2_R1200_U80, P2_U3060);
  nand ginst14491 (P2_R1200_U431, P2_R1200_U316, P2_R1200_U94);
  nand ginst14492 (P2_R1200_U432, P2_R1200_U170, P2_R1200_U308);
  nand ginst14493 (P2_R1200_U433, P2_R1200_U84, P2_U3902);
  nand ginst14494 (P2_R1200_U434, P2_R1200_U81, P2_U3074);
  nand ginst14495 (P2_R1200_U435, P2_R1200_U172, P2_R1200_U317);
  nand ginst14496 (P2_R1200_U436, P2_R1200_U171, P2_R1200_U280);
  nand ginst14497 (P2_R1200_U437, P2_R1200_U78, P2_U3903);
  nand ginst14498 (P2_R1200_U438, P2_R1200_U77, P2_U3075);
  not ginst14499 (P2_R1200_U439, P2_R1200_U145);
  nand ginst14500 (P2_R1200_U44, P2_R1200_U31, P2_U3059);
  nand ginst14501 (P2_R1200_U440, P2_R1200_U276, P2_R1200_U439);
  nand ginst14502 (P2_R1200_U441, P2_R1200_U145, P2_R1200_U173);
  nand ginst14503 (P2_R1200_U442, P2_R1200_U39, P2_U3392);
  nand ginst14504 (P2_R1200_U443, P2_R1200_U174, P2_U3077);
  not ginst14505 (P2_R1200_U444, P2_R1200_U146);
  nand ginst14506 (P2_R1200_U445, P2_R1200_U203, P2_R1200_U444);
  nand ginst14507 (P2_R1200_U446, P2_R1200_U146, P2_R1200_U175);
  nand ginst14508 (P2_R1200_U447, P2_R1200_U76, P2_U3445);
  nand ginst14509 (P2_R1200_U448, P2_R1200_U75, P2_U3080);
  not ginst14510 (P2_R1200_U449, P2_R1200_U147);
  nand ginst14511 (P2_R1200_U45, P2_R1200_U214, P2_R1200_U216);
  nand ginst14512 (P2_R1200_U450, P2_R1200_U272, P2_R1200_U449);
  nand ginst14513 (P2_R1200_U451, P2_R1200_U147, P2_R1200_U176);
  nand ginst14514 (P2_R1200_U452, P2_R1200_U74, P2_U3443);
  nand ginst14515 (P2_R1200_U453, P2_R1200_U177, P2_U3081);
  not ginst14516 (P2_R1200_U454, P2_R1200_U148);
  nand ginst14517 (P2_R1200_U455, P2_R1200_U270, P2_R1200_U454);
  nand ginst14518 (P2_R1200_U456, P2_R1200_U148, P2_R1200_U178);
  nand ginst14519 (P2_R1200_U457, P2_R1200_U73, P2_U3440);
  nand ginst14520 (P2_R1200_U458, P2_R1200_U72, P2_U3068);
  not ginst14521 (P2_R1200_U459, P2_R1200_U149);
  not ginst14522 (P2_R1200_U46, P2_U3416);
  nand ginst14523 (P2_R1200_U460, P2_R1200_U266, P2_R1200_U459);
  nand ginst14524 (P2_R1200_U461, P2_R1200_U149, P2_R1200_U179);
  nand ginst14525 (P2_R1200_U462, P2_R1200_U68, P2_U3437);
  nand ginst14526 (P2_R1200_U463, P2_R1200_U65, P2_U3072);
  nand ginst14527 (P2_R1200_U464, P2_R1200_U462, P2_R1200_U463);
  nand ginst14528 (P2_R1200_U465, P2_R1200_U69, P2_U3434);
  nand ginst14529 (P2_R1200_U466, P2_R1200_U66, P2_U3073);
  nand ginst14530 (P2_R1200_U467, P2_R1200_U327, P2_R1200_U95);
  nand ginst14531 (P2_R1200_U468, P2_R1200_U180, P2_R1200_U319);
  nand ginst14532 (P2_R1200_U469, P2_R1200_U70, P2_U3431);
  not ginst14533 (P2_R1200_U47, P2_U3082);
  nand ginst14534 (P2_R1200_U470, P2_R1200_U67, P2_U3078);
  nand ginst14535 (P2_R1200_U471, P2_R1200_U182, P2_R1200_U328);
  nand ginst14536 (P2_R1200_U472, P2_R1200_U181, P2_R1200_U256);
  nand ginst14537 (P2_R1200_U473, P2_R1200_U64, P2_U3428);
  nand ginst14538 (P2_R1200_U474, P2_R1200_U63, P2_U3079);
  not ginst14539 (P2_R1200_U475, P2_R1200_U152);
  nand ginst14540 (P2_R1200_U476, P2_R1200_U354, P2_R1200_U475);
  nand ginst14541 (P2_R1200_U477, P2_R1200_U152, P2_R1200_U183);
  nand ginst14542 (P2_R1200_U478, P2_R1200_U55, P2_U3425);
  nand ginst14543 (P2_R1200_U479, P2_R1200_U61, P2_U3071);
  nand ginst14544 (P2_R1200_U48, P2_R1200_U217, P2_R1200_U45);
  not ginst14545 (P2_R1200_U480, P2_R1200_U153);
  nand ginst14546 (P2_R1200_U481, P2_R1200_U352, P2_R1200_U480);
  nand ginst14547 (P2_R1200_U482, P2_R1200_U153, P2_R1200_U184);
  nand ginst14548 (P2_R1200_U483, P2_R1200_U56, P2_U3422);
  nand ginst14549 (P2_R1200_U484, P2_R1200_U60, P2_U3062);
  nand ginst14550 (P2_R1200_U485, P2_R1200_U483, P2_R1200_U484);
  nand ginst14551 (P2_R1200_U486, P2_R1200_U57, P2_U3419);
  nand ginst14552 (P2_R1200_U487, P2_R1200_U58, P2_U3061);
  nand ginst14553 (P2_R1200_U488, P2_R1200_U336, P2_R1200_U96);
  nand ginst14554 (P2_R1200_U489, P2_R1200_U185, P2_R1200_U350);
  nand ginst14555 (P2_R1200_U49, P2_R1200_U231, P2_R1200_U44);
  nand ginst14556 (P2_R1200_U50, P2_R1200_U188, P2_R1200_U204, P2_R1200_U338);
  not ginst14557 (P2_R1200_U51, P2_U3895);
  not ginst14558 (P2_R1200_U52, P2_U3056);
  nand ginst14559 (P2_R1200_U53, P2_R1200_U90, P2_U3056);
  not ginst14560 (P2_R1200_U54, P2_U3052);
  not ginst14561 (P2_R1200_U55, P2_U3071);
  not ginst14562 (P2_R1200_U56, P2_U3062);
  not ginst14563 (P2_R1200_U57, P2_U3061);
  not ginst14564 (P2_R1200_U58, P2_U3419);
  nand ginst14565 (P2_R1200_U59, P2_R1200_U46, P2_U3082);
  and ginst14566 (P2_R1200_U6, P2_R1200_U211, P2_R1200_U212);
  not ginst14567 (P2_R1200_U60, P2_U3422);
  not ginst14568 (P2_R1200_U61, P2_U3425);
  nand ginst14569 (P2_R1200_U62, P2_R1200_U248, P2_R1200_U249);
  not ginst14570 (P2_R1200_U63, P2_U3428);
  not ginst14571 (P2_R1200_U64, P2_U3079);
  not ginst14572 (P2_R1200_U65, P2_U3437);
  not ginst14573 (P2_R1200_U66, P2_U3434);
  not ginst14574 (P2_R1200_U67, P2_U3431);
  not ginst14575 (P2_R1200_U68, P2_U3072);
  not ginst14576 (P2_R1200_U69, P2_U3073);
  and ginst14577 (P2_R1200_U7, P2_R1200_U245, P2_R1200_U246);
  not ginst14578 (P2_R1200_U70, P2_U3078);
  nand ginst14579 (P2_R1200_U71, P2_R1200_U67, P2_U3078);
  not ginst14580 (P2_R1200_U72, P2_U3440);
  not ginst14581 (P2_R1200_U73, P2_U3068);
  not ginst14582 (P2_R1200_U74, P2_U3081);
  not ginst14583 (P2_R1200_U75, P2_U3445);
  not ginst14584 (P2_R1200_U76, P2_U3080);
  not ginst14585 (P2_R1200_U77, P2_U3903);
  not ginst14586 (P2_R1200_U78, P2_U3075);
  not ginst14587 (P2_R1200_U79, P2_U3900);
  and ginst14588 (P2_R1200_U8, P2_R1200_U193, P2_R1200_U257);
  not ginst14589 (P2_R1200_U80, P2_U3901);
  not ginst14590 (P2_R1200_U81, P2_U3902);
  not ginst14591 (P2_R1200_U82, P2_U3065);
  not ginst14592 (P2_R1200_U83, P2_U3060);
  not ginst14593 (P2_R1200_U84, P2_U3074);
  nand ginst14594 (P2_R1200_U85, P2_R1200_U81, P2_U3074);
  not ginst14595 (P2_R1200_U86, P2_U3899);
  not ginst14596 (P2_R1200_U87, P2_U3064);
  not ginst14597 (P2_R1200_U88, P2_U3898);
  not ginst14598 (P2_R1200_U89, P2_U3057);
  and ginst14599 (P2_R1200_U9, P2_R1200_U258, P2_R1200_U259);
  not ginst14600 (P2_R1200_U90, P2_U3897);
  not ginst14601 (P2_R1200_U91, P2_U3896);
  not ginst14602 (P2_R1200_U92, P2_U3053);
  nand ginst14603 (P2_R1200_U93, P2_R1200_U296, P2_R1200_U297);
  nand ginst14604 (P2_R1200_U94, P2_R1200_U307, P2_R1200_U85);
  nand ginst14605 (P2_R1200_U95, P2_R1200_U318, P2_R1200_U71);
  nand ginst14606 (P2_R1200_U96, P2_R1200_U349, P2_R1200_U59);
  not ginst14607 (P2_R1200_U97, P2_U3076);
  nand ginst14608 (P2_R1200_U98, P2_R1200_U405, P2_R1200_U406);
  nand ginst14609 (P2_R1200_U99, P2_R1200_U419, P2_R1200_U420);
  not ginst14610 (P2_R1209_U10, P2_REG1_REG_1__SCAN_IN);
  nand ginst14611 (P2_R1209_U100, P2_R1209_U150, P2_R1209_U151);
  nand ginst14612 (P2_R1209_U101, P2_R1209_U146, P2_R1209_U147);
  nand ginst14613 (P2_R1209_U102, P2_R1209_U142, P2_R1209_U143);
  nand ginst14614 (P2_R1209_U103, P2_R1209_U138, P2_R1209_U139);
  not ginst14615 (P2_R1209_U104, P2_R1209_U9);
  nand ginst14616 (P2_R1209_U105, P2_REG1_REG_1__SCAN_IN, P2_R1209_U104);
  nand ginst14617 (P2_R1209_U106, P2_R1209_U105, P2_U3391);
  nand ginst14618 (P2_R1209_U107, P2_R1209_U10, P2_R1209_U9);
  not ginst14619 (P2_R1209_U108, P2_R1209_U94);
  nand ginst14620 (P2_R1209_U109, P2_REG1_REG_2__SCAN_IN, P2_R1209_U13);
  not ginst14621 (P2_R1209_U11, P2_U3391);
  nand ginst14622 (P2_R1209_U110, P2_R1209_U109, P2_R1209_U94);
  nand ginst14623 (P2_R1209_U111, P2_R1209_U12, P2_U3394);
  not ginst14624 (P2_R1209_U112, P2_R1209_U93);
  nand ginst14625 (P2_R1209_U113, P2_REG1_REG_3__SCAN_IN, P2_R1209_U15);
  nand ginst14626 (P2_R1209_U114, P2_R1209_U113, P2_R1209_U93);
  nand ginst14627 (P2_R1209_U115, P2_R1209_U14, P2_U3397);
  not ginst14628 (P2_R1209_U116, P2_R1209_U92);
  nand ginst14629 (P2_R1209_U117, P2_REG1_REG_4__SCAN_IN, P2_R1209_U17);
  nand ginst14630 (P2_R1209_U118, P2_R1209_U117, P2_R1209_U92);
  nand ginst14631 (P2_R1209_U119, P2_R1209_U16, P2_U3400);
  not ginst14632 (P2_R1209_U12, P2_REG1_REG_2__SCAN_IN);
  not ginst14633 (P2_R1209_U120, P2_R1209_U91);
  nand ginst14634 (P2_R1209_U121, P2_REG1_REG_5__SCAN_IN, P2_R1209_U19);
  nand ginst14635 (P2_R1209_U122, P2_R1209_U121, P2_R1209_U91);
  nand ginst14636 (P2_R1209_U123, P2_R1209_U18, P2_U3403);
  not ginst14637 (P2_R1209_U124, P2_R1209_U90);
  nand ginst14638 (P2_R1209_U125, P2_REG1_REG_6__SCAN_IN, P2_R1209_U21);
  nand ginst14639 (P2_R1209_U126, P2_R1209_U125, P2_R1209_U90);
  nand ginst14640 (P2_R1209_U127, P2_R1209_U20, P2_U3406);
  not ginst14641 (P2_R1209_U128, P2_R1209_U89);
  nand ginst14642 (P2_R1209_U129, P2_REG1_REG_7__SCAN_IN, P2_R1209_U23);
  not ginst14643 (P2_R1209_U13, P2_U3394);
  nand ginst14644 (P2_R1209_U130, P2_R1209_U129, P2_R1209_U89);
  nand ginst14645 (P2_R1209_U131, P2_R1209_U22, P2_U3409);
  not ginst14646 (P2_R1209_U132, P2_R1209_U88);
  nand ginst14647 (P2_R1209_U133, P2_REG1_REG_8__SCAN_IN, P2_R1209_U25);
  nand ginst14648 (P2_R1209_U134, P2_R1209_U133, P2_R1209_U88);
  nand ginst14649 (P2_R1209_U135, P2_R1209_U24, P2_U3412);
  not ginst14650 (P2_R1209_U136, P2_R1209_U87);
  nand ginst14651 (P2_R1209_U137, P2_REG1_REG_9__SCAN_IN, P2_R1209_U27);
  nand ginst14652 (P2_R1209_U138, P2_R1209_U137, P2_R1209_U87);
  nand ginst14653 (P2_R1209_U139, P2_R1209_U26, P2_U3415);
  not ginst14654 (P2_R1209_U14, P2_REG1_REG_3__SCAN_IN);
  not ginst14655 (P2_R1209_U140, P2_R1209_U103);
  nand ginst14656 (P2_R1209_U141, P2_REG1_REG_10__SCAN_IN, P2_R1209_U29);
  nand ginst14657 (P2_R1209_U142, P2_R1209_U103, P2_R1209_U141);
  nand ginst14658 (P2_R1209_U143, P2_R1209_U28, P2_U3418);
  not ginst14659 (P2_R1209_U144, P2_R1209_U102);
  nand ginst14660 (P2_R1209_U145, P2_REG1_REG_11__SCAN_IN, P2_R1209_U31);
  nand ginst14661 (P2_R1209_U146, P2_R1209_U102, P2_R1209_U145);
  nand ginst14662 (P2_R1209_U147, P2_R1209_U30, P2_U3421);
  not ginst14663 (P2_R1209_U148, P2_R1209_U101);
  nand ginst14664 (P2_R1209_U149, P2_REG1_REG_12__SCAN_IN, P2_R1209_U33);
  not ginst14665 (P2_R1209_U15, P2_U3397);
  nand ginst14666 (P2_R1209_U150, P2_R1209_U101, P2_R1209_U149);
  nand ginst14667 (P2_R1209_U151, P2_R1209_U32, P2_U3424);
  not ginst14668 (P2_R1209_U152, P2_R1209_U100);
  nand ginst14669 (P2_R1209_U153, P2_REG1_REG_13__SCAN_IN, P2_R1209_U35);
  nand ginst14670 (P2_R1209_U154, P2_R1209_U100, P2_R1209_U153);
  nand ginst14671 (P2_R1209_U155, P2_R1209_U34, P2_U3427);
  not ginst14672 (P2_R1209_U156, P2_R1209_U99);
  nand ginst14673 (P2_R1209_U157, P2_REG1_REG_14__SCAN_IN, P2_R1209_U37);
  nand ginst14674 (P2_R1209_U158, P2_R1209_U157, P2_R1209_U99);
  nand ginst14675 (P2_R1209_U159, P2_R1209_U36, P2_U3430);
  not ginst14676 (P2_R1209_U16, P2_REG1_REG_4__SCAN_IN);
  not ginst14677 (P2_R1209_U160, P2_R1209_U38);
  nand ginst14678 (P2_R1209_U161, P2_REG1_REG_15__SCAN_IN, P2_R1209_U160);
  nand ginst14679 (P2_R1209_U162, P2_R1209_U161, P2_U3433);
  nand ginst14680 (P2_R1209_U163, P2_R1209_U38, P2_R1209_U39);
  not ginst14681 (P2_R1209_U164, P2_R1209_U98);
  nand ginst14682 (P2_R1209_U165, P2_REG1_REG_16__SCAN_IN, P2_R1209_U42);
  nand ginst14683 (P2_R1209_U166, P2_R1209_U165, P2_R1209_U98);
  nand ginst14684 (P2_R1209_U167, P2_R1209_U41, P2_U3436);
  not ginst14685 (P2_R1209_U168, P2_R1209_U97);
  nand ginst14686 (P2_R1209_U169, P2_REG1_REG_17__SCAN_IN, P2_R1209_U44);
  not ginst14687 (P2_R1209_U17, P2_U3400);
  nand ginst14688 (P2_R1209_U170, P2_R1209_U169, P2_R1209_U97);
  nand ginst14689 (P2_R1209_U171, P2_R1209_U43, P2_U3439);
  not ginst14690 (P2_R1209_U172, P2_R1209_U47);
  nand ginst14691 (P2_R1209_U173, P2_R1209_U45, P2_U3442);
  nand ginst14692 (P2_R1209_U174, P2_R1209_U172, P2_R1209_U173);
  nand ginst14693 (P2_R1209_U175, P2_REG1_REG_18__SCAN_IN, P2_R1209_U46);
  nand ginst14694 (P2_R1209_U176, P2_R1209_U174, P2_R1209_U77);
  nand ginst14695 (P2_R1209_U177, P2_REG1_REG_18__SCAN_IN, P2_R1209_U46);
  nand ginst14696 (P2_R1209_U178, P2_R1209_U177, P2_R1209_U47);
  nand ginst14697 (P2_R1209_U179, P2_R1209_U45, P2_U3442);
  not ginst14698 (P2_R1209_U18, P2_REG1_REG_5__SCAN_IN);
  nand ginst14699 (P2_R1209_U180, P2_R1209_U178, P2_R1209_U76);
  nand ginst14700 (P2_R1209_U181, P2_R1209_U8, P2_U3386);
  nand ginst14701 (P2_R1209_U182, P2_REG1_REG_9__SCAN_IN, P2_R1209_U27);
  nand ginst14702 (P2_R1209_U183, P2_R1209_U26, P2_U3415);
  not ginst14703 (P2_R1209_U184, P2_R1209_U67);
  nand ginst14704 (P2_R1209_U185, P2_R1209_U136, P2_R1209_U184);
  nand ginst14705 (P2_R1209_U186, P2_R1209_U67, P2_R1209_U87);
  nand ginst14706 (P2_R1209_U187, P2_REG1_REG_8__SCAN_IN, P2_R1209_U25);
  nand ginst14707 (P2_R1209_U188, P2_R1209_U24, P2_U3412);
  not ginst14708 (P2_R1209_U189, P2_R1209_U68);
  not ginst14709 (P2_R1209_U19, P2_U3403);
  nand ginst14710 (P2_R1209_U190, P2_R1209_U132, P2_R1209_U189);
  nand ginst14711 (P2_R1209_U191, P2_R1209_U68, P2_R1209_U88);
  nand ginst14712 (P2_R1209_U192, P2_REG1_REG_7__SCAN_IN, P2_R1209_U23);
  nand ginst14713 (P2_R1209_U193, P2_R1209_U22, P2_U3409);
  not ginst14714 (P2_R1209_U194, P2_R1209_U69);
  nand ginst14715 (P2_R1209_U195, P2_R1209_U128, P2_R1209_U194);
  nand ginst14716 (P2_R1209_U196, P2_R1209_U69, P2_R1209_U89);
  nand ginst14717 (P2_R1209_U197, P2_REG1_REG_6__SCAN_IN, P2_R1209_U21);
  nand ginst14718 (P2_R1209_U198, P2_R1209_U20, P2_U3406);
  not ginst14719 (P2_R1209_U199, P2_R1209_U70);
  not ginst14720 (P2_R1209_U20, P2_REG1_REG_6__SCAN_IN);
  nand ginst14721 (P2_R1209_U200, P2_R1209_U124, P2_R1209_U199);
  nand ginst14722 (P2_R1209_U201, P2_R1209_U70, P2_R1209_U90);
  nand ginst14723 (P2_R1209_U202, P2_REG1_REG_5__SCAN_IN, P2_R1209_U19);
  nand ginst14724 (P2_R1209_U203, P2_R1209_U18, P2_U3403);
  not ginst14725 (P2_R1209_U204, P2_R1209_U71);
  nand ginst14726 (P2_R1209_U205, P2_R1209_U120, P2_R1209_U204);
  nand ginst14727 (P2_R1209_U206, P2_R1209_U71, P2_R1209_U91);
  nand ginst14728 (P2_R1209_U207, P2_REG1_REG_4__SCAN_IN, P2_R1209_U17);
  nand ginst14729 (P2_R1209_U208, P2_R1209_U16, P2_U3400);
  not ginst14730 (P2_R1209_U209, P2_R1209_U72);
  not ginst14731 (P2_R1209_U21, P2_U3406);
  nand ginst14732 (P2_R1209_U210, P2_R1209_U116, P2_R1209_U209);
  nand ginst14733 (P2_R1209_U211, P2_R1209_U72, P2_R1209_U92);
  nand ginst14734 (P2_R1209_U212, P2_REG1_REG_3__SCAN_IN, P2_R1209_U15);
  nand ginst14735 (P2_R1209_U213, P2_R1209_U14, P2_U3397);
  not ginst14736 (P2_R1209_U214, P2_R1209_U73);
  nand ginst14737 (P2_R1209_U215, P2_R1209_U112, P2_R1209_U214);
  nand ginst14738 (P2_R1209_U216, P2_R1209_U73, P2_R1209_U93);
  nand ginst14739 (P2_R1209_U217, P2_REG1_REG_2__SCAN_IN, P2_R1209_U13);
  nand ginst14740 (P2_R1209_U218, P2_R1209_U12, P2_U3394);
  not ginst14741 (P2_R1209_U219, P2_R1209_U74);
  not ginst14742 (P2_R1209_U22, P2_REG1_REG_7__SCAN_IN);
  nand ginst14743 (P2_R1209_U220, P2_R1209_U108, P2_R1209_U219);
  nand ginst14744 (P2_R1209_U221, P2_R1209_U74, P2_R1209_U94);
  nand ginst14745 (P2_R1209_U222, P2_R1209_U10, P2_R1209_U104);
  nand ginst14746 (P2_R1209_U223, P2_REG1_REG_1__SCAN_IN, P2_R1209_U9);
  not ginst14747 (P2_R1209_U224, P2_R1209_U75);
  nand ginst14748 (P2_R1209_U225, P2_R1209_U224, P2_U3391);
  nand ginst14749 (P2_R1209_U226, P2_R1209_U11, P2_R1209_U75);
  nand ginst14750 (P2_R1209_U227, P2_REG1_REG_19__SCAN_IN, P2_R1209_U96);
  nand ginst14751 (P2_R1209_U228, P2_R1209_U95, P2_U3379);
  nand ginst14752 (P2_R1209_U229, P2_REG1_REG_19__SCAN_IN, P2_R1209_U96);
  not ginst14753 (P2_R1209_U23, P2_U3409);
  nand ginst14754 (P2_R1209_U230, P2_R1209_U95, P2_U3379);
  nand ginst14755 (P2_R1209_U231, P2_R1209_U229, P2_R1209_U230);
  nand ginst14756 (P2_R1209_U232, P2_REG1_REG_18__SCAN_IN, P2_R1209_U46);
  nand ginst14757 (P2_R1209_U233, P2_R1209_U45, P2_U3442);
  not ginst14758 (P2_R1209_U234, P2_R1209_U78);
  nand ginst14759 (P2_R1209_U235, P2_R1209_U172, P2_R1209_U234);
  nand ginst14760 (P2_R1209_U236, P2_R1209_U47, P2_R1209_U78);
  nand ginst14761 (P2_R1209_U237, P2_REG1_REG_17__SCAN_IN, P2_R1209_U44);
  nand ginst14762 (P2_R1209_U238, P2_R1209_U43, P2_U3439);
  not ginst14763 (P2_R1209_U239, P2_R1209_U79);
  not ginst14764 (P2_R1209_U24, P2_REG1_REG_8__SCAN_IN);
  nand ginst14765 (P2_R1209_U240, P2_R1209_U168, P2_R1209_U239);
  nand ginst14766 (P2_R1209_U241, P2_R1209_U79, P2_R1209_U97);
  nand ginst14767 (P2_R1209_U242, P2_REG1_REG_16__SCAN_IN, P2_R1209_U42);
  nand ginst14768 (P2_R1209_U243, P2_R1209_U41, P2_U3436);
  not ginst14769 (P2_R1209_U244, P2_R1209_U80);
  nand ginst14770 (P2_R1209_U245, P2_R1209_U164, P2_R1209_U244);
  nand ginst14771 (P2_R1209_U246, P2_R1209_U80, P2_R1209_U98);
  nand ginst14772 (P2_R1209_U247, P2_R1209_U39, P2_U3433);
  nand ginst14773 (P2_R1209_U248, P2_REG1_REG_15__SCAN_IN, P2_R1209_U40);
  not ginst14774 (P2_R1209_U249, P2_R1209_U81);
  not ginst14775 (P2_R1209_U25, P2_U3412);
  nand ginst14776 (P2_R1209_U250, P2_R1209_U160, P2_R1209_U249);
  nand ginst14777 (P2_R1209_U251, P2_R1209_U38, P2_R1209_U81);
  nand ginst14778 (P2_R1209_U252, P2_REG1_REG_14__SCAN_IN, P2_R1209_U37);
  nand ginst14779 (P2_R1209_U253, P2_R1209_U36, P2_U3430);
  not ginst14780 (P2_R1209_U254, P2_R1209_U82);
  nand ginst14781 (P2_R1209_U255, P2_R1209_U156, P2_R1209_U254);
  nand ginst14782 (P2_R1209_U256, P2_R1209_U82, P2_R1209_U99);
  nand ginst14783 (P2_R1209_U257, P2_REG1_REG_13__SCAN_IN, P2_R1209_U35);
  nand ginst14784 (P2_R1209_U258, P2_R1209_U34, P2_U3427);
  not ginst14785 (P2_R1209_U259, P2_R1209_U83);
  not ginst14786 (P2_R1209_U26, P2_REG1_REG_9__SCAN_IN);
  nand ginst14787 (P2_R1209_U260, P2_R1209_U152, P2_R1209_U259);
  nand ginst14788 (P2_R1209_U261, P2_R1209_U100, P2_R1209_U83);
  nand ginst14789 (P2_R1209_U262, P2_REG1_REG_12__SCAN_IN, P2_R1209_U33);
  nand ginst14790 (P2_R1209_U263, P2_R1209_U32, P2_U3424);
  not ginst14791 (P2_R1209_U264, P2_R1209_U84);
  nand ginst14792 (P2_R1209_U265, P2_R1209_U148, P2_R1209_U264);
  nand ginst14793 (P2_R1209_U266, P2_R1209_U101, P2_R1209_U84);
  nand ginst14794 (P2_R1209_U267, P2_REG1_REG_11__SCAN_IN, P2_R1209_U31);
  nand ginst14795 (P2_R1209_U268, P2_R1209_U30, P2_U3421);
  not ginst14796 (P2_R1209_U269, P2_R1209_U85);
  not ginst14797 (P2_R1209_U27, P2_U3415);
  nand ginst14798 (P2_R1209_U270, P2_R1209_U144, P2_R1209_U269);
  nand ginst14799 (P2_R1209_U271, P2_R1209_U102, P2_R1209_U85);
  nand ginst14800 (P2_R1209_U272, P2_REG1_REG_10__SCAN_IN, P2_R1209_U29);
  nand ginst14801 (P2_R1209_U273, P2_R1209_U28, P2_U3418);
  not ginst14802 (P2_R1209_U274, P2_R1209_U86);
  nand ginst14803 (P2_R1209_U275, P2_R1209_U140, P2_R1209_U274);
  nand ginst14804 (P2_R1209_U276, P2_R1209_U103, P2_R1209_U86);
  not ginst14805 (P2_R1209_U28, P2_REG1_REG_10__SCAN_IN);
  not ginst14806 (P2_R1209_U29, P2_U3418);
  not ginst14807 (P2_R1209_U30, P2_REG1_REG_11__SCAN_IN);
  not ginst14808 (P2_R1209_U31, P2_U3421);
  not ginst14809 (P2_R1209_U32, P2_REG1_REG_12__SCAN_IN);
  not ginst14810 (P2_R1209_U33, P2_U3424);
  not ginst14811 (P2_R1209_U34, P2_REG1_REG_13__SCAN_IN);
  not ginst14812 (P2_R1209_U35, P2_U3427);
  not ginst14813 (P2_R1209_U36, P2_REG1_REG_14__SCAN_IN);
  not ginst14814 (P2_R1209_U37, P2_U3430);
  nand ginst14815 (P2_R1209_U38, P2_R1209_U158, P2_R1209_U159);
  not ginst14816 (P2_R1209_U39, P2_REG1_REG_15__SCAN_IN);
  not ginst14817 (P2_R1209_U40, P2_U3433);
  not ginst14818 (P2_R1209_U41, P2_REG1_REG_16__SCAN_IN);
  not ginst14819 (P2_R1209_U42, P2_U3436);
  not ginst14820 (P2_R1209_U43, P2_REG1_REG_17__SCAN_IN);
  not ginst14821 (P2_R1209_U44, P2_U3439);
  not ginst14822 (P2_R1209_U45, P2_REG1_REG_18__SCAN_IN);
  not ginst14823 (P2_R1209_U46, P2_U3442);
  nand ginst14824 (P2_R1209_U47, P2_R1209_U170, P2_R1209_U171);
  not ginst14825 (P2_R1209_U48, P2_U3386);
  nand ginst14826 (P2_R1209_U49, P2_R1209_U185, P2_R1209_U186);
  nand ginst14827 (P2_R1209_U50, P2_R1209_U190, P2_R1209_U191);
  nand ginst14828 (P2_R1209_U51, P2_R1209_U195, P2_R1209_U196);
  nand ginst14829 (P2_R1209_U52, P2_R1209_U200, P2_R1209_U201);
  nand ginst14830 (P2_R1209_U53, P2_R1209_U205, P2_R1209_U206);
  nand ginst14831 (P2_R1209_U54, P2_R1209_U210, P2_R1209_U211);
  nand ginst14832 (P2_R1209_U55, P2_R1209_U215, P2_R1209_U216);
  nand ginst14833 (P2_R1209_U56, P2_R1209_U220, P2_R1209_U221);
  nand ginst14834 (P2_R1209_U57, P2_R1209_U225, P2_R1209_U226);
  nand ginst14835 (P2_R1209_U58, P2_R1209_U235, P2_R1209_U236);
  nand ginst14836 (P2_R1209_U59, P2_R1209_U240, P2_R1209_U241);
  nand ginst14837 (P2_R1209_U6, P2_R1209_U176, P2_R1209_U180);
  nand ginst14838 (P2_R1209_U60, P2_R1209_U245, P2_R1209_U246);
  nand ginst14839 (P2_R1209_U61, P2_R1209_U250, P2_R1209_U251);
  nand ginst14840 (P2_R1209_U62, P2_R1209_U255, P2_R1209_U256);
  nand ginst14841 (P2_R1209_U63, P2_R1209_U260, P2_R1209_U261);
  nand ginst14842 (P2_R1209_U64, P2_R1209_U265, P2_R1209_U266);
  nand ginst14843 (P2_R1209_U65, P2_R1209_U270, P2_R1209_U271);
  nand ginst14844 (P2_R1209_U66, P2_R1209_U275, P2_R1209_U276);
  nand ginst14845 (P2_R1209_U67, P2_R1209_U182, P2_R1209_U183);
  nand ginst14846 (P2_R1209_U68, P2_R1209_U187, P2_R1209_U188);
  nand ginst14847 (P2_R1209_U69, P2_R1209_U192, P2_R1209_U193);
  nand ginst14848 (P2_R1209_U7, P2_R1209_U181, P2_R1209_U9);
  nand ginst14849 (P2_R1209_U70, P2_R1209_U197, P2_R1209_U198);
  nand ginst14850 (P2_R1209_U71, P2_R1209_U202, P2_R1209_U203);
  nand ginst14851 (P2_R1209_U72, P2_R1209_U207, P2_R1209_U208);
  nand ginst14852 (P2_R1209_U73, P2_R1209_U212, P2_R1209_U213);
  nand ginst14853 (P2_R1209_U74, P2_R1209_U217, P2_R1209_U218);
  nand ginst14854 (P2_R1209_U75, P2_R1209_U222, P2_R1209_U223);
  and ginst14855 (P2_R1209_U76, P2_R1209_U179, P2_R1209_U227, P2_R1209_U228);
  and ginst14856 (P2_R1209_U77, P2_R1209_U175, P2_R1209_U231);
  nand ginst14857 (P2_R1209_U78, P2_R1209_U232, P2_R1209_U233);
  nand ginst14858 (P2_R1209_U79, P2_R1209_U237, P2_R1209_U238);
  not ginst14859 (P2_R1209_U8, P2_REG1_REG_0__SCAN_IN);
  nand ginst14860 (P2_R1209_U80, P2_R1209_U242, P2_R1209_U243);
  nand ginst14861 (P2_R1209_U81, P2_R1209_U247, P2_R1209_U248);
  nand ginst14862 (P2_R1209_U82, P2_R1209_U252, P2_R1209_U253);
  nand ginst14863 (P2_R1209_U83, P2_R1209_U257, P2_R1209_U258);
  nand ginst14864 (P2_R1209_U84, P2_R1209_U262, P2_R1209_U263);
  nand ginst14865 (P2_R1209_U85, P2_R1209_U267, P2_R1209_U268);
  nand ginst14866 (P2_R1209_U86, P2_R1209_U272, P2_R1209_U273);
  nand ginst14867 (P2_R1209_U87, P2_R1209_U134, P2_R1209_U135);
  nand ginst14868 (P2_R1209_U88, P2_R1209_U130, P2_R1209_U131);
  nand ginst14869 (P2_R1209_U89, P2_R1209_U126, P2_R1209_U127);
  nand ginst14870 (P2_R1209_U9, P2_REG1_REG_0__SCAN_IN, P2_R1209_U48);
  nand ginst14871 (P2_R1209_U90, P2_R1209_U122, P2_R1209_U123);
  nand ginst14872 (P2_R1209_U91, P2_R1209_U118, P2_R1209_U119);
  nand ginst14873 (P2_R1209_U92, P2_R1209_U114, P2_R1209_U115);
  nand ginst14874 (P2_R1209_U93, P2_R1209_U110, P2_R1209_U111);
  nand ginst14875 (P2_R1209_U94, P2_R1209_U106, P2_R1209_U107);
  not ginst14876 (P2_R1209_U95, P2_REG1_REG_19__SCAN_IN);
  not ginst14877 (P2_R1209_U96, P2_U3379);
  nand ginst14878 (P2_R1209_U97, P2_R1209_U166, P2_R1209_U167);
  nand ginst14879 (P2_R1209_U98, P2_R1209_U162, P2_R1209_U163);
  nand ginst14880 (P2_R1209_U99, P2_R1209_U154, P2_R1209_U155);
  not ginst14881 (P2_R1212_U10, P2_REG2_REG_1__SCAN_IN);
  nand ginst14882 (P2_R1212_U100, P2_R1212_U150, P2_R1212_U151);
  nand ginst14883 (P2_R1212_U101, P2_R1212_U146, P2_R1212_U147);
  nand ginst14884 (P2_R1212_U102, P2_R1212_U142, P2_R1212_U143);
  nand ginst14885 (P2_R1212_U103, P2_R1212_U138, P2_R1212_U139);
  not ginst14886 (P2_R1212_U104, P2_R1212_U9);
  nand ginst14887 (P2_R1212_U105, P2_REG2_REG_1__SCAN_IN, P2_R1212_U104);
  nand ginst14888 (P2_R1212_U106, P2_R1212_U105, P2_U3391);
  nand ginst14889 (P2_R1212_U107, P2_R1212_U10, P2_R1212_U9);
  not ginst14890 (P2_R1212_U108, P2_R1212_U94);
  nand ginst14891 (P2_R1212_U109, P2_REG2_REG_2__SCAN_IN, P2_R1212_U13);
  not ginst14892 (P2_R1212_U11, P2_U3391);
  nand ginst14893 (P2_R1212_U110, P2_R1212_U109, P2_R1212_U94);
  nand ginst14894 (P2_R1212_U111, P2_R1212_U12, P2_U3394);
  not ginst14895 (P2_R1212_U112, P2_R1212_U93);
  nand ginst14896 (P2_R1212_U113, P2_REG2_REG_3__SCAN_IN, P2_R1212_U15);
  nand ginst14897 (P2_R1212_U114, P2_R1212_U113, P2_R1212_U93);
  nand ginst14898 (P2_R1212_U115, P2_R1212_U14, P2_U3397);
  not ginst14899 (P2_R1212_U116, P2_R1212_U92);
  nand ginst14900 (P2_R1212_U117, P2_REG2_REG_4__SCAN_IN, P2_R1212_U17);
  nand ginst14901 (P2_R1212_U118, P2_R1212_U117, P2_R1212_U92);
  nand ginst14902 (P2_R1212_U119, P2_R1212_U16, P2_U3400);
  not ginst14903 (P2_R1212_U12, P2_REG2_REG_2__SCAN_IN);
  not ginst14904 (P2_R1212_U120, P2_R1212_U91);
  nand ginst14905 (P2_R1212_U121, P2_REG2_REG_5__SCAN_IN, P2_R1212_U19);
  nand ginst14906 (P2_R1212_U122, P2_R1212_U121, P2_R1212_U91);
  nand ginst14907 (P2_R1212_U123, P2_R1212_U18, P2_U3403);
  not ginst14908 (P2_R1212_U124, P2_R1212_U90);
  nand ginst14909 (P2_R1212_U125, P2_REG2_REG_6__SCAN_IN, P2_R1212_U21);
  nand ginst14910 (P2_R1212_U126, P2_R1212_U125, P2_R1212_U90);
  nand ginst14911 (P2_R1212_U127, P2_R1212_U20, P2_U3406);
  not ginst14912 (P2_R1212_U128, P2_R1212_U89);
  nand ginst14913 (P2_R1212_U129, P2_REG2_REG_7__SCAN_IN, P2_R1212_U23);
  not ginst14914 (P2_R1212_U13, P2_U3394);
  nand ginst14915 (P2_R1212_U130, P2_R1212_U129, P2_R1212_U89);
  nand ginst14916 (P2_R1212_U131, P2_R1212_U22, P2_U3409);
  not ginst14917 (P2_R1212_U132, P2_R1212_U88);
  nand ginst14918 (P2_R1212_U133, P2_REG2_REG_8__SCAN_IN, P2_R1212_U25);
  nand ginst14919 (P2_R1212_U134, P2_R1212_U133, P2_R1212_U88);
  nand ginst14920 (P2_R1212_U135, P2_R1212_U24, P2_U3412);
  not ginst14921 (P2_R1212_U136, P2_R1212_U87);
  nand ginst14922 (P2_R1212_U137, P2_REG2_REG_9__SCAN_IN, P2_R1212_U27);
  nand ginst14923 (P2_R1212_U138, P2_R1212_U137, P2_R1212_U87);
  nand ginst14924 (P2_R1212_U139, P2_R1212_U26, P2_U3415);
  not ginst14925 (P2_R1212_U14, P2_REG2_REG_3__SCAN_IN);
  not ginst14926 (P2_R1212_U140, P2_R1212_U103);
  nand ginst14927 (P2_R1212_U141, P2_REG2_REG_10__SCAN_IN, P2_R1212_U29);
  nand ginst14928 (P2_R1212_U142, P2_R1212_U103, P2_R1212_U141);
  nand ginst14929 (P2_R1212_U143, P2_R1212_U28, P2_U3418);
  not ginst14930 (P2_R1212_U144, P2_R1212_U102);
  nand ginst14931 (P2_R1212_U145, P2_REG2_REG_11__SCAN_IN, P2_R1212_U31);
  nand ginst14932 (P2_R1212_U146, P2_R1212_U102, P2_R1212_U145);
  nand ginst14933 (P2_R1212_U147, P2_R1212_U30, P2_U3421);
  not ginst14934 (P2_R1212_U148, P2_R1212_U101);
  nand ginst14935 (P2_R1212_U149, P2_REG2_REG_12__SCAN_IN, P2_R1212_U33);
  not ginst14936 (P2_R1212_U15, P2_U3397);
  nand ginst14937 (P2_R1212_U150, P2_R1212_U101, P2_R1212_U149);
  nand ginst14938 (P2_R1212_U151, P2_R1212_U32, P2_U3424);
  not ginst14939 (P2_R1212_U152, P2_R1212_U100);
  nand ginst14940 (P2_R1212_U153, P2_REG2_REG_13__SCAN_IN, P2_R1212_U35);
  nand ginst14941 (P2_R1212_U154, P2_R1212_U100, P2_R1212_U153);
  nand ginst14942 (P2_R1212_U155, P2_R1212_U34, P2_U3427);
  not ginst14943 (P2_R1212_U156, P2_R1212_U99);
  nand ginst14944 (P2_R1212_U157, P2_REG2_REG_14__SCAN_IN, P2_R1212_U37);
  nand ginst14945 (P2_R1212_U158, P2_R1212_U157, P2_R1212_U99);
  nand ginst14946 (P2_R1212_U159, P2_R1212_U36, P2_U3430);
  not ginst14947 (P2_R1212_U16, P2_REG2_REG_4__SCAN_IN);
  not ginst14948 (P2_R1212_U160, P2_R1212_U38);
  nand ginst14949 (P2_R1212_U161, P2_REG2_REG_15__SCAN_IN, P2_R1212_U160);
  nand ginst14950 (P2_R1212_U162, P2_R1212_U161, P2_U3433);
  nand ginst14951 (P2_R1212_U163, P2_R1212_U38, P2_R1212_U39);
  not ginst14952 (P2_R1212_U164, P2_R1212_U98);
  nand ginst14953 (P2_R1212_U165, P2_REG2_REG_16__SCAN_IN, P2_R1212_U42);
  nand ginst14954 (P2_R1212_U166, P2_R1212_U165, P2_R1212_U98);
  nand ginst14955 (P2_R1212_U167, P2_R1212_U41, P2_U3436);
  not ginst14956 (P2_R1212_U168, P2_R1212_U97);
  nand ginst14957 (P2_R1212_U169, P2_REG2_REG_17__SCAN_IN, P2_R1212_U44);
  not ginst14958 (P2_R1212_U17, P2_U3400);
  nand ginst14959 (P2_R1212_U170, P2_R1212_U169, P2_R1212_U97);
  nand ginst14960 (P2_R1212_U171, P2_R1212_U43, P2_U3439);
  not ginst14961 (P2_R1212_U172, P2_R1212_U47);
  nand ginst14962 (P2_R1212_U173, P2_R1212_U45, P2_U3442);
  nand ginst14963 (P2_R1212_U174, P2_R1212_U172, P2_R1212_U173);
  nand ginst14964 (P2_R1212_U175, P2_REG2_REG_18__SCAN_IN, P2_R1212_U46);
  nand ginst14965 (P2_R1212_U176, P2_R1212_U174, P2_R1212_U77);
  nand ginst14966 (P2_R1212_U177, P2_REG2_REG_18__SCAN_IN, P2_R1212_U46);
  nand ginst14967 (P2_R1212_U178, P2_R1212_U177, P2_R1212_U47);
  nand ginst14968 (P2_R1212_U179, P2_R1212_U45, P2_U3442);
  not ginst14969 (P2_R1212_U18, P2_REG2_REG_5__SCAN_IN);
  nand ginst14970 (P2_R1212_U180, P2_R1212_U178, P2_R1212_U76);
  nand ginst14971 (P2_R1212_U181, P2_R1212_U8, P2_U3386);
  nand ginst14972 (P2_R1212_U182, P2_REG2_REG_9__SCAN_IN, P2_R1212_U27);
  nand ginst14973 (P2_R1212_U183, P2_R1212_U26, P2_U3415);
  not ginst14974 (P2_R1212_U184, P2_R1212_U67);
  nand ginst14975 (P2_R1212_U185, P2_R1212_U136, P2_R1212_U184);
  nand ginst14976 (P2_R1212_U186, P2_R1212_U67, P2_R1212_U87);
  nand ginst14977 (P2_R1212_U187, P2_REG2_REG_8__SCAN_IN, P2_R1212_U25);
  nand ginst14978 (P2_R1212_U188, P2_R1212_U24, P2_U3412);
  not ginst14979 (P2_R1212_U189, P2_R1212_U68);
  not ginst14980 (P2_R1212_U19, P2_U3403);
  nand ginst14981 (P2_R1212_U190, P2_R1212_U132, P2_R1212_U189);
  nand ginst14982 (P2_R1212_U191, P2_R1212_U68, P2_R1212_U88);
  nand ginst14983 (P2_R1212_U192, P2_REG2_REG_7__SCAN_IN, P2_R1212_U23);
  nand ginst14984 (P2_R1212_U193, P2_R1212_U22, P2_U3409);
  not ginst14985 (P2_R1212_U194, P2_R1212_U69);
  nand ginst14986 (P2_R1212_U195, P2_R1212_U128, P2_R1212_U194);
  nand ginst14987 (P2_R1212_U196, P2_R1212_U69, P2_R1212_U89);
  nand ginst14988 (P2_R1212_U197, P2_REG2_REG_6__SCAN_IN, P2_R1212_U21);
  nand ginst14989 (P2_R1212_U198, P2_R1212_U20, P2_U3406);
  not ginst14990 (P2_R1212_U199, P2_R1212_U70);
  not ginst14991 (P2_R1212_U20, P2_REG2_REG_6__SCAN_IN);
  nand ginst14992 (P2_R1212_U200, P2_R1212_U124, P2_R1212_U199);
  nand ginst14993 (P2_R1212_U201, P2_R1212_U70, P2_R1212_U90);
  nand ginst14994 (P2_R1212_U202, P2_REG2_REG_5__SCAN_IN, P2_R1212_U19);
  nand ginst14995 (P2_R1212_U203, P2_R1212_U18, P2_U3403);
  not ginst14996 (P2_R1212_U204, P2_R1212_U71);
  nand ginst14997 (P2_R1212_U205, P2_R1212_U120, P2_R1212_U204);
  nand ginst14998 (P2_R1212_U206, P2_R1212_U71, P2_R1212_U91);
  nand ginst14999 (P2_R1212_U207, P2_REG2_REG_4__SCAN_IN, P2_R1212_U17);
  nand ginst15000 (P2_R1212_U208, P2_R1212_U16, P2_U3400);
  not ginst15001 (P2_R1212_U209, P2_R1212_U72);
  not ginst15002 (P2_R1212_U21, P2_U3406);
  nand ginst15003 (P2_R1212_U210, P2_R1212_U116, P2_R1212_U209);
  nand ginst15004 (P2_R1212_U211, P2_R1212_U72, P2_R1212_U92);
  nand ginst15005 (P2_R1212_U212, P2_REG2_REG_3__SCAN_IN, P2_R1212_U15);
  nand ginst15006 (P2_R1212_U213, P2_R1212_U14, P2_U3397);
  not ginst15007 (P2_R1212_U214, P2_R1212_U73);
  nand ginst15008 (P2_R1212_U215, P2_R1212_U112, P2_R1212_U214);
  nand ginst15009 (P2_R1212_U216, P2_R1212_U73, P2_R1212_U93);
  nand ginst15010 (P2_R1212_U217, P2_REG2_REG_2__SCAN_IN, P2_R1212_U13);
  nand ginst15011 (P2_R1212_U218, P2_R1212_U12, P2_U3394);
  not ginst15012 (P2_R1212_U219, P2_R1212_U74);
  not ginst15013 (P2_R1212_U22, P2_REG2_REG_7__SCAN_IN);
  nand ginst15014 (P2_R1212_U220, P2_R1212_U108, P2_R1212_U219);
  nand ginst15015 (P2_R1212_U221, P2_R1212_U74, P2_R1212_U94);
  nand ginst15016 (P2_R1212_U222, P2_R1212_U10, P2_R1212_U104);
  nand ginst15017 (P2_R1212_U223, P2_REG2_REG_1__SCAN_IN, P2_R1212_U9);
  not ginst15018 (P2_R1212_U224, P2_R1212_U75);
  nand ginst15019 (P2_R1212_U225, P2_R1212_U224, P2_U3391);
  nand ginst15020 (P2_R1212_U226, P2_R1212_U11, P2_R1212_U75);
  nand ginst15021 (P2_R1212_U227, P2_REG2_REG_19__SCAN_IN, P2_R1212_U96);
  nand ginst15022 (P2_R1212_U228, P2_R1212_U95, P2_U3379);
  nand ginst15023 (P2_R1212_U229, P2_REG2_REG_19__SCAN_IN, P2_R1212_U96);
  not ginst15024 (P2_R1212_U23, P2_U3409);
  nand ginst15025 (P2_R1212_U230, P2_R1212_U95, P2_U3379);
  nand ginst15026 (P2_R1212_U231, P2_R1212_U229, P2_R1212_U230);
  nand ginst15027 (P2_R1212_U232, P2_REG2_REG_18__SCAN_IN, P2_R1212_U46);
  nand ginst15028 (P2_R1212_U233, P2_R1212_U45, P2_U3442);
  not ginst15029 (P2_R1212_U234, P2_R1212_U78);
  nand ginst15030 (P2_R1212_U235, P2_R1212_U172, P2_R1212_U234);
  nand ginst15031 (P2_R1212_U236, P2_R1212_U47, P2_R1212_U78);
  nand ginst15032 (P2_R1212_U237, P2_REG2_REG_17__SCAN_IN, P2_R1212_U44);
  nand ginst15033 (P2_R1212_U238, P2_R1212_U43, P2_U3439);
  not ginst15034 (P2_R1212_U239, P2_R1212_U79);
  not ginst15035 (P2_R1212_U24, P2_REG2_REG_8__SCAN_IN);
  nand ginst15036 (P2_R1212_U240, P2_R1212_U168, P2_R1212_U239);
  nand ginst15037 (P2_R1212_U241, P2_R1212_U79, P2_R1212_U97);
  nand ginst15038 (P2_R1212_U242, P2_REG2_REG_16__SCAN_IN, P2_R1212_U42);
  nand ginst15039 (P2_R1212_U243, P2_R1212_U41, P2_U3436);
  not ginst15040 (P2_R1212_U244, P2_R1212_U80);
  nand ginst15041 (P2_R1212_U245, P2_R1212_U164, P2_R1212_U244);
  nand ginst15042 (P2_R1212_U246, P2_R1212_U80, P2_R1212_U98);
  nand ginst15043 (P2_R1212_U247, P2_R1212_U39, P2_U3433);
  nand ginst15044 (P2_R1212_U248, P2_REG2_REG_15__SCAN_IN, P2_R1212_U40);
  not ginst15045 (P2_R1212_U249, P2_R1212_U81);
  not ginst15046 (P2_R1212_U25, P2_U3412);
  nand ginst15047 (P2_R1212_U250, P2_R1212_U160, P2_R1212_U249);
  nand ginst15048 (P2_R1212_U251, P2_R1212_U38, P2_R1212_U81);
  nand ginst15049 (P2_R1212_U252, P2_REG2_REG_14__SCAN_IN, P2_R1212_U37);
  nand ginst15050 (P2_R1212_U253, P2_R1212_U36, P2_U3430);
  not ginst15051 (P2_R1212_U254, P2_R1212_U82);
  nand ginst15052 (P2_R1212_U255, P2_R1212_U156, P2_R1212_U254);
  nand ginst15053 (P2_R1212_U256, P2_R1212_U82, P2_R1212_U99);
  nand ginst15054 (P2_R1212_U257, P2_REG2_REG_13__SCAN_IN, P2_R1212_U35);
  nand ginst15055 (P2_R1212_U258, P2_R1212_U34, P2_U3427);
  not ginst15056 (P2_R1212_U259, P2_R1212_U83);
  not ginst15057 (P2_R1212_U26, P2_REG2_REG_9__SCAN_IN);
  nand ginst15058 (P2_R1212_U260, P2_R1212_U152, P2_R1212_U259);
  nand ginst15059 (P2_R1212_U261, P2_R1212_U100, P2_R1212_U83);
  nand ginst15060 (P2_R1212_U262, P2_REG2_REG_12__SCAN_IN, P2_R1212_U33);
  nand ginst15061 (P2_R1212_U263, P2_R1212_U32, P2_U3424);
  not ginst15062 (P2_R1212_U264, P2_R1212_U84);
  nand ginst15063 (P2_R1212_U265, P2_R1212_U148, P2_R1212_U264);
  nand ginst15064 (P2_R1212_U266, P2_R1212_U101, P2_R1212_U84);
  nand ginst15065 (P2_R1212_U267, P2_REG2_REG_11__SCAN_IN, P2_R1212_U31);
  nand ginst15066 (P2_R1212_U268, P2_R1212_U30, P2_U3421);
  not ginst15067 (P2_R1212_U269, P2_R1212_U85);
  not ginst15068 (P2_R1212_U27, P2_U3415);
  nand ginst15069 (P2_R1212_U270, P2_R1212_U144, P2_R1212_U269);
  nand ginst15070 (P2_R1212_U271, P2_R1212_U102, P2_R1212_U85);
  nand ginst15071 (P2_R1212_U272, P2_REG2_REG_10__SCAN_IN, P2_R1212_U29);
  nand ginst15072 (P2_R1212_U273, P2_R1212_U28, P2_U3418);
  not ginst15073 (P2_R1212_U274, P2_R1212_U86);
  nand ginst15074 (P2_R1212_U275, P2_R1212_U140, P2_R1212_U274);
  nand ginst15075 (P2_R1212_U276, P2_R1212_U103, P2_R1212_U86);
  not ginst15076 (P2_R1212_U28, P2_REG2_REG_10__SCAN_IN);
  not ginst15077 (P2_R1212_U29, P2_U3418);
  not ginst15078 (P2_R1212_U30, P2_REG2_REG_11__SCAN_IN);
  not ginst15079 (P2_R1212_U31, P2_U3421);
  not ginst15080 (P2_R1212_U32, P2_REG2_REG_12__SCAN_IN);
  not ginst15081 (P2_R1212_U33, P2_U3424);
  not ginst15082 (P2_R1212_U34, P2_REG2_REG_13__SCAN_IN);
  not ginst15083 (P2_R1212_U35, P2_U3427);
  not ginst15084 (P2_R1212_U36, P2_REG2_REG_14__SCAN_IN);
  not ginst15085 (P2_R1212_U37, P2_U3430);
  nand ginst15086 (P2_R1212_U38, P2_R1212_U158, P2_R1212_U159);
  not ginst15087 (P2_R1212_U39, P2_REG2_REG_15__SCAN_IN);
  not ginst15088 (P2_R1212_U40, P2_U3433);
  not ginst15089 (P2_R1212_U41, P2_REG2_REG_16__SCAN_IN);
  not ginst15090 (P2_R1212_U42, P2_U3436);
  not ginst15091 (P2_R1212_U43, P2_REG2_REG_17__SCAN_IN);
  not ginst15092 (P2_R1212_U44, P2_U3439);
  not ginst15093 (P2_R1212_U45, P2_REG2_REG_18__SCAN_IN);
  not ginst15094 (P2_R1212_U46, P2_U3442);
  nand ginst15095 (P2_R1212_U47, P2_R1212_U170, P2_R1212_U171);
  not ginst15096 (P2_R1212_U48, P2_U3386);
  nand ginst15097 (P2_R1212_U49, P2_R1212_U185, P2_R1212_U186);
  nand ginst15098 (P2_R1212_U50, P2_R1212_U190, P2_R1212_U191);
  nand ginst15099 (P2_R1212_U51, P2_R1212_U195, P2_R1212_U196);
  nand ginst15100 (P2_R1212_U52, P2_R1212_U200, P2_R1212_U201);
  nand ginst15101 (P2_R1212_U53, P2_R1212_U205, P2_R1212_U206);
  nand ginst15102 (P2_R1212_U54, P2_R1212_U210, P2_R1212_U211);
  nand ginst15103 (P2_R1212_U55, P2_R1212_U215, P2_R1212_U216);
  nand ginst15104 (P2_R1212_U56, P2_R1212_U220, P2_R1212_U221);
  nand ginst15105 (P2_R1212_U57, P2_R1212_U225, P2_R1212_U226);
  nand ginst15106 (P2_R1212_U58, P2_R1212_U235, P2_R1212_U236);
  nand ginst15107 (P2_R1212_U59, P2_R1212_U240, P2_R1212_U241);
  nand ginst15108 (P2_R1212_U6, P2_R1212_U176, P2_R1212_U180);
  nand ginst15109 (P2_R1212_U60, P2_R1212_U245, P2_R1212_U246);
  nand ginst15110 (P2_R1212_U61, P2_R1212_U250, P2_R1212_U251);
  nand ginst15111 (P2_R1212_U62, P2_R1212_U255, P2_R1212_U256);
  nand ginst15112 (P2_R1212_U63, P2_R1212_U260, P2_R1212_U261);
  nand ginst15113 (P2_R1212_U64, P2_R1212_U265, P2_R1212_U266);
  nand ginst15114 (P2_R1212_U65, P2_R1212_U270, P2_R1212_U271);
  nand ginst15115 (P2_R1212_U66, P2_R1212_U275, P2_R1212_U276);
  nand ginst15116 (P2_R1212_U67, P2_R1212_U182, P2_R1212_U183);
  nand ginst15117 (P2_R1212_U68, P2_R1212_U187, P2_R1212_U188);
  nand ginst15118 (P2_R1212_U69, P2_R1212_U192, P2_R1212_U193);
  nand ginst15119 (P2_R1212_U7, P2_R1212_U181, P2_R1212_U9);
  nand ginst15120 (P2_R1212_U70, P2_R1212_U197, P2_R1212_U198);
  nand ginst15121 (P2_R1212_U71, P2_R1212_U202, P2_R1212_U203);
  nand ginst15122 (P2_R1212_U72, P2_R1212_U207, P2_R1212_U208);
  nand ginst15123 (P2_R1212_U73, P2_R1212_U212, P2_R1212_U213);
  nand ginst15124 (P2_R1212_U74, P2_R1212_U217, P2_R1212_U218);
  nand ginst15125 (P2_R1212_U75, P2_R1212_U222, P2_R1212_U223);
  and ginst15126 (P2_R1212_U76, P2_R1212_U179, P2_R1212_U227, P2_R1212_U228);
  and ginst15127 (P2_R1212_U77, P2_R1212_U175, P2_R1212_U231);
  nand ginst15128 (P2_R1212_U78, P2_R1212_U232, P2_R1212_U233);
  nand ginst15129 (P2_R1212_U79, P2_R1212_U237, P2_R1212_U238);
  not ginst15130 (P2_R1212_U8, P2_REG2_REG_0__SCAN_IN);
  nand ginst15131 (P2_R1212_U80, P2_R1212_U242, P2_R1212_U243);
  nand ginst15132 (P2_R1212_U81, P2_R1212_U247, P2_R1212_U248);
  nand ginst15133 (P2_R1212_U82, P2_R1212_U252, P2_R1212_U253);
  nand ginst15134 (P2_R1212_U83, P2_R1212_U257, P2_R1212_U258);
  nand ginst15135 (P2_R1212_U84, P2_R1212_U262, P2_R1212_U263);
  nand ginst15136 (P2_R1212_U85, P2_R1212_U267, P2_R1212_U268);
  nand ginst15137 (P2_R1212_U86, P2_R1212_U272, P2_R1212_U273);
  nand ginst15138 (P2_R1212_U87, P2_R1212_U134, P2_R1212_U135);
  nand ginst15139 (P2_R1212_U88, P2_R1212_U130, P2_R1212_U131);
  nand ginst15140 (P2_R1212_U89, P2_R1212_U126, P2_R1212_U127);
  nand ginst15141 (P2_R1212_U9, P2_REG2_REG_0__SCAN_IN, P2_R1212_U48);
  nand ginst15142 (P2_R1212_U90, P2_R1212_U122, P2_R1212_U123);
  nand ginst15143 (P2_R1212_U91, P2_R1212_U118, P2_R1212_U119);
  nand ginst15144 (P2_R1212_U92, P2_R1212_U114, P2_R1212_U115);
  nand ginst15145 (P2_R1212_U93, P2_R1212_U110, P2_R1212_U111);
  nand ginst15146 (P2_R1212_U94, P2_R1212_U106, P2_R1212_U107);
  not ginst15147 (P2_R1212_U95, P2_REG2_REG_19__SCAN_IN);
  not ginst15148 (P2_R1212_U96, P2_U3379);
  nand ginst15149 (P2_R1212_U97, P2_R1212_U166, P2_R1212_U167);
  nand ginst15150 (P2_R1212_U98, P2_R1212_U162, P2_R1212_U163);
  nand ginst15151 (P2_R1212_U99, P2_R1212_U154, P2_R1212_U155);
  and ginst15152 (P2_R1269_U10, P2_R1269_U146, P2_R1269_U147);
  and ginst15153 (P2_R1269_U100, P2_R1269_U55, P2_U3146);
  and ginst15154 (P2_R1269_U101, P2_R1269_U54, P2_U3145);
  and ginst15155 (P2_R1269_U102, P2_R1269_U103, P2_R1269_U13);
  and ginst15156 (P2_R1269_U103, P2_R1269_U168, P2_R1269_U169);
  and ginst15157 (P2_R1269_U104, P2_R1269_U102, P2_R1269_U167);
  and ginst15158 (P2_R1269_U105, P2_R1269_U56, P2_U3104);
  and ginst15159 (P2_R1269_U106, P2_R1269_U65, P2_U3105);
  and ginst15160 (P2_R1269_U107, P2_R1269_U109, P2_R1269_U172);
  and ginst15161 (P2_R1269_U108, P2_R1269_U107, P2_R1269_U173);
  and ginst15162 (P2_R1269_U109, P2_R1269_U174, P2_R1269_U175);
  and ginst15163 (P2_R1269_U11, P2_R1269_U148, P2_R1269_U94, P2_R1269_U95);
  and ginst15164 (P2_R1269_U110, P2_R1269_U139, P2_R1269_U185, P2_R1269_U186);
  and ginst15165 (P2_R1269_U111, P2_R1269_U189, P2_R1269_U190);
  and ginst15166 (P2_R1269_U112, P2_R1269_U73, P2_U3093);
  and ginst15167 (P2_R1269_U113, P2_R1269_U196, P2_R1269_U197);
  and ginst15168 (P2_R1269_U114, P2_R1269_U76, P2_U3122);
  and ginst15169 (P2_R1269_U115, P2_R1269_U79, P2_U3121);
  and ginst15170 (P2_R1269_U116, P2_R1269_U80, P2_U3120);
  and ginst15171 (P2_R1269_U117, P2_R1269_U116, P2_R1269_U123);
  and ginst15172 (P2_R1269_U118, P2_R1269_U78, P2_U3119);
  and ginst15173 (P2_R1269_U119, P2_R1269_U201, P2_R1269_U202);
  and ginst15174 (P2_R1269_U12, P2_R1269_U11, P2_R1269_U96);
  and ginst15175 (P2_R1269_U120, P2_R1269_U15, P2_R1269_U203, P2_R1269_U204);
  nand ginst15176 (P2_R1269_U121, P2_R1269_U198, P2_R1269_U199);
  nand ginst15177 (P2_R1269_U122, P2_R1269_U26, P2_U3086);
  nand ginst15178 (P2_R1269_U123, P2_R1269_U84, P2_U3087);
  nand ginst15179 (P2_R1269_U124, P2_R1269_U82, P2_U3089);
  nand ginst15180 (P2_R1269_U125, P2_R1269_U83, P2_U3088);
  nand ginst15181 (P2_R1269_U126, P2_R1269_U27, P2_U3085);
  nand ginst15182 (P2_R1269_U127, P2_R1269_U126, P2_R1269_U21, P2_R1269_U85);
  nand ginst15183 (P2_R1269_U128, P2_R1269_U205, P2_R1269_U208, P2_R1269_U209);
  nand ginst15184 (P2_R1269_U129, P2_R1269_U21, P2_R1269_U23, P2_U3117);
  and ginst15185 (P2_R1269_U13, P2_R1269_U162, P2_R1269_U163);
  nand ginst15186 (P2_R1269_U130, P2_R1269_U39, P2_U3129);
  nand ginst15187 (P2_R1269_U131, P2_R1269_U36, P2_U3130);
  nand ginst15188 (P2_R1269_U132, P2_R1269_U72, P2_U3094);
  nand ginst15189 (P2_R1269_U133, P2_R1269_U32, P2_U3095);
  nand ginst15190 (P2_R1269_U134, P2_R1269_U130, P2_R1269_U89);
  nand ginst15191 (P2_R1269_U135, P2_R1269_U6, P2_R1269_U90);
  nand ginst15192 (P2_R1269_U136, P2_R1269_U35, P2_U3097);
  nand ginst15193 (P2_R1269_U137, P2_R1269_U34, P2_U3096);
  nand ginst15194 (P2_R1269_U138, P2_R1269_U42, P2_U3100);
  nand ginst15195 (P2_R1269_U139, P2_R1269_U75, P2_U3124);
  and ginst15196 (P2_R1269_U14, P2_R1269_U113, P2_R1269_U191, P2_R1269_U195, P2_R1269_U20, P2_R1269_U21);
  nand ginst15197 (P2_R1269_U140, P2_R1269_U77, P2_U3123);
  nand ginst15198 (P2_R1269_U141, P2_R1269_U71, P2_U3101);
  nand ginst15199 (P2_R1269_U142, P2_R1269_U51, P2_U3141);
  nand ginst15200 (P2_R1269_U143, P2_R1269_U142, P2_R1269_U92);
  nand ginst15201 (P2_R1269_U144, P2_R1269_U64, P2_U3106);
  nand ginst15202 (P2_R1269_U145, P2_R1269_U58, P2_U3107);
  nand ginst15203 (P2_R1269_U146, P2_R1269_U46, P2_U3142);
  nand ginst15204 (P2_R1269_U147, P2_R1269_U51, P2_U3141);
  nand ginst15205 (P2_R1269_U148, P2_R1269_U10, P2_R1269_U93);
  nand ginst15206 (P2_R1269_U149, P2_R1269_U45, P2_U3109);
  and ginst15207 (P2_R1269_U15, P2_R1269_U128, P2_R1269_U129);
  nand ginst15208 (P2_R1269_U150, P2_R1269_U59, P2_U3108);
  nand ginst15209 (P2_R1269_U151, P2_R1269_U63, P2_U3112);
  nand ginst15210 (P2_R1269_U152, P2_R1269_U61, P2_U3113);
  nand ginst15211 (P2_R1269_U153, P2_U3147, P2_U3148);
  nand ginst15212 (P2_R1269_U154, P2_R1269_U153, P2_U3115);
  or ginst15213 (P2_R1269_U155, P2_U3147, P2_U3148);
  nand ginst15214 (P2_R1269_U156, P2_R1269_U60, P2_U3114);
  nand ginst15215 (P2_R1269_U157, P2_R1269_U12, P2_R1269_U97);
  nand ginst15216 (P2_R1269_U158, P2_R1269_U101, P2_R1269_U151);
  nand ginst15217 (P2_R1269_U159, P2_R1269_U50, P2_U3143);
  and ginst15218 (P2_R1269_U16, P2_R1269_U114, P2_R1269_U20, P2_R1269_U21);
  nand ginst15219 (P2_R1269_U160, P2_R1269_U53, P2_U3144);
  nand ginst15220 (P2_R1269_U161, P2_R1269_U10, P2_R1269_U158, P2_R1269_U159, P2_R1269_U160);
  nand ginst15221 (P2_R1269_U162, P2_R1269_U66, P2_U3136);
  nand ginst15222 (P2_R1269_U163, P2_R1269_U69, P2_U3135);
  nand ginst15223 (P2_R1269_U164, P2_R1269_U144, P2_R1269_U98);
  nand ginst15224 (P2_R1269_U165, P2_R1269_U9, P2_R1269_U99);
  nand ginst15225 (P2_R1269_U166, P2_R1269_U100, P2_R1269_U12);
  nand ginst15226 (P2_R1269_U167, P2_R1269_U11, P2_R1269_U161);
  nand ginst15227 (P2_R1269_U168, P2_R1269_U48, P2_U3138);
  nand ginst15228 (P2_R1269_U169, P2_R1269_U67, P2_U3137);
  and ginst15229 (P2_R1269_U17, P2_R1269_U115, P2_R1269_U20, P2_R1269_U21);
  nand ginst15230 (P2_R1269_U170, P2_R1269_U104, P2_R1269_U157, P2_R1269_U164, P2_R1269_U165, P2_R1269_U166);
  nand ginst15231 (P2_R1269_U171, P2_R1269_U69, P2_U3135);
  nand ginst15232 (P2_R1269_U172, P2_R1269_U105, P2_R1269_U171);
  nand ginst15233 (P2_R1269_U173, P2_R1269_U106, P2_R1269_U13);
  nand ginst15234 (P2_R1269_U174, P2_R1269_U70, P2_U3102);
  nand ginst15235 (P2_R1269_U175, P2_R1269_U57, P2_U3103);
  nand ginst15236 (P2_R1269_U176, P2_R1269_U108, P2_R1269_U170);
  nand ginst15237 (P2_R1269_U177, P2_R1269_U68, P2_U3134);
  nand ginst15238 (P2_R1269_U178, P2_R1269_U176, P2_R1269_U177);
  nand ginst15239 (P2_R1269_U179, P2_R1269_U141, P2_R1269_U178);
  and ginst15240 (P2_R1269_U18, P2_R1269_U117, P2_R1269_U21);
  nand ginst15241 (P2_R1269_U180, P2_R1269_U44, P2_U3133);
  nand ginst15242 (P2_R1269_U181, P2_R1269_U179, P2_R1269_U180);
  nand ginst15243 (P2_R1269_U182, P2_R1269_U38, P2_U3131);
  nand ginst15244 (P2_R1269_U183, P2_R1269_U43, P2_U3132);
  nand ginst15245 (P2_R1269_U184, P2_R1269_U6, P2_R1269_U88);
  nand ginst15246 (P2_R1269_U185, P2_R1269_U132, P2_R1269_U86);
  nand ginst15247 (P2_R1269_U186, P2_R1269_U7, P2_R1269_U87);
  nand ginst15248 (P2_R1269_U187, P2_R1269_U184, P2_R1269_U8);
  nand ginst15249 (P2_R1269_U188, P2_R1269_U138, P2_R1269_U181, P2_R1269_U8);
  nand ginst15250 (P2_R1269_U189, P2_R1269_U31, P2_U3126);
  and ginst15251 (P2_R1269_U19, P2_R1269_U118, P2_R1269_U21);
  nand ginst15252 (P2_R1269_U190, P2_R1269_U74, P2_U3125);
  nand ginst15253 (P2_R1269_U191, P2_R1269_U110, P2_R1269_U111, P2_R1269_U140, P2_R1269_U187, P2_R1269_U188);
  nand ginst15254 (P2_R1269_U192, P2_R1269_U112, P2_R1269_U139);
  nand ginst15255 (P2_R1269_U193, P2_R1269_U29, P2_U3092);
  nand ginst15256 (P2_R1269_U194, P2_R1269_U192, P2_R1269_U193);
  nand ginst15257 (P2_R1269_U195, P2_R1269_U140, P2_R1269_U194);
  nand ginst15258 (P2_R1269_U196, P2_R1269_U81, P2_U3090);
  nand ginst15259 (P2_R1269_U197, P2_R1269_U30, P2_U3091);
  nand ginst15260 (P2_R1269_U198, P2_R1269_U122, P2_U3117);
  nand ginst15261 (P2_R1269_U199, P2_R1269_U122, P2_R1269_U23);
  and ginst15262 (P2_R1269_U20, P2_R1269_U123, P2_R1269_U124, P2_R1269_U125);
  nand ginst15263 (P2_R1269_U200, P2_R1269_U121, P2_R1269_U14);
  nand ginst15264 (P2_R1269_U201, P2_R1269_U121, P2_R1269_U16);
  nand ginst15265 (P2_R1269_U202, P2_R1269_U121, P2_R1269_U17);
  nand ginst15266 (P2_R1269_U203, P2_R1269_U121, P2_R1269_U18);
  nand ginst15267 (P2_R1269_U204, P2_R1269_U121, P2_R1269_U19);
  nand ginst15268 (P2_R1269_U205, P2_U3084, P2_U3116);
  nand ginst15269 (P2_R1269_U206, P2_R1269_U25, P2_U3084);
  nand ginst15270 (P2_R1269_U207, P2_R1269_U24, P2_U3116);
  or ginst15271 (P2_R1269_U208, P2_U3116, P2_U3149);
  nand ginst15272 (P2_R1269_U209, P2_R1269_U24, P2_U3149);
  and ginst15273 (P2_R1269_U21, P2_R1269_U206, P2_R1269_U207);
  nand ginst15274 (P2_R1269_U22, P2_R1269_U119, P2_R1269_U120, P2_R1269_U127, P2_R1269_U200);
  not ginst15275 (P2_R1269_U23, P2_U3085);
  not ginst15276 (P2_R1269_U24, P2_U3084);
  not ginst15277 (P2_R1269_U25, P2_U3116);
  not ginst15278 (P2_R1269_U26, P2_U3118);
  not ginst15279 (P2_R1269_U27, P2_U3117);
  not ginst15280 (P2_R1269_U28, P2_U3086);
  not ginst15281 (P2_R1269_U29, P2_U3124);
  not ginst15282 (P2_R1269_U30, P2_U3123);
  not ginst15283 (P2_R1269_U31, P2_U3094);
  not ginst15284 (P2_R1269_U32, P2_U3127);
  not ginst15285 (P2_R1269_U33, P2_U3095);
  not ginst15286 (P2_R1269_U34, P2_U3128);
  not ginst15287 (P2_R1269_U35, P2_U3129);
  not ginst15288 (P2_R1269_U36, P2_U3098);
  not ginst15289 (P2_R1269_U37, P2_U3130);
  not ginst15290 (P2_R1269_U38, P2_U3099);
  not ginst15291 (P2_R1269_U39, P2_U3097);
  not ginst15292 (P2_R1269_U40, P2_U3096);
  not ginst15293 (P2_R1269_U41, P2_U3131);
  not ginst15294 (P2_R1269_U42, P2_U3132);
  not ginst15295 (P2_R1269_U43, P2_U3100);
  not ginst15296 (P2_R1269_U44, P2_U3101);
  not ginst15297 (P2_R1269_U45, P2_U3141);
  not ginst15298 (P2_R1269_U46, P2_U3110);
  not ginst15299 (P2_R1269_U47, P2_U3107);
  not ginst15300 (P2_R1269_U48, P2_U3106);
  not ginst15301 (P2_R1269_U49, P2_U3142);
  not ginst15302 (P2_R1269_U50, P2_U3111);
  not ginst15303 (P2_R1269_U51, P2_U3109);
  not ginst15304 (P2_R1269_U52, P2_U3108);
  not ginst15305 (P2_R1269_U53, P2_U3112);
  not ginst15306 (P2_R1269_U54, P2_U3113);
  not ginst15307 (P2_R1269_U55, P2_U3114);
  not ginst15308 (P2_R1269_U56, P2_U3136);
  not ginst15309 (P2_R1269_U57, P2_U3135);
  not ginst15310 (P2_R1269_U58, P2_U3139);
  not ginst15311 (P2_R1269_U59, P2_U3140);
  and ginst15312 (P2_R1269_U6, P2_R1269_U130, P2_R1269_U131);
  not ginst15313 (P2_R1269_U60, P2_U3146);
  not ginst15314 (P2_R1269_U61, P2_U3145);
  not ginst15315 (P2_R1269_U62, P2_U3143);
  not ginst15316 (P2_R1269_U63, P2_U3144);
  not ginst15317 (P2_R1269_U64, P2_U3138);
  not ginst15318 (P2_R1269_U65, P2_U3137);
  not ginst15319 (P2_R1269_U66, P2_U3104);
  not ginst15320 (P2_R1269_U67, P2_U3105);
  not ginst15321 (P2_R1269_U68, P2_U3102);
  not ginst15322 (P2_R1269_U69, P2_U3103);
  and ginst15323 (P2_R1269_U7, P2_R1269_U132, P2_R1269_U133);
  not ginst15324 (P2_R1269_U70, P2_U3134);
  not ginst15325 (P2_R1269_U71, P2_U3133);
  not ginst15326 (P2_R1269_U72, P2_U3126);
  not ginst15327 (P2_R1269_U73, P2_U3125);
  not ginst15328 (P2_R1269_U74, P2_U3093);
  not ginst15329 (P2_R1269_U75, P2_U3092);
  not ginst15330 (P2_R1269_U76, P2_U3090);
  not ginst15331 (P2_R1269_U77, P2_U3091);
  not ginst15332 (P2_R1269_U78, P2_U3087);
  not ginst15333 (P2_R1269_U79, P2_U3089);
  and ginst15334 (P2_R1269_U8, P2_R1269_U135, P2_R1269_U137, P2_R1269_U7, P2_R1269_U91);
  not ginst15335 (P2_R1269_U80, P2_U3088);
  not ginst15336 (P2_R1269_U81, P2_U3122);
  not ginst15337 (P2_R1269_U82, P2_U3121);
  not ginst15338 (P2_R1269_U83, P2_U3120);
  not ginst15339 (P2_R1269_U84, P2_U3119);
  and ginst15340 (P2_R1269_U85, P2_R1269_U28, P2_U3118);
  and ginst15341 (P2_R1269_U86, P2_R1269_U33, P2_U3127);
  and ginst15342 (P2_R1269_U87, P2_R1269_U40, P2_U3128);
  and ginst15343 (P2_R1269_U88, P2_R1269_U182, P2_R1269_U183);
  and ginst15344 (P2_R1269_U89, P2_R1269_U37, P2_U3098);
  and ginst15345 (P2_R1269_U9, P2_R1269_U144, P2_R1269_U145);
  and ginst15346 (P2_R1269_U90, P2_R1269_U41, P2_U3099);
  and ginst15347 (P2_R1269_U91, P2_R1269_U134, P2_R1269_U136);
  and ginst15348 (P2_R1269_U92, P2_R1269_U49, P2_U3110);
  and ginst15349 (P2_R1269_U93, P2_R1269_U62, P2_U3111);
  and ginst15350 (P2_R1269_U94, P2_R1269_U143, P2_R1269_U149);
  and ginst15351 (P2_R1269_U95, P2_R1269_U150, P2_R1269_U9);
  and ginst15352 (P2_R1269_U96, P2_R1269_U151, P2_R1269_U152);
  and ginst15353 (P2_R1269_U97, P2_R1269_U154, P2_R1269_U155, P2_R1269_U156);
  and ginst15354 (P2_R1269_U98, P2_R1269_U47, P2_U3139);
  and ginst15355 (P2_R1269_U99, P2_R1269_U52, P2_U3140);
  and ginst15356 (P2_R1297_U6, P2_R1297_U7, P2_U3058);
  not ginst15357 (P2_R1297_U7, P2_U3055);
  nand ginst15358 (P2_R1300_U10, P2_R1300_U7, P2_U3058);
  not ginst15359 (P2_R1300_U6, P2_U3058);
  not ginst15360 (P2_R1300_U7, P2_U3055);
  and ginst15361 (P2_R1300_U8, P2_R1300_U10, P2_R1300_U9);
  nand ginst15362 (P2_R1300_U9, P2_R1300_U6, P2_U3055);
  and ginst15363 (P2_R693_U10, P2_R693_U130, P2_R693_U132, P2_R693_U133, P2_R693_U134);
  and ginst15364 (P2_R693_U100, P2_R693_U187, P2_R693_U188);
  and ginst15365 (P2_R693_U101, P2_R693_U100, P2_R693_U6);
  and ginst15366 (P2_R693_U102, P2_R693_U103, P2_R693_U191);
  and ginst15367 (P2_R693_U103, P2_R693_U18, P2_U3533);
  and ginst15368 (P2_R693_U104, P2_R693_U114, P2_R693_U115, P2_R693_U116, P2_R693_U117);
  and ginst15369 (P2_R693_U105, P2_R693_U190, P2_R693_U192);
  not ginst15370 (P2_R693_U106, P2_U3869);
  not ginst15371 (P2_R693_U107, P2_U3554);
  nand ginst15372 (P2_R693_U108, P2_R693_U113, P2_R693_U193);
  nand ginst15373 (P2_R693_U109, P2_R693_U20, P2_U3904);
  and ginst15374 (P2_R693_U11, P2_R693_U10, P2_R693_U83);
  nand ginst15375 (P2_R693_U110, P2_R693_U21, P2_U3896);
  nand ginst15376 (P2_R693_U111, P2_R693_U74, P2_U3895);
  nand ginst15377 (P2_R693_U112, P2_R693_U73, P2_U3529);
  nand ginst15378 (P2_R693_U113, P2_R693_U106, P2_R693_U112);
  nand ginst15379 (P2_R693_U114, P2_R693_U108, P2_R693_U6, P2_R693_U72, P2_U3535);
  nand ginst15380 (P2_R693_U115, P2_R693_U106, P2_R693_U112, P2_U3530);
  nand ginst15381 (P2_R693_U116, P2_R693_U108, P2_R693_U75);
  nand ginst15382 (P2_R693_U117, P2_R693_U108, P2_R693_U17, P2_R693_U6, P2_U3534);
  nand ginst15383 (P2_R693_U118, P2_R693_U32, P2_U3543);
  nand ginst15384 (P2_R693_U119, P2_R693_U29, P2_U3544);
  and ginst15385 (P2_R693_U12, P2_R693_U11, P2_R693_U138);
  nand ginst15386 (P2_R693_U120, P2_R693_U67, P2_U3901);
  nand ginst15387 (P2_R693_U121, P2_R693_U25, P2_U3902);
  nand ginst15388 (P2_R693_U122, P2_R693_U118, P2_R693_U79);
  nand ginst15389 (P2_R693_U123, P2_R693_U7, P2_R693_U80);
  nand ginst15390 (P2_R693_U124, P2_R693_U28, P2_U3445);
  nand ginst15391 (P2_R693_U125, P2_R693_U27, P2_U3903);
  nand ginst15392 (P2_R693_U126, P2_R693_U35, P2_U3437);
  nand ginst15393 (P2_R693_U127, P2_R693_U70, P2_U3537);
  nand ginst15394 (P2_R693_U128, P2_R693_U71, P2_U3536);
  nand ginst15395 (P2_R693_U129, P2_R693_U66, P2_U3434);
  and ginst15396 (P2_R693_U13, P2_R693_U143, P2_R693_U144);
  nand ginst15397 (P2_R693_U130, P2_R693_U59, P2_U3419);
  nand ginst15398 (P2_R693_U131, P2_R693_U48, P2_U3553);
  nand ginst15399 (P2_R693_U132, P2_R693_U58, P2_U3416);
  nand ginst15400 (P2_R693_U133, P2_R693_U56, P2_U3410);
  nand ginst15401 (P2_R693_U134, P2_R693_U57, P2_U3413);
  nand ginst15402 (P2_R693_U135, P2_R693_U55, P2_U3407);
  nand ginst15403 (P2_R693_U136, P2_R693_U54, P2_U3404);
  nand ginst15404 (P2_R693_U137, P2_R693_U53, P2_U3401);
  nand ginst15405 (P2_R693_U138, P2_R693_U52, P2_U3398);
  nand ginst15406 (P2_R693_U139, P2_R693_U131, P2_R693_U82);
  and ginst15407 (P2_R693_U14, P2_R693_U104, P2_R693_U105, P2_R693_U189);
  nand ginst15408 (P2_R693_U140, P2_R693_U51, P2_U3395);
  nand ginst15409 (P2_R693_U141, P2_R693_U46, P2_U3392);
  nand ginst15410 (P2_R693_U142, P2_R693_U12, P2_R693_U85);
  nand ginst15411 (P2_R693_U143, P2_R693_U61, P2_U3550);
  nand ginst15412 (P2_R693_U144, P2_R693_U64, P2_U3549);
  nand ginst15413 (P2_R693_U145, P2_R693_U41, P2_U3524);
  nand ginst15414 (P2_R693_U146, P2_R693_U39, P2_U3523);
  nand ginst15415 (P2_R693_U147, P2_R693_U145, P2_R693_U146);
  nand ginst15416 (P2_R693_U148, P2_R693_U44, P2_U3528);
  nand ginst15417 (P2_R693_U149, P2_R693_U43, P2_U3527);
  not ginst15418 (P2_R693_U15, P2_U3529);
  nand ginst15419 (P2_R693_U150, P2_R693_U148, P2_R693_U149);
  nand ginst15420 (P2_R693_U151, P2_R693_U150, P2_R693_U88);
  nand ginst15421 (P2_R693_U152, P2_R693_U42, P2_U3526);
  nand ginst15422 (P2_R693_U153, P2_R693_U40, P2_U3525);
  nand ginst15423 (P2_R693_U154, P2_R693_U151, P2_R693_U89);
  nand ginst15424 (P2_R693_U155, P2_R693_U12, P2_R693_U86);
  nand ginst15425 (P2_R693_U156, P2_R693_U11, P2_R693_U87);
  nand ginst15426 (P2_R693_U157, P2_R693_U10, P2_R693_U154);
  nand ginst15427 (P2_R693_U158, P2_R693_U147, P2_R693_U90);
  nand ginst15428 (P2_R693_U159, P2_R693_U38, P2_U3552);
  not ginst15429 (P2_R693_U16, P2_U3904);
  nand ginst15430 (P2_R693_U160, P2_R693_U62, P2_U3551);
  nand ginst15431 (P2_R693_U161, P2_R693_U142, P2_R693_U155, P2_R693_U156, P2_R693_U157, P2_R693_U92);
  nand ginst15432 (P2_R693_U162, P2_R693_U64, P2_U3549);
  nand ginst15433 (P2_R693_U163, P2_R693_U162, P2_R693_U93);
  nand ginst15434 (P2_R693_U164, P2_R693_U13, P2_R693_U94);
  nand ginst15435 (P2_R693_U165, P2_R693_U65, P2_U3431);
  nand ginst15436 (P2_R693_U166, P2_R693_U50, P2_U3428);
  nand ginst15437 (P2_R693_U167, P2_R693_U161, P2_R693_U96);
  nand ginst15438 (P2_R693_U168, P2_R693_U63, P2_U3548);
  nand ginst15439 (P2_R693_U169, P2_R693_U167, P2_R693_U168);
  not ginst15440 (P2_R693_U17, P2_U3896);
  nand ginst15441 (P2_R693_U170, P2_R693_U129, P2_R693_U169);
  nand ginst15442 (P2_R693_U171, P2_R693_U37, P2_U3547);
  nand ginst15443 (P2_R693_U172, P2_R693_U170, P2_R693_U171);
  nand ginst15444 (P2_R693_U173, P2_R693_U31, P2_U3545);
  nand ginst15445 (P2_R693_U174, P2_R693_U36, P2_U3546);
  nand ginst15446 (P2_R693_U175, P2_R693_U7, P2_R693_U78);
  nand ginst15447 (P2_R693_U176, P2_R693_U120, P2_R693_U76);
  nand ginst15448 (P2_R693_U177, P2_R693_U77, P2_R693_U8);
  nand ginst15449 (P2_R693_U178, P2_R693_U175, P2_R693_U9);
  nand ginst15450 (P2_R693_U179, P2_R693_U126, P2_R693_U172, P2_R693_U9);
  not ginst15451 (P2_R693_U18, P2_U3895);
  nand ginst15452 (P2_R693_U180, P2_R693_U24, P2_U3539);
  nand ginst15453 (P2_R693_U181, P2_R693_U69, P2_U3538);
  nand ginst15454 (P2_R693_U182, P2_R693_U178, P2_R693_U179, P2_R693_U98, P2_R693_U99);
  nand ginst15455 (P2_R693_U183, P2_R693_U68, P2_U3900);
  nand ginst15456 (P2_R693_U184, P2_R693_U22, P2_U3899);
  nand ginst15457 (P2_R693_U185, P2_R693_U183, P2_R693_U184);
  nand ginst15458 (P2_R693_U186, P2_R693_U127, P2_R693_U128, P2_R693_U185);
  nand ginst15459 (P2_R693_U187, P2_R693_U23, P2_U3898);
  nand ginst15460 (P2_R693_U188, P2_R693_U19, P2_U3897);
  nand ginst15461 (P2_R693_U189, P2_R693_U101, P2_R693_U108, P2_R693_U182, P2_R693_U186);
  not ginst15462 (P2_R693_U19, P2_U3535);
  nand ginst15463 (P2_R693_U190, P2_R693_U15, P2_U3868);
  nand ginst15464 (P2_R693_U191, P2_R693_U20, P2_U3904);
  nand ginst15465 (P2_R693_U192, P2_R693_U102, P2_R693_U108);
  nand ginst15466 (P2_R693_U193, P2_R693_U112, P2_U3530);
  not ginst15467 (P2_R693_U20, P2_U3532);
  not ginst15468 (P2_R693_U21, P2_U3534);
  not ginst15469 (P2_R693_U22, P2_U3537);
  not ginst15470 (P2_R693_U23, P2_U3536);
  not ginst15471 (P2_R693_U24, P2_U3901);
  not ginst15472 (P2_R693_U25, P2_U3540);
  not ginst15473 (P2_R693_U26, P2_U3902);
  not ginst15474 (P2_R693_U27, P2_U3541);
  not ginst15475 (P2_R693_U28, P2_U3543);
  not ginst15476 (P2_R693_U29, P2_U3443);
  not ginst15477 (P2_R693_U30, P2_U3544);
  not ginst15478 (P2_R693_U31, P2_U3440);
  not ginst15479 (P2_R693_U32, P2_U3445);
  not ginst15480 (P2_R693_U33, P2_U3903);
  not ginst15481 (P2_R693_U34, P2_U3545);
  not ginst15482 (P2_R693_U35, P2_U3546);
  not ginst15483 (P2_R693_U36, P2_U3437);
  not ginst15484 (P2_R693_U37, P2_U3434);
  not ginst15485 (P2_R693_U38, P2_U3419);
  not ginst15486 (P2_R693_U39, P2_U3416);
  not ginst15487 (P2_R693_U40, P2_U3410);
  not ginst15488 (P2_R693_U41, P2_U3413);
  not ginst15489 (P2_R693_U42, P2_U3407);
  not ginst15490 (P2_R693_U43, P2_U3404);
  not ginst15491 (P2_R693_U44, P2_U3401);
  not ginst15492 (P2_R693_U45, P2_U3398);
  not ginst15493 (P2_R693_U46, P2_U3553);
  not ginst15494 (P2_R693_U47, P2_U3395);
  not ginst15495 (P2_R693_U48, P2_U3392);
  not ginst15496 (P2_R693_U49, P2_U3550);
  not ginst15497 (P2_R693_U50, P2_U3549);
  not ginst15498 (P2_R693_U51, P2_U3542);
  not ginst15499 (P2_R693_U52, P2_U3531);
  not ginst15500 (P2_R693_U53, P2_U3528);
  not ginst15501 (P2_R693_U54, P2_U3527);
  not ginst15502 (P2_R693_U55, P2_U3526);
  not ginst15503 (P2_R693_U56, P2_U3525);
  not ginst15504 (P2_R693_U57, P2_U3524);
  not ginst15505 (P2_R693_U58, P2_U3523);
  not ginst15506 (P2_R693_U59, P2_U3552);
  and ginst15507 (P2_R693_U6, P2_R693_U109, P2_R693_U110, P2_R693_U111);
  not ginst15508 (P2_R693_U60, P2_U3551);
  not ginst15509 (P2_R693_U61, P2_U3425);
  not ginst15510 (P2_R693_U62, P2_U3422);
  not ginst15511 (P2_R693_U63, P2_U3431);
  not ginst15512 (P2_R693_U64, P2_U3428);
  not ginst15513 (P2_R693_U65, P2_U3548);
  not ginst15514 (P2_R693_U66, P2_U3547);
  not ginst15515 (P2_R693_U67, P2_U3539);
  not ginst15516 (P2_R693_U68, P2_U3538);
  not ginst15517 (P2_R693_U69, P2_U3900);
  and ginst15518 (P2_R693_U7, P2_R693_U118, P2_R693_U119);
  not ginst15519 (P2_R693_U70, P2_U3899);
  not ginst15520 (P2_R693_U71, P2_U3898);
  not ginst15521 (P2_R693_U72, P2_U3897);
  not ginst15522 (P2_R693_U73, P2_U3868);
  not ginst15523 (P2_R693_U74, P2_U3533);
  and ginst15524 (P2_R693_U75, P2_R693_U16, P2_U3532);
  and ginst15525 (P2_R693_U76, P2_R693_U26, P2_U3540);
  and ginst15526 (P2_R693_U77, P2_R693_U33, P2_U3541);
  and ginst15527 (P2_R693_U78, P2_R693_U173, P2_R693_U174);
  and ginst15528 (P2_R693_U79, P2_R693_U30, P2_U3443);
  and ginst15529 (P2_R693_U8, P2_R693_U120, P2_R693_U121);
  and ginst15530 (P2_R693_U80, P2_R693_U34, P2_U3440);
  and ginst15531 (P2_R693_U81, P2_R693_U122, P2_R693_U124);
  and ginst15532 (P2_R693_U82, P2_R693_U107, P2_U3387);
  and ginst15533 (P2_R693_U83, P2_R693_U135, P2_R693_U136, P2_R693_U137);
  and ginst15534 (P2_R693_U84, P2_R693_U140, P2_R693_U141);
  and ginst15535 (P2_R693_U85, P2_R693_U139, P2_R693_U84);
  and ginst15536 (P2_R693_U86, P2_R693_U47, P2_U3542);
  and ginst15537 (P2_R693_U87, P2_R693_U45, P2_U3531);
  and ginst15538 (P2_R693_U88, P2_R693_U135, P2_R693_U136);
  and ginst15539 (P2_R693_U89, P2_R693_U152, P2_R693_U153);
  and ginst15540 (P2_R693_U9, P2_R693_U123, P2_R693_U125, P2_R693_U8, P2_R693_U81);
  and ginst15541 (P2_R693_U90, P2_R693_U130, P2_R693_U132);
  and ginst15542 (P2_R693_U91, P2_R693_U13, P2_R693_U160);
  and ginst15543 (P2_R693_U92, P2_R693_U158, P2_R693_U159, P2_R693_U91);
  and ginst15544 (P2_R693_U93, P2_R693_U49, P2_U3425);
  and ginst15545 (P2_R693_U94, P2_R693_U60, P2_U3422);
  and ginst15546 (P2_R693_U95, P2_R693_U163, P2_R693_U97);
  and ginst15547 (P2_R693_U96, P2_R693_U164, P2_R693_U95);
  and ginst15548 (P2_R693_U97, P2_R693_U165, P2_R693_U166);
  and ginst15549 (P2_R693_U98, P2_R693_U127, P2_R693_U128, P2_R693_U176, P2_R693_U177);
  and ginst15550 (P2_R693_U99, P2_R693_U180, P2_R693_U181);
  and ginst15551 (P2_SUB_594_U10, P2_SUB_594_U132, P2_SUB_594_U47);
  not ginst15552 (P2_SUB_594_U100, P2_SUB_594_U51);
  nand ginst15553 (P2_SUB_594_U101, P2_SUB_594_U100, P2_SUB_594_U52);
  not ginst15554 (P2_SUB_594_U102, P2_SUB_594_U47);
  not ginst15555 (P2_SUB_594_U103, P2_SUB_594_U48);
  nand ginst15556 (P2_SUB_594_U104, P2_SUB_594_U103, P2_SUB_594_U50);
  not ginst15557 (P2_SUB_594_U105, P2_SUB_594_U35);
  not ginst15558 (P2_SUB_594_U106, P2_SUB_594_U45);
  nand ginst15559 (P2_SUB_594_U107, P2_SUB_594_U106, P2_SUB_594_U46);
  not ginst15560 (P2_SUB_594_U108, P2_SUB_594_U41);
  not ginst15561 (P2_SUB_594_U109, P2_SUB_594_U42);
  and ginst15562 (P2_SUB_594_U11, P2_SUB_594_U131, P2_SUB_594_U48);
  nand ginst15563 (P2_SUB_594_U110, P2_SUB_594_U109, P2_SUB_594_U44);
  not ginst15564 (P2_SUB_594_U111, P2_SUB_594_U36);
  not ginst15565 (P2_SUB_594_U112, P2_SUB_594_U76);
  not ginst15566 (P2_SUB_594_U113, P2_SUB_594_U37);
  not ginst15567 (P2_SUB_594_U114, P2_SUB_594_U38);
  or ginst15568 (P2_SUB_594_U115, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN);
  nand ginst15569 (P2_SUB_594_U116, P2_IR_REG_2__SCAN_IN, P2_SUB_594_U115);
  nand ginst15570 (P2_SUB_594_U117, P2_IR_REG_29__SCAN_IN, P2_SUB_594_U37);
  nand ginst15571 (P2_SUB_594_U118, P2_SUB_594_U111, P2_SUB_594_U78);
  nand ginst15572 (P2_SUB_594_U119, P2_IR_REG_26__SCAN_IN, P2_SUB_594_U118);
  and ginst15573 (P2_SUB_594_U12, P2_SUB_594_U104, P2_SUB_594_U129);
  nand ginst15574 (P2_SUB_594_U120, P2_IR_REG_24__SCAN_IN, P2_SUB_594_U110);
  nand ginst15575 (P2_SUB_594_U121, P2_IR_REG_23__SCAN_IN, P2_SUB_594_U42);
  nand ginst15576 (P2_SUB_594_U122, P2_SUB_594_U108, P2_SUB_594_U80);
  nand ginst15577 (P2_SUB_594_U123, P2_IR_REG_22__SCAN_IN, P2_SUB_594_U122);
  nand ginst15578 (P2_SUB_594_U124, P2_IR_REG_20__SCAN_IN, P2_SUB_594_U107);
  nand ginst15579 (P2_SUB_594_U125, P2_IR_REG_19__SCAN_IN, P2_SUB_594_U45);
  nand ginst15580 (P2_SUB_594_U126, P2_SUB_594_U105, P2_SUB_594_U84);
  nand ginst15581 (P2_SUB_594_U127, P2_IR_REG_18__SCAN_IN, P2_SUB_594_U126);
  nand ginst15582 (P2_SUB_594_U128, P2_IR_REG_16__SCAN_IN, P2_SUB_594_U104);
  nand ginst15583 (P2_SUB_594_U129, P2_IR_REG_15__SCAN_IN, P2_SUB_594_U48);
  and ginst15584 (P2_SUB_594_U13, P2_SUB_594_U128, P2_SUB_594_U35);
  nand ginst15585 (P2_SUB_594_U130, P2_SUB_594_U102, P2_SUB_594_U86);
  nand ginst15586 (P2_SUB_594_U131, P2_IR_REG_14__SCAN_IN, P2_SUB_594_U130);
  nand ginst15587 (P2_SUB_594_U132, P2_IR_REG_12__SCAN_IN, P2_SUB_594_U101);
  nand ginst15588 (P2_SUB_594_U133, P2_IR_REG_11__SCAN_IN, P2_SUB_594_U51);
  nand ginst15589 (P2_SUB_594_U134, P2_SUB_594_U69, P2_SUB_594_U93);
  nand ginst15590 (P2_SUB_594_U135, P2_IR_REG_10__SCAN_IN, P2_SUB_594_U134);
  nand ginst15591 (P2_SUB_594_U136, P2_SUB_594_U114, P2_SUB_594_U74);
  nand ginst15592 (P2_SUB_594_U137, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN);
  nand ginst15593 (P2_SUB_594_U138, P2_IR_REG_28__SCAN_IN, P2_SUB_594_U76);
  nand ginst15594 (P2_SUB_594_U139, P2_IR_REG_9__SCAN_IN, P2_SUB_594_U29);
  and ginst15595 (P2_SUB_594_U14, P2_SUB_594_U127, P2_SUB_594_U45);
  nand ginst15596 (P2_SUB_594_U140, P2_SUB_594_U69, P2_SUB_594_U93);
  nand ginst15597 (P2_SUB_594_U141, P2_IR_REG_5__SCAN_IN, P2_SUB_594_U30);
  nand ginst15598 (P2_SUB_594_U142, P2_SUB_594_U71, P2_SUB_594_U90);
  nand ginst15599 (P2_SUB_594_U143, P2_SUB_594_U136, P2_SUB_594_U73);
  nand ginst15600 (P2_SUB_594_U144, P2_IR_REG_31__SCAN_IN, P2_SUB_594_U114, P2_SUB_594_U74);
  nand ginst15601 (P2_SUB_594_U145, P2_IR_REG_30__SCAN_IN, P2_SUB_594_U38);
  nand ginst15602 (P2_SUB_594_U146, P2_SUB_594_U114, P2_SUB_594_U74);
  nand ginst15603 (P2_SUB_594_U147, P2_IR_REG_27__SCAN_IN, P2_SUB_594_U76);
  nand ginst15604 (P2_SUB_594_U148, P2_SUB_594_U112, P2_SUB_594_U40);
  nand ginst15605 (P2_SUB_594_U149, P2_IR_REG_25__SCAN_IN, P2_SUB_594_U36);
  and ginst15606 (P2_SUB_594_U15, P2_SUB_594_U107, P2_SUB_594_U125);
  nand ginst15607 (P2_SUB_594_U150, P2_SUB_594_U111, P2_SUB_594_U78);
  nand ginst15608 (P2_SUB_594_U151, P2_IR_REG_21__SCAN_IN, P2_SUB_594_U41);
  nand ginst15609 (P2_SUB_594_U152, P2_SUB_594_U108, P2_SUB_594_U80);
  nand ginst15610 (P2_SUB_594_U153, P2_IR_REG_1__SCAN_IN, P2_SUB_594_U83);
  nand ginst15611 (P2_SUB_594_U154, P2_IR_REG_0__SCAN_IN, P2_SUB_594_U82);
  nand ginst15612 (P2_SUB_594_U155, P2_IR_REG_17__SCAN_IN, P2_SUB_594_U35);
  nand ginst15613 (P2_SUB_594_U156, P2_SUB_594_U105, P2_SUB_594_U84);
  nand ginst15614 (P2_SUB_594_U157, P2_IR_REG_13__SCAN_IN, P2_SUB_594_U47);
  nand ginst15615 (P2_SUB_594_U158, P2_SUB_594_U102, P2_SUB_594_U86);
  and ginst15616 (P2_SUB_594_U16, P2_SUB_594_U124, P2_SUB_594_U41);
  and ginst15617 (P2_SUB_594_U17, P2_SUB_594_U123, P2_SUB_594_U42);
  and ginst15618 (P2_SUB_594_U18, P2_SUB_594_U110, P2_SUB_594_U121);
  and ginst15619 (P2_SUB_594_U19, P2_SUB_594_U120, P2_SUB_594_U36);
  and ginst15620 (P2_SUB_594_U20, P2_SUB_594_U119, P2_SUB_594_U76);
  and ginst15621 (P2_SUB_594_U21, P2_SUB_594_U138, P2_SUB_594_U64);
  and ginst15622 (P2_SUB_594_U22, P2_SUB_594_U117, P2_SUB_594_U38);
  and ginst15623 (P2_SUB_594_U23, P2_SUB_594_U116, P2_SUB_594_U33);
  and ginst15624 (P2_SUB_594_U24, P2_SUB_594_U89, P2_SUB_594_U99);
  and ginst15625 (P2_SUB_594_U25, P2_SUB_594_U30, P2_SUB_594_U98);
  and ginst15626 (P2_SUB_594_U26, P2_SUB_594_U31, P2_SUB_594_U97);
  and ginst15627 (P2_SUB_594_U27, P2_SUB_594_U92, P2_SUB_594_U95);
  and ginst15628 (P2_SUB_594_U28, P2_SUB_594_U29, P2_SUB_594_U94);
  nand ginst15629 (P2_SUB_594_U29, P2_SUB_594_U55, P2_SUB_594_U56);
  or ginst15630 (P2_SUB_594_U30, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN, P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN);
  nand ginst15631 (P2_SUB_594_U31, P2_SUB_594_U57, P2_SUB_594_U90);
  not ginst15632 (P2_SUB_594_U32, P2_IR_REG_7__SCAN_IN);
  or ginst15633 (P2_SUB_594_U33, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN, P2_IR_REG_2__SCAN_IN);
  not ginst15634 (P2_SUB_594_U34, P2_IR_REG_3__SCAN_IN);
  nand ginst15635 (P2_SUB_594_U35, P2_SUB_594_U59, P2_SUB_594_U93);
  nand ginst15636 (P2_SUB_594_U36, P2_SUB_594_U105, P2_SUB_594_U61);
  nand ginst15637 (P2_SUB_594_U37, P2_SUB_594_U111, P2_SUB_594_U62);
  nand ginst15638 (P2_SUB_594_U38, P2_SUB_594_U113, P2_SUB_594_U39);
  not ginst15639 (P2_SUB_594_U39, P2_IR_REG_29__SCAN_IN);
  not ginst15640 (P2_SUB_594_U40, P2_IR_REG_27__SCAN_IN);
  nand ginst15641 (P2_SUB_594_U41, P2_SUB_594_U105, P2_SUB_594_U7);
  nand ginst15642 (P2_SUB_594_U42, P2_SUB_594_U108, P2_SUB_594_U65);
  not ginst15643 (P2_SUB_594_U43, P2_IR_REG_24__SCAN_IN);
  not ginst15644 (P2_SUB_594_U44, P2_IR_REG_23__SCAN_IN);
  nand ginst15645 (P2_SUB_594_U45, P2_SUB_594_U105, P2_SUB_594_U66);
  not ginst15646 (P2_SUB_594_U46, P2_IR_REG_19__SCAN_IN);
  nand ginst15647 (P2_SUB_594_U47, P2_SUB_594_U6, P2_SUB_594_U93);
  nand ginst15648 (P2_SUB_594_U48, P2_SUB_594_U102, P2_SUB_594_U67);
  not ginst15649 (P2_SUB_594_U49, P2_IR_REG_16__SCAN_IN);
  not ginst15650 (P2_SUB_594_U50, P2_IR_REG_15__SCAN_IN);
  nand ginst15651 (P2_SUB_594_U51, P2_SUB_594_U68, P2_SUB_594_U93);
  not ginst15652 (P2_SUB_594_U52, P2_IR_REG_11__SCAN_IN);
  nand ginst15653 (P2_SUB_594_U53, P2_SUB_594_U153, P2_SUB_594_U154);
  nand ginst15654 (P2_SUB_594_U54, P2_SUB_594_U143, P2_SUB_594_U144);
  nor ginst15655 (P2_SUB_594_U55, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN, P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN);
  nor ginst15656 (P2_SUB_594_U56, P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN, P2_IR_REG_8__SCAN_IN);
  nor ginst15657 (P2_SUB_594_U57, P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN);
  nor ginst15658 (P2_SUB_594_U58, P2_IR_REG_13__SCAN_IN, P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN);
  and ginst15659 (P2_SUB_594_U59, P2_SUB_594_U49, P2_SUB_594_U58, P2_SUB_594_U6);
  nor ginst15660 (P2_SUB_594_U6, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN, P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN);
  nor ginst15661 (P2_SUB_594_U60, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN, P2_IR_REG_23__SCAN_IN);
  and ginst15662 (P2_SUB_594_U61, P2_SUB_594_U43, P2_SUB_594_U60, P2_SUB_594_U7);
  nor ginst15663 (P2_SUB_594_U62, P2_IR_REG_25__SCAN_IN, P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN);
  nor ginst15664 (P2_SUB_594_U63, P2_IR_REG_25__SCAN_IN, P2_IR_REG_26__SCAN_IN);
  and ginst15665 (P2_SUB_594_U64, P2_SUB_594_U137, P2_SUB_594_U37);
  nor ginst15666 (P2_SUB_594_U65, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN);
  nor ginst15667 (P2_SUB_594_U66, P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN);
  nor ginst15668 (P2_SUB_594_U67, P2_IR_REG_13__SCAN_IN, P2_IR_REG_14__SCAN_IN);
  nor ginst15669 (P2_SUB_594_U68, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN);
  not ginst15670 (P2_SUB_594_U69, P2_IR_REG_9__SCAN_IN);
  nor ginst15671 (P2_SUB_594_U7, P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN, P2_IR_REG_20__SCAN_IN);
  and ginst15672 (P2_SUB_594_U70, P2_SUB_594_U139, P2_SUB_594_U140);
  not ginst15673 (P2_SUB_594_U71, P2_IR_REG_5__SCAN_IN);
  and ginst15674 (P2_SUB_594_U72, P2_SUB_594_U141, P2_SUB_594_U142);
  not ginst15675 (P2_SUB_594_U73, P2_IR_REG_31__SCAN_IN);
  not ginst15676 (P2_SUB_594_U74, P2_IR_REG_30__SCAN_IN);
  and ginst15677 (P2_SUB_594_U75, P2_SUB_594_U145, P2_SUB_594_U146);
  nand ginst15678 (P2_SUB_594_U76, P2_SUB_594_U111, P2_SUB_594_U63);
  and ginst15679 (P2_SUB_594_U77, P2_SUB_594_U147, P2_SUB_594_U148);
  not ginst15680 (P2_SUB_594_U78, P2_IR_REG_25__SCAN_IN);
  and ginst15681 (P2_SUB_594_U79, P2_SUB_594_U149, P2_SUB_594_U150);
  and ginst15682 (P2_SUB_594_U8, P2_SUB_594_U135, P2_SUB_594_U51);
  not ginst15683 (P2_SUB_594_U80, P2_IR_REG_21__SCAN_IN);
  and ginst15684 (P2_SUB_594_U81, P2_SUB_594_U151, P2_SUB_594_U152);
  not ginst15685 (P2_SUB_594_U82, P2_IR_REG_1__SCAN_IN);
  not ginst15686 (P2_SUB_594_U83, P2_IR_REG_0__SCAN_IN);
  not ginst15687 (P2_SUB_594_U84, P2_IR_REG_17__SCAN_IN);
  and ginst15688 (P2_SUB_594_U85, P2_SUB_594_U155, P2_SUB_594_U156);
  not ginst15689 (P2_SUB_594_U86, P2_IR_REG_13__SCAN_IN);
  and ginst15690 (P2_SUB_594_U87, P2_SUB_594_U157, P2_SUB_594_U158);
  not ginst15691 (P2_SUB_594_U88, P2_SUB_594_U33);
  nand ginst15692 (P2_SUB_594_U89, P2_SUB_594_U34, P2_SUB_594_U88);
  and ginst15693 (P2_SUB_594_U9, P2_SUB_594_U101, P2_SUB_594_U133);
  not ginst15694 (P2_SUB_594_U90, P2_SUB_594_U30);
  not ginst15695 (P2_SUB_594_U91, P2_SUB_594_U31);
  nand ginst15696 (P2_SUB_594_U92, P2_SUB_594_U32, P2_SUB_594_U91);
  not ginst15697 (P2_SUB_594_U93, P2_SUB_594_U29);
  nand ginst15698 (P2_SUB_594_U94, P2_IR_REG_8__SCAN_IN, P2_SUB_594_U92);
  nand ginst15699 (P2_SUB_594_U95, P2_IR_REG_7__SCAN_IN, P2_SUB_594_U31);
  nand ginst15700 (P2_SUB_594_U96, P2_SUB_594_U71, P2_SUB_594_U90);
  nand ginst15701 (P2_SUB_594_U97, P2_IR_REG_6__SCAN_IN, P2_SUB_594_U96);
  nand ginst15702 (P2_SUB_594_U98, P2_IR_REG_4__SCAN_IN, P2_SUB_594_U89);
  nand ginst15703 (P2_SUB_594_U99, P2_IR_REG_3__SCAN_IN, P2_SUB_594_U33);
  nand ginst15704 (P2_SUB_605_U10, P2_SUB_605_U89, P2_SUB_605_U99);
  nand ginst15705 (P2_SUB_605_U100, P2_REG3_REG_23__SCAN_IN, P2_SUB_605_U87);
  nand ginst15706 (P2_SUB_605_U101, P2_REG3_REG_22__SCAN_IN, P2_SUB_605_U38);
  nand ginst15707 (P2_SUB_605_U102, P2_REG3_REG_21__SCAN_IN, P2_SUB_605_U85);
  nand ginst15708 (P2_SUB_605_U103, P2_REG3_REG_20__SCAN_IN, P2_SUB_605_U37);
  nand ginst15709 (P2_SUB_605_U104, P2_REG3_REG_19__SCAN_IN, P2_SUB_605_U83);
  nand ginst15710 (P2_SUB_605_U105, P2_REG3_REG_18__SCAN_IN, P2_SUB_605_U36);
  nand ginst15711 (P2_SUB_605_U106, P2_REG3_REG_17__SCAN_IN, P2_SUB_605_U81);
  nand ginst15712 (P2_SUB_605_U107, P2_REG3_REG_16__SCAN_IN, P2_SUB_605_U35);
  nand ginst15713 (P2_SUB_605_U108, P2_REG3_REG_15__SCAN_IN, P2_SUB_605_U79);
  nand ginst15714 (P2_SUB_605_U109, P2_REG3_REG_14__SCAN_IN, P2_SUB_605_U49);
  nand ginst15715 (P2_SUB_605_U11, P2_SUB_605_U105, P2_SUB_605_U83);
  nand ginst15716 (P2_SUB_605_U110, P2_REG3_REG_13__SCAN_IN, P2_SUB_605_U77);
  nand ginst15717 (P2_SUB_605_U111, P2_REG3_REG_12__SCAN_IN, P2_SUB_605_U34);
  nand ginst15718 (P2_SUB_605_U112, P2_REG3_REG_11__SCAN_IN, P2_SUB_605_U75);
  nand ginst15719 (P2_SUB_605_U113, P2_REG3_REG_10__SCAN_IN, P2_SUB_605_U68);
  nand ginst15720 (P2_SUB_605_U12, P2_SUB_605_U67, P2_SUB_605_U70);
  nand ginst15721 (P2_SUB_605_U13, P2_SUB_605_U113, P2_SUB_605_U75);
  nand ginst15722 (P2_SUB_605_U14, P2_SUB_605_U68, P2_SUB_605_U69);
  nand ginst15723 (P2_SUB_605_U15, P2_SUB_605_U104, P2_SUB_605_U37);
  nand ginst15724 (P2_SUB_605_U16, P2_SUB_605_U40, P2_SUB_605_U98);
  nand ginst15725 (P2_SUB_605_U17, P2_SUB_605_U101, P2_SUB_605_U87);
  nand ginst15726 (P2_SUB_605_U18, P2_SUB_605_U32, P2_SUB_605_U71);
  nand ginst15727 (P2_SUB_605_U19, P2_SUB_605_U106, P2_SUB_605_U36);
  nand ginst15728 (P2_SUB_605_U20, P2_SUB_605_U103, P2_SUB_605_U85);
  nand ginst15729 (P2_SUB_605_U21, P2_SUB_605_U108, P2_SUB_605_U35);
  nand ginst15730 (P2_SUB_605_U22, P2_SUB_605_U64, P2_SUB_605_U73);
  nand ginst15731 (P2_SUB_605_U23, P2_SUB_605_U41, P2_SUB_605_U96);
  nand ginst15732 (P2_SUB_605_U24, P2_SUB_605_U111, P2_SUB_605_U77);
  nand ginst15733 (P2_SUB_605_U25, P2_SUB_605_U110, P2_SUB_605_U49);
  not ginst15734 (P2_SUB_605_U26, P2_REG3_REG_3__SCAN_IN);
  nand ginst15735 (P2_SUB_605_U27, P2_SUB_605_U91, P2_SUB_605_U97);
  nand ginst15736 (P2_SUB_605_U28, P2_SUB_605_U102, P2_SUB_605_U38);
  nand ginst15737 (P2_SUB_605_U29, P2_SUB_605_U93, P2_SUB_605_U95);
  nand ginst15738 (P2_SUB_605_U30, P2_SUB_605_U63, P2_SUB_605_U74);
  nand ginst15739 (P2_SUB_605_U31, P2_SUB_605_U109, P2_SUB_605_U79);
  or ginst15740 (P2_SUB_605_U32, P2_REG3_REG_7__SCAN_IN, P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_5__SCAN_IN, P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_6__SCAN_IN);
  not ginst15741 (P2_SUB_605_U33, P2_REG3_REG_8__SCAN_IN);
  nand ginst15742 (P2_SUB_605_U34, P2_SUB_605_U53, P2_SUB_605_U66);
  nand ginst15743 (P2_SUB_605_U35, P2_SUB_605_U54, P2_SUB_605_U76);
  nand ginst15744 (P2_SUB_605_U36, P2_SUB_605_U55, P2_SUB_605_U80);
  nand ginst15745 (P2_SUB_605_U37, P2_SUB_605_U56, P2_SUB_605_U82);
  nand ginst15746 (P2_SUB_605_U38, P2_SUB_605_U57, P2_SUB_605_U84);
  nand ginst15747 (P2_SUB_605_U39, P2_SUB_605_U58, P2_SUB_605_U86);
  nand ginst15748 (P2_SUB_605_U40, P2_SUB_605_U59, P2_SUB_605_U88);
  nand ginst15749 (P2_SUB_605_U41, P2_SUB_605_U60, P2_SUB_605_U90);
  not ginst15750 (P2_SUB_605_U42, P2_REG3_REG_28__SCAN_IN);
  not ginst15751 (P2_SUB_605_U43, P2_REG3_REG_26__SCAN_IN);
  not ginst15752 (P2_SUB_605_U44, P2_REG3_REG_24__SCAN_IN);
  not ginst15753 (P2_SUB_605_U45, P2_REG3_REG_22__SCAN_IN);
  not ginst15754 (P2_SUB_605_U46, P2_REG3_REG_20__SCAN_IN);
  not ginst15755 (P2_SUB_605_U47, P2_REG3_REG_18__SCAN_IN);
  not ginst15756 (P2_SUB_605_U48, P2_REG3_REG_16__SCAN_IN);
  nand ginst15757 (P2_SUB_605_U49, P2_SUB_605_U61, P2_SUB_605_U76);
  not ginst15758 (P2_SUB_605_U50, P2_REG3_REG_14__SCAN_IN);
  not ginst15759 (P2_SUB_605_U51, P2_REG3_REG_12__SCAN_IN);
  nor ginst15760 (P2_SUB_605_U52, P2_REG3_REG_8__SCAN_IN, P2_REG3_REG_9__SCAN_IN);
  nor ginst15761 (P2_SUB_605_U53, P2_REG3_REG_10__SCAN_IN, P2_REG3_REG_8__SCAN_IN, P2_REG3_REG_9__SCAN_IN, P2_REG3_REG_11__SCAN_IN);
  nor ginst15762 (P2_SUB_605_U54, P2_REG3_REG_14__SCAN_IN, P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_13__SCAN_IN, P2_REG3_REG_15__SCAN_IN);
  nor ginst15763 (P2_SUB_605_U55, P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_17__SCAN_IN);
  nor ginst15764 (P2_SUB_605_U56, P2_REG3_REG_19__SCAN_IN, P2_REG3_REG_18__SCAN_IN);
  nor ginst15765 (P2_SUB_605_U57, P2_REG3_REG_21__SCAN_IN, P2_REG3_REG_20__SCAN_IN);
  nor ginst15766 (P2_SUB_605_U58, P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_22__SCAN_IN);
  nor ginst15767 (P2_SUB_605_U59, P2_REG3_REG_25__SCAN_IN, P2_REG3_REG_24__SCAN_IN);
  nand ginst15768 (P2_SUB_605_U6, P2_SUB_605_U100, P2_SUB_605_U39);
  nor ginst15769 (P2_SUB_605_U60, P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_26__SCAN_IN);
  nor ginst15770 (P2_SUB_605_U61, P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_13__SCAN_IN);
  nor ginst15771 (P2_SUB_605_U62, P2_REG3_REG_10__SCAN_IN, P2_REG3_REG_8__SCAN_IN, P2_REG3_REG_9__SCAN_IN);
  or ginst15772 (P2_SUB_605_U63, P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_4__SCAN_IN);
  or ginst15773 (P2_SUB_605_U64, P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_5__SCAN_IN, P2_REG3_REG_4__SCAN_IN);
  or ginst15774 (P2_SUB_605_U65, P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_5__SCAN_IN, P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_6__SCAN_IN);
  not ginst15775 (P2_SUB_605_U66, P2_SUB_605_U32);
  nand ginst15776 (P2_SUB_605_U67, P2_SUB_605_U33, P2_SUB_605_U66);
  nand ginst15777 (P2_SUB_605_U68, P2_SUB_605_U52, P2_SUB_605_U66);
  nand ginst15778 (P2_SUB_605_U69, P2_REG3_REG_9__SCAN_IN, P2_SUB_605_U67);
  nand ginst15779 (P2_SUB_605_U7, P2_SUB_605_U107, P2_SUB_605_U81);
  nand ginst15780 (P2_SUB_605_U70, P2_REG3_REG_8__SCAN_IN, P2_SUB_605_U32);
  nand ginst15781 (P2_SUB_605_U71, P2_REG3_REG_7__SCAN_IN, P2_SUB_605_U65);
  nand ginst15782 (P2_SUB_605_U72, P2_REG3_REG_6__SCAN_IN, P2_SUB_605_U64);
  nand ginst15783 (P2_SUB_605_U73, P2_REG3_REG_5__SCAN_IN, P2_SUB_605_U63);
  nand ginst15784 (P2_SUB_605_U74, P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_4__SCAN_IN);
  nand ginst15785 (P2_SUB_605_U75, P2_SUB_605_U62, P2_SUB_605_U66);
  not ginst15786 (P2_SUB_605_U76, P2_SUB_605_U34);
  nand ginst15787 (P2_SUB_605_U77, P2_SUB_605_U51, P2_SUB_605_U76);
  not ginst15788 (P2_SUB_605_U78, P2_SUB_605_U49);
  nand ginst15789 (P2_SUB_605_U79, P2_SUB_605_U50, P2_SUB_605_U78);
  nand ginst15790 (P2_SUB_605_U8, P2_SUB_605_U65, P2_SUB_605_U72);
  not ginst15791 (P2_SUB_605_U80, P2_SUB_605_U35);
  nand ginst15792 (P2_SUB_605_U81, P2_SUB_605_U48, P2_SUB_605_U80);
  not ginst15793 (P2_SUB_605_U82, P2_SUB_605_U36);
  nand ginst15794 (P2_SUB_605_U83, P2_SUB_605_U47, P2_SUB_605_U82);
  not ginst15795 (P2_SUB_605_U84, P2_SUB_605_U37);
  nand ginst15796 (P2_SUB_605_U85, P2_SUB_605_U46, P2_SUB_605_U84);
  not ginst15797 (P2_SUB_605_U86, P2_SUB_605_U38);
  nand ginst15798 (P2_SUB_605_U87, P2_SUB_605_U45, P2_SUB_605_U86);
  not ginst15799 (P2_SUB_605_U88, P2_SUB_605_U39);
  nand ginst15800 (P2_SUB_605_U89, P2_SUB_605_U44, P2_SUB_605_U88);
  nand ginst15801 (P2_SUB_605_U9, P2_SUB_605_U112, P2_SUB_605_U34);
  not ginst15802 (P2_SUB_605_U90, P2_SUB_605_U40);
  nand ginst15803 (P2_SUB_605_U91, P2_SUB_605_U43, P2_SUB_605_U90);
  not ginst15804 (P2_SUB_605_U92, P2_SUB_605_U41);
  nand ginst15805 (P2_SUB_605_U93, P2_SUB_605_U42, P2_SUB_605_U92);
  not ginst15806 (P2_SUB_605_U94, P2_SUB_605_U93);
  nand ginst15807 (P2_SUB_605_U95, P2_REG3_REG_28__SCAN_IN, P2_SUB_605_U41);
  nand ginst15808 (P2_SUB_605_U96, P2_REG3_REG_27__SCAN_IN, P2_SUB_605_U91);
  nand ginst15809 (P2_SUB_605_U97, P2_REG3_REG_26__SCAN_IN, P2_SUB_605_U40);
  nand ginst15810 (P2_SUB_605_U98, P2_REG3_REG_25__SCAN_IN, P2_SUB_605_U89);
  nand ginst15811 (P2_SUB_605_U99, P2_REG3_REG_24__SCAN_IN, P2_SUB_605_U39);
  and ginst15812 (P2_U3013, P2_U3380, P2_U5446);
  and ginst15813 (P2_U3014, P2_U3379, P2_U3380);
  and ginst15814 (P2_U3015, P2_U3379, P2_U5449);
  and ginst15815 (P2_U3016, P2_U5446, P2_U5449);
  and ginst15816 (P2_U3017, P2_U3870, P2_U5443);
  and ginst15817 (P2_U3018, P2_U3582, P2_U3587);
  and ginst15818 (P2_U3019, P2_U3381, P2_U3382);
  and ginst15819 (P2_U3020, P2_U3381, P2_U5458);
  and ginst15820 (P2_U3021, P2_U3382, P2_U5455);
  and ginst15821 (P2_U3022, P2_U5455, P2_U5458);
  and ginst15822 (P2_U3023, P2_STATE_REG_SCAN_IN, P2_U3046);
  and ginst15823 (P2_U3024, P2_U3366, P2_U3701);
  and ginst15824 (P2_U3025, P2_U3907, P2_U4069);
  and ginst15825 (P2_U3026, P2_U3015, P2_U5443);
  and ginst15826 (P2_U3027, P2_STATE_REG_SCAN_IN, P2_U3297);
  and ginst15827 (P2_U3028, P2_U3882, P2_U3908);
  and ginst15828 (P2_U3029, P2_U3365, P2_U3908);
  and ginst15829 (P2_U3030, P2_U3698, P2_U3908);
  and ginst15830 (P2_U3031, P2_U3023, P2_U3886);
  and ginst15831 (P2_U3032, P2_U3891, P2_U4069);
  and ginst15832 (P2_U3033, P2_U3907, P2_U4085);
  and ginst15833 (P2_U3034, P2_U3025, P2_U3908);
  and ginst15834 (P2_U3035, P2_U3023, P2_U4985);
  and ginst15835 (P2_U3036, P2_U3891, P2_U4085);
  and ginst15836 (P2_U3037, P2_U4750, P2_U5464);
  and ginst15837 (P2_U3038, P2_U3024, P2_U5464);
  and ginst15838 (P2_U3039, P2_U4750, P2_U5461);
  and ginst15839 (P2_U3040, P2_U3888, P2_U4750);
  and ginst15840 (P2_U3041, P2_U3024, P2_U3888);
  and ginst15841 (P2_U3042, P2_U3023, P2_U3366);
  and ginst15842 (P2_U3043, P2_U3023, P2_U3365);
  and ginst15843 (P2_U3044, P2_STATE_REG_SCAN_IN, P2_U5000);
  and ginst15844 (P2_U3045, P2_U3023, P2_U5002);
  and ginst15845 (P2_U3046, P2_U3362, P2_U5436);
  and ginst15846 (P2_U3047, P2_U3018, P2_U3697);
  and ginst15847 (P2_U3048, P2_U3018, P2_U3696);
  and ginst15848 (P2_U3049, P2_U4744, P2_U4745);
  and ginst15849 (P2_U3050, P2_STATE_REG_SCAN_IN, P2_U4755);
  and ginst15850 (P2_U3051, P2_U3893, P2_U4757);
  nand ginst15851 (P2_U3052, P2_U4531, P2_U4532, P2_U4533, P2_U4534);
  nand ginst15852 (P2_U3053, P2_U4549, P2_U4550, P2_U4551, P2_U4552);
  nand ginst15853 (P2_U3054, P2_U4567, P2_U4568, P2_U4569, P2_U4570);
  nand ginst15854 (P2_U3055, P2_U4605, P2_U4606, P2_U4607, P2_U4608);
  nand ginst15855 (P2_U3056, P2_U4513, P2_U4514, P2_U4515, P2_U4516);
  nand ginst15856 (P2_U3057, P2_U4495, P2_U4496, P2_U4497, P2_U4498);
  nand ginst15857 (P2_U3058, P2_U4585, P2_U4586, P2_U4587, P2_U4588);
  nand ginst15858 (P2_U3059, P2_U4117, P2_U4118, P2_U4119, P2_U4120);
  nand ginst15859 (P2_U3060, P2_U4441, P2_U4442, P2_U4443, P2_U4444);
  nand ginst15860 (P2_U3061, P2_U4225, P2_U4226, P2_U4227, P2_U4228);
  nand ginst15861 (P2_U3062, P2_U4243, P2_U4244, P2_U4245, P2_U4246);
  nand ginst15862 (P2_U3063, P2_U4099, P2_U4100, P2_U4101, P2_U4102);
  nand ginst15863 (P2_U3064, P2_U4477, P2_U4478, P2_U4479, P2_U4480);
  nand ginst15864 (P2_U3065, P2_U4459, P2_U4460, P2_U4461, P2_U4462);
  nand ginst15865 (P2_U3066, P2_U4135, P2_U4136, P2_U4137, P2_U4138);
  nand ginst15866 (P2_U3067, P2_U4074, P2_U4075, P2_U4076, P2_U4077);
  nand ginst15867 (P2_U3068, P2_U4351, P2_U4352, P2_U4353, P2_U4354);
  nand ginst15868 (P2_U3069, P2_U4171, P2_U4172, P2_U4173, P2_U4174);
  nand ginst15869 (P2_U3070, P2_U4153, P2_U4154, P2_U4155, P2_U4156);
  nand ginst15870 (P2_U3071, P2_U4261, P2_U4262, P2_U4263, P2_U4264);
  nand ginst15871 (P2_U3072, P2_U4333, P2_U4334, P2_U4335, P2_U4336);
  nand ginst15872 (P2_U3073, P2_U4315, P2_U4316, P2_U4317, P2_U4318);
  nand ginst15873 (P2_U3074, P2_U4423, P2_U4424, P2_U4425, P2_U4426);
  nand ginst15874 (P2_U3075, P2_U4405, P2_U4406, P2_U4407, P2_U4408);
  nand ginst15875 (P2_U3076, P2_U4079, P2_U4080, P2_U4081, P2_U4082);
  nand ginst15876 (P2_U3077, P2_U4055, P2_U4056, P2_U4057, P2_U4058);
  nand ginst15877 (P2_U3078, P2_U4297, P2_U4298, P2_U4299, P2_U4300);
  nand ginst15878 (P2_U3079, P2_U4279, P2_U4280, P2_U4281, P2_U4282);
  nand ginst15879 (P2_U3080, P2_U4387, P2_U4388, P2_U4389, P2_U4390);
  nand ginst15880 (P2_U3081, P2_U4369, P2_U4370, P2_U4371, P2_U4372);
  nand ginst15881 (P2_U3082, P2_U4207, P2_U4208, P2_U4209, P2_U4210);
  nand ginst15882 (P2_U3083, P2_U4189, P2_U4190, P2_U4191, P2_U4192);
  nand ginst15883 (P2_U3084, P2_U5336, P2_U5337);
  nand ginst15884 (P2_U3085, P2_U5338, P2_U5339);
  nand ginst15885 (P2_U3086, P2_U5343, P2_U5344, P2_U5345);
  nand ginst15886 (P2_U3087, P2_U5346, P2_U5347, P2_U5348);
  nand ginst15887 (P2_U3088, P2_U5349, P2_U5350, P2_U5351);
  nand ginst15888 (P2_U3089, P2_U5352, P2_U5353, P2_U5354);
  nand ginst15889 (P2_U3090, P2_U5355, P2_U5356, P2_U5357);
  nand ginst15890 (P2_U3091, P2_U5358, P2_U5359, P2_U5360);
  nand ginst15891 (P2_U3092, P2_U5361, P2_U5362, P2_U5363);
  nand ginst15892 (P2_U3093, P2_U5364, P2_U5365, P2_U5366);
  nand ginst15893 (P2_U3094, P2_U5367, P2_U5368, P2_U5369);
  nand ginst15894 (P2_U3095, P2_U5370, P2_U5371, P2_U5372);
  nand ginst15895 (P2_U3096, P2_U5376, P2_U5377, P2_U5378);
  nand ginst15896 (P2_U3097, P2_U5379, P2_U5380, P2_U5381);
  nand ginst15897 (P2_U3098, P2_U5382, P2_U5383, P2_U5384);
  nand ginst15898 (P2_U3099, P2_U5385, P2_U5386, P2_U5387);
  nand ginst15899 (P2_U3100, P2_U5388, P2_U5389, P2_U5390);
  nand ginst15900 (P2_U3101, P2_U5391, P2_U5392, P2_U5393);
  nand ginst15901 (P2_U3102, P2_U5394, P2_U5395, P2_U5396);
  nand ginst15902 (P2_U3103, P2_U5397, P2_U5398, P2_U5399);
  nand ginst15903 (P2_U3104, P2_U5400, P2_U5401, P2_U5402);
  nand ginst15904 (P2_U3105, P2_U5403, P2_U5404, P2_U5405);
  nand ginst15905 (P2_U3106, P2_U5318, P2_U5319, P2_U5320);
  nand ginst15906 (P2_U3107, P2_U5321, P2_U5322, P2_U5323);
  nand ginst15907 (P2_U3108, P2_U5324, P2_U5325, P2_U5326);
  nand ginst15908 (P2_U3109, P2_U5327, P2_U5328, P2_U5329);
  nand ginst15909 (P2_U3110, P2_U5330, P2_U5331, P2_U5332);
  nand ginst15910 (P2_U3111, P2_U5333, P2_U5334, P2_U5335);
  nand ginst15911 (P2_U3112, P2_U5340, P2_U5341, P2_U5342);
  nand ginst15912 (P2_U3113, P2_U5373, P2_U5374, P2_U5375);
  nand ginst15913 (P2_U3114, P2_U5406, P2_U5407, P2_U5408);
  nand ginst15914 (P2_U3115, P2_U5409, P2_U5410);
  nand ginst15915 (P2_U3116, P2_U5266, P2_U5267);
  nand ginst15916 (P2_U3117, P2_U5268, P2_U5269);
  nand ginst15917 (P2_U3118, P2_U3375, P2_U5272, P2_U5273);
  nand ginst15918 (P2_U3119, P2_U3375, P2_U5274, P2_U5275);
  nand ginst15919 (P2_U3120, P2_U3375, P2_U5276, P2_U5277);
  nand ginst15920 (P2_U3121, P2_U3375, P2_U5278, P2_U5279);
  nand ginst15921 (P2_U3122, P2_U3375, P2_U5280, P2_U5281);
  nand ginst15922 (P2_U3123, P2_U3375, P2_U5282, P2_U5283);
  nand ginst15923 (P2_U3124, P2_U3375, P2_U5284, P2_U5285);
  nand ginst15924 (P2_U3125, P2_U3375, P2_U5286, P2_U5287);
  nand ginst15925 (P2_U3126, P2_U3375, P2_U5288, P2_U5289);
  nand ginst15926 (P2_U3127, P2_U3375, P2_U5290, P2_U5291);
  nand ginst15927 (P2_U3128, P2_U3375, P2_U5294, P2_U5295);
  nand ginst15928 (P2_U3129, P2_U3375, P2_U5296, P2_U5297);
  nand ginst15929 (P2_U3130, P2_U3375, P2_U5298, P2_U5299);
  nand ginst15930 (P2_U3131, P2_U3375, P2_U5300, P2_U5301);
  nand ginst15931 (P2_U3132, P2_U3375, P2_U5302, P2_U5303);
  nand ginst15932 (P2_U3133, P2_U3375, P2_U5304, P2_U5305);
  nand ginst15933 (P2_U3134, P2_U3375, P2_U5306, P2_U5307);
  nand ginst15934 (P2_U3135, P2_U3375, P2_U5308, P2_U5309);
  nand ginst15935 (P2_U3136, P2_U3375, P2_U5310, P2_U5311);
  nand ginst15936 (P2_U3137, P2_U3375, P2_U5312, P2_U5313);
  nand ginst15937 (P2_U3138, P2_U3375, P2_U5254, P2_U5255);
  nand ginst15938 (P2_U3139, P2_U3375, P2_U5256, P2_U5257);
  nand ginst15939 (P2_U3140, P2_U3375, P2_U5258, P2_U5259);
  nand ginst15940 (P2_U3141, P2_U3375, P2_U5260, P2_U5261);
  nand ginst15941 (P2_U3142, P2_U3375, P2_U5262, P2_U5263);
  nand ginst15942 (P2_U3143, P2_U3822, P2_U5265);
  nand ginst15943 (P2_U3144, P2_U3823, P2_U5271);
  nand ginst15944 (P2_U3145, P2_U3824, P2_U5293);
  nand ginst15945 (P2_U3146, P2_U3825, P2_U5315);
  nand ginst15946 (P2_U3147, P2_U3826, P2_U5317);
  nand ginst15947 (P2_U3148, P2_U3375, P2_U3385, P2_U5449);
  nand ginst15948 (P2_U3149, P2_U3013, P2_U3818);
  nand ginst15949 (P2_U3150, P2_U3817, P2_U5249);
  not ginst15950 (P2_U3151, P2_STATE_REG_SCAN_IN);
  nand ginst15951 (P2_U3152, P2_U3359, P2_U5939, P2_U5940);
  nand ginst15952 (P2_U3153, P2_U3816, P2_U5244, P2_U5245, P2_U5246);
  nand ginst15953 (P2_U3154, P2_U3815, P2_U5235, P2_U5236, P2_U5237);
  nand ginst15954 (P2_U3155, P2_U3814, P2_U5226, P2_U5227, P2_U5228);
  nand ginst15955 (P2_U3156, P2_U3813, P2_U5217, P2_U5218, P2_U5219);
  nand ginst15956 (P2_U3157, P2_U3812, P2_U5208, P2_U5209, P2_U5210);
  nand ginst15957 (P2_U3158, P2_U3810, P2_U3811, P2_U5200);
  nand ginst15958 (P2_U3159, P2_U3809, P2_U5190, P2_U5191, P2_U5192);
  nand ginst15959 (P2_U3160, P2_U3808, P2_U5181, P2_U5182, P2_U5183);
  nand ginst15960 (P2_U3161, P2_U3807, P2_U5172, P2_U5173, P2_U5174);
  nand ginst15961 (P2_U3162, P2_U3805, P2_U3806, P2_U5164);
  nand ginst15962 (P2_U3163, P2_U3804, P2_U5154, P2_U5155, P2_U5156);
  nand ginst15963 (P2_U3164, P2_U3803, P2_U5145, P2_U5146, P2_U5147);
  nand ginst15964 (P2_U3165, P2_U3802, P2_U5136, P2_U5137, P2_U5138);
  nand ginst15965 (P2_U3166, P2_U3801, P2_U5127, P2_U5128, P2_U5129);
  nand ginst15966 (P2_U3167, P2_U3800, P2_U5118, P2_U5119, P2_U5120);
  nand ginst15967 (P2_U3168, P2_U3799, P2_U5109, P2_U5110, P2_U5111);
  nand ginst15968 (P2_U3169, P2_U3798, P2_U5100, P2_U5101, P2_U5102);
  nand ginst15969 (P2_U3170, P2_U3796, P2_U3797, P2_U5092);
  nand ginst15970 (P2_U3171, P2_U3795, P2_U5082, P2_U5083, P2_U5084);
  nand ginst15971 (P2_U3172, P2_U3794, P2_U5075);
  nand ginst15972 (P2_U3173, P2_U3791, P2_U5066, P2_U5067, P2_U5068);
  nand ginst15973 (P2_U3174, P2_U3790, P2_U5057, P2_U5058, P2_U5059);
  nand ginst15974 (P2_U3175, P2_U3789, P2_U5048, P2_U5049, P2_U5050);
  nand ginst15975 (P2_U3176, P2_U3788, P2_U5039, P2_U5040, P2_U5041);
  nand ginst15976 (P2_U3177, P2_U3786, P2_U3787, P2_U5031);
  nand ginst15977 (P2_U3178, P2_U3785, P2_U5021, P2_U5022, P2_U5023);
  nand ginst15978 (P2_U3179, P2_U3784, P2_U5012, P2_U5013, P2_U5014);
  nand ginst15979 (P2_U3180, P2_U3783, P2_U5003, P2_U5004, P2_U5005);
  nand ginst15980 (P2_U3181, P2_U3782, P2_U4990, P2_U4991, P2_U4992);
  nand ginst15981 (P2_U3182, P2_U3761, P2_U4969);
  nand ginst15982 (P2_U3183, P2_U3758, P2_U4958);
  nand ginst15983 (P2_U3184, P2_U3755, P2_U4947);
  nand ginst15984 (P2_U3185, P2_U3752, P2_U4936, P2_U4937);
  nand ginst15985 (P2_U3186, P2_U3749, P2_U4925, P2_U4926);
  nand ginst15986 (P2_U3187, P2_U3746, P2_U3748, P2_U4912, P2_U4914);
  nand ginst15987 (P2_U3188, P2_U3743, P2_U4901, P2_U4903);
  nand ginst15988 (P2_U3189, P2_U3740, P2_U3741, P2_U4892);
  nand ginst15989 (P2_U3190, P2_U3737, P2_U3738, P2_U4881);
  nand ginst15990 (P2_U3191, P2_U3734, P2_U4870);
  nand ginst15991 (P2_U3192, P2_U3731, P2_U4859);
  nand ginst15992 (P2_U3193, P2_U3728, P2_U4848);
  nand ginst15993 (P2_U3194, P2_U3725, P2_U4837);
  nand ginst15994 (P2_U3195, P2_U3722, P2_U4826);
  nand ginst15995 (P2_U3196, P2_U3719, P2_U4815);
  nand ginst15996 (P2_U3197, P2_U3716, P2_U4804);
  nand ginst15997 (P2_U3198, P2_U3713, P2_U4793);
  nand ginst15998 (P2_U3199, P2_U3710, P2_U4782);
  nand ginst15999 (P2_U3200, P2_U3707, P2_U4771);
  nand ginst16000 (P2_U3201, P2_U3704, P2_U4760);
  nand ginst16001 (P2_U3202, P2_U3049, P2_U4748, P2_U4749);
  nand ginst16002 (P2_U3203, P2_U3049, P2_U4746, P2_U4747);
  nand ginst16003 (P2_U3204, P2_U3862, P2_U4741, P2_U4742, P2_U4743);
  nand ginst16004 (P2_U3205, P2_U3861, P2_U4737, P2_U4738, P2_U4739, P2_U4740);
  nand ginst16005 (P2_U3206, P2_U3860, P2_U4733, P2_U4734, P2_U4735, P2_U4736);
  nand ginst16006 (P2_U3207, P2_U3859, P2_U4729, P2_U4730, P2_U4731, P2_U4732);
  nand ginst16007 (P2_U3208, P2_U3858, P2_U4725, P2_U4726, P2_U4727, P2_U4728);
  nand ginst16008 (P2_U3209, P2_U3857, P2_U4721, P2_U4722, P2_U4723, P2_U4724);
  nand ginst16009 (P2_U3210, P2_U3856, P2_U4717, P2_U4718, P2_U4719, P2_U4720);
  nand ginst16010 (P2_U3211, P2_U3855, P2_U4713, P2_U4714, P2_U4715, P2_U4716);
  nand ginst16011 (P2_U3212, P2_U3854, P2_U4709, P2_U4710, P2_U4711, P2_U4712);
  nand ginst16012 (P2_U3213, P2_U3853, P2_U4705, P2_U4706, P2_U4707, P2_U4708);
  nand ginst16013 (P2_U3214, P2_U3852, P2_U4701, P2_U4702, P2_U4703, P2_U4704);
  nand ginst16014 (P2_U3215, P2_U3851, P2_U4697, P2_U4698, P2_U4699, P2_U4700);
  nand ginst16015 (P2_U3216, P2_U3850, P2_U4693, P2_U4694, P2_U4695, P2_U4696);
  nand ginst16016 (P2_U3217, P2_U3849, P2_U4689, P2_U4690, P2_U4691, P2_U4692);
  nand ginst16017 (P2_U3218, P2_U3848, P2_U4685, P2_U4686, P2_U4687, P2_U4688);
  nand ginst16018 (P2_U3219, P2_U3847, P2_U4681, P2_U4682, P2_U4683, P2_U4684);
  nand ginst16019 (P2_U3220, P2_U3846, P2_U4677, P2_U4678, P2_U4679, P2_U4680);
  nand ginst16020 (P2_U3221, P2_U3845, P2_U4673, P2_U4674, P2_U4675, P2_U4676);
  nand ginst16021 (P2_U3222, P2_U3844, P2_U4669, P2_U4670, P2_U4671, P2_U4672);
  nand ginst16022 (P2_U3223, P2_U3843, P2_U4665, P2_U4666, P2_U4667, P2_U4668);
  nand ginst16023 (P2_U3224, P2_U3842, P2_U4661, P2_U4662, P2_U4663, P2_U4664);
  nand ginst16024 (P2_U3225, P2_U3841, P2_U4657, P2_U4658, P2_U4659, P2_U4660);
  nand ginst16025 (P2_U3226, P2_U3840, P2_U4653, P2_U4654, P2_U4655, P2_U4656);
  nand ginst16026 (P2_U3227, P2_U3839, P2_U4649, P2_U4650, P2_U4651, P2_U4652);
  nand ginst16027 (P2_U3228, P2_U3838, P2_U4645, P2_U4646, P2_U4647, P2_U4648);
  nand ginst16028 (P2_U3229, P2_U3837, P2_U4641, P2_U4642, P2_U4643, P2_U4644);
  nand ginst16029 (P2_U3230, P2_U3836, P2_U4637, P2_U4638, P2_U4639, P2_U4640);
  nand ginst16030 (P2_U3231, P2_U3835, P2_U4633, P2_U4634, P2_U4635, P2_U4636);
  nand ginst16031 (P2_U3232, P2_U3834, P2_U4629, P2_U4630, P2_U4631, P2_U4632);
  nand ginst16032 (P2_U3233, P2_U3833, P2_U4625, P2_U4626, P2_U4627, P2_U4628);
  and ginst16033 (P2_U3234, P2_D_REG_31__SCAN_IN, P2_U3828);
  and ginst16034 (P2_U3235, P2_D_REG_30__SCAN_IN, P2_U3828);
  and ginst16035 (P2_U3236, P2_D_REG_29__SCAN_IN, P2_U3828);
  and ginst16036 (P2_U3237, P2_D_REG_28__SCAN_IN, P2_U3828);
  and ginst16037 (P2_U3238, P2_D_REG_27__SCAN_IN, P2_U3828);
  and ginst16038 (P2_U3239, P2_D_REG_26__SCAN_IN, P2_U3828);
  and ginst16039 (P2_U3240, P2_D_REG_25__SCAN_IN, P2_U3828);
  and ginst16040 (P2_U3241, P2_D_REG_24__SCAN_IN, P2_U3828);
  and ginst16041 (P2_U3242, P2_D_REG_23__SCAN_IN, P2_U3828);
  and ginst16042 (P2_U3243, P2_D_REG_22__SCAN_IN, P2_U3828);
  and ginst16043 (P2_U3244, P2_D_REG_21__SCAN_IN, P2_U3828);
  and ginst16044 (P2_U3245, P2_D_REG_20__SCAN_IN, P2_U3828);
  and ginst16045 (P2_U3246, P2_D_REG_19__SCAN_IN, P2_U3828);
  and ginst16046 (P2_U3247, P2_D_REG_18__SCAN_IN, P2_U3828);
  and ginst16047 (P2_U3248, P2_D_REG_17__SCAN_IN, P2_U3828);
  and ginst16048 (P2_U3249, P2_D_REG_16__SCAN_IN, P2_U3828);
  and ginst16049 (P2_U3250, P2_D_REG_15__SCAN_IN, P2_U3828);
  and ginst16050 (P2_U3251, P2_D_REG_14__SCAN_IN, P2_U3828);
  and ginst16051 (P2_U3252, P2_D_REG_13__SCAN_IN, P2_U3828);
  and ginst16052 (P2_U3253, P2_D_REG_12__SCAN_IN, P2_U3828);
  and ginst16053 (P2_U3254, P2_D_REG_11__SCAN_IN, P2_U3828);
  and ginst16054 (P2_U3255, P2_D_REG_10__SCAN_IN, P2_U3828);
  and ginst16055 (P2_U3256, P2_D_REG_9__SCAN_IN, P2_U3828);
  and ginst16056 (P2_U3257, P2_D_REG_8__SCAN_IN, P2_U3828);
  and ginst16057 (P2_U3258, P2_D_REG_7__SCAN_IN, P2_U3828);
  and ginst16058 (P2_U3259, P2_D_REG_6__SCAN_IN, P2_U3828);
  and ginst16059 (P2_U3260, P2_D_REG_5__SCAN_IN, P2_U3828);
  and ginst16060 (P2_U3261, P2_D_REG_4__SCAN_IN, P2_U3828);
  and ginst16061 (P2_U3262, P2_D_REG_3__SCAN_IN, P2_U3828);
  and ginst16062 (P2_U3263, P2_D_REG_2__SCAN_IN, P2_U3828);
  nand ginst16063 (P2_U3264, P2_U4011, P2_U4012, P2_U4013);
  nand ginst16064 (P2_U3265, P2_U4008, P2_U4009, P2_U4010);
  nand ginst16065 (P2_U3266, P2_U4005, P2_U4006, P2_U4007);
  nand ginst16066 (P2_U3267, P2_U4002, P2_U4003, P2_U4004);
  nand ginst16067 (P2_U3268, P2_U3999, P2_U4000, P2_U4001);
  nand ginst16068 (P2_U3269, P2_U3996, P2_U3997, P2_U3998);
  nand ginst16069 (P2_U3270, P2_U3993, P2_U3994, P2_U3995);
  nand ginst16070 (P2_U3271, P2_U3990, P2_U3991, P2_U3992);
  nand ginst16071 (P2_U3272, P2_U3987, P2_U3988, P2_U3989);
  nand ginst16072 (P2_U3273, P2_U3984, P2_U3985, P2_U3986);
  nand ginst16073 (P2_U3274, P2_U3981, P2_U3982, P2_U3983);
  nand ginst16074 (P2_U3275, P2_U3978, P2_U3979, P2_U3980);
  nand ginst16075 (P2_U3276, P2_U3975, P2_U3976, P2_U3977);
  nand ginst16076 (P2_U3277, P2_U3972, P2_U3973, P2_U3974);
  nand ginst16077 (P2_U3278, P2_U3969, P2_U3970, P2_U3971);
  nand ginst16078 (P2_U3279, P2_U3966, P2_U3967, P2_U3968);
  nand ginst16079 (P2_U3280, P2_U3963, P2_U3964, P2_U3965);
  nand ginst16080 (P2_U3281, P2_U3960, P2_U3961, P2_U3962);
  nand ginst16081 (P2_U3282, P2_U3957, P2_U3958, P2_U3959);
  nand ginst16082 (P2_U3283, P2_U3954, P2_U3955, P2_U3956);
  nand ginst16083 (P2_U3284, P2_U3951, P2_U3952, P2_U3953);
  nand ginst16084 (P2_U3285, P2_U3948, P2_U3949, P2_U3950);
  nand ginst16085 (P2_U3286, P2_U3945, P2_U3946, P2_U3947);
  nand ginst16086 (P2_U3287, P2_U3942, P2_U3943, P2_U3944);
  nand ginst16087 (P2_U3288, P2_U3939, P2_U3940, P2_U3941);
  nand ginst16088 (P2_U3289, P2_U3936, P2_U3937, P2_U3938);
  nand ginst16089 (P2_U3290, P2_U3933, P2_U3934, P2_U3935);
  nand ginst16090 (P2_U3291, P2_U3930, P2_U3931, P2_U3932);
  nand ginst16091 (P2_U3292, P2_U3927, P2_U3928, P2_U3929);
  nand ginst16092 (P2_U3293, P2_U3924, P2_U3925, P2_U3926);
  nand ginst16093 (P2_U3294, P2_U3921, P2_U3922, P2_U3923);
  nand ginst16094 (P2_U3295, P2_U3918, P2_U3919, P2_U3920);
  and ginst16095 (P2_U3296, P2_U3780, P2_U5417);
  nand ginst16096 (P2_U3297, P2_STATE_REG_SCAN_IN, P2_U3827);
  not ginst16097 (P2_U3298, P2_B_REG_SCAN_IN);
  nand ginst16098 (P2_U3299, P2_U3374, P2_U5427);
  nand ginst16099 (P2_U3300, P2_U3374, P2_U4014);
  nand ginst16100 (P2_U3301, P2_U3013, P2_U5443);
  nand ginst16101 (P2_U3302, P2_U3014, P2_U5452);
  nand ginst16102 (P2_U3303, P2_U3018, P2_U3588);
  nand ginst16103 (P2_U3304, P2_U3018, P2_U3589);
  nand ginst16104 (P2_U3305, P2_U3014, P2_U5443);
  nand ginst16105 (P2_U3306, P2_U3014, P2_U3378);
  nand ginst16106 (P2_U3307, P2_U3013, P2_U3378);
  nand ginst16107 (P2_U3308, P2_U3378, P2_U3379, P2_U3385);
  nand ginst16108 (P2_U3309, P2_U3378, P2_U3385, P2_U5446);
  nand ginst16109 (P2_U3310, P2_U3013, P2_U5452);
  nand ginst16110 (P2_U3311, P2_U3874, P2_U5443);
  nand ginst16111 (P2_U3312, P2_U3016, P2_U3385);
  nand ginst16112 (P2_U3313, P2_U3380, P2_U3385);
  nand ginst16113 (P2_U3314, P2_U3575, P2_U3576, P2_U4065, P2_U4066, P2_U4067);
  nand ginst16114 (P2_U3315, P2_U3590, P2_U3592, P2_U4086, P2_U4087);
  nand ginst16115 (P2_U3316, P2_U3594, P2_U3596, P2_U4104, P2_U4105);
  nand ginst16116 (P2_U3317, P2_U3598, P2_U3600, P2_U4122, P2_U4123);
  nand ginst16117 (P2_U3318, P2_U3602, P2_U3604, P2_U4140, P2_U4141);
  nand ginst16118 (P2_U3319, P2_U3606, P2_U3608, P2_U4158, P2_U4159);
  nand ginst16119 (P2_U3320, P2_U3610, P2_U3612, P2_U4176, P2_U4177);
  nand ginst16120 (P2_U3321, P2_U3614, P2_U3616, P2_U4194, P2_U4195);
  nand ginst16121 (P2_U3322, P2_U3619, P2_U4212, P2_U4213, P2_U4214, P2_U4215);
  nand ginst16122 (P2_U3323, P2_U3622, P2_U4230, P2_U4231, P2_U4232, P2_U4233);
  nand ginst16123 (P2_U3324, P2_U3625, P2_U4248, P2_U4249, P2_U4250, P2_U4251);
  nand ginst16124 (P2_U3325, P2_U3628, P2_U4266, P2_U4267, P2_U4268, P2_U4269);
  nand ginst16125 (P2_U3326, P2_U3630, P2_U3632, P2_U4284, P2_U4285);
  nand ginst16126 (P2_U3327, P2_U3634, P2_U3636, P2_U4302, P2_U4303);
  nand ginst16127 (P2_U3328, P2_U3639, P2_U4320, P2_U4321, P2_U4322, P2_U4323);
  nand ginst16128 (P2_U3329, P2_U3642, P2_U4338, P2_U4339, P2_U4340, P2_U4341);
  nand ginst16129 (P2_U3330, P2_U3645, P2_U4356, P2_U4357, P2_U4358, P2_U4359);
  nand ginst16130 (P2_U3331, P2_U3647, P2_U3649, P2_U4374, P2_U4375);
  nand ginst16131 (P2_U3332, P2_U3651, P2_U3653, P2_U4392, P2_U4393);
  nand ginst16132 (P2_U3333, P2_U3655, P2_U3657, P2_U4410, P2_U4411);
  nand ginst16133 (P2_U3334, P2_U3829, U44);
  nand ginst16134 (P2_U3335, P2_U3659, P2_U3661, P2_U4428, P2_U4429);
  nand ginst16135 (P2_U3336, P2_U3829, U43);
  nand ginst16136 (P2_U3337, P2_U3664, P2_U4446, P2_U4447, P2_U4448, P2_U4449);
  nand ginst16137 (P2_U3338, P2_U3829, U42);
  nand ginst16138 (P2_U3339, P2_U3667, P2_U4464, P2_U4465, P2_U4466, P2_U4467);
  nand ginst16139 (P2_U3340, P2_U3829, U41);
  nand ginst16140 (P2_U3341, P2_U3670, P2_U4482, P2_U4483, P2_U4484, P2_U4485);
  nand ginst16141 (P2_U3342, P2_U3829, U40);
  nand ginst16142 (P2_U3343, P2_U3672, P2_U3674, P2_U4500, P2_U4501);
  nand ginst16143 (P2_U3344, P2_U3829, U39);
  nand ginst16144 (P2_U3345, P2_U3676, P2_U3678, P2_U4518, P2_U4519);
  nand ginst16145 (P2_U3346, P2_U3829, U38);
  nand ginst16146 (P2_U3347, P2_U3680, P2_U3682, P2_U4536, P2_U4537);
  nand ginst16147 (P2_U3348, P2_U3829, U37);
  nand ginst16148 (P2_U3349, P2_U3684, P2_U3686, P2_U4554, P2_U4555);
  nand ginst16149 (P2_U3350, P2_U3829, U36);
  nand ginst16150 (P2_U3351, P2_U3688, P2_U3690, P2_U4572, P2_U4573);
  nand ginst16151 (P2_U3352, P2_U3383, P2_U3384);
  nand ginst16152 (P2_U3353, P2_U3829, U35);
  nand ginst16153 (P2_U3354, P2_U3692, P2_U3694);
  nand ginst16154 (P2_U3355, P2_U3829, U33);
  nand ginst16155 (P2_U3356, P2_U3829, U32);
  nand ginst16156 (P2_U3357, P2_U3015, P2_U5452);
  nand ginst16157 (P2_U3358, P2_U3023, P2_U4623);
  nand ginst16158 (P2_U3359, P2_U3385, P2_U5443);
  nand ginst16159 (P2_U3360, P2_U3875, P2_U5443);
  nand ginst16160 (P2_U3361, P2_U3055, P2_U3907, P2_U4591);
  nand ginst16161 (P2_U3362, P2_U3372, P2_U3373, P2_U3374);
  nand ginst16162 (P2_U3363, P2_U3699, P2_U3906);
  nand ginst16163 (P2_U3364, P2_U3313, P2_U3829);
  nand ginst16164 (P2_U3365, P2_U3873, P2_U5419);
  nand ginst16165 (P2_U3366, P2_U3050, P2_U3700);
  nand ginst16166 (P2_U3367, P2_U3385, P2_U3878);
  nand ginst16167 (P2_U3368, P2_U3764, P2_U3886);
  nand ginst16168 (P2_U3369, P2_U3378, P2_U3872);
  nand ginst16169 (P2_U3370, P2_U3781, P2_U4987, P2_U4988);
  nand ginst16170 (P2_U3371, P2_U3913, P2_U5413);
  nand ginst16171 (P2_U3372, P2_U5422, P2_U5423);
  nand ginst16172 (P2_U3373, P2_U5425, P2_U5426);
  nand ginst16173 (P2_U3374, P2_U5428, P2_U5429);
  nand ginst16174 (P2_U3375, P2_U5434, P2_U5435);
  nand ginst16175 (P2_U3376, P2_U5437, P2_U5438);
  nand ginst16176 (P2_U3377, P2_U5439, P2_U5440);
  nand ginst16177 (P2_U3378, P2_U5441, P2_U5442);
  nand ginst16178 (P2_U3379, P2_U5444, P2_U5445);
  nand ginst16179 (P2_U3380, P2_U5447, P2_U5448);
  nand ginst16180 (P2_U3381, P2_U5453, P2_U5454);
  nand ginst16181 (P2_U3382, P2_U5456, P2_U5457);
  nand ginst16182 (P2_U3383, P2_U5459, P2_U5460);
  nand ginst16183 (P2_U3384, P2_U5462, P2_U5463);
  nand ginst16184 (P2_U3385, P2_U5450, P2_U5451);
  nand ginst16185 (P2_U3386, P2_U5465, P2_U5466);
  nand ginst16186 (P2_U3387, P2_U5467, P2_U5468);
  nand ginst16187 (P2_U3388, P2_U5470, P2_U5471);
  nand ginst16188 (P2_U3389, P2_U5473, P2_U5474);
  nand ginst16189 (P2_U3390, P2_U5479, P2_U5480);
  nand ginst16190 (P2_U3391, P2_U5481, P2_U5482);
  nand ginst16191 (P2_U3392, P2_U5483, P2_U5484);
  nand ginst16192 (P2_U3393, P2_U5486, P2_U5487);
  nand ginst16193 (P2_U3394, P2_U5488, P2_U5489);
  nand ginst16194 (P2_U3395, P2_U5490, P2_U5491);
  nand ginst16195 (P2_U3396, P2_U5493, P2_U5494);
  nand ginst16196 (P2_U3397, P2_U5495, P2_U5496);
  nand ginst16197 (P2_U3398, P2_U5497, P2_U5498);
  nand ginst16198 (P2_U3399, P2_U5500, P2_U5501);
  nand ginst16199 (P2_U3400, P2_U5502, P2_U5503);
  nand ginst16200 (P2_U3401, P2_U5504, P2_U5505);
  nand ginst16201 (P2_U3402, P2_U5507, P2_U5508);
  nand ginst16202 (P2_U3403, P2_U5509, P2_U5510);
  nand ginst16203 (P2_U3404, P2_U5511, P2_U5512);
  nand ginst16204 (P2_U3405, P2_U5514, P2_U5515);
  nand ginst16205 (P2_U3406, P2_U5516, P2_U5517);
  nand ginst16206 (P2_U3407, P2_U5518, P2_U5519);
  nand ginst16207 (P2_U3408, P2_U5521, P2_U5522);
  nand ginst16208 (P2_U3409, P2_U5523, P2_U5524);
  nand ginst16209 (P2_U3410, P2_U5525, P2_U5526);
  nand ginst16210 (P2_U3411, P2_U5528, P2_U5529);
  nand ginst16211 (P2_U3412, P2_U5530, P2_U5531);
  nand ginst16212 (P2_U3413, P2_U5532, P2_U5533);
  nand ginst16213 (P2_U3414, P2_U5535, P2_U5536);
  nand ginst16214 (P2_U3415, P2_U5537, P2_U5538);
  nand ginst16215 (P2_U3416, P2_U5539, P2_U5540);
  nand ginst16216 (P2_U3417, P2_U5542, P2_U5543);
  nand ginst16217 (P2_U3418, P2_U5544, P2_U5545);
  nand ginst16218 (P2_U3419, P2_U5546, P2_U5547);
  nand ginst16219 (P2_U3420, P2_U5549, P2_U5550);
  nand ginst16220 (P2_U3421, P2_U5551, P2_U5552);
  nand ginst16221 (P2_U3422, P2_U5553, P2_U5554);
  nand ginst16222 (P2_U3423, P2_U5556, P2_U5557);
  nand ginst16223 (P2_U3424, P2_U5558, P2_U5559);
  nand ginst16224 (P2_U3425, P2_U5560, P2_U5561);
  nand ginst16225 (P2_U3426, P2_U5563, P2_U5564);
  nand ginst16226 (P2_U3427, P2_U5565, P2_U5566);
  nand ginst16227 (P2_U3428, P2_U5567, P2_U5568);
  nand ginst16228 (P2_U3429, P2_U5570, P2_U5571);
  nand ginst16229 (P2_U3430, P2_U5572, P2_U5573);
  nand ginst16230 (P2_U3431, P2_U5574, P2_U5575);
  nand ginst16231 (P2_U3432, P2_U5577, P2_U5578);
  nand ginst16232 (P2_U3433, P2_U5579, P2_U5580);
  nand ginst16233 (P2_U3434, P2_U5581, P2_U5582);
  nand ginst16234 (P2_U3435, P2_U5584, P2_U5585);
  nand ginst16235 (P2_U3436, P2_U5586, P2_U5587);
  nand ginst16236 (P2_U3437, P2_U5588, P2_U5589);
  nand ginst16237 (P2_U3438, P2_U5591, P2_U5592);
  nand ginst16238 (P2_U3439, P2_U5593, P2_U5594);
  nand ginst16239 (P2_U3440, P2_U5595, P2_U5596);
  nand ginst16240 (P2_U3441, P2_U5598, P2_U5599);
  nand ginst16241 (P2_U3442, P2_U5600, P2_U5601);
  nand ginst16242 (P2_U3443, P2_U5602, P2_U5603);
  nand ginst16243 (P2_U3444, P2_U5605, P2_U5606);
  nand ginst16244 (P2_U3445, P2_U5607, P2_U5608);
  nand ginst16245 (P2_U3446, P2_U5610, P2_U5611);
  nand ginst16246 (P2_U3447, P2_U5612, P2_U5613);
  nand ginst16247 (P2_U3448, P2_U5614, P2_U5615);
  nand ginst16248 (P2_U3449, P2_U5616, P2_U5617);
  nand ginst16249 (P2_U3450, P2_U5618, P2_U5619);
  nand ginst16250 (P2_U3451, P2_U5620, P2_U5621);
  nand ginst16251 (P2_U3452, P2_U5622, P2_U5623);
  nand ginst16252 (P2_U3453, P2_U5624, P2_U5625);
  nand ginst16253 (P2_U3454, P2_U5626, P2_U5627);
  nand ginst16254 (P2_U3455, P2_U5628, P2_U5629);
  nand ginst16255 (P2_U3456, P2_U5630, P2_U5631);
  nand ginst16256 (P2_U3457, P2_U5632, P2_U5633);
  nand ginst16257 (P2_U3458, P2_U5634, P2_U5635);
  nand ginst16258 (P2_U3459, P2_U5638, P2_U5639);
  nand ginst16259 (P2_U3460, P2_U5640, P2_U5641);
  nand ginst16260 (P2_U3461, P2_U5642, P2_U5643);
  nand ginst16261 (P2_U3462, P2_U5644, P2_U5645);
  nand ginst16262 (P2_U3463, P2_U5646, P2_U5647);
  nand ginst16263 (P2_U3464, P2_U5648, P2_U5649);
  nand ginst16264 (P2_U3465, P2_U5650, P2_U5651);
  nand ginst16265 (P2_U3466, P2_U5652, P2_U5653);
  nand ginst16266 (P2_U3467, P2_U5654, P2_U5655);
  nand ginst16267 (P2_U3468, P2_U5656, P2_U5657);
  nand ginst16268 (P2_U3469, P2_U5658, P2_U5659);
  nand ginst16269 (P2_U3470, P2_U5660, P2_U5661);
  nand ginst16270 (P2_U3471, P2_U5662, P2_U5663);
  nand ginst16271 (P2_U3472, P2_U5664, P2_U5665);
  nand ginst16272 (P2_U3473, P2_U5666, P2_U5667);
  nand ginst16273 (P2_U3474, P2_U5668, P2_U5669);
  nand ginst16274 (P2_U3475, P2_U5670, P2_U5671);
  nand ginst16275 (P2_U3476, P2_U5672, P2_U5673);
  nand ginst16276 (P2_U3477, P2_U5674, P2_U5675);
  nand ginst16277 (P2_U3478, P2_U5676, P2_U5677);
  nand ginst16278 (P2_U3479, P2_U5678, P2_U5679);
  nand ginst16279 (P2_U3480, P2_U5680, P2_U5681);
  nand ginst16280 (P2_U3481, P2_U5682, P2_U5683);
  nand ginst16281 (P2_U3482, P2_U5684, P2_U5685);
  nand ginst16282 (P2_U3483, P2_U5686, P2_U5687);
  nand ginst16283 (P2_U3484, P2_U5688, P2_U5689);
  nand ginst16284 (P2_U3485, P2_U5690, P2_U5691);
  nand ginst16285 (P2_U3486, P2_U5692, P2_U5693);
  nand ginst16286 (P2_U3487, P2_U5694, P2_U5695);
  nand ginst16287 (P2_U3488, P2_U5696, P2_U5697);
  nand ginst16288 (P2_U3489, P2_U5698, P2_U5699);
  nand ginst16289 (P2_U3490, P2_U5700, P2_U5701);
  nand ginst16290 (P2_U3491, P2_U5765, P2_U5766);
  nand ginst16291 (P2_U3492, P2_U5767, P2_U5768);
  nand ginst16292 (P2_U3493, P2_U5769, P2_U5770);
  nand ginst16293 (P2_U3494, P2_U5771, P2_U5772);
  nand ginst16294 (P2_U3495, P2_U5773, P2_U5774);
  nand ginst16295 (P2_U3496, P2_U5775, P2_U5776);
  nand ginst16296 (P2_U3497, P2_U5777, P2_U5778);
  nand ginst16297 (P2_U3498, P2_U5779, P2_U5780);
  nand ginst16298 (P2_U3499, P2_U5781, P2_U5782);
  nand ginst16299 (P2_U3500, P2_U5783, P2_U5784);
  nand ginst16300 (P2_U3501, P2_U5785, P2_U5786);
  nand ginst16301 (P2_U3502, P2_U5787, P2_U5788);
  nand ginst16302 (P2_U3503, P2_U5789, P2_U5790);
  nand ginst16303 (P2_U3504, P2_U5791, P2_U5792);
  nand ginst16304 (P2_U3505, P2_U5793, P2_U5794);
  nand ginst16305 (P2_U3506, P2_U5795, P2_U5796);
  nand ginst16306 (P2_U3507, P2_U5797, P2_U5798);
  nand ginst16307 (P2_U3508, P2_U5799, P2_U5800);
  nand ginst16308 (P2_U3509, P2_U5801, P2_U5802);
  nand ginst16309 (P2_U3510, P2_U5803, P2_U5804);
  nand ginst16310 (P2_U3511, P2_U5805, P2_U5806);
  nand ginst16311 (P2_U3512, P2_U5807, P2_U5808);
  nand ginst16312 (P2_U3513, P2_U5809, P2_U5810);
  nand ginst16313 (P2_U3514, P2_U5811, P2_U5812);
  nand ginst16314 (P2_U3515, P2_U5813, P2_U5814);
  nand ginst16315 (P2_U3516, P2_U5815, P2_U5816);
  nand ginst16316 (P2_U3517, P2_U5817, P2_U5818);
  nand ginst16317 (P2_U3518, P2_U5819, P2_U5820);
  nand ginst16318 (P2_U3519, P2_U5821, P2_U5822);
  nand ginst16319 (P2_U3520, P2_U5823, P2_U5824);
  nand ginst16320 (P2_U3521, P2_U5825, P2_U5826);
  nand ginst16321 (P2_U3522, P2_U5827, P2_U5828);
  nand ginst16322 (P2_U3523, P2_U5941, P2_U5942);
  nand ginst16323 (P2_U3524, P2_U5943, P2_U5944);
  nand ginst16324 (P2_U3525, P2_U5945, P2_U5946);
  nand ginst16325 (P2_U3526, P2_U5947, P2_U5948);
  nand ginst16326 (P2_U3527, P2_U5949, P2_U5950);
  nand ginst16327 (P2_U3528, P2_U5951, P2_U5952);
  nand ginst16328 (P2_U3529, P2_U5953, P2_U5954);
  nand ginst16329 (P2_U3530, P2_U5955, P2_U5956);
  nand ginst16330 (P2_U3531, P2_U5957, P2_U5958);
  nand ginst16331 (P2_U3532, P2_U5959, P2_U5960);
  nand ginst16332 (P2_U3533, P2_U5961, P2_U5962);
  nand ginst16333 (P2_U3534, P2_U5963, P2_U5964);
  nand ginst16334 (P2_U3535, P2_U5965, P2_U5966);
  nand ginst16335 (P2_U3536, P2_U5967, P2_U5968);
  nand ginst16336 (P2_U3537, P2_U5969, P2_U5970);
  nand ginst16337 (P2_U3538, P2_U5971, P2_U5972);
  nand ginst16338 (P2_U3539, P2_U5973, P2_U5974);
  nand ginst16339 (P2_U3540, P2_U5975, P2_U5976);
  nand ginst16340 (P2_U3541, P2_U5977, P2_U5978);
  nand ginst16341 (P2_U3542, P2_U5979, P2_U5980);
  nand ginst16342 (P2_U3543, P2_U5981, P2_U5982);
  nand ginst16343 (P2_U3544, P2_U5983, P2_U5984);
  nand ginst16344 (P2_U3545, P2_U5985, P2_U5986);
  nand ginst16345 (P2_U3546, P2_U5987, P2_U5988);
  nand ginst16346 (P2_U3547, P2_U5989, P2_U5990);
  nand ginst16347 (P2_U3548, P2_U5991, P2_U5992);
  nand ginst16348 (P2_U3549, P2_U5993, P2_U5994);
  nand ginst16349 (P2_U3550, P2_U5995, P2_U5996);
  nand ginst16350 (P2_U3551, P2_U5997, P2_U5998);
  nand ginst16351 (P2_U3552, P2_U5999, P2_U6000);
  nand ginst16352 (P2_U3553, P2_U6001, P2_U6002);
  nand ginst16353 (P2_U3554, P2_U6003, P2_U6004);
  nand ginst16354 (P2_U3555, P2_U6005, P2_U6006);
  nand ginst16355 (P2_U3556, P2_U6007, P2_U6008);
  nand ginst16356 (P2_U3557, P2_U6009, P2_U6010);
  nand ginst16357 (P2_U3558, P2_U6011, P2_U6012);
  nand ginst16358 (P2_U3559, P2_U6013, P2_U6014);
  nand ginst16359 (P2_U3560, P2_U6015, P2_U6016);
  nand ginst16360 (P2_U3561, P2_U6017, P2_U6018);
  nand ginst16361 (P2_U3562, P2_U6019, P2_U6020);
  nand ginst16362 (P2_U3563, P2_U6021, P2_U6022);
  nand ginst16363 (P2_U3564, P2_U6023, P2_U6024);
  nand ginst16364 (P2_U3565, P2_U6025, P2_U6026);
  nand ginst16365 (P2_U3566, P2_U6027, P2_U6028);
  nand ginst16366 (P2_U3567, P2_U6029, P2_U6030);
  nand ginst16367 (P2_U3568, P2_U6031, P2_U6032);
  nand ginst16368 (P2_U3569, P2_U6033, P2_U6034);
  nand ginst16369 (P2_U3570, P2_U6035, P2_U6036);
  nand ginst16370 (P2_U3571, P2_U6037, P2_U6038);
  nand ginst16371 (P2_U3572, P2_U6039, P2_U6040);
  nand ginst16372 (P2_U3573, P2_U6041, P2_U6042);
  nand ginst16373 (P2_U3574, P2_U6043, P2_U6044);
  and ginst16374 (P2_U3575, P2_U4061, P2_U4062);
  and ginst16375 (P2_U3576, P2_U4063, P2_U4064);
  and ginst16376 (P2_U3577, P2_U4070, P2_U4071, P2_U4072);
  and ginst16377 (P2_U3578, P2_U4018, P2_U4019, P2_U4020, P2_U4021);
  and ginst16378 (P2_U3579, P2_U4022, P2_U4023, P2_U4024, P2_U4025);
  and ginst16379 (P2_U3580, P2_U4026, P2_U4027, P2_U4028, P2_U4029);
  and ginst16380 (P2_U3581, P2_U4030, P2_U4031, P2_U4032);
  and ginst16381 (P2_U3582, P2_U3578, P2_U3579, P2_U3580, P2_U3581);
  and ginst16382 (P2_U3583, P2_U4033, P2_U4034, P2_U4035, P2_U4036);
  and ginst16383 (P2_U3584, P2_U4037, P2_U4038, P2_U4039, P2_U4040);
  and ginst16384 (P2_U3585, P2_U4041, P2_U4042, P2_U4043, P2_U4044);
  and ginst16385 (P2_U3586, P2_U4045, P2_U4046, P2_U4047);
  and ginst16386 (P2_U3587, P2_U3583, P2_U3584, P2_U3585, P2_U3586);
  and ginst16387 (P2_U3588, P2_U3388, P2_U3389);
  and ginst16388 (P2_U3589, P2_U5472, P2_U5475);
  and ginst16389 (P2_U3590, P2_U4088, P2_U4089);
  and ginst16390 (P2_U3591, P2_U4090, P2_U4091);
  and ginst16391 (P2_U3592, P2_U3591, P2_U4092, P2_U4093);
  and ginst16392 (P2_U3593, P2_U4095, P2_U4096, P2_U4097);
  and ginst16393 (P2_U3594, P2_U4106, P2_U4107);
  and ginst16394 (P2_U3595, P2_U4108, P2_U4109);
  and ginst16395 (P2_U3596, P2_U3595, P2_U4110, P2_U4111);
  and ginst16396 (P2_U3597, P2_U4113, P2_U4114, P2_U4115);
  and ginst16397 (P2_U3598, P2_U4124, P2_U4125);
  and ginst16398 (P2_U3599, P2_U4126, P2_U4127);
  and ginst16399 (P2_U3600, P2_U3599, P2_U4128, P2_U4129);
  and ginst16400 (P2_U3601, P2_U4131, P2_U4132, P2_U4133);
  and ginst16401 (P2_U3602, P2_U4142, P2_U4143);
  and ginst16402 (P2_U3603, P2_U4144, P2_U4145);
  and ginst16403 (P2_U3604, P2_U3603, P2_U4146, P2_U4147);
  and ginst16404 (P2_U3605, P2_U4149, P2_U4150, P2_U4151);
  and ginst16405 (P2_U3606, P2_U4160, P2_U4161);
  and ginst16406 (P2_U3607, P2_U4162, P2_U4163);
  and ginst16407 (P2_U3608, P2_U3607, P2_U4164, P2_U4165);
  and ginst16408 (P2_U3609, P2_U4167, P2_U4168, P2_U4169);
  and ginst16409 (P2_U3610, P2_U4178, P2_U4179);
  and ginst16410 (P2_U3611, P2_U4180, P2_U4181);
  and ginst16411 (P2_U3612, P2_U3611, P2_U4182, P2_U4183);
  and ginst16412 (P2_U3613, P2_U4185, P2_U4186, P2_U4187);
  and ginst16413 (P2_U3614, P2_U4196, P2_U4197);
  and ginst16414 (P2_U3615, P2_U4198, P2_U4199);
  and ginst16415 (P2_U3616, P2_U3615, P2_U4200, P2_U4201);
  and ginst16416 (P2_U3617, P2_U4203, P2_U4204, P2_U4205);
  and ginst16417 (P2_U3618, P2_U4216, P2_U4217);
  and ginst16418 (P2_U3619, P2_U3618, P2_U4218, P2_U4219);
  and ginst16419 (P2_U3620, P2_U4221, P2_U4222, P2_U4223);
  and ginst16420 (P2_U3621, P2_U4234, P2_U4235);
  and ginst16421 (P2_U3622, P2_U3621, P2_U4236, P2_U4237);
  and ginst16422 (P2_U3623, P2_U4239, P2_U4240, P2_U4241);
  and ginst16423 (P2_U3624, P2_U4252, P2_U4253);
  and ginst16424 (P2_U3625, P2_U3624, P2_U4254, P2_U4255);
  and ginst16425 (P2_U3626, P2_U4257, P2_U4258, P2_U4259);
  and ginst16426 (P2_U3627, P2_U4270, P2_U4271);
  and ginst16427 (P2_U3628, P2_U3627, P2_U4272, P2_U4273);
  and ginst16428 (P2_U3629, P2_U4275, P2_U4276, P2_U4277);
  and ginst16429 (P2_U3630, P2_U4286, P2_U4287);
  and ginst16430 (P2_U3631, P2_U4288, P2_U4289);
  and ginst16431 (P2_U3632, P2_U3631, P2_U4290, P2_U4291);
  and ginst16432 (P2_U3633, P2_U4293, P2_U4294, P2_U4295);
  and ginst16433 (P2_U3634, P2_U4304, P2_U4305);
  and ginst16434 (P2_U3635, P2_U4306, P2_U4307);
  and ginst16435 (P2_U3636, P2_U3635, P2_U4308, P2_U4309);
  and ginst16436 (P2_U3637, P2_U4311, P2_U4312, P2_U4313);
  and ginst16437 (P2_U3638, P2_U4324, P2_U4325);
  and ginst16438 (P2_U3639, P2_U3638, P2_U4326, P2_U4327);
  and ginst16439 (P2_U3640, P2_U4329, P2_U4330, P2_U4331);
  and ginst16440 (P2_U3641, P2_U4342, P2_U4343);
  and ginst16441 (P2_U3642, P2_U3641, P2_U4344, P2_U4345);
  and ginst16442 (P2_U3643, P2_U4347, P2_U4348, P2_U4349);
  and ginst16443 (P2_U3644, P2_U4360, P2_U4361);
  and ginst16444 (P2_U3645, P2_U3644, P2_U4362, P2_U4363);
  and ginst16445 (P2_U3646, P2_U4365, P2_U4366, P2_U4367);
  and ginst16446 (P2_U3647, P2_U4376, P2_U4377);
  and ginst16447 (P2_U3648, P2_U4378, P2_U4379);
  and ginst16448 (P2_U3649, P2_U3648, P2_U4380, P2_U4381);
  and ginst16449 (P2_U3650, P2_U4383, P2_U4384, P2_U4385);
  and ginst16450 (P2_U3651, P2_U4394, P2_U4395);
  and ginst16451 (P2_U3652, P2_U4396, P2_U4397);
  and ginst16452 (P2_U3653, P2_U3652, P2_U4398, P2_U4399);
  and ginst16453 (P2_U3654, P2_U4401, P2_U4402, P2_U4403);
  and ginst16454 (P2_U3655, P2_U4412, P2_U4413);
  and ginst16455 (P2_U3656, P2_U4414, P2_U4415);
  and ginst16456 (P2_U3657, P2_U3656, P2_U4416, P2_U4417);
  and ginst16457 (P2_U3658, P2_U4419, P2_U4420, P2_U4421);
  and ginst16458 (P2_U3659, P2_U4430, P2_U4431);
  and ginst16459 (P2_U3660, P2_U4432, P2_U4433);
  and ginst16460 (P2_U3661, P2_U3660, P2_U4434, P2_U4435);
  and ginst16461 (P2_U3662, P2_U4437, P2_U4438, P2_U4439);
  and ginst16462 (P2_U3663, P2_U4450, P2_U4451);
  and ginst16463 (P2_U3664, P2_U3663, P2_U4452, P2_U4453);
  and ginst16464 (P2_U3665, P2_U4455, P2_U4456, P2_U4457);
  and ginst16465 (P2_U3666, P2_U4468, P2_U4469);
  and ginst16466 (P2_U3667, P2_U3666, P2_U4470, P2_U4471);
  and ginst16467 (P2_U3668, P2_U4473, P2_U4474, P2_U4475);
  and ginst16468 (P2_U3669, P2_U4486, P2_U4487);
  and ginst16469 (P2_U3670, P2_U3669, P2_U4488, P2_U4489);
  and ginst16470 (P2_U3671, P2_U4491, P2_U4492, P2_U4493);
  and ginst16471 (P2_U3672, P2_U4502, P2_U4503);
  and ginst16472 (P2_U3673, P2_U4504, P2_U4505);
  and ginst16473 (P2_U3674, P2_U3673, P2_U4506, P2_U4507);
  and ginst16474 (P2_U3675, P2_U4509, P2_U4510, P2_U4511);
  and ginst16475 (P2_U3676, P2_U4520, P2_U4521);
  and ginst16476 (P2_U3677, P2_U4522, P2_U4523);
  and ginst16477 (P2_U3678, P2_U3677, P2_U4524, P2_U4525);
  and ginst16478 (P2_U3679, P2_U4527, P2_U4528, P2_U4529);
  and ginst16479 (P2_U3680, P2_U4538, P2_U4539);
  and ginst16480 (P2_U3681, P2_U4540, P2_U4541);
  and ginst16481 (P2_U3682, P2_U3681, P2_U4542, P2_U4543);
  and ginst16482 (P2_U3683, P2_U4545, P2_U4546, P2_U4547);
  and ginst16483 (P2_U3684, P2_U4556, P2_U4557);
  and ginst16484 (P2_U3685, P2_U4558, P2_U4559);
  and ginst16485 (P2_U3686, P2_U3685, P2_U4560, P2_U4561);
  and ginst16486 (P2_U3687, P2_U4563, P2_U4564, P2_U4565);
  and ginst16487 (P2_U3688, P2_U4574, P2_U4575);
  and ginst16488 (P2_U3689, P2_U4576, P2_U4577);
  and ginst16489 (P2_U3690, P2_U3689, P2_U4578, P2_U4579);
  and ginst16490 (P2_U3691, P2_U4581, P2_U4582, P2_U4583);
  and ginst16491 (P2_U3692, P2_U4592, P2_U4593, P2_U4594, P2_U4595, P2_U4596);
  and ginst16492 (P2_U3693, P2_U4597, P2_U4598);
  and ginst16493 (P2_U3694, P2_U3693, P2_U4599, P2_U4600);
  and ginst16494 (P2_U3695, P2_U4602, P2_U4603);
  and ginst16495 (P2_U3696, P2_U3389, P2_U5472);
  and ginst16496 (P2_U3697, P2_U3388, P2_U5475);
  and ginst16497 (P2_U3698, P2_U3379, P2_U3916);
  and ginst16498 (P2_U3699, P2_STATE_REG_SCAN_IN, P2_U5436);
  and ginst16499 (P2_U3700, P2_U3364, P2_U5420);
  and ginst16500 (P2_U3701, P2_STATE_REG_SCAN_IN, P2_U3375);
  and ginst16501 (P2_U3702, P2_U3301, P2_U3305, P2_U3306, P2_U3307, P2_U3308);
  and ginst16502 (P2_U3703, P2_U3309, P2_U3360);
  and ginst16503 (P2_U3704, P2_U3706, P2_U4758, P2_U4759, P2_U4761);
  and ginst16504 (P2_U3705, P2_U4762, P2_U4764);
  and ginst16505 (P2_U3706, P2_U3705, P2_U4763);
  and ginst16506 (P2_U3707, P2_U3709, P2_U4769, P2_U4770, P2_U4772);
  and ginst16507 (P2_U3708, P2_U4773, P2_U4775);
  and ginst16508 (P2_U3709, P2_U3708, P2_U4774);
  and ginst16509 (P2_U3710, P2_U3712, P2_U4780, P2_U4781, P2_U4783);
  and ginst16510 (P2_U3711, P2_U4784, P2_U4786);
  and ginst16511 (P2_U3712, P2_U3711, P2_U4785);
  and ginst16512 (P2_U3713, P2_U3715, P2_U4791, P2_U4792, P2_U4794);
  and ginst16513 (P2_U3714, P2_U4795, P2_U4797);
  and ginst16514 (P2_U3715, P2_U3714, P2_U4796);
  and ginst16515 (P2_U3716, P2_U3718, P2_U4802, P2_U4803, P2_U4805);
  and ginst16516 (P2_U3717, P2_U4806, P2_U4808);
  and ginst16517 (P2_U3718, P2_U3717, P2_U4807);
  and ginst16518 (P2_U3719, P2_U3721, P2_U4813, P2_U4814, P2_U4816);
  and ginst16519 (P2_U3720, P2_U4817, P2_U4819);
  and ginst16520 (P2_U3721, P2_U3720, P2_U4818);
  and ginst16521 (P2_U3722, P2_U3724, P2_U4824, P2_U4825, P2_U4827);
  and ginst16522 (P2_U3723, P2_U4828, P2_U4830);
  and ginst16523 (P2_U3724, P2_U3723, P2_U4829);
  and ginst16524 (P2_U3725, P2_U3727, P2_U4835, P2_U4836, P2_U4838);
  and ginst16525 (P2_U3726, P2_U4839, P2_U4841);
  and ginst16526 (P2_U3727, P2_U3726, P2_U4840);
  and ginst16527 (P2_U3728, P2_U3730, P2_U4846, P2_U4847, P2_U4849);
  and ginst16528 (P2_U3729, P2_U4850, P2_U4852);
  and ginst16529 (P2_U3730, P2_U3729, P2_U4851);
  and ginst16530 (P2_U3731, P2_U3733, P2_U4857, P2_U4858, P2_U4860);
  and ginst16531 (P2_U3732, P2_U4861, P2_U4863);
  and ginst16532 (P2_U3733, P2_U3732, P2_U4862);
  and ginst16533 (P2_U3734, P2_U3736, P2_U4868, P2_U4869, P2_U4871);
  and ginst16534 (P2_U3735, P2_U4872, P2_U4874);
  and ginst16535 (P2_U3736, P2_U3735, P2_U4873);
  and ginst16536 (P2_U3737, P2_U4879, P2_U4880);
  and ginst16537 (P2_U3738, P2_U3739, P2_U4882, P2_U4884);
  and ginst16538 (P2_U3739, P2_U4883, P2_U4885);
  and ginst16539 (P2_U3740, P2_U4890, P2_U4891);
  and ginst16540 (P2_U3741, P2_U3742, P2_U4893, P2_U4895);
  and ginst16541 (P2_U3742, P2_U4894, P2_U4896);
  and ginst16542 (P2_U3743, P2_U3745, P2_U4902, P2_U4904);
  and ginst16543 (P2_U3744, P2_U4905, P2_U4907);
  and ginst16544 (P2_U3745, P2_U3744, P2_U4906);
  and ginst16545 (P2_U3746, P2_U4913, P2_U4915);
  and ginst16546 (P2_U3747, P2_U4916, P2_U4918);
  and ginst16547 (P2_U3748, P2_U3747, P2_U4917);
  and ginst16548 (P2_U3749, P2_U3751, P2_U4923, P2_U4924);
  and ginst16549 (P2_U3750, P2_U4927, P2_U4929);
  and ginst16550 (P2_U3751, P2_U3750, P2_U4928);
  and ginst16551 (P2_U3752, P2_U3754, P2_U4934, P2_U4935);
  and ginst16552 (P2_U3753, P2_U4938, P2_U4940);
  and ginst16553 (P2_U3754, P2_U3753, P2_U4939);
  and ginst16554 (P2_U3755, P2_U3757, P2_U4945, P2_U4946, P2_U4948);
  and ginst16555 (P2_U3756, P2_U4949, P2_U4951);
  and ginst16556 (P2_U3757, P2_U3756, P2_U4950);
  and ginst16557 (P2_U3758, P2_U3760, P2_U4956, P2_U4957, P2_U4959);
  and ginst16558 (P2_U3759, P2_U4960, P2_U4962);
  and ginst16559 (P2_U3760, P2_U3759, P2_U4961);
  and ginst16560 (P2_U3761, P2_U3763, P2_U4967, P2_U4968, P2_U4970);
  and ginst16561 (P2_U3762, P2_U4971, P2_U4973);
  and ginst16562 (P2_U3763, P2_U3762, P2_U4972);
  and ginst16563 (P2_U3764, P2_U3383, P2_U5464);
  nand ginst16564 (P2_U3765, P2_U5829, P2_U5830);
  and ginst16565 (P2_U3766, P2_U5908, P2_U5911);
  and ginst16566 (P2_U3767, P2_U3766, P2_U3768, P2_U3769, P2_U5893);
  and ginst16567 (P2_U3768, P2_U5896, P2_U5899);
  and ginst16568 (P2_U3769, P2_U5902, P2_U5905);
  and ginst16569 (P2_U3770, P2_U5872, P2_U5875, P2_U5878);
  and ginst16570 (P2_U3771, P2_U5881, P2_U5884, P2_U5887, P2_U5890);
  and ginst16571 (P2_U3772, P2_U3770, P2_U3771, P2_U5869);
  and ginst16572 (P2_U3773, P2_U5854, P2_U5857, P2_U5860, P2_U5863);
  and ginst16573 (P2_U3774, P2_U5848, P2_U5851);
  and ginst16574 (P2_U3775, P2_U5917, P2_U5920, P2_U5923, P2_U5926);
  and ginst16575 (P2_U3776, P2_U5836, P2_U5839, P2_U5842);
  and ginst16576 (P2_U3777, P2_U3773, P2_U3774, P2_U3776, P2_U5845, P2_U5866);
  and ginst16577 (P2_U3778, P2_U3767, P2_U3772, P2_U3775, P2_U5914, P2_U5929);
  and ginst16578 (P2_U3779, P2_U3866, P2_U4976, P2_U4977);
  and ginst16579 (P2_U3780, P2_U5411, P2_U5412);
  and ginst16580 (P2_U3781, P2_U3362, P2_U3876, P2_U4986, P2_U5436);
  and ginst16581 (P2_U3782, P2_U4993, P2_U4994);
  and ginst16582 (P2_U3783, P2_U5006, P2_U5007);
  and ginst16583 (P2_U3784, P2_U5015, P2_U5016);
  and ginst16584 (P2_U3785, P2_U5024, P2_U5025);
  and ginst16585 (P2_U3786, P2_U5030, P2_U5032);
  and ginst16586 (P2_U3787, P2_U5033, P2_U5034);
  and ginst16587 (P2_U3788, P2_U5042, P2_U5043);
  and ginst16588 (P2_U3789, P2_U5051, P2_U5052);
  and ginst16589 (P2_U3790, P2_U5060, P2_U5061);
  and ginst16590 (P2_U3791, P2_U5069, P2_U5070);
  and ginst16591 (P2_U3792, P2_U3031, P2_U3077);
  and ginst16592 (P2_U3793, P2_U5073, P2_U5074);
  and ginst16593 (P2_U3794, P2_U3793, P2_U5076, P2_U5077);
  and ginst16594 (P2_U3795, P2_U5085, P2_U5086);
  and ginst16595 (P2_U3796, P2_U5091, P2_U5093);
  and ginst16596 (P2_U3797, P2_U5094, P2_U5095);
  and ginst16597 (P2_U3798, P2_U5103, P2_U5104);
  and ginst16598 (P2_U3799, P2_U5112, P2_U5113);
  and ginst16599 (P2_U3800, P2_U5121, P2_U5122);
  and ginst16600 (P2_U3801, P2_U5130, P2_U5131);
  and ginst16601 (P2_U3802, P2_U5139, P2_U5140);
  and ginst16602 (P2_U3803, P2_U5148, P2_U5149);
  and ginst16603 (P2_U3804, P2_U5157, P2_U5158);
  and ginst16604 (P2_U3805, P2_U5163, P2_U5165);
  and ginst16605 (P2_U3806, P2_U5166, P2_U5167);
  and ginst16606 (P2_U3807, P2_U5175, P2_U5176);
  and ginst16607 (P2_U3808, P2_U5184, P2_U5185);
  and ginst16608 (P2_U3809, P2_U5193, P2_U5194);
  and ginst16609 (P2_U3810, P2_U5199, P2_U5201);
  and ginst16610 (P2_U3811, P2_U5202, P2_U5203);
  and ginst16611 (P2_U3812, P2_U5211, P2_U5212);
  and ginst16612 (P2_U3813, P2_U5220, P2_U5221);
  and ginst16613 (P2_U3814, P2_U5229, P2_U5230);
  and ginst16614 (P2_U3815, P2_U5238, P2_U5239);
  and ginst16615 (P2_U3816, P2_U5247, P2_U5248);
  and ginst16616 (P2_U3817, P2_STATE_REG_SCAN_IN, P2_U5250);
  and ginst16617 (P2_U3818, P2_U3385, P2_U5436);
  and ginst16618 (P2_U3819, P2_U3375, P2_U3385);
  and ginst16619 (P2_U3820, P2_U3302, P2_U3312, P2_U3871);
  and ginst16620 (P2_U3821, P2_U3310, P2_U3357, P2_U3873);
  and ginst16621 (P2_U3822, P2_U3375, P2_U5264);
  and ginst16622 (P2_U3823, P2_U3375, P2_U5270);
  and ginst16623 (P2_U3824, P2_U3375, P2_U5292);
  and ginst16624 (P2_U3825, P2_U3375, P2_U5314);
  and ginst16625 (P2_U3826, P2_U3375, P2_U5316);
  not ginst16626 (P2_U3827, P2_IR_REG_31__SCAN_IN);
  nand ginst16627 (P2_U3828, P2_U3023, P2_U3300);
  nand ginst16628 (P2_U3829, P2_U5461, P2_U5464);
  nand ginst16629 (P2_U3830, P2_U5443, P2_U5452);
  nand ginst16630 (P2_U3831, P2_U3023, P2_U4054);
  nand ginst16631 (P2_U3832, P2_U3023, P2_U4618);
  and ginst16632 (P2_U3833, P2_U5702, P2_U5703);
  and ginst16633 (P2_U3834, P2_U5704, P2_U5705);
  and ginst16634 (P2_U3835, P2_U5706, P2_U5707);
  and ginst16635 (P2_U3836, P2_U5708, P2_U5709);
  and ginst16636 (P2_U3837, P2_U5710, P2_U5711);
  and ginst16637 (P2_U3838, P2_U5712, P2_U5713);
  and ginst16638 (P2_U3839, P2_U5714, P2_U5715);
  and ginst16639 (P2_U3840, P2_U5716, P2_U5717);
  and ginst16640 (P2_U3841, P2_U5718, P2_U5719);
  and ginst16641 (P2_U3842, P2_U5720, P2_U5721);
  and ginst16642 (P2_U3843, P2_U5722, P2_U5723);
  and ginst16643 (P2_U3844, P2_U5724, P2_U5725);
  and ginst16644 (P2_U3845, P2_U5726, P2_U5727);
  and ginst16645 (P2_U3846, P2_U5728, P2_U5729);
  and ginst16646 (P2_U3847, P2_U5730, P2_U5731);
  and ginst16647 (P2_U3848, P2_U5732, P2_U5733);
  and ginst16648 (P2_U3849, P2_U5734, P2_U5735);
  and ginst16649 (P2_U3850, P2_U5736, P2_U5737);
  and ginst16650 (P2_U3851, P2_U5738, P2_U5739);
  and ginst16651 (P2_U3852, P2_U5740, P2_U5741);
  and ginst16652 (P2_U3853, P2_U5742, P2_U5743);
  and ginst16653 (P2_U3854, P2_U5744, P2_U5745);
  and ginst16654 (P2_U3855, P2_U5746, P2_U5747);
  and ginst16655 (P2_U3856, P2_U5748, P2_U5749);
  and ginst16656 (P2_U3857, P2_U5750, P2_U5751);
  and ginst16657 (P2_U3858, P2_U5752, P2_U5753);
  and ginst16658 (P2_U3859, P2_U5754, P2_U5755);
  and ginst16659 (P2_U3860, P2_U5756, P2_U5757);
  and ginst16660 (P2_U3861, P2_U5758, P2_U5759);
  and ginst16661 (P2_U3862, P2_U5760, P2_U5761);
  not ginst16662 (P2_U3863, P2_R1269_U22);
  nand ginst16663 (P2_U3864, P2_U3777, P2_U3778);
  not ginst16664 (P2_U3865, P2_R693_U14);
  and ginst16665 (P2_U3866, P2_U5935, P2_U5936);
  not ginst16666 (P2_U3867, P2_R1297_U6);
  not ginst16667 (P2_U3868, P2_U3356);
  not ginst16668 (P2_U3869, P2_U3355);
  not ginst16669 (P2_U3870, P2_U3312);
  nand ginst16670 (P2_U3871, P2_U3015, P2_U3385);
  not ginst16671 (P2_U3872, P2_U3302);
  nand ginst16672 (P2_U3873, P2_U3016, P2_U5452);
  not ginst16673 (P2_U3874, P2_U3310);
  not ginst16674 (P2_U3875, P2_U3357);
  nand ginst16675 (P2_U3876, P2_U3014, P2_U3385);
  not ginst16676 (P2_U3877, P2_U3308);
  not ginst16677 (P2_U3878, P2_U3301);
  not ginst16678 (P2_U3879, P2_U3305);
  not ginst16679 (P2_U3880, P2_U3307);
  not ginst16680 (P2_U3881, P2_U3306);
  not ginst16681 (P2_U3882, P2_U3360);
  not ginst16682 (P2_U3883, P2_U3311);
  nand ginst16683 (P2_U3884, P2_U3378, P2_U3874);
  not ginst16684 (P2_U3885, P2_U3369);
  not ginst16685 (P2_U3886, P2_U3367);
  not ginst16686 (P2_U3887, P2_U3309);
  not ginst16687 (P2_U3888, P2_U3352);
  not ginst16688 (P2_U3889, P2_U3829);
  not ginst16689 (P2_U3890, P2_U3303);
  not ginst16690 (P2_U3891, P2_U3304);
  nand ginst16691 (P2_U3892, P2_U3384, P2_U5461);
  not ginst16692 (P2_U3893, P2_U3363);
  not ginst16693 (P2_U3894, P2_U3364);
  not ginst16694 (P2_U3895, P2_U3350);
  not ginst16695 (P2_U3896, P2_U3348);
  not ginst16696 (P2_U3897, P2_U3346);
  not ginst16697 (P2_U3898, P2_U3344);
  not ginst16698 (P2_U3899, P2_U3342);
  not ginst16699 (P2_U3900, P2_U3340);
  not ginst16700 (P2_U3901, P2_U3338);
  not ginst16701 (P2_U3902, P2_U3336);
  not ginst16702 (P2_U3903, P2_U3334);
  not ginst16703 (P2_U3904, P2_U3353);
  not ginst16704 (P2_U3905, P2_U3368);
  not ginst16705 (P2_U3906, P2_U3362);
  not ginst16706 (P2_U3907, P2_U3313);
  not ginst16707 (P2_U3908, P2_U3358);
  not ginst16708 (P2_U3909, P2_U3832);
  not ginst16709 (P2_U3910, P2_U3831);
  not ginst16710 (P2_U3911, P2_U3828);
  not ginst16711 (P2_U3912, P2_U3361);
  nand ginst16712 (P2_U3913, P2_STATE_REG_SCAN_IN, P2_U3370);
  nand ginst16713 (P2_U3914, P2_U3023, P2_U3882);
  not ginst16714 (P2_U3915, P2_U3299);
  not ginst16715 (P2_U3916, P2_U3359);
  not ginst16716 (P2_U3917, P2_U3297);
  nand ginst16717 (P2_U3918, P2_U3151, U56);
  nand ginst16718 (P2_U3919, P2_IR_REG_0__SCAN_IN, P2_U3027);
  nand ginst16719 (P2_U3920, P2_IR_REG_0__SCAN_IN, P2_U3917);
  nand ginst16720 (P2_U3921, P2_U3151, U45);
  nand ginst16721 (P2_U3922, P2_SUB_594_U53, P2_U3027);
  nand ginst16722 (P2_U3923, P2_IR_REG_1__SCAN_IN, P2_U3917);
  nand ginst16723 (P2_U3924, P2_U3151, U34);
  nand ginst16724 (P2_U3925, P2_SUB_594_U23, P2_U3027);
  nand ginst16725 (P2_U3926, P2_IR_REG_2__SCAN_IN, P2_U3917);
  nand ginst16726 (P2_U3927, P2_U3151, U31);
  nand ginst16727 (P2_U3928, P2_SUB_594_U24, P2_U3027);
  nand ginst16728 (P2_U3929, P2_IR_REG_3__SCAN_IN, P2_U3917);
  nand ginst16729 (P2_U3930, P2_U3151, U30);
  nand ginst16730 (P2_U3931, P2_SUB_594_U25, P2_U3027);
  nand ginst16731 (P2_U3932, P2_IR_REG_4__SCAN_IN, P2_U3917);
  nand ginst16732 (P2_U3933, P2_U3151, U29);
  nand ginst16733 (P2_U3934, P2_SUB_594_U72, P2_U3027);
  nand ginst16734 (P2_U3935, P2_IR_REG_5__SCAN_IN, P2_U3917);
  nand ginst16735 (P2_U3936, P2_U3151, U28);
  nand ginst16736 (P2_U3937, P2_SUB_594_U26, P2_U3027);
  nand ginst16737 (P2_U3938, P2_IR_REG_6__SCAN_IN, P2_U3917);
  nand ginst16738 (P2_U3939, P2_U3151, U27);
  nand ginst16739 (P2_U3940, P2_SUB_594_U27, P2_U3027);
  nand ginst16740 (P2_U3941, P2_IR_REG_7__SCAN_IN, P2_U3917);
  nand ginst16741 (P2_U3942, P2_U3151, U26);
  nand ginst16742 (P2_U3943, P2_SUB_594_U28, P2_U3027);
  nand ginst16743 (P2_U3944, P2_IR_REG_8__SCAN_IN, P2_U3917);
  nand ginst16744 (P2_U3945, P2_U3151, U25);
  nand ginst16745 (P2_U3946, P2_SUB_594_U70, P2_U3027);
  nand ginst16746 (P2_U3947, P2_IR_REG_9__SCAN_IN, P2_U3917);
  nand ginst16747 (P2_U3948, P2_U3151, U55);
  nand ginst16748 (P2_U3949, P2_SUB_594_U8, P2_U3027);
  nand ginst16749 (P2_U3950, P2_IR_REG_10__SCAN_IN, P2_U3917);
  nand ginst16750 (P2_U3951, P2_U3151, U54);
  nand ginst16751 (P2_U3952, P2_SUB_594_U9, P2_U3027);
  nand ginst16752 (P2_U3953, P2_IR_REG_11__SCAN_IN, P2_U3917);
  nand ginst16753 (P2_U3954, P2_U3151, U53);
  nand ginst16754 (P2_U3955, P2_SUB_594_U10, P2_U3027);
  nand ginst16755 (P2_U3956, P2_IR_REG_12__SCAN_IN, P2_U3917);
  nand ginst16756 (P2_U3957, P2_U3151, U52);
  nand ginst16757 (P2_U3958, P2_SUB_594_U87, P2_U3027);
  nand ginst16758 (P2_U3959, P2_IR_REG_13__SCAN_IN, P2_U3917);
  nand ginst16759 (P2_U3960, P2_U3151, U51);
  nand ginst16760 (P2_U3961, P2_SUB_594_U11, P2_U3027);
  nand ginst16761 (P2_U3962, P2_IR_REG_14__SCAN_IN, P2_U3917);
  nand ginst16762 (P2_U3963, P2_U3151, U50);
  nand ginst16763 (P2_U3964, P2_SUB_594_U12, P2_U3027);
  nand ginst16764 (P2_U3965, P2_IR_REG_15__SCAN_IN, P2_U3917);
  nand ginst16765 (P2_U3966, P2_U3151, U49);
  nand ginst16766 (P2_U3967, P2_SUB_594_U13, P2_U3027);
  nand ginst16767 (P2_U3968, P2_IR_REG_16__SCAN_IN, P2_U3917);
  nand ginst16768 (P2_U3969, P2_U3151, U48);
  nand ginst16769 (P2_U3970, P2_SUB_594_U85, P2_U3027);
  nand ginst16770 (P2_U3971, P2_IR_REG_17__SCAN_IN, P2_U3917);
  nand ginst16771 (P2_U3972, P2_U3151, U47);
  nand ginst16772 (P2_U3973, P2_SUB_594_U14, P2_U3027);
  nand ginst16773 (P2_U3974, P2_IR_REG_18__SCAN_IN, P2_U3917);
  nand ginst16774 (P2_U3975, P2_U3151, U46);
  nand ginst16775 (P2_U3976, P2_SUB_594_U15, P2_U3027);
  nand ginst16776 (P2_U3977, P2_IR_REG_19__SCAN_IN, P2_U3917);
  nand ginst16777 (P2_U3978, P2_U3151, U44);
  nand ginst16778 (P2_U3979, P2_SUB_594_U16, P2_U3027);
  nand ginst16779 (P2_U3980, P2_IR_REG_20__SCAN_IN, P2_U3917);
  nand ginst16780 (P2_U3981, P2_U3151, U43);
  nand ginst16781 (P2_U3982, P2_SUB_594_U81, P2_U3027);
  nand ginst16782 (P2_U3983, P2_IR_REG_21__SCAN_IN, P2_U3917);
  nand ginst16783 (P2_U3984, P2_U3151, U42);
  nand ginst16784 (P2_U3985, P2_SUB_594_U17, P2_U3027);
  nand ginst16785 (P2_U3986, P2_IR_REG_22__SCAN_IN, P2_U3917);
  nand ginst16786 (P2_U3987, P2_U3151, U41);
  nand ginst16787 (P2_U3988, P2_SUB_594_U18, P2_U3027);
  nand ginst16788 (P2_U3989, P2_IR_REG_23__SCAN_IN, P2_U3917);
  nand ginst16789 (P2_U3990, P2_U3151, U40);
  nand ginst16790 (P2_U3991, P2_SUB_594_U19, P2_U3027);
  nand ginst16791 (P2_U3992, P2_IR_REG_24__SCAN_IN, P2_U3917);
  nand ginst16792 (P2_U3993, P2_U3151, U39);
  nand ginst16793 (P2_U3994, P2_SUB_594_U79, P2_U3027);
  nand ginst16794 (P2_U3995, P2_IR_REG_25__SCAN_IN, P2_U3917);
  nand ginst16795 (P2_U3996, P2_U3151, U38);
  nand ginst16796 (P2_U3997, P2_SUB_594_U20, P2_U3027);
  nand ginst16797 (P2_U3998, P2_IR_REG_26__SCAN_IN, P2_U3917);
  nand ginst16798 (P2_U3999, P2_U3151, U37);
  nand ginst16799 (P2_U4000, P2_SUB_594_U77, P2_U3027);
  nand ginst16800 (P2_U4001, P2_IR_REG_27__SCAN_IN, P2_U3917);
  nand ginst16801 (P2_U4002, P2_U3151, U36);
  nand ginst16802 (P2_U4003, P2_SUB_594_U21, P2_U3027);
  nand ginst16803 (P2_U4004, P2_IR_REG_28__SCAN_IN, P2_U3917);
  nand ginst16804 (P2_U4005, P2_U3151, U35);
  nand ginst16805 (P2_U4006, P2_SUB_594_U22, P2_U3027);
  nand ginst16806 (P2_U4007, P2_IR_REG_29__SCAN_IN, P2_U3917);
  nand ginst16807 (P2_U4008, P2_U3151, U33);
  nand ginst16808 (P2_U4009, P2_SUB_594_U75, P2_U3027);
  nand ginst16809 (P2_U4010, P2_IR_REG_30__SCAN_IN, P2_U3917);
  nand ginst16810 (P2_U4011, P2_U3151, U32);
  nand ginst16811 (P2_U4012, P2_SUB_594_U54, P2_U3027);
  nand ginst16812 (P2_U4013, P2_IR_REG_31__SCAN_IN, P2_U3917);
  nand ginst16813 (P2_U4014, P2_U3915, P2_U5433);
  not ginst16814 (P2_U4015, P2_U3300);
  nand ginst16815 (P2_U4016, P2_U3299, P2_U5424);
  nand ginst16816 (P2_U4017, P2_U3299, P2_U5427);
  nand ginst16817 (P2_U4018, P2_D_REG_10__SCAN_IN, P2_U4015);
  nand ginst16818 (P2_U4019, P2_D_REG_11__SCAN_IN, P2_U4015);
  nand ginst16819 (P2_U4020, P2_D_REG_12__SCAN_IN, P2_U4015);
  nand ginst16820 (P2_U4021, P2_D_REG_13__SCAN_IN, P2_U4015);
  nand ginst16821 (P2_U4022, P2_D_REG_14__SCAN_IN, P2_U4015);
  nand ginst16822 (P2_U4023, P2_D_REG_15__SCAN_IN, P2_U4015);
  nand ginst16823 (P2_U4024, P2_D_REG_16__SCAN_IN, P2_U4015);
  nand ginst16824 (P2_U4025, P2_D_REG_17__SCAN_IN, P2_U4015);
  nand ginst16825 (P2_U4026, P2_D_REG_18__SCAN_IN, P2_U4015);
  nand ginst16826 (P2_U4027, P2_D_REG_19__SCAN_IN, P2_U4015);
  nand ginst16827 (P2_U4028, P2_D_REG_20__SCAN_IN, P2_U4015);
  nand ginst16828 (P2_U4029, P2_D_REG_21__SCAN_IN, P2_U4015);
  nand ginst16829 (P2_U4030, P2_D_REG_22__SCAN_IN, P2_U4015);
  nand ginst16830 (P2_U4031, P2_D_REG_23__SCAN_IN, P2_U4015);
  nand ginst16831 (P2_U4032, P2_D_REG_24__SCAN_IN, P2_U4015);
  nand ginst16832 (P2_U4033, P2_D_REG_25__SCAN_IN, P2_U4015);
  nand ginst16833 (P2_U4034, P2_D_REG_26__SCAN_IN, P2_U4015);
  nand ginst16834 (P2_U4035, P2_D_REG_27__SCAN_IN, P2_U4015);
  nand ginst16835 (P2_U4036, P2_D_REG_28__SCAN_IN, P2_U4015);
  nand ginst16836 (P2_U4037, P2_D_REG_29__SCAN_IN, P2_U4015);
  nand ginst16837 (P2_U4038, P2_D_REG_2__SCAN_IN, P2_U4015);
  nand ginst16838 (P2_U4039, P2_D_REG_30__SCAN_IN, P2_U4015);
  nand ginst16839 (P2_U4040, P2_D_REG_31__SCAN_IN, P2_U4015);
  nand ginst16840 (P2_U4041, P2_D_REG_3__SCAN_IN, P2_U4015);
  nand ginst16841 (P2_U4042, P2_D_REG_4__SCAN_IN, P2_U4015);
  nand ginst16842 (P2_U4043, P2_D_REG_5__SCAN_IN, P2_U4015);
  nand ginst16843 (P2_U4044, P2_D_REG_6__SCAN_IN, P2_U4015);
  nand ginst16844 (P2_U4045, P2_D_REG_7__SCAN_IN, P2_U4015);
  nand ginst16845 (P2_U4046, P2_D_REG_8__SCAN_IN, P2_U4015);
  nand ginst16846 (P2_U4047, P2_D_REG_9__SCAN_IN, P2_U4015);
  not ginst16847 (P2_U4048, P2_U3830);
  nand ginst16848 (P2_U4049, P2_U5446, P2_U5452);
  nand ginst16849 (P2_U4050, P2_U4049, P2_U5478);
  nand ginst16850 (P2_U4051, P2_U3367, P2_U3369);
  nand ginst16851 (P2_U4052, P2_U3890, P2_U4051);
  nand ginst16852 (P2_U4053, P2_U3891, P2_U4050);
  nand ginst16853 (P2_U4054, P2_U4052, P2_U4053);
  nand ginst16854 (P2_U4055, P2_REG0_REG_1__SCAN_IN, P2_U3022);
  nand ginst16855 (P2_U4056, P2_REG1_REG_1__SCAN_IN, P2_U3021);
  nand ginst16856 (P2_U4057, P2_REG2_REG_1__SCAN_IN, P2_U3020);
  nand ginst16857 (P2_U4058, P2_REG3_REG_1__SCAN_IN, P2_U3019);
  not ginst16858 (P2_U4059, P2_U3077);
  nand ginst16859 (P2_U4060, P2_U3357, P2_U3873);
  nand ginst16860 (P2_U4061, P2_R1110_U95, P2_U3879);
  nand ginst16861 (P2_U4062, P2_R1077_U95, P2_U3881);
  nand ginst16862 (P2_U4063, P2_R1095_U25, P2_U3880);
  nand ginst16863 (P2_U4064, P2_R1143_U95, P2_U3877);
  nand ginst16864 (P2_U4065, P2_R1161_U95, P2_U3887);
  nand ginst16865 (P2_U4066, P2_R1131_U25, P2_U3883);
  nand ginst16866 (P2_U4067, P2_R1200_U25, P2_U3017);
  not ginst16867 (P2_U4068, P2_U3314);
  nand ginst16868 (P2_U4069, P2_U3352, P2_U3829);
  nand ginst16869 (P2_U4070, P2_R1179_U25, P2_U3026);
  nand ginst16870 (P2_U4071, P2_U3025, P2_U3077);
  nand ginst16871 (P2_U4072, P2_U3387, P2_U4060);
  nand ginst16872 (P2_U4073, P2_U3577, P2_U4068);
  nand ginst16873 (P2_U4074, P2_REG0_REG_2__SCAN_IN, P2_U3022);
  nand ginst16874 (P2_U4075, P2_REG1_REG_2__SCAN_IN, P2_U3021);
  nand ginst16875 (P2_U4076, P2_REG2_REG_2__SCAN_IN, P2_U3020);
  nand ginst16876 (P2_U4077, P2_REG3_REG_2__SCAN_IN, P2_U3019);
  not ginst16877 (P2_U4078, P2_U3067);
  nand ginst16878 (P2_U4079, P2_REG0_REG_0__SCAN_IN, P2_U3022);
  nand ginst16879 (P2_U4080, P2_REG1_REG_0__SCAN_IN, P2_U3021);
  nand ginst16880 (P2_U4081, P2_REG2_REG_0__SCAN_IN, P2_U3020);
  nand ginst16881 (P2_U4082, P2_REG3_REG_0__SCAN_IN, P2_U3019);
  not ginst16882 (P2_U4083, P2_U3076);
  nand ginst16883 (P2_U4084, P2_U3383, P2_U5464);
  nand ginst16884 (P2_U4085, P2_U3892, P2_U4084);
  nand ginst16885 (P2_U4086, P2_U3033, P2_U3076);
  nand ginst16886 (P2_U4087, P2_R1110_U94, P2_U3879);
  nand ginst16887 (P2_U4088, P2_R1077_U94, P2_U3881);
  nand ginst16888 (P2_U4089, P2_R1095_U102, P2_U3880);
  nand ginst16889 (P2_U4090, P2_R1143_U94, P2_U3877);
  nand ginst16890 (P2_U4091, P2_R1161_U94, P2_U3887);
  nand ginst16891 (P2_U4092, P2_R1131_U102, P2_U3883);
  nand ginst16892 (P2_U4093, P2_R1200_U102, P2_U3017);
  not ginst16893 (P2_U4094, P2_U3315);
  nand ginst16894 (P2_U4095, P2_R1179_U102, P2_U3026);
  nand ginst16895 (P2_U4096, P2_U3025, P2_U3067);
  nand ginst16896 (P2_U4097, P2_U3392, P2_U4060);
  nand ginst16897 (P2_U4098, P2_U3593, P2_U4094);
  nand ginst16898 (P2_U4099, P2_REG0_REG_3__SCAN_IN, P2_U3022);
  nand ginst16899 (P2_U4100, P2_REG1_REG_3__SCAN_IN, P2_U3021);
  nand ginst16900 (P2_U4101, P2_REG2_REG_3__SCAN_IN, P2_U3020);
  nand ginst16901 (P2_U4102, P2_SUB_605_U26, P2_U3019);
  not ginst16902 (P2_U4103, P2_U3063);
  nand ginst16903 (P2_U4104, P2_U3033, P2_U3077);
  nand ginst16904 (P2_U4105, P2_R1110_U16, P2_U3879);
  nand ginst16905 (P2_U4106, P2_R1077_U16, P2_U3881);
  nand ginst16906 (P2_U4107, P2_R1095_U112, P2_U3880);
  nand ginst16907 (P2_U4108, P2_R1143_U16, P2_U3877);
  nand ginst16908 (P2_U4109, P2_R1161_U16, P2_U3887);
  nand ginst16909 (P2_U4110, P2_R1131_U112, P2_U3883);
  nand ginst16910 (P2_U4111, P2_R1200_U112, P2_U3017);
  not ginst16911 (P2_U4112, P2_U3316);
  nand ginst16912 (P2_U4113, P2_R1179_U112, P2_U3026);
  nand ginst16913 (P2_U4114, P2_U3025, P2_U3063);
  nand ginst16914 (P2_U4115, P2_U3395, P2_U4060);
  nand ginst16915 (P2_U4116, P2_U3597, P2_U4112);
  nand ginst16916 (P2_U4117, P2_REG0_REG_4__SCAN_IN, P2_U3022);
  nand ginst16917 (P2_U4118, P2_REG1_REG_4__SCAN_IN, P2_U3021);
  nand ginst16918 (P2_U4119, P2_REG2_REG_4__SCAN_IN, P2_U3020);
  nand ginst16919 (P2_U4120, P2_SUB_605_U30, P2_U3019);
  not ginst16920 (P2_U4121, P2_U3059);
  nand ginst16921 (P2_U4122, P2_U3033, P2_U3067);
  nand ginst16922 (P2_U4123, P2_R1110_U100, P2_U3879);
  nand ginst16923 (P2_U4124, P2_R1077_U100, P2_U3881);
  nand ginst16924 (P2_U4125, P2_R1095_U22, P2_U3880);
  nand ginst16925 (P2_U4126, P2_R1143_U100, P2_U3877);
  nand ginst16926 (P2_U4127, P2_R1161_U100, P2_U3887);
  nand ginst16927 (P2_U4128, P2_R1131_U22, P2_U3883);
  nand ginst16928 (P2_U4129, P2_R1200_U22, P2_U3017);
  not ginst16929 (P2_U4130, P2_U3317);
  nand ginst16930 (P2_U4131, P2_R1179_U22, P2_U3026);
  nand ginst16931 (P2_U4132, P2_U3025, P2_U3059);
  nand ginst16932 (P2_U4133, P2_U3398, P2_U4060);
  nand ginst16933 (P2_U4134, P2_U3601, P2_U4130);
  nand ginst16934 (P2_U4135, P2_REG0_REG_5__SCAN_IN, P2_U3022);
  nand ginst16935 (P2_U4136, P2_REG1_REG_5__SCAN_IN, P2_U3021);
  nand ginst16936 (P2_U4137, P2_REG2_REG_5__SCAN_IN, P2_U3020);
  nand ginst16937 (P2_U4138, P2_SUB_605_U22, P2_U3019);
  not ginst16938 (P2_U4139, P2_U3066);
  nand ginst16939 (P2_U4140, P2_U3033, P2_U3063);
  nand ginst16940 (P2_U4141, P2_R1110_U99, P2_U3879);
  nand ginst16941 (P2_U4142, P2_R1077_U99, P2_U3881);
  nand ginst16942 (P2_U4143, P2_R1095_U111, P2_U3880);
  nand ginst16943 (P2_U4144, P2_R1143_U99, P2_U3877);
  nand ginst16944 (P2_U4145, P2_R1161_U99, P2_U3887);
  nand ginst16945 (P2_U4146, P2_R1131_U111, P2_U3883);
  nand ginst16946 (P2_U4147, P2_R1200_U111, P2_U3017);
  not ginst16947 (P2_U4148, P2_U3318);
  nand ginst16948 (P2_U4149, P2_R1179_U111, P2_U3026);
  nand ginst16949 (P2_U4150, P2_U3025, P2_U3066);
  nand ginst16950 (P2_U4151, P2_U3401, P2_U4060);
  nand ginst16951 (P2_U4152, P2_U3605, P2_U4148);
  nand ginst16952 (P2_U4153, P2_REG0_REG_6__SCAN_IN, P2_U3022);
  nand ginst16953 (P2_U4154, P2_REG1_REG_6__SCAN_IN, P2_U3021);
  nand ginst16954 (P2_U4155, P2_REG2_REG_6__SCAN_IN, P2_U3020);
  nand ginst16955 (P2_U4156, P2_SUB_605_U8, P2_U3019);
  not ginst16956 (P2_U4157, P2_U3070);
  nand ginst16957 (P2_U4158, P2_U3033, P2_U3059);
  nand ginst16958 (P2_U4159, P2_R1110_U17, P2_U3879);
  nand ginst16959 (P2_U4160, P2_R1077_U17, P2_U3881);
  nand ginst16960 (P2_U4161, P2_R1095_U110, P2_U3880);
  nand ginst16961 (P2_U4162, P2_R1143_U17, P2_U3877);
  nand ginst16962 (P2_U4163, P2_R1161_U17, P2_U3887);
  nand ginst16963 (P2_U4164, P2_R1131_U110, P2_U3883);
  nand ginst16964 (P2_U4165, P2_R1200_U110, P2_U3017);
  not ginst16965 (P2_U4166, P2_U3319);
  nand ginst16966 (P2_U4167, P2_R1179_U110, P2_U3026);
  nand ginst16967 (P2_U4168, P2_U3025, P2_U3070);
  nand ginst16968 (P2_U4169, P2_U3404, P2_U4060);
  nand ginst16969 (P2_U4170, P2_U3609, P2_U4166);
  nand ginst16970 (P2_U4171, P2_REG0_REG_7__SCAN_IN, P2_U3022);
  nand ginst16971 (P2_U4172, P2_REG1_REG_7__SCAN_IN, P2_U3021);
  nand ginst16972 (P2_U4173, P2_REG2_REG_7__SCAN_IN, P2_U3020);
  nand ginst16973 (P2_U4174, P2_SUB_605_U18, P2_U3019);
  not ginst16974 (P2_U4175, P2_U3069);
  nand ginst16975 (P2_U4176, P2_U3033, P2_U3066);
  nand ginst16976 (P2_U4177, P2_R1110_U98, P2_U3879);
  nand ginst16977 (P2_U4178, P2_R1077_U98, P2_U3881);
  nand ginst16978 (P2_U4179, P2_R1095_U23, P2_U3880);
  nand ginst16979 (P2_U4180, P2_R1143_U98, P2_U3877);
  nand ginst16980 (P2_U4181, P2_R1161_U98, P2_U3887);
  nand ginst16981 (P2_U4182, P2_R1131_U23, P2_U3883);
  nand ginst16982 (P2_U4183, P2_R1200_U23, P2_U3017);
  not ginst16983 (P2_U4184, P2_U3320);
  nand ginst16984 (P2_U4185, P2_R1179_U23, P2_U3026);
  nand ginst16985 (P2_U4186, P2_U3025, P2_U3069);
  nand ginst16986 (P2_U4187, P2_U3407, P2_U4060);
  nand ginst16987 (P2_U4188, P2_U3613, P2_U4184);
  nand ginst16988 (P2_U4189, P2_REG0_REG_8__SCAN_IN, P2_U3022);
  nand ginst16989 (P2_U4190, P2_REG1_REG_8__SCAN_IN, P2_U3021);
  nand ginst16990 (P2_U4191, P2_REG2_REG_8__SCAN_IN, P2_U3020);
  nand ginst16991 (P2_U4192, P2_SUB_605_U12, P2_U3019);
  not ginst16992 (P2_U4193, P2_U3083);
  nand ginst16993 (P2_U4194, P2_U3033, P2_U3070);
  nand ginst16994 (P2_U4195, P2_R1110_U18, P2_U3879);
  nand ginst16995 (P2_U4196, P2_R1077_U18, P2_U3881);
  nand ginst16996 (P2_U4197, P2_R1095_U109, P2_U3880);
  nand ginst16997 (P2_U4198, P2_R1143_U18, P2_U3877);
  nand ginst16998 (P2_U4199, P2_R1161_U18, P2_U3887);
  nand ginst16999 (P2_U4200, P2_R1131_U109, P2_U3883);
  nand ginst17000 (P2_U4201, P2_R1200_U109, P2_U3017);
  not ginst17001 (P2_U4202, P2_U3321);
  nand ginst17002 (P2_U4203, P2_R1179_U109, P2_U3026);
  nand ginst17003 (P2_U4204, P2_U3025, P2_U3083);
  nand ginst17004 (P2_U4205, P2_U3410, P2_U4060);
  nand ginst17005 (P2_U4206, P2_U3617, P2_U4202);
  nand ginst17006 (P2_U4207, P2_REG0_REG_9__SCAN_IN, P2_U3022);
  nand ginst17007 (P2_U4208, P2_REG1_REG_9__SCAN_IN, P2_U3021);
  nand ginst17008 (P2_U4209, P2_REG2_REG_9__SCAN_IN, P2_U3020);
  nand ginst17009 (P2_U4210, P2_SUB_605_U14, P2_U3019);
  not ginst17010 (P2_U4211, P2_U3082);
  nand ginst17011 (P2_U4212, P2_U3033, P2_U3069);
  nand ginst17012 (P2_U4213, P2_R1110_U97, P2_U3879);
  nand ginst17013 (P2_U4214, P2_R1077_U97, P2_U3881);
  nand ginst17014 (P2_U4215, P2_R1095_U24, P2_U3880);
  nand ginst17015 (P2_U4216, P2_R1143_U97, P2_U3877);
  nand ginst17016 (P2_U4217, P2_R1161_U97, P2_U3887);
  nand ginst17017 (P2_U4218, P2_R1131_U24, P2_U3883);
  nand ginst17018 (P2_U4219, P2_R1200_U24, P2_U3017);
  not ginst17019 (P2_U4220, P2_U3322);
  nand ginst17020 (P2_U4221, P2_R1179_U24, P2_U3026);
  nand ginst17021 (P2_U4222, P2_U3025, P2_U3082);
  nand ginst17022 (P2_U4223, P2_U3413, P2_U4060);
  nand ginst17023 (P2_U4224, P2_U3620, P2_U4220);
  nand ginst17024 (P2_U4225, P2_REG0_REG_10__SCAN_IN, P2_U3022);
  nand ginst17025 (P2_U4226, P2_REG1_REG_10__SCAN_IN, P2_U3021);
  nand ginst17026 (P2_U4227, P2_REG2_REG_10__SCAN_IN, P2_U3020);
  nand ginst17027 (P2_U4228, P2_SUB_605_U13, P2_U3019);
  not ginst17028 (P2_U4229, P2_U3061);
  nand ginst17029 (P2_U4230, P2_U3033, P2_U3083);
  nand ginst17030 (P2_U4231, P2_R1110_U96, P2_U3879);
  nand ginst17031 (P2_U4232, P2_R1077_U96, P2_U3881);
  nand ginst17032 (P2_U4233, P2_R1095_U108, P2_U3880);
  nand ginst17033 (P2_U4234, P2_R1143_U96, P2_U3877);
  nand ginst17034 (P2_U4235, P2_R1161_U96, P2_U3887);
  nand ginst17035 (P2_U4236, P2_R1131_U108, P2_U3883);
  nand ginst17036 (P2_U4237, P2_R1200_U108, P2_U3017);
  not ginst17037 (P2_U4238, P2_U3323);
  nand ginst17038 (P2_U4239, P2_R1179_U108, P2_U3026);
  nand ginst17039 (P2_U4240, P2_U3025, P2_U3061);
  nand ginst17040 (P2_U4241, P2_U3416, P2_U4060);
  nand ginst17041 (P2_U4242, P2_U3623, P2_U4238);
  nand ginst17042 (P2_U4243, P2_REG0_REG_11__SCAN_IN, P2_U3022);
  nand ginst17043 (P2_U4244, P2_REG1_REG_11__SCAN_IN, P2_U3021);
  nand ginst17044 (P2_U4245, P2_REG2_REG_11__SCAN_IN, P2_U3020);
  nand ginst17045 (P2_U4246, P2_SUB_605_U9, P2_U3019);
  not ginst17046 (P2_U4247, P2_U3062);
  nand ginst17047 (P2_U4248, P2_U3033, P2_U3082);
  nand ginst17048 (P2_U4249, P2_R1110_U10, P2_U3879);
  nand ginst17049 (P2_U4250, P2_R1077_U10, P2_U3881);
  nand ginst17050 (P2_U4251, P2_R1095_U118, P2_U3880);
  nand ginst17051 (P2_U4252, P2_R1143_U10, P2_U3877);
  nand ginst17052 (P2_U4253, P2_R1161_U10, P2_U3887);
  nand ginst17053 (P2_U4254, P2_R1131_U118, P2_U3883);
  nand ginst17054 (P2_U4255, P2_R1200_U118, P2_U3017);
  not ginst17055 (P2_U4256, P2_U3324);
  nand ginst17056 (P2_U4257, P2_R1179_U118, P2_U3026);
  nand ginst17057 (P2_U4258, P2_U3025, P2_U3062);
  nand ginst17058 (P2_U4259, P2_U3419, P2_U4060);
  nand ginst17059 (P2_U4260, P2_U3626, P2_U4256);
  nand ginst17060 (P2_U4261, P2_REG0_REG_12__SCAN_IN, P2_U3022);
  nand ginst17061 (P2_U4262, P2_REG1_REG_12__SCAN_IN, P2_U3021);
  nand ginst17062 (P2_U4263, P2_REG2_REG_12__SCAN_IN, P2_U3020);
  nand ginst17063 (P2_U4264, P2_SUB_605_U24, P2_U3019);
  not ginst17064 (P2_U4265, P2_U3071);
  nand ginst17065 (P2_U4266, P2_U3033, P2_U3061);
  nand ginst17066 (P2_U4267, P2_R1110_U114, P2_U3879);
  nand ginst17067 (P2_U4268, P2_R1077_U114, P2_U3881);
  nand ginst17068 (P2_U4269, P2_R1095_U17, P2_U3880);
  nand ginst17069 (P2_U4270, P2_R1143_U114, P2_U3877);
  nand ginst17070 (P2_U4271, P2_R1161_U114, P2_U3887);
  nand ginst17071 (P2_U4272, P2_R1131_U17, P2_U3883);
  nand ginst17072 (P2_U4273, P2_R1200_U17, P2_U3017);
  not ginst17073 (P2_U4274, P2_U3325);
  nand ginst17074 (P2_U4275, P2_R1179_U17, P2_U3026);
  nand ginst17075 (P2_U4276, P2_U3025, P2_U3071);
  nand ginst17076 (P2_U4277, P2_U3422, P2_U4060);
  nand ginst17077 (P2_U4278, P2_U3629, P2_U4274);
  nand ginst17078 (P2_U4279, P2_REG0_REG_13__SCAN_IN, P2_U3022);
  nand ginst17079 (P2_U4280, P2_REG1_REG_13__SCAN_IN, P2_U3021);
  nand ginst17080 (P2_U4281, P2_REG2_REG_13__SCAN_IN, P2_U3020);
  nand ginst17081 (P2_U4282, P2_SUB_605_U25, P2_U3019);
  not ginst17082 (P2_U4283, P2_U3079);
  nand ginst17083 (P2_U4284, P2_U3033, P2_U3062);
  nand ginst17084 (P2_U4285, P2_R1110_U113, P2_U3879);
  nand ginst17085 (P2_U4286, P2_R1077_U113, P2_U3881);
  nand ginst17086 (P2_U4287, P2_R1095_U107, P2_U3880);
  nand ginst17087 (P2_U4288, P2_R1143_U113, P2_U3877);
  nand ginst17088 (P2_U4289, P2_R1161_U113, P2_U3887);
  nand ginst17089 (P2_U4290, P2_R1131_U107, P2_U3883);
  nand ginst17090 (P2_U4291, P2_R1200_U107, P2_U3017);
  not ginst17091 (P2_U4292, P2_U3326);
  nand ginst17092 (P2_U4293, P2_R1179_U107, P2_U3026);
  nand ginst17093 (P2_U4294, P2_U3025, P2_U3079);
  nand ginst17094 (P2_U4295, P2_U3425, P2_U4060);
  nand ginst17095 (P2_U4296, P2_U3633, P2_U4292);
  nand ginst17096 (P2_U4297, P2_REG0_REG_14__SCAN_IN, P2_U3022);
  nand ginst17097 (P2_U4298, P2_REG1_REG_14__SCAN_IN, P2_U3021);
  nand ginst17098 (P2_U4299, P2_REG2_REG_14__SCAN_IN, P2_U3020);
  nand ginst17099 (P2_U4300, P2_SUB_605_U31, P2_U3019);
  not ginst17100 (P2_U4301, P2_U3078);
  nand ginst17101 (P2_U4302, P2_U3033, P2_U3071);
  nand ginst17102 (P2_U4303, P2_R1110_U11, P2_U3879);
  nand ginst17103 (P2_U4304, P2_R1077_U11, P2_U3881);
  nand ginst17104 (P2_U4305, P2_R1095_U106, P2_U3880);
  nand ginst17105 (P2_U4306, P2_R1143_U11, P2_U3877);
  nand ginst17106 (P2_U4307, P2_R1161_U11, P2_U3887);
  nand ginst17107 (P2_U4308, P2_R1131_U106, P2_U3883);
  nand ginst17108 (P2_U4309, P2_R1200_U106, P2_U3017);
  not ginst17109 (P2_U4310, P2_U3327);
  nand ginst17110 (P2_U4311, P2_R1179_U106, P2_U3026);
  nand ginst17111 (P2_U4312, P2_U3025, P2_U3078);
  nand ginst17112 (P2_U4313, P2_U3428, P2_U4060);
  nand ginst17113 (P2_U4314, P2_U3637, P2_U4310);
  nand ginst17114 (P2_U4315, P2_REG0_REG_15__SCAN_IN, P2_U3022);
  nand ginst17115 (P2_U4316, P2_REG1_REG_15__SCAN_IN, P2_U3021);
  nand ginst17116 (P2_U4317, P2_REG2_REG_15__SCAN_IN, P2_U3020);
  nand ginst17117 (P2_U4318, P2_SUB_605_U21, P2_U3019);
  not ginst17118 (P2_U4319, P2_U3073);
  nand ginst17119 (P2_U4320, P2_U3033, P2_U3079);
  nand ginst17120 (P2_U4321, P2_R1110_U112, P2_U3879);
  nand ginst17121 (P2_U4322, P2_R1077_U112, P2_U3881);
  nand ginst17122 (P2_U4323, P2_R1095_U117, P2_U3880);
  nand ginst17123 (P2_U4324, P2_R1143_U112, P2_U3877);
  nand ginst17124 (P2_U4325, P2_R1161_U112, P2_U3887);
  nand ginst17125 (P2_U4326, P2_R1131_U117, P2_U3883);
  nand ginst17126 (P2_U4327, P2_R1200_U117, P2_U3017);
  not ginst17127 (P2_U4328, P2_U3328);
  nand ginst17128 (P2_U4329, P2_R1179_U117, P2_U3026);
  nand ginst17129 (P2_U4330, P2_U3025, P2_U3073);
  nand ginst17130 (P2_U4331, P2_U3431, P2_U4060);
  nand ginst17131 (P2_U4332, P2_U3640, P2_U4328);
  nand ginst17132 (P2_U4333, P2_REG0_REG_16__SCAN_IN, P2_U3022);
  nand ginst17133 (P2_U4334, P2_REG1_REG_16__SCAN_IN, P2_U3021);
  nand ginst17134 (P2_U4335, P2_REG2_REG_16__SCAN_IN, P2_U3020);
  nand ginst17135 (P2_U4336, P2_SUB_605_U7, P2_U3019);
  not ginst17136 (P2_U4337, P2_U3072);
  nand ginst17137 (P2_U4338, P2_U3033, P2_U3078);
  nand ginst17138 (P2_U4339, P2_R1110_U111, P2_U3879);
  nand ginst17139 (P2_U4340, P2_R1077_U111, P2_U3881);
  nand ginst17140 (P2_U4341, P2_R1095_U116, P2_U3880);
  nand ginst17141 (P2_U4342, P2_R1143_U111, P2_U3877);
  nand ginst17142 (P2_U4343, P2_R1161_U111, P2_U3887);
  nand ginst17143 (P2_U4344, P2_R1131_U116, P2_U3883);
  nand ginst17144 (P2_U4345, P2_R1200_U116, P2_U3017);
  not ginst17145 (P2_U4346, P2_U3329);
  nand ginst17146 (P2_U4347, P2_R1179_U116, P2_U3026);
  nand ginst17147 (P2_U4348, P2_U3025, P2_U3072);
  nand ginst17148 (P2_U4349, P2_U3434, P2_U4060);
  nand ginst17149 (P2_U4350, P2_U3643, P2_U4346);
  nand ginst17150 (P2_U4351, P2_REG0_REG_17__SCAN_IN, P2_U3022);
  nand ginst17151 (P2_U4352, P2_REG1_REG_17__SCAN_IN, P2_U3021);
  nand ginst17152 (P2_U4353, P2_REG2_REG_17__SCAN_IN, P2_U3020);
  nand ginst17153 (P2_U4354, P2_SUB_605_U19, P2_U3019);
  not ginst17154 (P2_U4355, P2_U3068);
  nand ginst17155 (P2_U4356, P2_U3033, P2_U3073);
  nand ginst17156 (P2_U4357, P2_R1110_U110, P2_U3879);
  nand ginst17157 (P2_U4358, P2_R1077_U110, P2_U3881);
  nand ginst17158 (P2_U4359, P2_R1095_U18, P2_U3880);
  nand ginst17159 (P2_U4360, P2_R1143_U110, P2_U3877);
  nand ginst17160 (P2_U4361, P2_R1161_U110, P2_U3887);
  nand ginst17161 (P2_U4362, P2_R1131_U18, P2_U3883);
  nand ginst17162 (P2_U4363, P2_R1200_U18, P2_U3017);
  not ginst17163 (P2_U4364, P2_U3330);
  nand ginst17164 (P2_U4365, P2_R1179_U18, P2_U3026);
  nand ginst17165 (P2_U4366, P2_U3025, P2_U3068);
  nand ginst17166 (P2_U4367, P2_U3437, P2_U4060);
  nand ginst17167 (P2_U4368, P2_U3646, P2_U4364);
  nand ginst17168 (P2_U4369, P2_REG0_REG_18__SCAN_IN, P2_U3022);
  nand ginst17169 (P2_U4370, P2_REG1_REG_18__SCAN_IN, P2_U3021);
  nand ginst17170 (P2_U4371, P2_REG2_REG_18__SCAN_IN, P2_U3020);
  nand ginst17171 (P2_U4372, P2_SUB_605_U11, P2_U3019);
  not ginst17172 (P2_U4373, P2_U3081);
  nand ginst17173 (P2_U4374, P2_U3033, P2_U3072);
  nand ginst17174 (P2_U4375, P2_R1110_U12, P2_U3879);
  nand ginst17175 (P2_U4376, P2_R1077_U12, P2_U3881);
  nand ginst17176 (P2_U4377, P2_R1095_U105, P2_U3880);
  nand ginst17177 (P2_U4378, P2_R1143_U12, P2_U3877);
  nand ginst17178 (P2_U4379, P2_R1161_U12, P2_U3887);
  nand ginst17179 (P2_U4380, P2_R1131_U105, P2_U3883);
  nand ginst17180 (P2_U4381, P2_R1200_U105, P2_U3017);
  not ginst17181 (P2_U4382, P2_U3331);
  nand ginst17182 (P2_U4383, P2_R1179_U105, P2_U3026);
  nand ginst17183 (P2_U4384, P2_U3025, P2_U3081);
  nand ginst17184 (P2_U4385, P2_U3440, P2_U4060);
  nand ginst17185 (P2_U4386, P2_U3650, P2_U4382);
  nand ginst17186 (P2_U4387, P2_REG0_REG_19__SCAN_IN, P2_U3022);
  nand ginst17187 (P2_U4388, P2_REG1_REG_19__SCAN_IN, P2_U3021);
  nand ginst17188 (P2_U4389, P2_REG2_REG_19__SCAN_IN, P2_U3020);
  nand ginst17189 (P2_U4390, P2_SUB_605_U15, P2_U3019);
  not ginst17190 (P2_U4391, P2_U3080);
  nand ginst17191 (P2_U4392, P2_U3033, P2_U3068);
  nand ginst17192 (P2_U4393, P2_R1110_U109, P2_U3879);
  nand ginst17193 (P2_U4394, P2_R1077_U109, P2_U3881);
  nand ginst17194 (P2_U4395, P2_R1095_U104, P2_U3880);
  nand ginst17195 (P2_U4396, P2_R1143_U109, P2_U3877);
  nand ginst17196 (P2_U4397, P2_R1161_U109, P2_U3887);
  nand ginst17197 (P2_U4398, P2_R1131_U104, P2_U3883);
  nand ginst17198 (P2_U4399, P2_R1200_U104, P2_U3017);
  not ginst17199 (P2_U4400, P2_U3332);
  nand ginst17200 (P2_U4401, P2_R1179_U104, P2_U3026);
  nand ginst17201 (P2_U4402, P2_U3025, P2_U3080);
  nand ginst17202 (P2_U4403, P2_U3443, P2_U4060);
  nand ginst17203 (P2_U4404, P2_U3654, P2_U4400);
  nand ginst17204 (P2_U4405, P2_REG2_REG_20__SCAN_IN, P2_U3020);
  nand ginst17205 (P2_U4406, P2_REG1_REG_20__SCAN_IN, P2_U3021);
  nand ginst17206 (P2_U4407, P2_REG0_REG_20__SCAN_IN, P2_U3022);
  nand ginst17207 (P2_U4408, P2_SUB_605_U20, P2_U3019);
  not ginst17208 (P2_U4409, P2_U3075);
  nand ginst17209 (P2_U4410, P2_U3033, P2_U3081);
  nand ginst17210 (P2_U4411, P2_R1110_U108, P2_U3879);
  nand ginst17211 (P2_U4412, P2_R1077_U108, P2_U3881);
  nand ginst17212 (P2_U4413, P2_R1095_U103, P2_U3880);
  nand ginst17213 (P2_U4414, P2_R1143_U108, P2_U3877);
  nand ginst17214 (P2_U4415, P2_R1161_U108, P2_U3887);
  nand ginst17215 (P2_U4416, P2_R1131_U103, P2_U3883);
  nand ginst17216 (P2_U4417, P2_R1200_U103, P2_U3017);
  not ginst17217 (P2_U4418, P2_U3333);
  nand ginst17218 (P2_U4419, P2_R1179_U103, P2_U3026);
  nand ginst17219 (P2_U4420, P2_U3025, P2_U3075);
  nand ginst17220 (P2_U4421, P2_U3445, P2_U4060);
  nand ginst17221 (P2_U4422, P2_U3658, P2_U4418);
  nand ginst17222 (P2_U4423, P2_REG2_REG_21__SCAN_IN, P2_U3020);
  nand ginst17223 (P2_U4424, P2_REG1_REG_21__SCAN_IN, P2_U3021);
  nand ginst17224 (P2_U4425, P2_REG0_REG_21__SCAN_IN, P2_U3022);
  nand ginst17225 (P2_U4426, P2_SUB_605_U28, P2_U3019);
  not ginst17226 (P2_U4427, P2_U3074);
  nand ginst17227 (P2_U4428, P2_U3033, P2_U3080);
  nand ginst17228 (P2_U4429, P2_R1110_U13, P2_U3879);
  nand ginst17229 (P2_U4430, P2_R1077_U13, P2_U3881);
  nand ginst17230 (P2_U4431, P2_R1095_U101, P2_U3880);
  nand ginst17231 (P2_U4432, P2_R1143_U13, P2_U3877);
  nand ginst17232 (P2_U4433, P2_R1161_U13, P2_U3887);
  nand ginst17233 (P2_U4434, P2_R1131_U101, P2_U3883);
  nand ginst17234 (P2_U4435, P2_R1200_U101, P2_U3017);
  not ginst17235 (P2_U4436, P2_U3335);
  nand ginst17236 (P2_U4437, P2_R1179_U101, P2_U3026);
  nand ginst17237 (P2_U4438, P2_U3025, P2_U3074);
  nand ginst17238 (P2_U4439, P2_U3903, P2_U4060);
  nand ginst17239 (P2_U4440, P2_U3662, P2_U4436);
  nand ginst17240 (P2_U4441, P2_REG2_REG_22__SCAN_IN, P2_U3020);
  nand ginst17241 (P2_U4442, P2_REG1_REG_22__SCAN_IN, P2_U3021);
  nand ginst17242 (P2_U4443, P2_REG0_REG_22__SCAN_IN, P2_U3022);
  nand ginst17243 (P2_U4444, P2_SUB_605_U17, P2_U3019);
  not ginst17244 (P2_U4445, P2_U3060);
  nand ginst17245 (P2_U4446, P2_U3033, P2_U3075);
  nand ginst17246 (P2_U4447, P2_R1110_U14, P2_U3879);
  nand ginst17247 (P2_U4448, P2_R1077_U14, P2_U3881);
  nand ginst17248 (P2_U4449, P2_R1095_U115, P2_U3880);
  nand ginst17249 (P2_U4450, P2_R1143_U14, P2_U3877);
  nand ginst17250 (P2_U4451, P2_R1161_U14, P2_U3887);
  nand ginst17251 (P2_U4452, P2_R1131_U115, P2_U3883);
  nand ginst17252 (P2_U4453, P2_R1200_U115, P2_U3017);
  not ginst17253 (P2_U4454, P2_U3337);
  nand ginst17254 (P2_U4455, P2_R1179_U115, P2_U3026);
  nand ginst17255 (P2_U4456, P2_U3025, P2_U3060);
  nand ginst17256 (P2_U4457, P2_U3902, P2_U4060);
  nand ginst17257 (P2_U4458, P2_U3665, P2_U4454);
  nand ginst17258 (P2_U4459, P2_REG2_REG_23__SCAN_IN, P2_U3020);
  nand ginst17259 (P2_U4460, P2_REG1_REG_23__SCAN_IN, P2_U3021);
  nand ginst17260 (P2_U4461, P2_REG0_REG_23__SCAN_IN, P2_U3022);
  nand ginst17261 (P2_U4462, P2_SUB_605_U6, P2_U3019);
  not ginst17262 (P2_U4463, P2_U3065);
  nand ginst17263 (P2_U4464, P2_U3033, P2_U3074);
  nand ginst17264 (P2_U4465, P2_R1110_U107, P2_U3879);
  nand ginst17265 (P2_U4466, P2_R1077_U107, P2_U3881);
  nand ginst17266 (P2_U4467, P2_R1095_U114, P2_U3880);
  nand ginst17267 (P2_U4468, P2_R1143_U107, P2_U3877);
  nand ginst17268 (P2_U4469, P2_R1161_U107, P2_U3887);
  nand ginst17269 (P2_U4470, P2_R1131_U114, P2_U3883);
  nand ginst17270 (P2_U4471, P2_R1200_U114, P2_U3017);
  not ginst17271 (P2_U4472, P2_U3339);
  nand ginst17272 (P2_U4473, P2_R1179_U114, P2_U3026);
  nand ginst17273 (P2_U4474, P2_U3025, P2_U3065);
  nand ginst17274 (P2_U4475, P2_U3901, P2_U4060);
  nand ginst17275 (P2_U4476, P2_U3668, P2_U4472);
  nand ginst17276 (P2_U4477, P2_REG2_REG_24__SCAN_IN, P2_U3020);
  nand ginst17277 (P2_U4478, P2_REG1_REG_24__SCAN_IN, P2_U3021);
  nand ginst17278 (P2_U4479, P2_REG0_REG_24__SCAN_IN, P2_U3022);
  nand ginst17279 (P2_U4480, P2_SUB_605_U10, P2_U3019);
  not ginst17280 (P2_U4481, P2_U3064);
  nand ginst17281 (P2_U4482, P2_U3033, P2_U3060);
  nand ginst17282 (P2_U4483, P2_R1110_U106, P2_U3879);
  nand ginst17283 (P2_U4484, P2_R1077_U106, P2_U3881);
  nand ginst17284 (P2_U4485, P2_R1095_U19, P2_U3880);
  nand ginst17285 (P2_U4486, P2_R1143_U106, P2_U3877);
  nand ginst17286 (P2_U4487, P2_R1161_U106, P2_U3887);
  nand ginst17287 (P2_U4488, P2_R1131_U19, P2_U3883);
  nand ginst17288 (P2_U4489, P2_R1200_U19, P2_U3017);
  not ginst17289 (P2_U4490, P2_U3341);
  nand ginst17290 (P2_U4491, P2_R1179_U19, P2_U3026);
  nand ginst17291 (P2_U4492, P2_U3025, P2_U3064);
  nand ginst17292 (P2_U4493, P2_U3900, P2_U4060);
  nand ginst17293 (P2_U4494, P2_U3671, P2_U4490);
  nand ginst17294 (P2_U4495, P2_REG2_REG_25__SCAN_IN, P2_U3020);
  nand ginst17295 (P2_U4496, P2_REG1_REG_25__SCAN_IN, P2_U3021);
  nand ginst17296 (P2_U4497, P2_REG0_REG_25__SCAN_IN, P2_U3022);
  nand ginst17297 (P2_U4498, P2_SUB_605_U16, P2_U3019);
  not ginst17298 (P2_U4499, P2_U3057);
  nand ginst17299 (P2_U4500, P2_U3033, P2_U3065);
  nand ginst17300 (P2_U4501, P2_R1110_U105, P2_U3879);
  nand ginst17301 (P2_U4502, P2_R1077_U105, P2_U3881);
  nand ginst17302 (P2_U4503, P2_R1095_U100, P2_U3880);
  nand ginst17303 (P2_U4504, P2_R1143_U105, P2_U3877);
  nand ginst17304 (P2_U4505, P2_R1161_U105, P2_U3887);
  nand ginst17305 (P2_U4506, P2_R1131_U100, P2_U3883);
  nand ginst17306 (P2_U4507, P2_R1200_U100, P2_U3017);
  not ginst17307 (P2_U4508, P2_U3343);
  nand ginst17308 (P2_U4509, P2_R1179_U100, P2_U3026);
  nand ginst17309 (P2_U4510, P2_U3025, P2_U3057);
  nand ginst17310 (P2_U4511, P2_U3899, P2_U4060);
  nand ginst17311 (P2_U4512, P2_U3675, P2_U4508);
  nand ginst17312 (P2_U4513, P2_REG2_REG_26__SCAN_IN, P2_U3020);
  nand ginst17313 (P2_U4514, P2_REG1_REG_26__SCAN_IN, P2_U3021);
  nand ginst17314 (P2_U4515, P2_REG0_REG_26__SCAN_IN, P2_U3022);
  nand ginst17315 (P2_U4516, P2_SUB_605_U27, P2_U3019);
  not ginst17316 (P2_U4517, P2_U3056);
  nand ginst17317 (P2_U4518, P2_U3033, P2_U3064);
  nand ginst17318 (P2_U4519, P2_R1110_U104, P2_U3879);
  nand ginst17319 (P2_U4520, P2_R1077_U104, P2_U3881);
  nand ginst17320 (P2_U4521, P2_R1095_U99, P2_U3880);
  nand ginst17321 (P2_U4522, P2_R1143_U104, P2_U3877);
  nand ginst17322 (P2_U4523, P2_R1161_U104, P2_U3887);
  nand ginst17323 (P2_U4524, P2_R1131_U99, P2_U3883);
  nand ginst17324 (P2_U4525, P2_R1200_U99, P2_U3017);
  not ginst17325 (P2_U4526, P2_U3345);
  nand ginst17326 (P2_U4527, P2_R1179_U99, P2_U3026);
  nand ginst17327 (P2_U4528, P2_U3025, P2_U3056);
  nand ginst17328 (P2_U4529, P2_U3898, P2_U4060);
  nand ginst17329 (P2_U4530, P2_U3679, P2_U4526);
  nand ginst17330 (P2_U4531, P2_REG2_REG_27__SCAN_IN, P2_U3020);
  nand ginst17331 (P2_U4532, P2_REG1_REG_27__SCAN_IN, P2_U3021);
  nand ginst17332 (P2_U4533, P2_REG0_REG_27__SCAN_IN, P2_U3022);
  nand ginst17333 (P2_U4534, P2_SUB_605_U23, P2_U3019);
  not ginst17334 (P2_U4535, P2_U3052);
  nand ginst17335 (P2_U4536, P2_U3033, P2_U3057);
  nand ginst17336 (P2_U4537, P2_R1110_U15, P2_U3879);
  nand ginst17337 (P2_U4538, P2_R1077_U15, P2_U3881);
  nand ginst17338 (P2_U4539, P2_R1095_U113, P2_U3880);
  nand ginst17339 (P2_U4540, P2_R1143_U15, P2_U3877);
  nand ginst17340 (P2_U4541, P2_R1161_U15, P2_U3887);
  nand ginst17341 (P2_U4542, P2_R1131_U113, P2_U3883);
  nand ginst17342 (P2_U4543, P2_R1200_U113, P2_U3017);
  not ginst17343 (P2_U4544, P2_U3347);
  nand ginst17344 (P2_U4545, P2_R1179_U113, P2_U3026);
  nand ginst17345 (P2_U4546, P2_U3025, P2_U3052);
  nand ginst17346 (P2_U4547, P2_U3897, P2_U4060);
  nand ginst17347 (P2_U4548, P2_U3683, P2_U4544);
  nand ginst17348 (P2_U4549, P2_REG2_REG_28__SCAN_IN, P2_U3020);
  nand ginst17349 (P2_U4550, P2_REG1_REG_28__SCAN_IN, P2_U3021);
  nand ginst17350 (P2_U4551, P2_REG0_REG_28__SCAN_IN, P2_U3022);
  nand ginst17351 (P2_U4552, P2_SUB_605_U29, P2_U3019);
  not ginst17352 (P2_U4553, P2_U3053);
  nand ginst17353 (P2_U4554, P2_U3033, P2_U3056);
  nand ginst17354 (P2_U4555, P2_R1110_U103, P2_U3879);
  nand ginst17355 (P2_U4556, P2_R1077_U103, P2_U3881);
  nand ginst17356 (P2_U4557, P2_R1095_U20, P2_U3880);
  nand ginst17357 (P2_U4558, P2_R1143_U103, P2_U3877);
  nand ginst17358 (P2_U4559, P2_R1161_U103, P2_U3887);
  nand ginst17359 (P2_U4560, P2_R1131_U20, P2_U3883);
  nand ginst17360 (P2_U4561, P2_R1200_U20, P2_U3017);
  not ginst17361 (P2_U4562, P2_U3349);
  nand ginst17362 (P2_U4563, P2_R1179_U20, P2_U3026);
  nand ginst17363 (P2_U4564, P2_U3025, P2_U3053);
  nand ginst17364 (P2_U4565, P2_U3896, P2_U4060);
  nand ginst17365 (P2_U4566, P2_U3687, P2_U4562);
  nand ginst17366 (P2_U4567, P2_SUB_605_U94, P2_U3019);
  nand ginst17367 (P2_U4568, P2_REG2_REG_29__SCAN_IN, P2_U3020);
  nand ginst17368 (P2_U4569, P2_REG1_REG_29__SCAN_IN, P2_U3021);
  nand ginst17369 (P2_U4570, P2_REG0_REG_29__SCAN_IN, P2_U3022);
  not ginst17370 (P2_U4571, P2_U3054);
  nand ginst17371 (P2_U4572, P2_U3033, P2_U3052);
  nand ginst17372 (P2_U4573, P2_R1110_U102, P2_U3879);
  nand ginst17373 (P2_U4574, P2_R1077_U102, P2_U3881);
  nand ginst17374 (P2_U4575, P2_R1095_U98, P2_U3880);
  nand ginst17375 (P2_U4576, P2_R1143_U102, P2_U3877);
  nand ginst17376 (P2_U4577, P2_R1161_U102, P2_U3887);
  nand ginst17377 (P2_U4578, P2_R1131_U98, P2_U3883);
  nand ginst17378 (P2_U4579, P2_R1200_U98, P2_U3017);
  not ginst17379 (P2_U4580, P2_U3351);
  nand ginst17380 (P2_U4581, P2_R1179_U98, P2_U3026);
  nand ginst17381 (P2_U4582, P2_U3025, P2_U3054);
  nand ginst17382 (P2_U4583, P2_U3895, P2_U4060);
  nand ginst17383 (P2_U4584, P2_U3691, P2_U4580);
  nand ginst17384 (P2_U4585, P2_REG2_REG_30__SCAN_IN, P2_U3020);
  nand ginst17385 (P2_U4586, P2_REG1_REG_30__SCAN_IN, P2_U3021);
  nand ginst17386 (P2_U4587, P2_REG0_REG_30__SCAN_IN, P2_U3022);
  nand ginst17387 (P2_U4588, P2_SUB_605_U94, P2_U3019);
  not ginst17388 (P2_U4589, P2_U3058);
  nand ginst17389 (P2_U4590, P2_U3298, P2_U3888);
  nand ginst17390 (P2_U4591, P2_U3829, P2_U4590);
  nand ginst17391 (P2_U4592, P2_U3058, P2_U3907, P2_U4591);
  nand ginst17392 (P2_U4593, P2_U3033, P2_U3053);
  nand ginst17393 (P2_U4594, P2_R1110_U101, P2_U3879);
  nand ginst17394 (P2_U4595, P2_R1077_U101, P2_U3881);
  nand ginst17395 (P2_U4596, P2_R1095_U21, P2_U3880);
  nand ginst17396 (P2_U4597, P2_R1143_U101, P2_U3877);
  nand ginst17397 (P2_U4598, P2_R1161_U101, P2_U3887);
  nand ginst17398 (P2_U4599, P2_R1131_U21, P2_U3883);
  nand ginst17399 (P2_U4600, P2_R1200_U21, P2_U3017);
  not ginst17400 (P2_U4601, P2_U3354);
  nand ginst17401 (P2_U4602, P2_R1179_U21, P2_U3026);
  nand ginst17402 (P2_U4603, P2_U3904, P2_U4060);
  nand ginst17403 (P2_U4604, P2_U3695, P2_U4601);
  nand ginst17404 (P2_U4605, P2_SUB_605_U94, P2_U3019);
  nand ginst17405 (P2_U4606, P2_REG2_REG_31__SCAN_IN, P2_U3020);
  nand ginst17406 (P2_U4607, P2_REG1_REG_31__SCAN_IN, P2_U3021);
  nand ginst17407 (P2_U4608, P2_REG0_REG_31__SCAN_IN, P2_U3022);
  not ginst17408 (P2_U4609, P2_U3055);
  nand ginst17409 (P2_U4610, P2_U3869, P2_U4060);
  nand ginst17410 (P2_U4611, P2_U3361, P2_U4610);
  nand ginst17411 (P2_U4612, P2_U3868, P2_U4060);
  nand ginst17412 (P2_U4613, P2_U3361, P2_U4612);
  nand ginst17413 (P2_U4614, P2_U3302, P2_U5636, P2_U5637);
  nand ginst17414 (P2_U4615, P2_U3367, P2_U3884);
  nand ginst17415 (P2_U4616, P2_U3048, P2_U4615);
  nand ginst17416 (P2_U4617, P2_U3047, P2_U4614);
  nand ginst17417 (P2_U4618, P2_U4616, P2_U4617);
  nand ginst17418 (P2_U4619, P2_U3379, P2_U5452);
  nand ginst17419 (P2_U4620, P2_U3380, P2_U3830, P2_U4619);
  nand ginst17420 (P2_U4621, P2_U3048, P2_U4620);
  nand ginst17421 (P2_U4622, P2_U3047, P2_U4615);
  nand ginst17422 (P2_U4623, P2_U3360, P2_U4621, P2_U4622);
  not ginst17423 (P2_U4624, P2_U3365);
  nand ginst17424 (P2_U4625, P2_U3034, P2_U3077);
  nand ginst17425 (P2_U4626, P2_R1179_U25, P2_U3030);
  nand ginst17426 (P2_U4627, P2_U3029, P2_U3387);
  nand ginst17427 (P2_U4628, P2_REG3_REG_0__SCAN_IN, P2_U3028);
  nand ginst17428 (P2_U4629, P2_U3034, P2_U3067);
  nand ginst17429 (P2_U4630, P2_R1179_U102, P2_U3030);
  nand ginst17430 (P2_U4631, P2_U3029, P2_U3392);
  nand ginst17431 (P2_U4632, P2_REG3_REG_1__SCAN_IN, P2_U3028);
  nand ginst17432 (P2_U4633, P2_U3034, P2_U3063);
  nand ginst17433 (P2_U4634, P2_R1179_U112, P2_U3030);
  nand ginst17434 (P2_U4635, P2_U3029, P2_U3395);
  nand ginst17435 (P2_U4636, P2_REG3_REG_2__SCAN_IN, P2_U3028);
  nand ginst17436 (P2_U4637, P2_U3034, P2_U3059);
  nand ginst17437 (P2_U4638, P2_R1179_U22, P2_U3030);
  nand ginst17438 (P2_U4639, P2_U3029, P2_U3398);
  nand ginst17439 (P2_U4640, P2_SUB_605_U26, P2_U3028);
  nand ginst17440 (P2_U4641, P2_U3034, P2_U3066);
  nand ginst17441 (P2_U4642, P2_R1179_U111, P2_U3030);
  nand ginst17442 (P2_U4643, P2_U3029, P2_U3401);
  nand ginst17443 (P2_U4644, P2_SUB_605_U30, P2_U3028);
  nand ginst17444 (P2_U4645, P2_U3034, P2_U3070);
  nand ginst17445 (P2_U4646, P2_R1179_U110, P2_U3030);
  nand ginst17446 (P2_U4647, P2_U3029, P2_U3404);
  nand ginst17447 (P2_U4648, P2_SUB_605_U22, P2_U3028);
  nand ginst17448 (P2_U4649, P2_U3034, P2_U3069);
  nand ginst17449 (P2_U4650, P2_R1179_U23, P2_U3030);
  nand ginst17450 (P2_U4651, P2_U3029, P2_U3407);
  nand ginst17451 (P2_U4652, P2_SUB_605_U8, P2_U3028);
  nand ginst17452 (P2_U4653, P2_U3034, P2_U3083);
  nand ginst17453 (P2_U4654, P2_R1179_U109, P2_U3030);
  nand ginst17454 (P2_U4655, P2_U3029, P2_U3410);
  nand ginst17455 (P2_U4656, P2_SUB_605_U18, P2_U3028);
  nand ginst17456 (P2_U4657, P2_U3034, P2_U3082);
  nand ginst17457 (P2_U4658, P2_R1179_U24, P2_U3030);
  nand ginst17458 (P2_U4659, P2_U3029, P2_U3413);
  nand ginst17459 (P2_U4660, P2_SUB_605_U12, P2_U3028);
  nand ginst17460 (P2_U4661, P2_U3034, P2_U3061);
  nand ginst17461 (P2_U4662, P2_R1179_U108, P2_U3030);
  nand ginst17462 (P2_U4663, P2_U3029, P2_U3416);
  nand ginst17463 (P2_U4664, P2_SUB_605_U14, P2_U3028);
  nand ginst17464 (P2_U4665, P2_U3034, P2_U3062);
  nand ginst17465 (P2_U4666, P2_R1179_U118, P2_U3030);
  nand ginst17466 (P2_U4667, P2_U3029, P2_U3419);
  nand ginst17467 (P2_U4668, P2_SUB_605_U13, P2_U3028);
  nand ginst17468 (P2_U4669, P2_U3034, P2_U3071);
  nand ginst17469 (P2_U4670, P2_R1179_U17, P2_U3030);
  nand ginst17470 (P2_U4671, P2_U3029, P2_U3422);
  nand ginst17471 (P2_U4672, P2_SUB_605_U9, P2_U3028);
  nand ginst17472 (P2_U4673, P2_U3034, P2_U3079);
  nand ginst17473 (P2_U4674, P2_R1179_U107, P2_U3030);
  nand ginst17474 (P2_U4675, P2_U3029, P2_U3425);
  nand ginst17475 (P2_U4676, P2_SUB_605_U24, P2_U3028);
  nand ginst17476 (P2_U4677, P2_U3034, P2_U3078);
  nand ginst17477 (P2_U4678, P2_R1179_U106, P2_U3030);
  nand ginst17478 (P2_U4679, P2_U3029, P2_U3428);
  nand ginst17479 (P2_U4680, P2_SUB_605_U25, P2_U3028);
  nand ginst17480 (P2_U4681, P2_U3034, P2_U3073);
  nand ginst17481 (P2_U4682, P2_R1179_U117, P2_U3030);
  nand ginst17482 (P2_U4683, P2_U3029, P2_U3431);
  nand ginst17483 (P2_U4684, P2_SUB_605_U31, P2_U3028);
  nand ginst17484 (P2_U4685, P2_U3034, P2_U3072);
  nand ginst17485 (P2_U4686, P2_R1179_U116, P2_U3030);
  nand ginst17486 (P2_U4687, P2_U3029, P2_U3434);
  nand ginst17487 (P2_U4688, P2_SUB_605_U21, P2_U3028);
  nand ginst17488 (P2_U4689, P2_U3034, P2_U3068);
  nand ginst17489 (P2_U4690, P2_R1179_U18, P2_U3030);
  nand ginst17490 (P2_U4691, P2_U3029, P2_U3437);
  nand ginst17491 (P2_U4692, P2_SUB_605_U7, P2_U3028);
  nand ginst17492 (P2_U4693, P2_U3034, P2_U3081);
  nand ginst17493 (P2_U4694, P2_R1179_U105, P2_U3030);
  nand ginst17494 (P2_U4695, P2_U3029, P2_U3440);
  nand ginst17495 (P2_U4696, P2_SUB_605_U19, P2_U3028);
  nand ginst17496 (P2_U4697, P2_U3034, P2_U3080);
  nand ginst17497 (P2_U4698, P2_R1179_U104, P2_U3030);
  nand ginst17498 (P2_U4699, P2_U3029, P2_U3443);
  nand ginst17499 (P2_U4700, P2_SUB_605_U11, P2_U3028);
  nand ginst17500 (P2_U4701, P2_U3034, P2_U3075);
  nand ginst17501 (P2_U4702, P2_R1179_U103, P2_U3030);
  nand ginst17502 (P2_U4703, P2_U3029, P2_U3445);
  nand ginst17503 (P2_U4704, P2_SUB_605_U15, P2_U3028);
  nand ginst17504 (P2_U4705, P2_U3034, P2_U3074);
  nand ginst17505 (P2_U4706, P2_R1179_U101, P2_U3030);
  nand ginst17506 (P2_U4707, P2_U3029, P2_U3903);
  nand ginst17507 (P2_U4708, P2_SUB_605_U20, P2_U3028);
  nand ginst17508 (P2_U4709, P2_U3034, P2_U3060);
  nand ginst17509 (P2_U4710, P2_R1179_U115, P2_U3030);
  nand ginst17510 (P2_U4711, P2_U3029, P2_U3902);
  nand ginst17511 (P2_U4712, P2_SUB_605_U28, P2_U3028);
  nand ginst17512 (P2_U4713, P2_U3034, P2_U3065);
  nand ginst17513 (P2_U4714, P2_R1179_U114, P2_U3030);
  nand ginst17514 (P2_U4715, P2_U3029, P2_U3901);
  nand ginst17515 (P2_U4716, P2_SUB_605_U17, P2_U3028);
  nand ginst17516 (P2_U4717, P2_U3034, P2_U3064);
  nand ginst17517 (P2_U4718, P2_R1179_U19, P2_U3030);
  nand ginst17518 (P2_U4719, P2_U3029, P2_U3900);
  nand ginst17519 (P2_U4720, P2_SUB_605_U6, P2_U3028);
  nand ginst17520 (P2_U4721, P2_U3034, P2_U3057);
  nand ginst17521 (P2_U4722, P2_R1179_U100, P2_U3030);
  nand ginst17522 (P2_U4723, P2_U3029, P2_U3899);
  nand ginst17523 (P2_U4724, P2_SUB_605_U10, P2_U3028);
  nand ginst17524 (P2_U4725, P2_U3034, P2_U3056);
  nand ginst17525 (P2_U4726, P2_R1179_U99, P2_U3030);
  nand ginst17526 (P2_U4727, P2_U3029, P2_U3898);
  nand ginst17527 (P2_U4728, P2_SUB_605_U16, P2_U3028);
  nand ginst17528 (P2_U4729, P2_U3034, P2_U3052);
  nand ginst17529 (P2_U4730, P2_R1179_U113, P2_U3030);
  nand ginst17530 (P2_U4731, P2_U3029, P2_U3897);
  nand ginst17531 (P2_U4732, P2_SUB_605_U27, P2_U3028);
  nand ginst17532 (P2_U4733, P2_U3034, P2_U3053);
  nand ginst17533 (P2_U4734, P2_R1179_U20, P2_U3030);
  nand ginst17534 (P2_U4735, P2_U3029, P2_U3896);
  nand ginst17535 (P2_U4736, P2_SUB_605_U23, P2_U3028);
  nand ginst17536 (P2_U4737, P2_U3034, P2_U3054);
  nand ginst17537 (P2_U4738, P2_R1179_U98, P2_U3030);
  nand ginst17538 (P2_U4739, P2_U3029, P2_U3895);
  nand ginst17539 (P2_U4740, P2_SUB_605_U29, P2_U3028);
  nand ginst17540 (P2_U4741, P2_R1179_U21, P2_U3030);
  nand ginst17541 (P2_U4742, P2_U3029, P2_U3904);
  nand ginst17542 (P2_U4743, P2_SUB_605_U94, P2_U3028);
  nand ginst17543 (P2_U4744, P2_SUB_605_U94, P2_U3028);
  nand ginst17544 (P2_U4745, P2_U3908, P2_U3912);
  nand ginst17545 (P2_U4746, P2_U3029, P2_U3869);
  nand ginst17546 (P2_U4747, P2_REG2_REG_30__SCAN_IN, P2_U3358);
  nand ginst17547 (P2_U4748, P2_U3029, P2_U3868);
  nand ginst17548 (P2_U4749, P2_REG2_REG_31__SCAN_IN, P2_U3358);
  nand ginst17549 (P2_U4750, P2_U3359, P2_U3702, P2_U3703, P2_U4624);
  nand ginst17550 (P2_U4751, P2_R1212_U6, P2_U3040);
  nand ginst17551 (P2_U4752, P2_U3039, P2_U3379);
  nand ginst17552 (P2_U4753, P2_R1209_U6, P2_U3037);
  nand ginst17553 (P2_U4754, P2_U4751, P2_U4752, P2_U4753);
  nand ginst17554 (P2_U4755, P2_U3906, P2_U5436);
  not ginst17555 (P2_U4756, P2_U3366);
  nand ginst17556 (P2_U4757, P2_U3829, P2_U3892);
  nand ginst17557 (P2_U4758, P2_R1054_U67, P2_U3051);
  nand ginst17558 (P2_U4759, P2_U3379, P2_U5764);
  nand ginst17559 (P2_U4760, P2_U3042, P2_U4754);
  nand ginst17560 (P2_U4761, P2_R1212_U6, P2_U3041);
  nand ginst17561 (P2_U4762, P2_REG3_REG_19__SCAN_IN, P2_U3151);
  nand ginst17562 (P2_U4763, P2_R1209_U6, P2_U3038);
  nand ginst17563 (P2_U4764, P2_ADDR_REG_19__SCAN_IN, P2_U4756);
  nand ginst17564 (P2_U4765, P2_R1212_U58, P2_U3040);
  nand ginst17565 (P2_U4766, P2_U3039, P2_U3442);
  nand ginst17566 (P2_U4767, P2_R1209_U58, P2_U3037);
  nand ginst17567 (P2_U4768, P2_U4765, P2_U4766, P2_U4767);
  nand ginst17568 (P2_U4769, P2_R1054_U68, P2_U3051);
  nand ginst17569 (P2_U4770, P2_U3442, P2_U5764);
  nand ginst17570 (P2_U4771, P2_U3042, P2_U4768);
  nand ginst17571 (P2_U4772, P2_R1212_U58, P2_U3041);
  nand ginst17572 (P2_U4773, P2_REG3_REG_18__SCAN_IN, P2_U3151);
  nand ginst17573 (P2_U4774, P2_R1209_U58, P2_U3038);
  nand ginst17574 (P2_U4775, P2_ADDR_REG_18__SCAN_IN, P2_U4756);
  nand ginst17575 (P2_U4776, P2_R1212_U59, P2_U3040);
  nand ginst17576 (P2_U4777, P2_U3039, P2_U3439);
  nand ginst17577 (P2_U4778, P2_R1209_U59, P2_U3037);
  nand ginst17578 (P2_U4779, P2_U4776, P2_U4777, P2_U4778);
  nand ginst17579 (P2_U4780, P2_R1054_U69, P2_U3051);
  nand ginst17580 (P2_U4781, P2_U3439, P2_U5764);
  nand ginst17581 (P2_U4782, P2_U3042, P2_U4779);
  nand ginst17582 (P2_U4783, P2_R1212_U59, P2_U3041);
  nand ginst17583 (P2_U4784, P2_REG3_REG_17__SCAN_IN, P2_U3151);
  nand ginst17584 (P2_U4785, P2_R1209_U59, P2_U3038);
  nand ginst17585 (P2_U4786, P2_ADDR_REG_17__SCAN_IN, P2_U4756);
  nand ginst17586 (P2_U4787, P2_R1212_U60, P2_U3040);
  nand ginst17587 (P2_U4788, P2_U3039, P2_U3436);
  nand ginst17588 (P2_U4789, P2_R1209_U60, P2_U3037);
  nand ginst17589 (P2_U4790, P2_U4787, P2_U4788, P2_U4789);
  nand ginst17590 (P2_U4791, P2_R1054_U13, P2_U3051);
  nand ginst17591 (P2_U4792, P2_U3436, P2_U5764);
  nand ginst17592 (P2_U4793, P2_U3042, P2_U4790);
  nand ginst17593 (P2_U4794, P2_R1212_U60, P2_U3041);
  nand ginst17594 (P2_U4795, P2_REG3_REG_16__SCAN_IN, P2_U3151);
  nand ginst17595 (P2_U4796, P2_R1209_U60, P2_U3038);
  nand ginst17596 (P2_U4797, P2_ADDR_REG_16__SCAN_IN, P2_U4756);
  nand ginst17597 (P2_U4798, P2_R1212_U61, P2_U3040);
  nand ginst17598 (P2_U4799, P2_U3039, P2_U3433);
  nand ginst17599 (P2_U4800, P2_R1209_U61, P2_U3037);
  nand ginst17600 (P2_U4801, P2_U4798, P2_U4799, P2_U4800);
  nand ginst17601 (P2_U4802, P2_R1054_U77, P2_U3051);
  nand ginst17602 (P2_U4803, P2_U3433, P2_U5764);
  nand ginst17603 (P2_U4804, P2_U3042, P2_U4801);
  nand ginst17604 (P2_U4805, P2_R1212_U61, P2_U3041);
  nand ginst17605 (P2_U4806, P2_REG3_REG_15__SCAN_IN, P2_U3151);
  nand ginst17606 (P2_U4807, P2_R1209_U61, P2_U3038);
  nand ginst17607 (P2_U4808, P2_ADDR_REG_15__SCAN_IN, P2_U4756);
  nand ginst17608 (P2_U4809, P2_R1212_U62, P2_U3040);
  nand ginst17609 (P2_U4810, P2_U3039, P2_U3430);
  nand ginst17610 (P2_U4811, P2_R1209_U62, P2_U3037);
  nand ginst17611 (P2_U4812, P2_U4809, P2_U4810, P2_U4811);
  nand ginst17612 (P2_U4813, P2_R1054_U78, P2_U3051);
  nand ginst17613 (P2_U4814, P2_U3430, P2_U5764);
  nand ginst17614 (P2_U4815, P2_U3042, P2_U4812);
  nand ginst17615 (P2_U4816, P2_R1212_U62, P2_U3041);
  nand ginst17616 (P2_U4817, P2_REG3_REG_14__SCAN_IN, P2_U3151);
  nand ginst17617 (P2_U4818, P2_R1209_U62, P2_U3038);
  nand ginst17618 (P2_U4819, P2_ADDR_REG_14__SCAN_IN, P2_U4756);
  nand ginst17619 (P2_U4820, P2_R1212_U63, P2_U3040);
  nand ginst17620 (P2_U4821, P2_U3039, P2_U3427);
  nand ginst17621 (P2_U4822, P2_R1209_U63, P2_U3037);
  nand ginst17622 (P2_U4823, P2_U4820, P2_U4821, P2_U4822);
  nand ginst17623 (P2_U4824, P2_R1054_U70, P2_U3051);
  nand ginst17624 (P2_U4825, P2_U3427, P2_U5764);
  nand ginst17625 (P2_U4826, P2_U3042, P2_U4823);
  nand ginst17626 (P2_U4827, P2_R1212_U63, P2_U3041);
  nand ginst17627 (P2_U4828, P2_REG3_REG_13__SCAN_IN, P2_U3151);
  nand ginst17628 (P2_U4829, P2_R1209_U63, P2_U3038);
  nand ginst17629 (P2_U4830, P2_ADDR_REG_13__SCAN_IN, P2_U4756);
  nand ginst17630 (P2_U4831, P2_R1212_U64, P2_U3040);
  nand ginst17631 (P2_U4832, P2_U3039, P2_U3424);
  nand ginst17632 (P2_U4833, P2_R1209_U64, P2_U3037);
  nand ginst17633 (P2_U4834, P2_U4831, P2_U4832, P2_U4833);
  nand ginst17634 (P2_U4835, P2_R1054_U71, P2_U3051);
  nand ginst17635 (P2_U4836, P2_U3424, P2_U5764);
  nand ginst17636 (P2_U4837, P2_U3042, P2_U4834);
  nand ginst17637 (P2_U4838, P2_R1212_U64, P2_U3041);
  nand ginst17638 (P2_U4839, P2_REG3_REG_12__SCAN_IN, P2_U3151);
  nand ginst17639 (P2_U4840, P2_R1209_U64, P2_U3038);
  nand ginst17640 (P2_U4841, P2_ADDR_REG_12__SCAN_IN, P2_U4756);
  nand ginst17641 (P2_U4842, P2_R1212_U65, P2_U3040);
  nand ginst17642 (P2_U4843, P2_U3039, P2_U3421);
  nand ginst17643 (P2_U4844, P2_R1209_U65, P2_U3037);
  nand ginst17644 (P2_U4845, P2_U4842, P2_U4843, P2_U4844);
  nand ginst17645 (P2_U4846, P2_R1054_U12, P2_U3051);
  nand ginst17646 (P2_U4847, P2_U3421, P2_U5764);
  nand ginst17647 (P2_U4848, P2_U3042, P2_U4845);
  nand ginst17648 (P2_U4849, P2_R1212_U65, P2_U3041);
  nand ginst17649 (P2_U4850, P2_REG3_REG_11__SCAN_IN, P2_U3151);
  nand ginst17650 (P2_U4851, P2_R1209_U65, P2_U3038);
  nand ginst17651 (P2_U4852, P2_ADDR_REG_11__SCAN_IN, P2_U4756);
  nand ginst17652 (P2_U4853, P2_R1212_U66, P2_U3040);
  nand ginst17653 (P2_U4854, P2_U3039, P2_U3418);
  nand ginst17654 (P2_U4855, P2_R1209_U66, P2_U3037);
  nand ginst17655 (P2_U4856, P2_U4853, P2_U4854, P2_U4855);
  nand ginst17656 (P2_U4857, P2_R1054_U79, P2_U3051);
  nand ginst17657 (P2_U4858, P2_U3418, P2_U5764);
  nand ginst17658 (P2_U4859, P2_U3042, P2_U4856);
  nand ginst17659 (P2_U4860, P2_R1212_U66, P2_U3041);
  nand ginst17660 (P2_U4861, P2_REG3_REG_10__SCAN_IN, P2_U3151);
  nand ginst17661 (P2_U4862, P2_R1209_U66, P2_U3038);
  nand ginst17662 (P2_U4863, P2_ADDR_REG_10__SCAN_IN, P2_U4756);
  nand ginst17663 (P2_U4864, P2_R1212_U49, P2_U3040);
  nand ginst17664 (P2_U4865, P2_U3039, P2_U3415);
  nand ginst17665 (P2_U4866, P2_R1209_U49, P2_U3037);
  nand ginst17666 (P2_U4867, P2_U4864, P2_U4865, P2_U4866);
  nand ginst17667 (P2_U4868, P2_R1054_U72, P2_U3051);
  nand ginst17668 (P2_U4869, P2_U3415, P2_U5764);
  nand ginst17669 (P2_U4870, P2_U3042, P2_U4867);
  nand ginst17670 (P2_U4871, P2_R1212_U49, P2_U3041);
  nand ginst17671 (P2_U4872, P2_REG3_REG_9__SCAN_IN, P2_U3151);
  nand ginst17672 (P2_U4873, P2_R1209_U49, P2_U3038);
  nand ginst17673 (P2_U4874, P2_ADDR_REG_9__SCAN_IN, P2_U4756);
  nand ginst17674 (P2_U4875, P2_R1212_U50, P2_U3040);
  nand ginst17675 (P2_U4876, P2_U3039, P2_U3412);
  nand ginst17676 (P2_U4877, P2_R1209_U50, P2_U3037);
  nand ginst17677 (P2_U4878, P2_U4875, P2_U4876, P2_U4877);
  nand ginst17678 (P2_U4879, P2_R1054_U16, P2_U3051);
  nand ginst17679 (P2_U4880, P2_U3412, P2_U5764);
  nand ginst17680 (P2_U4881, P2_U3042, P2_U4878);
  nand ginst17681 (P2_U4882, P2_R1212_U50, P2_U3041);
  nand ginst17682 (P2_U4883, P2_REG3_REG_8__SCAN_IN, P2_U3151);
  nand ginst17683 (P2_U4884, P2_R1209_U50, P2_U3038);
  nand ginst17684 (P2_U4885, P2_ADDR_REG_8__SCAN_IN, P2_U4756);
  nand ginst17685 (P2_U4886, P2_R1212_U51, P2_U3040);
  nand ginst17686 (P2_U4887, P2_U3039, P2_U3409);
  nand ginst17687 (P2_U4888, P2_R1209_U51, P2_U3037);
  nand ginst17688 (P2_U4889, P2_U4886, P2_U4887, P2_U4888);
  nand ginst17689 (P2_U4890, P2_R1054_U73, P2_U3051);
  nand ginst17690 (P2_U4891, P2_U3409, P2_U5764);
  nand ginst17691 (P2_U4892, P2_U3042, P2_U4889);
  nand ginst17692 (P2_U4893, P2_R1212_U51, P2_U3041);
  nand ginst17693 (P2_U4894, P2_REG3_REG_7__SCAN_IN, P2_U3151);
  nand ginst17694 (P2_U4895, P2_R1209_U51, P2_U3038);
  nand ginst17695 (P2_U4896, P2_ADDR_REG_7__SCAN_IN, P2_U4756);
  nand ginst17696 (P2_U4897, P2_R1212_U52, P2_U3040);
  nand ginst17697 (P2_U4898, P2_U3039, P2_U3406);
  nand ginst17698 (P2_U4899, P2_R1209_U52, P2_U3037);
  nand ginst17699 (P2_U4900, P2_U4897, P2_U4898, P2_U4899);
  nand ginst17700 (P2_U4901, P2_R1054_U15, P2_U3051);
  nand ginst17701 (P2_U4902, P2_U3406, P2_U5764);
  nand ginst17702 (P2_U4903, P2_U3042, P2_U4900);
  nand ginst17703 (P2_U4904, P2_R1212_U52, P2_U3041);
  nand ginst17704 (P2_U4905, P2_REG3_REG_6__SCAN_IN, P2_U3151);
  nand ginst17705 (P2_U4906, P2_R1209_U52, P2_U3038);
  nand ginst17706 (P2_U4907, P2_ADDR_REG_6__SCAN_IN, P2_U4756);
  nand ginst17707 (P2_U4908, P2_R1212_U53, P2_U3040);
  nand ginst17708 (P2_U4909, P2_U3039, P2_U3403);
  nand ginst17709 (P2_U4910, P2_R1209_U53, P2_U3037);
  nand ginst17710 (P2_U4911, P2_U4908, P2_U4909, P2_U4910);
  nand ginst17711 (P2_U4912, P2_R1054_U74, P2_U3051);
  nand ginst17712 (P2_U4913, P2_U3403, P2_U5764);
  nand ginst17713 (P2_U4914, P2_U3042, P2_U4911);
  nand ginst17714 (P2_U4915, P2_R1212_U53, P2_U3041);
  nand ginst17715 (P2_U4916, P2_REG3_REG_5__SCAN_IN, P2_U3151);
  nand ginst17716 (P2_U4917, P2_R1209_U53, P2_U3038);
  nand ginst17717 (P2_U4918, P2_ADDR_REG_5__SCAN_IN, P2_U4756);
  nand ginst17718 (P2_U4919, P2_R1212_U54, P2_U3040);
  nand ginst17719 (P2_U4920, P2_U3039, P2_U3400);
  nand ginst17720 (P2_U4921, P2_R1209_U54, P2_U3037);
  nand ginst17721 (P2_U4922, P2_U4919, P2_U4920, P2_U4921);
  nand ginst17722 (P2_U4923, P2_R1054_U75, P2_U3051);
  nand ginst17723 (P2_U4924, P2_U3400, P2_U5764);
  nand ginst17724 (P2_U4925, P2_U3042, P2_U4922);
  nand ginst17725 (P2_U4926, P2_R1212_U54, P2_U3041);
  nand ginst17726 (P2_U4927, P2_REG3_REG_4__SCAN_IN, P2_U3151);
  nand ginst17727 (P2_U4928, P2_R1209_U54, P2_U3038);
  nand ginst17728 (P2_U4929, P2_ADDR_REG_4__SCAN_IN, P2_U4756);
  nand ginst17729 (P2_U4930, P2_R1212_U55, P2_U3040);
  nand ginst17730 (P2_U4931, P2_U3039, P2_U3397);
  nand ginst17731 (P2_U4932, P2_R1209_U55, P2_U3037);
  nand ginst17732 (P2_U4933, P2_U4930, P2_U4931, P2_U4932);
  nand ginst17733 (P2_U4934, P2_R1054_U14, P2_U3051);
  nand ginst17734 (P2_U4935, P2_U3397, P2_U5764);
  nand ginst17735 (P2_U4936, P2_U3042, P2_U4933);
  nand ginst17736 (P2_U4937, P2_R1212_U55, P2_U3041);
  nand ginst17737 (P2_U4938, P2_REG3_REG_3__SCAN_IN, P2_U3151);
  nand ginst17738 (P2_U4939, P2_R1209_U55, P2_U3038);
  nand ginst17739 (P2_U4940, P2_ADDR_REG_3__SCAN_IN, P2_U4756);
  nand ginst17740 (P2_U4941, P2_R1212_U56, P2_U3040);
  nand ginst17741 (P2_U4942, P2_U3039, P2_U3394);
  nand ginst17742 (P2_U4943, P2_R1209_U56, P2_U3037);
  nand ginst17743 (P2_U4944, P2_U4941, P2_U4942, P2_U4943);
  nand ginst17744 (P2_U4945, P2_R1054_U76, P2_U3051);
  nand ginst17745 (P2_U4946, P2_U3394, P2_U5764);
  nand ginst17746 (P2_U4947, P2_U3042, P2_U4944);
  nand ginst17747 (P2_U4948, P2_R1212_U56, P2_U3041);
  nand ginst17748 (P2_U4949, P2_REG3_REG_2__SCAN_IN, P2_U3151);
  nand ginst17749 (P2_U4950, P2_R1209_U56, P2_U3038);
  nand ginst17750 (P2_U4951, P2_ADDR_REG_2__SCAN_IN, P2_U4756);
  nand ginst17751 (P2_U4952, P2_R1212_U57, P2_U3040);
  nand ginst17752 (P2_U4953, P2_U3039, P2_U3391);
  nand ginst17753 (P2_U4954, P2_R1209_U57, P2_U3037);
  nand ginst17754 (P2_U4955, P2_U4952, P2_U4953, P2_U4954);
  nand ginst17755 (P2_U4956, P2_R1054_U66, P2_U3051);
  nand ginst17756 (P2_U4957, P2_U3391, P2_U5764);
  nand ginst17757 (P2_U4958, P2_U3042, P2_U4955);
  nand ginst17758 (P2_U4959, P2_R1212_U57, P2_U3041);
  nand ginst17759 (P2_U4960, P2_REG3_REG_1__SCAN_IN, P2_U3151);
  nand ginst17760 (P2_U4961, P2_R1209_U57, P2_U3038);
  nand ginst17761 (P2_U4962, P2_ADDR_REG_1__SCAN_IN, P2_U4756);
  nand ginst17762 (P2_U4963, P2_R1212_U7, P2_U3040);
  nand ginst17763 (P2_U4964, P2_U3039, P2_U3386);
  nand ginst17764 (P2_U4965, P2_R1209_U7, P2_U3037);
  nand ginst17765 (P2_U4966, P2_U4963, P2_U4964, P2_U4965);
  nand ginst17766 (P2_U4967, P2_R1054_U17, P2_U3051);
  nand ginst17767 (P2_U4968, P2_U3386, P2_U5764);
  nand ginst17768 (P2_U4969, P2_U3042, P2_U4966);
  nand ginst17769 (P2_U4970, P2_R1212_U7, P2_U3041);
  nand ginst17770 (P2_U4971, P2_REG3_REG_0__SCAN_IN, P2_U3151);
  nand ginst17771 (P2_U4972, P2_R1209_U7, P2_U3038);
  nand ginst17772 (P2_U4973, P2_ADDR_REG_0__SCAN_IN, P2_U4756);
  not ginst17773 (P2_U4974, P2_U3864);
  nand ginst17774 (P2_U4975, P2_U3050, P2_U5937, P2_U5938);
  nand ginst17775 (P2_U4976, P2_U3023, P2_U3863, P2_U3905);
  nand ginst17776 (P2_U4977, P2_B_REG_SCAN_IN, P2_U4975);
  nand ginst17777 (P2_U4978, P2_U3036, P2_U3078);
  nand ginst17778 (P2_U4979, P2_U3032, P2_U3072);
  nand ginst17779 (P2_U4980, P2_SUB_605_U21, P2_U3304);
  nand ginst17780 (P2_U4981, P2_U4978, P2_U4979, P2_U4980);
  nand ginst17781 (P2_U4982, P2_U3311, P2_U3312, P2_U3871, P2_U3884, P2_U5421);
  nand ginst17782 (P2_U4983, P2_U3890, P2_U4982);
  nand ginst17783 (P2_U4984, P2_U3885, P2_U3891);
  nand ginst17784 (P2_U4985, P2_U4983, P2_U4984);
  nand ginst17785 (P2_U4986, P2_U3378, P2_U3907);
  nand ginst17786 (P2_U4987, P2_U3304, P2_U3885);
  nand ginst17787 (P2_U4988, P2_U3303, P2_U4982);
  not ginst17788 (P2_U4989, P2_U3370);
  nand ginst17789 (P2_U4990, P2_U3434, P2_U5416);
  nand ginst17790 (P2_U4991, P2_SUB_605_U21, P2_U3371);
  nand ginst17791 (P2_U4992, P2_R1158_U114, P2_U3035);
  nand ginst17792 (P2_U4993, P2_U3031, P2_U4981);
  nand ginst17793 (P2_U4994, P2_REG3_REG_15__SCAN_IN, P2_U3151);
  nand ginst17794 (P2_U4995, P2_U3036, P2_U3057);
  nand ginst17795 (P2_U4996, P2_U3032, P2_U3052);
  nand ginst17796 (P2_U4997, P2_SUB_605_U27, P2_U3304);
  nand ginst17797 (P2_U4998, P2_U4995, P2_U4996, P2_U4997);
  nand ginst17798 (P2_U4999, P2_U3303, P2_U3365);
  nand ginst17799 (P2_U5000, P2_U4989, P2_U4999);
  nand ginst17800 (P2_U5001, P2_U3365, P2_U3890);
  nand ginst17801 (P2_U5002, P2_U3360, P2_U5001);
  nand ginst17802 (P2_U5003, P2_U3045, P2_U3897);
  nand ginst17803 (P2_U5004, P2_SUB_605_U27, P2_U3044);
  nand ginst17804 (P2_U5005, P2_R1158_U17, P2_U3035);
  nand ginst17805 (P2_U5006, P2_U3031, P2_U4998);
  nand ginst17806 (P2_U5007, P2_REG3_REG_26__SCAN_IN, P2_U3151);
  nand ginst17807 (P2_U5008, P2_U3036, P2_U3066);
  nand ginst17808 (P2_U5009, P2_U3032, P2_U3069);
  nand ginst17809 (P2_U5010, P2_SUB_605_U8, P2_U3304);
  nand ginst17810 (P2_U5011, P2_U5008, P2_U5009, P2_U5010);
  nand ginst17811 (P2_U5012, P2_U3407, P2_U5416);
  nand ginst17812 (P2_U5013, P2_SUB_605_U8, P2_U3371);
  nand ginst17813 (P2_U5014, P2_R1158_U99, P2_U3035);
  nand ginst17814 (P2_U5015, P2_U3031, P2_U5011);
  nand ginst17815 (P2_U5016, P2_REG3_REG_6__SCAN_IN, P2_U3151);
  nand ginst17816 (P2_U5017, P2_U3036, P2_U3068);
  nand ginst17817 (P2_U5018, P2_U3032, P2_U3080);
  nand ginst17818 (P2_U5019, P2_SUB_605_U11, P2_U3304);
  nand ginst17819 (P2_U5020, P2_U5017, P2_U5018, P2_U5019);
  nand ginst17820 (P2_U5021, P2_U3443, P2_U5416);
  nand ginst17821 (P2_U5022, P2_SUB_605_U11, P2_U3371);
  nand ginst17822 (P2_U5023, P2_R1158_U112, P2_U3035);
  nand ginst17823 (P2_U5024, P2_U3031, P2_U5020);
  nand ginst17824 (P2_U5025, P2_REG3_REG_18__SCAN_IN, P2_U3151);
  nand ginst17825 (P2_U5026, P2_U3036, P2_U3077);
  nand ginst17826 (P2_U5027, P2_U3032, P2_U3063);
  nand ginst17827 (P2_U5028, P2_REG3_REG_2__SCAN_IN, P2_U3304);
  nand ginst17828 (P2_U5029, P2_U5026, P2_U5027, P2_U5028);
  nand ginst17829 (P2_U5030, P2_U3395, P2_U5416);
  nand ginst17830 (P2_U5031, P2_REG3_REG_2__SCAN_IN, P2_U3371);
  nand ginst17831 (P2_U5032, P2_R1158_U102, P2_U3035);
  nand ginst17832 (P2_U5033, P2_U3031, P2_U5029);
  nand ginst17833 (P2_U5034, P2_REG3_REG_2__SCAN_IN, P2_U3151);
  nand ginst17834 (P2_U5035, P2_U3036, P2_U3061);
  nand ginst17835 (P2_U5036, P2_U3032, P2_U3071);
  nand ginst17836 (P2_U5037, P2_SUB_605_U9, P2_U3304);
  nand ginst17837 (P2_U5038, P2_U5035, P2_U5036, P2_U5037);
  nand ginst17838 (P2_U5039, P2_U3422, P2_U5416);
  nand ginst17839 (P2_U5040, P2_SUB_605_U9, P2_U3371);
  nand ginst17840 (P2_U5041, P2_R1158_U117, P2_U3035);
  nand ginst17841 (P2_U5042, P2_U3031, P2_U5038);
  nand ginst17842 (P2_U5043, P2_REG3_REG_11__SCAN_IN, P2_U3151);
  nand ginst17843 (P2_U5044, P2_U3036, P2_U3074);
  nand ginst17844 (P2_U5045, P2_U3032, P2_U3065);
  nand ginst17845 (P2_U5046, P2_SUB_605_U17, P2_U3304);
  nand ginst17846 (P2_U5047, P2_U5044, P2_U5045, P2_U5046);
  nand ginst17847 (P2_U5048, P2_U3045, P2_U3901);
  nand ginst17848 (P2_U5049, P2_SUB_605_U17, P2_U3044);
  nand ginst17849 (P2_U5050, P2_R1158_U108, P2_U3035);
  nand ginst17850 (P2_U5051, P2_U3031, P2_U5047);
  nand ginst17851 (P2_U5052, P2_REG3_REG_22__SCAN_IN, P2_U3151);
  nand ginst17852 (P2_U5053, P2_U3036, P2_U3071);
  nand ginst17853 (P2_U5054, P2_U3032, P2_U3078);
  nand ginst17854 (P2_U5055, P2_SUB_605_U25, P2_U3304);
  nand ginst17855 (P2_U5056, P2_U5053, P2_U5054, P2_U5055);
  nand ginst17856 (P2_U5057, P2_U3428, P2_U5416);
  nand ginst17857 (P2_U5058, P2_SUB_605_U25, P2_U3371);
  nand ginst17858 (P2_U5059, P2_R1158_U14, P2_U3035);
  nand ginst17859 (P2_U5060, P2_U3031, P2_U5056);
  nand ginst17860 (P2_U5061, P2_REG3_REG_13__SCAN_IN, P2_U3151);
  nand ginst17861 (P2_U5062, P2_U3036, P2_U3080);
  nand ginst17862 (P2_U5063, P2_U3032, P2_U3074);
  nand ginst17863 (P2_U5064, P2_SUB_605_U20, P2_U3304);
  nand ginst17864 (P2_U5065, P2_U5062, P2_U5063, P2_U5064);
  nand ginst17865 (P2_U5066, P2_U3045, P2_U3903);
  nand ginst17866 (P2_U5067, P2_SUB_605_U20, P2_U3044);
  nand ginst17867 (P2_U5068, P2_R1158_U109, P2_U3035);
  nand ginst17868 (P2_U5069, P2_U3031, P2_U5065);
  nand ginst17869 (P2_U5070, P2_REG3_REG_20__SCAN_IN, P2_U3151);
  nand ginst17870 (P2_U5071, P2_U3031, P2_U3304);
  nand ginst17871 (P2_U5072, P2_U5071, P2_U5415);
  nand ginst17872 (P2_U5073, P2_U3032, P2_U3792);
  nand ginst17873 (P2_U5074, P2_U3387, P2_U5416);
  nand ginst17874 (P2_U5075, P2_REG3_REG_0__SCAN_IN, P2_U5072);
  nand ginst17875 (P2_U5076, P2_R1158_U96, P2_U3035);
  nand ginst17876 (P2_U5077, P2_REG3_REG_0__SCAN_IN, P2_U3151);
  nand ginst17877 (P2_U5078, P2_U3036, P2_U3083);
  nand ginst17878 (P2_U5079, P2_U3032, P2_U3061);
  nand ginst17879 (P2_U5080, P2_SUB_605_U14, P2_U3304);
  nand ginst17880 (P2_U5081, P2_U5078, P2_U5079, P2_U5080);
  nand ginst17881 (P2_U5082, P2_U3416, P2_U5416);
  nand ginst17882 (P2_U5083, P2_SUB_605_U14, P2_U3371);
  nand ginst17883 (P2_U5084, P2_R1158_U97, P2_U3035);
  nand ginst17884 (P2_U5085, P2_U3031, P2_U5081);
  nand ginst17885 (P2_U5086, P2_REG3_REG_9__SCAN_IN, P2_U3151);
  nand ginst17886 (P2_U5087, P2_U3036, P2_U3063);
  nand ginst17887 (P2_U5088, P2_U3032, P2_U3066);
  nand ginst17888 (P2_U5089, P2_SUB_605_U30, P2_U3304);
  nand ginst17889 (P2_U5090, P2_U5087, P2_U5088, P2_U5089);
  nand ginst17890 (P2_U5091, P2_U3401, P2_U5416);
  nand ginst17891 (P2_U5092, P2_SUB_605_U30, P2_U3371);
  nand ginst17892 (P2_U5093, P2_R1158_U101, P2_U3035);
  nand ginst17893 (P2_U5094, P2_U3031, P2_U5090);
  nand ginst17894 (P2_U5095, P2_REG3_REG_4__SCAN_IN, P2_U3151);
  nand ginst17895 (P2_U5096, P2_U3036, P2_U3065);
  nand ginst17896 (P2_U5097, P2_U3032, P2_U3057);
  nand ginst17897 (P2_U5098, P2_SUB_605_U10, P2_U3304);
  nand ginst17898 (P2_U5099, P2_U5096, P2_U5097, P2_U5098);
  nand ginst17899 (P2_U5100, P2_U3045, P2_U3899);
  nand ginst17900 (P2_U5101, P2_SUB_605_U10, P2_U3044);
  nand ginst17901 (P2_U5102, P2_R1158_U106, P2_U3035);
  nand ginst17902 (P2_U5103, P2_U3031, P2_U5099);
  nand ginst17903 (P2_U5104, P2_REG3_REG_24__SCAN_IN, P2_U3151);
  nand ginst17904 (P2_U5105, P2_U3036, P2_U3072);
  nand ginst17905 (P2_U5106, P2_U3032, P2_U3081);
  nand ginst17906 (P2_U5107, P2_SUB_605_U19, P2_U3304);
  nand ginst17907 (P2_U5108, P2_U5105, P2_U5106, P2_U5107);
  nand ginst17908 (P2_U5109, P2_U3440, P2_U5416);
  nand ginst17909 (P2_U5110, P2_SUB_605_U19, P2_U3371);
  nand ginst17910 (P2_U5111, P2_R1158_U15, P2_U3035);
  nand ginst17911 (P2_U5112, P2_U3031, P2_U5108);
  nand ginst17912 (P2_U5113, P2_REG3_REG_17__SCAN_IN, P2_U3151);
  nand ginst17913 (P2_U5114, P2_U3036, P2_U3059);
  nand ginst17914 (P2_U5115, P2_U3032, P2_U3070);
  nand ginst17915 (P2_U5116, P2_SUB_605_U22, P2_U3304);
  nand ginst17916 (P2_U5117, P2_U5114, P2_U5115, P2_U5116);
  nand ginst17917 (P2_U5118, P2_U3404, P2_U5416);
  nand ginst17918 (P2_U5119, P2_SUB_605_U22, P2_U3371);
  nand ginst17919 (P2_U5120, P2_R1158_U100, P2_U3035);
  nand ginst17920 (P2_U5121, P2_U3031, P2_U5117);
  nand ginst17921 (P2_U5122, P2_REG3_REG_5__SCAN_IN, P2_U3151);
  nand ginst17922 (P2_U5123, P2_U3036, P2_U3073);
  nand ginst17923 (P2_U5124, P2_U3032, P2_U3068);
  nand ginst17924 (P2_U5125, P2_SUB_605_U7, P2_U3304);
  nand ginst17925 (P2_U5126, P2_U5123, P2_U5124, P2_U5125);
  nand ginst17926 (P2_U5127, P2_U3437, P2_U5416);
  nand ginst17927 (P2_U5128, P2_SUB_605_U7, P2_U3371);
  nand ginst17928 (P2_U5129, P2_R1158_U113, P2_U3035);
  nand ginst17929 (P2_U5130, P2_U3031, P2_U5126);
  nand ginst17930 (P2_U5131, P2_REG3_REG_16__SCAN_IN, P2_U3151);
  nand ginst17931 (P2_U5132, P2_U3036, P2_U3064);
  nand ginst17932 (P2_U5133, P2_U3032, P2_U3056);
  nand ginst17933 (P2_U5134, P2_SUB_605_U16, P2_U3304);
  nand ginst17934 (P2_U5135, P2_U5132, P2_U5133, P2_U5134);
  nand ginst17935 (P2_U5136, P2_U3045, P2_U3898);
  nand ginst17936 (P2_U5137, P2_SUB_605_U16, P2_U3044);
  nand ginst17937 (P2_U5138, P2_R1158_U105, P2_U3035);
  nand ginst17938 (P2_U5139, P2_U3031, P2_U5135);
  nand ginst17939 (P2_U5140, P2_REG3_REG_25__SCAN_IN, P2_U3151);
  nand ginst17940 (P2_U5141, P2_U3036, P2_U3062);
  nand ginst17941 (P2_U5142, P2_U3032, P2_U3079);
  nand ginst17942 (P2_U5143, P2_SUB_605_U24, P2_U3304);
  nand ginst17943 (P2_U5144, P2_U5141, P2_U5142, P2_U5143);
  nand ginst17944 (P2_U5145, P2_U3425, P2_U5416);
  nand ginst17945 (P2_U5146, P2_SUB_605_U24, P2_U3371);
  nand ginst17946 (P2_U5147, P2_R1158_U116, P2_U3035);
  nand ginst17947 (P2_U5148, P2_U3031, P2_U5144);
  nand ginst17948 (P2_U5149, P2_REG3_REG_12__SCAN_IN, P2_U3151);
  nand ginst17949 (P2_U5150, P2_U3036, P2_U3075);
  nand ginst17950 (P2_U5151, P2_U3032, P2_U3060);
  nand ginst17951 (P2_U5152, P2_SUB_605_U28, P2_U3304);
  nand ginst17952 (P2_U5153, P2_U5150, P2_U5151, P2_U5152);
  nand ginst17953 (P2_U5154, P2_U3045, P2_U3902);
  nand ginst17954 (P2_U5155, P2_SUB_605_U28, P2_U3044);
  nand ginst17955 (P2_U5156, P2_R1158_U16, P2_U3035);
  nand ginst17956 (P2_U5157, P2_U3031, P2_U5153);
  nand ginst17957 (P2_U5158, P2_REG3_REG_21__SCAN_IN, P2_U3151);
  nand ginst17958 (P2_U5159, P2_U3036, P2_U3076);
  nand ginst17959 (P2_U5160, P2_U3032, P2_U3067);
  nand ginst17960 (P2_U5161, P2_REG3_REG_1__SCAN_IN, P2_U3304);
  nand ginst17961 (P2_U5162, P2_U5159, P2_U5160, P2_U5161);
  nand ginst17962 (P2_U5163, P2_U3392, P2_U5416);
  nand ginst17963 (P2_U5164, P2_REG3_REG_1__SCAN_IN, P2_U3371);
  nand ginst17964 (P2_U5165, P2_R1158_U110, P2_U3035);
  nand ginst17965 (P2_U5166, P2_U3031, P2_U5162);
  nand ginst17966 (P2_U5167, P2_REG3_REG_1__SCAN_IN, P2_U3151);
  nand ginst17967 (P2_U5168, P2_U3036, P2_U3069);
  nand ginst17968 (P2_U5169, P2_U3032, P2_U3082);
  nand ginst17969 (P2_U5170, P2_SUB_605_U12, P2_U3304);
  nand ginst17970 (P2_U5171, P2_U5168, P2_U5169, P2_U5170);
  nand ginst17971 (P2_U5172, P2_U3413, P2_U5416);
  nand ginst17972 (P2_U5173, P2_SUB_605_U12, P2_U3371);
  nand ginst17973 (P2_U5174, P2_R1158_U98, P2_U3035);
  nand ginst17974 (P2_U5175, P2_U3031, P2_U5171);
  nand ginst17975 (P2_U5176, P2_REG3_REG_8__SCAN_IN, P2_U3151);
  nand ginst17976 (P2_U5177, P2_U3036, P2_U3052);
  nand ginst17977 (P2_U5178, P2_U3032, P2_U3054);
  nand ginst17978 (P2_U5179, P2_SUB_605_U29, P2_U3304);
  nand ginst17979 (P2_U5180, P2_U5177, P2_U5178, P2_U5179);
  nand ginst17980 (P2_U5181, P2_U3045, P2_U3895);
  nand ginst17981 (P2_U5182, P2_SUB_605_U29, P2_U3044);
  nand ginst17982 (P2_U5183, P2_R1158_U103, P2_U3035);
  nand ginst17983 (P2_U5184, P2_U3031, P2_U5180);
  nand ginst17984 (P2_U5185, P2_REG3_REG_28__SCAN_IN, P2_U3151);
  nand ginst17985 (P2_U5186, P2_U3036, P2_U3081);
  nand ginst17986 (P2_U5187, P2_U3032, P2_U3075);
  nand ginst17987 (P2_U5188, P2_SUB_605_U15, P2_U3304);
  nand ginst17988 (P2_U5189, P2_U5186, P2_U5187, P2_U5188);
  nand ginst17989 (P2_U5190, P2_U3445, P2_U5416);
  nand ginst17990 (P2_U5191, P2_SUB_605_U15, P2_U3371);
  nand ginst17991 (P2_U5192, P2_R1158_U111, P2_U3035);
  nand ginst17992 (P2_U5193, P2_U3031, P2_U5189);
  nand ginst17993 (P2_U5194, P2_REG3_REG_19__SCAN_IN, P2_U3151);
  nand ginst17994 (P2_U5195, P2_U3036, P2_U3067);
  nand ginst17995 (P2_U5196, P2_U3032, P2_U3059);
  nand ginst17996 (P2_U5197, P2_SUB_605_U26, P2_U3304);
  nand ginst17997 (P2_U5198, P2_U5195, P2_U5196, P2_U5197);
  nand ginst17998 (P2_U5199, P2_U3398, P2_U5416);
  nand ginst17999 (P2_U5200, P2_SUB_605_U26, P2_U3371);
  nand ginst18000 (P2_U5201, P2_R1158_U18, P2_U3035);
  nand ginst18001 (P2_U5202, P2_U3031, P2_U5198);
  nand ginst18002 (P2_U5203, P2_REG3_REG_3__SCAN_IN, P2_U3151);
  nand ginst18003 (P2_U5204, P2_U3036, P2_U3082);
  nand ginst18004 (P2_U5205, P2_U3032, P2_U3062);
  nand ginst18005 (P2_U5206, P2_SUB_605_U13, P2_U3304);
  nand ginst18006 (P2_U5207, P2_U5204, P2_U5205, P2_U5206);
  nand ginst18007 (P2_U5208, P2_U3419, P2_U5416);
  nand ginst18008 (P2_U5209, P2_SUB_605_U13, P2_U3371);
  nand ginst18009 (P2_U5210, P2_R1158_U118, P2_U3035);
  nand ginst18010 (P2_U5211, P2_U3031, P2_U5207);
  nand ginst18011 (P2_U5212, P2_REG3_REG_10__SCAN_IN, P2_U3151);
  nand ginst18012 (P2_U5213, P2_U3036, P2_U3060);
  nand ginst18013 (P2_U5214, P2_U3032, P2_U3064);
  nand ginst18014 (P2_U5215, P2_SUB_605_U6, P2_U3304);
  nand ginst18015 (P2_U5216, P2_U5213, P2_U5214, P2_U5215);
  nand ginst18016 (P2_U5217, P2_U3045, P2_U3900);
  nand ginst18017 (P2_U5218, P2_SUB_605_U6, P2_U3044);
  nand ginst18018 (P2_U5219, P2_R1158_U107, P2_U3035);
  nand ginst18019 (P2_U5220, P2_U3031, P2_U5216);
  nand ginst18020 (P2_U5221, P2_REG3_REG_23__SCAN_IN, P2_U3151);
  nand ginst18021 (P2_U5222, P2_U3036, P2_U3079);
  nand ginst18022 (P2_U5223, P2_U3032, P2_U3073);
  nand ginst18023 (P2_U5224, P2_SUB_605_U31, P2_U3304);
  nand ginst18024 (P2_U5225, P2_U5222, P2_U5223, P2_U5224);
  nand ginst18025 (P2_U5226, P2_U3431, P2_U5416);
  nand ginst18026 (P2_U5227, P2_SUB_605_U31, P2_U3371);
  nand ginst18027 (P2_U5228, P2_R1158_U115, P2_U3035);
  nand ginst18028 (P2_U5229, P2_U3031, P2_U5225);
  nand ginst18029 (P2_U5230, P2_REG3_REG_14__SCAN_IN, P2_U3151);
  nand ginst18030 (P2_U5231, P2_U3036, P2_U3056);
  nand ginst18031 (P2_U5232, P2_U3032, P2_U3053);
  nand ginst18032 (P2_U5233, P2_SUB_605_U23, P2_U3304);
  nand ginst18033 (P2_U5234, P2_U5231, P2_U5232, P2_U5233);
  nand ginst18034 (P2_U5235, P2_U3045, P2_U3896);
  nand ginst18035 (P2_U5236, P2_SUB_605_U23, P2_U3044);
  nand ginst18036 (P2_U5237, P2_R1158_U104, P2_U3035);
  nand ginst18037 (P2_U5238, P2_U3031, P2_U5234);
  nand ginst18038 (P2_U5239, P2_REG3_REG_27__SCAN_IN, P2_U3151);
  nand ginst18039 (P2_U5240, P2_U3036, P2_U3070);
  nand ginst18040 (P2_U5241, P2_U3032, P2_U3083);
  nand ginst18041 (P2_U5242, P2_SUB_605_U18, P2_U3304);
  nand ginst18042 (P2_U5243, P2_U5240, P2_U5241, P2_U5242);
  nand ginst18043 (P2_U5244, P2_U3410, P2_U5416);
  nand ginst18044 (P2_U5245, P2_SUB_605_U18, P2_U3371);
  nand ginst18045 (P2_U5246, P2_R1158_U19, P2_U3035);
  nand ginst18046 (P2_U5247, P2_U3031, P2_U5243);
  nand ginst18047 (P2_U5248, P2_REG3_REG_7__SCAN_IN, P2_U3151);
  nand ginst18048 (P2_U5249, P2_U3046, P2_U3894);
  nand ginst18049 (P2_U5250, P2_U3375, P2_U3829);
  nand ginst18050 (P2_U5251, P2_U3820, P2_U3821);
  nand ginst18051 (P2_U5252, P2_U3013, P2_U3819);
  nand ginst18052 (P2_U5253, P2_U3876, P2_U5252);
  nand ginst18053 (P2_U5254, P2_U3416, P2_U5253);
  nand ginst18054 (P2_U5255, P2_U3082, P2_U5251);
  nand ginst18055 (P2_U5256, P2_U3413, P2_U5253);
  nand ginst18056 (P2_U5257, P2_U3083, P2_U5251);
  nand ginst18057 (P2_U5258, P2_U3410, P2_U5253);
  nand ginst18058 (P2_U5259, P2_U3069, P2_U5251);
  nand ginst18059 (P2_U5260, P2_U3407, P2_U5253);
  nand ginst18060 (P2_U5261, P2_U3070, P2_U5251);
  nand ginst18061 (P2_U5262, P2_U3404, P2_U5253);
  nand ginst18062 (P2_U5263, P2_U3066, P2_U5251);
  nand ginst18063 (P2_U5264, P2_U3401, P2_U5253);
  nand ginst18064 (P2_U5265, P2_U3059, P2_U5251);
  nand ginst18065 (P2_U5266, P2_U3868, P2_U5253);
  nand ginst18066 (P2_U5267, P2_U3055, P2_U5251);
  nand ginst18067 (P2_U5268, P2_U3869, P2_U5253);
  nand ginst18068 (P2_U5269, P2_U3058, P2_U5251);
  nand ginst18069 (P2_U5270, P2_U3398, P2_U5253);
  nand ginst18070 (P2_U5271, P2_U3063, P2_U5251);
  nand ginst18071 (P2_U5272, P2_U3904, P2_U5253);
  nand ginst18072 (P2_U5273, P2_U3054, P2_U5251);
  nand ginst18073 (P2_U5274, P2_U3895, P2_U5253);
  nand ginst18074 (P2_U5275, P2_U3053, P2_U5251);
  nand ginst18075 (P2_U5276, P2_U3896, P2_U5253);
  nand ginst18076 (P2_U5277, P2_U3052, P2_U5251);
  nand ginst18077 (P2_U5278, P2_U3897, P2_U5253);
  nand ginst18078 (P2_U5279, P2_U3056, P2_U5251);
  nand ginst18079 (P2_U5280, P2_U3898, P2_U5253);
  nand ginst18080 (P2_U5281, P2_U3057, P2_U5251);
  nand ginst18081 (P2_U5282, P2_U3899, P2_U5253);
  nand ginst18082 (P2_U5283, P2_U3064, P2_U5251);
  nand ginst18083 (P2_U5284, P2_U3900, P2_U5253);
  nand ginst18084 (P2_U5285, P2_U3065, P2_U5251);
  nand ginst18085 (P2_U5286, P2_U3901, P2_U5253);
  nand ginst18086 (P2_U5287, P2_U3060, P2_U5251);
  nand ginst18087 (P2_U5288, P2_U3902, P2_U5253);
  nand ginst18088 (P2_U5289, P2_U3074, P2_U5251);
  nand ginst18089 (P2_U5290, P2_U3903, P2_U5253);
  nand ginst18090 (P2_U5291, P2_U3075, P2_U5251);
  nand ginst18091 (P2_U5292, P2_U3395, P2_U5253);
  nand ginst18092 (P2_U5293, P2_U3067, P2_U5251);
  nand ginst18093 (P2_U5294, P2_U3445, P2_U5253);
  nand ginst18094 (P2_U5295, P2_U3080, P2_U5251);
  nand ginst18095 (P2_U5296, P2_U3443, P2_U5253);
  nand ginst18096 (P2_U5297, P2_U3081, P2_U5251);
  nand ginst18097 (P2_U5298, P2_U3440, P2_U5253);
  nand ginst18098 (P2_U5299, P2_U3068, P2_U5251);
  nand ginst18099 (P2_U5300, P2_U3437, P2_U5253);
  nand ginst18100 (P2_U5301, P2_U3072, P2_U5251);
  nand ginst18101 (P2_U5302, P2_U3434, P2_U5253);
  nand ginst18102 (P2_U5303, P2_U3073, P2_U5251);
  nand ginst18103 (P2_U5304, P2_U3431, P2_U5253);
  nand ginst18104 (P2_U5305, P2_U3078, P2_U5251);
  nand ginst18105 (P2_U5306, P2_U3428, P2_U5253);
  nand ginst18106 (P2_U5307, P2_U3079, P2_U5251);
  nand ginst18107 (P2_U5308, P2_U3425, P2_U5253);
  nand ginst18108 (P2_U5309, P2_U3071, P2_U5251);
  nand ginst18109 (P2_U5310, P2_U3422, P2_U5253);
  nand ginst18110 (P2_U5311, P2_U3062, P2_U5251);
  nand ginst18111 (P2_U5312, P2_U3419, P2_U5253);
  nand ginst18112 (P2_U5313, P2_U3061, P2_U5251);
  nand ginst18113 (P2_U5314, P2_U3392, P2_U5253);
  nand ginst18114 (P2_U5315, P2_U3077, P2_U5251);
  nand ginst18115 (P2_U5316, P2_U3387, P2_U5253);
  nand ginst18116 (P2_U5317, P2_U3076, P2_U5251);
  nand ginst18117 (P2_U5318, P2_U3416, P2_U5251);
  nand ginst18118 (P2_U5319, P2_U3082, P2_U5253);
  nand ginst18119 (P2_U5320, P2_U3083, P2_U5436);
  nand ginst18120 (P2_U5321, P2_U3413, P2_U5251);
  nand ginst18121 (P2_U5322, P2_U3083, P2_U5253);
  nand ginst18122 (P2_U5323, P2_U3069, P2_U5436);
  nand ginst18123 (P2_U5324, P2_U3410, P2_U5251);
  nand ginst18124 (P2_U5325, P2_U3069, P2_U5253);
  nand ginst18125 (P2_U5326, P2_U3070, P2_U5436);
  nand ginst18126 (P2_U5327, P2_U3407, P2_U5251);
  nand ginst18127 (P2_U5328, P2_U3070, P2_U5253);
  nand ginst18128 (P2_U5329, P2_U3066, P2_U5436);
  nand ginst18129 (P2_U5330, P2_U3404, P2_U5251);
  nand ginst18130 (P2_U5331, P2_U3066, P2_U5253);
  nand ginst18131 (P2_U5332, P2_U3059, P2_U5436);
  nand ginst18132 (P2_U5333, P2_U3401, P2_U5251);
  nand ginst18133 (P2_U5334, P2_U3059, P2_U5253);
  nand ginst18134 (P2_U5335, P2_U3063, P2_U5436);
  nand ginst18135 (P2_U5336, P2_U3055, P2_U5253);
  nand ginst18136 (P2_U5337, P2_U3868, P2_U5251);
  nand ginst18137 (P2_U5338, P2_U3058, P2_U5253);
  nand ginst18138 (P2_U5339, P2_U3869, P2_U5251);
  nand ginst18139 (P2_U5340, P2_U3398, P2_U5251);
  nand ginst18140 (P2_U5341, P2_U3063, P2_U5253);
  nand ginst18141 (P2_U5342, P2_U3067, P2_U5436);
  nand ginst18142 (P2_U5343, P2_U3054, P2_U5253);
  nand ginst18143 (P2_U5344, P2_U3904, P2_U5251);
  nand ginst18144 (P2_U5345, P2_U3053, P2_U5436);
  nand ginst18145 (P2_U5346, P2_U3053, P2_U5253);
  nand ginst18146 (P2_U5347, P2_U3895, P2_U5251);
  nand ginst18147 (P2_U5348, P2_U3052, P2_U5436);
  nand ginst18148 (P2_U5349, P2_U3052, P2_U5253);
  nand ginst18149 (P2_U5350, P2_U3896, P2_U5251);
  nand ginst18150 (P2_U5351, P2_U3056, P2_U5436);
  nand ginst18151 (P2_U5352, P2_U3056, P2_U5253);
  nand ginst18152 (P2_U5353, P2_U3897, P2_U5251);
  nand ginst18153 (P2_U5354, P2_U3057, P2_U5436);
  nand ginst18154 (P2_U5355, P2_U3057, P2_U5253);
  nand ginst18155 (P2_U5356, P2_U3898, P2_U5251);
  nand ginst18156 (P2_U5357, P2_U3064, P2_U5436);
  nand ginst18157 (P2_U5358, P2_U3064, P2_U5253);
  nand ginst18158 (P2_U5359, P2_U3899, P2_U5251);
  nand ginst18159 (P2_U5360, P2_U3065, P2_U5436);
  nand ginst18160 (P2_U5361, P2_U3065, P2_U5253);
  nand ginst18161 (P2_U5362, P2_U3900, P2_U5251);
  nand ginst18162 (P2_U5363, P2_U3060, P2_U5436);
  nand ginst18163 (P2_U5364, P2_U3060, P2_U5253);
  nand ginst18164 (P2_U5365, P2_U3901, P2_U5251);
  nand ginst18165 (P2_U5366, P2_U3074, P2_U5436);
  nand ginst18166 (P2_U5367, P2_U3074, P2_U5253);
  nand ginst18167 (P2_U5368, P2_U3902, P2_U5251);
  nand ginst18168 (P2_U5369, P2_U3075, P2_U5436);
  nand ginst18169 (P2_U5370, P2_U3075, P2_U5253);
  nand ginst18170 (P2_U5371, P2_U3903, P2_U5251);
  nand ginst18171 (P2_U5372, P2_U3080, P2_U5436);
  nand ginst18172 (P2_U5373, P2_U3395, P2_U5251);
  nand ginst18173 (P2_U5374, P2_U3067, P2_U5253);
  nand ginst18174 (P2_U5375, P2_U3077, P2_U5436);
  nand ginst18175 (P2_U5376, P2_U3445, P2_U5251);
  nand ginst18176 (P2_U5377, P2_U3080, P2_U5253);
  nand ginst18177 (P2_U5378, P2_U3081, P2_U5436);
  nand ginst18178 (P2_U5379, P2_U3443, P2_U5251);
  nand ginst18179 (P2_U5380, P2_U3081, P2_U5253);
  nand ginst18180 (P2_U5381, P2_U3068, P2_U5436);
  nand ginst18181 (P2_U5382, P2_U3440, P2_U5251);
  nand ginst18182 (P2_U5383, P2_U3068, P2_U5253);
  nand ginst18183 (P2_U5384, P2_U3072, P2_U5436);
  nand ginst18184 (P2_U5385, P2_U3437, P2_U5251);
  nand ginst18185 (P2_U5386, P2_U3072, P2_U5253);
  nand ginst18186 (P2_U5387, P2_U3073, P2_U5436);
  nand ginst18187 (P2_U5388, P2_U3434, P2_U5251);
  nand ginst18188 (P2_U5389, P2_U3073, P2_U5253);
  nand ginst18189 (P2_U5390, P2_U3078, P2_U5436);
  nand ginst18190 (P2_U5391, P2_U3431, P2_U5251);
  nand ginst18191 (P2_U5392, P2_U3078, P2_U5253);
  nand ginst18192 (P2_U5393, P2_U3079, P2_U5436);
  nand ginst18193 (P2_U5394, P2_U3428, P2_U5251);
  nand ginst18194 (P2_U5395, P2_U3079, P2_U5253);
  nand ginst18195 (P2_U5396, P2_U3071, P2_U5436);
  nand ginst18196 (P2_U5397, P2_U3425, P2_U5251);
  nand ginst18197 (P2_U5398, P2_U3071, P2_U5253);
  nand ginst18198 (P2_U5399, P2_U3062, P2_U5436);
  nand ginst18199 (P2_U5400, P2_U3422, P2_U5251);
  nand ginst18200 (P2_U5401, P2_U3062, P2_U5253);
  nand ginst18201 (P2_U5402, P2_U3061, P2_U5436);
  nand ginst18202 (P2_U5403, P2_U3419, P2_U5251);
  nand ginst18203 (P2_U5404, P2_U3061, P2_U5253);
  nand ginst18204 (P2_U5405, P2_U3082, P2_U5436);
  nand ginst18205 (P2_U5406, P2_U3392, P2_U5251);
  nand ginst18206 (P2_U5407, P2_U3077, P2_U5253);
  nand ginst18207 (P2_U5408, P2_U3076, P2_U5436);
  nand ginst18208 (P2_U5409, P2_U3387, P2_U5251);
  nand ginst18209 (P2_U5410, P2_U3076, P2_U5253);
  nand ginst18210 (P2_U5411, P2_U3151, P2_U4977);
  nand ginst18211 (P2_U5412, P2_U4976, P2_U4977, P2_U5436);
  nand ginst18212 (P2_U5413, P2_U3043, P2_U3303);
  nand ginst18213 (P2_U5414, P2_U3043, P2_U3890);
  not ginst18214 (P2_U5415, P2_U3371);
  nand ginst18215 (P2_U5416, P2_U3914, P2_U5414);
  nand ginst18216 (P2_U5417, P2_U3779, P2_U5933, P2_U5934);
  nand ginst18217 (P2_U5418, P2_U5424, P2_U5430);
  nand ginst18218 (P2_U5419, P2_U3378, P2_U3875);
  nand ginst18219 (P2_U5420, P2_U3375, P2_U3829);
  nand ginst18220 (P2_U5421, P2_U3872, P2_U5443);
  nand ginst18221 (P2_U5422, P2_IR_REG_24__SCAN_IN, P2_U3827);
  nand ginst18222 (P2_U5423, P2_IR_REG_31__SCAN_IN, P2_SUB_594_U19);
  not ginst18223 (P2_U5424, P2_U3372);
  nand ginst18224 (P2_U5425, P2_IR_REG_25__SCAN_IN, P2_U3827);
  nand ginst18225 (P2_U5426, P2_IR_REG_31__SCAN_IN, P2_SUB_594_U79);
  not ginst18226 (P2_U5427, P2_U3373);
  nand ginst18227 (P2_U5428, P2_IR_REG_26__SCAN_IN, P2_U3827);
  nand ginst18228 (P2_U5429, P2_IR_REG_31__SCAN_IN, P2_SUB_594_U20);
  not ginst18229 (P2_U5430, P2_U3374);
  nand ginst18230 (P2_U5431, P2_B_REG_SCAN_IN, P2_U5424);
  nand ginst18231 (P2_U5432, P2_U3298, P2_U3372);
  nand ginst18232 (P2_U5433, P2_U5431, P2_U5432);
  nand ginst18233 (P2_U5434, P2_IR_REG_23__SCAN_IN, P2_U3827);
  nand ginst18234 (P2_U5435, P2_IR_REG_31__SCAN_IN, P2_SUB_594_U18);
  not ginst18235 (P2_U5436, P2_U3375);
  nand ginst18236 (P2_U5437, P2_D_REG_0__SCAN_IN, P2_U3828);
  nand ginst18237 (P2_U5438, P2_U3911, P2_U4016);
  nand ginst18238 (P2_U5439, P2_D_REG_1__SCAN_IN, P2_U3828);
  nand ginst18239 (P2_U5440, P2_U3911, P2_U4017);
  nand ginst18240 (P2_U5441, P2_IR_REG_20__SCAN_IN, P2_U3827);
  nand ginst18241 (P2_U5442, P2_IR_REG_31__SCAN_IN, P2_SUB_594_U16);
  not ginst18242 (P2_U5443, P2_U3378);
  nand ginst18243 (P2_U5444, P2_IR_REG_19__SCAN_IN, P2_U3827);
  nand ginst18244 (P2_U5445, P2_IR_REG_31__SCAN_IN, P2_SUB_594_U15);
  not ginst18245 (P2_U5446, P2_U3379);
  nand ginst18246 (P2_U5447, P2_IR_REG_22__SCAN_IN, P2_U3827);
  nand ginst18247 (P2_U5448, P2_IR_REG_31__SCAN_IN, P2_SUB_594_U17);
  not ginst18248 (P2_U5449, P2_U3380);
  nand ginst18249 (P2_U5450, P2_IR_REG_21__SCAN_IN, P2_U3827);
  nand ginst18250 (P2_U5451, P2_IR_REG_31__SCAN_IN, P2_SUB_594_U81);
  not ginst18251 (P2_U5452, P2_U3385);
  nand ginst18252 (P2_U5453, P2_IR_REG_30__SCAN_IN, P2_U3827);
  nand ginst18253 (P2_U5454, P2_IR_REG_31__SCAN_IN, P2_SUB_594_U75);
  not ginst18254 (P2_U5455, P2_U3381);
  nand ginst18255 (P2_U5456, P2_IR_REG_29__SCAN_IN, P2_U3827);
  nand ginst18256 (P2_U5457, P2_IR_REG_31__SCAN_IN, P2_SUB_594_U22);
  not ginst18257 (P2_U5458, P2_U3382);
  nand ginst18258 (P2_U5459, P2_IR_REG_28__SCAN_IN, P2_U3827);
  nand ginst18259 (P2_U5460, P2_IR_REG_31__SCAN_IN, P2_SUB_594_U21);
  not ginst18260 (P2_U5461, P2_U3383);
  nand ginst18261 (P2_U5462, P2_IR_REG_27__SCAN_IN, P2_U3827);
  nand ginst18262 (P2_U5463, P2_IR_REG_31__SCAN_IN, P2_SUB_594_U77);
  not ginst18263 (P2_U5464, P2_U3384);
  nand ginst18264 (P2_U5465, P2_IR_REG_0__SCAN_IN, P2_U3827);
  nand ginst18265 (P2_U5466, P2_IR_REG_0__SCAN_IN, P2_IR_REG_31__SCAN_IN);
  nand ginst18266 (P2_U5467, P2_U3829, U56);
  nand ginst18267 (P2_U5468, P2_U3386, P2_U3889);
  not ginst18268 (P2_U5469, P2_U3387);
  nand ginst18269 (P2_U5470, P2_U3300, P2_U5418);
  nand ginst18270 (P2_U5471, P2_D_REG_0__SCAN_IN, P2_U4015);
  not ginst18271 (P2_U5472, P2_U3388);
  nand ginst18272 (P2_U5473, P2_D_REG_1__SCAN_IN, P2_U4015);
  nand ginst18273 (P2_U5474, P2_U3300, P2_U4017);
  not ginst18274 (P2_U5475, P2_U3389);
  nand ginst18275 (P2_U5476, P2_U4048, P2_U5449);
  nand ginst18276 (P2_U5477, P2_U3380, P2_U3830);
  nand ginst18277 (P2_U5478, P2_U5476, P2_U5477);
  nand ginst18278 (P2_U5479, P2_REG0_REG_0__SCAN_IN, P2_U3831);
  nand ginst18279 (P2_U5480, P2_U3910, P2_U4073);
  nand ginst18280 (P2_U5481, P2_IR_REG_1__SCAN_IN, P2_U3827);
  nand ginst18281 (P2_U5482, P2_IR_REG_31__SCAN_IN, P2_SUB_594_U53);
  nand ginst18282 (P2_U5483, P2_U3829, U45);
  nand ginst18283 (P2_U5484, P2_U3391, P2_U3889);
  not ginst18284 (P2_U5485, P2_U3392);
  nand ginst18285 (P2_U5486, P2_REG0_REG_1__SCAN_IN, P2_U3831);
  nand ginst18286 (P2_U5487, P2_U3910, P2_U4098);
  nand ginst18287 (P2_U5488, P2_IR_REG_2__SCAN_IN, P2_U3827);
  nand ginst18288 (P2_U5489, P2_IR_REG_31__SCAN_IN, P2_SUB_594_U23);
  nand ginst18289 (P2_U5490, P2_U3829, U34);
  nand ginst18290 (P2_U5491, P2_U3394, P2_U3889);
  not ginst18291 (P2_U5492, P2_U3395);
  nand ginst18292 (P2_U5493, P2_REG0_REG_2__SCAN_IN, P2_U3831);
  nand ginst18293 (P2_U5494, P2_U3910, P2_U4116);
  nand ginst18294 (P2_U5495, P2_IR_REG_3__SCAN_IN, P2_U3827);
  nand ginst18295 (P2_U5496, P2_IR_REG_31__SCAN_IN, P2_SUB_594_U24);
  nand ginst18296 (P2_U5497, P2_U3829, U31);
  nand ginst18297 (P2_U5498, P2_U3397, P2_U3889);
  not ginst18298 (P2_U5499, P2_U3398);
  nand ginst18299 (P2_U5500, P2_REG0_REG_3__SCAN_IN, P2_U3831);
  nand ginst18300 (P2_U5501, P2_U3910, P2_U4134);
  nand ginst18301 (P2_U5502, P2_IR_REG_4__SCAN_IN, P2_U3827);
  nand ginst18302 (P2_U5503, P2_IR_REG_31__SCAN_IN, P2_SUB_594_U25);
  nand ginst18303 (P2_U5504, P2_U3829, U30);
  nand ginst18304 (P2_U5505, P2_U3400, P2_U3889);
  not ginst18305 (P2_U5506, P2_U3401);
  nand ginst18306 (P2_U5507, P2_REG0_REG_4__SCAN_IN, P2_U3831);
  nand ginst18307 (P2_U5508, P2_U3910, P2_U4152);
  nand ginst18308 (P2_U5509, P2_IR_REG_5__SCAN_IN, P2_U3827);
  nand ginst18309 (P2_U5510, P2_IR_REG_31__SCAN_IN, P2_SUB_594_U72);
  nand ginst18310 (P2_U5511, P2_U3829, U29);
  nand ginst18311 (P2_U5512, P2_U3403, P2_U3889);
  not ginst18312 (P2_U5513, P2_U3404);
  nand ginst18313 (P2_U5514, P2_REG0_REG_5__SCAN_IN, P2_U3831);
  nand ginst18314 (P2_U5515, P2_U3910, P2_U4170);
  nand ginst18315 (P2_U5516, P2_IR_REG_6__SCAN_IN, P2_U3827);
  nand ginst18316 (P2_U5517, P2_IR_REG_31__SCAN_IN, P2_SUB_594_U26);
  nand ginst18317 (P2_U5518, P2_U3829, U28);
  nand ginst18318 (P2_U5519, P2_U3406, P2_U3889);
  not ginst18319 (P2_U5520, P2_U3407);
  nand ginst18320 (P2_U5521, P2_REG0_REG_6__SCAN_IN, P2_U3831);
  nand ginst18321 (P2_U5522, P2_U3910, P2_U4188);
  nand ginst18322 (P2_U5523, P2_IR_REG_7__SCAN_IN, P2_U3827);
  nand ginst18323 (P2_U5524, P2_IR_REG_31__SCAN_IN, P2_SUB_594_U27);
  nand ginst18324 (P2_U5525, P2_U3829, U27);
  nand ginst18325 (P2_U5526, P2_U3409, P2_U3889);
  not ginst18326 (P2_U5527, P2_U3410);
  nand ginst18327 (P2_U5528, P2_REG0_REG_7__SCAN_IN, P2_U3831);
  nand ginst18328 (P2_U5529, P2_U3910, P2_U4206);
  nand ginst18329 (P2_U5530, P2_IR_REG_8__SCAN_IN, P2_U3827);
  nand ginst18330 (P2_U5531, P2_IR_REG_31__SCAN_IN, P2_SUB_594_U28);
  nand ginst18331 (P2_U5532, P2_U3829, U26);
  nand ginst18332 (P2_U5533, P2_U3412, P2_U3889);
  not ginst18333 (P2_U5534, P2_U3413);
  nand ginst18334 (P2_U5535, P2_REG0_REG_8__SCAN_IN, P2_U3831);
  nand ginst18335 (P2_U5536, P2_U3910, P2_U4224);
  nand ginst18336 (P2_U5537, P2_IR_REG_9__SCAN_IN, P2_U3827);
  nand ginst18337 (P2_U5538, P2_IR_REG_31__SCAN_IN, P2_SUB_594_U70);
  nand ginst18338 (P2_U5539, P2_U3829, U25);
  nand ginst18339 (P2_U5540, P2_U3415, P2_U3889);
  not ginst18340 (P2_U5541, P2_U3416);
  nand ginst18341 (P2_U5542, P2_REG0_REG_9__SCAN_IN, P2_U3831);
  nand ginst18342 (P2_U5543, P2_U3910, P2_U4242);
  nand ginst18343 (P2_U5544, P2_IR_REG_10__SCAN_IN, P2_U3827);
  nand ginst18344 (P2_U5545, P2_IR_REG_31__SCAN_IN, P2_SUB_594_U8);
  nand ginst18345 (P2_U5546, P2_U3829, U55);
  nand ginst18346 (P2_U5547, P2_U3418, P2_U3889);
  not ginst18347 (P2_U5548, P2_U3419);
  nand ginst18348 (P2_U5549, P2_REG0_REG_10__SCAN_IN, P2_U3831);
  nand ginst18349 (P2_U5550, P2_U3910, P2_U4260);
  nand ginst18350 (P2_U5551, P2_IR_REG_11__SCAN_IN, P2_U3827);
  nand ginst18351 (P2_U5552, P2_IR_REG_31__SCAN_IN, P2_SUB_594_U9);
  nand ginst18352 (P2_U5553, P2_U3829, U54);
  nand ginst18353 (P2_U5554, P2_U3421, P2_U3889);
  not ginst18354 (P2_U5555, P2_U3422);
  nand ginst18355 (P2_U5556, P2_REG0_REG_11__SCAN_IN, P2_U3831);
  nand ginst18356 (P2_U5557, P2_U3910, P2_U4278);
  nand ginst18357 (P2_U5558, P2_IR_REG_12__SCAN_IN, P2_U3827);
  nand ginst18358 (P2_U5559, P2_IR_REG_31__SCAN_IN, P2_SUB_594_U10);
  nand ginst18359 (P2_U5560, P2_U3829, U53);
  nand ginst18360 (P2_U5561, P2_U3424, P2_U3889);
  not ginst18361 (P2_U5562, P2_U3425);
  nand ginst18362 (P2_U5563, P2_REG0_REG_12__SCAN_IN, P2_U3831);
  nand ginst18363 (P2_U5564, P2_U3910, P2_U4296);
  nand ginst18364 (P2_U5565, P2_IR_REG_13__SCAN_IN, P2_U3827);
  nand ginst18365 (P2_U5566, P2_IR_REG_31__SCAN_IN, P2_SUB_594_U87);
  nand ginst18366 (P2_U5567, P2_U3829, U52);
  nand ginst18367 (P2_U5568, P2_U3427, P2_U3889);
  not ginst18368 (P2_U5569, P2_U3428);
  nand ginst18369 (P2_U5570, P2_REG0_REG_13__SCAN_IN, P2_U3831);
  nand ginst18370 (P2_U5571, P2_U3910, P2_U4314);
  nand ginst18371 (P2_U5572, P2_IR_REG_14__SCAN_IN, P2_U3827);
  nand ginst18372 (P2_U5573, P2_IR_REG_31__SCAN_IN, P2_SUB_594_U11);
  nand ginst18373 (P2_U5574, P2_U3829, U51);
  nand ginst18374 (P2_U5575, P2_U3430, P2_U3889);
  not ginst18375 (P2_U5576, P2_U3431);
  nand ginst18376 (P2_U5577, P2_REG0_REG_14__SCAN_IN, P2_U3831);
  nand ginst18377 (P2_U5578, P2_U3910, P2_U4332);
  nand ginst18378 (P2_U5579, P2_IR_REG_15__SCAN_IN, P2_U3827);
  nand ginst18379 (P2_U5580, P2_IR_REG_31__SCAN_IN, P2_SUB_594_U12);
  nand ginst18380 (P2_U5581, P2_U3829, U50);
  nand ginst18381 (P2_U5582, P2_U3433, P2_U3889);
  not ginst18382 (P2_U5583, P2_U3434);
  nand ginst18383 (P2_U5584, P2_REG0_REG_15__SCAN_IN, P2_U3831);
  nand ginst18384 (P2_U5585, P2_U3910, P2_U4350);
  nand ginst18385 (P2_U5586, P2_IR_REG_16__SCAN_IN, P2_U3827);
  nand ginst18386 (P2_U5587, P2_IR_REG_31__SCAN_IN, P2_SUB_594_U13);
  nand ginst18387 (P2_U5588, P2_U3829, U49);
  nand ginst18388 (P2_U5589, P2_U3436, P2_U3889);
  not ginst18389 (P2_U5590, P2_U3437);
  nand ginst18390 (P2_U5591, P2_REG0_REG_16__SCAN_IN, P2_U3831);
  nand ginst18391 (P2_U5592, P2_U3910, P2_U4368);
  nand ginst18392 (P2_U5593, P2_IR_REG_17__SCAN_IN, P2_U3827);
  nand ginst18393 (P2_U5594, P2_IR_REG_31__SCAN_IN, P2_SUB_594_U85);
  nand ginst18394 (P2_U5595, P2_U3829, U48);
  nand ginst18395 (P2_U5596, P2_U3439, P2_U3889);
  not ginst18396 (P2_U5597, P2_U3440);
  nand ginst18397 (P2_U5598, P2_REG0_REG_17__SCAN_IN, P2_U3831);
  nand ginst18398 (P2_U5599, P2_U3910, P2_U4386);
  nand ginst18399 (P2_U5600, P2_IR_REG_18__SCAN_IN, P2_U3827);
  nand ginst18400 (P2_U5601, P2_IR_REG_31__SCAN_IN, P2_SUB_594_U14);
  nand ginst18401 (P2_U5602, P2_U3829, U47);
  nand ginst18402 (P2_U5603, P2_U3442, P2_U3889);
  not ginst18403 (P2_U5604, P2_U3443);
  nand ginst18404 (P2_U5605, P2_REG0_REG_18__SCAN_IN, P2_U3831);
  nand ginst18405 (P2_U5606, P2_U3910, P2_U4404);
  nand ginst18406 (P2_U5607, P2_U3829, U46);
  nand ginst18407 (P2_U5608, P2_U3379, P2_U3889);
  not ginst18408 (P2_U5609, P2_U3445);
  nand ginst18409 (P2_U5610, P2_REG0_REG_19__SCAN_IN, P2_U3831);
  nand ginst18410 (P2_U5611, P2_U3910, P2_U4422);
  nand ginst18411 (P2_U5612, P2_REG0_REG_20__SCAN_IN, P2_U3831);
  nand ginst18412 (P2_U5613, P2_U3910, P2_U4440);
  nand ginst18413 (P2_U5614, P2_REG0_REG_21__SCAN_IN, P2_U3831);
  nand ginst18414 (P2_U5615, P2_U3910, P2_U4458);
  nand ginst18415 (P2_U5616, P2_REG0_REG_22__SCAN_IN, P2_U3831);
  nand ginst18416 (P2_U5617, P2_U3910, P2_U4476);
  nand ginst18417 (P2_U5618, P2_REG0_REG_23__SCAN_IN, P2_U3831);
  nand ginst18418 (P2_U5619, P2_U3910, P2_U4494);
  nand ginst18419 (P2_U5620, P2_REG0_REG_24__SCAN_IN, P2_U3831);
  nand ginst18420 (P2_U5621, P2_U3910, P2_U4512);
  nand ginst18421 (P2_U5622, P2_REG0_REG_25__SCAN_IN, P2_U3831);
  nand ginst18422 (P2_U5623, P2_U3910, P2_U4530);
  nand ginst18423 (P2_U5624, P2_REG0_REG_26__SCAN_IN, P2_U3831);
  nand ginst18424 (P2_U5625, P2_U3910, P2_U4548);
  nand ginst18425 (P2_U5626, P2_REG0_REG_27__SCAN_IN, P2_U3831);
  nand ginst18426 (P2_U5627, P2_U3910, P2_U4566);
  nand ginst18427 (P2_U5628, P2_REG0_REG_28__SCAN_IN, P2_U3831);
  nand ginst18428 (P2_U5629, P2_U3910, P2_U4584);
  nand ginst18429 (P2_U5630, P2_REG0_REG_29__SCAN_IN, P2_U3831);
  nand ginst18430 (P2_U5631, P2_U3910, P2_U4604);
  nand ginst18431 (P2_U5632, P2_REG0_REG_30__SCAN_IN, P2_U3831);
  nand ginst18432 (P2_U5633, P2_U3910, P2_U4611);
  nand ginst18433 (P2_U5634, P2_REG0_REG_31__SCAN_IN, P2_U3831);
  nand ginst18434 (P2_U5635, P2_U3910, P2_U4613);
  nand ginst18435 (P2_U5636, P2_U3830, P2_U5449);
  nand ginst18436 (P2_U5637, P2_U4048, P2_U5446);
  nand ginst18437 (P2_U5638, P2_REG1_REG_0__SCAN_IN, P2_U3832);
  nand ginst18438 (P2_U5639, P2_U3909, P2_U4073);
  nand ginst18439 (P2_U5640, P2_REG1_REG_1__SCAN_IN, P2_U3832);
  nand ginst18440 (P2_U5641, P2_U3909, P2_U4098);
  nand ginst18441 (P2_U5642, P2_REG1_REG_2__SCAN_IN, P2_U3832);
  nand ginst18442 (P2_U5643, P2_U3909, P2_U4116);
  nand ginst18443 (P2_U5644, P2_REG1_REG_3__SCAN_IN, P2_U3832);
  nand ginst18444 (P2_U5645, P2_U3909, P2_U4134);
  nand ginst18445 (P2_U5646, P2_REG1_REG_4__SCAN_IN, P2_U3832);
  nand ginst18446 (P2_U5647, P2_U3909, P2_U4152);
  nand ginst18447 (P2_U5648, P2_REG1_REG_5__SCAN_IN, P2_U3832);
  nand ginst18448 (P2_U5649, P2_U3909, P2_U4170);
  nand ginst18449 (P2_U5650, P2_REG1_REG_6__SCAN_IN, P2_U3832);
  nand ginst18450 (P2_U5651, P2_U3909, P2_U4188);
  nand ginst18451 (P2_U5652, P2_REG1_REG_7__SCAN_IN, P2_U3832);
  nand ginst18452 (P2_U5653, P2_U3909, P2_U4206);
  nand ginst18453 (P2_U5654, P2_REG1_REG_8__SCAN_IN, P2_U3832);
  nand ginst18454 (P2_U5655, P2_U3909, P2_U4224);
  nand ginst18455 (P2_U5656, P2_REG1_REG_9__SCAN_IN, P2_U3832);
  nand ginst18456 (P2_U5657, P2_U3909, P2_U4242);
  nand ginst18457 (P2_U5658, P2_REG1_REG_10__SCAN_IN, P2_U3832);
  nand ginst18458 (P2_U5659, P2_U3909, P2_U4260);
  nand ginst18459 (P2_U5660, P2_REG1_REG_11__SCAN_IN, P2_U3832);
  nand ginst18460 (P2_U5661, P2_U3909, P2_U4278);
  nand ginst18461 (P2_U5662, P2_REG1_REG_12__SCAN_IN, P2_U3832);
  nand ginst18462 (P2_U5663, P2_U3909, P2_U4296);
  nand ginst18463 (P2_U5664, P2_REG1_REG_13__SCAN_IN, P2_U3832);
  nand ginst18464 (P2_U5665, P2_U3909, P2_U4314);
  nand ginst18465 (P2_U5666, P2_REG1_REG_14__SCAN_IN, P2_U3832);
  nand ginst18466 (P2_U5667, P2_U3909, P2_U4332);
  nand ginst18467 (P2_U5668, P2_REG1_REG_15__SCAN_IN, P2_U3832);
  nand ginst18468 (P2_U5669, P2_U3909, P2_U4350);
  nand ginst18469 (P2_U5670, P2_REG1_REG_16__SCAN_IN, P2_U3832);
  nand ginst18470 (P2_U5671, P2_U3909, P2_U4368);
  nand ginst18471 (P2_U5672, P2_REG1_REG_17__SCAN_IN, P2_U3832);
  nand ginst18472 (P2_U5673, P2_U3909, P2_U4386);
  nand ginst18473 (P2_U5674, P2_REG1_REG_18__SCAN_IN, P2_U3832);
  nand ginst18474 (P2_U5675, P2_U3909, P2_U4404);
  nand ginst18475 (P2_U5676, P2_REG1_REG_19__SCAN_IN, P2_U3832);
  nand ginst18476 (P2_U5677, P2_U3909, P2_U4422);
  nand ginst18477 (P2_U5678, P2_REG1_REG_20__SCAN_IN, P2_U3832);
  nand ginst18478 (P2_U5679, P2_U3909, P2_U4440);
  nand ginst18479 (P2_U5680, P2_REG1_REG_21__SCAN_IN, P2_U3832);
  nand ginst18480 (P2_U5681, P2_U3909, P2_U4458);
  nand ginst18481 (P2_U5682, P2_REG1_REG_22__SCAN_IN, P2_U3832);
  nand ginst18482 (P2_U5683, P2_U3909, P2_U4476);
  nand ginst18483 (P2_U5684, P2_REG1_REG_23__SCAN_IN, P2_U3832);
  nand ginst18484 (P2_U5685, P2_U3909, P2_U4494);
  nand ginst18485 (P2_U5686, P2_REG1_REG_24__SCAN_IN, P2_U3832);
  nand ginst18486 (P2_U5687, P2_U3909, P2_U4512);
  nand ginst18487 (P2_U5688, P2_REG1_REG_25__SCAN_IN, P2_U3832);
  nand ginst18488 (P2_U5689, P2_U3909, P2_U4530);
  nand ginst18489 (P2_U5690, P2_REG1_REG_26__SCAN_IN, P2_U3832);
  nand ginst18490 (P2_U5691, P2_U3909, P2_U4548);
  nand ginst18491 (P2_U5692, P2_REG1_REG_27__SCAN_IN, P2_U3832);
  nand ginst18492 (P2_U5693, P2_U3909, P2_U4566);
  nand ginst18493 (P2_U5694, P2_REG1_REG_28__SCAN_IN, P2_U3832);
  nand ginst18494 (P2_U5695, P2_U3909, P2_U4584);
  nand ginst18495 (P2_U5696, P2_REG1_REG_29__SCAN_IN, P2_U3832);
  nand ginst18496 (P2_U5697, P2_U3909, P2_U4604);
  nand ginst18497 (P2_U5698, P2_REG1_REG_30__SCAN_IN, P2_U3832);
  nand ginst18498 (P2_U5699, P2_U3909, P2_U4611);
  nand ginst18499 (P2_U5700, P2_REG1_REG_31__SCAN_IN, P2_U3832);
  nand ginst18500 (P2_U5701, P2_U3909, P2_U4613);
  nand ginst18501 (P2_U5702, P2_REG2_REG_0__SCAN_IN, P2_U3358);
  nand ginst18502 (P2_U5703, P2_U3314, P2_U3908);
  nand ginst18503 (P2_U5704, P2_REG2_REG_1__SCAN_IN, P2_U3358);
  nand ginst18504 (P2_U5705, P2_U3315, P2_U3908);
  nand ginst18505 (P2_U5706, P2_REG2_REG_2__SCAN_IN, P2_U3358);
  nand ginst18506 (P2_U5707, P2_U3316, P2_U3908);
  nand ginst18507 (P2_U5708, P2_REG2_REG_3__SCAN_IN, P2_U3358);
  nand ginst18508 (P2_U5709, P2_U3317, P2_U3908);
  nand ginst18509 (P2_U5710, P2_REG2_REG_4__SCAN_IN, P2_U3358);
  nand ginst18510 (P2_U5711, P2_U3318, P2_U3908);
  nand ginst18511 (P2_U5712, P2_REG2_REG_5__SCAN_IN, P2_U3358);
  nand ginst18512 (P2_U5713, P2_U3319, P2_U3908);
  nand ginst18513 (P2_U5714, P2_REG2_REG_6__SCAN_IN, P2_U3358);
  nand ginst18514 (P2_U5715, P2_U3320, P2_U3908);
  nand ginst18515 (P2_U5716, P2_REG2_REG_7__SCAN_IN, P2_U3358);
  nand ginst18516 (P2_U5717, P2_U3321, P2_U3908);
  nand ginst18517 (P2_U5718, P2_REG2_REG_8__SCAN_IN, P2_U3358);
  nand ginst18518 (P2_U5719, P2_U3322, P2_U3908);
  nand ginst18519 (P2_U5720, P2_REG2_REG_9__SCAN_IN, P2_U3358);
  nand ginst18520 (P2_U5721, P2_U3323, P2_U3908);
  nand ginst18521 (P2_U5722, P2_REG2_REG_10__SCAN_IN, P2_U3358);
  nand ginst18522 (P2_U5723, P2_U3324, P2_U3908);
  nand ginst18523 (P2_U5724, P2_REG2_REG_11__SCAN_IN, P2_U3358);
  nand ginst18524 (P2_U5725, P2_U3325, P2_U3908);
  nand ginst18525 (P2_U5726, P2_REG2_REG_12__SCAN_IN, P2_U3358);
  nand ginst18526 (P2_U5727, P2_U3326, P2_U3908);
  nand ginst18527 (P2_U5728, P2_REG2_REG_13__SCAN_IN, P2_U3358);
  nand ginst18528 (P2_U5729, P2_U3327, P2_U3908);
  nand ginst18529 (P2_U5730, P2_REG2_REG_14__SCAN_IN, P2_U3358);
  nand ginst18530 (P2_U5731, P2_U3328, P2_U3908);
  nand ginst18531 (P2_U5732, P2_REG2_REG_15__SCAN_IN, P2_U3358);
  nand ginst18532 (P2_U5733, P2_U3329, P2_U3908);
  nand ginst18533 (P2_U5734, P2_REG2_REG_16__SCAN_IN, P2_U3358);
  nand ginst18534 (P2_U5735, P2_U3330, P2_U3908);
  nand ginst18535 (P2_U5736, P2_REG2_REG_17__SCAN_IN, P2_U3358);
  nand ginst18536 (P2_U5737, P2_U3331, P2_U3908);
  nand ginst18537 (P2_U5738, P2_REG2_REG_18__SCAN_IN, P2_U3358);
  nand ginst18538 (P2_U5739, P2_U3332, P2_U3908);
  nand ginst18539 (P2_U5740, P2_REG2_REG_19__SCAN_IN, P2_U3358);
  nand ginst18540 (P2_U5741, P2_U3333, P2_U3908);
  nand ginst18541 (P2_U5742, P2_REG2_REG_20__SCAN_IN, P2_U3358);
  nand ginst18542 (P2_U5743, P2_U3335, P2_U3908);
  nand ginst18543 (P2_U5744, P2_REG2_REG_21__SCAN_IN, P2_U3358);
  nand ginst18544 (P2_U5745, P2_U3337, P2_U3908);
  nand ginst18545 (P2_U5746, P2_REG2_REG_22__SCAN_IN, P2_U3358);
  nand ginst18546 (P2_U5747, P2_U3339, P2_U3908);
  nand ginst18547 (P2_U5748, P2_REG2_REG_23__SCAN_IN, P2_U3358);
  nand ginst18548 (P2_U5749, P2_U3341, P2_U3908);
  nand ginst18549 (P2_U5750, P2_REG2_REG_24__SCAN_IN, P2_U3358);
  nand ginst18550 (P2_U5751, P2_U3343, P2_U3908);
  nand ginst18551 (P2_U5752, P2_REG2_REG_25__SCAN_IN, P2_U3358);
  nand ginst18552 (P2_U5753, P2_U3345, P2_U3908);
  nand ginst18553 (P2_U5754, P2_REG2_REG_26__SCAN_IN, P2_U3358);
  nand ginst18554 (P2_U5755, P2_U3347, P2_U3908);
  nand ginst18555 (P2_U5756, P2_REG2_REG_27__SCAN_IN, P2_U3358);
  nand ginst18556 (P2_U5757, P2_U3349, P2_U3908);
  nand ginst18557 (P2_U5758, P2_REG2_REG_28__SCAN_IN, P2_U3358);
  nand ginst18558 (P2_U5759, P2_U3351, P2_U3908);
  nand ginst18559 (P2_U5760, P2_REG2_REG_29__SCAN_IN, P2_U3358);
  nand ginst18560 (P2_U5761, P2_U3354, P2_U3908);
  nand ginst18561 (P2_U5762, P2_U3024, P2_U5461);
  nand ginst18562 (P2_U5763, P2_U3383, P2_U3893);
  nand ginst18563 (P2_U5764, P2_U5762, P2_U5763);
  nand ginst18564 (P2_U5765, P2_DATAO_REG_0__SCAN_IN, P2_U3363);
  nand ginst18565 (P2_U5766, P2_U3076, P2_U3893);
  nand ginst18566 (P2_U5767, P2_DATAO_REG_1__SCAN_IN, P2_U3363);
  nand ginst18567 (P2_U5768, P2_U3077, P2_U3893);
  nand ginst18568 (P2_U5769, P2_DATAO_REG_2__SCAN_IN, P2_U3363);
  nand ginst18569 (P2_U5770, P2_U3067, P2_U3893);
  nand ginst18570 (P2_U5771, P2_DATAO_REG_3__SCAN_IN, P2_U3363);
  nand ginst18571 (P2_U5772, P2_U3063, P2_U3893);
  nand ginst18572 (P2_U5773, P2_DATAO_REG_4__SCAN_IN, P2_U3363);
  nand ginst18573 (P2_U5774, P2_U3059, P2_U3893);
  nand ginst18574 (P2_U5775, P2_DATAO_REG_5__SCAN_IN, P2_U3363);
  nand ginst18575 (P2_U5776, P2_U3066, P2_U3893);
  nand ginst18576 (P2_U5777, P2_DATAO_REG_6__SCAN_IN, P2_U3363);
  nand ginst18577 (P2_U5778, P2_U3070, P2_U3893);
  nand ginst18578 (P2_U5779, P2_DATAO_REG_7__SCAN_IN, P2_U3363);
  nand ginst18579 (P2_U5780, P2_U3069, P2_U3893);
  nand ginst18580 (P2_U5781, P2_DATAO_REG_8__SCAN_IN, P2_U3363);
  nand ginst18581 (P2_U5782, P2_U3083, P2_U3893);
  nand ginst18582 (P2_U5783, P2_DATAO_REG_9__SCAN_IN, P2_U3363);
  nand ginst18583 (P2_U5784, P2_U3082, P2_U3893);
  nand ginst18584 (P2_U5785, P2_DATAO_REG_10__SCAN_IN, P2_U3363);
  nand ginst18585 (P2_U5786, P2_U3061, P2_U3893);
  nand ginst18586 (P2_U5787, P2_DATAO_REG_11__SCAN_IN, P2_U3363);
  nand ginst18587 (P2_U5788, P2_U3062, P2_U3893);
  nand ginst18588 (P2_U5789, P2_DATAO_REG_12__SCAN_IN, P2_U3363);
  nand ginst18589 (P2_U5790, P2_U3071, P2_U3893);
  nand ginst18590 (P2_U5791, P2_DATAO_REG_13__SCAN_IN, P2_U3363);
  nand ginst18591 (P2_U5792, P2_U3079, P2_U3893);
  nand ginst18592 (P2_U5793, P2_DATAO_REG_14__SCAN_IN, P2_U3363);
  nand ginst18593 (P2_U5794, P2_U3078, P2_U3893);
  nand ginst18594 (P2_U5795, P2_DATAO_REG_15__SCAN_IN, P2_U3363);
  nand ginst18595 (P2_U5796, P2_U3073, P2_U3893);
  nand ginst18596 (P2_U5797, P2_DATAO_REG_16__SCAN_IN, P2_U3363);
  nand ginst18597 (P2_U5798, P2_U3072, P2_U3893);
  nand ginst18598 (P2_U5799, P2_DATAO_REG_17__SCAN_IN, P2_U3363);
  nand ginst18599 (P2_U5800, P2_U3068, P2_U3893);
  nand ginst18600 (P2_U5801, P2_DATAO_REG_18__SCAN_IN, P2_U3363);
  nand ginst18601 (P2_U5802, P2_U3081, P2_U3893);
  nand ginst18602 (P2_U5803, P2_DATAO_REG_19__SCAN_IN, P2_U3363);
  nand ginst18603 (P2_U5804, P2_U3080, P2_U3893);
  nand ginst18604 (P2_U5805, P2_DATAO_REG_20__SCAN_IN, P2_U3363);
  nand ginst18605 (P2_U5806, P2_U3075, P2_U3893);
  nand ginst18606 (P2_U5807, P2_DATAO_REG_21__SCAN_IN, P2_U3363);
  nand ginst18607 (P2_U5808, P2_U3074, P2_U3893);
  nand ginst18608 (P2_U5809, P2_DATAO_REG_22__SCAN_IN, P2_U3363);
  nand ginst18609 (P2_U5810, P2_U3060, P2_U3893);
  nand ginst18610 (P2_U5811, P2_DATAO_REG_23__SCAN_IN, P2_U3363);
  nand ginst18611 (P2_U5812, P2_U3065, P2_U3893);
  nand ginst18612 (P2_U5813, P2_DATAO_REG_24__SCAN_IN, P2_U3363);
  nand ginst18613 (P2_U5814, P2_U3064, P2_U3893);
  nand ginst18614 (P2_U5815, P2_DATAO_REG_25__SCAN_IN, P2_U3363);
  nand ginst18615 (P2_U5816, P2_U3057, P2_U3893);
  nand ginst18616 (P2_U5817, P2_DATAO_REG_26__SCAN_IN, P2_U3363);
  nand ginst18617 (P2_U5818, P2_U3056, P2_U3893);
  nand ginst18618 (P2_U5819, P2_DATAO_REG_27__SCAN_IN, P2_U3363);
  nand ginst18619 (P2_U5820, P2_U3052, P2_U3893);
  nand ginst18620 (P2_U5821, P2_DATAO_REG_28__SCAN_IN, P2_U3363);
  nand ginst18621 (P2_U5822, P2_U3053, P2_U3893);
  nand ginst18622 (P2_U5823, P2_DATAO_REG_29__SCAN_IN, P2_U3363);
  nand ginst18623 (P2_U5824, P2_U3054, P2_U3893);
  nand ginst18624 (P2_U5825, P2_DATAO_REG_30__SCAN_IN, P2_U3363);
  nand ginst18625 (P2_U5826, P2_U3058, P2_U3893);
  nand ginst18626 (P2_U5827, P2_DATAO_REG_31__SCAN_IN, P2_U3363);
  nand ginst18627 (P2_U5828, P2_U3055, P2_U3893);
  nand ginst18628 (P2_U5829, P2_U3313, P2_U3379);
  nand ginst18629 (P2_U5830, P2_U3907, P2_U5446);
  not ginst18630 (P2_U5831, P2_U3765);
  nand ginst18631 (P2_U5832, P2_R1269_U22, P2_U5831);
  nand ginst18632 (P2_U5833, P2_U3765, P2_U3863);
  nand ginst18633 (P2_U5834, P2_U3052, P2_U3896);
  nand ginst18634 (P2_U5835, P2_U3348, P2_U4535);
  nand ginst18635 (P2_U5836, P2_U5834, P2_U5835);
  nand ginst18636 (P2_U5837, P2_U3053, P2_U3895);
  nand ginst18637 (P2_U5838, P2_U3350, P2_U4553);
  nand ginst18638 (P2_U5839, P2_U5837, P2_U5838);
  nand ginst18639 (P2_U5840, P2_U3055, P2_U3868);
  nand ginst18640 (P2_U5841, P2_U3356, P2_U4609);
  nand ginst18641 (P2_U5842, P2_U5840, P2_U5841);
  nand ginst18642 (P2_U5843, P2_U3054, P2_U3904);
  nand ginst18643 (P2_U5844, P2_U3353, P2_U4571);
  nand ginst18644 (P2_U5845, P2_U5843, P2_U5844);
  nand ginst18645 (P2_U5846, P2_U3074, P2_U3902);
  nand ginst18646 (P2_U5847, P2_U3336, P2_U4427);
  nand ginst18647 (P2_U5848, P2_U5846, P2_U5847);
  nand ginst18648 (P2_U5849, P2_U3075, P2_U3903);
  nand ginst18649 (P2_U5850, P2_U3334, P2_U4409);
  nand ginst18650 (P2_U5851, P2_U5849, P2_U5850);
  nand ginst18651 (P2_U5852, P2_U4103, P2_U5499);
  nand ginst18652 (P2_U5853, P2_U3063, P2_U3398);
  nand ginst18653 (P2_U5854, P2_U5852, P2_U5853);
  nand ginst18654 (P2_U5855, P2_U4247, P2_U5555);
  nand ginst18655 (P2_U5856, P2_U3062, P2_U3422);
  nand ginst18656 (P2_U5857, P2_U5855, P2_U5856);
  nand ginst18657 (P2_U5858, P2_U4229, P2_U5548);
  nand ginst18658 (P2_U5859, P2_U3061, P2_U3419);
  nand ginst18659 (P2_U5860, P2_U5858, P2_U5859);
  nand ginst18660 (P2_U5861, P2_U4121, P2_U5506);
  nand ginst18661 (P2_U5862, P2_U3059, P2_U3401);
  nand ginst18662 (P2_U5863, P2_U5861, P2_U5862);
  nand ginst18663 (P2_U5864, P2_U3060, P2_U3901);
  nand ginst18664 (P2_U5865, P2_U3338, P2_U4445);
  nand ginst18665 (P2_U5866, P2_U5864, P2_U5865);
  nand ginst18666 (P2_U5867, P2_U4355, P2_U5597);
  nand ginst18667 (P2_U5868, P2_U3068, P2_U3440);
  nand ginst18668 (P2_U5869, P2_U5867, P2_U5868);
  nand ginst18669 (P2_U5870, P2_U4319, P2_U5583);
  nand ginst18670 (P2_U5871, P2_U3073, P2_U3434);
  nand ginst18671 (P2_U5872, P2_U5870, P2_U5871);
  nand ginst18672 (P2_U5873, P2_U4265, P2_U5562);
  nand ginst18673 (P2_U5874, P2_U3071, P2_U3425);
  nand ginst18674 (P2_U5875, P2_U5873, P2_U5874);
  nand ginst18675 (P2_U5876, P2_U4157, P2_U5520);
  nand ginst18676 (P2_U5877, P2_U3070, P2_U3407);
  nand ginst18677 (P2_U5878, P2_U5876, P2_U5877);
  nand ginst18678 (P2_U5879, P2_U4175, P2_U5527);
  nand ginst18679 (P2_U5880, P2_U3069, P2_U3410);
  nand ginst18680 (P2_U5881, P2_U5879, P2_U5880);
  nand ginst18681 (P2_U5882, P2_U4078, P2_U5492);
  nand ginst18682 (P2_U5883, P2_U3067, P2_U3395);
  nand ginst18683 (P2_U5884, P2_U5882, P2_U5883);
  nand ginst18684 (P2_U5885, P2_U4139, P2_U5513);
  nand ginst18685 (P2_U5886, P2_U3066, P2_U3404);
  nand ginst18686 (P2_U5887, P2_U5885, P2_U5886);
  nand ginst18687 (P2_U5888, P2_U4337, P2_U5590);
  nand ginst18688 (P2_U5889, P2_U3072, P2_U3437);
  nand ginst18689 (P2_U5890, P2_U5888, P2_U5889);
  nand ginst18690 (P2_U5891, P2_U4373, P2_U5604);
  nand ginst18691 (P2_U5892, P2_U3081, P2_U3443);
  nand ginst18692 (P2_U5893, P2_U5891, P2_U5892);
  nand ginst18693 (P2_U5894, P2_U4283, P2_U5569);
  nand ginst18694 (P2_U5895, P2_U3079, P2_U3428);
  nand ginst18695 (P2_U5896, P2_U5894, P2_U5895);
  nand ginst18696 (P2_U5897, P2_U4301, P2_U5576);
  nand ginst18697 (P2_U5898, P2_U3078, P2_U3431);
  nand ginst18698 (P2_U5899, P2_U5897, P2_U5898);
  nand ginst18699 (P2_U5900, P2_U4059, P2_U5485);
  nand ginst18700 (P2_U5901, P2_U3077, P2_U3392);
  nand ginst18701 (P2_U5902, P2_U5900, P2_U5901);
  nand ginst18702 (P2_U5903, P2_U4083, P2_U5469);
  nand ginst18703 (P2_U5904, P2_U3076, P2_U3387);
  nand ginst18704 (P2_U5905, P2_U5903, P2_U5904);
  nand ginst18705 (P2_U5906, P2_U4193, P2_U5534);
  nand ginst18706 (P2_U5907, P2_U3083, P2_U3413);
  nand ginst18707 (P2_U5908, P2_U5906, P2_U5907);
  nand ginst18708 (P2_U5909, P2_U4211, P2_U5541);
  nand ginst18709 (P2_U5910, P2_U3082, P2_U3416);
  nand ginst18710 (P2_U5911, P2_U5909, P2_U5910);
  nand ginst18711 (P2_U5912, P2_U4391, P2_U5609);
  nand ginst18712 (P2_U5913, P2_U3080, P2_U3445);
  nand ginst18713 (P2_U5914, P2_U5912, P2_U5913);
  nand ginst18714 (P2_U5915, P2_U3056, P2_U3897);
  nand ginst18715 (P2_U5916, P2_U3346, P2_U4517);
  nand ginst18716 (P2_U5917, P2_U5915, P2_U5916);
  nand ginst18717 (P2_U5918, P2_U3057, P2_U3898);
  nand ginst18718 (P2_U5919, P2_U3344, P2_U4499);
  nand ginst18719 (P2_U5920, P2_U5918, P2_U5919);
  nand ginst18720 (P2_U5921, P2_U3065, P2_U3900);
  nand ginst18721 (P2_U5922, P2_U3340, P2_U4463);
  nand ginst18722 (P2_U5923, P2_U5921, P2_U5922);
  nand ginst18723 (P2_U5924, P2_U3064, P2_U3899);
  nand ginst18724 (P2_U5925, P2_U3342, P2_U4481);
  nand ginst18725 (P2_U5926, P2_U5924, P2_U5925);
  nand ginst18726 (P2_U5927, P2_U3058, P2_U3869);
  nand ginst18727 (P2_U5928, P2_U3355, P2_U4589);
  nand ginst18728 (P2_U5929, P2_U5927, P2_U5928);
  nand ginst18729 (P2_U5930, P2_U4974, P2_U5446);
  nand ginst18730 (P2_U5931, P2_U3379, P2_U3864);
  nand ginst18731 (P2_U5932, P2_U5930, P2_U5931);
  nand ginst18732 (P2_U5933, P2_U5443, P2_U5832, P2_U5833);
  nand ginst18733 (P2_U5934, P2_U3378, P2_U5452, P2_U5932);
  nand ginst18734 (P2_U5935, P2_U3865, P2_U3877);
  nand ginst18735 (P2_U5936, P2_R693_U14, P2_U3887);
  nand ginst18736 (P2_U5937, P2_U3368, P2_U5436);
  nand ginst18737 (P2_U5938, P2_U3375, P2_U3380);
  nand ginst18738 (P2_U5939, P2_U5443, P2_U5446);
  nand ginst18739 (P2_U5940, P2_U3378, P2_U3388, P2_U5452);
  nand ginst18740 (P2_U5941, P2_R1297_U6, P2_U3082);
  nand ginst18741 (P2_U5942, P2_U3082, P2_U3867);
  nand ginst18742 (P2_U5943, P2_R1297_U6, P2_U3083);
  nand ginst18743 (P2_U5944, P2_U3083, P2_U3867);
  nand ginst18744 (P2_U5945, P2_R1297_U6, P2_U3069);
  nand ginst18745 (P2_U5946, P2_U3069, P2_U3867);
  nand ginst18746 (P2_U5947, P2_R1297_U6, P2_U3070);
  nand ginst18747 (P2_U5948, P2_U3070, P2_U3867);
  nand ginst18748 (P2_U5949, P2_R1297_U6, P2_U3066);
  nand ginst18749 (P2_U5950, P2_U3066, P2_U3867);
  nand ginst18750 (P2_U5951, P2_R1297_U6, P2_U3059);
  nand ginst18751 (P2_U5952, P2_U3059, P2_U3867);
  nand ginst18752 (P2_U5953, P2_R1297_U6, P2_R1300_U8);
  nand ginst18753 (P2_U5954, P2_U3055, P2_U3867);
  nand ginst18754 (P2_U5955, P2_R1297_U6, P2_R1300_U6);
  nand ginst18755 (P2_U5956, P2_U3058, P2_U3867);
  nand ginst18756 (P2_U5957, P2_R1297_U6, P2_U3063);
  nand ginst18757 (P2_U5958, P2_U3063, P2_U3867);
  nand ginst18758 (P2_U5959, P2_R1297_U6, P2_U3054);
  nand ginst18759 (P2_U5960, P2_U3054, P2_U3867);
  nand ginst18760 (P2_U5961, P2_R1297_U6, P2_U3053);
  nand ginst18761 (P2_U5962, P2_U3053, P2_U3867);
  nand ginst18762 (P2_U5963, P2_R1297_U6, P2_U3052);
  nand ginst18763 (P2_U5964, P2_U3052, P2_U3867);
  nand ginst18764 (P2_U5965, P2_R1297_U6, P2_U3056);
  nand ginst18765 (P2_U5966, P2_U3056, P2_U3867);
  nand ginst18766 (P2_U5967, P2_R1297_U6, P2_U3057);
  nand ginst18767 (P2_U5968, P2_U3057, P2_U3867);
  nand ginst18768 (P2_U5969, P2_R1297_U6, P2_U3064);
  nand ginst18769 (P2_U5970, P2_U3064, P2_U3867);
  nand ginst18770 (P2_U5971, P2_R1297_U6, P2_U3065);
  nand ginst18771 (P2_U5972, P2_U3065, P2_U3867);
  nand ginst18772 (P2_U5973, P2_R1297_U6, P2_U3060);
  nand ginst18773 (P2_U5974, P2_U3060, P2_U3867);
  nand ginst18774 (P2_U5975, P2_R1297_U6, P2_U3074);
  nand ginst18775 (P2_U5976, P2_U3074, P2_U3867);
  nand ginst18776 (P2_U5977, P2_R1297_U6, P2_U3075);
  nand ginst18777 (P2_U5978, P2_U3075, P2_U3867);
  nand ginst18778 (P2_U5979, P2_R1297_U6, P2_U3067);
  nand ginst18779 (P2_U5980, P2_U3067, P2_U3867);
  nand ginst18780 (P2_U5981, P2_R1297_U6, P2_U3080);
  nand ginst18781 (P2_U5982, P2_U3080, P2_U3867);
  nand ginst18782 (P2_U5983, P2_R1297_U6, P2_U3081);
  nand ginst18783 (P2_U5984, P2_U3081, P2_U3867);
  nand ginst18784 (P2_U5985, P2_R1297_U6, P2_U3068);
  nand ginst18785 (P2_U5986, P2_U3068, P2_U3867);
  nand ginst18786 (P2_U5987, P2_R1297_U6, P2_U3072);
  nand ginst18787 (P2_U5988, P2_U3072, P2_U3867);
  nand ginst18788 (P2_U5989, P2_R1297_U6, P2_U3073);
  nand ginst18789 (P2_U5990, P2_U3073, P2_U3867);
  nand ginst18790 (P2_U5991, P2_R1297_U6, P2_U3078);
  nand ginst18791 (P2_U5992, P2_U3078, P2_U3867);
  nand ginst18792 (P2_U5993, P2_R1297_U6, P2_U3079);
  nand ginst18793 (P2_U5994, P2_U3079, P2_U3867);
  nand ginst18794 (P2_U5995, P2_R1297_U6, P2_U3071);
  nand ginst18795 (P2_U5996, P2_U3071, P2_U3867);
  nand ginst18796 (P2_U5997, P2_R1297_U6, P2_U3062);
  nand ginst18797 (P2_U5998, P2_U3062, P2_U3867);
  nand ginst18798 (P2_U5999, P2_R1297_U6, P2_U3061);
  nand ginst18799 (P2_U6000, P2_U3061, P2_U3867);
  nand ginst18800 (P2_U6001, P2_R1297_U6, P2_U3077);
  nand ginst18801 (P2_U6002, P2_U3077, P2_U3867);
  nand ginst18802 (P2_U6003, P2_R1297_U6, P2_U3076);
  nand ginst18803 (P2_U6004, P2_U3076, P2_U3867);
  nand ginst18804 (P2_U6005, P2_REG1_REG_9__SCAN_IN, P2_U5464);
  nand ginst18805 (P2_U6006, P2_REG2_REG_9__SCAN_IN, P2_U3384);
  nand ginst18806 (P2_U6007, P2_REG1_REG_8__SCAN_IN, P2_U5464);
  nand ginst18807 (P2_U6008, P2_REG2_REG_8__SCAN_IN, P2_U3384);
  nand ginst18808 (P2_U6009, P2_REG1_REG_7__SCAN_IN, P2_U5464);
  nand ginst18809 (P2_U6010, P2_REG2_REG_7__SCAN_IN, P2_U3384);
  nand ginst18810 (P2_U6011, P2_REG1_REG_6__SCAN_IN, P2_U5464);
  nand ginst18811 (P2_U6012, P2_REG2_REG_6__SCAN_IN, P2_U3384);
  nand ginst18812 (P2_U6013, P2_REG1_REG_5__SCAN_IN, P2_U5464);
  nand ginst18813 (P2_U6014, P2_REG2_REG_5__SCAN_IN, P2_U3384);
  nand ginst18814 (P2_U6015, P2_REG1_REG_4__SCAN_IN, P2_U5464);
  nand ginst18815 (P2_U6016, P2_REG2_REG_4__SCAN_IN, P2_U3384);
  nand ginst18816 (P2_U6017, P2_REG1_REG_3__SCAN_IN, P2_U5464);
  nand ginst18817 (P2_U6018, P2_REG2_REG_3__SCAN_IN, P2_U3384);
  nand ginst18818 (P2_U6019, P2_REG1_REG_2__SCAN_IN, P2_U5464);
  nand ginst18819 (P2_U6020, P2_REG2_REG_2__SCAN_IN, P2_U3384);
  nand ginst18820 (P2_U6021, P2_REG1_REG_19__SCAN_IN, P2_U5464);
  nand ginst18821 (P2_U6022, P2_REG2_REG_19__SCAN_IN, P2_U3384);
  nand ginst18822 (P2_U6023, P2_REG1_REG_18__SCAN_IN, P2_U5464);
  nand ginst18823 (P2_U6024, P2_REG2_REG_18__SCAN_IN, P2_U3384);
  nand ginst18824 (P2_U6025, P2_REG1_REG_17__SCAN_IN, P2_U5464);
  nand ginst18825 (P2_U6026, P2_REG2_REG_17__SCAN_IN, P2_U3384);
  nand ginst18826 (P2_U6027, P2_REG1_REG_16__SCAN_IN, P2_U5464);
  nand ginst18827 (P2_U6028, P2_REG2_REG_16__SCAN_IN, P2_U3384);
  nand ginst18828 (P2_U6029, P2_REG1_REG_15__SCAN_IN, P2_U5464);
  nand ginst18829 (P2_U6030, P2_REG2_REG_15__SCAN_IN, P2_U3384);
  nand ginst18830 (P2_U6031, P2_REG1_REG_14__SCAN_IN, P2_U5464);
  nand ginst18831 (P2_U6032, P2_REG2_REG_14__SCAN_IN, P2_U3384);
  nand ginst18832 (P2_U6033, P2_REG1_REG_13__SCAN_IN, P2_U5464);
  nand ginst18833 (P2_U6034, P2_REG2_REG_13__SCAN_IN, P2_U3384);
  nand ginst18834 (P2_U6035, P2_REG1_REG_12__SCAN_IN, P2_U5464);
  nand ginst18835 (P2_U6036, P2_REG2_REG_12__SCAN_IN, P2_U3384);
  nand ginst18836 (P2_U6037, P2_REG1_REG_11__SCAN_IN, P2_U5464);
  nand ginst18837 (P2_U6038, P2_REG2_REG_11__SCAN_IN, P2_U3384);
  nand ginst18838 (P2_U6039, P2_REG1_REG_10__SCAN_IN, P2_U5464);
  nand ginst18839 (P2_U6040, P2_REG2_REG_10__SCAN_IN, P2_U3384);
  nand ginst18840 (P2_U6041, P2_REG1_REG_1__SCAN_IN, P2_U5464);
  nand ginst18841 (P2_U6042, P2_REG2_REG_1__SCAN_IN, P2_U3384);
  nand ginst18842 (P2_U6043, P2_REG1_REG_0__SCAN_IN, P2_U5464);
  nand ginst18843 (P2_U6044, P2_REG2_REG_0__SCAN_IN, P2_U3384);
  nand ginst18844 (R140_U10, R140_U324, R140_U468, R140_U469);
  nand ginst18845 (R140_U100, R140_U449, R140_U450);
  nand ginst18846 (R140_U101, R140_U456, R140_U457);
  nand ginst18847 (R140_U102, R140_U463, R140_U464);
  nand ginst18848 (R140_U103, R140_U475, R140_U476);
  nand ginst18849 (R140_U104, R140_U482, R140_U483);
  nand ginst18850 (R140_U105, R140_U489, R140_U490);
  nand ginst18851 (R140_U106, R140_U496, R140_U497);
  nand ginst18852 (R140_U107, R140_U503, R140_U504);
  nand ginst18853 (R140_U108, R140_U510, R140_U511);
  nand ginst18854 (R140_U109, R140_U517, R140_U518);
  and ginst18855 (R140_U11, R140_U124, R140_U323);
  nand ginst18856 (R140_U110, R140_U524, R140_U525);
  nand ginst18857 (R140_U111, R140_U531, R140_U532);
  nand ginst18858 (R140_U112, R140_U538, R140_U539);
  and ginst18859 (R140_U113, R140_U189, R140_U193);
  and ginst18860 (R140_U114, R140_U194, R140_U287);
  and ginst18861 (R140_U115, R140_U199, R140_U4);
  and ginst18862 (R140_U116, R140_U200, R140_U290);
  and ginst18863 (R140_U117, R140_U204, R140_U291);
  and ginst18864 (R140_U118, R140_U207, R140_U6);
  and ginst18865 (R140_U119, R140_U208, R140_U295);
  not ginst18866 (R140_U12, SI_8_);
  and ginst18867 (R140_U120, R140_U219, R140_U8);
  and ginst18868 (R140_U121, R140_U220, R140_U303);
  and ginst18869 (R140_U122, R140_U280, R140_U282, R140_U9);
  and ginst18870 (R140_U123, R140_U283, R140_U376);
  and ginst18871 (R140_U124, R140_U141, R140_U284);
  and ginst18872 (R140_U125, R140_U325, R140_U326);
  nand ginst18873 (R140_U126, R140_U117, R140_U309);
  and ginst18874 (R140_U127, R140_U332, R140_U333);
  nand ginst18875 (R140_U128, R140_U16, R140_U307);
  and ginst18876 (R140_U129, R140_U339, R140_U340);
  not ginst18877 (R140_U13, U90);
  nand ginst18878 (R140_U130, R140_U116, R140_U319);
  and ginst18879 (R140_U131, R140_U346, R140_U347);
  nand ginst18880 (R140_U132, R140_U289, R140_U317);
  and ginst18881 (R140_U133, R140_U353, R140_U354);
  nand ginst18882 (R140_U134, R140_U23, R140_U315);
  and ginst18883 (R140_U135, R140_U360, R140_U361);
  nand ginst18884 (R140_U136, R140_U114, R140_U321);
  and ginst18885 (R140_U137, R140_U367, R140_U368);
  nand ginst18886 (R140_U138, R140_U190, R140_U28);
  not ginst18887 (R140_U139, U95);
  not ginst18888 (R140_U14, SI_7_);
  not ginst18889 (R140_U140, SI_31_);
  and ginst18890 (R140_U141, R140_U379, R140_U380);
  and ginst18891 (R140_U142, R140_U381, R140_U382);
  nand ginst18892 (R140_U143, R140_U279, R140_U280);
  nand ginst18893 (R140_U144, R140_U285, R140_U286, R140_U79);
  and ginst18894 (R140_U145, R140_U395, R140_U396);
  nand ginst18895 (R140_U146, R140_U275, R140_U276);
  and ginst18896 (R140_U147, R140_U402, R140_U403);
  nand ginst18897 (R140_U148, R140_U271, R140_U272);
  and ginst18898 (R140_U149, R140_U409, R140_U410);
  not ginst18899 (R140_U15, U91);
  nand ginst18900 (R140_U150, R140_U267, R140_U268);
  and ginst18901 (R140_U151, R140_U416, R140_U417);
  nand ginst18902 (R140_U152, R140_U263, R140_U264);
  and ginst18903 (R140_U153, R140_U423, R140_U424);
  nand ginst18904 (R140_U154, R140_U259, R140_U260);
  and ginst18905 (R140_U155, R140_U430, R140_U431);
  nand ginst18906 (R140_U156, R140_U255, R140_U256);
  and ginst18907 (R140_U157, R140_U437, R140_U438);
  nand ginst18908 (R140_U158, R140_U251, R140_U252);
  and ginst18909 (R140_U159, R140_U444, R140_U445);
  nand ginst18910 (R140_U16, SI_7_, U91);
  nand ginst18911 (R140_U160, R140_U247, R140_U248);
  and ginst18912 (R140_U161, R140_U451, R140_U452);
  nand ginst18913 (R140_U162, R140_U243, R140_U244);
  and ginst18914 (R140_U163, R140_U458, R140_U459);
  nand ginst18915 (R140_U164, R140_U239, R140_U240);
  nand ginst18916 (R140_U165, SI_0_, U120);
  and ginst18917 (R140_U166, R140_U470, R140_U471);
  nand ginst18918 (R140_U167, R140_U235, R140_U236);
  and ginst18919 (R140_U168, R140_U477, R140_U478);
  nand ginst18920 (R140_U169, R140_U231, R140_U232);
  not ginst18921 (R140_U17, SI_6_);
  and ginst18922 (R140_U170, R140_U484, R140_U485);
  nand ginst18923 (R140_U171, R140_U227, R140_U228);
  and ginst18924 (R140_U172, R140_U491, R140_U492);
  nand ginst18925 (R140_U173, R140_U223, R140_U224);
  and ginst18926 (R140_U174, R140_U498, R140_U499);
  nand ginst18927 (R140_U175, R140_U121, R140_U302);
  and ginst18928 (R140_U176, R140_U505, R140_U506);
  nand ginst18929 (R140_U177, R140_U299, R140_U301);
  and ginst18930 (R140_U178, R140_U512, R140_U513);
  nand ginst18931 (R140_U179, R140_U296, R140_U298);
  not ginst18932 (R140_U18, U92);
  and ginst18933 (R140_U180, R140_U519, R140_U520);
  nand ginst18934 (R140_U181, R140_U210, R140_U46);
  and ginst18935 (R140_U182, R140_U526, R140_U527);
  nand ginst18936 (R140_U183, R140_U119, R140_U313);
  and ginst18937 (R140_U184, R140_U533, R140_U534);
  nand ginst18938 (R140_U185, R140_U294, R140_U311);
  not ginst18939 (R140_U186, R140_U79);
  not ginst18940 (R140_U187, R140_U165);
  not ginst18941 (R140_U188, R140_U144);
  or ginst18942 (R140_U189, SI_2_, U108);
  not ginst18943 (R140_U19, SI_5_);
  nand ginst18944 (R140_U190, R140_U189, R140_U304);
  not ginst18945 (R140_U191, R140_U28);
  not ginst18946 (R140_U192, R140_U138);
  or ginst18947 (R140_U193, SI_3_, U97);
  nand ginst18948 (R140_U194, SI_3_, U97);
  or ginst18949 (R140_U195, SI_4_, U94);
  not ginst18950 (R140_U196, R140_U23);
  or ginst18951 (R140_U197, SI_5_, U93);
  nand ginst18952 (R140_U198, SI_5_, U93);
  or ginst18953 (R140_U199, SI_6_, U92);
  not ginst18954 (R140_U20, U93);
  nand ginst18955 (R140_U200, SI_6_, U92);
  or ginst18956 (R140_U201, SI_7_, U91);
  not ginst18957 (R140_U202, R140_U16);
  or ginst18958 (R140_U203, SI_8_, U90);
  nand ginst18959 (R140_U204, SI_8_, U90);
  or ginst18960 (R140_U205, SI_9_, U89);
  nand ginst18961 (R140_U206, SI_9_, U89);
  or ginst18962 (R140_U207, SI_10_, U118);
  nand ginst18963 (R140_U208, SI_10_, U118);
  or ginst18964 (R140_U209, SI_11_, U117);
  not ginst18965 (R140_U21, SI_4_);
  nand ginst18966 (R140_U210, R140_U183, R140_U209);
  not ginst18967 (R140_U211, R140_U46);
  not ginst18968 (R140_U212, R140_U181);
  or ginst18969 (R140_U213, SI_12_, U116);
  nand ginst18970 (R140_U214, SI_12_, U116);
  not ginst18971 (R140_U215, R140_U179);
  or ginst18972 (R140_U216, SI_13_, U115);
  nand ginst18973 (R140_U217, SI_13_, U115);
  not ginst18974 (R140_U218, R140_U177);
  or ginst18975 (R140_U219, SI_14_, U114);
  not ginst18976 (R140_U22, U94);
  nand ginst18977 (R140_U220, SI_14_, U114);
  not ginst18978 (R140_U221, R140_U175);
  or ginst18979 (R140_U222, SI_15_, U113);
  nand ginst18980 (R140_U223, R140_U175, R140_U222);
  nand ginst18981 (R140_U224, SI_15_, U113);
  not ginst18982 (R140_U225, R140_U173);
  or ginst18983 (R140_U226, SI_16_, U112);
  nand ginst18984 (R140_U227, R140_U173, R140_U226);
  nand ginst18985 (R140_U228, SI_16_, U112);
  not ginst18986 (R140_U229, R140_U171);
  nand ginst18987 (R140_U23, SI_4_, U94);
  or ginst18988 (R140_U230, SI_17_, U111);
  nand ginst18989 (R140_U231, R140_U171, R140_U230);
  nand ginst18990 (R140_U232, SI_17_, U111);
  not ginst18991 (R140_U233, R140_U169);
  or ginst18992 (R140_U234, SI_18_, U110);
  nand ginst18993 (R140_U235, R140_U169, R140_U234);
  nand ginst18994 (R140_U236, SI_18_, U110);
  not ginst18995 (R140_U237, R140_U167);
  or ginst18996 (R140_U238, SI_19_, U109);
  nand ginst18997 (R140_U239, R140_U167, R140_U238);
  not ginst18998 (R140_U24, SI_3_);
  nand ginst18999 (R140_U240, SI_19_, U109);
  not ginst19000 (R140_U241, R140_U164);
  or ginst19001 (R140_U242, SI_20_, U107);
  nand ginst19002 (R140_U243, R140_U164, R140_U242);
  nand ginst19003 (R140_U244, SI_20_, U107);
  not ginst19004 (R140_U245, R140_U162);
  or ginst19005 (R140_U246, SI_21_, U106);
  nand ginst19006 (R140_U247, R140_U162, R140_U246);
  nand ginst19007 (R140_U248, SI_21_, U106);
  not ginst19008 (R140_U249, R140_U160);
  not ginst19009 (R140_U25, U97);
  or ginst19010 (R140_U250, SI_22_, U105);
  nand ginst19011 (R140_U251, R140_U160, R140_U250);
  nand ginst19012 (R140_U252, SI_22_, U105);
  not ginst19013 (R140_U253, R140_U158);
  or ginst19014 (R140_U254, SI_23_, U104);
  nand ginst19015 (R140_U255, R140_U158, R140_U254);
  nand ginst19016 (R140_U256, SI_23_, U104);
  not ginst19017 (R140_U257, R140_U156);
  or ginst19018 (R140_U258, SI_24_, U103);
  nand ginst19019 (R140_U259, R140_U156, R140_U258);
  not ginst19020 (R140_U26, SI_2_);
  nand ginst19021 (R140_U260, SI_24_, U103);
  not ginst19022 (R140_U261, R140_U154);
  or ginst19023 (R140_U262, SI_25_, U102);
  nand ginst19024 (R140_U263, R140_U154, R140_U262);
  nand ginst19025 (R140_U264, SI_25_, U102);
  not ginst19026 (R140_U265, R140_U152);
  or ginst19027 (R140_U266, SI_26_, U101);
  nand ginst19028 (R140_U267, R140_U152, R140_U266);
  nand ginst19029 (R140_U268, SI_26_, U101);
  not ginst19030 (R140_U269, R140_U150);
  not ginst19031 (R140_U27, U108);
  or ginst19032 (R140_U270, SI_27_, U100);
  nand ginst19033 (R140_U271, R140_U150, R140_U270);
  nand ginst19034 (R140_U272, SI_27_, U100);
  not ginst19035 (R140_U273, R140_U148);
  or ginst19036 (R140_U274, SI_28_, U99);
  nand ginst19037 (R140_U275, R140_U148, R140_U274);
  nand ginst19038 (R140_U276, SI_28_, U99);
  not ginst19039 (R140_U277, R140_U146);
  or ginst19040 (R140_U278, SI_29_, U98);
  nand ginst19041 (R140_U279, R140_U146, R140_U278);
  nand ginst19042 (R140_U28, SI_2_, U108);
  nand ginst19043 (R140_U280, SI_29_, U98);
  not ginst19044 (R140_U281, R140_U143);
  nand ginst19045 (R140_U282, SI_30_, U96);
  or ginst19046 (R140_U283, SI_30_, U96);
  nand ginst19047 (R140_U284, R140_U122, R140_U279);
  nand ginst19048 (R140_U285, SI_0_, U119, U120);
  nand ginst19049 (R140_U286, SI_1_, U119);
  nand ginst19050 (R140_U287, R140_U191, R140_U193);
  nand ginst19051 (R140_U288, R140_U196, R140_U197);
  not ginst19052 (R140_U289, R140_U35);
  not ginst19053 (R140_U29, SI_1_);
  nand ginst19054 (R140_U290, R140_U199, R140_U35);
  nand ginst19055 (R140_U291, R140_U202, R140_U203);
  nand ginst19056 (R140_U292, R140_U204, R140_U291);
  nand ginst19057 (R140_U293, R140_U205, R140_U292);
  not ginst19058 (R140_U294, R140_U82);
  nand ginst19059 (R140_U295, R140_U207, R140_U82);
  nand ginst19060 (R140_U296, R140_U183, R140_U7);
  nand ginst19061 (R140_U297, R140_U211, R140_U213);
  not ginst19062 (R140_U298, R140_U81);
  nand ginst19063 (R140_U299, R140_U183, R140_U8);
  not ginst19064 (R140_U30, SI_0_);
  nand ginst19065 (R140_U300, R140_U216, R140_U81);
  not ginst19066 (R140_U301, R140_U80);
  nand ginst19067 (R140_U302, R140_U120, R140_U183);
  nand ginst19068 (R140_U303, R140_U219, R140_U80);
  nand ginst19069 (R140_U304, R140_U286, R140_U305, R140_U306);
  nand ginst19070 (R140_U305, SI_0_, U119, U120);
  nand ginst19071 (R140_U306, SI_1_, SI_0_, U120);
  nand ginst19072 (R140_U307, R140_U130, R140_U201);
  not ginst19073 (R140_U308, R140_U128);
  nand ginst19074 (R140_U309, R140_U130, R140_U5);
  not ginst19075 (R140_U31, U120);
  not ginst19076 (R140_U310, R140_U126);
  nand ginst19077 (R140_U311, R140_U130, R140_U6);
  not ginst19078 (R140_U312, R140_U185);
  nand ginst19079 (R140_U313, R140_U118, R140_U130);
  not ginst19080 (R140_U314, R140_U183);
  nand ginst19081 (R140_U315, R140_U136, R140_U195);
  not ginst19082 (R140_U316, R140_U134);
  nand ginst19083 (R140_U317, R140_U136, R140_U4);
  not ginst19084 (R140_U318, R140_U132);
  nand ginst19085 (R140_U319, R140_U115, R140_U136);
  not ginst19086 (R140_U32, U119);
  not ginst19087 (R140_U320, R140_U130);
  nand ginst19088 (R140_U321, R140_U113, R140_U144);
  not ginst19089 (R140_U322, R140_U136);
  nand ginst19090 (R140_U323, R140_U123, R140_U143);
  nand ginst19091 (R140_U324, R140_U186, U119);
  nand ginst19092 (R140_U325, R140_U34, U89);
  nand ginst19093 (R140_U326, SI_9_, R140_U33);
  nand ginst19094 (R140_U327, R140_U34, U89);
  nand ginst19095 (R140_U328, SI_9_, R140_U33);
  nand ginst19096 (R140_U329, R140_U327, R140_U328);
  not ginst19097 (R140_U33, U89);
  nand ginst19098 (R140_U330, R140_U125, R140_U126);
  nand ginst19099 (R140_U331, R140_U310, R140_U329);
  nand ginst19100 (R140_U332, R140_U12, U90);
  nand ginst19101 (R140_U333, SI_8_, R140_U13);
  nand ginst19102 (R140_U334, R140_U12, U90);
  nand ginst19103 (R140_U335, SI_8_, R140_U13);
  nand ginst19104 (R140_U336, R140_U334, R140_U335);
  nand ginst19105 (R140_U337, R140_U127, R140_U128);
  nand ginst19106 (R140_U338, R140_U308, R140_U336);
  nand ginst19107 (R140_U339, R140_U14, U91);
  not ginst19108 (R140_U34, SI_9_);
  nand ginst19109 (R140_U340, SI_7_, R140_U15);
  nand ginst19110 (R140_U341, R140_U14, U91);
  nand ginst19111 (R140_U342, SI_7_, R140_U15);
  nand ginst19112 (R140_U343, R140_U341, R140_U342);
  nand ginst19113 (R140_U344, R140_U129, R140_U130);
  nand ginst19114 (R140_U345, R140_U320, R140_U343);
  nand ginst19115 (R140_U346, R140_U17, U92);
  nand ginst19116 (R140_U347, SI_6_, R140_U18);
  nand ginst19117 (R140_U348, R140_U17, U92);
  nand ginst19118 (R140_U349, SI_6_, R140_U18);
  nand ginst19119 (R140_U35, R140_U198, R140_U288);
  nand ginst19120 (R140_U350, R140_U348, R140_U349);
  nand ginst19121 (R140_U351, R140_U131, R140_U132);
  nand ginst19122 (R140_U352, R140_U318, R140_U350);
  nand ginst19123 (R140_U353, R140_U19, U93);
  nand ginst19124 (R140_U354, SI_5_, R140_U20);
  nand ginst19125 (R140_U355, R140_U19, U93);
  nand ginst19126 (R140_U356, SI_5_, R140_U20);
  nand ginst19127 (R140_U357, R140_U355, R140_U356);
  nand ginst19128 (R140_U358, R140_U133, R140_U134);
  nand ginst19129 (R140_U359, R140_U316, R140_U357);
  not ginst19130 (R140_U36, SI_14_);
  nand ginst19131 (R140_U360, R140_U21, U94);
  nand ginst19132 (R140_U361, SI_4_, R140_U22);
  nand ginst19133 (R140_U362, R140_U21, U94);
  nand ginst19134 (R140_U363, SI_4_, R140_U22);
  nand ginst19135 (R140_U364, R140_U362, R140_U363);
  nand ginst19136 (R140_U365, R140_U135, R140_U136);
  nand ginst19137 (R140_U366, R140_U322, R140_U364);
  nand ginst19138 (R140_U367, R140_U24, U97);
  nand ginst19139 (R140_U368, SI_3_, R140_U25);
  nand ginst19140 (R140_U369, R140_U24, U97);
  not ginst19141 (R140_U37, U114);
  nand ginst19142 (R140_U370, SI_3_, R140_U25);
  nand ginst19143 (R140_U371, R140_U369, R140_U370);
  nand ginst19144 (R140_U372, R140_U137, R140_U138);
  nand ginst19145 (R140_U373, R140_U192, R140_U371);
  nand ginst19146 (R140_U374, R140_U140, U95);
  nand ginst19147 (R140_U375, SI_31_, R140_U139);
  nand ginst19148 (R140_U376, R140_U374, R140_U375);
  nand ginst19149 (R140_U377, R140_U140, U95);
  nand ginst19150 (R140_U378, SI_31_, R140_U139);
  nand ginst19151 (R140_U379, R140_U77, R140_U78, R140_U9);
  not ginst19152 (R140_U38, SI_10_);
  nand ginst19153 (R140_U380, SI_30_, R140_U376, U96);
  nand ginst19154 (R140_U381, R140_U77, U96);
  nand ginst19155 (R140_U382, SI_30_, R140_U78);
  nand ginst19156 (R140_U383, R140_U77, U96);
  nand ginst19157 (R140_U384, SI_30_, R140_U78);
  nand ginst19158 (R140_U385, R140_U383, R140_U384);
  nand ginst19159 (R140_U386, R140_U142, R140_U143);
  nand ginst19160 (R140_U387, R140_U281, R140_U385);
  nand ginst19161 (R140_U388, R140_U26, U108);
  nand ginst19162 (R140_U389, SI_2_, R140_U27);
  not ginst19163 (R140_U39, U118);
  nand ginst19164 (R140_U390, R140_U26, U108);
  nand ginst19165 (R140_U391, SI_2_, R140_U27);
  nand ginst19166 (R140_U392, R140_U390, R140_U391);
  nand ginst19167 (R140_U393, R140_U144, R140_U388, R140_U389);
  nand ginst19168 (R140_U394, R140_U188, R140_U392);
  nand ginst19169 (R140_U395, R140_U75, U98);
  nand ginst19170 (R140_U396, SI_29_, R140_U76);
  nand ginst19171 (R140_U397, R140_U75, U98);
  nand ginst19172 (R140_U398, SI_29_, R140_U76);
  nand ginst19173 (R140_U399, R140_U397, R140_U398);
  and ginst19174 (R140_U4, R140_U195, R140_U197);
  not ginst19175 (R140_U40, SI_13_);
  nand ginst19176 (R140_U400, R140_U145, R140_U146);
  nand ginst19177 (R140_U401, R140_U277, R140_U399);
  nand ginst19178 (R140_U402, R140_U73, U99);
  nand ginst19179 (R140_U403, SI_28_, R140_U74);
  nand ginst19180 (R140_U404, R140_U73, U99);
  nand ginst19181 (R140_U405, SI_28_, R140_U74);
  nand ginst19182 (R140_U406, R140_U404, R140_U405);
  nand ginst19183 (R140_U407, R140_U147, R140_U148);
  nand ginst19184 (R140_U408, R140_U273, R140_U406);
  nand ginst19185 (R140_U409, R140_U71, U100);
  not ginst19186 (R140_U41, U115);
  nand ginst19187 (R140_U410, SI_27_, R140_U72);
  nand ginst19188 (R140_U411, R140_U71, U100);
  nand ginst19189 (R140_U412, SI_27_, R140_U72);
  nand ginst19190 (R140_U413, R140_U411, R140_U412);
  nand ginst19191 (R140_U414, R140_U149, R140_U150);
  nand ginst19192 (R140_U415, R140_U269, R140_U413);
  nand ginst19193 (R140_U416, R140_U69, U101);
  nand ginst19194 (R140_U417, SI_26_, R140_U70);
  nand ginst19195 (R140_U418, R140_U69, U101);
  nand ginst19196 (R140_U419, SI_26_, R140_U70);
  not ginst19197 (R140_U42, SI_12_);
  nand ginst19198 (R140_U420, R140_U418, R140_U419);
  nand ginst19199 (R140_U421, R140_U151, R140_U152);
  nand ginst19200 (R140_U422, R140_U265, R140_U420);
  nand ginst19201 (R140_U423, R140_U67, U102);
  nand ginst19202 (R140_U424, SI_25_, R140_U68);
  nand ginst19203 (R140_U425, R140_U67, U102);
  nand ginst19204 (R140_U426, SI_25_, R140_U68);
  nand ginst19205 (R140_U427, R140_U425, R140_U426);
  nand ginst19206 (R140_U428, R140_U153, R140_U154);
  nand ginst19207 (R140_U429, R140_U261, R140_U427);
  not ginst19208 (R140_U43, U116);
  nand ginst19209 (R140_U430, R140_U65, U103);
  nand ginst19210 (R140_U431, SI_24_, R140_U66);
  nand ginst19211 (R140_U432, R140_U65, U103);
  nand ginst19212 (R140_U433, SI_24_, R140_U66);
  nand ginst19213 (R140_U434, R140_U432, R140_U433);
  nand ginst19214 (R140_U435, R140_U155, R140_U156);
  nand ginst19215 (R140_U436, R140_U257, R140_U434);
  nand ginst19216 (R140_U437, R140_U63, U104);
  nand ginst19217 (R140_U438, SI_23_, R140_U64);
  nand ginst19218 (R140_U439, R140_U63, U104);
  not ginst19219 (R140_U44, SI_11_);
  nand ginst19220 (R140_U440, SI_23_, R140_U64);
  nand ginst19221 (R140_U441, R140_U439, R140_U440);
  nand ginst19222 (R140_U442, R140_U157, R140_U158);
  nand ginst19223 (R140_U443, R140_U253, R140_U441);
  nand ginst19224 (R140_U444, R140_U61, U105);
  nand ginst19225 (R140_U445, SI_22_, R140_U62);
  nand ginst19226 (R140_U446, R140_U61, U105);
  nand ginst19227 (R140_U447, SI_22_, R140_U62);
  nand ginst19228 (R140_U448, R140_U446, R140_U447);
  nand ginst19229 (R140_U449, R140_U159, R140_U160);
  not ginst19230 (R140_U45, U117);
  nand ginst19231 (R140_U450, R140_U249, R140_U448);
  nand ginst19232 (R140_U451, R140_U59, U106);
  nand ginst19233 (R140_U452, SI_21_, R140_U60);
  nand ginst19234 (R140_U453, R140_U59, U106);
  nand ginst19235 (R140_U454, SI_21_, R140_U60);
  nand ginst19236 (R140_U455, R140_U453, R140_U454);
  nand ginst19237 (R140_U456, R140_U161, R140_U162);
  nand ginst19238 (R140_U457, R140_U245, R140_U455);
  nand ginst19239 (R140_U458, R140_U57, U107);
  nand ginst19240 (R140_U459, SI_20_, R140_U58);
  nand ginst19241 (R140_U46, SI_11_, U117);
  nand ginst19242 (R140_U460, R140_U57, U107);
  nand ginst19243 (R140_U461, SI_20_, R140_U58);
  nand ginst19244 (R140_U462, R140_U460, R140_U461);
  nand ginst19245 (R140_U463, R140_U163, R140_U164);
  nand ginst19246 (R140_U464, R140_U241, R140_U462);
  nand ginst19247 (R140_U465, R140_U165, U119);
  nand ginst19248 (R140_U466, R140_U187, R140_U32);
  nand ginst19249 (R140_U467, R140_U465, R140_U466);
  nand ginst19250 (R140_U468, SI_1_, R140_U165, R140_U32);
  nand ginst19251 (R140_U469, R140_U29, R140_U467);
  not ginst19252 (R140_U47, SI_15_);
  nand ginst19253 (R140_U470, R140_U55, U109);
  nand ginst19254 (R140_U471, SI_19_, R140_U56);
  nand ginst19255 (R140_U472, R140_U55, U109);
  nand ginst19256 (R140_U473, SI_19_, R140_U56);
  nand ginst19257 (R140_U474, R140_U472, R140_U473);
  nand ginst19258 (R140_U475, R140_U166, R140_U167);
  nand ginst19259 (R140_U476, R140_U237, R140_U474);
  nand ginst19260 (R140_U477, R140_U53, U110);
  nand ginst19261 (R140_U478, SI_18_, R140_U54);
  nand ginst19262 (R140_U479, R140_U53, U110);
  not ginst19263 (R140_U48, U113);
  nand ginst19264 (R140_U480, SI_18_, R140_U54);
  nand ginst19265 (R140_U481, R140_U479, R140_U480);
  nand ginst19266 (R140_U482, R140_U168, R140_U169);
  nand ginst19267 (R140_U483, R140_U233, R140_U481);
  nand ginst19268 (R140_U484, R140_U51, U111);
  nand ginst19269 (R140_U485, SI_17_, R140_U52);
  nand ginst19270 (R140_U486, R140_U51, U111);
  nand ginst19271 (R140_U487, SI_17_, R140_U52);
  nand ginst19272 (R140_U488, R140_U486, R140_U487);
  nand ginst19273 (R140_U489, R140_U170, R140_U171);
  not ginst19274 (R140_U49, SI_16_);
  nand ginst19275 (R140_U490, R140_U229, R140_U488);
  nand ginst19276 (R140_U491, R140_U49, U112);
  nand ginst19277 (R140_U492, SI_16_, R140_U50);
  nand ginst19278 (R140_U493, R140_U49, U112);
  nand ginst19279 (R140_U494, SI_16_, R140_U50);
  nand ginst19280 (R140_U495, R140_U493, R140_U494);
  nand ginst19281 (R140_U496, R140_U172, R140_U173);
  nand ginst19282 (R140_U497, R140_U225, R140_U495);
  nand ginst19283 (R140_U498, R140_U47, U113);
  nand ginst19284 (R140_U499, SI_15_, R140_U48);
  and ginst19285 (R140_U5, R140_U201, R140_U203);
  not ginst19286 (R140_U50, U112);
  nand ginst19287 (R140_U500, R140_U47, U113);
  nand ginst19288 (R140_U501, SI_15_, R140_U48);
  nand ginst19289 (R140_U502, R140_U500, R140_U501);
  nand ginst19290 (R140_U503, R140_U174, R140_U175);
  nand ginst19291 (R140_U504, R140_U221, R140_U502);
  nand ginst19292 (R140_U505, R140_U36, U114);
  nand ginst19293 (R140_U506, SI_14_, R140_U37);
  nand ginst19294 (R140_U507, R140_U36, U114);
  nand ginst19295 (R140_U508, SI_14_, R140_U37);
  nand ginst19296 (R140_U509, R140_U507, R140_U508);
  not ginst19297 (R140_U51, SI_17_);
  nand ginst19298 (R140_U510, R140_U176, R140_U177);
  nand ginst19299 (R140_U511, R140_U218, R140_U509);
  nand ginst19300 (R140_U512, R140_U40, U115);
  nand ginst19301 (R140_U513, SI_13_, R140_U41);
  nand ginst19302 (R140_U514, R140_U40, U115);
  nand ginst19303 (R140_U515, SI_13_, R140_U41);
  nand ginst19304 (R140_U516, R140_U514, R140_U515);
  nand ginst19305 (R140_U517, R140_U178, R140_U179);
  nand ginst19306 (R140_U518, R140_U215, R140_U516);
  nand ginst19307 (R140_U519, R140_U42, U116);
  not ginst19308 (R140_U52, U111);
  nand ginst19309 (R140_U520, SI_12_, R140_U43);
  nand ginst19310 (R140_U521, R140_U42, U116);
  nand ginst19311 (R140_U522, SI_12_, R140_U43);
  nand ginst19312 (R140_U523, R140_U521, R140_U522);
  nand ginst19313 (R140_U524, R140_U180, R140_U181);
  nand ginst19314 (R140_U525, R140_U212, R140_U523);
  nand ginst19315 (R140_U526, R140_U44, U117);
  nand ginst19316 (R140_U527, SI_11_, R140_U45);
  nand ginst19317 (R140_U528, R140_U44, U117);
  nand ginst19318 (R140_U529, SI_11_, R140_U45);
  not ginst19319 (R140_U53, SI_18_);
  nand ginst19320 (R140_U530, R140_U528, R140_U529);
  nand ginst19321 (R140_U531, R140_U182, R140_U183);
  nand ginst19322 (R140_U532, R140_U314, R140_U530);
  nand ginst19323 (R140_U533, R140_U38, U118);
  nand ginst19324 (R140_U534, SI_10_, R140_U39);
  nand ginst19325 (R140_U535, R140_U38, U118);
  nand ginst19326 (R140_U536, SI_10_, R140_U39);
  nand ginst19327 (R140_U537, R140_U535, R140_U536);
  nand ginst19328 (R140_U538, R140_U184, R140_U185);
  nand ginst19329 (R140_U539, R140_U312, R140_U537);
  not ginst19330 (R140_U54, U110);
  nand ginst19331 (R140_U540, R140_U30, U120);
  nand ginst19332 (R140_U541, SI_0_, R140_U31);
  not ginst19333 (R140_U55, SI_19_);
  not ginst19334 (R140_U56, U109);
  not ginst19335 (R140_U57, SI_20_);
  not ginst19336 (R140_U58, U107);
  not ginst19337 (R140_U59, SI_21_);
  and ginst19338 (R140_U6, R140_U205, R140_U5);
  not ginst19339 (R140_U60, U106);
  not ginst19340 (R140_U61, SI_22_);
  not ginst19341 (R140_U62, U105);
  not ginst19342 (R140_U63, SI_23_);
  not ginst19343 (R140_U64, U104);
  not ginst19344 (R140_U65, SI_24_);
  not ginst19345 (R140_U66, U103);
  not ginst19346 (R140_U67, SI_25_);
  not ginst19347 (R140_U68, U102);
  not ginst19348 (R140_U69, SI_26_);
  and ginst19349 (R140_U7, R140_U209, R140_U213);
  not ginst19350 (R140_U70, U101);
  not ginst19351 (R140_U71, SI_27_);
  not ginst19352 (R140_U72, U100);
  not ginst19353 (R140_U73, SI_28_);
  not ginst19354 (R140_U74, U99);
  not ginst19355 (R140_U75, SI_29_);
  not ginst19356 (R140_U76, U98);
  not ginst19357 (R140_U77, SI_30_);
  not ginst19358 (R140_U78, U96);
  nand ginst19359 (R140_U79, SI_1_, SI_0_, U120);
  and ginst19360 (R140_U8, R140_U216, R140_U7);
  nand ginst19361 (R140_U80, R140_U217, R140_U300);
  nand ginst19362 (R140_U81, R140_U214, R140_U297);
  nand ginst19363 (R140_U82, R140_U206, R140_U293);
  nand ginst19364 (R140_U83, R140_U540, R140_U541);
  nand ginst19365 (R140_U84, R140_U330, R140_U331);
  nand ginst19366 (R140_U85, R140_U337, R140_U338);
  nand ginst19367 (R140_U86, R140_U344, R140_U345);
  nand ginst19368 (R140_U87, R140_U351, R140_U352);
  nand ginst19369 (R140_U88, R140_U358, R140_U359);
  nand ginst19370 (R140_U89, R140_U365, R140_U366);
  and ginst19371 (R140_U9, R140_U377, R140_U378);
  nand ginst19372 (R140_U90, R140_U372, R140_U373);
  nand ginst19373 (R140_U91, R140_U386, R140_U387);
  nand ginst19374 (R140_U92, R140_U393, R140_U394);
  nand ginst19375 (R140_U93, R140_U400, R140_U401);
  nand ginst19376 (R140_U94, R140_U407, R140_U408);
  nand ginst19377 (R140_U95, R140_U414, R140_U415);
  nand ginst19378 (R140_U96, R140_U421, R140_U422);
  nand ginst19379 (R140_U97, R140_U428, R140_U429);
  nand ginst19380 (R140_U98, R140_U435, R140_U436);
  nand ginst19381 (R140_U99, R140_U442, R140_U443);
  nand ginst19382 (U100, U285, U286);
  nand ginst19383 (U101, U287, U288);
  nand ginst19384 (U102, U289, U290);
  nand ginst19385 (U103, U291, U292);
  nand ginst19386 (U104, U293, U294);
  nand ginst19387 (U105, U295, U296);
  nand ginst19388 (U106, U297, U298);
  nand ginst19389 (U107, U299, U300);
  nand ginst19390 (U108, U301, U302);
  nand ginst19391 (U109, U303, U304);
  nand ginst19392 (U110, U305, U306);
  nand ginst19393 (U111, U307, U308);
  nand ginst19394 (U112, U309, U310);
  nand ginst19395 (U113, U311, U312);
  nand ginst19396 (U114, U313, U314);
  nand ginst19397 (U115, U315, U316);
  nand ginst19398 (U116, U317, U318);
  nand ginst19399 (U117, U319, U320);
  nand ginst19400 (U118, U321, U322);
  nand ginst19401 (U119, U323, U324);
  nand ginst19402 (U120, U325, U326);
  not ginst19403 (U121, P2_WR_REG_SCAN_IN);
  not ginst19404 (U122, P1_WR_REG_SCAN_IN);
  and ginst19405 (U123, U131, U132);
  not ginst19406 (U124, P2_RD_REG_SCAN_IN);
  not ginst19407 (U125, P1_RD_REG_SCAN_IN);
  and ginst19408 (U126, U133, U134);
  nand ginst19409 (U127, U128, U129);
  nand ginst19410 (U128, LT_1075_19_U6, LT_1075_U6, U125);
  nand ginst19411 (U129, P1_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_19__SCAN_IN, U124);
  not ginst19412 (U130, U127);
  nand ginst19413 (U131, P2_WR_REG_SCAN_IN, U122);
  nand ginst19414 (U132, P1_WR_REG_SCAN_IN, U121);
  nand ginst19415 (U133, P2_RD_REG_SCAN_IN, U125);
  nand ginst19416 (U134, P1_RD_REG_SCAN_IN, U124);
  nand ginst19417 (U135, P1_DATAO_REG_9__SCAN_IN, U127);
  nand ginst19418 (U136, R140_U84, U130);
  nand ginst19419 (U137, P1_DATAO_REG_8__SCAN_IN, U127);
  nand ginst19420 (U138, R140_U85, U130);
  nand ginst19421 (U139, P1_DATAO_REG_7__SCAN_IN, U127);
  nand ginst19422 (U140, R140_U86, U130);
  nand ginst19423 (U141, P1_DATAO_REG_6__SCAN_IN, U127);
  nand ginst19424 (U142, R140_U87, U130);
  nand ginst19425 (U143, P1_DATAO_REG_5__SCAN_IN, U127);
  nand ginst19426 (U144, R140_U88, U130);
  nand ginst19427 (U145, P1_DATAO_REG_4__SCAN_IN, U127);
  nand ginst19428 (U146, R140_U89, U130);
  nand ginst19429 (U147, P1_DATAO_REG_3__SCAN_IN, U127);
  nand ginst19430 (U148, R140_U90, U130);
  nand ginst19431 (U149, P1_DATAO_REG_31__SCAN_IN, U127);
  nand ginst19432 (U150, R140_U11, U130);
  nand ginst19433 (U151, P1_DATAO_REG_30__SCAN_IN, U127);
  nand ginst19434 (U152, R140_U91, U130);
  nand ginst19435 (U153, P1_DATAO_REG_2__SCAN_IN, U127);
  nand ginst19436 (U154, R140_U92, U130);
  nand ginst19437 (U155, P1_DATAO_REG_29__SCAN_IN, U127);
  nand ginst19438 (U156, R140_U93, U130);
  nand ginst19439 (U157, P1_DATAO_REG_28__SCAN_IN, U127);
  nand ginst19440 (U158, R140_U94, U130);
  nand ginst19441 (U159, P1_DATAO_REG_27__SCAN_IN, U127);
  nand ginst19442 (U160, R140_U95, U130);
  nand ginst19443 (U161, P1_DATAO_REG_26__SCAN_IN, U127);
  nand ginst19444 (U162, R140_U96, U130);
  nand ginst19445 (U163, P1_DATAO_REG_25__SCAN_IN, U127);
  nand ginst19446 (U164, R140_U97, U130);
  nand ginst19447 (U165, P1_DATAO_REG_24__SCAN_IN, U127);
  nand ginst19448 (U166, R140_U98, U130);
  nand ginst19449 (U167, P1_DATAO_REG_23__SCAN_IN, U127);
  nand ginst19450 (U168, R140_U99, U130);
  nand ginst19451 (U169, P1_DATAO_REG_22__SCAN_IN, U127);
  nand ginst19452 (U170, R140_U100, U130);
  nand ginst19453 (U171, P1_DATAO_REG_21__SCAN_IN, U127);
  nand ginst19454 (U172, R140_U101, U130);
  nand ginst19455 (U173, P1_DATAO_REG_20__SCAN_IN, U127);
  nand ginst19456 (U174, R140_U102, U130);
  nand ginst19457 (U175, P1_DATAO_REG_1__SCAN_IN, U127);
  nand ginst19458 (U176, R140_U10, U130);
  nand ginst19459 (U177, P1_DATAO_REG_19__SCAN_IN, U127);
  nand ginst19460 (U178, R140_U103, U130);
  nand ginst19461 (U179, P1_DATAO_REG_18__SCAN_IN, U127);
  nand ginst19462 (U180, R140_U104, U130);
  nand ginst19463 (U181, P1_DATAO_REG_17__SCAN_IN, U127);
  nand ginst19464 (U182, R140_U105, U130);
  nand ginst19465 (U183, P1_DATAO_REG_16__SCAN_IN, U127);
  nand ginst19466 (U184, R140_U106, U130);
  nand ginst19467 (U185, P1_DATAO_REG_15__SCAN_IN, U127);
  nand ginst19468 (U186, R140_U107, U130);
  nand ginst19469 (U187, P1_DATAO_REG_14__SCAN_IN, U127);
  nand ginst19470 (U188, R140_U108, U130);
  nand ginst19471 (U189, P1_DATAO_REG_13__SCAN_IN, U127);
  nand ginst19472 (U190, R140_U109, U130);
  nand ginst19473 (U191, P1_DATAO_REG_12__SCAN_IN, U127);
  nand ginst19474 (U192, R140_U110, U130);
  nand ginst19475 (U193, P1_DATAO_REG_11__SCAN_IN, U127);
  nand ginst19476 (U194, R140_U111, U130);
  nand ginst19477 (U195, P1_DATAO_REG_10__SCAN_IN, U127);
  nand ginst19478 (U196, R140_U112, U130);
  nand ginst19479 (U197, P1_DATAO_REG_0__SCAN_IN, U127);
  nand ginst19480 (U198, R140_U83, U130);
  nand ginst19481 (U199, R140_U84, U127);
  nand ginst19482 (U200, P2_DATAO_REG_9__SCAN_IN, U130);
  nand ginst19483 (U201, R140_U85, U127);
  nand ginst19484 (U202, P2_DATAO_REG_8__SCAN_IN, U130);
  nand ginst19485 (U203, R140_U86, U127);
  nand ginst19486 (U204, P2_DATAO_REG_7__SCAN_IN, U130);
  nand ginst19487 (U205, R140_U87, U127);
  nand ginst19488 (U206, P2_DATAO_REG_6__SCAN_IN, U130);
  nand ginst19489 (U207, R140_U88, U127);
  nand ginst19490 (U208, P2_DATAO_REG_5__SCAN_IN, U130);
  nand ginst19491 (U209, R140_U89, U127);
  nand ginst19492 (U210, P2_DATAO_REG_4__SCAN_IN, U130);
  nand ginst19493 (U211, R140_U90, U127);
  nand ginst19494 (U212, P2_DATAO_REG_3__SCAN_IN, U130);
  nand ginst19495 (U213, R140_U11, U127);
  nand ginst19496 (U214, P2_DATAO_REG_31__SCAN_IN, U130);
  nand ginst19497 (U215, R140_U91, U127);
  nand ginst19498 (U216, P2_DATAO_REG_30__SCAN_IN, U130);
  nand ginst19499 (U217, R140_U92, U127);
  nand ginst19500 (U218, P2_DATAO_REG_2__SCAN_IN, U130);
  nand ginst19501 (U219, R140_U93, U127);
  nand ginst19502 (U220, P2_DATAO_REG_29__SCAN_IN, U130);
  nand ginst19503 (U221, R140_U94, U127);
  nand ginst19504 (U222, P2_DATAO_REG_28__SCAN_IN, U130);
  nand ginst19505 (U223, R140_U95, U127);
  nand ginst19506 (U224, P2_DATAO_REG_27__SCAN_IN, U130);
  nand ginst19507 (U225, R140_U96, U127);
  nand ginst19508 (U226, P2_DATAO_REG_26__SCAN_IN, U130);
  nand ginst19509 (U227, R140_U97, U127);
  nand ginst19510 (U228, P2_DATAO_REG_25__SCAN_IN, U130);
  nand ginst19511 (U229, R140_U98, U127);
  nand ginst19512 (U230, P2_DATAO_REG_24__SCAN_IN, U130);
  nand ginst19513 (U231, R140_U99, U127);
  nand ginst19514 (U232, P2_DATAO_REG_23__SCAN_IN, U130);
  nand ginst19515 (U233, R140_U100, U127);
  nand ginst19516 (U234, P2_DATAO_REG_22__SCAN_IN, U130);
  nand ginst19517 (U235, R140_U101, U127);
  nand ginst19518 (U236, P2_DATAO_REG_21__SCAN_IN, U130);
  nand ginst19519 (U237, R140_U102, U127);
  nand ginst19520 (U238, P2_DATAO_REG_20__SCAN_IN, U130);
  nand ginst19521 (U239, R140_U10, U127);
  nand ginst19522 (U240, P2_DATAO_REG_1__SCAN_IN, U130);
  nand ginst19523 (U241, R140_U103, U127);
  nand ginst19524 (U242, P2_DATAO_REG_19__SCAN_IN, U130);
  nand ginst19525 (U243, R140_U104, U127);
  nand ginst19526 (U244, P2_DATAO_REG_18__SCAN_IN, U130);
  nand ginst19527 (U245, R140_U105, U127);
  nand ginst19528 (U246, P2_DATAO_REG_17__SCAN_IN, U130);
  nand ginst19529 (U247, R140_U106, U127);
  nand ginst19530 (U248, P2_DATAO_REG_16__SCAN_IN, U130);
  nand ginst19531 (U249, R140_U107, U127);
  nand ginst19532 (U25, U135, U136);
  nand ginst19533 (U250, P2_DATAO_REG_15__SCAN_IN, U130);
  nand ginst19534 (U251, R140_U108, U127);
  nand ginst19535 (U252, P2_DATAO_REG_14__SCAN_IN, U130);
  nand ginst19536 (U253, R140_U109, U127);
  nand ginst19537 (U254, P2_DATAO_REG_13__SCAN_IN, U130);
  nand ginst19538 (U255, R140_U110, U127);
  nand ginst19539 (U256, P2_DATAO_REG_12__SCAN_IN, U130);
  nand ginst19540 (U257, R140_U111, U127);
  nand ginst19541 (U258, P2_DATAO_REG_11__SCAN_IN, U130);
  nand ginst19542 (U259, R140_U112, U127);
  nand ginst19543 (U26, U137, U138);
  nand ginst19544 (U260, P2_DATAO_REG_10__SCAN_IN, U130);
  nand ginst19545 (U261, R140_U83, U127);
  nand ginst19546 (U262, P2_DATAO_REG_0__SCAN_IN, U130);
  nand ginst19547 (U263, P2_DATAO_REG_9__SCAN_IN, U127);
  nand ginst19548 (U264, P1_DATAO_REG_9__SCAN_IN, U130);
  nand ginst19549 (U265, P2_DATAO_REG_8__SCAN_IN, U127);
  nand ginst19550 (U266, P1_DATAO_REG_8__SCAN_IN, U130);
  nand ginst19551 (U267, P2_DATAO_REG_7__SCAN_IN, U127);
  nand ginst19552 (U268, P1_DATAO_REG_7__SCAN_IN, U130);
  nand ginst19553 (U269, P2_DATAO_REG_6__SCAN_IN, U127);
  nand ginst19554 (U27, U139, U140);
  nand ginst19555 (U270, P1_DATAO_REG_6__SCAN_IN, U130);
  nand ginst19556 (U271, P2_DATAO_REG_5__SCAN_IN, U127);
  nand ginst19557 (U272, P1_DATAO_REG_5__SCAN_IN, U130);
  nand ginst19558 (U273, P2_DATAO_REG_4__SCAN_IN, U127);
  nand ginst19559 (U274, P1_DATAO_REG_4__SCAN_IN, U130);
  nand ginst19560 (U275, P2_DATAO_REG_31__SCAN_IN, U127);
  nand ginst19561 (U276, P1_DATAO_REG_31__SCAN_IN, U130);
  nand ginst19562 (U277, P2_DATAO_REG_30__SCAN_IN, U127);
  nand ginst19563 (U278, P1_DATAO_REG_30__SCAN_IN, U130);
  nand ginst19564 (U279, P2_DATAO_REG_3__SCAN_IN, U127);
  nand ginst19565 (U28, U141, U142);
  nand ginst19566 (U280, P1_DATAO_REG_3__SCAN_IN, U130);
  nand ginst19567 (U281, P2_DATAO_REG_29__SCAN_IN, U127);
  nand ginst19568 (U282, P1_DATAO_REG_29__SCAN_IN, U130);
  nand ginst19569 (U283, P2_DATAO_REG_28__SCAN_IN, U127);
  nand ginst19570 (U284, P1_DATAO_REG_28__SCAN_IN, U130);
  nand ginst19571 (U285, P2_DATAO_REG_27__SCAN_IN, U127);
  nand ginst19572 (U286, P1_DATAO_REG_27__SCAN_IN, U130);
  nand ginst19573 (U287, P2_DATAO_REG_26__SCAN_IN, U127);
  nand ginst19574 (U288, P1_DATAO_REG_26__SCAN_IN, U130);
  nand ginst19575 (U289, P2_DATAO_REG_25__SCAN_IN, U127);
  nand ginst19576 (U29, U143, U144);
  nand ginst19577 (U290, P1_DATAO_REG_25__SCAN_IN, U130);
  nand ginst19578 (U291, P2_DATAO_REG_24__SCAN_IN, U127);
  nand ginst19579 (U292, P1_DATAO_REG_24__SCAN_IN, U130);
  nand ginst19580 (U293, P2_DATAO_REG_23__SCAN_IN, U127);
  nand ginst19581 (U294, P1_DATAO_REG_23__SCAN_IN, U130);
  nand ginst19582 (U295, P2_DATAO_REG_22__SCAN_IN, U127);
  nand ginst19583 (U296, P1_DATAO_REG_22__SCAN_IN, U130);
  nand ginst19584 (U297, P2_DATAO_REG_21__SCAN_IN, U127);
  nand ginst19585 (U298, P1_DATAO_REG_21__SCAN_IN, U130);
  nand ginst19586 (U299, P2_DATAO_REG_20__SCAN_IN, U127);
  nand ginst19587 (U30, U145, U146);
  nand ginst19588 (U300, P1_DATAO_REG_20__SCAN_IN, U130);
  nand ginst19589 (U301, P2_DATAO_REG_2__SCAN_IN, U127);
  nand ginst19590 (U302, P1_DATAO_REG_2__SCAN_IN, U130);
  nand ginst19591 (U303, P2_DATAO_REG_19__SCAN_IN, U127);
  nand ginst19592 (U304, P1_DATAO_REG_19__SCAN_IN, U130);
  nand ginst19593 (U305, P2_DATAO_REG_18__SCAN_IN, U127);
  nand ginst19594 (U306, P1_DATAO_REG_18__SCAN_IN, U130);
  nand ginst19595 (U307, P2_DATAO_REG_17__SCAN_IN, U127);
  nand ginst19596 (U308, P1_DATAO_REG_17__SCAN_IN, U130);
  nand ginst19597 (U309, P2_DATAO_REG_16__SCAN_IN, U127);
  nand ginst19598 (U31, U147, U148);
  nand ginst19599 (U310, P1_DATAO_REG_16__SCAN_IN, U130);
  nand ginst19600 (U311, P2_DATAO_REG_15__SCAN_IN, U127);
  nand ginst19601 (U312, P1_DATAO_REG_15__SCAN_IN, U130);
  nand ginst19602 (U313, P2_DATAO_REG_14__SCAN_IN, U127);
  nand ginst19603 (U314, P1_DATAO_REG_14__SCAN_IN, U130);
  nand ginst19604 (U315, P2_DATAO_REG_13__SCAN_IN, U127);
  nand ginst19605 (U316, P1_DATAO_REG_13__SCAN_IN, U130);
  nand ginst19606 (U317, P2_DATAO_REG_12__SCAN_IN, U127);
  nand ginst19607 (U318, P1_DATAO_REG_12__SCAN_IN, U130);
  nand ginst19608 (U319, P2_DATAO_REG_11__SCAN_IN, U127);
  nand ginst19609 (U32, U149, U150);
  nand ginst19610 (U320, P1_DATAO_REG_11__SCAN_IN, U130);
  nand ginst19611 (U321, P2_DATAO_REG_10__SCAN_IN, U127);
  nand ginst19612 (U322, P1_DATAO_REG_10__SCAN_IN, U130);
  nand ginst19613 (U323, P2_DATAO_REG_1__SCAN_IN, U127);
  nand ginst19614 (U324, P1_DATAO_REG_1__SCAN_IN, U130);
  nand ginst19615 (U325, P2_DATAO_REG_0__SCAN_IN, U127);
  nand ginst19616 (U326, P1_DATAO_REG_0__SCAN_IN, U130);
  nand ginst19617 (U33, U151, U152);
  nand ginst19618 (U34, U153, U154);
  nand ginst19619 (U35, U155, U156);
  nand ginst19620 (U36, U157, U158);
  nand ginst19621 (U37, U159, U160);
  nand ginst19622 (U38, U161, U162);
  nand ginst19623 (U39, U163, U164);
  nand ginst19624 (U40, U165, U166);
  nand ginst19625 (U41, U167, U168);
  nand ginst19626 (U42, U169, U170);
  nand ginst19627 (U43, U171, U172);
  nand ginst19628 (U44, U173, U174);
  nand ginst19629 (U45, U175, U176);
  nand ginst19630 (U46, U177, U178);
  nand ginst19631 (U47, U179, U180);
  nand ginst19632 (U48, U181, U182);
  nand ginst19633 (U49, U183, U184);
  nand ginst19634 (U50, U185, U186);
  nand ginst19635 (U51, U187, U188);
  nand ginst19636 (U52, U189, U190);
  nand ginst19637 (U53, U191, U192);
  nand ginst19638 (U54, U193, U194);
  nand ginst19639 (U55, U195, U196);
  nand ginst19640 (U56, U197, U198);
  nand ginst19641 (U57, U199, U200);
  nand ginst19642 (U58, U201, U202);
  nand ginst19643 (U59, U203, U204);
  nand ginst19644 (U60, U205, U206);
  nand ginst19645 (U61, U207, U208);
  nand ginst19646 (U62, U209, U210);
  nand ginst19647 (U63, U211, U212);
  nand ginst19648 (U64, U213, U214);
  nand ginst19649 (U65, U215, U216);
  nand ginst19650 (U66, U217, U218);
  nand ginst19651 (U67, U219, U220);
  nand ginst19652 (U68, U221, U222);
  nand ginst19653 (U69, U223, U224);
  nand ginst19654 (U70, U225, U226);
  nand ginst19655 (U71, U227, U228);
  nand ginst19656 (U72, U229, U230);
  nand ginst19657 (U73, U231, U232);
  nand ginst19658 (U74, U233, U234);
  nand ginst19659 (U75, U235, U236);
  nand ginst19660 (U76, U237, U238);
  nand ginst19661 (U77, U239, U240);
  nand ginst19662 (U78, U241, U242);
  nand ginst19663 (U79, U243, U244);
  nand ginst19664 (U80, U245, U246);
  nand ginst19665 (U81, U247, U248);
  nand ginst19666 (U82, U249, U250);
  nand ginst19667 (U83, U251, U252);
  nand ginst19668 (U84, U253, U254);
  nand ginst19669 (U85, U255, U256);
  nand ginst19670 (U86, U257, U258);
  nand ginst19671 (U87, U259, U260);
  nand ginst19672 (U88, U261, U262);
  nand ginst19673 (U89, U263, U264);
  nand ginst19674 (U90, U265, U266);
  nand ginst19675 (U91, U267, U268);
  nand ginst19676 (U92, U269, U270);
  nand ginst19677 (U93, U271, U272);
  nand ginst19678 (U94, U273, U274);
  nand ginst19679 (U95, U275, U276);
  nand ginst19680 (U96, U277, U278);
  nand ginst19681 (U97, U279, U280);
  nand ginst19682 (U98, U281, U282);
  nand ginst19683 (U99, U283, U284);

SatHard block1 (flip_signal, P1_U4199, U211, P1_R1117_U43, P1_R1282_U101, P1_SUB_84_U84, P1_SUB_84_U40, P1_R1207_U39, P1_R1192_U200, P1_IR_REG_20__SCAN_IN, P1_R1117_U91, P1_R1192_U145, P1_SUB_84_U224, P1_U3363, P1_R1150_U237, P1_R1282_U28, R140_U536, P1_U5731, P1_R1138_U251, P1_R1207_U51, P1_SUB_84_U72, SI_3_, P1_R1192_U191, P1_ADD_95_U89, P1_SUB_84_U243, P1_ADD_95_U151, P1_R1150_U38, P1_R1192_U185, U314, P1_IR_REG_25__SCAN_IN, R140_U31, P1_R1150_U190, P1_U5684, keyinput0, keyinput1, keyinput2, keyinput3, keyinput4, keyinput5, keyinput6, keyinput7, keyinput8, keyinput9, keyinput10, keyinput11, keyinput12, keyinput13, keyinput14, keyinput15, keyinput16, keyinput17, keyinput18, keyinput19, keyinput20, keyinput21, keyinput22, keyinput23, keyinput24, keyinput25, keyinput26, keyinput27, keyinput28, keyinput29, keyinput30, keyinput31);

endmodule
/*************** SatHard block ***************/
module SatHard (flip_signal, P1_U4199, U211, P1_R1117_U43, P1_R1282_U101, P1_SUB_84_U84, P1_SUB_84_U40, P1_R1207_U39, P1_R1192_U200, P1_IR_REG_20__SCAN_IN, P1_R1117_U91, P1_R1192_U145, P1_SUB_84_U224, P1_U3363, P1_R1150_U237, P1_R1282_U28, R140_U536, P1_U5731, P1_R1138_U251, P1_R1207_U51, P1_SUB_84_U72, SI_3_, P1_R1192_U191, P1_ADD_95_U89, P1_SUB_84_U243, P1_ADD_95_U151, P1_R1150_U38, P1_R1192_U185, U314, P1_IR_REG_25__SCAN_IN, R140_U31, P1_R1150_U190, P1_U5684, keyinput0, keyinput1, keyinput2, keyinput3, keyinput4, keyinput5, keyinput6, keyinput7, keyinput8, keyinput9, keyinput10, keyinput11, keyinput12, keyinput13, keyinput14, keyinput15, keyinput16, keyinput17, keyinput18, keyinput19, keyinput20, keyinput21, keyinput22, keyinput23, keyinput24, keyinput25, keyinput26, keyinput27, keyinput28, keyinput29, keyinput30, keyinput31);

  input P1_U4199, U211, P1_R1117_U43, P1_R1282_U101, P1_SUB_84_U84, P1_SUB_84_U40, P1_R1207_U39, P1_R1192_U200, P1_IR_REG_20__SCAN_IN, P1_R1117_U91, P1_R1192_U145, P1_SUB_84_U224, P1_U3363, P1_R1150_U237, P1_R1282_U28, R140_U536, P1_U5731, P1_R1138_U251, P1_R1207_U51, P1_SUB_84_U72, SI_3_, P1_R1192_U191, P1_ADD_95_U89, P1_SUB_84_U243, P1_ADD_95_U151, P1_R1150_U38, P1_R1192_U185, U314, P1_IR_REG_25__SCAN_IN, R140_U31, P1_R1150_U190, P1_U5684, keyinput0, keyinput1, keyinput2, keyinput3, keyinput4, keyinput5, keyinput6, keyinput7, keyinput8, keyinput9, keyinput10, keyinput11, keyinput12, keyinput13, keyinput14, keyinput15, keyinput16, keyinput17, keyinput18, keyinput19, keyinput20, keyinput21, keyinput22, keyinput23, keyinput24, keyinput25, keyinput26, keyinput27, keyinput28, keyinput29, keyinput30, keyinput31;
  output flip_signal;
  //SatHard key=10011010110001101101000011100100
  wire [31:0] sat_res_inputs;
  assign sat_res_inputs[31:0] = {P1_U4199, U211, P1_R1117_U43, P1_R1282_U101, P1_SUB_84_U84, P1_SUB_84_U40, P1_R1207_U39, P1_R1192_U200, P1_IR_REG_20__SCAN_IN, P1_R1117_U91, P1_R1192_U145, P1_SUB_84_U224, P1_U3363, P1_R1150_U237, P1_R1282_U28, R140_U536, P1_U5731, P1_R1138_U251, P1_R1207_U51, P1_SUB_84_U72, SI_3_, P1_R1192_U191, P1_ADD_95_U89, P1_SUB_84_U243, P1_ADD_95_U151, P1_R1150_U38, P1_R1192_U185, U314, P1_IR_REG_25__SCAN_IN, R140_U31, P1_R1150_U190, P1_U5684};
  wire [31:0] keyinputs, keyvalue;
  assign keyinputs[31:0] = {keyinput0, keyinput1, keyinput2, keyinput3, keyinput4, keyinput5, keyinput6, keyinput7, keyinput8, keyinput9, keyinput10, keyinput11, keyinput12, keyinput13, keyinput14, keyinput15, keyinput16, keyinput17, keyinput18, keyinput19, keyinput20, keyinput21, keyinput22, keyinput23, keyinput24, keyinput25, keyinput26, keyinput27, keyinput28, keyinput29, keyinput30, keyinput31};
  assign keyvalue[31:0] = 32'b10011010110001101101000011100100;

  integer ham_dist_peturb, idx;
  wire [31:0] diff;
  assign diff = sat_res_inputs ^ keyvalue;

  always@* begin
    ham_dist_peturb = 0;
    for(idx=0; idx<32; idx=idx+1) ham_dist_peturb = ham_dist_peturb + diff[idx];
  end

  integer ham_dist_restore, idx;
  wire [31:0] diff;
  assign diff = sat_res_inputs ^ keyinputs;

  always@* begin
    ham_dist_restore = 0;
    for(idx=0; idx<32; idx=idx+1) ham_dist_restore = ham_dist_restore + diff[idx];
  end

  assign flip_signal = ( (ham_dist_peturb==0) ^ (ham_dist_restore==0) ) ? 'b1 : 'b0;
endmodule
/*************** SatHard block ***************/
