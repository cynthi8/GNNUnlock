// Main module
module c2670(1, 2, 3, 4, 5, 6, 7, 8, 11, 14, 15, 16, 19, 20, 21, 22, 23, 24, 25, 26, 27, 28, 29, 32, 33, 34, 35, 36, 37, 40, 43, 44, 47, 48, 49, 50, 51, 52, 53, 54, 55, 56, 57, 60, 61, 62, 63, 64, 65, 66, 67, 68, 69, 72, 73, 74, 75, 76, 77, 78, 79, 80, 81, 82, 85, 86, 87, 88, 89, 90, 91, 92, 93, 94, 95, 96, 99, 100, 101, 102, 103, 104, 105, 106, 107, 108, 111, 112, 113, 114, 115, 116, 117, 118, 119, 120, 123, 124, 125, 126, 127, 128, 129, 130, 131, 132, 135, 136, 137, 138, 139, 140, 141, 142, 143, 144, 145, 146, 147, 148, 149, 150, 151, 152, 153, 154, 155, 156, 157, 158, 159, 160, 161, 162, 163, 164, 165, 166, 167, 168, 169, 170, 171, 172, 173, 174, 175, 176, 177, 178, 179, 180, 181, 182, 183, 184, 185, 186, 187, 188, 189, 190, 191, 192, 193, 194, 195, 196, 197, 198, 199, 200, 201, 202, 203, 204, 205, 206, 207, 208, 209, 210, 211, 212, 213, 214, 215, 216, 217, 218, 219, 224, 227, 230, 231, 234, 237, 241, 246, 253, 256, 259, 262, 263, 266, 269, 272, 275, 278, 281, 284, 287, 290, 294, 297, 301, 305, 309, 313, 316, 319, 322, 325, 328, 331, 334, 337, 340, 343, 346, 349, 352, 355, 143, 144, 145, 146, 147, 148, 149, 150, 151, 152, 153, 154, 155, 156, 157, 158, 159, 160, 161, 162, 163, 164, 165, 166, 167, 168, 169, 170, 171, 172, 173, 174, 175, 176, 177, 178, 179, 180, 181, 182, 183, 184, 185, 186, 187, 188, 189, 190, 191, 192, 193, 194, 195, 196, 197, 198, 199, 200, 201, 202, 203, 204, 205, 206, 207, 208, 209, 210, 211, 212, 213, 214, 215, 216, 217, 218, 398, 400, 401, 419, 420, 456, 457, 458, 487, 488, 489, 490, 491, 492, 493, 494, 792, 799, 805, 1026, 1028, 1029, 1269, 1277, 1448, 1726, 1816, 1817, 1818, 1819, 1820, 1821, 1969, 1970, 1971, 2010, 2012, 2014, 2016, 2018, 2020, 2022, 2387, 2388, 2389, 2390, 2496, 2643, 2644, 2891, 2925, 2970, 2971, 3038, 3079, 3546, 3671, 3803, 3804, 3809, 3851, 3875, 3881, 3882);

  input 1, 2, 3, 4, 5, 6, 7, 8, 11, 14, 15, 16, 19, 20, 21, 22, 23, 24, 25, 26, 27, 28, 29, 32, 33, 34, 35, 36, 37, 40, 43, 44, 47, 48, 49, 50, 51, 52, 53, 54, 55, 56, 57, 60, 61, 62, 63, 64, 65, 66, 67, 68, 69, 72, 73, 74, 75, 76, 77, 78, 79, 80, 81, 82, 85, 86, 87, 88, 89, 90, 91, 92, 93, 94, 95, 96, 99, 100, 101, 102, 103, 104, 105, 106, 107, 108, 111, 112, 113, 114, 115, 116, 117, 118, 119, 120, 123, 124, 125, 126, 127, 128, 129, 130, 131, 132, 135, 136, 137, 138, 139, 140, 141, 142, 143, 144, 145, 146, 147, 148, 149, 150, 151, 152, 153, 154, 155, 156, 157, 158, 159, 160, 161, 162, 163, 164, 165, 166, 167, 168, 169, 170, 171, 172, 173, 174, 175, 176, 177, 178, 179, 180, 181, 182, 183, 184, 185, 186, 187, 188, 189, 190, 191, 192, 193, 194, 195, 196, 197, 198, 199, 200, 201, 202, 203, 204, 205, 206, 207, 208, 209, 210, 211, 212, 213, 214, 215, 216, 217, 218, 219, 224, 227, 230, 231, 234, 237, 241, 246, 253, 256, 259, 262, 263, 266, 269, 272, 275, 278, 281, 284, 287, 290, 294, 297, 301, 305, 309, 313, 316, 319, 322, 325, 328, 331, 334, 337, 340, 343, 346, 349, 352, 355;
  output 143, 144, 145, 146, 147, 148, 149, 150, 151, 152, 153, 154, 155, 156, 157, 158, 159, 160, 161, 162, 163, 164, 165, 166, 167, 168, 169, 170, 171, 172, 173, 174, 175, 176, 177, 178, 179, 180, 181, 182, 183, 184, 185, 186, 187, 188, 189, 190, 191, 192, 193, 194, 195, 196, 197, 198, 199, 200, 201, 202, 203, 204, 205, 206, 207, 208, 209, 210, 211, 212, 213, 214, 215, 216, 217, 218, 398, 400, 401, 419, 420, 456, 457, 458, 487, 488, 489, 490, 491, 492, 493, 494, 792, 799, 805, 1026, 1028, 1029, 1269, 1277, 1448, 1726, 1816, 1817, 1818, 1819, 1820, 1821, 1969, 1970, 1971, 2010, 2012, 2014, 2016, 2018, 2020, 2022, 2387, 2388, 2389, 2390, 2496, 2643, 2644, 2891, 2925, 2970, 2971, 3038, 3079, 3546, 3671, 3803, 3804, 3809, 3851, 3875, 3881, 3882;
  wire 405, 408, 425, 485, 486, 495, 496, 499, 500, 503, 506, 509, 521, 533, 537, 543, 544, 547, 550, 562, 574, 578, 582, 594, 606, 607, 608, 609, 610, 611, 612, 613, 625, 637, 643, 650, 651, 655, 659, 663, 667, 671, 675, 679, 683, 687, 693, 699, 705, 711, 715, 719, 723, 727, 730, 733, 734, 735, 738, 741, 744, 747, 750, 753, 756, 759, 762, 765, 768, 771, 774, 777, 780, 783, 786, 800, 900, 901, 902, 903, 904, 905, 998, 999, 1027, 1032, 1033, 1034, 1037, 1042, 1053, 1064, 1065, 1066, 1067, 1068, 1069, 1070, 1075, 1086, 1097, 1098, 1099, 1100, 1101, 1102, 1113, 1124, 1125, 1126, 1127, 1128, 1129, 1133, 1137, 1140, 1141, 1142, 1143, 1144, 1145, 1146, 1157, 1168, 1169, 1170, 1171, 1172, 1173, 1178, 1184, 1185, 1186, 1187, 1188, 1189, 1190, 1195, 1200, 1205, 1210, 1211, 1212, 1213, 1214, 1215, 1216, 1219, 1222, 1225, 1228, 1231, 1234, 1237, 1240, 1243, 1246, 1249, 1250, 1251, 1254, 1257, 1260, 1263, 1266, 1275, 1276, 1302, 1351, 1352, 1353, 1354, 1355, 1395, 1396, 1397, 1398, 1399, 1422, 1423, 1424, 1425, 1426, 1427, 1440, 1441, 1449, 1450, 1451, 1452, 1453, 1454, 1455, 1456, 1457, 1458, 1459, 1460, 1461, 1462, 1463, 1464, 1465, 1466, 1467, 1468, 1469, 1470, 1471, 1472, 1473, 1474, 1475, 1476, 1477, 1478, 1479, 1480, 1481, 1482, 1483, 1484, 1485, 1486, 1487, 1488, 1489, 1490, 1491, 1492, 1493, 1494, 1495, 1496, 1499, 1502, 1506, 1510, 1513, 1516, 1519, 1520, 1521, 1522, 1523, 1524, 1525, 1526, 1527, 1528, 1529, 1530, 1531, 1532, 1533, 1534, 1535, 1536, 1537, 1538, 1539, 1540, 1541, 1542, 1543, 1544, 1545, 1546, 1547, 1548, 1549, 1550, 1551, 1552, 1553, 1557, 1561, 1564, 1565, 1566, 1567, 1568, 1569, 1570, 1571, 1572, 1573, 1574, 1575, 1576, 1577, 1578, 1581, 1582, 1585, 1588, 1591, 1596, 1600, 1606, 1612, 1615, 1619, 1624, 1628, 1631, 1634, 1637, 1642, 1647, 1651, 1656, 1676, 1681, 1686, 1690, 1708, 1770, 1773, 1776, 1777, 1778, 1781, 1784, 1785, 1795, 1798, 1801, 1804, 1807, 1808, 1809, 1810, 1811, 1813, 1814, 1815, 1822, 1823, 1824, 1827, 1830, 1831, 1832, 1833, 1836, 1841, 1848, 1852, 1856, 1863, 1870, 1875, 1880, 1885, 1888, 1891, 1894, 1897, 1908, 1909, 1910, 1911, 1912, 1913, 1914, 1915, 1916, 1917, 1918, 1919, 1928, 1929, 1930, 1931, 1932, 1933, 1934, 1935, 1936, 1939, 1940, 1941, 1942, 1945, 1948, 1951, 1954, 1957, 1960, 1963, 1966, 2028, 2029, 2030, 2031, 2032, 2033, 2034, 2040, 2041, 2042, 2043, 2046, 2049, 2052, 2055, 2058, 2061, 2064, 2067, 2070, 2073, 2076, 2079, 2095, 2098, 2101, 2104, 2107, 2110, 2113, 2119, 2120, 2125, 2126, 2127, 2128, 2135, 2141, 2144, 2147, 2150, 2153, 2154, 2155, 2156, 2157, 2158, 2171, 2172, 2173, 2174, 2175, 2176, 2177, 2178, 2185, 2188, 2191, 2194, 2197, 2200, 2201, 2204, 2207, 2210, 2213, 2216, 2219, 2234, 2235, 2236, 2237, 2250, 2266, 2269, 2291, 2294, 2297, 2298, 2300, 2301, 2302, 2303, 2304, 2305, 2306, 2307, 2308, 2309, 2310, 2311, 2312, 2313, 2314, 2315, 2316, 2317, 2318, 2319, 2320, 2321, 2322, 2323, 2324, 2325, 2326, 2327, 2328, 2329, 2330, 2331, 2332, 2333, 2334, 2335, 2336, 2337, 2338, 2339, 2340, 2354, 2355, 2356, 2357, 2358, 2359, 2364, 2365, 2366, 2367, 2368, 2372, 2373, 2374, 2375, 2376, 2377, 2382, 2386, 2391, 2395, 2400, 2403, 2406, 2407, 2408, 2409, 2410, 2411, 2412, 2413, 2414, 2415, 2416, 2417, 2421, 2425, 2428, 2429, 2430, 2431, 2432, 2433, 2434, 2437, 2440, 2443, 2446, 2449, 2452, 2453, 2454, 2457, 2460, 2463, 2466, 2469, 2472, 2475, 2478, 2481, 2484, 2487, 2490, 2493, 2503, 2504, 2510, 2511, 2521, 2528, 2531, 2534, 2537, 2540, 2544, 2545, 2546, 2547, 2548, 2549, 2550, 2551, 2552, 2553, 2563, 2564, 2565, 2566, 2567, 2568, 2579, 2603, 2607, 2608, 2609, 2610, 2611, 2612, 2613, 2617, 2618, 2619, 2620, 2621, 2624, 2628, 2629, 2630, 2631, 2632, 2633, 2634, 2635, 2636, 2638, 2645, 2646, 2652, 2655, 2656, 2659, 2663, 2664, 2665, 2666, 2667, 2668, 2669, 2670, 2671, 2672, 2673, 2674, 2675, 2676, 2677, 2678, 2679, 2680, 2681, 2684, 2687, 2690, 2693, 2694, 2695, 2696, 2697, 2698, 2699, 2700, 2701, 2702, 2703, 2706, 2707, 2708, 2709, 2710, 2719, 2720, 2726, 2729, 2738, 2743, 2747, 2748, 2749, 2750, 2751, 2760, 2761, 2766, 2771, 2772, 2773, 2774, 2775, 2776, 2777, 2778, 2781, 2782, 2783, 2784, 2789, 2790, 2791, 2792, 2793, 2796, 2800, 2803, 2806, 2809, 2810, 2811, 2812, 2817, 2820, 2826, 2829, 2830, 2831, 2837, 2838, 2839, 2840, 2841, 2844, 2854, 2859, 2869, 2874, 2877, 2880, 2881, 2882, 2885, 2888, 2894, 2895, 2896, 2897, 2898, 2899, 2900, 2901, 2914, 2915, 2916, 2917, 2918, 2919, 2920, 2921, 2931, 2938, 2939, 2963, 2972, 2975, 2978, 2981, 2984, 2985, 2986, 2989, 2992, 2995, 2998, 3001, 3004, 3007, 3008, 3009, 3010, 3013, 3016, 3019, 3022, 3025, 3028, 3029, 3030, 3035, 3036, 3037, 3039, 3044, 3045, 3046, 3047, 3048, 3049, 3050, 3053, 3054, 3055, 3056, 3057, 3058, 3059, 3060, 3061, 3064, 3065, 3066, 3067, 3068, 3069, 3070, 3071, 3072, 3073, 3074, 3075, 3076, 3088, 3091, 3110, 3113, 3137, 3140, 3143, 3146, 3149, 3152, 3157, 3160, 3163, 3166, 3169, 3172, 3175, 3176, 3177, 3178, 3180, 3187, 3188, 3189, 3190, 3191, 3192, 3193, 3194, 3195, 3196, 3197, 3208, 3215, 3216, 3217, 3218, 3219, 3220, 3222, 3223, 3230, 3231, 3238, 3241, 3244, 3247, 3250, 3253, 3256, 3259, 3262, 3265, 3268, 3271, 3274, 3277, 3281, 3282, 3283, 3284, 3286, 3288, 3289, 3291, 3293, 3295, 3296, 3299, 3301, 3302, 3304, 3306, 3308, 3309, 3312, 3314, 3315, 3318, 3321, 3324, 3327, 3330, 3333, 3334, 3335, 3336, 3337, 3340, 3344, 3348, 3352, 3356, 3360, 3364, 3367, 3370, 3374, 3378, 3382, 3386, 3390, 3394, 3397, 3400, 3401, 3402, 3403, 3404, 3405, 3406, 3409, 3410, 3412, 3414, 3416, 3418, 3420, 3422, 3428, 3430, 3432, 3434, 3436, 3438, 3440, 3450, 3453, 3456, 3459, 3478, 3479, 3480, 3481, 3482, 3483, 3484, 3485, 3486, 3487, 3488, 3489, 3490, 3491, 3492, 3493, 3494, 3496, 3498, 3499, 3500, 3501, 3502, 3503, 3504, 3505, 3506, 3507, 3508, 3509, 3510, 3511, 3512, 3513, 3515, 3517, 3522, 3525, 3528, 3531, 3534, 3537, 3540, 3543, 3551, 3552, 3553, 3554, 3555, 3556, 3557, 3558, 3559, 3563, 3564, 3565, 3566, 3567, 3568, 3569, 3570, 3576, 3579, 3585, 3588, 3592, 3593, 3594, 3595, 3596, 3597, 3598, 3599, 3600, 3603, 3608, 3612, 3615, 3616, 3622, 3629, 3630, 3631, 3632, 3633, 3634, 3635, 3640, 3644, 3647, 3648, 3654, 3661, 3662, 3667, 3668, 3669, 3670, 3691, 3692, 3693, 3694, 3695, 3696, 3697, 3716, 3717, 3718, 3719, 3720, 3721, 3722, 3723, 3726, 3727, 3728, 3729, 3730, 3731, 3732, 3733, 3734, 3735, 3736, 3737, 3740, 3741, 3742, 3743, 3744, 3745, 3746, 3747, 3748, 3749, 3750, 3753, 3754, 3758, 3761, 3762, 3767, 3771, 3774, 3775, 3778, 3779, 3780, 3790, 3793, 3794, 3802, 3805, 3806, 3807, 3808, 3811, 3812, 3813, 3814, 3815, 3816, 3817, 3818, 3819, 3820, 3821, 3822, 3823, 3826, 3827, 3834, 3835, 3836, 3837, 3838, 3839, 3840, 3843, 3852, 3857, 3858, 3859, 3864, 3869, 3870, 3876, 3877;

  and ginst1 (1026, 94, 500);
  and ginst2 (1027, 325, 651);
  not ginst3 (1028, 651);
  nand ginst4 (1029, 231, 651);
  not ginst5 (1032, 544);
  not ginst6 (1033, 547);
  and ginst7 (1034, 547, 544);
  buf ginst8 (1037, 503);
  not ginst9 (1042, 509);
  not ginst10 (1053, 521);
  and ginst11 (1064, 80, 509, 521);
  and ginst12 (1065, 68, 509, 521);
  and ginst13 (1066, 79, 509, 521);
  and ginst14 (1067, 78, 509, 521);
  and ginst15 (1068, 77, 509, 521);
  and ginst16 (1069, 11, 537);
  buf ginst17 (1070, 503);
  not ginst18 (1075, 550);
  not ginst19 (1086, 562);
  and ginst20 (1097, 76, 550, 562);
  and ginst21 (1098, 75, 550, 562);
  and ginst22 (1099, 74, 550, 562);
  and ginst23 (1100, 73, 550, 562);
  and ginst24 (1101, 72, 550, 562);
  not ginst25 (1102, 582);
  not ginst26 (1113, 594);
  and ginst27 (1124, 114, 582, 594);
  and ginst28 (1125, 113, 582, 594);
  and ginst29 (1126, 112, 582, 594);
  and ginst30 (1127, 111, 582, 594);
  and ginst31 (1128, 582, 594);
  nand ginst32 (1129, 900, 901);
  nand ginst33 (1133, 902, 903);
  nand ginst34 (1137, 904, 905);
  not ginst35 (1140, 741);
  nand ginst36 (1141, 741, 612);
  not ginst37 (1142, 744);
  not ginst38 (1143, 747);
  not ginst39 (1144, 750);
  not ginst40 (1145, 753);
  not ginst41 (1146, 613);
  not ginst42 (1157, 625);
  and ginst43 (1168, 118, 613, 625);
  and ginst44 (1169, 107, 613, 625);
  and ginst45 (1170, 117, 613, 625);
  and ginst46 (1171, 116, 613, 625);
  and ginst47 (1172, 115, 613, 625);
  not ginst48 (1173, 637);
  not ginst49 (1178, 643);
  not ginst50 (1184, 768);
  nand ginst51 (1185, 768, 650);
  not ginst52 (1186, 771);
  not ginst53 (1187, 774);
  not ginst54 (1188, 777);
  not ginst55 (1189, 780);
  buf ginst56 (1190, 506);
  buf ginst57 (1195, 506);
  not ginst58 (1200, 693);
  not ginst59 (1205, 699);
  not ginst60 (1210, 735);
  not ginst61 (1211, 738);
  not ginst62 (1212, 756);
  not ginst63 (1213, 759);
  not ginst64 (1214, 762);
  not ginst65 (1215, 765);
  nand ginst66 (1216, 998, 999);
  buf ginst67 (1219, 574);
  buf ginst68 (1222, 578);
  buf ginst69 (1225, 655);
  buf ginst70 (1228, 659);
  buf ginst71 (1231, 663);
  buf ginst72 (1234, 667);
  buf ginst73 (1237, 671);
  buf ginst74 (1240, 675);
  buf ginst75 (1243, 679);
  buf ginst76 (1246, 683);
  not ginst77 (1249, 783);
  not ginst78 (1250, 786);
  buf ginst79 (1251, 687);
  buf ginst80 (1254, 705);
  buf ginst81 (1257, 711);
  buf ginst82 (1260, 715);
  buf ginst83 (1263, 719);
  buf ginst84 (1266, 723);
  not ginst85 (1269, 1027);
  and ginst86 (1275, 325, 1032);
  and ginst87 (1276, 231, 1033);
  buf ginst88 (1277, 1034);
  or ginst89 (1302, 1069, 543);
  nand ginst90 (1351, 352, 1140);
  nand ginst91 (1352, 747, 1142);
  nand ginst92 (1353, 744, 1143);
  nand ginst93 (1354, 753, 1144);
  nand ginst94 (1355, 750, 1145);
  nand ginst95 (1395, 355, 1184);
  nand ginst96 (1396, 774, 1186);
  nand ginst97 (1397, 771, 1187);
  nand ginst98 (1398, 780, 1188);
  nand ginst99 (1399, 777, 1189);
  nand ginst100 (1422, 738, 1210);
  nand ginst101 (1423, 735, 1211);
  nand ginst102 (1424, 759, 1212);
  nand ginst103 (1425, 756, 1213);
  nand ginst104 (1426, 765, 1214);
  nand ginst105 (1427, 762, 1215);
  nand ginst106 (1440, 786, 1249);
  nand ginst107 (1441, 783, 1250);
  not ginst108 (1448, 1034);
  not ginst109 (1449, 1275);
  not ginst110 (1450, 1276);
  and ginst111 (1451, 93, 1042, 1053);
  and ginst112 (1452, 55, 509, 1053);
  and ginst113 (1453, 67, 1042, 521);
  and ginst114 (1454, 81, 1042, 1053);
  and ginst115 (1455, 43, 509, 1053);
  and ginst116 (1456, 56, 1042, 521);
  and ginst117 (1457, 92, 1042, 1053);
  and ginst118 (1458, 54, 509, 1053);
  and ginst119 (1459, 66, 1042, 521);
  and ginst120 (1460, 91, 1042, 1053);
  and ginst121 (1461, 53, 509, 1053);
  and ginst122 (1462, 65, 1042, 521);
  and ginst123 (1463, 90, 1042, 1053);
  and ginst124 (1464, 52, 509, 1053);
  and ginst125 (1465, 64, 1042, 521);
  and ginst126 (1466, 89, 1075, 1086);
  and ginst127 (1467, 51, 550, 1086);
  and ginst128 (1468, 63, 1075, 562);
  and ginst129 (1469, 88, 1075, 1086);
  and ginst130 (1470, 50, 550, 1086);
  and ginst131 (1471, 62, 1075, 562);
  and ginst132 (1472, 87, 1075, 1086);
  and ginst133 (1473, 49, 550, 1086);
  and ginst134 (1474, 1075, 562);
  and ginst135 (1475, 86, 1075, 1086);
  and ginst136 (1476, 48, 550, 1086);
  and ginst137 (1477, 61, 1075, 562);
  and ginst138 (1478, 85, 1075, 1086);
  and ginst139 (1479, 47, 550, 1086);
  and ginst140 (1480, 60, 1075, 562);
  and ginst141 (1481, 138, 1102, 1113);
  and ginst142 (1482, 102, 582, 1113);
  and ginst143 (1483, 126, 1102, 594);
  and ginst144 (1484, 137, 1102, 1113);
  and ginst145 (1485, 101, 582, 1113);
  and ginst146 (1486, 125, 1102, 594);
  and ginst147 (1487, 136, 1102, 1113);
  and ginst148 (1488, 100, 582, 1113);
  and ginst149 (1489, 124, 1102, 594);
  and ginst150 (1490, 135, 1102, 1113);
  and ginst151 (1491, 99, 582, 1113);
  and ginst152 (1492, 123, 1102, 594);
  and ginst153 (1493, 1102, 1113);
  and ginst154 (1494, 582, 1113);
  and ginst155 (1495, 1102, 594);
  not ginst156 (1496, 1129);
  not ginst157 (1499, 1133);
  nand ginst158 (1502, 1351, 1141);
  nand ginst159 (1506, 1352, 1353);
  nand ginst160 (1510, 1354, 1355);
  buf ginst161 (1513, 1137);
  buf ginst162 (1516, 1137);
  not ginst163 (1519, 1219);
  not ginst164 (1520, 1222);
  not ginst165 (1521, 1225);
  not ginst166 (1522, 1228);
  not ginst167 (1523, 1231);
  not ginst168 (1524, 1234);
  not ginst169 (1525, 1237);
  not ginst170 (1526, 1240);
  not ginst171 (1527, 1243);
  not ginst172 (1528, 1246);
  and ginst173 (1529, 142, 1146, 1157);
  and ginst174 (1530, 106, 613, 1157);
  and ginst175 (1531, 130, 1146, 625);
  and ginst176 (1532, 131, 1146, 1157);
  and ginst177 (1533, 95, 613, 1157);
  and ginst178 (1534, 119, 1146, 625);
  and ginst179 (1535, 141, 1146, 1157);
  and ginst180 (1536, 105, 613, 1157);
  and ginst181 (1537, 129, 1146, 625);
  and ginst182 (1538, 140, 1146, 1157);
  and ginst183 (1539, 104, 613, 1157);
  and ginst184 (1540, 128, 1146, 625);
  and ginst185 (1541, 139, 1146, 1157);
  and ginst186 (1542, 103, 613, 1157);
  and ginst187 (1543, 127, 1146, 625);
  and ginst188 (1544, 19, 1173);
  and ginst189 (1545, 4, 1173);
  and ginst190 (1546, 20, 1173);
  and ginst191 (1547, 5, 1173);
  and ginst192 (1548, 21, 1178);
  and ginst193 (1549, 22, 1178);
  and ginst194 (1550, 23, 1178);
  and ginst195 (1551, 6, 1178);
  and ginst196 (1552, 24, 1178);
  nand ginst197 (1553, 1395, 1185);
  nand ginst198 (1557, 1396, 1397);
  nand ginst199 (1561, 1398, 1399);
  and ginst200 (1564, 25, 1200);
  and ginst201 (1565, 32, 1200);
  and ginst202 (1566, 26, 1200);
  and ginst203 (1567, 33, 1200);
  and ginst204 (1568, 27, 1205);
  and ginst205 (1569, 34, 1205);
  and ginst206 (1570, 35, 1205);
  and ginst207 (1571, 28, 1205);
  not ginst208 (1572, 1251);
  not ginst209 (1573, 1254);
  not ginst210 (1574, 1257);
  not ginst211 (1575, 1260);
  not ginst212 (1576, 1263);
  not ginst213 (1577, 1266);
  nand ginst214 (1578, 1422, 1423);
  not ginst215 (1581, 1216);
  nand ginst216 (1582, 1426, 1427);
  nand ginst217 (1585, 1424, 1425);
  nand ginst218 (1588, 1440, 1441);
  and ginst219 (1591, 1449, 1450);
  or ginst220 (1596, 1451, 1452, 1453, 1064);
  or ginst221 (1600, 1454, 1455, 1456, 1065);
  or ginst222 (1606, 1457, 1458, 1459, 1066);
  or ginst223 (1612, 1460, 1461, 1462, 1067);
  or ginst224 (1615, 1463, 1464, 1465, 1068);
  or ginst225 (1619, 1466, 1467, 1468, 1097);
  or ginst226 (1624, 1469, 1470, 1471, 1098);
  or ginst227 (1628, 1472, 1473, 1474, 1099);
  or ginst228 (1631, 1475, 1476, 1477, 1100);
  or ginst229 (1634, 1478, 1479, 1480, 1101);
  or ginst230 (1637, 1481, 1482, 1483, 1124);
  or ginst231 (1642, 1484, 1485, 1486, 1125);
  or ginst232 (1647, 1487, 1488, 1489, 1126);
  or ginst233 (1651, 1490, 1491, 1492, 1127);
  or ginst234 (1656, 1493, 1494, 1495, 1128);
  or ginst235 (1676, 1532, 1533, 1534, 1169);
  or ginst236 (1681, 1535, 1536, 1537, 1170);
  or ginst237 (1686, 1538, 1539, 1540, 1171);
  or ginst238 (1690, 1541, 1542, 1543, 1172);
  or ginst239 (1708, 1529, 1530, 1531, 1168);
  buf ginst240 (1726, 1591);
  not ginst241 (1770, 1502);
  not ginst242 (1773, 1506);
  not ginst243 (1776, 1513);
  not ginst244 (1777, 1516);
  buf ginst245 (1778, 1510);
  buf ginst246 (1781, 1510);
  and ginst247 (1784, 1133, 1129, 1513);
  and ginst248 (1785, 1499, 1496, 1516);
  not ginst249 (1795, 1553);
  not ginst250 (1798, 1557);
  buf ginst251 (1801, 1561);
  buf ginst252 (1804, 1561);
  not ginst253 (1807, 1588);
  not ginst254 (1808, 1578);
  nand ginst255 (1809, 1578, 1581);
  not ginst256 (1810, 1582);
  not ginst257 (1811, 1585);
  and ginst258 (1813, 1596, 241);
  and ginst259 (1814, 1606, 241);
  and ginst260 (1815, 1600, 241);
  not ginst261 (1816, 1642);
  not ginst262 (1817, 1647);
  not ginst263 (1818, 1637);
  not ginst264 (1819, 1624);
  not ginst265 (1820, 1619);
  not ginst266 (1821, 1615);
  and ginst267 (1822, 496, 224, 36, 1591);
  and ginst268 (1823, 496, 224, 1591, 486);
  buf ginst269 (1824, 1596);
  not ginst270 (1827, 1606);
  and ginst271 (1830, 1600, 537);
  and ginst272 (1831, 1606, 537);
  and ginst273 (1832, 1619, 246);
  not ginst274 (1833, 1596);
  not ginst275 (1836, 1600);
  not ginst276 (1841, 1606);
  buf ginst277 (1848, 1612);
  buf ginst278 (1852, 1615);
  buf ginst279 (1856, 1619);
  buf ginst280 (1863, 1624);
  buf ginst281 (1870, 1628);
  buf ginst282 (1875, 1631);
  buf ginst283 (1880, 1634);
  nand ginst284 (1885, 727, 1651);
  nand ginst285 (1888, 730, 1656);
  buf ginst286 (1891, 1686);
  and ginst287 (1894, 1637, 425);
  not ginst288 (1897, 1642);
  and ginst289 (1908, 1496, 1133, 1776);
  and ginst290 (1909, 1129, 1499, 1777);
  and ginst291 (1910, 1600, 637);
  and ginst292 (1911, 1606, 637);
  and ginst293 (1912, 1612, 637);
  and ginst294 (1913, 1615, 637);
  and ginst295 (1914, 1619, 643);
  and ginst296 (1915, 1624, 643);
  and ginst297 (1916, 1628, 643);
  and ginst298 (1917, 1631, 643);
  and ginst299 (1918, 1634, 643);
  not ginst300 (1919, 1708);
  and ginst301 (1928, 1676, 693);
  and ginst302 (1929, 1681, 693);
  and ginst303 (1930, 1686, 693);
  and ginst304 (1931, 1690, 693);
  and ginst305 (1932, 1637, 699);
  and ginst306 (1933, 1642, 699);
  and ginst307 (1934, 1647, 699);
  and ginst308 (1935, 1651, 699);
  buf ginst309 (1936, 1600);
  nand ginst310 (1939, 1216, 1808);
  nand ginst311 (1940, 1585, 1810);
  nand ginst312 (1941, 1582, 1811);
  buf ginst313 (1942, 1676);
  buf ginst314 (1945, 1686);
  buf ginst315 (1948, 1681);
  buf ginst316 (1951, 1637);
  buf ginst317 (1954, 1690);
  buf ginst318 (1957, 1647);
  buf ginst319 (1960, 1642);
  buf ginst320 (1963, 1656);
  buf ginst321 (1966, 1651);
  or ginst322 (1969, 533, 1815);
  not ginst323 (1970, 1822);
  not ginst324 (1971, 1823);
  buf ginst325 (2010, 1848);
  buf ginst326 (2012, 1852);
  buf ginst327 (2014, 1856);
  buf ginst328 (2016, 1863);
  buf ginst329 (2018, 1870);
  buf ginst330 (2020, 1875);
  buf ginst331 (2022, 1880);
  not ginst332 (2028, 1778);
  not ginst333 (2029, 1781);
  nor ginst334 (2030, 1908, 1784);
  nor ginst335 (2031, 1909, 1785);
  and ginst336 (2032, 1506, 1502, 1778);
  and ginst337 (2033, 1773, 1770, 1781);
  or ginst338 (2034, 1571, 1935);
  not ginst339 (2040, 1801);
  not ginst340 (2041, 1804);
  and ginst341 (2042, 1557, 1553, 1801);
  and ginst342 (2043, 1798, 1795, 1804);
  nand ginst343 (2046, 1939, 1809);
  nand ginst344 (2049, 1940, 1941);
  or ginst345 (2052, 1544, 1910);
  or ginst346 (2055, 1545, 1911);
  or ginst347 (2058, 1546, 1912);
  or ginst348 (2061, 1547, 1913);
  or ginst349 (2064, 1548, 1914);
  or ginst350 (2067, 1549, 1915);
  or ginst351 (2070, 1550, 1916);
  or ginst352 (2073, 1551, 1917);
  or ginst353 (2076, 1552, 1918);
  or ginst354 (2079, 1564, 1928);
  or ginst355 (2095, 1565, 1929);
  or ginst356 (2098, 1566, 1930);
  or ginst357 (2101, 1567, 1931);
  or ginst358 (2104, 1568, 1932);
  or ginst359 (2107, 1569, 1933);
  or ginst360 (2110, 1570, 1934);
  and ginst361 (2113, 1897, 1894, 40);
  not ginst362 (2119, 1894);
  nand ginst363 (2120, 408, 1827);
  and ginst364 (2125, 1824, 537);
  and ginst365 (2126, 1852, 246);
  and ginst366 (2127, 1848, 537);
  not ginst367 (2128, 1848);
  not ginst368 (2135, 1852);
  not ginst369 (2141, 1863);
  not ginst370 (2144, 1870);
  not ginst371 (2147, 1875);
  not ginst372 (2150, 1880);
  and ginst373 (2153, 727, 1885);
  and ginst374 (2154, 1885, 1651);
  and ginst375 (2155, 730, 1888);
  and ginst376 (2156, 1888, 1656);
  and ginst377 (2157, 1770, 1506, 2028);
  and ginst378 (2158, 1502, 1773, 2029);
  not ginst379 (2171, 1942);
  nand ginst380 (2172, 1942, 1919);
  not ginst381 (2173, 1945);
  not ginst382 (2174, 1948);
  not ginst383 (2175, 1951);
  not ginst384 (2176, 1954);
  and ginst385 (2177, 1795, 1557, 2040);
  and ginst386 (2178, 1553, 1798, 2041);
  buf ginst387 (2185, 1836);
  buf ginst388 (2188, 1833);
  buf ginst389 (2191, 1841);
  not ginst390 (2194, 1856);
  not ginst391 (2197, 1827);
  not ginst392 (2200, 1936);
  buf ginst393 (2201, 1836);
  buf ginst394 (2204, 1833);
  buf ginst395 (2207, 1841);
  buf ginst396 (2210, 1824);
  buf ginst397 (2213, 1841);
  buf ginst398 (2216, 1841);
  nand ginst399 (2219, 2031, 2030);
  not ginst400 (2234, 1957);
  not ginst401 (2235, 1960);
  not ginst402 (2236, 1963);
  not ginst403 (2237, 1966);
  and ginst404 (2250, 40, 1897, 2119);
  or ginst405 (2266, 1831, 2126);
  or ginst406 (2269, 2127, 1832);
  or ginst407 (2291, 2153, 2154);
  or ginst408 (2294, 2155, 2156);
  nor ginst409 (2297, 2157, 2032);
  nor ginst410 (2298, 2158, 2033);
  not ginst411 (2300, 2046);
  not ginst412 (2301, 2049);
  nand ginst413 (2302, 2052, 1519);
  not ginst414 (2303, 2052);
  nand ginst415 (2304, 2055, 1520);
  not ginst416 (2305, 2055);
  nand ginst417 (2306, 2058, 1521);
  not ginst418 (2307, 2058);
  nand ginst419 (2308, 2061, 1522);
  not ginst420 (2309, 2061);
  nand ginst421 (2310, 2064, 1523);
  not ginst422 (2311, 2064);
  nand ginst423 (2312, 2067, 1524);
  not ginst424 (2313, 2067);
  nand ginst425 (2314, 2070, 1525);
  not ginst426 (2315, 2070);
  nand ginst427 (2316, 2073, 1526);
  not ginst428 (2317, 2073);
  nand ginst429 (2318, 2076, 1527);
  not ginst430 (2319, 2076);
  nand ginst431 (2320, 2079, 1528);
  not ginst432 (2321, 2079);
  nand ginst433 (2322, 1708, 2171);
  nand ginst434 (2323, 1948, 2173);
  nand ginst435 (2324, 1945, 2174);
  nand ginst436 (2325, 1954, 2175);
  nand ginst437 (2326, 1951, 2176);
  nor ginst438 (2327, 2177, 2042);
  nor ginst439 (2328, 2178, 2043);
  nand ginst440 (2329, 2095, 1572);
  not ginst441 (2330, 2095);
  nand ginst442 (2331, 2098, 1573);
  not ginst443 (2332, 2098);
  nand ginst444 (2333, 2101, 1574);
  not ginst445 (2334, 2101);
  nand ginst446 (2335, 2104, 1575);
  not ginst447 (2336, 2104);
  nand ginst448 (2337, 2107, 1576);
  not ginst449 (2338, 2107);
  nand ginst450 (2339, 2110, 1577);
  not ginst451 (2340, 2110);
  nand ginst452 (2354, 1960, 2234);
  nand ginst453 (2355, 1957, 2235);
  nand ginst454 (2356, 1966, 2236);
  nand ginst455 (2357, 1963, 2237);
  and ginst456 (2358, 2120, 533);
  not ginst457 (2359, 2113);
  not ginst458 (2364, 2185);
  not ginst459 (2365, 2188);
  not ginst460 (2366, 2191);
  not ginst461 (2367, 2194);
  buf ginst462 (2368, 2120);
  not ginst463 (2372, 2201);
  not ginst464 (2373, 2204);
  not ginst465 (2374, 2207);
  not ginst466 (2375, 2210);
  not ginst467 (2376, 2213);
  not ginst468 (2377, 2113);
  buf ginst469 (2382, 2113);
  and ginst470 (2386, 2120, 246);
  buf ginst471 (2387, 2266);
  buf ginst472 (2388, 2266);
  buf ginst473 (2389, 2269);
  buf ginst474 (2390, 2269);
  buf ginst475 (2391, 2113);
  not ginst476 (2395, 2113);
  nand ginst477 (2400, 2219, 2300);
  not ginst478 (2403, 2216);
  not ginst479 (2406, 2219);
  nand ginst480 (2407, 1219, 2303);
  nand ginst481 (2408, 1222, 2305);
  nand ginst482 (2409, 1225, 2307);
  nand ginst483 (2410, 1228, 2309);
  nand ginst484 (2411, 1231, 2311);
  nand ginst485 (2412, 1234, 2313);
  nand ginst486 (2413, 1237, 2315);
  nand ginst487 (2414, 1240, 2317);
  nand ginst488 (2415, 1243, 2319);
  nand ginst489 (2416, 1246, 2321);
  nand ginst490 (2417, 2322, 2172);
  nand ginst491 (2421, 2323, 2324);
  nand ginst492 (2425, 2325, 2326);
  nand ginst493 (2428, 1251, 2330);
  nand ginst494 (2429, 1254, 2332);
  nand ginst495 (2430, 1257, 2334);
  nand ginst496 (2431, 1260, 2336);
  nand ginst497 (2432, 1263, 2338);
  nand ginst498 (2433, 1266, 2340);
  buf ginst499 (2434, 2128);
  buf ginst500 (2437, 2135);
  buf ginst501 (2440, 2144);
  buf ginst502 (2443, 2141);
  buf ginst503 (2446, 2150);
  buf ginst504 (2449, 2147);
  not ginst505 (2452, 2197);
  nand ginst506 (2453, 2197, 2200);
  buf ginst507 (2454, 2128);
  buf ginst508 (2457, 2144);
  buf ginst509 (2460, 2141);
  buf ginst510 (2463, 2150);
  buf ginst511 (2466, 2147);
  not ginst512 (2469, 2120);
  buf ginst513 (2472, 2128);
  buf ginst514 (2475, 2135);
  buf ginst515 (2478, 2128);
  buf ginst516 (2481, 2135);
  nand ginst517 (2484, 2298, 2297);
  nand ginst518 (2487, 2356, 2357);
  nand ginst519 (2490, 2354, 2355);
  nand ginst520 (2493, 2328, 2327);
  or ginst521 (2496, 2358, 1814);
  nand ginst522 (2503, 2188, 2364);
  nand ginst523 (2504, 2185, 2365);
  nand ginst524 (2510, 2204, 2372);
  nand ginst525 (2511, 2201, 2373);
  or ginst526 (2521, 1830, 2386);
  nand ginst527 (2528, 2046, 2406);
  not ginst528 (2531, 2291);
  not ginst529 (2534, 2294);
  buf ginst530 (2537, 2250);
  buf ginst531 (2540, 2250);
  nand ginst532 (2544, 2302, 2407);
  nand ginst533 (2545, 2304, 2408);
  nand ginst534 (2546, 2306, 2409);
  nand ginst535 (2547, 2308, 2410);
  nand ginst536 (2548, 2310, 2411);
  nand ginst537 (2549, 2312, 2412);
  nand ginst538 (2550, 2314, 2413);
  nand ginst539 (2551, 2316, 2414);
  nand ginst540 (2552, 2318, 2415);
  nand ginst541 (2553, 2320, 2416);
  nand ginst542 (2563, 2329, 2428);
  nand ginst543 (2564, 2331, 2429);
  nand ginst544 (2565, 2333, 2430);
  nand ginst545 (2566, 2335, 2431);
  nand ginst546 (2567, 2337, 2432);
  nand ginst547 (2568, 2339, 2433);
  nand ginst548 (2579, 1936, 2452);
  buf ginst549 (2603, 2359);
  and ginst550 (2607, 1880, 2377);
  and ginst551 (2608, 1676, 2377);
  and ginst552 (2609, 1681, 2377);
  and ginst553 (2610, 1891, 2377);
  and ginst554 (2611, 1856, 2382);
  and ginst555 (2612, 1863, 2382);
  nand ginst556 (2613, 2503, 2504);
  not ginst557 (2617, 2434);
  nand ginst558 (2618, 2434, 2366);
  nand ginst559 (2619, 2437, 2367);
  not ginst560 (2620, 2437);
  not ginst561 (2621, 2368);
  nand ginst562 (2624, 2510, 2511);
  not ginst563 (2628, 2454);
  nand ginst564 (2629, 2454, 2374);
  not ginst565 (2630, 2472);
  and ginst566 (2631, 1856, 2391);
  and ginst567 (2632, 1863, 2391);
  and ginst568 (2633, 1880, 2395);
  and ginst569 (2634, 1676, 2395);
  and ginst570 (2635, 1681, 2395);
  and ginst571 (2636, 1891, 2395);
  not ginst572 (2638, 2382);
  buf ginst573 (2643, 2521);
  buf ginst574 (2644, 2521);
  not ginst575 (2645, 2475);
  not ginst576 (2646, 2391);
  nand ginst577 (2652, 2528, 2400);
  not ginst578 (2655, 2478);
  not ginst579 (2656, 2481);
  buf ginst580 (2659, 2359);
  not ginst581 (2663, 2484);
  nand ginst582 (2664, 2484, 2301);
  not ginst583 (2665, 2553);
  not ginst584 (2666, 2552);
  not ginst585 (2667, 2551);
  not ginst586 (2668, 2550);
  not ginst587 (2669, 2549);
  not ginst588 (2670, 2548);
  not ginst589 (2671, 2547);
  not ginst590 (2672, 2546);
  not ginst591 (2673, 2545);
  not ginst592 (2674, 2544);
  not ginst593 (2675, 2568);
  not ginst594 (2676, 2567);
  not ginst595 (2677, 2566);
  not ginst596 (2678, 2565);
  not ginst597 (2679, 2564);
  not ginst598 (2680, 2563);
  not ginst599 (2681, 2417);
  not ginst600 (2684, 2421);
  buf ginst601 (2687, 2425);
  buf ginst602 (2690, 2425);
  not ginst603 (2693, 2493);
  nand ginst604 (2694, 2493, 1807);
  not ginst605 (2695, 2440);
  not ginst606 (2696, 2443);
  not ginst607 (2697, 2446);
  not ginst608 (2698, 2449);
  not ginst609 (2699, 2457);
  not ginst610 (2700, 2460);
  not ginst611 (2701, 2463);
  not ginst612 (2702, 2466);
  nand ginst613 (2703, 2579, 2453);
  not ginst614 (2706, 2469);
  not ginst615 (2707, 2487);
  not ginst616 (2708, 2490);
  and ginst617 (2709, 2294, 2534);
  and ginst618 (2710, 2291, 2531);
  nand ginst619 (2719, 2191, 2617);
  nand ginst620 (2720, 2194, 2620);
  nand ginst621 (2726, 2207, 2628);
  buf ginst622 (2729, 2537);
  buf ginst623 (2738, 2537);
  not ginst624 (2743, 2652);
  nand ginst625 (2747, 2049, 2663);
  and ginst626 (2748, 2665, 2666, 2667, 2668, 2669);
  and ginst627 (2749, 2670, 2671, 2672, 2673, 2674);
  and ginst628 (2750, 2034, 2675);
  and ginst629 (2751, 2676, 2677, 2678, 2679, 2680);
  nand ginst630 (2760, 1588, 2693);
  buf ginst631 (2761, 2540);
  buf ginst632 (2766, 2540);
  nand ginst633 (2771, 2443, 2695);
  nand ginst634 (2772, 2440, 2696);
  nand ginst635 (2773, 2449, 2697);
  nand ginst636 (2774, 2446, 2698);
  nand ginst637 (2775, 2460, 2699);
  nand ginst638 (2776, 2457, 2700);
  nand ginst639 (2777, 2466, 2701);
  nand ginst640 (2778, 2463, 2702);
  nand ginst641 (2781, 2490, 2707);
  nand ginst642 (2782, 2487, 2708);
  or ginst643 (2783, 2709, 2534);
  or ginst644 (2784, 2710, 2531);
  and ginst645 (2789, 1856, 2638);
  and ginst646 (2790, 1863, 2638);
  and ginst647 (2791, 1870, 2638);
  and ginst648 (2792, 1875, 2638);
  not ginst649 (2793, 2613);
  nand ginst650 (2796, 2719, 2618);
  nand ginst651 (2800, 2619, 2720);
  not ginst652 (2803, 2624);
  nand ginst653 (2806, 2726, 2629);
  and ginst654 (2809, 1856, 2646);
  and ginst655 (2810, 1863, 2646);
  and ginst656 (2811, 1870, 2646);
  and ginst657 (2812, 1875, 2646);
  and ginst658 (2817, 2743, 14);
  buf ginst659 (2820, 2603);
  nand ginst660 (2826, 2747, 2664);
  and ginst661 (2829, 2748, 2749);
  and ginst662 (2830, 2750, 2751);
  buf ginst663 (2831, 2659);
  not ginst664 (2837, 2687);
  not ginst665 (2838, 2690);
  and ginst666 (2839, 2421, 2417, 2687);
  and ginst667 (2840, 2684, 2681, 2690);
  nand ginst668 (2841, 2760, 2694);
  buf ginst669 (2844, 2603);
  buf ginst670 (2854, 2603);
  buf ginst671 (2859, 2659);
  buf ginst672 (2869, 2659);
  nand ginst673 (2874, 2773, 2774);
  nand ginst674 (2877, 2771, 2772);
  not ginst675 (2880, 2703);
  nand ginst676 (2881, 2703, 2706);
  nand ginst677 (2882, 2777, 2778);
  nand ginst678 (2885, 2775, 2776);
  nand ginst679 (2888, 2781, 2782);
  nand ginst680 (2891, 2783, 2784);
  and ginst681 (2894, 2607, 2729);
  and ginst682 (2895, 2608, 2729);
  and ginst683 (2896, 2609, 2729);
  and ginst684 (2897, 2610, 2729);
  or ginst685 (2898, 2789, 2611);
  or ginst686 (2899, 2790, 2612);
  and ginst687 (2900, 2791, 1037);
  and ginst688 (2901, 2792, 1037);
  or ginst689 (2914, 2809, 2631);
  or ginst690 (2915, 2810, 2632);
  and ginst691 (2916, 2811, 1070);
  and ginst692 (2917, 2812, 1070);
  and ginst693 (2918, 2633, 2738);
  and ginst694 (2919, 2634, 2738);
  and ginst695 (2920, 2635, 2738);
  and ginst696 (2921, 2636, 2738);
  buf ginst697 (2925, 2817);
  and ginst698 (2931, 2829, 2830, 1302);
  and ginst699 (2938, 2681, 2421, 2837);
  and ginst700 (2939, 2417, 2684, 2838);
  nand ginst701 (2963, 2469, 2880);
  not ginst702 (2970, 2841);
  not ginst703 (2971, 2826);
  not ginst704 (2972, 2894);
  not ginst705 (2975, 2895);
  not ginst706 (2978, 2896);
  not ginst707 (2981, 2897);
  and ginst708 (2984, 2898, 1037);
  and ginst709 (2985, 2899, 1037);
  not ginst710 (2986, 2900);
  not ginst711 (2989, 2901);
  not ginst712 (2992, 2796);
  buf ginst713 (2995, 2800);
  buf ginst714 (2998, 2800);
  buf ginst715 (3001, 2806);
  buf ginst716 (3004, 2806);
  and ginst717 (3007, 574, 2820);
  and ginst718 (3008, 2914, 1070);
  and ginst719 (3009, 2915, 1070);
  not ginst720 (3010, 2916);
  not ginst721 (3013, 2917);
  not ginst722 (3016, 2918);
  not ginst723 (3019, 2919);
  not ginst724 (3022, 2920);
  not ginst725 (3025, 2921);
  not ginst726 (3028, 2817);
  and ginst727 (3029, 574, 2831);
  not ginst728 (3030, 2820);
  and ginst729 (3035, 578, 2820);
  and ginst730 (3036, 655, 2820);
  and ginst731 (3037, 659, 2820);
  buf ginst732 (3038, 2931);
  not ginst733 (3039, 2831);
  and ginst734 (3044, 578, 2831);
  and ginst735 (3045, 655, 2831);
  and ginst736 (3046, 659, 2831);
  nor ginst737 (3047, 2938, 2839);
  nor ginst738 (3048, 2939, 2840);
  not ginst739 (3049, 2888);
  not ginst740 (3050, 2844);
  and ginst741 (3053, 663, 2844);
  and ginst742 (3054, 667, 2844);
  and ginst743 (3055, 671, 2844);
  and ginst744 (3056, 675, 2844);
  and ginst745 (3057, 679, 2854);
  and ginst746 (3058, 683, 2854);
  and ginst747 (3059, 687, 2854);
  and ginst748 (3060, 705, 2854);
  not ginst749 (3061, 2859);
  and ginst750 (3064, 663, 2859);
  and ginst751 (3065, 667, 2859);
  and ginst752 (3066, 671, 2859);
  and ginst753 (3067, 675, 2859);
  and ginst754 (3068, 679, 2869);
  and ginst755 (3069, 683, 2869);
  and ginst756 (3070, 687, 2869);
  and ginst757 (3071, 705, 2869);
  not ginst758 (3072, 2874);
  not ginst759 (3073, 2877);
  not ginst760 (3074, 2882);
  not ginst761 (3075, 2885);
  nand ginst762 (3076, 2881, 2963);
  not ginst763 (3079, 2931);
  not ginst764 (3088, 2984);
  not ginst765 (3091, 2985);
  not ginst766 (3110, 3008);
  not ginst767 (3113, 3009);
  and ginst768 (3137, 3055, 1190);
  and ginst769 (3140, 3056, 1190);
  and ginst770 (3143, 3057, 2761);
  and ginst771 (3146, 3058, 2761);
  and ginst772 (3149, 3059, 2761);
  and ginst773 (3152, 3060, 2761);
  and ginst774 (3157, 3066, 1195);
  and ginst775 (3160, 3067, 1195);
  and ginst776 (3163, 3068, 2766);
  and ginst777 (3166, 3069, 2766);
  and ginst778 (3169, 3070, 2766);
  and ginst779 (3172, 3071, 2766);
  nand ginst780 (3175, 2877, 3072);
  nand ginst781 (3176, 2874, 3073);
  nand ginst782 (3177, 2885, 3074);
  nand ginst783 (3178, 2882, 3075);
  nand ginst784 (3180, 3048, 3047);
  not ginst785 (3187, 2995);
  not ginst786 (3188, 2998);
  not ginst787 (3189, 3001);
  not ginst788 (3190, 3004);
  and ginst789 (3191, 2796, 2613, 2995);
  and ginst790 (3192, 2992, 2793, 2998);
  and ginst791 (3193, 2624, 2368, 3001);
  and ginst792 (3194, 2803, 2621, 3004);
  nand ginst793 (3195, 3076, 2375);
  not ginst794 (3196, 3076);
  and ginst795 (3197, 687, 3030);
  and ginst796 (3208, 687, 3039);
  and ginst797 (3215, 705, 3030);
  and ginst798 (3216, 711, 3030);
  and ginst799 (3217, 715, 3030);
  and ginst800 (3218, 705, 3039);
  and ginst801 (3219, 711, 3039);
  and ginst802 (3220, 715, 3039);
  and ginst803 (3222, 719, 3050);
  and ginst804 (3223, 723, 3050);
  and ginst805 (3230, 719, 3061);
  and ginst806 (3231, 723, 3061);
  nand ginst807 (3238, 3175, 3176);
  nand ginst808 (3241, 3177, 3178);
  buf ginst809 (3244, 2981);
  buf ginst810 (3247, 2978);
  buf ginst811 (3250, 2975);
  buf ginst812 (3253, 2972);
  buf ginst813 (3256, 2989);
  buf ginst814 (3259, 2986);
  buf ginst815 (3262, 3025);
  buf ginst816 (3265, 3022);
  buf ginst817 (3268, 3019);
  buf ginst818 (3271, 3016);
  buf ginst819 (3274, 3013);
  buf ginst820 (3277, 3010);
  and ginst821 (3281, 2793, 2796, 3187);
  and ginst822 (3282, 2613, 2992, 3188);
  and ginst823 (3283, 2621, 2624, 3189);
  and ginst824 (3284, 2368, 2803, 3190);
  nand ginst825 (3286, 2210, 3196);
  or ginst826 (3288, 3197, 3007);
  nand ginst827 (3289, 3180, 3049);
  and ginst828 (3291, 3152, 2981);
  and ginst829 (3293, 3149, 2978);
  and ginst830 (3295, 3146, 2975);
  and ginst831 (3296, 2972, 3143);
  and ginst832 (3299, 3140, 2989);
  and ginst833 (3301, 3137, 2986);
  or ginst834 (3302, 3208, 3029);
  and ginst835 (3304, 3172, 3025);
  and ginst836 (3306, 3169, 3022);
  and ginst837 (3308, 3166, 3019);
  and ginst838 (3309, 3016, 3163);
  and ginst839 (3312, 3160, 3013);
  and ginst840 (3314, 3157, 3010);
  or ginst841 (3315, 3215, 3035);
  or ginst842 (3318, 3216, 3036);
  or ginst843 (3321, 3217, 3037);
  or ginst844 (3324, 3218, 3044);
  or ginst845 (3327, 3219, 3045);
  or ginst846 (3330, 3220, 3046);
  not ginst847 (3333, 3180);
  or ginst848 (3334, 3222, 3053);
  or ginst849 (3335, 3223, 3054);
  or ginst850 (3336, 3230, 3064);
  or ginst851 (3337, 3231, 3065);
  buf ginst852 (3340, 3152);
  buf ginst853 (3344, 3149);
  buf ginst854 (3348, 3146);
  buf ginst855 (3352, 3143);
  buf ginst856 (3356, 3140);
  buf ginst857 (3360, 3137);
  buf ginst858 (3364, 3091);
  buf ginst859 (3367, 3088);
  buf ginst860 (3370, 3172);
  buf ginst861 (3374, 3169);
  buf ginst862 (3378, 3166);
  buf ginst863 (3382, 3163);
  buf ginst864 (3386, 3160);
  buf ginst865 (3390, 3157);
  buf ginst866 (3394, 3113);
  buf ginst867 (3397, 3110);
  nand ginst868 (3400, 3195, 3286);
  nor ginst869 (3401, 3281, 3191);
  nor ginst870 (3402, 3282, 3192);
  nor ginst871 (3403, 3283, 3193);
  nor ginst872 (3404, 3284, 3194);
  not ginst873 (3405, 3238);
  not ginst874 (3406, 3241);
  and ginst875 (3409, 3288, 1836);
  nand ginst876 (3410, 2888, 3333);
  not ginst877 (3412, 3244);
  not ginst878 (3414, 3247);
  not ginst879 (3416, 3250);
  not ginst880 (3418, 3253);
  not ginst881 (3420, 3256);
  not ginst882 (3422, 3259);
  and ginst883 (3428, 3302, 1836);
  not ginst884 (3430, 3262);
  not ginst885 (3432, 3265);
  not ginst886 (3434, 3268);
  not ginst887 (3436, 3271);
  not ginst888 (3438, 3274);
  not ginst889 (3440, 3277);
  and ginst890 (3450, 3334, 1190);
  and ginst891 (3453, 3335, 1190);
  and ginst892 (3456, 3336, 1195);
  and ginst893 (3459, 3337, 1195);
  and ginst894 (3478, 3400, 533);
  and ginst895 (3479, 3318, 2128);
  and ginst896 (3480, 3315, 1841);
  nand ginst897 (3481, 3410, 3289);
  not ginst898 (3482, 3340);
  nand ginst899 (3483, 3340, 3412);
  not ginst900 (3484, 3344);
  nand ginst901 (3485, 3344, 3414);
  not ginst902 (3486, 3348);
  nand ginst903 (3487, 3348, 3416);
  not ginst904 (3488, 3352);
  nand ginst905 (3489, 3352, 3418);
  not ginst906 (3490, 3356);
  nand ginst907 (3491, 3356, 3420);
  not ginst908 (3492, 3360);
  nand ginst909 (3493, 3360, 3422);
  not ginst910 (3494, 3364);
  not ginst911 (3496, 3367);
  and ginst912 (3498, 3321, 2135);
  and ginst913 (3499, 3327, 2128);
  and ginst914 (3500, 3324, 1841);
  not ginst915 (3501, 3370);
  nand ginst916 (3502, 3370, 3430);
  not ginst917 (3503, 3374);
  nand ginst918 (3504, 3374, 3432);
  not ginst919 (3505, 3378);
  nand ginst920 (3506, 3378, 3434);
  not ginst921 (3507, 3382);
  nand ginst922 (3508, 3382, 3436);
  not ginst923 (3509, 3386);
  nand ginst924 (3510, 3386, 3438);
  not ginst925 (3511, 3390);
  nand ginst926 (3512, 3390, 3440);
  not ginst927 (3513, 3394);
  not ginst928 (3515, 3397);
  and ginst929 (3517, 3330, 2135);
  nand ginst930 (3522, 3402, 3401);
  nand ginst931 (3525, 3404, 3403);
  buf ginst932 (3528, 3318);
  buf ginst933 (3531, 3315);
  buf ginst934 (3534, 3321);
  buf ginst935 (3537, 3327);
  buf ginst936 (3540, 3324);
  buf ginst937 (3543, 3330);
  or ginst938 (3546, 3478, 1813);
  not ginst939 (3551, 3481);
  nand ginst940 (3552, 3244, 3482);
  nand ginst941 (3553, 3247, 3484);
  nand ginst942 (3554, 3250, 3486);
  nand ginst943 (3555, 3253, 3488);
  nand ginst944 (3556, 3256, 3490);
  nand ginst945 (3557, 3259, 3492);
  and ginst946 (3558, 3453, 3091);
  and ginst947 (3559, 3450, 3088);
  nand ginst948 (3563, 3262, 3501);
  nand ginst949 (3564, 3265, 3503);
  nand ginst950 (3565, 3268, 3505);
  nand ginst951 (3566, 3271, 3507);
  nand ginst952 (3567, 3274, 3509);
  nand ginst953 (3568, 3277, 3511);
  and ginst954 (3569, 3459, 3113);
  and ginst955 (3570, 3456, 3110);
  buf ginst956 (3576, 3453);
  buf ginst957 (3579, 3450);
  buf ginst958 (3585, 3459);
  buf ginst959 (3588, 3456);
  not ginst960 (3592, 3522);
  nand ginst961 (3593, 3522, 3405);
  not ginst962 (3594, 3525);
  nand ginst963 (3595, 3525, 3406);
  not ginst964 (3596, 3528);
  nand ginst965 (3597, 3528, 2630);
  nand ginst966 (3598, 3531, 2376);
  not ginst967 (3599, 3531);
  and ginst968 (3600, 3551, 800);
  nand ginst969 (3603, 3552, 3483);
  nand ginst970 (3608, 3553, 3485);
  nand ginst971 (3612, 3554, 3487);
  nand ginst972 (3615, 3555, 3489);
  nand ginst973 (3616, 3556, 3491);
  nand ginst974 (3622, 3557, 3493);
  not ginst975 (3629, 3534);
  nand ginst976 (3630, 3534, 2645);
  not ginst977 (3631, 3537);
  nand ginst978 (3632, 3537, 2655);
  nand ginst979 (3633, 3540, 2403);
  not ginst980 (3634, 3540);
  nand ginst981 (3635, 3563, 3502);
  nand ginst982 (3640, 3564, 3504);
  nand ginst983 (3644, 3565, 3506);
  nand ginst984 (3647, 3566, 3508);
  nand ginst985 (3648, 3567, 3510);
  nand ginst986 (3654, 3568, 3512);
  not ginst987 (3661, 3543);
  nand ginst988 (3662, 3543, 2656);
  nand ginst989 (3667, 3238, 3592);
  nand ginst990 (3668, 3241, 3594);
  nand ginst991 (3669, 2472, 3596);
  nand ginst992 (3670, 2213, 3599);
  buf ginst993 (3671, 3600);
  not ginst994 (3691, 3576);
  nand ginst995 (3692, 3576, 3494);
  not ginst996 (3693, 3579);
  nand ginst997 (3694, 3579, 3496);
  nand ginst998 (3695, 2475, 3629);
  nand ginst999 (3696, 2478, 3631);
  nand ginst1000 (3697, 2216, 3634);
  not ginst1001 (3716, 3585);
  nand ginst1002 (3717, 3585, 3513);
  not ginst1003 (3718, 3588);
  nand ginst1004 (3719, 3588, 3515);
  nand ginst1005 (3720, 2481, 3661);
  nand ginst1006 (3721, 3667, 3593);
  nand ginst1007 (3722, 3668, 3595);
  nand ginst1008 (3723, 3669, 3597);
  nand ginst1009 (3726, 3670, 3598);
  not ginst1010 (3727, 3600);
  nand ginst1011 (3728, 3364, 3691);
  nand ginst1012 (3729, 3367, 3693);
  nand ginst1013 (3730, 3695, 3630);
  and ginst1014 (3731, 3608, 3615, 3612, 3603);
  and ginst1015 (3732, 3603, 3293);
  and ginst1016 (3733, 3608, 3603, 3295);
  and ginst1017 (3734, 3612, 3603, 3296, 3608);
  and ginst1018 (3735, 3616, 3301);
  and ginst1019 (3736, 3622, 3616, 3558);
  nand ginst1020 (3737, 3696, 3632);
  nand ginst1021 (3740, 3697, 3633);
  nand ginst1022 (3741, 3394, 3716);
  nand ginst1023 (3742, 3397, 3718);
  nand ginst1024 (3743, 3720, 3662);
  and ginst1025 (3744, 3640, 3647, 3644, 3635);
  and ginst1026 (3745, 3635, 3306);
  and ginst1027 (3746, 3640, 3635, 3308);
  and ginst1028 (3747, 3644, 3635, 3309, 3640);
  and ginst1029 (3748, 3648, 3314);
  and ginst1030 (3749, 3654, 3648, 3569);
  not ginst1031 (3750, 3721);
  and ginst1032 (3753, 3722, 246);
  nand ginst1033 (3754, 3728, 3692);
  nand ginst1034 (3758, 3729, 3694);
  not ginst1035 (3761, 3731);
  or ginst1036 (3762, 3291, 3732, 3733, 3734);
  nand ginst1037 (3767, 3741, 3717);
  nand ginst1038 (3771, 3742, 3719);
  not ginst1039 (3774, 3744);
  or ginst1040 (3775, 3304, 3745, 3746, 3747);
  and ginst1041 (3778, 3723, 3480);
  and ginst1042 (3779, 3726, 3723, 3409);
  or ginst1043 (3780, 2125, 3753);
  and ginst1044 (3790, 3750, 800);
  and ginst1045 (3793, 3737, 3500);
  and ginst1046 (3794, 3740, 3737, 3428);
  or ginst1047 (3802, 3479, 3778, 3779);
  buf ginst1048 (3803, 3780);
  buf ginst1049 (3804, 3780);
  not ginst1050 (3805, 3762);
  and ginst1051 (3806, 3622, 3730, 3754, 3616, 3758);
  and ginst1052 (3807, 3754, 3616, 3559, 3622);
  and ginst1053 (3808, 3758, 3754, 3616, 3498, 3622);
  buf ginst1054 (3809, 3790);
  or ginst1055 (3811, 3499, 3793, 3794);
  not ginst1056 (3812, 3775);
  and ginst1057 (3813, 3654, 3743, 3767, 3648, 3771);
  and ginst1058 (3814, 3767, 3648, 3570, 3654);
  and ginst1059 (3815, 3771, 3767, 3648, 3517, 3654);
  or ginst1060 (3816, 3299, 3735, 3736, 3807, 3808);
  and ginst1061 (3817, 3806, 3802);
  nand ginst1062 (3818, 3805, 3761);
  not ginst1063 (3819, 3790);
  or ginst1064 (3820, 3312, 3748, 3749, 3814, 3815);
  and ginst1065 (3821, 3813, 3811);
  nand ginst1066 (3822, 3812, 3774);
  or ginst1067 (3823, 3816, 3817);
  and ginst1068 (3826, 3727, 3819, 2841);
  or ginst1069 (3827, 3820, 3821);
  not ginst1070 (3834, 3823);
  and ginst1071 (3835, 3818, 3823);
  not ginst1072 (3836, 3827);
  and ginst1073 (3837, 3822, 3827);
  and ginst1074 (3838, 3762, 3834);
  and ginst1075 (3839, 3775, 3836);
  or ginst1076 (3840, 3838, 3835);
  or ginst1077 (3843, 3839, 3837);
  buf ginst1078 (3851, 3843);
  nand ginst1079 (3852, 3843, 3840);
  and ginst1080 (3857, 3843, 3852);
  and ginst1081 (3858, 3852, 3840);
  or ginst1082 (3859, 3857, 3858);
  not ginst1083 (3864, 3859);
  and ginst1084 (3869, 3859, 3864);
  or ginst1085 (3870, 3869, 3864);
  not ginst1086 (3875, 3870);
  and ginst1087 (3876, 2826, 3028, 3870);
  and ginst1088 (3877, 3826, 3876, 1591);
  buf ginst1089 (3881, 3877);
  not ginst1090 (3882, 3877);
  buf ginst1091 (398, 219);
  buf ginst1092 (400, 219);
  buf ginst1093 (401, 219);
  and ginst1094 (405, 1, 3);
  not ginst1095 (408, 230);
  buf ginst1096 (419, 253);
  buf ginst1097 (420, 253);
  not ginst1098 (425, 262);
  buf ginst1099 (456, 290);
  buf ginst1100 (457, 290);
  buf ginst1101 (458, 290);
  and ginst1102 (485, 309, 305, 301, 297);
  not ginst1103 (486, 405);
  not ginst1104 (487, 44);
  not ginst1105 (488, 132);
  not ginst1106 (489, 82);
  not ginst1107 (490, 96);
  not ginst1108 (491, 69);
  not ginst1109 (492, 120);
  not ginst1110 (493, 57);
  not ginst1111 (494, 108);
  and ginst1112 (495, 2, 15, 237);
  buf ginst1113 (496, 237);
  and ginst1114 (499, 37, 37);
  buf ginst1115 (500, 219);
  buf ginst1116 (503, 8);
  buf ginst1117 (506, 8);
  buf ginst1118 (509, 227);
  buf ginst1119 (521, 234);
  not ginst1120 (533, 241);
  not ginst1121 (537, 246);
  and ginst1122 (543, 11, 246);
  and ginst1123 (544, 132, 82, 96, 44);
  and ginst1124 (547, 120, 57, 108, 69);
  buf ginst1125 (550, 227);
  buf ginst1126 (562, 234);
  not ginst1127 (574, 256);
  not ginst1128 (578, 259);
  buf ginst1129 (582, 319);
  buf ginst1130 (594, 322);
  not ginst1131 (606, 328);
  not ginst1132 (607, 331);
  not ginst1133 (608, 334);
  not ginst1134 (609, 337);
  not ginst1135 (610, 340);
  not ginst1136 (611, 343);
  not ginst1137 (612, 352);
  buf ginst1138 (613, 319);
  buf ginst1139 (625, 322);
  buf ginst1140 (637, 16);
  buf ginst1141 (643, 16);
  not ginst1142 (650, 355);
  and ginst1143 (651, 7, 237);
  not ginst1144 (655, 263);
  not ginst1145 (659, 266);
  not ginst1146 (663, 269);
  not ginst1147 (667, 272);
  not ginst1148 (671, 275);
  not ginst1149 (675, 278);
  not ginst1150 (679, 281);
  not ginst1151 (683, 284);
  not ginst1152 (687, 287);
  buf ginst1153 (693, 29);
  buf ginst1154 (699, 29);
  not ginst1155 (705, 294);
  not ginst1156 (711, 297);
  not ginst1157 (715, 301);
  not ginst1158 (719, 305);
  not ginst1159 (723, 309);
  not ginst1160 (727, 313);
  not ginst1161 (730, 316);
  not ginst1162 (733, 346);
  not ginst1163 (734, 349);
  buf ginst1164 (735, 259);
  buf ginst1165 (738, 256);
  buf ginst1166 (741, 263);
  buf ginst1167 (744, 269);
  buf ginst1168 (747, 266);
  buf ginst1169 (750, 275);
  buf ginst1170 (753, 272);
  buf ginst1171 (756, 281);
  buf ginst1172 (759, 278);
  buf ginst1173 (762, 287);
  buf ginst1174 (765, 284);
  buf ginst1175 (768, 294);
  buf ginst1176 (771, 301);
  buf ginst1177 (774, 297);
  buf ginst1178 (777, 309);
  buf ginst1179 (780, 305);
  buf ginst1180 (783, 316);
  buf ginst1181 (786, 313);
  not ginst1182 (792, 485);
  not ginst1183 (799, 495);
  not ginst1184 (800, 499);
  buf ginst1185 (805, 500);
  nand ginst1186 (900, 331, 606);
  nand ginst1187 (901, 328, 607);
  nand ginst1188 (902, 337, 608);
  nand ginst1189 (903, 334, 609);
  nand ginst1190 (904, 343, 610);
  nand ginst1191 (905, 340, 611);
  nand ginst1192 (998, 349, 733);
  nand ginst1193 (999, 346, 734);

endmodule
