// Main module
module temp(N1, N2, N3, N4);

  input N1, N2;
  output N3, N4;
  wire ;

  buf ginst1 (N3, N1);
  not ginst2 (N4, N2);

endmodule
