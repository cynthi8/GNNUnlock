/*************** Top Level ***************/
module c2670_AntiSAT_8_0_top (N145, N153, N162, N168, N172, N210, N190, N212, N167, N185, N173, N174, N183, N196, N151, N200, N187, N195, N155, N193, N146, N163, N178, N211, N208, N177, N182, N213, N191, N216, N204, N170, N165, N179, N189, N207, N184, N148, N154, N157, N158, N164, N149, N180, N192, N156, N194, N203, N199, N171, N205, N161, N160, N176, N197, N209, N201, N202, N188, N218, N143, N175, N169, N166, N186, N159, N217, N147, N144, N181, N150, N215, N206, N198, N152, N214, N1, N2, N3, N4, N5, N6, N7, N8, N11, N14, N15, N16, N19, N20, N21, N22, N23, N24, N25, N26, N27, N28, N29, N32, N33, N34, N35, N36, N37, N40, N43, N44, N47, N48, N49, N50, N51, N52, N53, N54, N55, N56, N57, N60, N61, N62, N63, N64, N65, N66, N67, N68, N69, N72, N73, N74, N75, N76, N77, N78, N79, N80, N81, N82, N85, N86, N87, N88, N89, N90, N91, N92, N93, N94, N95, N96, N99, N100, N101, N102, N103, N104, N105, N106, N107, N108, N111, N112, N113, N114, N115, N116, N117, N118, N119, N120, N123, N124, N125, N126, N127, N128, N129, N130, N131, N132, N135, N136, N137, N138, N139, N140, N141, N142, N219, N224, N227, N230, N231, N234, N237, N241, N246, N253, N256, N259, N262, N263, N266, N269, N272, N275, N278, N281, N284, N287, N290, N294, N297, N301, N305, N309, N313, N316, N319, N322, N325, N328, N331, N334, N337, N340, N343, N346, N349, N352, N355, keyinput0, keyinput1, keyinput2, keyinput3, keyinput4, keyinput5, keyinput6, keyinput7, N2016, N3803, N214_BUFF, N217_BUFF, N160_BUFF, N2496, N2022, N173_BUFF, N3809, N213_BUFF, N190_BUFF, N799, N215_BUFF, N183_BUFF, N164_BUFF, N1269, N3851, N192_BUFF, N218_BUFF, N2925, N188_BUFF, N1726, N148_BUFF, N1448, N159_BUFF, N494, N2644, N1026, N2014, N158_BUFF, N2389, N492, N152_BUFF, N162_BUFF, N167_BUFF, N199_BUFF, N145_BUFF, N144_BUFF, N489, N1816, N1969, N458, N206_BUFF, N1029, N2012, N202_BUFF, N156_BUFF, N210_BUFF, N488, N2018, N3038, N487, N2390, N1970, N208_BUFF, N2643, N401, N490, N197_BUFF, N194_BUFF, N189_BUFF, N491, N155_BUFF, N1028, N151_BUFF, N186_BUFF, N3079, N198_BUFF, N398, N178_BUFF, N212_BUFF, N1818, N203_BUFF, N182_BUFF, N196_BUFF, N419, N143_BUFF, N201_BUFF, N193_BUFF, N187_BUFF, N161_BUFF, N1819, N3882, N170_BUFF, N792, N166_BUFF, N1817, N157_BUFF, N456, N2388, N195_BUFF, N3881, N805, N154_BUFF, N176_BUFF, N169_BUFF, N205_BUFF, N184_BUFF, N179_BUFF, N3804, N146_BUFF, N1820, N200_BUFF, N149_BUFF, N3875, N150_BUFF, N153_BUFF, N204_BUFF, N2387, N400, N191_BUFF, N207_BUFF, N420, N163_BUFF, N2970, N172_BUFF, N180_BUFF, N2971, N2010, N177_BUFF, N209_BUFF, N174_BUFF, N2891, N147_BUFF, N165_BUFF, N457, N185_BUFF, N3671, N211_BUFF, N171_BUFF, N168_BUFF, N2020, N216_BUFF, N1277, N1821, N3546, N175_BUFF, N493, N1971, N181_BUFF);

  input N145, N153, N162, N168, N172, N210, N190, N212, N167, N185, N173, N174, N183, N196, N151, N200, N187, N195, N155, N193, N146, N163, N178, N211, N208, N177, N182, N213, N191, N216, N204, N170, N165, N179, N189, N207, N184, N148, N154, N157, N158, N164, N149, N180, N192, N156, N194, N203, N199, N171, N205, N161, N160, N176, N197, N209, N201, N202, N188, N218, N143, N175, N169, N166, N186, N159, N217, N147, N144, N181, N150, N215, N206, N198, N152, N214, N1, N2, N3, N4, N5, N6, N7, N8, N11, N14, N15, N16, N19, N20, N21, N22, N23, N24, N25, N26, N27, N28, N29, N32, N33, N34, N35, N36, N37, N40, N43, N44, N47, N48, N49, N50, N51, N52, N53, N54, N55, N56, N57, N60, N61, N62, N63, N64, N65, N66, N67, N68, N69, N72, N73, N74, N75, N76, N77, N78, N79, N80, N81, N82, N85, N86, N87, N88, N89, N90, N91, N92, N93, N94, N95, N96, N99, N100, N101, N102, N103, N104, N105, N106, N107, N108, N111, N112, N113, N114, N115, N116, N117, N118, N119, N120, N123, N124, N125, N126, N127, N128, N129, N130, N131, N132, N135, N136, N137, N138, N139, N140, N141, N142, N219, N224, N227, N230, N231, N234, N237, N241, N246, N253, N256, N259, N262, N263, N266, N269, N272, N275, N278, N281, N284, N287, N290, N294, N297, N301, N305, N309, N313, N316, N319, N322, N325, N328, N331, N334, N337, N340, N343, N346, N349, N352, N355, keyinput0, keyinput1, keyinput2, keyinput3, keyinput4, keyinput5, keyinput6, keyinput7;
  output N2016, N3803, N214_BUFF, N217_BUFF, N160_BUFF, N2496, N2022, N173_BUFF, N3809, N213_BUFF, N190_BUFF, N799, N215_BUFF, N183_BUFF, N164_BUFF, N1269, N3851, N192_BUFF, N218_BUFF, N2925, N188_BUFF, N1726, N148_BUFF, N1448, N159_BUFF, N494, N2644, N1026, N2014, N158_BUFF, N2389, N492, N152_BUFF, N162_BUFF, N167_BUFF, N199_BUFF, N145_BUFF, N144_BUFF, N489, N1816, N1969, N458, N206_BUFF, N1029, N2012, N202_BUFF, N156_BUFF, N210_BUFF, N488, N2018, N3038, N487, N2390, N1970, N208_BUFF, N2643, N401, N490, N197_BUFF, N194_BUFF, N189_BUFF, N491, N155_BUFF, N1028, N151_BUFF, N186_BUFF, N3079, N198_BUFF, N398, N178_BUFF, N212_BUFF, N1818, N203_BUFF, N182_BUFF, N196_BUFF, N419, N143_BUFF, N201_BUFF, N193_BUFF, N187_BUFF, N161_BUFF, N1819, N3882, N170_BUFF, N792, N166_BUFF, N1817, N157_BUFF, N456, N2388, N195_BUFF, N3881, N805, N154_BUFF, N176_BUFF, N169_BUFF, N205_BUFF, N184_BUFF, N179_BUFF, N3804, N146_BUFF, N1820, N200_BUFF, N149_BUFF, N3875, N150_BUFF, N153_BUFF, N204_BUFF, N2387, N400, N191_BUFF, N207_BUFF, N420, N163_BUFF, N2970, N172_BUFF, N180_BUFF, N2971, N2010, N177_BUFF, N209_BUFF, N174_BUFF, N2891, N147_BUFF, N165_BUFF, N457, N185_BUFF, N3671, N211_BUFF, N171_BUFF, N168_BUFF, N2020, N216_BUFF, N1277, N1821, N3546, N175_BUFF, N493, N1971, N181_BUFF;
  wire flip_signal;

  c2670_AntiSAT_8_0 main (N145, N153, N162, N168, N172, N210, N190, N212, N167, N185, N173, N174, N183, N196, N151, N200, N187, N195, N155, N193, N146, N163, N178, N211, N208, N177, N182, N213, N191, N216, N204, N170, N165, N179, N189, N207, N184, N148, N154, N157, N158, N164, N149, N180, N192, N156, N194, N203, N199, N171, N205, N161, N160, N176, N197, N209, N201, N202, N188, N218, N143, N175, N169, N166, N186, N159, N217, N147, N144, N181, N150, N215, N206, N198, N152, N214, N1, N2, N3, N4, N5, N6, N7, N8, N11, N14, N15, N16, N19, N20, N21, N22, N23, N24, N25, N26, N27, N28, N29, N32, N33, N34, N35, N36, N37, N40, N43, N44, N47, N48, N49, N50, N51, N52, N53, N54, N55, N56, N57, N60, N61, N62, N63, N64, N65, N66, N67, N68, N69, N72, N73, N74, N75, N76, N77, N78, N79, N80, N81, N82, N85, N86, N87, N88, N89, N90, N91, N92, N93, N94, N95, N96, N99, N100, N101, N102, N103, N104, N105, N106, N107, N108, N111, N112, N113, N114, N115, N116, N117, N118, N119, N120, N123, N124, N125, N126, N127, N128, N129, N130, N131, N132, N135, N136, N137, N138, N139, N140, N141, N142, N219, N224, N227, N230, N231, N234, N237, N241, N246, N253, N256, N259, N262, N263, N266, N269, N272, N275, N278, N281, N284, N287, N290, N294, N297, N301, N305, N309, N313, N316, N319, N322, N325, N328, N331, N334, N337, N340, N343, N346, N349, N352, N355, flip_signal, N145_BUFF, N153_BUFF, N162_BUFF, N168_BUFF, N172_BUFF, N210_BUFF, N190_BUFF, N212_BUFF, N167_BUFF, N185_BUFF, N173_BUFF, N174_BUFF, N183_BUFF, N196_BUFF, N151_BUFF, N200_BUFF, N187_BUFF, N195_BUFF, N155_BUFF, N193_BUFF, N146_BUFF, N163_BUFF, N178_BUFF, N211_BUFF, N208_BUFF, N177_BUFF, N182_BUFF, N213_BUFF, N191_BUFF, N216_BUFF, N204_BUFF, N170_BUFF, N165_BUFF, N179_BUFF, N189_BUFF, N207_BUFF, N184_BUFF, N148_BUFF, N154_BUFF, N157_BUFF, N158_BUFF, N164_BUFF, N149_BUFF, N180_BUFF, N192_BUFF, N156_BUFF, N194_BUFF, N203_BUFF, N199_BUFF, N171_BUFF, N205_BUFF, N161_BUFF, N160_BUFF, N176_BUFF, N197_BUFF, N209_BUFF, N201_BUFF, N202_BUFF, N188_BUFF, N218_BUFF, N143_BUFF, N175_BUFF, N169_BUFF, N166_BUFF, N186_BUFF, N159_BUFF, N217_BUFF, N147_BUFF, N144_BUFF, N181_BUFF, N150_BUFF, N215_BUFF, N206_BUFF, N198_BUFF, N152_BUFF, N214_BUFF, N398, N400, N401, N419, N420, N456, N457, N458, N487, N488, N489, N490, N491, N492, N493, N494, N792, N799, N805, N1026, N1028, N1029, N1269, N1277, N1448, N1726, N1816, N1817, N1818, N1819, N1820, N1821, N1969, N1970, N1971, N2010, N2012, N2014, N2016, N2018, N2020, N2022, N2387, N2388, N2389, N2390, N2496, N2643, N2644, N2891, N2925, N2970, N2971, N3038, N3079, N3546, N3671, N3803, N3804, N3809, N3851, N3875, N3881, N3882);
  SatHard flip (N96, N231, N82, N120, keyinput0, keyinput1, keyinput2, keyinput3, keyinput4, keyinput5, keyinput6, keyinput7, flip_signal);
endmodule
/*************** Top Level ***************/

// Main module
module c2670_AntiSAT_8_0(N145, N153, N162, N168, N172, N210, N190, N212, N167, N185, N173, N174, N183, N196, N151, N200, N187, N195, N155, N193, N146, N163, N178, N211, N208, N177, N182, N213, N191, N216, N204, N170, N165, N179, N189, N207, N184, N148, N154, N157, N158, N164, N149, N180, N192, N156, N194, N203, N199, N171, N205, N161, N160, N176, N197, N209, N201, N202, N188, N218, N143, N175, N169, N166, N186, N159, N217, N147, N144, N181, N150, N215, N206, N198, N152, N214, N1, N2, N3, N4, N5, N6, N7, N8, N11, N14, N15, N16, N19, N20, N21, N22, N23, N24, N25, N26, N27, N28, N29, N32, N33, N34, N35, N36, N37, N40, N43, N44, N47, N48, N49, N50, N51, N52, N53, N54, N55, N56, N57, N60, N61, N62, N63, N64, N65, N66, N67, N68, N69, N72, N73, N74, N75, N76, N77, N78, N79, N80, N81, N82, N85, N86, N87, N88, N89, N90, N91, N92, N93, N94, N95, N96, N99, N100, N101, N102, N103, N104, N105, N106, N107, N108, N111, N112, N113, N114, N115, N116, N117, N118, N119, N120, N123, N124, N125, N126, N127, N128, N129, N130, N131, N132, N135, N136, N137, N138, N139, N140, N141, N142, N219, N224, N227, N230, N231, N234, N237, N241, N246, N253, N256, N259, N262, N263, N266, N269, N272, N275, N278, N281, N284, N287, N290, N294, N297, N301, N305, N309, N313, N316, N319, N322, N325, N328, N331, N334, N337, N340, N343, N346, N349, N352, N355, flip_signal, N145_BUFF, N153_BUFF, N162_BUFF, N168_BUFF, N172_BUFF, N210_BUFF, N190_BUFF, N212_BUFF, N167_BUFF, N185_BUFF, N173_BUFF, N174_BUFF, N183_BUFF, N196_BUFF, N151_BUFF, N200_BUFF, N187_BUFF, N195_BUFF, N155_BUFF, N193_BUFF, N146_BUFF, N163_BUFF, N178_BUFF, N211_BUFF, N208_BUFF, N177_BUFF, N182_BUFF, N213_BUFF, N191_BUFF, N216_BUFF, N204_BUFF, N170_BUFF, N165_BUFF, N179_BUFF, N189_BUFF, N207_BUFF, N184_BUFF, N148_BUFF, N154_BUFF, N157_BUFF, N158_BUFF, N164_BUFF, N149_BUFF, N180_BUFF, N192_BUFF, N156_BUFF, N194_BUFF, N203_BUFF, N199_BUFF, N171_BUFF, N205_BUFF, N161_BUFF, N160_BUFF, N176_BUFF, N197_BUFF, N209_BUFF, N201_BUFF, N202_BUFF, N188_BUFF, N218_BUFF, N143_BUFF, N175_BUFF, N169_BUFF, N166_BUFF, N186_BUFF, N159_BUFF, N217_BUFF, N147_BUFF, N144_BUFF, N181_BUFF, N150_BUFF, N215_BUFF, N206_BUFF, N198_BUFF, N152_BUFF, N214_BUFF, N398, N400, N401, N419, N420, N456, N457, N458, N487, N488, N489, N490, N491, N492, N493, N494, N792, N799, N805, N1026, N1028, N1029, N1269, N1277, N1448, N1726, N1816, N1817, N1818, N1819, N1820, N1821, N1969, N1970, N1971, N2010, N2012, N2014, N2016, N2018, N2020, N2022, N2387, N2388, N2389, N2390, N2496, N2643, N2644, N2891, N2925, N2970, N2971, N3038, N3079, N3546, N3671, N3803, N3804, N3809, N3851, N3875, N3881, N3882);

  input N145, N153, N162, N168, N172, N210, N190, N212, N167, N185, N173, N174, N183, N196, N151, N200, N187, N195, N155, N193, N146, N163, N178, N211, N208, N177, N182, N213, N191, N216, N204, N170, N165, N179, N189, N207, N184, N148, N154, N157, N158, N164, N149, N180, N192, N156, N194, N203, N199, N171, N205, N161, N160, N176, N197, N209, N201, N202, N188, N218, N143, N175, N169, N166, N186, N159, N217, N147, N144, N181, N150, N215, N206, N198, N152, N214, N1, N2, N3, N4, N5, N6, N7, N8, N11, N14, N15, N16, N19, N20, N21, N22, N23, N24, N25, N26, N27, N28, N29, N32, N33, N34, N35, N36, N37, N40, N43, N44, N47, N48, N49, N50, N51, N52, N53, N54, N55, N56, N57, N60, N61, N62, N63, N64, N65, N66, N67, N68, N69, N72, N73, N74, N75, N76, N77, N78, N79, N80, N81, N82, N85, N86, N87, N88, N89, N90, N91, N92, N93, N94, N95, N96, N99, N100, N101, N102, N103, N104, N105, N106, N107, N108, N111, N112, N113, N114, N115, N116, N117, N118, N119, N120, N123, N124, N125, N126, N127, N128, N129, N130, N131, N132, N135, N136, N137, N138, N139, N140, N141, N142, N219, N224, N227, N230, N231, N234, N237, N241, N246, N253, N256, N259, N262, N263, N266, N269, N272, N275, N278, N281, N284, N287, N290, N294, N297, N301, N305, N309, N313, N316, N319, N322, N325, N328, N331, N334, N337, N340, N343, N346, N349, N352, N355, flip_signal;
  output N145_BUFF, N153_BUFF, N162_BUFF, N168_BUFF, N172_BUFF, N210_BUFF, N190_BUFF, N212_BUFF, N167_BUFF, N185_BUFF, N173_BUFF, N174_BUFF, N183_BUFF, N196_BUFF, N151_BUFF, N200_BUFF, N187_BUFF, N195_BUFF, N155_BUFF, N193_BUFF, N146_BUFF, N163_BUFF, N178_BUFF, N211_BUFF, N208_BUFF, N177_BUFF, N182_BUFF, N213_BUFF, N191_BUFF, N216_BUFF, N204_BUFF, N170_BUFF, N165_BUFF, N179_BUFF, N189_BUFF, N207_BUFF, N184_BUFF, N148_BUFF, N154_BUFF, N157_BUFF, N158_BUFF, N164_BUFF, N149_BUFF, N180_BUFF, N192_BUFF, N156_BUFF, N194_BUFF, N203_BUFF, N199_BUFF, N171_BUFF, N205_BUFF, N161_BUFF, N160_BUFF, N176_BUFF, N197_BUFF, N209_BUFF, N201_BUFF, N202_BUFF, N188_BUFF, N218_BUFF, N143_BUFF, N175_BUFF, N169_BUFF, N166_BUFF, N186_BUFF, N159_BUFF, N217_BUFF, N147_BUFF, N144_BUFF, N181_BUFF, N150_BUFF, N215_BUFF, N206_BUFF, N198_BUFF, N152_BUFF, N214_BUFF, N398, N400, N401, N419, N420, N456, N457, N458, N487, N488, N489, N490, N491, N492, N493, N494, N792, N799, N805, N1026, N1028, N1029, N1269, N1277, N1448, N1726, N1816, N1817, N1818, N1819, N1820, N1821, N1969, N1970, N1971, N2010, N2012, N2014, N2016, N2018, N2020, N2022, N2387, N2388, N2389, N2390, N2496, N2643, N2644, N2891, N2925, N2970, N2971, N3038, N3079, N3546, N3671, N3803, N3804, N3809, N3851, N3875, N3881, N3882;
  wire N1027, N1032, N1033, N1034, N1037, N1042, N1053, N1064, N1065, N1066, N1067, N1068, N1069, N1070, N1075, N1086, N1097, N1098, N1099, N1100, N1101, N1102, N1113, N1124, N1125, N1126, N1127, N1128, N1129, N1133, N1137, N1140, N1141, N1142, N1143, N1144, N1145, N1146, N1157, N1168, N1169, N1170, N1171, N1172, N1173, N1178, N1184, N1185, N1186, N1187, N1188, N1189, N1190, N1195, N1200, N1205, N1210, N1211, N1212, N1213, N1214, N1215, N1216, N1219, N1222, N1225, N1228, N1231, N1234, N1237, N1240, N1243, N1246, N1249, N1250, N1251, N1254, N1257, N1260, N1263, N1266, N1275, N1276, N1302, N1351, N1352, N1353, N1354, N1355, N1395, N1396, N1397, N1398, N1399, N1422, N1423, N1424, N1425, N1426, N1427, N1440, N1441, N1449, N1450, N1451, N1452, N1453, N1454, N1455, N1456, N1457, N1458, N1459, N1460, N1461, N1462, N1463, N1464, N1465, N1466, N1467, N1468, N1469, N1470, N1471, N1472, N1473, N1474, N1475, N1476, N1477, N1478, N1479, N1480, N1481, N1482, N1483, N1484, N1485, N1486, N1487, N1488, N1489, N1490, N1491, N1492, N1493, N1494, N1495, N1496, N1499, N1502, N1506, N1510, N1513, N1516, N1519, N1520, N1521, N1522, N1523, N1524, N1525, N1526, N1527, N1528, N1529, N1530, N1531, N1532, N1533, N1534, N1535, N1536, N1537, N1538, N1539, N1540, N1541, N1542, N1543, N1544, N1545, N1546, N1547, N1548, N1549, N1550, N1551, N1552, N1553, N1557, N1561, N1564, N1565, N1566, N1567, N1568, N1569, N1570, N1571, N1572, N1573, N1574, N1575, N1576, N1577, N1578, N1581, N1582, N1585, N1588, N1591, N1596, N1600, N1606, N1612, N1615, N1619, N1624, N1628, N1631, N1634, N1637, N1642, N1647, N1651, N1656, N1676, N1681, N1686, N1690, N1708, N1770, N1773, N1776, N1777, N1778, N1781, N1784, N1785, N1795, N1798, N1801, N1804, N1807, N1808, N1809, N1810, N1811, N1813, N1814, N1815, N1822, N1823, N1824, N1827, N1830, N1831, N1832, N1833, N1836, N1841, N1848, N1852, N1856, N1863, N1870, N1875, N1880, N1885, N1888, N1891, N1894, N1897, N1908, N1909, N1910, N1911, N1912, N1913, N1914, N1915, N1916, N1917, N1918, N1919, N1928, N1929, N1930, N1931, N1932, N1933, N1934, N1935, N1936, N1939, N1940, N1941, N1942, N1945, N1948, N1951, N1954, N1957, N1960, N1963, N1966, N2028, N2029, N2030, N2031, N2032, N2033, N2034, N2040, N2041, N2042, N2043, N2046, N2049, N2052, N2055, N2058, N2061, N2064, N2067, N2070, N2073, N2076, N2079, N2095, N2098, N2101, N2104, N2107, N2110, N2113, N2119, N2120, N2125, N2126, N2127, N2128, N2135, N2141, N2144, N2147, N2150, N2153, N2154, N2155, N2156, N2157, N2158, N2171, N2172, N2173, N2174, N2175, N2176, N2177, N2178, N2185, N2188, N2191, N2194, N2197, N2200, N2201, N2204, N2207, N2210, N2213, N2216, N2219, N2234, N2235, N2236, N2237, N2250, N2266, N2269, N2291, N2294, N2297, N2298, N2300, N2301, N2302, N2303, N2304, N2305, N2306, N2307, N2308, N2309, N2310, N2311, N2312, N2313, N2314, N2315, N2316, N2317, N2318, N2319, N2320, N2321, N2322, N2323, N2324, N2325, N2326, N2327, N2328, N2329, N2330, N2331, N2332, N2333, N2334, N2335, N2336, N2337, N2338, N2339, N2340, N2354, N2355, N2356, N2357, N2358, N2359, N2364, N2365, N2366, N2367, N2368, N2372, N2373, N2374, N2375, N2376, N2377, N2382, N2386, N2391, N2395, N2400, N2403, N2406, N2407, N2408, N2409, N2410, N2411, N2412, N2413, N2414, N2415, N2416, N2417, N2421, N2425, N2428, N2429, N2430, N2431, N2432, N2433, N2434, N2437, N2440, N2443, N2446, N2449, N2452, N2453, N2454, N2457, N2460, N2463, N2466, N2469, N2472, N2475, N2478, N2481, N2484, N2487, N2490, N2493, N2503, N2504, N2510, N2511, N2521, N2528, N2531, N2534, N2537, N2540, N2544, N2545, N2546, N2547, N2548, N2549, N2550, N2551, N2552, N2553, N2563, N2564, N2565, N2566, N2567, N2568, N2579, N2603, N2607, N2608, N2609, N2610, N2611, N2612, N2613, N2617, N2618, N2619, N2620, N2621, N2624, N2628, N2629, N2630, N2631, N2632, N2633, N2634, N2635, N2636, N2638, N2645, N2646, N2652, N2655, N2656, N2659, N2663, N2664, N2665, N2666, N2667, N2668, N2669, N2670, N2671, N2672, N2673, N2674, N2675, N2676, N2677, N2678, N2679, N2680, N2681, N2684, N2687, N2690, N2693, N2694, N2695, N2696, N2697, N2698, N2699, N2700, N2701, N2702, N2703, N2706, N2707, N2708, N2709, N2710, N2719, N2720, N2726, N2729, N2738, N2743, N2747, N2748, N2749, N2750, N2751, N2760, N2761, N2766, N2771, N2772, N2773, N2774, N2775, N2776, N2777, N2778, N2781, N2782, N2783, N2784, N2789, N2790, N2791, N2792, N2793, N2796, N2800, N2803, N2806, N2809, N2810, N2811, N2812, N2817, N2820, N2826, N2829, N2830, N2831, N2837, N2838, N2839, N2840, N2841, N2844, N2854, N2859, N2869, N2874, N2877, N2880, N2881, N2882, N2885, N2888, N2894, N2895, N2896, N2897, N2898, N2899, N2900, N2901, N2914, N2915, N2916, N2917, N2918, N2919, N2920, N2921, N2931, N2938, N2939, N2963, N2972, N2975, N2978, N2981, N2984, N2985, N2986, N2989, N2992, N2995, N2998, N3001, N3004, N3007, N3008, N3009, N3010, N3013, N3016, N3019, N3022, N3025, N3028, N3029, N3030, N3035, N3036, N3037, N3039, N3044, N3045, N3046, N3047, N3048, N3049, N3050, N3053, N3054, N3055, N3056, N3057, N3058, N3059, N3060, N3061, N3064, N3065, N3066, N3067, N3068, N3069, N3070, N3071, N3072, N3073, N3074, N3075, N3076, N3088, N3091, N3110, N3113, N3137, N3140, N3143, N3146, N3149, N3152, N3157, N3160, N3163, N3166, N3169, N3172, N3175, N3176, N3177, N3178, N3180, N3187, N3188, N3189, N3190, N3191, N3192, N3193, N3194, N3195, N3196, N3197, N3208, N3215, N3216, N3217, N3218, N3219, N3220, N3222, N3223, N3230, N3231, N3238, N3241, N3244, N3247, N3250, N3253, N3256, N3259, N3262, N3265, N3268, N3271, N3274, N3277, N3281, N3282, N3283, N3284, N3286, N3288, N3289, N3291, N3293, N3295, N3296, N3299, N3301, N3302, N3304, N3306, N3308, N3309, N3312, N3314, N3315, N3318, N3321, N3324, N3327, N3330, N3333, N3334, N3335, N3336, N3337, N3340, N3344, N3348, N3352, N3356, N3360, N3364, N3367, N3370, N3374, N3378, N3382, N3386, N3390, N3394, N3397, N3400, N3401, N3402, N3403, N3404, N3405, N3406, N3409, N3410, N3412, N3414, N3416, N3418, N3420, N3422, N3428, N3430, N3432, N3434, N3436, N3438, N3440, N3450, N3453, N3456, N3459, N3478, N3479, N3480, N3481, N3482, N3483, N3484, N3485, N3486, N3487, N3488, N3489, N3490, N3491, N3492, N3493, N3494, N3496, N3498, N3499, N3500, N3501, N3502, N3503, N3504, N3505, N3506, N3507, N3508, N3509, N3510, N3511, N3512, N3513, N3515, N3517, N3522, N3525, N3528, N3531, N3534, N3537, N3540, N3543, N3551, N3552, N3553, N3554, N3555, N3556, N3557, N3558, N3559, N3563, N3564, N3565, N3566, N3567, N3568, N3569, N3570, N3576, N3579, N3585, N3588, N3592, N3593, N3594, N3595, N3596, N3597, N3598, N3599, N3600, N3603, N3608, N3612, N3615, N3616, N3622, N3629, N3630, N3631, N3632, N3633, N3634, N3635, N3640, N3644, N3647, N3648, N3654, N3661, N3662, N3667, N3668, N3669, N3670, N3691, N3692, N3693, N3694, N3695, N3696, N3697, N3716, N3717, N3718, N3719, N3720, N3721, N3722, N3723, N3726, N3727, N3728, N3729, N3730, N3731, N3732, N3733, N3734, N3735, N3736, N3737, N3740, N3741, N3742, N3743, N3744, N3745, N3746, N3747, N3748, N3749, N3750, N3753, N3754, N3758, N3761, N3762, N3767, N3771, N3774, N3775, N3778, N3779, N3780, N3790, N3793, N3794, N3802, N3805, N3806, N3807, N3808, N3811, N3812, N3813, N3814, N3815, N3816, N3817, N3818, N3819, N3820, N3821, N3822, N3823, N3826, N3827, N3834, N3835, N3836, N3837, N3838, N3839, N3840, N3843, N3852, N3857, N3858, N3859, N3864, N3869, N3870, N3876, N3877, N405, N408, N425, N485, N486, N495, N496, N499, N500, N503, N506, N509, N521, N533, N537, N543, N544, N547, N550, N562, N574, N578, N582, N594, N606, N607, N608, N609, N610, N611, N612, N613, N625, N637, N643, N650, N651, N655, N659, N663, N667, N671, N675, N679, N683, N687, N693, N699, N705, N711, N715, N719, N723, N727, N730, N733, N734, N735, N738, N741, N744, N747, N750, N753, N756, N759, N762, N765, N768, N771, N774, N777, N780, N783, N786, N800, N900, N901, N902, N903, N904, N905, N998, N999, N1726_in;

  and ginst1 (N1026, N94, N500);
  and ginst2 (N1027, N325, N651);
  not ginst3 (N1028, N651);
  nand ginst4 (N1029, N231, N651);
  not ginst5 (N1032, N544);
  not ginst6 (N1033, N547);
  and ginst7 (N1034, N544, N547);
  buf ginst8 (N1037, N503);
  not ginst9 (N1042, N509);
  not ginst10 (N1053, N521);
  and ginst11 (N1064, N80, N509, N521);
  and ginst12 (N1065, N68, N509, N521);
  and ginst13 (N1066, N79, N509, N521);
  and ginst14 (N1067, N78, N509, N521);
  and ginst15 (N1068, N77, N509, N521);
  and ginst16 (N1069, N11, N537);
  buf ginst17 (N1070, N503);
  not ginst18 (N1075, N550);
  not ginst19 (N1086, N562);
  and ginst20 (N1097, N76, N550, N562);
  and ginst21 (N1098, N75, N550, N562);
  and ginst22 (N1099, N74, N550, N562);
  and ginst23 (N1100, N73, N550, N562);
  and ginst24 (N1101, N72, N550, N562);
  not ginst25 (N1102, N582);
  not ginst26 (N1113, N594);
  and ginst27 (N1124, N114, N582, N594);
  and ginst28 (N1125, N113, N582, N594);
  and ginst29 (N1126, N112, N582, N594);
  and ginst30 (N1127, N111, N582, N594);
  and ginst31 (N1128, N582, N594);
  nand ginst32 (N1129, N900, N901);
  nand ginst33 (N1133, N902, N903);
  nand ginst34 (N1137, N904, N905);
  not ginst35 (N1140, N741);
  nand ginst36 (N1141, N612, N741);
  not ginst37 (N1142, N744);
  not ginst38 (N1143, N747);
  not ginst39 (N1144, N750);
  not ginst40 (N1145, N753);
  not ginst41 (N1146, N613);
  not ginst42 (N1157, N625);
  and ginst43 (N1168, N118, N613, N625);
  and ginst44 (N1169, N107, N613, N625);
  and ginst45 (N1170, N117, N613, N625);
  and ginst46 (N1171, N116, N613, N625);
  and ginst47 (N1172, N115, N613, N625);
  not ginst48 (N1173, N637);
  not ginst49 (N1178, N643);
  not ginst50 (N1184, N768);
  nand ginst51 (N1185, N650, N768);
  not ginst52 (N1186, N771);
  not ginst53 (N1187, N774);
  not ginst54 (N1188, N777);
  not ginst55 (N1189, N780);
  buf ginst56 (N1190, N506);
  buf ginst57 (N1195, N506);
  not ginst58 (N1200, N693);
  not ginst59 (N1205, N699);
  not ginst60 (N1210, N735);
  not ginst61 (N1211, N738);
  not ginst62 (N1212, N756);
  not ginst63 (N1213, N759);
  not ginst64 (N1214, N762);
  not ginst65 (N1215, N765);
  nand ginst66 (N1216, N998, N999);
  buf ginst67 (N1219, N574);
  buf ginst68 (N1222, N578);
  buf ginst69 (N1225, N655);
  buf ginst70 (N1228, N659);
  buf ginst71 (N1231, N663);
  buf ginst72 (N1234, N667);
  buf ginst73 (N1237, N671);
  buf ginst74 (N1240, N675);
  buf ginst75 (N1243, N679);
  buf ginst76 (N1246, N683);
  not ginst77 (N1249, N783);
  not ginst78 (N1250, N786);
  buf ginst79 (N1251, N687);
  buf ginst80 (N1254, N705);
  buf ginst81 (N1257, N711);
  buf ginst82 (N1260, N715);
  buf ginst83 (N1263, N719);
  buf ginst84 (N1266, N723);
  not ginst85 (N1269, N1027);
  and ginst86 (N1275, N325, N1032);
  and ginst87 (N1276, N231, N1033);
  buf ginst88 (N1277, N1034);
  or ginst89 (N1302, N1069, N543);
  nand ginst90 (N1351, N352, N1140);
  nand ginst91 (N1352, N1142, N747);
  nand ginst92 (N1353, N1143, N744);
  nand ginst93 (N1354, N1144, N753);
  nand ginst94 (N1355, N1145, N750);
  nand ginst95 (N1395, N355, N1184);
  nand ginst96 (N1396, N1186, N774);
  nand ginst97 (N1397, N1187, N771);
  nand ginst98 (N1398, N1188, N780);
  nand ginst99 (N1399, N1189, N777);
  nand ginst100 (N1422, N1210, N738);
  nand ginst101 (N1423, N1211, N735);
  nand ginst102 (N1424, N1212, N759);
  nand ginst103 (N1425, N1213, N756);
  nand ginst104 (N1426, N1214, N765);
  nand ginst105 (N1427, N1215, N762);
  buf ginst106 (N143_BUFF, N143);
  nand ginst107 (N1440, N1249, N786);
  nand ginst108 (N1441, N1250, N783);
  not ginst109 (N1448, N1034);
  not ginst110 (N1449, N1275);
  buf ginst111 (N144_BUFF, N144);
  not ginst112 (N1450, N1276);
  and ginst113 (N1451, N93, N1042, N1053);
  and ginst114 (N1452, N55, N1053, N509);
  and ginst115 (N1453, N67, N1042, N521);
  and ginst116 (N1454, N81, N1042, N1053);
  and ginst117 (N1455, N43, N1053, N509);
  and ginst118 (N1456, N56, N1042, N521);
  and ginst119 (N1457, N92, N1042, N1053);
  and ginst120 (N1458, N54, N1053, N509);
  and ginst121 (N1459, N66, N1042, N521);
  buf ginst122 (N145_BUFF, N145);
  and ginst123 (N1460, N91, N1042, N1053);
  and ginst124 (N1461, N53, N1053, N509);
  and ginst125 (N1462, N65, N1042, N521);
  and ginst126 (N1463, N90, N1042, N1053);
  and ginst127 (N1464, N52, N1053, N509);
  and ginst128 (N1465, N64, N1042, N521);
  and ginst129 (N1466, N89, N1075, N1086);
  and ginst130 (N1467, N51, N1086, N550);
  and ginst131 (N1468, N63, N1075, N562);
  and ginst132 (N1469, N88, N1075, N1086);
  buf ginst133 (N146_BUFF, N146);
  and ginst134 (N1470, N50, N1086, N550);
  and ginst135 (N1471, N62, N1075, N562);
  and ginst136 (N1472, N87, N1075, N1086);
  and ginst137 (N1473, N49, N1086, N550);
  and ginst138 (N1474, N1075, N562);
  and ginst139 (N1475, N86, N1075, N1086);
  and ginst140 (N1476, N48, N1086, N550);
  and ginst141 (N1477, N61, N1075, N562);
  and ginst142 (N1478, N85, N1075, N1086);
  and ginst143 (N1479, N47, N1086, N550);
  buf ginst144 (N147_BUFF, N147);
  and ginst145 (N1480, N60, N1075, N562);
  and ginst146 (N1481, N138, N1102, N1113);
  and ginst147 (N1482, N102, N1113, N582);
  and ginst148 (N1483, N126, N1102, N594);
  and ginst149 (N1484, N137, N1102, N1113);
  and ginst150 (N1485, N101, N1113, N582);
  and ginst151 (N1486, N125, N1102, N594);
  and ginst152 (N1487, N136, N1102, N1113);
  and ginst153 (N1488, N100, N1113, N582);
  and ginst154 (N1489, N124, N1102, N594);
  buf ginst155 (N148_BUFF, N148);
  and ginst156 (N1490, N135, N1102, N1113);
  and ginst157 (N1491, N99, N1113, N582);
  and ginst158 (N1492, N123, N1102, N594);
  and ginst159 (N1493, N1102, N1113);
  and ginst160 (N1494, N1113, N582);
  and ginst161 (N1495, N1102, N594);
  not ginst162 (N1496, N1129);
  not ginst163 (N1499, N1133);
  buf ginst164 (N149_BUFF, N149);
  nand ginst165 (N1502, N1141, N1351);
  nand ginst166 (N1506, N1352, N1353);
  buf ginst167 (N150_BUFF, N150);
  nand ginst168 (N1510, N1354, N1355);
  buf ginst169 (N1513, N1137);
  buf ginst170 (N1516, N1137);
  not ginst171 (N1519, N1219);
  buf ginst172 (N151_BUFF, N151);
  not ginst173 (N1520, N1222);
  not ginst174 (N1521, N1225);
  not ginst175 (N1522, N1228);
  not ginst176 (N1523, N1231);
  not ginst177 (N1524, N1234);
  not ginst178 (N1525, N1237);
  not ginst179 (N1526, N1240);
  not ginst180 (N1527, N1243);
  not ginst181 (N1528, N1246);
  and ginst182 (N1529, N142, N1146, N1157);
  buf ginst183 (N152_BUFF, N152);
  and ginst184 (N1530, N106, N1157, N613);
  and ginst185 (N1531, N130, N1146, N625);
  and ginst186 (N1532, N131, N1146, N1157);
  and ginst187 (N1533, N95, N1157, N613);
  and ginst188 (N1534, N119, N1146, N625);
  and ginst189 (N1535, N141, N1146, N1157);
  and ginst190 (N1536, N105, N1157, N613);
  and ginst191 (N1537, N129, N1146, N625);
  and ginst192 (N1538, N140, N1146, N1157);
  and ginst193 (N1539, N104, N1157, N613);
  buf ginst194 (N153_BUFF, N153);
  and ginst195 (N1540, N128, N1146, N625);
  and ginst196 (N1541, N139, N1146, N1157);
  and ginst197 (N1542, N103, N1157, N613);
  and ginst198 (N1543, N127, N1146, N625);
  and ginst199 (N1544, N19, N1173);
  and ginst200 (N1545, N4, N1173);
  and ginst201 (N1546, N20, N1173);
  and ginst202 (N1547, N5, N1173);
  and ginst203 (N1548, N21, N1178);
  and ginst204 (N1549, N22, N1178);
  buf ginst205 (N154_BUFF, N154);
  and ginst206 (N1550, N23, N1178);
  and ginst207 (N1551, N6, N1178);
  and ginst208 (N1552, N24, N1178);
  nand ginst209 (N1553, N1185, N1395);
  nand ginst210 (N1557, N1396, N1397);
  buf ginst211 (N155_BUFF, N155);
  nand ginst212 (N1561, N1398, N1399);
  and ginst213 (N1564, N25, N1200);
  and ginst214 (N1565, N32, N1200);
  and ginst215 (N1566, N26, N1200);
  and ginst216 (N1567, N33, N1200);
  and ginst217 (N1568, N27, N1205);
  and ginst218 (N1569, N34, N1205);
  buf ginst219 (N156_BUFF, N156);
  and ginst220 (N1570, N35, N1205);
  and ginst221 (N1571, N28, N1205);
  not ginst222 (N1572, N1251);
  not ginst223 (N1573, N1254);
  not ginst224 (N1574, N1257);
  not ginst225 (N1575, N1260);
  not ginst226 (N1576, N1263);
  not ginst227 (N1577, N1266);
  nand ginst228 (N1578, N1422, N1423);
  buf ginst229 (N157_BUFF, N157);
  not ginst230 (N1581, N1216);
  nand ginst231 (N1582, N1426, N1427);
  nand ginst232 (N1585, N1424, N1425);
  nand ginst233 (N1588, N1440, N1441);
  buf ginst234 (N158_BUFF, N158);
  and ginst235 (N1591, N1449, N1450);
  or ginst236 (N1596, N1064, N1451, N1452, N1453);
  buf ginst237 (N159_BUFF, N159);
  or ginst238 (N1600, N1065, N1454, N1455, N1456);
  or ginst239 (N1606, N1066, N1457, N1458, N1459);
  buf ginst240 (N160_BUFF, N160);
  or ginst241 (N1612, N1067, N1460, N1461, N1462);
  or ginst242 (N1615, N1068, N1463, N1464, N1465);
  or ginst243 (N1619, N1097, N1466, N1467, N1468);
  buf ginst244 (N161_BUFF, N161);
  or ginst245 (N1624, N1098, N1469, N1470, N1471);
  or ginst246 (N1628, N1099, N1472, N1473, N1474);
  buf ginst247 (N162_BUFF, N162);
  or ginst248 (N1631, N1100, N1475, N1476, N1477);
  or ginst249 (N1634, N1101, N1478, N1479, N1480);
  or ginst250 (N1637, N1124, N1481, N1482, N1483);
  buf ginst251 (N163_BUFF, N163);
  or ginst252 (N1642, N1125, N1484, N1485, N1486);
  or ginst253 (N1647, N1126, N1487, N1488, N1489);
  buf ginst254 (N164_BUFF, N164);
  or ginst255 (N1651, N1127, N1490, N1491, N1492);
  or ginst256 (N1656, N1128, N1493, N1494, N1495);
  buf ginst257 (N165_BUFF, N165);
  buf ginst258 (N166_BUFF, N166);
  or ginst259 (N1676, N1169, N1532, N1533, N1534);
  buf ginst260 (N167_BUFF, N167);
  or ginst261 (N1681, N1170, N1535, N1536, N1537);
  or ginst262 (N1686, N1171, N1538, N1539, N1540);
  buf ginst263 (N168_BUFF, N168);
  or ginst264 (N1690, N1172, N1541, N1542, N1543);
  buf ginst265 (N169_BUFF, N169);
  or ginst266 (N1708, N1168, N1529, N1530, N1531);
  buf ginst267 (N170_BUFF, N170);
  buf ginst268 (N171_BUFF, N171);
  xor ginst269 (N1726, N1726_in, flip_signal);
  buf ginst270 (N1726_in, N1591);
  buf ginst271 (N172_BUFF, N172);
  buf ginst272 (N173_BUFF, N173);
  buf ginst273 (N174_BUFF, N174);
  buf ginst274 (N175_BUFF, N175);
  buf ginst275 (N176_BUFF, N176);
  not ginst276 (N1770, N1502);
  not ginst277 (N1773, N1506);
  not ginst278 (N1776, N1513);
  not ginst279 (N1777, N1516);
  buf ginst280 (N1778, N1510);
  buf ginst281 (N177_BUFF, N177);
  buf ginst282 (N1781, N1510);
  and ginst283 (N1784, N1129, N1133, N1513);
  and ginst284 (N1785, N1496, N1499, N1516);
  buf ginst285 (N178_BUFF, N178);
  not ginst286 (N1795, N1553);
  not ginst287 (N1798, N1557);
  buf ginst288 (N179_BUFF, N179);
  buf ginst289 (N1801, N1561);
  buf ginst290 (N1804, N1561);
  not ginst291 (N1807, N1588);
  not ginst292 (N1808, N1578);
  nand ginst293 (N1809, N1578, N1581);
  buf ginst294 (N180_BUFF, N180);
  not ginst295 (N1810, N1582);
  not ginst296 (N1811, N1585);
  and ginst297 (N1813, N241, N1596);
  and ginst298 (N1814, N241, N1606);
  and ginst299 (N1815, N241, N1600);
  not ginst300 (N1816, N1642);
  not ginst301 (N1817, N1647);
  not ginst302 (N1818, N1637);
  not ginst303 (N1819, N1624);
  buf ginst304 (N181_BUFF, N181);
  not ginst305 (N1820, N1619);
  not ginst306 (N1821, N1615);
  and ginst307 (N1822, N36, N224, N1591, N496);
  and ginst308 (N1823, N224, N1591, N486, N496);
  buf ginst309 (N1824, N1596);
  not ginst310 (N1827, N1606);
  buf ginst311 (N182_BUFF, N182);
  and ginst312 (N1830, N1600, N537);
  and ginst313 (N1831, N1606, N537);
  and ginst314 (N1832, N246, N1619);
  not ginst315 (N1833, N1596);
  not ginst316 (N1836, N1600);
  buf ginst317 (N183_BUFF, N183);
  not ginst318 (N1841, N1606);
  buf ginst319 (N1848, N1612);
  buf ginst320 (N184_BUFF, N184);
  buf ginst321 (N1852, N1615);
  buf ginst322 (N1856, N1619);
  buf ginst323 (N185_BUFF, N185);
  buf ginst324 (N1863, N1624);
  buf ginst325 (N186_BUFF, N186);
  buf ginst326 (N1870, N1628);
  buf ginst327 (N1875, N1631);
  buf ginst328 (N187_BUFF, N187);
  buf ginst329 (N1880, N1634);
  nand ginst330 (N1885, N1651, N727);
  nand ginst331 (N1888, N1656, N730);
  buf ginst332 (N188_BUFF, N188);
  buf ginst333 (N1891, N1686);
  and ginst334 (N1894, N1637, N425);
  not ginst335 (N1897, N1642);
  buf ginst336 (N189_BUFF, N189);
  and ginst337 (N1908, N1133, N1496, N1776);
  and ginst338 (N1909, N1129, N1499, N1777);
  buf ginst339 (N190_BUFF, N190);
  and ginst340 (N1910, N1600, N637);
  and ginst341 (N1911, N1606, N637);
  and ginst342 (N1912, N1612, N637);
  and ginst343 (N1913, N1615, N637);
  and ginst344 (N1914, N1619, N643);
  and ginst345 (N1915, N1624, N643);
  and ginst346 (N1916, N1628, N643);
  and ginst347 (N1917, N1631, N643);
  and ginst348 (N1918, N1634, N643);
  not ginst349 (N1919, N1708);
  buf ginst350 (N191_BUFF, N191);
  and ginst351 (N1928, N1676, N693);
  and ginst352 (N1929, N1681, N693);
  buf ginst353 (N192_BUFF, N192);
  and ginst354 (N1930, N1686, N693);
  and ginst355 (N1931, N1690, N693);
  and ginst356 (N1932, N1637, N699);
  and ginst357 (N1933, N1642, N699);
  and ginst358 (N1934, N1647, N699);
  and ginst359 (N1935, N1651, N699);
  buf ginst360 (N1936, N1600);
  nand ginst361 (N1939, N1216, N1808);
  buf ginst362 (N193_BUFF, N193);
  nand ginst363 (N1940, N1585, N1810);
  nand ginst364 (N1941, N1582, N1811);
  buf ginst365 (N1942, N1676);
  buf ginst366 (N1945, N1686);
  buf ginst367 (N1948, N1681);
  buf ginst368 (N194_BUFF, N194);
  buf ginst369 (N1951, N1637);
  buf ginst370 (N1954, N1690);
  buf ginst371 (N1957, N1647);
  buf ginst372 (N195_BUFF, N195);
  buf ginst373 (N1960, N1642);
  buf ginst374 (N1963, N1656);
  buf ginst375 (N1966, N1651);
  or ginst376 (N1969, N1815, N533);
  buf ginst377 (N196_BUFF, N196);
  not ginst378 (N1970, N1822);
  not ginst379 (N1971, N1823);
  buf ginst380 (N197_BUFF, N197);
  buf ginst381 (N198_BUFF, N198);
  buf ginst382 (N199_BUFF, N199);
  buf ginst383 (N200_BUFF, N200);
  buf ginst384 (N2010, N1848);
  buf ginst385 (N2012, N1852);
  buf ginst386 (N2014, N1856);
  buf ginst387 (N2016, N1863);
  buf ginst388 (N2018, N1870);
  buf ginst389 (N201_BUFF, N201);
  buf ginst390 (N2020, N1875);
  buf ginst391 (N2022, N1880);
  not ginst392 (N2028, N1778);
  not ginst393 (N2029, N1781);
  buf ginst394 (N202_BUFF, N202);
  nor ginst395 (N2030, N1784, N1908);
  nor ginst396 (N2031, N1785, N1909);
  and ginst397 (N2032, N1502, N1506, N1778);
  and ginst398 (N2033, N1770, N1773, N1781);
  or ginst399 (N2034, N1571, N1935);
  buf ginst400 (N203_BUFF, N203);
  not ginst401 (N2040, N1801);
  not ginst402 (N2041, N1804);
  and ginst403 (N2042, N1553, N1557, N1801);
  and ginst404 (N2043, N1795, N1798, N1804);
  nand ginst405 (N2046, N1809, N1939);
  nand ginst406 (N2049, N1940, N1941);
  buf ginst407 (N204_BUFF, N204);
  or ginst408 (N2052, N1544, N1910);
  or ginst409 (N2055, N1545, N1911);
  or ginst410 (N2058, N1546, N1912);
  buf ginst411 (N205_BUFF, N205);
  or ginst412 (N2061, N1547, N1913);
  or ginst413 (N2064, N1548, N1914);
  or ginst414 (N2067, N1549, N1915);
  buf ginst415 (N206_BUFF, N206);
  or ginst416 (N2070, N1550, N1916);
  or ginst417 (N2073, N1551, N1917);
  or ginst418 (N2076, N1552, N1918);
  or ginst419 (N2079, N1564, N1928);
  buf ginst420 (N207_BUFF, N207);
  buf ginst421 (N208_BUFF, N208);
  or ginst422 (N2095, N1565, N1929);
  or ginst423 (N2098, N1566, N1930);
  buf ginst424 (N209_BUFF, N209);
  or ginst425 (N2101, N1567, N1931);
  or ginst426 (N2104, N1568, N1932);
  or ginst427 (N2107, N1569, N1933);
  buf ginst428 (N210_BUFF, N210);
  or ginst429 (N2110, N1570, N1934);
  and ginst430 (N2113, N40, N1894, N1897);
  not ginst431 (N2119, N1894);
  buf ginst432 (N211_BUFF, N211);
  nand ginst433 (N2120, N1827, N408);
  and ginst434 (N2125, N1824, N537);
  and ginst435 (N2126, N246, N1852);
  and ginst436 (N2127, N1848, N537);
  not ginst437 (N2128, N1848);
  buf ginst438 (N212_BUFF, N212);
  not ginst439 (N2135, N1852);
  buf ginst440 (N213_BUFF, N213);
  not ginst441 (N2141, N1863);
  not ginst442 (N2144, N1870);
  not ginst443 (N2147, N1875);
  buf ginst444 (N214_BUFF, N214);
  not ginst445 (N2150, N1880);
  and ginst446 (N2153, N1885, N727);
  and ginst447 (N2154, N1651, N1885);
  and ginst448 (N2155, N1888, N730);
  and ginst449 (N2156, N1656, N1888);
  and ginst450 (N2157, N1506, N1770, N2028);
  and ginst451 (N2158, N1502, N1773, N2029);
  buf ginst452 (N215_BUFF, N215);
  buf ginst453 (N216_BUFF, N216);
  not ginst454 (N2171, N1942);
  nand ginst455 (N2172, N1919, N1942);
  not ginst456 (N2173, N1945);
  not ginst457 (N2174, N1948);
  not ginst458 (N2175, N1951);
  not ginst459 (N2176, N1954);
  and ginst460 (N2177, N1557, N1795, N2040);
  and ginst461 (N2178, N1553, N1798, N2041);
  buf ginst462 (N217_BUFF, N217);
  buf ginst463 (N2185, N1836);
  buf ginst464 (N2188, N1833);
  buf ginst465 (N218_BUFF, N218);
  buf ginst466 (N2191, N1841);
  not ginst467 (N2194, N1856);
  not ginst468 (N2197, N1827);
  not ginst469 (N2200, N1936);
  buf ginst470 (N2201, N1836);
  buf ginst471 (N2204, N1833);
  buf ginst472 (N2207, N1841);
  buf ginst473 (N2210, N1824);
  buf ginst474 (N2213, N1841);
  buf ginst475 (N2216, N1841);
  nand ginst476 (N2219, N2030, N2031);
  not ginst477 (N2234, N1957);
  not ginst478 (N2235, N1960);
  not ginst479 (N2236, N1963);
  not ginst480 (N2237, N1966);
  and ginst481 (N2250, N40, N1897, N2119);
  or ginst482 (N2266, N1831, N2126);
  or ginst483 (N2269, N1832, N2127);
  or ginst484 (N2291, N2153, N2154);
  or ginst485 (N2294, N2155, N2156);
  nor ginst486 (N2297, N2032, N2157);
  nor ginst487 (N2298, N2033, N2158);
  not ginst488 (N2300, N2046);
  not ginst489 (N2301, N2049);
  nand ginst490 (N2302, N1519, N2052);
  not ginst491 (N2303, N2052);
  nand ginst492 (N2304, N1520, N2055);
  not ginst493 (N2305, N2055);
  nand ginst494 (N2306, N1521, N2058);
  not ginst495 (N2307, N2058);
  nand ginst496 (N2308, N1522, N2061);
  not ginst497 (N2309, N2061);
  nand ginst498 (N2310, N1523, N2064);
  not ginst499 (N2311, N2064);
  nand ginst500 (N2312, N1524, N2067);
  not ginst501 (N2313, N2067);
  nand ginst502 (N2314, N1525, N2070);
  not ginst503 (N2315, N2070);
  nand ginst504 (N2316, N1526, N2073);
  not ginst505 (N2317, N2073);
  nand ginst506 (N2318, N1527, N2076);
  not ginst507 (N2319, N2076);
  nand ginst508 (N2320, N1528, N2079);
  not ginst509 (N2321, N2079);
  nand ginst510 (N2322, N1708, N2171);
  nand ginst511 (N2323, N1948, N2173);
  nand ginst512 (N2324, N1945, N2174);
  nand ginst513 (N2325, N1954, N2175);
  nand ginst514 (N2326, N1951, N2176);
  nor ginst515 (N2327, N2042, N2177);
  nor ginst516 (N2328, N2043, N2178);
  nand ginst517 (N2329, N1572, N2095);
  not ginst518 (N2330, N2095);
  nand ginst519 (N2331, N1573, N2098);
  not ginst520 (N2332, N2098);
  nand ginst521 (N2333, N1574, N2101);
  not ginst522 (N2334, N2101);
  nand ginst523 (N2335, N1575, N2104);
  not ginst524 (N2336, N2104);
  nand ginst525 (N2337, N1576, N2107);
  not ginst526 (N2338, N2107);
  nand ginst527 (N2339, N1577, N2110);
  not ginst528 (N2340, N2110);
  nand ginst529 (N2354, N1960, N2234);
  nand ginst530 (N2355, N1957, N2235);
  nand ginst531 (N2356, N1966, N2236);
  nand ginst532 (N2357, N1963, N2237);
  and ginst533 (N2358, N2120, N533);
  not ginst534 (N2359, N2113);
  not ginst535 (N2364, N2185);
  not ginst536 (N2365, N2188);
  not ginst537 (N2366, N2191);
  not ginst538 (N2367, N2194);
  buf ginst539 (N2368, N2120);
  not ginst540 (N2372, N2201);
  not ginst541 (N2373, N2204);
  not ginst542 (N2374, N2207);
  not ginst543 (N2375, N2210);
  not ginst544 (N2376, N2213);
  not ginst545 (N2377, N2113);
  buf ginst546 (N2382, N2113);
  and ginst547 (N2386, N246, N2120);
  buf ginst548 (N2387, N2266);
  buf ginst549 (N2388, N2266);
  buf ginst550 (N2389, N2269);
  buf ginst551 (N2390, N2269);
  buf ginst552 (N2391, N2113);
  not ginst553 (N2395, N2113);
  nand ginst554 (N2400, N2219, N2300);
  not ginst555 (N2403, N2216);
  not ginst556 (N2406, N2219);
  nand ginst557 (N2407, N1219, N2303);
  nand ginst558 (N2408, N1222, N2305);
  nand ginst559 (N2409, N1225, N2307);
  nand ginst560 (N2410, N1228, N2309);
  nand ginst561 (N2411, N1231, N2311);
  nand ginst562 (N2412, N1234, N2313);
  nand ginst563 (N2413, N1237, N2315);
  nand ginst564 (N2414, N1240, N2317);
  nand ginst565 (N2415, N1243, N2319);
  nand ginst566 (N2416, N1246, N2321);
  nand ginst567 (N2417, N2172, N2322);
  nand ginst568 (N2421, N2323, N2324);
  nand ginst569 (N2425, N2325, N2326);
  nand ginst570 (N2428, N1251, N2330);
  nand ginst571 (N2429, N1254, N2332);
  nand ginst572 (N2430, N1257, N2334);
  nand ginst573 (N2431, N1260, N2336);
  nand ginst574 (N2432, N1263, N2338);
  nand ginst575 (N2433, N1266, N2340);
  buf ginst576 (N2434, N2128);
  buf ginst577 (N2437, N2135);
  buf ginst578 (N2440, N2144);
  buf ginst579 (N2443, N2141);
  buf ginst580 (N2446, N2150);
  buf ginst581 (N2449, N2147);
  not ginst582 (N2452, N2197);
  nand ginst583 (N2453, N2197, N2200);
  buf ginst584 (N2454, N2128);
  buf ginst585 (N2457, N2144);
  buf ginst586 (N2460, N2141);
  buf ginst587 (N2463, N2150);
  buf ginst588 (N2466, N2147);
  not ginst589 (N2469, N2120);
  buf ginst590 (N2472, N2128);
  buf ginst591 (N2475, N2135);
  buf ginst592 (N2478, N2128);
  buf ginst593 (N2481, N2135);
  nand ginst594 (N2484, N2297, N2298);
  nand ginst595 (N2487, N2356, N2357);
  nand ginst596 (N2490, N2354, N2355);
  nand ginst597 (N2493, N2327, N2328);
  or ginst598 (N2496, N1814, N2358);
  nand ginst599 (N2503, N2188, N2364);
  nand ginst600 (N2504, N2185, N2365);
  nand ginst601 (N2510, N2204, N2372);
  nand ginst602 (N2511, N2201, N2373);
  or ginst603 (N2521, N1830, N2386);
  nand ginst604 (N2528, N2046, N2406);
  not ginst605 (N2531, N2291);
  not ginst606 (N2534, N2294);
  buf ginst607 (N2537, N2250);
  buf ginst608 (N2540, N2250);
  nand ginst609 (N2544, N2302, N2407);
  nand ginst610 (N2545, N2304, N2408);
  nand ginst611 (N2546, N2306, N2409);
  nand ginst612 (N2547, N2308, N2410);
  nand ginst613 (N2548, N2310, N2411);
  nand ginst614 (N2549, N2312, N2412);
  nand ginst615 (N2550, N2314, N2413);
  nand ginst616 (N2551, N2316, N2414);
  nand ginst617 (N2552, N2318, N2415);
  nand ginst618 (N2553, N2320, N2416);
  nand ginst619 (N2563, N2329, N2428);
  nand ginst620 (N2564, N2331, N2429);
  nand ginst621 (N2565, N2333, N2430);
  nand ginst622 (N2566, N2335, N2431);
  nand ginst623 (N2567, N2337, N2432);
  nand ginst624 (N2568, N2339, N2433);
  nand ginst625 (N2579, N1936, N2452);
  buf ginst626 (N2603, N2359);
  and ginst627 (N2607, N1880, N2377);
  and ginst628 (N2608, N1676, N2377);
  and ginst629 (N2609, N1681, N2377);
  and ginst630 (N2610, N1891, N2377);
  and ginst631 (N2611, N1856, N2382);
  and ginst632 (N2612, N1863, N2382);
  nand ginst633 (N2613, N2503, N2504);
  not ginst634 (N2617, N2434);
  nand ginst635 (N2618, N2366, N2434);
  nand ginst636 (N2619, N2367, N2437);
  not ginst637 (N2620, N2437);
  not ginst638 (N2621, N2368);
  nand ginst639 (N2624, N2510, N2511);
  not ginst640 (N2628, N2454);
  nand ginst641 (N2629, N2374, N2454);
  not ginst642 (N2630, N2472);
  and ginst643 (N2631, N1856, N2391);
  and ginst644 (N2632, N1863, N2391);
  and ginst645 (N2633, N1880, N2395);
  and ginst646 (N2634, N1676, N2395);
  and ginst647 (N2635, N1681, N2395);
  and ginst648 (N2636, N1891, N2395);
  not ginst649 (N2638, N2382);
  buf ginst650 (N2643, N2521);
  buf ginst651 (N2644, N2521);
  not ginst652 (N2645, N2475);
  not ginst653 (N2646, N2391);
  nand ginst654 (N2652, N2400, N2528);
  not ginst655 (N2655, N2478);
  not ginst656 (N2656, N2481);
  buf ginst657 (N2659, N2359);
  not ginst658 (N2663, N2484);
  nand ginst659 (N2664, N2301, N2484);
  not ginst660 (N2665, N2553);
  not ginst661 (N2666, N2552);
  not ginst662 (N2667, N2551);
  not ginst663 (N2668, N2550);
  not ginst664 (N2669, N2549);
  not ginst665 (N2670, N2548);
  not ginst666 (N2671, N2547);
  not ginst667 (N2672, N2546);
  not ginst668 (N2673, N2545);
  not ginst669 (N2674, N2544);
  not ginst670 (N2675, N2568);
  not ginst671 (N2676, N2567);
  not ginst672 (N2677, N2566);
  not ginst673 (N2678, N2565);
  not ginst674 (N2679, N2564);
  not ginst675 (N2680, N2563);
  not ginst676 (N2681, N2417);
  not ginst677 (N2684, N2421);
  buf ginst678 (N2687, N2425);
  buf ginst679 (N2690, N2425);
  not ginst680 (N2693, N2493);
  nand ginst681 (N2694, N1807, N2493);
  not ginst682 (N2695, N2440);
  not ginst683 (N2696, N2443);
  not ginst684 (N2697, N2446);
  not ginst685 (N2698, N2449);
  not ginst686 (N2699, N2457);
  not ginst687 (N2700, N2460);
  not ginst688 (N2701, N2463);
  not ginst689 (N2702, N2466);
  nand ginst690 (N2703, N2453, N2579);
  not ginst691 (N2706, N2469);
  not ginst692 (N2707, N2487);
  not ginst693 (N2708, N2490);
  and ginst694 (N2709, N2294, N2534);
  and ginst695 (N2710, N2291, N2531);
  nand ginst696 (N2719, N2191, N2617);
  nand ginst697 (N2720, N2194, N2620);
  nand ginst698 (N2726, N2207, N2628);
  buf ginst699 (N2729, N2537);
  buf ginst700 (N2738, N2537);
  not ginst701 (N2743, N2652);
  nand ginst702 (N2747, N2049, N2663);
  and ginst703 (N2748, N2665, N2666, N2667, N2668, N2669);
  and ginst704 (N2749, N2670, N2671, N2672, N2673, N2674);
  and ginst705 (N2750, N2034, N2675);
  and ginst706 (N2751, N2676, N2677, N2678, N2679, N2680);
  nand ginst707 (N2760, N1588, N2693);
  buf ginst708 (N2761, N2540);
  buf ginst709 (N2766, N2540);
  nand ginst710 (N2771, N2443, N2695);
  nand ginst711 (N2772, N2440, N2696);
  nand ginst712 (N2773, N2449, N2697);
  nand ginst713 (N2774, N2446, N2698);
  nand ginst714 (N2775, N2460, N2699);
  nand ginst715 (N2776, N2457, N2700);
  nand ginst716 (N2777, N2466, N2701);
  nand ginst717 (N2778, N2463, N2702);
  nand ginst718 (N2781, N2490, N2707);
  nand ginst719 (N2782, N2487, N2708);
  or ginst720 (N2783, N2534, N2709);
  or ginst721 (N2784, N2531, N2710);
  and ginst722 (N2789, N1856, N2638);
  and ginst723 (N2790, N1863, N2638);
  and ginst724 (N2791, N1870, N2638);
  and ginst725 (N2792, N1875, N2638);
  not ginst726 (N2793, N2613);
  nand ginst727 (N2796, N2618, N2719);
  nand ginst728 (N2800, N2619, N2720);
  not ginst729 (N2803, N2624);
  nand ginst730 (N2806, N2629, N2726);
  and ginst731 (N2809, N1856, N2646);
  and ginst732 (N2810, N1863, N2646);
  and ginst733 (N2811, N1870, N2646);
  and ginst734 (N2812, N1875, N2646);
  and ginst735 (N2817, N14, N2743);
  buf ginst736 (N2820, N2603);
  nand ginst737 (N2826, N2664, N2747);
  and ginst738 (N2829, N2748, N2749);
  and ginst739 (N2830, N2750, N2751);
  buf ginst740 (N2831, N2659);
  not ginst741 (N2837, N2687);
  not ginst742 (N2838, N2690);
  and ginst743 (N2839, N2417, N2421, N2687);
  and ginst744 (N2840, N2681, N2684, N2690);
  nand ginst745 (N2841, N2694, N2760);
  buf ginst746 (N2844, N2603);
  buf ginst747 (N2854, N2603);
  buf ginst748 (N2859, N2659);
  buf ginst749 (N2869, N2659);
  nand ginst750 (N2874, N2773, N2774);
  nand ginst751 (N2877, N2771, N2772);
  not ginst752 (N2880, N2703);
  nand ginst753 (N2881, N2703, N2706);
  nand ginst754 (N2882, N2777, N2778);
  nand ginst755 (N2885, N2775, N2776);
  nand ginst756 (N2888, N2781, N2782);
  nand ginst757 (N2891, N2783, N2784);
  and ginst758 (N2894, N2607, N2729);
  and ginst759 (N2895, N2608, N2729);
  and ginst760 (N2896, N2609, N2729);
  and ginst761 (N2897, N2610, N2729);
  or ginst762 (N2898, N2611, N2789);
  or ginst763 (N2899, N2612, N2790);
  and ginst764 (N2900, N1037, N2791);
  and ginst765 (N2901, N1037, N2792);
  or ginst766 (N2914, N2631, N2809);
  or ginst767 (N2915, N2632, N2810);
  and ginst768 (N2916, N1070, N2811);
  and ginst769 (N2917, N1070, N2812);
  and ginst770 (N2918, N2633, N2738);
  and ginst771 (N2919, N2634, N2738);
  and ginst772 (N2920, N2635, N2738);
  and ginst773 (N2921, N2636, N2738);
  buf ginst774 (N2925, N2817);
  and ginst775 (N2931, N1302, N2829, N2830);
  and ginst776 (N2938, N2421, N2681, N2837);
  and ginst777 (N2939, N2417, N2684, N2838);
  nand ginst778 (N2963, N2469, N2880);
  not ginst779 (N2970, N2841);
  not ginst780 (N2971, N2826);
  not ginst781 (N2972, N2894);
  not ginst782 (N2975, N2895);
  not ginst783 (N2978, N2896);
  not ginst784 (N2981, N2897);
  and ginst785 (N2984, N1037, N2898);
  and ginst786 (N2985, N1037, N2899);
  not ginst787 (N2986, N2900);
  not ginst788 (N2989, N2901);
  not ginst789 (N2992, N2796);
  buf ginst790 (N2995, N2800);
  buf ginst791 (N2998, N2800);
  buf ginst792 (N3001, N2806);
  buf ginst793 (N3004, N2806);
  and ginst794 (N3007, N2820, N574);
  and ginst795 (N3008, N1070, N2914);
  and ginst796 (N3009, N1070, N2915);
  not ginst797 (N3010, N2916);
  not ginst798 (N3013, N2917);
  not ginst799 (N3016, N2918);
  not ginst800 (N3019, N2919);
  not ginst801 (N3022, N2920);
  not ginst802 (N3025, N2921);
  not ginst803 (N3028, N2817);
  and ginst804 (N3029, N2831, N574);
  not ginst805 (N3030, N2820);
  and ginst806 (N3035, N2820, N578);
  and ginst807 (N3036, N2820, N655);
  and ginst808 (N3037, N2820, N659);
  buf ginst809 (N3038, N2931);
  not ginst810 (N3039, N2831);
  and ginst811 (N3044, N2831, N578);
  and ginst812 (N3045, N2831, N655);
  and ginst813 (N3046, N2831, N659);
  nor ginst814 (N3047, N2839, N2938);
  nor ginst815 (N3048, N2840, N2939);
  not ginst816 (N3049, N2888);
  not ginst817 (N3050, N2844);
  and ginst818 (N3053, N2844, N663);
  and ginst819 (N3054, N2844, N667);
  and ginst820 (N3055, N2844, N671);
  and ginst821 (N3056, N2844, N675);
  and ginst822 (N3057, N2854, N679);
  and ginst823 (N3058, N2854, N683);
  and ginst824 (N3059, N2854, N687);
  and ginst825 (N3060, N2854, N705);
  not ginst826 (N3061, N2859);
  and ginst827 (N3064, N2859, N663);
  and ginst828 (N3065, N2859, N667);
  and ginst829 (N3066, N2859, N671);
  and ginst830 (N3067, N2859, N675);
  and ginst831 (N3068, N2869, N679);
  and ginst832 (N3069, N2869, N683);
  and ginst833 (N3070, N2869, N687);
  and ginst834 (N3071, N2869, N705);
  not ginst835 (N3072, N2874);
  not ginst836 (N3073, N2877);
  not ginst837 (N3074, N2882);
  not ginst838 (N3075, N2885);
  nand ginst839 (N3076, N2881, N2963);
  not ginst840 (N3079, N2931);
  not ginst841 (N3088, N2984);
  not ginst842 (N3091, N2985);
  not ginst843 (N3110, N3008);
  not ginst844 (N3113, N3009);
  and ginst845 (N3137, N1190, N3055);
  and ginst846 (N3140, N1190, N3056);
  and ginst847 (N3143, N2761, N3057);
  and ginst848 (N3146, N2761, N3058);
  and ginst849 (N3149, N2761, N3059);
  and ginst850 (N3152, N2761, N3060);
  and ginst851 (N3157, N1195, N3066);
  and ginst852 (N3160, N1195, N3067);
  and ginst853 (N3163, N2766, N3068);
  and ginst854 (N3166, N2766, N3069);
  and ginst855 (N3169, N2766, N3070);
  and ginst856 (N3172, N2766, N3071);
  nand ginst857 (N3175, N2877, N3072);
  nand ginst858 (N3176, N2874, N3073);
  nand ginst859 (N3177, N2885, N3074);
  nand ginst860 (N3178, N2882, N3075);
  nand ginst861 (N3180, N3047, N3048);
  not ginst862 (N3187, N2995);
  not ginst863 (N3188, N2998);
  not ginst864 (N3189, N3001);
  not ginst865 (N3190, N3004);
  and ginst866 (N3191, N2613, N2796, N2995);
  and ginst867 (N3192, N2793, N2992, N2998);
  and ginst868 (N3193, N2368, N2624, N3001);
  and ginst869 (N3194, N2621, N2803, N3004);
  nand ginst870 (N3195, N2375, N3076);
  not ginst871 (N3196, N3076);
  and ginst872 (N3197, N3030, N687);
  and ginst873 (N3208, N3039, N687);
  and ginst874 (N3215, N3030, N705);
  and ginst875 (N3216, N3030, N711);
  and ginst876 (N3217, N3030, N715);
  and ginst877 (N3218, N3039, N705);
  and ginst878 (N3219, N3039, N711);
  and ginst879 (N3220, N3039, N715);
  and ginst880 (N3222, N3050, N719);
  and ginst881 (N3223, N3050, N723);
  and ginst882 (N3230, N3061, N719);
  and ginst883 (N3231, N3061, N723);
  nand ginst884 (N3238, N3175, N3176);
  nand ginst885 (N3241, N3177, N3178);
  buf ginst886 (N3244, N2981);
  buf ginst887 (N3247, N2978);
  buf ginst888 (N3250, N2975);
  buf ginst889 (N3253, N2972);
  buf ginst890 (N3256, N2989);
  buf ginst891 (N3259, N2986);
  buf ginst892 (N3262, N3025);
  buf ginst893 (N3265, N3022);
  buf ginst894 (N3268, N3019);
  buf ginst895 (N3271, N3016);
  buf ginst896 (N3274, N3013);
  buf ginst897 (N3277, N3010);
  and ginst898 (N3281, N2793, N2796, N3187);
  and ginst899 (N3282, N2613, N2992, N3188);
  and ginst900 (N3283, N2621, N2624, N3189);
  and ginst901 (N3284, N2368, N2803, N3190);
  nand ginst902 (N3286, N2210, N3196);
  or ginst903 (N3288, N3007, N3197);
  nand ginst904 (N3289, N3049, N3180);
  and ginst905 (N3291, N2981, N3152);
  and ginst906 (N3293, N2978, N3149);
  and ginst907 (N3295, N2975, N3146);
  and ginst908 (N3296, N2972, N3143);
  and ginst909 (N3299, N2989, N3140);
  and ginst910 (N3301, N2986, N3137);
  or ginst911 (N3302, N3029, N3208);
  and ginst912 (N3304, N3025, N3172);
  and ginst913 (N3306, N3022, N3169);
  and ginst914 (N3308, N3019, N3166);
  and ginst915 (N3309, N3016, N3163);
  and ginst916 (N3312, N3013, N3160);
  and ginst917 (N3314, N3010, N3157);
  or ginst918 (N3315, N3035, N3215);
  or ginst919 (N3318, N3036, N3216);
  or ginst920 (N3321, N3037, N3217);
  or ginst921 (N3324, N3044, N3218);
  or ginst922 (N3327, N3045, N3219);
  or ginst923 (N3330, N3046, N3220);
  not ginst924 (N3333, N3180);
  or ginst925 (N3334, N3053, N3222);
  or ginst926 (N3335, N3054, N3223);
  or ginst927 (N3336, N3064, N3230);
  or ginst928 (N3337, N3065, N3231);
  buf ginst929 (N3340, N3152);
  buf ginst930 (N3344, N3149);
  buf ginst931 (N3348, N3146);
  buf ginst932 (N3352, N3143);
  buf ginst933 (N3356, N3140);
  buf ginst934 (N3360, N3137);
  buf ginst935 (N3364, N3091);
  buf ginst936 (N3367, N3088);
  buf ginst937 (N3370, N3172);
  buf ginst938 (N3374, N3169);
  buf ginst939 (N3378, N3166);
  buf ginst940 (N3382, N3163);
  buf ginst941 (N3386, N3160);
  buf ginst942 (N3390, N3157);
  buf ginst943 (N3394, N3113);
  buf ginst944 (N3397, N3110);
  nand ginst945 (N3400, N3195, N3286);
  nor ginst946 (N3401, N3191, N3281);
  nor ginst947 (N3402, N3192, N3282);
  nor ginst948 (N3403, N3193, N3283);
  nor ginst949 (N3404, N3194, N3284);
  not ginst950 (N3405, N3238);
  not ginst951 (N3406, N3241);
  and ginst952 (N3409, N1836, N3288);
  nand ginst953 (N3410, N2888, N3333);
  not ginst954 (N3412, N3244);
  not ginst955 (N3414, N3247);
  not ginst956 (N3416, N3250);
  not ginst957 (N3418, N3253);
  not ginst958 (N3420, N3256);
  not ginst959 (N3422, N3259);
  and ginst960 (N3428, N1836, N3302);
  not ginst961 (N3430, N3262);
  not ginst962 (N3432, N3265);
  not ginst963 (N3434, N3268);
  not ginst964 (N3436, N3271);
  not ginst965 (N3438, N3274);
  not ginst966 (N3440, N3277);
  and ginst967 (N3450, N1190, N3334);
  and ginst968 (N3453, N1190, N3335);
  and ginst969 (N3456, N1195, N3336);
  and ginst970 (N3459, N1195, N3337);
  and ginst971 (N3478, N3400, N533);
  and ginst972 (N3479, N2128, N3318);
  and ginst973 (N3480, N1841, N3315);
  nand ginst974 (N3481, N3289, N3410);
  not ginst975 (N3482, N3340);
  nand ginst976 (N3483, N3340, N3412);
  not ginst977 (N3484, N3344);
  nand ginst978 (N3485, N3344, N3414);
  not ginst979 (N3486, N3348);
  nand ginst980 (N3487, N3348, N3416);
  not ginst981 (N3488, N3352);
  nand ginst982 (N3489, N3352, N3418);
  not ginst983 (N3490, N3356);
  nand ginst984 (N3491, N3356, N3420);
  not ginst985 (N3492, N3360);
  nand ginst986 (N3493, N3360, N3422);
  not ginst987 (N3494, N3364);
  not ginst988 (N3496, N3367);
  and ginst989 (N3498, N2135, N3321);
  and ginst990 (N3499, N2128, N3327);
  and ginst991 (N3500, N1841, N3324);
  not ginst992 (N3501, N3370);
  nand ginst993 (N3502, N3370, N3430);
  not ginst994 (N3503, N3374);
  nand ginst995 (N3504, N3374, N3432);
  not ginst996 (N3505, N3378);
  nand ginst997 (N3506, N3378, N3434);
  not ginst998 (N3507, N3382);
  nand ginst999 (N3508, N3382, N3436);
  not ginst1000 (N3509, N3386);
  nand ginst1001 (N3510, N3386, N3438);
  not ginst1002 (N3511, N3390);
  nand ginst1003 (N3512, N3390, N3440);
  not ginst1004 (N3513, N3394);
  not ginst1005 (N3515, N3397);
  and ginst1006 (N3517, N2135, N3330);
  nand ginst1007 (N3522, N3401, N3402);
  nand ginst1008 (N3525, N3403, N3404);
  buf ginst1009 (N3528, N3318);
  buf ginst1010 (N3531, N3315);
  buf ginst1011 (N3534, N3321);
  buf ginst1012 (N3537, N3327);
  buf ginst1013 (N3540, N3324);
  buf ginst1014 (N3543, N3330);
  or ginst1015 (N3546, N1813, N3478);
  not ginst1016 (N3551, N3481);
  nand ginst1017 (N3552, N3244, N3482);
  nand ginst1018 (N3553, N3247, N3484);
  nand ginst1019 (N3554, N3250, N3486);
  nand ginst1020 (N3555, N3253, N3488);
  nand ginst1021 (N3556, N3256, N3490);
  nand ginst1022 (N3557, N3259, N3492);
  and ginst1023 (N3558, N3091, N3453);
  and ginst1024 (N3559, N3088, N3450);
  nand ginst1025 (N3563, N3262, N3501);
  nand ginst1026 (N3564, N3265, N3503);
  nand ginst1027 (N3565, N3268, N3505);
  nand ginst1028 (N3566, N3271, N3507);
  nand ginst1029 (N3567, N3274, N3509);
  nand ginst1030 (N3568, N3277, N3511);
  and ginst1031 (N3569, N3113, N3459);
  and ginst1032 (N3570, N3110, N3456);
  buf ginst1033 (N3576, N3453);
  buf ginst1034 (N3579, N3450);
  buf ginst1035 (N3585, N3459);
  buf ginst1036 (N3588, N3456);
  not ginst1037 (N3592, N3522);
  nand ginst1038 (N3593, N3405, N3522);
  not ginst1039 (N3594, N3525);
  nand ginst1040 (N3595, N3406, N3525);
  not ginst1041 (N3596, N3528);
  nand ginst1042 (N3597, N2630, N3528);
  nand ginst1043 (N3598, N2376, N3531);
  not ginst1044 (N3599, N3531);
  and ginst1045 (N3600, N3551, N800);
  nand ginst1046 (N3603, N3483, N3552);
  nand ginst1047 (N3608, N3485, N3553);
  nand ginst1048 (N3612, N3487, N3554);
  nand ginst1049 (N3615, N3489, N3555);
  nand ginst1050 (N3616, N3491, N3556);
  nand ginst1051 (N3622, N3493, N3557);
  not ginst1052 (N3629, N3534);
  nand ginst1053 (N3630, N2645, N3534);
  not ginst1054 (N3631, N3537);
  nand ginst1055 (N3632, N2655, N3537);
  nand ginst1056 (N3633, N2403, N3540);
  not ginst1057 (N3634, N3540);
  nand ginst1058 (N3635, N3502, N3563);
  nand ginst1059 (N3640, N3504, N3564);
  nand ginst1060 (N3644, N3506, N3565);
  nand ginst1061 (N3647, N3508, N3566);
  nand ginst1062 (N3648, N3510, N3567);
  nand ginst1063 (N3654, N3512, N3568);
  not ginst1064 (N3661, N3543);
  nand ginst1065 (N3662, N2656, N3543);
  nand ginst1066 (N3667, N3238, N3592);
  nand ginst1067 (N3668, N3241, N3594);
  nand ginst1068 (N3669, N2472, N3596);
  nand ginst1069 (N3670, N2213, N3599);
  buf ginst1070 (N3671, N3600);
  not ginst1071 (N3691, N3576);
  nand ginst1072 (N3692, N3494, N3576);
  not ginst1073 (N3693, N3579);
  nand ginst1074 (N3694, N3496, N3579);
  nand ginst1075 (N3695, N2475, N3629);
  nand ginst1076 (N3696, N2478, N3631);
  nand ginst1077 (N3697, N2216, N3634);
  not ginst1078 (N3716, N3585);
  nand ginst1079 (N3717, N3513, N3585);
  not ginst1080 (N3718, N3588);
  nand ginst1081 (N3719, N3515, N3588);
  nand ginst1082 (N3720, N2481, N3661);
  nand ginst1083 (N3721, N3593, N3667);
  nand ginst1084 (N3722, N3595, N3668);
  nand ginst1085 (N3723, N3597, N3669);
  nand ginst1086 (N3726, N3598, N3670);
  not ginst1087 (N3727, N3600);
  nand ginst1088 (N3728, N3364, N3691);
  nand ginst1089 (N3729, N3367, N3693);
  nand ginst1090 (N3730, N3630, N3695);
  and ginst1091 (N3731, N3603, N3608, N3612, N3615);
  and ginst1092 (N3732, N3293, N3603);
  and ginst1093 (N3733, N3295, N3603, N3608);
  and ginst1094 (N3734, N3296, N3603, N3608, N3612);
  and ginst1095 (N3735, N3301, N3616);
  and ginst1096 (N3736, N3558, N3616, N3622);
  nand ginst1097 (N3737, N3632, N3696);
  nand ginst1098 (N3740, N3633, N3697);
  nand ginst1099 (N3741, N3394, N3716);
  nand ginst1100 (N3742, N3397, N3718);
  nand ginst1101 (N3743, N3662, N3720);
  and ginst1102 (N3744, N3635, N3640, N3644, N3647);
  and ginst1103 (N3745, N3306, N3635);
  and ginst1104 (N3746, N3308, N3635, N3640);
  and ginst1105 (N3747, N3309, N3635, N3640, N3644);
  and ginst1106 (N3748, N3314, N3648);
  and ginst1107 (N3749, N3569, N3648, N3654);
  not ginst1108 (N3750, N3721);
  and ginst1109 (N3753, N246, N3722);
  nand ginst1110 (N3754, N3692, N3728);
  nand ginst1111 (N3758, N3694, N3729);
  not ginst1112 (N3761, N3731);
  or ginst1113 (N3762, N3291, N3732, N3733, N3734);
  nand ginst1114 (N3767, N3717, N3741);
  nand ginst1115 (N3771, N3719, N3742);
  not ginst1116 (N3774, N3744);
  or ginst1117 (N3775, N3304, N3745, N3746, N3747);
  and ginst1118 (N3778, N3480, N3723);
  and ginst1119 (N3779, N3409, N3723, N3726);
  or ginst1120 (N3780, N2125, N3753);
  and ginst1121 (N3790, N3750, N800);
  and ginst1122 (N3793, N3500, N3737);
  and ginst1123 (N3794, N3428, N3737, N3740);
  or ginst1124 (N3802, N3479, N3778, N3779);
  buf ginst1125 (N3803, N3780);
  buf ginst1126 (N3804, N3780);
  not ginst1127 (N3805, N3762);
  and ginst1128 (N3806, N3616, N3622, N3730, N3754, N3758);
  and ginst1129 (N3807, N3559, N3616, N3622, N3754);
  and ginst1130 (N3808, N3498, N3616, N3622, N3754, N3758);
  buf ginst1131 (N3809, N3790);
  or ginst1132 (N3811, N3499, N3793, N3794);
  not ginst1133 (N3812, N3775);
  and ginst1134 (N3813, N3648, N3654, N3743, N3767, N3771);
  and ginst1135 (N3814, N3570, N3648, N3654, N3767);
  and ginst1136 (N3815, N3517, N3648, N3654, N3767, N3771);
  or ginst1137 (N3816, N3299, N3735, N3736, N3807, N3808);
  and ginst1138 (N3817, N3802, N3806);
  nand ginst1139 (N3818, N3761, N3805);
  not ginst1140 (N3819, N3790);
  or ginst1141 (N3820, N3312, N3748, N3749, N3814, N3815);
  and ginst1142 (N3821, N3811, N3813);
  nand ginst1143 (N3822, N3774, N3812);
  or ginst1144 (N3823, N3816, N3817);
  and ginst1145 (N3826, N2841, N3727, N3819);
  or ginst1146 (N3827, N3820, N3821);
  not ginst1147 (N3834, N3823);
  and ginst1148 (N3835, N3818, N3823);
  not ginst1149 (N3836, N3827);
  and ginst1150 (N3837, N3822, N3827);
  and ginst1151 (N3838, N3762, N3834);
  and ginst1152 (N3839, N3775, N3836);
  or ginst1153 (N3840, N3835, N3838);
  or ginst1154 (N3843, N3837, N3839);
  buf ginst1155 (N3851, N3843);
  nand ginst1156 (N3852, N3840, N3843);
  and ginst1157 (N3857, N3843, N3852);
  and ginst1158 (N3858, N3840, N3852);
  or ginst1159 (N3859, N3857, N3858);
  not ginst1160 (N3864, N3859);
  and ginst1161 (N3869, N3859, N3864);
  or ginst1162 (N3870, N3864, N3869);
  not ginst1163 (N3875, N3870);
  and ginst1164 (N3876, N2826, N3028, N3870);
  and ginst1165 (N3877, N1591, N3826, N3876);
  buf ginst1166 (N3881, N3877);
  not ginst1167 (N3882, N3877);
  buf ginst1168 (N398, N219);
  buf ginst1169 (N400, N219);
  buf ginst1170 (N401, N219);
  and ginst1171 (N405, N1, N3);
  not ginst1172 (N408, N230);
  buf ginst1173 (N419, N253);
  buf ginst1174 (N420, N253);
  not ginst1175 (N425, N262);
  buf ginst1176 (N456, N290);
  buf ginst1177 (N457, N290);
  buf ginst1178 (N458, N290);
  and ginst1179 (N485, N297, N301, N305, N309);
  not ginst1180 (N486, N405);
  not ginst1181 (N487, N44);
  not ginst1182 (N488, N132);
  not ginst1183 (N489, N82);
  not ginst1184 (N490, N96);
  not ginst1185 (N491, N69);
  not ginst1186 (N492, N120);
  not ginst1187 (N493, N57);
  not ginst1188 (N494, N108);
  and ginst1189 (N495, N2, N15, N237);
  buf ginst1190 (N496, N237);
  and ginst1191 (N499, N37, N37);
  buf ginst1192 (N500, N219);
  buf ginst1193 (N503, N8);
  buf ginst1194 (N506, N8);
  buf ginst1195 (N509, N227);
  buf ginst1196 (N521, N234);
  not ginst1197 (N533, N241);
  not ginst1198 (N537, N246);
  and ginst1199 (N543, N11, N246);
  and ginst1200 (N544, N44, N82, N96, N132);
  and ginst1201 (N547, N57, N69, N108, N120);
  buf ginst1202 (N550, N227);
  buf ginst1203 (N562, N234);
  not ginst1204 (N574, N256);
  not ginst1205 (N578, N259);
  buf ginst1206 (N582, N319);
  buf ginst1207 (N594, N322);
  not ginst1208 (N606, N328);
  not ginst1209 (N607, N331);
  not ginst1210 (N608, N334);
  not ginst1211 (N609, N337);
  not ginst1212 (N610, N340);
  not ginst1213 (N611, N343);
  not ginst1214 (N612, N352);
  buf ginst1215 (N613, N319);
  buf ginst1216 (N625, N322);
  buf ginst1217 (N637, N16);
  buf ginst1218 (N643, N16);
  not ginst1219 (N650, N355);
  and ginst1220 (N651, N7, N237);
  not ginst1221 (N655, N263);
  not ginst1222 (N659, N266);
  not ginst1223 (N663, N269);
  not ginst1224 (N667, N272);
  not ginst1225 (N671, N275);
  not ginst1226 (N675, N278);
  not ginst1227 (N679, N281);
  not ginst1228 (N683, N284);
  not ginst1229 (N687, N287);
  buf ginst1230 (N693, N29);
  buf ginst1231 (N699, N29);
  not ginst1232 (N705, N294);
  not ginst1233 (N711, N297);
  not ginst1234 (N715, N301);
  not ginst1235 (N719, N305);
  not ginst1236 (N723, N309);
  not ginst1237 (N727, N313);
  not ginst1238 (N730, N316);
  not ginst1239 (N733, N346);
  not ginst1240 (N734, N349);
  buf ginst1241 (N735, N259);
  buf ginst1242 (N738, N256);
  buf ginst1243 (N741, N263);
  buf ginst1244 (N744, N269);
  buf ginst1245 (N747, N266);
  buf ginst1246 (N750, N275);
  buf ginst1247 (N753, N272);
  buf ginst1248 (N756, N281);
  buf ginst1249 (N759, N278);
  buf ginst1250 (N762, N287);
  buf ginst1251 (N765, N284);
  buf ginst1252 (N768, N294);
  buf ginst1253 (N771, N301);
  buf ginst1254 (N774, N297);
  buf ginst1255 (N777, N309);
  buf ginst1256 (N780, N305);
  buf ginst1257 (N783, N316);
  buf ginst1258 (N786, N313);
  not ginst1259 (N792, N485);
  not ginst1260 (N799, N495);
  not ginst1261 (N800, N499);
  buf ginst1262 (N805, N500);
  nand ginst1263 (N900, N331, N606);
  nand ginst1264 (N901, N328, N607);
  nand ginst1265 (N902, N337, N608);
  nand ginst1266 (N903, N334, N609);
  nand ginst1267 (N904, N343, N610);
  nand ginst1268 (N905, N340, N611);
  nand ginst1269 (N998, N349, N733);
  nand ginst1270 (N999, N346, N734);

endmodule

/*************** SatHard block ***************/
module SatHard (N96, N231, N82, N120, keyinput0, keyinput1, keyinput2, keyinput3, keyinput4, keyinput5, keyinput6, keyinput7, flip_signal);

  input N96, N231, N82, N120, keyinput0, keyinput1, keyinput2, keyinput3, keyinput4, keyinput5, keyinput6, keyinput7;
  output flip_signal;
  //SatHard key=10010100
  wire [3:0] sat_res_inputs;
  wire [7:0] keyinputs, keyvalue;
  assign sat_res_inputs[3:0] = {N96, N231, N82, N120};
  assign keyinputs[7:0] = {keyinput0, keyinput1, keyinput2, keyinput3, keyinput4, keyinput5, keyinput6, keyinput7};
  assign keyvalue[7:0] = 8'b10010100;

  wire g, g_bar;
  assign g = &(keyinputs[3:0] ^ sat_res_inputs ^ keyvalue[3:0]);
  assign g_bar = ~&(keyinputs[7:4] ^ sat_res_inputs ^ keyvalue[7:4]);
  assign flip_signal = g & g_bar;

endmodule
/*************** SatHard block ***************/
