//key=0011110010011111110011011101100011100110100000110010100100111110
// Main module
module b14_C_AntiSAT_64_0(WR_REG_SCAN_IN, DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, DATAI_27_, DATAI_26_, DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, DATAI_21_, DATAI_20_, DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, DATAI_15_, DATAI_14_, DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, DATAI_9_, DATAI_8_, DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, DATAI_2_, DATAI_1_, DATAI_0_, RD_REG_SCAN_IN, STATE_REG_SCAN_IN, REG3_REG_7__SCAN_IN, REG3_REG_27__SCAN_IN, REG3_REG_14__SCAN_IN, REG3_REG_23__SCAN_IN, REG3_REG_10__SCAN_IN, REG3_REG_3__SCAN_IN, REG3_REG_19__SCAN_IN, REG3_REG_28__SCAN_IN, REG3_REG_8__SCAN_IN, REG3_REG_1__SCAN_IN, REG3_REG_21__SCAN_IN, REG3_REG_12__SCAN_IN, REG3_REG_25__SCAN_IN, REG3_REG_16__SCAN_IN, REG3_REG_5__SCAN_IN, REG3_REG_17__SCAN_IN, REG3_REG_24__SCAN_IN, REG3_REG_4__SCAN_IN, REG3_REG_9__SCAN_IN, REG3_REG_0__SCAN_IN, REG3_REG_20__SCAN_IN, REG3_REG_13__SCAN_IN, IR_REG_0__SCAN_IN, IR_REG_1__SCAN_IN, IR_REG_2__SCAN_IN, IR_REG_3__SCAN_IN, IR_REG_4__SCAN_IN, IR_REG_5__SCAN_IN, IR_REG_6__SCAN_IN, IR_REG_7__SCAN_IN, IR_REG_8__SCAN_IN, IR_REG_9__SCAN_IN, IR_REG_10__SCAN_IN, IR_REG_11__SCAN_IN, IR_REG_12__SCAN_IN, IR_REG_13__SCAN_IN, IR_REG_14__SCAN_IN, IR_REG_15__SCAN_IN, IR_REG_16__SCAN_IN, IR_REG_17__SCAN_IN, IR_REG_18__SCAN_IN, IR_REG_19__SCAN_IN, IR_REG_20__SCAN_IN, IR_REG_21__SCAN_IN, IR_REG_22__SCAN_IN, IR_REG_23__SCAN_IN, IR_REG_24__SCAN_IN, IR_REG_25__SCAN_IN, IR_REG_26__SCAN_IN, IR_REG_27__SCAN_IN, IR_REG_28__SCAN_IN, IR_REG_29__SCAN_IN, IR_REG_30__SCAN_IN, IR_REG_31__SCAN_IN, D_REG_0__SCAN_IN, D_REG_1__SCAN_IN, D_REG_2__SCAN_IN, D_REG_3__SCAN_IN, D_REG_4__SCAN_IN, D_REG_5__SCAN_IN, D_REG_6__SCAN_IN, D_REG_7__SCAN_IN, D_REG_8__SCAN_IN, D_REG_9__SCAN_IN, D_REG_10__SCAN_IN, D_REG_11__SCAN_IN, D_REG_12__SCAN_IN, D_REG_13__SCAN_IN, D_REG_14__SCAN_IN, D_REG_15__SCAN_IN, D_REG_16__SCAN_IN, D_REG_17__SCAN_IN, D_REG_18__SCAN_IN, D_REG_19__SCAN_IN, D_REG_20__SCAN_IN, D_REG_21__SCAN_IN, D_REG_22__SCAN_IN, D_REG_23__SCAN_IN, D_REG_24__SCAN_IN, D_REG_25__SCAN_IN, D_REG_26__SCAN_IN, D_REG_27__SCAN_IN, D_REG_28__SCAN_IN, D_REG_29__SCAN_IN, D_REG_30__SCAN_IN, D_REG_31__SCAN_IN, REG0_REG_0__SCAN_IN, REG0_REG_1__SCAN_IN, REG0_REG_2__SCAN_IN, REG0_REG_3__SCAN_IN, REG0_REG_4__SCAN_IN, REG0_REG_5__SCAN_IN, REG0_REG_6__SCAN_IN, REG0_REG_7__SCAN_IN, REG0_REG_8__SCAN_IN, REG0_REG_9__SCAN_IN, REG0_REG_10__SCAN_IN, REG0_REG_11__SCAN_IN, REG0_REG_12__SCAN_IN, REG0_REG_13__SCAN_IN, REG0_REG_14__SCAN_IN, REG0_REG_15__SCAN_IN, REG0_REG_16__SCAN_IN, REG0_REG_17__SCAN_IN, REG0_REG_18__SCAN_IN, REG0_REG_19__SCAN_IN, REG0_REG_20__SCAN_IN, REG0_REG_21__SCAN_IN, REG0_REG_22__SCAN_IN, REG0_REG_23__SCAN_IN, REG0_REG_24__SCAN_IN, REG0_REG_25__SCAN_IN, REG0_REG_26__SCAN_IN, REG0_REG_27__SCAN_IN, REG0_REG_28__SCAN_IN, REG0_REG_29__SCAN_IN, REG0_REG_30__SCAN_IN, REG0_REG_31__SCAN_IN, REG1_REG_0__SCAN_IN, REG1_REG_1__SCAN_IN, REG1_REG_2__SCAN_IN, REG1_REG_3__SCAN_IN, REG1_REG_4__SCAN_IN, REG1_REG_5__SCAN_IN, REG1_REG_6__SCAN_IN, REG1_REG_7__SCAN_IN, REG1_REG_8__SCAN_IN, REG1_REG_9__SCAN_IN, REG1_REG_10__SCAN_IN, REG1_REG_11__SCAN_IN, REG1_REG_12__SCAN_IN, REG1_REG_13__SCAN_IN, REG1_REG_14__SCAN_IN, REG1_REG_15__SCAN_IN, REG1_REG_16__SCAN_IN, REG1_REG_17__SCAN_IN, REG1_REG_18__SCAN_IN, REG1_REG_19__SCAN_IN, REG1_REG_20__SCAN_IN, REG1_REG_21__SCAN_IN, REG1_REG_22__SCAN_IN, REG1_REG_23__SCAN_IN, REG1_REG_24__SCAN_IN, REG1_REG_25__SCAN_IN, REG1_REG_26__SCAN_IN, REG1_REG_27__SCAN_IN, REG1_REG_28__SCAN_IN, REG1_REG_29__SCAN_IN, REG1_REG_30__SCAN_IN, REG1_REG_31__SCAN_IN, REG2_REG_0__SCAN_IN, REG2_REG_1__SCAN_IN, REG2_REG_2__SCAN_IN, REG2_REG_3__SCAN_IN, REG2_REG_4__SCAN_IN, REG2_REG_5__SCAN_IN, REG2_REG_6__SCAN_IN, REG2_REG_7__SCAN_IN, REG2_REG_8__SCAN_IN, REG2_REG_9__SCAN_IN, REG2_REG_10__SCAN_IN, REG2_REG_11__SCAN_IN, REG2_REG_12__SCAN_IN, REG2_REG_13__SCAN_IN, REG2_REG_14__SCAN_IN, REG2_REG_15__SCAN_IN, REG2_REG_16__SCAN_IN, REG2_REG_17__SCAN_IN, REG2_REG_18__SCAN_IN, REG2_REG_19__SCAN_IN, REG2_REG_20__SCAN_IN, REG2_REG_21__SCAN_IN, REG2_REG_22__SCAN_IN, REG2_REG_23__SCAN_IN, REG2_REG_24__SCAN_IN, REG2_REG_25__SCAN_IN, REG2_REG_26__SCAN_IN, REG2_REG_27__SCAN_IN, REG2_REG_28__SCAN_IN, REG2_REG_29__SCAN_IN, REG2_REG_30__SCAN_IN, REG2_REG_31__SCAN_IN, ADDR_REG_19__SCAN_IN, ADDR_REG_18__SCAN_IN, ADDR_REG_17__SCAN_IN, ADDR_REG_16__SCAN_IN, ADDR_REG_15__SCAN_IN, ADDR_REG_14__SCAN_IN, ADDR_REG_13__SCAN_IN, ADDR_REG_12__SCAN_IN, ADDR_REG_11__SCAN_IN, ADDR_REG_10__SCAN_IN, ADDR_REG_9__SCAN_IN, ADDR_REG_8__SCAN_IN, ADDR_REG_7__SCAN_IN, ADDR_REG_6__SCAN_IN, ADDR_REG_5__SCAN_IN, ADDR_REG_4__SCAN_IN, ADDR_REG_3__SCAN_IN, ADDR_REG_2__SCAN_IN, ADDR_REG_1__SCAN_IN, ADDR_REG_0__SCAN_IN, DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN, DATAO_REG_2__SCAN_IN, DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN, DATAO_REG_5__SCAN_IN, DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN, DATAO_REG_8__SCAN_IN, DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN, DATAO_REG_11__SCAN_IN, DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN, DATAO_REG_14__SCAN_IN, DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN, DATAO_REG_17__SCAN_IN, DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN, DATAO_REG_20__SCAN_IN, DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN, DATAO_REG_23__SCAN_IN, DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN, DATAO_REG_26__SCAN_IN, DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN, DATAO_REG_29__SCAN_IN, DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN, B_REG_SCAN_IN, REG3_REG_15__SCAN_IN, REG3_REG_26__SCAN_IN, REG3_REG_6__SCAN_IN, REG3_REG_18__SCAN_IN, REG3_REG_2__SCAN_IN, REG3_REG_11__SCAN_IN, REG3_REG_22__SCAN_IN, keyinput0, keyinput1, keyinput2, keyinput3, keyinput4, keyinput5, keyinput6, keyinput7, keyinput8, keyinput9, keyinput10, keyinput11, keyinput12, keyinput13, keyinput14, keyinput15, keyinput16, keyinput17, keyinput18, keyinput19, keyinput20, keyinput21, keyinput22, keyinput23, keyinput24, keyinput25, keyinput26, keyinput27, keyinput28, keyinput29, keyinput30, keyinput31, keyinput32, keyinput33, keyinput34, keyinput35, keyinput36, keyinput37, keyinput38, keyinput39, keyinput40, keyinput41, keyinput42, keyinput43, keyinput44, keyinput45, keyinput46, keyinput47, keyinput48, keyinput49, keyinput50, keyinput51, keyinput52, keyinput53, keyinput54, keyinput55, keyinput56, keyinput57, keyinput58, keyinput59, keyinput60, keyinput61, keyinput62, keyinput63, ADDR_REG_19__SCAN_IN, ADDR_REG_18__SCAN_IN, ADDR_REG_17__SCAN_IN, ADDR_REG_16__SCAN_IN, ADDR_REG_15__SCAN_IN, ADDR_REG_14__SCAN_IN, ADDR_REG_13__SCAN_IN, ADDR_REG_12__SCAN_IN, ADDR_REG_11__SCAN_IN, ADDR_REG_10__SCAN_IN, ADDR_REG_9__SCAN_IN, ADDR_REG_8__SCAN_IN, ADDR_REG_7__SCAN_IN, ADDR_REG_6__SCAN_IN, ADDR_REG_5__SCAN_IN, ADDR_REG_4__SCAN_IN, ADDR_REG_3__SCAN_IN, ADDR_REG_2__SCAN_IN, ADDR_REG_1__SCAN_IN, ADDR_REG_0__SCAN_IN, DATAO_REG_31__SCAN_IN, DATAO_REG_30__SCAN_IN, DATAO_REG_29__SCAN_IN, DATAO_REG_28__SCAN_IN, DATAO_REG_27__SCAN_IN, DATAO_REG_26__SCAN_IN, DATAO_REG_25__SCAN_IN, DATAO_REG_24__SCAN_IN, DATAO_REG_23__SCAN_IN, DATAO_REG_22__SCAN_IN, DATAO_REG_21__SCAN_IN, DATAO_REG_20__SCAN_IN, DATAO_REG_19__SCAN_IN, DATAO_REG_18__SCAN_IN, DATAO_REG_17__SCAN_IN, DATAO_REG_16__SCAN_IN, DATAO_REG_15__SCAN_IN, DATAO_REG_14__SCAN_IN, DATAO_REG_13__SCAN_IN, DATAO_REG_12__SCAN_IN, DATAO_REG_11__SCAN_IN, DATAO_REG_10__SCAN_IN, DATAO_REG_9__SCAN_IN, DATAO_REG_8__SCAN_IN, DATAO_REG_7__SCAN_IN, DATAO_REG_6__SCAN_IN, DATAO_REG_5__SCAN_IN, DATAO_REG_4__SCAN_IN, DATAO_REG_3__SCAN_IN, DATAO_REG_2__SCAN_IN, DATAO_REG_1__SCAN_IN, DATAO_REG_0__SCAN_IN, RD_REG_SCAN_IN, WR_REG_SCAN_IN, U3352, U3351, U3350, U3349, U3348, U3347, U3346, U3345, U3344, U3343, U3342, U3341, U3340, U3339, U3338, U3337, U3336, U3335, U3334, U3333, U3332, U3331, U3330, U3329, U3328, U3327, U3326, U3325, U3324, U3323, U3322, U3321, U3458, U3459, U3320, U3319, U3318, U3317, U3316, U3315, U3314, U3313, U3312, U3311, U3310, U3309, U3308, U3307, U3306, U3305, U3304, U3303, U3302, U3301, U3300, U3299, U3298, U3297, U3296, U3295, U3294, U3293, U3292, U3291, U3467, U3469, U3471, U3473, U3475, U3477, U3479, U3481, U3483, U3485, U3487, U3489, U3491, U3493, U3495, U3497, U3499, U3501, U3503, U3505, U3506, U3507, U3508, U3509, U3510, U3511, U3512, U3513, U3514, U3515, U3516, U3517, U3518, U3519, U3520, U3521, U3522, U3523, U3524, U3525, U3526, U3527, U3528, U3529, U3530, U3531, U3532, U3533, U3534, U3535, U3536, U3537, U3538, U3539, U3540, U3541, U3542, U3543, U3544, U3545, U3546, U3547, U3548, U3549, U3290, U3289, U3288, U3287, U3286, U3285, U3284, U3283, U3282, U3281, U3280, U3279, U3278, U3277, U3276, U3275, U3274, U3273, U3272, U3271, U3270, U3269, U3268, U3267, U3266, U3265, U3264, U3263, U3262, U3354, U3261, U3260, U3259, U3258, U3257, U3256, U3255, U3254, U3253, U3252, U3251, U3250, U3249, U3248, U3247, U3246, U3245, U3244, U3243, U3242, U3241, U3240, U3550, U3551, U3552, U3553, U3554, U3555, U3556, U3557, U3558, U3559, U3560, U3561, U3562, U3563, U3564, U3565, U3566, U3567, U3568, U3569, U3570, U3571, U3572, U3573, U3574, U3575, U3576, U3577, U3578, U3579, U3580, U3581, U3239, U3238, U3237, U3236, U3235, U3234, U3233, U3232, U3231, U3230, U3229, U3228, U3227, U3226, U3225, U3224, U3223, U3222, U3221, U3220, U3219, U3218, U3217, U3216, U3215, U3214, U3213, U3212, U3211, U3210, U3149, U3148, U4043);

  input WR_REG_SCAN_IN, DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, DATAI_27_, DATAI_26_, DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, DATAI_21_, DATAI_20_, DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, DATAI_15_, DATAI_14_, DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, DATAI_9_, DATAI_8_, DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, DATAI_2_, DATAI_1_, DATAI_0_, RD_REG_SCAN_IN, STATE_REG_SCAN_IN, REG3_REG_7__SCAN_IN, REG3_REG_27__SCAN_IN, REG3_REG_14__SCAN_IN, REG3_REG_23__SCAN_IN, REG3_REG_10__SCAN_IN, REG3_REG_3__SCAN_IN, REG3_REG_19__SCAN_IN, REG3_REG_28__SCAN_IN, REG3_REG_8__SCAN_IN, REG3_REG_1__SCAN_IN, REG3_REG_21__SCAN_IN, REG3_REG_12__SCAN_IN, REG3_REG_25__SCAN_IN, REG3_REG_16__SCAN_IN, REG3_REG_5__SCAN_IN, REG3_REG_17__SCAN_IN, REG3_REG_24__SCAN_IN, REG3_REG_4__SCAN_IN, REG3_REG_9__SCAN_IN, REG3_REG_0__SCAN_IN, REG3_REG_20__SCAN_IN, REG3_REG_13__SCAN_IN, IR_REG_0__SCAN_IN, IR_REG_1__SCAN_IN, IR_REG_2__SCAN_IN, IR_REG_3__SCAN_IN, IR_REG_4__SCAN_IN, IR_REG_5__SCAN_IN, IR_REG_6__SCAN_IN, IR_REG_7__SCAN_IN, IR_REG_8__SCAN_IN, IR_REG_9__SCAN_IN, IR_REG_10__SCAN_IN, IR_REG_11__SCAN_IN, IR_REG_12__SCAN_IN, IR_REG_13__SCAN_IN, IR_REG_14__SCAN_IN, IR_REG_15__SCAN_IN, IR_REG_16__SCAN_IN, IR_REG_17__SCAN_IN, IR_REG_18__SCAN_IN, IR_REG_19__SCAN_IN, IR_REG_20__SCAN_IN, IR_REG_21__SCAN_IN, IR_REG_22__SCAN_IN, IR_REG_23__SCAN_IN, IR_REG_24__SCAN_IN, IR_REG_25__SCAN_IN, IR_REG_26__SCAN_IN, IR_REG_27__SCAN_IN, IR_REG_28__SCAN_IN, IR_REG_29__SCAN_IN, IR_REG_30__SCAN_IN, IR_REG_31__SCAN_IN, D_REG_0__SCAN_IN, D_REG_1__SCAN_IN, D_REG_2__SCAN_IN, D_REG_3__SCAN_IN, D_REG_4__SCAN_IN, D_REG_5__SCAN_IN, D_REG_6__SCAN_IN, D_REG_7__SCAN_IN, D_REG_8__SCAN_IN, D_REG_9__SCAN_IN, D_REG_10__SCAN_IN, D_REG_11__SCAN_IN, D_REG_12__SCAN_IN, D_REG_13__SCAN_IN, D_REG_14__SCAN_IN, D_REG_15__SCAN_IN, D_REG_16__SCAN_IN, D_REG_17__SCAN_IN, D_REG_18__SCAN_IN, D_REG_19__SCAN_IN, D_REG_20__SCAN_IN, D_REG_21__SCAN_IN, D_REG_22__SCAN_IN, D_REG_23__SCAN_IN, D_REG_24__SCAN_IN, D_REG_25__SCAN_IN, D_REG_26__SCAN_IN, D_REG_27__SCAN_IN, D_REG_28__SCAN_IN, D_REG_29__SCAN_IN, D_REG_30__SCAN_IN, D_REG_31__SCAN_IN, REG0_REG_0__SCAN_IN, REG0_REG_1__SCAN_IN, REG0_REG_2__SCAN_IN, REG0_REG_3__SCAN_IN, REG0_REG_4__SCAN_IN, REG0_REG_5__SCAN_IN, REG0_REG_6__SCAN_IN, REG0_REG_7__SCAN_IN, REG0_REG_8__SCAN_IN, REG0_REG_9__SCAN_IN, REG0_REG_10__SCAN_IN, REG0_REG_11__SCAN_IN, REG0_REG_12__SCAN_IN, REG0_REG_13__SCAN_IN, REG0_REG_14__SCAN_IN, REG0_REG_15__SCAN_IN, REG0_REG_16__SCAN_IN, REG0_REG_17__SCAN_IN, REG0_REG_18__SCAN_IN, REG0_REG_19__SCAN_IN, REG0_REG_20__SCAN_IN, REG0_REG_21__SCAN_IN, REG0_REG_22__SCAN_IN, REG0_REG_23__SCAN_IN, REG0_REG_24__SCAN_IN, REG0_REG_25__SCAN_IN, REG0_REG_26__SCAN_IN, REG0_REG_27__SCAN_IN, REG0_REG_28__SCAN_IN, REG0_REG_29__SCAN_IN, REG0_REG_30__SCAN_IN, REG0_REG_31__SCAN_IN, REG1_REG_0__SCAN_IN, REG1_REG_1__SCAN_IN, REG1_REG_2__SCAN_IN, REG1_REG_3__SCAN_IN, REG1_REG_4__SCAN_IN, REG1_REG_5__SCAN_IN, REG1_REG_6__SCAN_IN, REG1_REG_7__SCAN_IN, REG1_REG_8__SCAN_IN, REG1_REG_9__SCAN_IN, REG1_REG_10__SCAN_IN, REG1_REG_11__SCAN_IN, REG1_REG_12__SCAN_IN, REG1_REG_13__SCAN_IN, REG1_REG_14__SCAN_IN, REG1_REG_15__SCAN_IN, REG1_REG_16__SCAN_IN, REG1_REG_17__SCAN_IN, REG1_REG_18__SCAN_IN, REG1_REG_19__SCAN_IN, REG1_REG_20__SCAN_IN, REG1_REG_21__SCAN_IN, REG1_REG_22__SCAN_IN, REG1_REG_23__SCAN_IN, REG1_REG_24__SCAN_IN, REG1_REG_25__SCAN_IN, REG1_REG_26__SCAN_IN, REG1_REG_27__SCAN_IN, REG1_REG_28__SCAN_IN, REG1_REG_29__SCAN_IN, REG1_REG_30__SCAN_IN, REG1_REG_31__SCAN_IN, REG2_REG_0__SCAN_IN, REG2_REG_1__SCAN_IN, REG2_REG_2__SCAN_IN, REG2_REG_3__SCAN_IN, REG2_REG_4__SCAN_IN, REG2_REG_5__SCAN_IN, REG2_REG_6__SCAN_IN, REG2_REG_7__SCAN_IN, REG2_REG_8__SCAN_IN, REG2_REG_9__SCAN_IN, REG2_REG_10__SCAN_IN, REG2_REG_11__SCAN_IN, REG2_REG_12__SCAN_IN, REG2_REG_13__SCAN_IN, REG2_REG_14__SCAN_IN, REG2_REG_15__SCAN_IN, REG2_REG_16__SCAN_IN, REG2_REG_17__SCAN_IN, REG2_REG_18__SCAN_IN, REG2_REG_19__SCAN_IN, REG2_REG_20__SCAN_IN, REG2_REG_21__SCAN_IN, REG2_REG_22__SCAN_IN, REG2_REG_23__SCAN_IN, REG2_REG_24__SCAN_IN, REG2_REG_25__SCAN_IN, REG2_REG_26__SCAN_IN, REG2_REG_27__SCAN_IN, REG2_REG_28__SCAN_IN, REG2_REG_29__SCAN_IN, REG2_REG_30__SCAN_IN, REG2_REG_31__SCAN_IN, ADDR_REG_19__SCAN_IN, ADDR_REG_18__SCAN_IN, ADDR_REG_17__SCAN_IN, ADDR_REG_16__SCAN_IN, ADDR_REG_15__SCAN_IN, ADDR_REG_14__SCAN_IN, ADDR_REG_13__SCAN_IN, ADDR_REG_12__SCAN_IN, ADDR_REG_11__SCAN_IN, ADDR_REG_10__SCAN_IN, ADDR_REG_9__SCAN_IN, ADDR_REG_8__SCAN_IN, ADDR_REG_7__SCAN_IN, ADDR_REG_6__SCAN_IN, ADDR_REG_5__SCAN_IN, ADDR_REG_4__SCAN_IN, ADDR_REG_3__SCAN_IN, ADDR_REG_2__SCAN_IN, ADDR_REG_1__SCAN_IN, ADDR_REG_0__SCAN_IN, DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN, DATAO_REG_2__SCAN_IN, DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN, DATAO_REG_5__SCAN_IN, DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN, DATAO_REG_8__SCAN_IN, DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN, DATAO_REG_11__SCAN_IN, DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN, DATAO_REG_14__SCAN_IN, DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN, DATAO_REG_17__SCAN_IN, DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN, DATAO_REG_20__SCAN_IN, DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN, DATAO_REG_23__SCAN_IN, DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN, DATAO_REG_26__SCAN_IN, DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN, DATAO_REG_29__SCAN_IN, DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN, B_REG_SCAN_IN, REG3_REG_15__SCAN_IN, REG3_REG_26__SCAN_IN, REG3_REG_6__SCAN_IN, REG3_REG_18__SCAN_IN, REG3_REG_2__SCAN_IN, REG3_REG_11__SCAN_IN, REG3_REG_22__SCAN_IN, keyinput0, keyinput1, keyinput2, keyinput3, keyinput4, keyinput5, keyinput6, keyinput7, keyinput8, keyinput9, keyinput10, keyinput11, keyinput12, keyinput13, keyinput14, keyinput15, keyinput16, keyinput17, keyinput18, keyinput19, keyinput20, keyinput21, keyinput22, keyinput23, keyinput24, keyinput25, keyinput26, keyinput27, keyinput28, keyinput29, keyinput30, keyinput31, keyinput32, keyinput33, keyinput34, keyinput35, keyinput36, keyinput37, keyinput38, keyinput39, keyinput40, keyinput41, keyinput42, keyinput43, keyinput44, keyinput45, keyinput46, keyinput47, keyinput48, keyinput49, keyinput50, keyinput51, keyinput52, keyinput53, keyinput54, keyinput55, keyinput56, keyinput57, keyinput58, keyinput59, keyinput60, keyinput61, keyinput62, keyinput63;
  output ADDR_REG_19__SCAN_IN, ADDR_REG_18__SCAN_IN, ADDR_REG_17__SCAN_IN, ADDR_REG_16__SCAN_IN, ADDR_REG_15__SCAN_IN, ADDR_REG_14__SCAN_IN, ADDR_REG_13__SCAN_IN, ADDR_REG_12__SCAN_IN, ADDR_REG_11__SCAN_IN, ADDR_REG_10__SCAN_IN, ADDR_REG_9__SCAN_IN, ADDR_REG_8__SCAN_IN, ADDR_REG_7__SCAN_IN, ADDR_REG_6__SCAN_IN, ADDR_REG_5__SCAN_IN, ADDR_REG_4__SCAN_IN, ADDR_REG_3__SCAN_IN, ADDR_REG_2__SCAN_IN, ADDR_REG_1__SCAN_IN, ADDR_REG_0__SCAN_IN, DATAO_REG_31__SCAN_IN, DATAO_REG_30__SCAN_IN, DATAO_REG_29__SCAN_IN, DATAO_REG_28__SCAN_IN, DATAO_REG_27__SCAN_IN, DATAO_REG_26__SCAN_IN, DATAO_REG_25__SCAN_IN, DATAO_REG_24__SCAN_IN, DATAO_REG_23__SCAN_IN, DATAO_REG_22__SCAN_IN, DATAO_REG_21__SCAN_IN, DATAO_REG_20__SCAN_IN, DATAO_REG_19__SCAN_IN, DATAO_REG_18__SCAN_IN, DATAO_REG_17__SCAN_IN, DATAO_REG_16__SCAN_IN, DATAO_REG_15__SCAN_IN, DATAO_REG_14__SCAN_IN, DATAO_REG_13__SCAN_IN, DATAO_REG_12__SCAN_IN, DATAO_REG_11__SCAN_IN, DATAO_REG_10__SCAN_IN, DATAO_REG_9__SCAN_IN, DATAO_REG_8__SCAN_IN, DATAO_REG_7__SCAN_IN, DATAO_REG_6__SCAN_IN, DATAO_REG_5__SCAN_IN, DATAO_REG_4__SCAN_IN, DATAO_REG_3__SCAN_IN, DATAO_REG_2__SCAN_IN, DATAO_REG_1__SCAN_IN, DATAO_REG_0__SCAN_IN, RD_REG_SCAN_IN, WR_REG_SCAN_IN, U3352, U3351, U3350, U3349, U3348, U3347, U3346, U3345, U3344, U3343, U3342, U3341, U3340, U3339, U3338, U3337, U3336, U3335, U3334, U3333, U3332, U3331, U3330, U3329, U3328, U3327, U3326, U3325, U3324, U3323, U3322, U3321, U3458, U3459, U3320, U3319, U3318, U3317, U3316, U3315, U3314, U3313, U3312, U3311, U3310, U3309, U3308, U3307, U3306, U3305, U3304, U3303, U3302, U3301, U3300, U3299, U3298, U3297, U3296, U3295, U3294, U3293, U3292, U3291, U3467, U3469, U3471, U3473, U3475, U3477, U3479, U3481, U3483, U3485, U3487, U3489, U3491, U3493, U3495, U3497, U3499, U3501, U3503, U3505, U3506, U3507, U3508, U3509, U3510, U3511, U3512, U3513, U3514, U3515, U3516, U3517, U3518, U3519, U3520, U3521, U3522, U3523, U3524, U3525, U3526, U3527, U3528, U3529, U3530, U3531, U3532, U3533, U3534, U3535, U3536, U3537, U3538, U3539, U3540, U3541, U3542, U3543, U3544, U3545, U3546, U3547, U3548, U3549, U3290, U3289, U3288, U3287, U3286, U3285, U3284, U3283, U3282, U3281, U3280, U3279, U3278, U3277, U3276, U3275, U3274, U3273, U3272, U3271, U3270, U3269, U3268, U3267, U3266, U3265, U3264, U3263, U3262, U3354, U3261, U3260, U3259, U3258, U3257, U3256, U3255, U3254, U3253, U3252, U3251, U3250, U3249, U3248, U3247, U3246, U3245, U3244, U3243, U3242, U3241, U3240, U3550, U3551, U3552, U3553, U3554, U3555, U3556, U3557, U3558, U3559, U3560, U3561, U3562, U3563, U3564, U3565, U3566, U3567, U3568, U3569, U3570, U3571, U3572, U3573, U3574, U3575, U3576, U3577, U3578, U3579, U3580, U3581, U3239, U3238, U3237, U3236, U3235, U3234, U3233, U3232, U3231, U3230, U3229, U3228, U3227, U3226, U3225, U3224, U3223, U3222, U3221, U3220, U3219, U3218, U3217, U3216, U3215, U3214, U3213, U3212, U3211, U3210, U3149, U3148, U4043;
  wire ADD_95_U10, ADD_95_U100, ADD_95_U101, ADD_95_U102, ADD_95_U103, ADD_95_U104, ADD_95_U105, ADD_95_U106, ADD_95_U107, ADD_95_U108, ADD_95_U109, ADD_95_U11, ADD_95_U110, ADD_95_U111, ADD_95_U112, ADD_95_U113, ADD_95_U114, ADD_95_U115, ADD_95_U116, ADD_95_U117, ADD_95_U118, ADD_95_U119, ADD_95_U12, ADD_95_U120, ADD_95_U121, ADD_95_U122, ADD_95_U123, ADD_95_U124, ADD_95_U125, ADD_95_U126, ADD_95_U127, ADD_95_U128, ADD_95_U129, ADD_95_U13, ADD_95_U130, ADD_95_U131, ADD_95_U132, ADD_95_U133, ADD_95_U134, ADD_95_U135, ADD_95_U136, ADD_95_U137, ADD_95_U138, ADD_95_U139, ADD_95_U14, ADD_95_U140, ADD_95_U141, ADD_95_U142, ADD_95_U143, ADD_95_U144, ADD_95_U145, ADD_95_U146, ADD_95_U147, ADD_95_U148, ADD_95_U149, ADD_95_U15, ADD_95_U150, ADD_95_U151, ADD_95_U152, ADD_95_U153, ADD_95_U154, ADD_95_U155, ADD_95_U156, ADD_95_U157, ADD_95_U158, ADD_95_U159, ADD_95_U16, ADD_95_U17, ADD_95_U18, ADD_95_U19, ADD_95_U20, ADD_95_U21, ADD_95_U22, ADD_95_U23, ADD_95_U24, ADD_95_U25, ADD_95_U26, ADD_95_U27, ADD_95_U28, ADD_95_U29, ADD_95_U30, ADD_95_U31, ADD_95_U32, ADD_95_U33, ADD_95_U34, ADD_95_U35, ADD_95_U36, ADD_95_U37, ADD_95_U38, ADD_95_U39, ADD_95_U4, ADD_95_U40, ADD_95_U41, ADD_95_U42, ADD_95_U43, ADD_95_U44, ADD_95_U45, ADD_95_U46, ADD_95_U47, ADD_95_U48, ADD_95_U49, ADD_95_U5, ADD_95_U50, ADD_95_U51, ADD_95_U52, ADD_95_U53, ADD_95_U54, ADD_95_U55, ADD_95_U56, ADD_95_U57, ADD_95_U58, ADD_95_U59, ADD_95_U6, ADD_95_U60, ADD_95_U61, ADD_95_U62, ADD_95_U63, ADD_95_U64, ADD_95_U65, ADD_95_U66, ADD_95_U67, ADD_95_U68, ADD_95_U69, ADD_95_U7, ADD_95_U70, ADD_95_U71, ADD_95_U72, ADD_95_U73, ADD_95_U74, ADD_95_U75, ADD_95_U76, ADD_95_U77, ADD_95_U78, ADD_95_U79, ADD_95_U8, ADD_95_U80, ADD_95_U81, ADD_95_U82, ADD_95_U83, ADD_95_U84, ADD_95_U85, ADD_95_U86, ADD_95_U87, ADD_95_U88, ADD_95_U89, ADD_95_U9, ADD_95_U90, ADD_95_U91, ADD_95_U92, ADD_95_U93, ADD_95_U94, ADD_95_U95, ADD_95_U96, ADD_95_U97, ADD_95_U98, ADD_95_U99, R1105_U10, R1105_U100, R1105_U101, R1105_U102, R1105_U103, R1105_U104, R1105_U105, R1105_U106, R1105_U107, R1105_U108, R1105_U109, R1105_U11, R1105_U110, R1105_U111, R1105_U112, R1105_U113, R1105_U114, R1105_U115, R1105_U116, R1105_U117, R1105_U118, R1105_U119, R1105_U12, R1105_U120, R1105_U121, R1105_U122, R1105_U123, R1105_U124, R1105_U125, R1105_U126, R1105_U127, R1105_U128, R1105_U129, R1105_U13, R1105_U130, R1105_U131, R1105_U132, R1105_U133, R1105_U134, R1105_U135, R1105_U136, R1105_U137, R1105_U138, R1105_U139, R1105_U14, R1105_U140, R1105_U141, R1105_U142, R1105_U143, R1105_U144, R1105_U145, R1105_U146, R1105_U147, R1105_U148, R1105_U149, R1105_U15, R1105_U150, R1105_U151, R1105_U152, R1105_U153, R1105_U154, R1105_U155, R1105_U156, R1105_U157, R1105_U158, R1105_U159, R1105_U16, R1105_U160, R1105_U161, R1105_U162, R1105_U163, R1105_U164, R1105_U165, R1105_U166, R1105_U167, R1105_U168, R1105_U169, R1105_U17, R1105_U170, R1105_U171, R1105_U172, R1105_U173, R1105_U174, R1105_U175, R1105_U176, R1105_U177, R1105_U178, R1105_U179, R1105_U18, R1105_U180, R1105_U181, R1105_U182, R1105_U183, R1105_U184, R1105_U185, R1105_U186, R1105_U187, R1105_U188, R1105_U189, R1105_U19, R1105_U190, R1105_U191, R1105_U192, R1105_U193, R1105_U194, R1105_U195, R1105_U196, R1105_U197, R1105_U198, R1105_U199, R1105_U20, R1105_U200, R1105_U201, R1105_U202, R1105_U203, R1105_U204, R1105_U205, R1105_U206, R1105_U207, R1105_U208, R1105_U209, R1105_U21, R1105_U210, R1105_U211, R1105_U212, R1105_U213, R1105_U214, R1105_U215, R1105_U216, R1105_U217, R1105_U218, R1105_U219, R1105_U22, R1105_U220, R1105_U221, R1105_U222, R1105_U223, R1105_U224, R1105_U225, R1105_U226, R1105_U227, R1105_U228, R1105_U229, R1105_U23, R1105_U230, R1105_U231, R1105_U232, R1105_U233, R1105_U234, R1105_U235, R1105_U236, R1105_U237, R1105_U238, R1105_U239, R1105_U24, R1105_U240, R1105_U241, R1105_U242, R1105_U243, R1105_U244, R1105_U245, R1105_U246, R1105_U247, R1105_U248, R1105_U249, R1105_U25, R1105_U250, R1105_U251, R1105_U252, R1105_U253, R1105_U254, R1105_U255, R1105_U256, R1105_U257, R1105_U258, R1105_U259, R1105_U26, R1105_U260, R1105_U261, R1105_U262, R1105_U263, R1105_U264, R1105_U265, R1105_U266, R1105_U267, R1105_U268, R1105_U269, R1105_U27, R1105_U270, R1105_U271, R1105_U272, R1105_U273, R1105_U274, R1105_U275, R1105_U276, R1105_U277, R1105_U278, R1105_U279, R1105_U28, R1105_U280, R1105_U281, R1105_U282, R1105_U283, R1105_U284, R1105_U285, R1105_U286, R1105_U287, R1105_U288, R1105_U289, R1105_U29, R1105_U290, R1105_U291, R1105_U292, R1105_U293, R1105_U294, R1105_U295, R1105_U296, R1105_U297, R1105_U298, R1105_U299, R1105_U30, R1105_U300, R1105_U301, R1105_U302, R1105_U303, R1105_U304, R1105_U305, R1105_U306, R1105_U307, R1105_U308, R1105_U309, R1105_U31, R1105_U310, R1105_U311, R1105_U32, R1105_U33, R1105_U34, R1105_U35, R1105_U36, R1105_U37, R1105_U38, R1105_U39, R1105_U4, R1105_U40, R1105_U41, R1105_U42, R1105_U43, R1105_U44, R1105_U45, R1105_U46, R1105_U47, R1105_U48, R1105_U49, R1105_U5, R1105_U50, R1105_U51, R1105_U52, R1105_U53, R1105_U54, R1105_U55, R1105_U56, R1105_U57, R1105_U58, R1105_U59, R1105_U6, R1105_U60, R1105_U61, R1105_U62, R1105_U63, R1105_U64, R1105_U65, R1105_U66, R1105_U67, R1105_U68, R1105_U69, R1105_U7, R1105_U70, R1105_U71, R1105_U72, R1105_U73, R1105_U74, R1105_U75, R1105_U76, R1105_U77, R1105_U78, R1105_U79, R1105_U8, R1105_U80, R1105_U81, R1105_U82, R1105_U83, R1105_U84, R1105_U85, R1105_U86, R1105_U87, R1105_U88, R1105_U89, R1105_U9, R1105_U90, R1105_U91, R1105_U92, R1105_U93, R1105_U94, R1105_U95, R1105_U96, R1105_U97, R1105_U98, R1105_U99, R1117_U10, R1117_U100, R1117_U101, R1117_U102, R1117_U103, R1117_U104, R1117_U105, R1117_U106, R1117_U107, R1117_U108, R1117_U109, R1117_U11, R1117_U110, R1117_U111, R1117_U112, R1117_U113, R1117_U114, R1117_U115, R1117_U116, R1117_U117, R1117_U118, R1117_U119, R1117_U12, R1117_U120, R1117_U121, R1117_U122, R1117_U123, R1117_U124, R1117_U125, R1117_U126, R1117_U127, R1117_U128, R1117_U129, R1117_U13, R1117_U130, R1117_U131, R1117_U132, R1117_U133, R1117_U134, R1117_U135, R1117_U136, R1117_U137, R1117_U138, R1117_U139, R1117_U14, R1117_U140, R1117_U141, R1117_U142, R1117_U143, R1117_U144, R1117_U145, R1117_U146, R1117_U147, R1117_U148, R1117_U149, R1117_U15, R1117_U150, R1117_U151, R1117_U152, R1117_U153, R1117_U154, R1117_U155, R1117_U156, R1117_U157, R1117_U158, R1117_U159, R1117_U16, R1117_U160, R1117_U161, R1117_U162, R1117_U163, R1117_U164, R1117_U165, R1117_U166, R1117_U167, R1117_U168, R1117_U169, R1117_U17, R1117_U170, R1117_U171, R1117_U172, R1117_U173, R1117_U174, R1117_U175, R1117_U176, R1117_U177, R1117_U178, R1117_U179, R1117_U18, R1117_U180, R1117_U181, R1117_U182, R1117_U183, R1117_U184, R1117_U185, R1117_U186, R1117_U187, R1117_U188, R1117_U189, R1117_U19, R1117_U190, R1117_U191, R1117_U192, R1117_U193, R1117_U194, R1117_U195, R1117_U196, R1117_U197, R1117_U198, R1117_U199, R1117_U20, R1117_U200, R1117_U201, R1117_U202, R1117_U203, R1117_U204, R1117_U205, R1117_U206, R1117_U207, R1117_U208, R1117_U209, R1117_U21, R1117_U210, R1117_U211, R1117_U212, R1117_U213, R1117_U214, R1117_U215, R1117_U216, R1117_U217, R1117_U218, R1117_U219, R1117_U22, R1117_U220, R1117_U221, R1117_U222, R1117_U223, R1117_U224, R1117_U225, R1117_U226, R1117_U227, R1117_U228, R1117_U229, R1117_U23, R1117_U230, R1117_U231, R1117_U232, R1117_U233, R1117_U234, R1117_U235, R1117_U236, R1117_U237, R1117_U238, R1117_U239, R1117_U24, R1117_U240, R1117_U241, R1117_U242, R1117_U243, R1117_U244, R1117_U245, R1117_U246, R1117_U247, R1117_U248, R1117_U249, R1117_U25, R1117_U250, R1117_U251, R1117_U252, R1117_U253, R1117_U254, R1117_U255, R1117_U256, R1117_U257, R1117_U258, R1117_U259, R1117_U26, R1117_U260, R1117_U261, R1117_U262, R1117_U263, R1117_U264, R1117_U265, R1117_U266, R1117_U267, R1117_U268, R1117_U269, R1117_U27, R1117_U270, R1117_U271, R1117_U272, R1117_U273, R1117_U274, R1117_U275, R1117_U276, R1117_U277, R1117_U278, R1117_U279, R1117_U28, R1117_U280, R1117_U281, R1117_U282, R1117_U283, R1117_U284, R1117_U285, R1117_U286, R1117_U287, R1117_U288, R1117_U289, R1117_U29, R1117_U290, R1117_U291, R1117_U292, R1117_U293, R1117_U294, R1117_U295, R1117_U296, R1117_U297, R1117_U298, R1117_U299, R1117_U30, R1117_U300, R1117_U301, R1117_U302, R1117_U303, R1117_U304, R1117_U305, R1117_U306, R1117_U307, R1117_U308, R1117_U309, R1117_U31, R1117_U310, R1117_U311, R1117_U312, R1117_U313, R1117_U314, R1117_U315, R1117_U316, R1117_U317, R1117_U318, R1117_U319, R1117_U32, R1117_U320, R1117_U321, R1117_U322, R1117_U323, R1117_U324, R1117_U325, R1117_U326, R1117_U327, R1117_U328, R1117_U329, R1117_U33, R1117_U330, R1117_U331, R1117_U332, R1117_U333, R1117_U334, R1117_U335, R1117_U336, R1117_U337, R1117_U338, R1117_U339, R1117_U34, R1117_U340, R1117_U341, R1117_U342, R1117_U343, R1117_U344, R1117_U345, R1117_U346, R1117_U347, R1117_U348, R1117_U349, R1117_U35, R1117_U350, R1117_U351, R1117_U352, R1117_U353, R1117_U354, R1117_U355, R1117_U356, R1117_U357, R1117_U358, R1117_U359, R1117_U36, R1117_U360, R1117_U361, R1117_U362, R1117_U363, R1117_U364, R1117_U365, R1117_U366, R1117_U367, R1117_U368, R1117_U369, R1117_U37, R1117_U370, R1117_U371, R1117_U372, R1117_U373, R1117_U374, R1117_U375, R1117_U376, R1117_U377, R1117_U378, R1117_U379, R1117_U38, R1117_U380, R1117_U381, R1117_U382, R1117_U383, R1117_U384, R1117_U385, R1117_U386, R1117_U387, R1117_U388, R1117_U389, R1117_U39, R1117_U390, R1117_U391, R1117_U392, R1117_U393, R1117_U394, R1117_U395, R1117_U396, R1117_U397, R1117_U398, R1117_U399, R1117_U40, R1117_U400, R1117_U401, R1117_U402, R1117_U403, R1117_U404, R1117_U405, R1117_U406, R1117_U407, R1117_U408, R1117_U409, R1117_U41, R1117_U410, R1117_U411, R1117_U412, R1117_U413, R1117_U414, R1117_U415, R1117_U416, R1117_U417, R1117_U418, R1117_U419, R1117_U42, R1117_U420, R1117_U421, R1117_U422, R1117_U423, R1117_U424, R1117_U425, R1117_U426, R1117_U427, R1117_U428, R1117_U429, R1117_U43, R1117_U430, R1117_U431, R1117_U432, R1117_U433, R1117_U434, R1117_U435, R1117_U436, R1117_U437, R1117_U438, R1117_U439, R1117_U44, R1117_U440, R1117_U441, R1117_U442, R1117_U443, R1117_U444, R1117_U445, R1117_U446, R1117_U447, R1117_U448, R1117_U449, R1117_U45, R1117_U450, R1117_U451, R1117_U452, R1117_U453, R1117_U454, R1117_U455, R1117_U456, R1117_U457, R1117_U458, R1117_U459, R1117_U46, R1117_U460, R1117_U461, R1117_U462, R1117_U463, R1117_U464, R1117_U465, R1117_U466, R1117_U467, R1117_U468, R1117_U469, R1117_U47, R1117_U470, R1117_U471, R1117_U472, R1117_U473, R1117_U474, R1117_U475, R1117_U476, R1117_U477, R1117_U478, R1117_U479, R1117_U48, R1117_U480, R1117_U481, R1117_U482, R1117_U483, R1117_U484, R1117_U485, R1117_U486, R1117_U487, R1117_U488, R1117_U489, R1117_U49, R1117_U490, R1117_U491, R1117_U492, R1117_U493, R1117_U494, R1117_U495, R1117_U496, R1117_U497, R1117_U498, R1117_U499, R1117_U50, R1117_U500, R1117_U501, R1117_U502, R1117_U503, R1117_U504, R1117_U505, R1117_U506, R1117_U507, R1117_U508, R1117_U509, R1117_U51, R1117_U510, R1117_U511, R1117_U512, R1117_U513, R1117_U514, R1117_U515, R1117_U52, R1117_U53, R1117_U54, R1117_U55, R1117_U56, R1117_U57, R1117_U58, R1117_U59, R1117_U6, R1117_U60, R1117_U61, R1117_U62, R1117_U63, R1117_U64, R1117_U65, R1117_U66, R1117_U67, R1117_U68, R1117_U69, R1117_U7, R1117_U70, R1117_U71, R1117_U72, R1117_U73, R1117_U74, R1117_U75, R1117_U76, R1117_U77, R1117_U78, R1117_U79, R1117_U8, R1117_U80, R1117_U81, R1117_U82, R1117_U83, R1117_U84, R1117_U85, R1117_U86, R1117_U87, R1117_U88, R1117_U89, R1117_U9, R1117_U90, R1117_U91, R1117_U92, R1117_U93, R1117_U94, R1117_U95, R1117_U96, R1117_U97, R1117_U98, R1117_U99, R1138_U10, R1138_U100, R1138_U101, R1138_U102, R1138_U103, R1138_U104, R1138_U105, R1138_U106, R1138_U107, R1138_U108, R1138_U109, R1138_U11, R1138_U110, R1138_U111, R1138_U112, R1138_U113, R1138_U114, R1138_U115, R1138_U116, R1138_U117, R1138_U118, R1138_U119, R1138_U12, R1138_U120, R1138_U121, R1138_U122, R1138_U123, R1138_U124, R1138_U125, R1138_U126, R1138_U127, R1138_U128, R1138_U129, R1138_U13, R1138_U130, R1138_U131, R1138_U132, R1138_U133, R1138_U134, R1138_U135, R1138_U136, R1138_U137, R1138_U138, R1138_U139, R1138_U14, R1138_U140, R1138_U141, R1138_U142, R1138_U143, R1138_U144, R1138_U145, R1138_U146, R1138_U147, R1138_U148, R1138_U149, R1138_U15, R1138_U150, R1138_U151, R1138_U152, R1138_U153, R1138_U154, R1138_U155, R1138_U156, R1138_U157, R1138_U158, R1138_U159, R1138_U16, R1138_U160, R1138_U161, R1138_U162, R1138_U163, R1138_U164, R1138_U165, R1138_U166, R1138_U167, R1138_U168, R1138_U169, R1138_U17, R1138_U170, R1138_U171, R1138_U172, R1138_U173, R1138_U174, R1138_U175, R1138_U176, R1138_U177, R1138_U178, R1138_U179, R1138_U18, R1138_U180, R1138_U181, R1138_U182, R1138_U183, R1138_U184, R1138_U185, R1138_U186, R1138_U187, R1138_U188, R1138_U189, R1138_U19, R1138_U190, R1138_U191, R1138_U192, R1138_U193, R1138_U194, R1138_U195, R1138_U196, R1138_U197, R1138_U198, R1138_U199, R1138_U20, R1138_U200, R1138_U201, R1138_U202, R1138_U203, R1138_U204, R1138_U205, R1138_U206, R1138_U207, R1138_U208, R1138_U209, R1138_U21, R1138_U210, R1138_U211, R1138_U212, R1138_U213, R1138_U214, R1138_U215, R1138_U216, R1138_U217, R1138_U218, R1138_U219, R1138_U22, R1138_U220, R1138_U221, R1138_U222, R1138_U223, R1138_U224, R1138_U225, R1138_U226, R1138_U227, R1138_U228, R1138_U229, R1138_U23, R1138_U230, R1138_U231, R1138_U232, R1138_U233, R1138_U234, R1138_U235, R1138_U236, R1138_U237, R1138_U238, R1138_U239, R1138_U24, R1138_U240, R1138_U241, R1138_U242, R1138_U243, R1138_U244, R1138_U245, R1138_U246, R1138_U247, R1138_U248, R1138_U249, R1138_U25, R1138_U250, R1138_U251, R1138_U252, R1138_U253, R1138_U254, R1138_U255, R1138_U256, R1138_U257, R1138_U258, R1138_U259, R1138_U26, R1138_U260, R1138_U261, R1138_U262, R1138_U263, R1138_U264, R1138_U265, R1138_U266, R1138_U267, R1138_U268, R1138_U269, R1138_U27, R1138_U270, R1138_U271, R1138_U272, R1138_U273, R1138_U274, R1138_U275, R1138_U276, R1138_U277, R1138_U278, R1138_U279, R1138_U28, R1138_U280, R1138_U281, R1138_U282, R1138_U283, R1138_U284, R1138_U285, R1138_U286, R1138_U287, R1138_U288, R1138_U289, R1138_U29, R1138_U290, R1138_U291, R1138_U292, R1138_U293, R1138_U294, R1138_U295, R1138_U296, R1138_U297, R1138_U298, R1138_U299, R1138_U30, R1138_U300, R1138_U301, R1138_U302, R1138_U303, R1138_U304, R1138_U305, R1138_U306, R1138_U307, R1138_U308, R1138_U309, R1138_U31, R1138_U310, R1138_U311, R1138_U312, R1138_U313, R1138_U314, R1138_U315, R1138_U316, R1138_U317, R1138_U318, R1138_U319, R1138_U32, R1138_U320, R1138_U321, R1138_U322, R1138_U323, R1138_U324, R1138_U325, R1138_U326, R1138_U327, R1138_U328, R1138_U329, R1138_U33, R1138_U330, R1138_U331, R1138_U332, R1138_U333, R1138_U334, R1138_U335, R1138_U336, R1138_U337, R1138_U338, R1138_U339, R1138_U34, R1138_U340, R1138_U341, R1138_U342, R1138_U343, R1138_U344, R1138_U345, R1138_U346, R1138_U347, R1138_U348, R1138_U349, R1138_U35, R1138_U350, R1138_U351, R1138_U352, R1138_U353, R1138_U354, R1138_U355, R1138_U356, R1138_U357, R1138_U358, R1138_U359, R1138_U36, R1138_U360, R1138_U361, R1138_U362, R1138_U363, R1138_U364, R1138_U365, R1138_U366, R1138_U367, R1138_U368, R1138_U369, R1138_U37, R1138_U370, R1138_U371, R1138_U372, R1138_U373, R1138_U374, R1138_U375, R1138_U376, R1138_U377, R1138_U378, R1138_U379, R1138_U38, R1138_U380, R1138_U381, R1138_U382, R1138_U383, R1138_U384, R1138_U385, R1138_U386, R1138_U387, R1138_U388, R1138_U389, R1138_U39, R1138_U390, R1138_U391, R1138_U392, R1138_U393, R1138_U394, R1138_U395, R1138_U396, R1138_U397, R1138_U398, R1138_U399, R1138_U4, R1138_U40, R1138_U400, R1138_U401, R1138_U402, R1138_U403, R1138_U404, R1138_U405, R1138_U406, R1138_U407, R1138_U408, R1138_U409, R1138_U41, R1138_U410, R1138_U411, R1138_U412, R1138_U413, R1138_U414, R1138_U415, R1138_U416, R1138_U417, R1138_U418, R1138_U419, R1138_U42, R1138_U420, R1138_U421, R1138_U422, R1138_U423, R1138_U424, R1138_U425, R1138_U426, R1138_U427, R1138_U428, R1138_U429, R1138_U43, R1138_U430, R1138_U431, R1138_U432, R1138_U433, R1138_U434, R1138_U435, R1138_U436, R1138_U437, R1138_U438, R1138_U439, R1138_U44, R1138_U440, R1138_U441, R1138_U442, R1138_U443, R1138_U444, R1138_U445, R1138_U446, R1138_U447, R1138_U448, R1138_U449, R1138_U45, R1138_U450, R1138_U451, R1138_U452, R1138_U453, R1138_U454, R1138_U455, R1138_U456, R1138_U457, R1138_U458, R1138_U459, R1138_U46, R1138_U460, R1138_U461, R1138_U462, R1138_U463, R1138_U464, R1138_U465, R1138_U466, R1138_U467, R1138_U468, R1138_U469, R1138_U47, R1138_U470, R1138_U471, R1138_U472, R1138_U473, R1138_U474, R1138_U475, R1138_U476, R1138_U477, R1138_U478, R1138_U479, R1138_U48, R1138_U480, R1138_U481, R1138_U482, R1138_U483, R1138_U484, R1138_U485, R1138_U486, R1138_U487, R1138_U488, R1138_U489, R1138_U49, R1138_U490, R1138_U491, R1138_U492, R1138_U493, R1138_U494, R1138_U495, R1138_U496, R1138_U497, R1138_U498, R1138_U499, R1138_U5, R1138_U50, R1138_U500, R1138_U501, R1138_U502, R1138_U503, R1138_U504, R1138_U505, R1138_U506, R1138_U507, R1138_U508, R1138_U509, R1138_U51, R1138_U510, R1138_U511, R1138_U512, R1138_U513, R1138_U514, R1138_U515, R1138_U516, R1138_U517, R1138_U518, R1138_U519, R1138_U52, R1138_U520, R1138_U521, R1138_U522, R1138_U523, R1138_U524, R1138_U525, R1138_U526, R1138_U527, R1138_U528, R1138_U529, R1138_U53, R1138_U530, R1138_U531, R1138_U54, R1138_U55, R1138_U56, R1138_U57, R1138_U58, R1138_U59, R1138_U6, R1138_U60, R1138_U61, R1138_U62, R1138_U63, R1138_U64, R1138_U65, R1138_U66, R1138_U67, R1138_U68, R1138_U69, R1138_U7, R1138_U70, R1138_U71, R1138_U72, R1138_U73, R1138_U74, R1138_U75, R1138_U76, R1138_U77, R1138_U78, R1138_U79, R1138_U8, R1138_U80, R1138_U81, R1138_U82, R1138_U83, R1138_U84, R1138_U85, R1138_U86, R1138_U87, R1138_U88, R1138_U89, R1138_U9, R1138_U90, R1138_U91, R1138_U92, R1138_U93, R1138_U94, R1138_U95, R1138_U96, R1138_U97, R1138_U98, R1138_U99, R1150_U10, R1150_U100, R1150_U101, R1150_U102, R1150_U103, R1150_U104, R1150_U105, R1150_U106, R1150_U107, R1150_U108, R1150_U109, R1150_U11, R1150_U110, R1150_U111, R1150_U112, R1150_U113, R1150_U114, R1150_U115, R1150_U116, R1150_U117, R1150_U118, R1150_U119, R1150_U12, R1150_U120, R1150_U121, R1150_U122, R1150_U123, R1150_U124, R1150_U125, R1150_U126, R1150_U127, R1150_U128, R1150_U129, R1150_U13, R1150_U130, R1150_U131, R1150_U132, R1150_U133, R1150_U134, R1150_U135, R1150_U136, R1150_U137, R1150_U138, R1150_U139, R1150_U14, R1150_U140, R1150_U141, R1150_U142, R1150_U143, R1150_U144, R1150_U145, R1150_U146, R1150_U147, R1150_U148, R1150_U149, R1150_U15, R1150_U150, R1150_U151, R1150_U152, R1150_U153, R1150_U154, R1150_U155, R1150_U156, R1150_U157, R1150_U158, R1150_U159, R1150_U16, R1150_U160, R1150_U161, R1150_U162, R1150_U163, R1150_U164, R1150_U165, R1150_U166, R1150_U167, R1150_U168, R1150_U169, R1150_U17, R1150_U170, R1150_U171, R1150_U172, R1150_U173, R1150_U174, R1150_U175, R1150_U176, R1150_U177, R1150_U178, R1150_U179, R1150_U18, R1150_U180, R1150_U181, R1150_U182, R1150_U183, R1150_U184, R1150_U185, R1150_U186, R1150_U187, R1150_U188, R1150_U189, R1150_U19, R1150_U190, R1150_U191, R1150_U192, R1150_U193, R1150_U194, R1150_U195, R1150_U196, R1150_U197, R1150_U198, R1150_U199, R1150_U20, R1150_U200, R1150_U201, R1150_U202, R1150_U203, R1150_U204, R1150_U205, R1150_U206, R1150_U207, R1150_U208, R1150_U209, R1150_U21, R1150_U210, R1150_U211, R1150_U212, R1150_U213, R1150_U214, R1150_U215, R1150_U216, R1150_U217, R1150_U218, R1150_U219, R1150_U22, R1150_U220, R1150_U221, R1150_U222, R1150_U223, R1150_U224, R1150_U225, R1150_U226, R1150_U227, R1150_U228, R1150_U229, R1150_U23, R1150_U230, R1150_U231, R1150_U232, R1150_U233, R1150_U234, R1150_U235, R1150_U236, R1150_U237, R1150_U238, R1150_U239, R1150_U24, R1150_U240, R1150_U241, R1150_U242, R1150_U243, R1150_U244, R1150_U245, R1150_U246, R1150_U247, R1150_U248, R1150_U249, R1150_U25, R1150_U250, R1150_U251, R1150_U252, R1150_U253, R1150_U254, R1150_U255, R1150_U256, R1150_U257, R1150_U258, R1150_U259, R1150_U26, R1150_U260, R1150_U261, R1150_U262, R1150_U263, R1150_U264, R1150_U265, R1150_U266, R1150_U267, R1150_U268, R1150_U269, R1150_U27, R1150_U270, R1150_U271, R1150_U272, R1150_U273, R1150_U274, R1150_U275, R1150_U276, R1150_U277, R1150_U278, R1150_U279, R1150_U28, R1150_U280, R1150_U281, R1150_U282, R1150_U283, R1150_U284, R1150_U285, R1150_U286, R1150_U287, R1150_U288, R1150_U289, R1150_U29, R1150_U290, R1150_U291, R1150_U292, R1150_U293, R1150_U294, R1150_U295, R1150_U296, R1150_U297, R1150_U298, R1150_U299, R1150_U30, R1150_U300, R1150_U301, R1150_U302, R1150_U303, R1150_U304, R1150_U305, R1150_U306, R1150_U307, R1150_U308, R1150_U309, R1150_U31, R1150_U310, R1150_U311, R1150_U312, R1150_U313, R1150_U314, R1150_U315, R1150_U316, R1150_U317, R1150_U318, R1150_U319, R1150_U32, R1150_U320, R1150_U321, R1150_U322, R1150_U323, R1150_U324, R1150_U325, R1150_U326, R1150_U327, R1150_U328, R1150_U329, R1150_U33, R1150_U330, R1150_U331, R1150_U332, R1150_U333, R1150_U334, R1150_U335, R1150_U336, R1150_U337, R1150_U338, R1150_U339, R1150_U34, R1150_U340, R1150_U341, R1150_U342, R1150_U343, R1150_U344, R1150_U345, R1150_U346, R1150_U347, R1150_U348, R1150_U349, R1150_U35, R1150_U350, R1150_U351, R1150_U352, R1150_U353, R1150_U354, R1150_U355, R1150_U356, R1150_U357, R1150_U358, R1150_U359, R1150_U36, R1150_U360, R1150_U361, R1150_U362, R1150_U363, R1150_U364, R1150_U365, R1150_U366, R1150_U367, R1150_U368, R1150_U369, R1150_U37, R1150_U370, R1150_U371, R1150_U372, R1150_U373, R1150_U374, R1150_U375, R1150_U376, R1150_U377, R1150_U378, R1150_U379, R1150_U38, R1150_U380, R1150_U381, R1150_U382, R1150_U383, R1150_U384, R1150_U385, R1150_U386, R1150_U387, R1150_U388, R1150_U389, R1150_U39, R1150_U390, R1150_U391, R1150_U392, R1150_U393, R1150_U394, R1150_U395, R1150_U396, R1150_U397, R1150_U398, R1150_U399, R1150_U40, R1150_U400, R1150_U401, R1150_U402, R1150_U403, R1150_U404, R1150_U405, R1150_U406, R1150_U407, R1150_U408, R1150_U409, R1150_U41, R1150_U410, R1150_U411, R1150_U412, R1150_U413, R1150_U414, R1150_U415, R1150_U416, R1150_U417, R1150_U418, R1150_U419, R1150_U42, R1150_U420, R1150_U421, R1150_U422, R1150_U423, R1150_U424, R1150_U425, R1150_U426, R1150_U427, R1150_U428, R1150_U429, R1150_U43, R1150_U430, R1150_U431, R1150_U432, R1150_U433, R1150_U434, R1150_U435, R1150_U436, R1150_U437, R1150_U438, R1150_U439, R1150_U44, R1150_U440, R1150_U441, R1150_U442, R1150_U443, R1150_U444, R1150_U445, R1150_U446, R1150_U447, R1150_U448, R1150_U449, R1150_U45, R1150_U450, R1150_U451, R1150_U452, R1150_U453, R1150_U454, R1150_U455, R1150_U456, R1150_U457, R1150_U458, R1150_U459, R1150_U46, R1150_U460, R1150_U461, R1150_U462, R1150_U463, R1150_U464, R1150_U465, R1150_U466, R1150_U467, R1150_U468, R1150_U469, R1150_U47, R1150_U470, R1150_U471, R1150_U472, R1150_U473, R1150_U474, R1150_U475, R1150_U476, R1150_U477, R1150_U478, R1150_U479, R1150_U48, R1150_U480, R1150_U481, R1150_U482, R1150_U483, R1150_U484, R1150_U485, R1150_U486, R1150_U487, R1150_U488, R1150_U489, R1150_U49, R1150_U490, R1150_U491, R1150_U492, R1150_U493, R1150_U494, R1150_U495, R1150_U496, R1150_U497, R1150_U498, R1150_U499, R1150_U50, R1150_U500, R1150_U501, R1150_U502, R1150_U503, R1150_U504, R1150_U505, R1150_U506, R1150_U507, R1150_U508, R1150_U509, R1150_U51, R1150_U510, R1150_U511, R1150_U52, R1150_U53, R1150_U54, R1150_U55, R1150_U56, R1150_U57, R1150_U58, R1150_U59, R1150_U6, R1150_U60, R1150_U61, R1150_U62, R1150_U63, R1150_U64, R1150_U65, R1150_U66, R1150_U67, R1150_U68, R1150_U69, R1150_U7, R1150_U70, R1150_U71, R1150_U72, R1150_U73, R1150_U74, R1150_U75, R1150_U76, R1150_U77, R1150_U78, R1150_U79, R1150_U8, R1150_U80, R1150_U81, R1150_U82, R1150_U83, R1150_U84, R1150_U85, R1150_U86, R1150_U87, R1150_U88, R1150_U89, R1150_U9, R1150_U90, R1150_U91, R1150_U92, R1150_U93, R1150_U94, R1150_U95, R1150_U96, R1150_U97, R1150_U98, R1150_U99, R1162_U10, R1162_U100, R1162_U101, R1162_U102, R1162_U103, R1162_U104, R1162_U105, R1162_U106, R1162_U107, R1162_U108, R1162_U109, R1162_U11, R1162_U110, R1162_U111, R1162_U112, R1162_U113, R1162_U114, R1162_U115, R1162_U116, R1162_U117, R1162_U118, R1162_U119, R1162_U12, R1162_U120, R1162_U121, R1162_U122, R1162_U123, R1162_U124, R1162_U125, R1162_U126, R1162_U127, R1162_U128, R1162_U129, R1162_U13, R1162_U130, R1162_U131, R1162_U132, R1162_U133, R1162_U134, R1162_U135, R1162_U136, R1162_U137, R1162_U138, R1162_U139, R1162_U14, R1162_U140, R1162_U141, R1162_U142, R1162_U143, R1162_U144, R1162_U145, R1162_U146, R1162_U147, R1162_U148, R1162_U149, R1162_U15, R1162_U150, R1162_U151, R1162_U152, R1162_U153, R1162_U154, R1162_U155, R1162_U156, R1162_U157, R1162_U158, R1162_U159, R1162_U16, R1162_U160, R1162_U161, R1162_U162, R1162_U163, R1162_U164, R1162_U165, R1162_U166, R1162_U167, R1162_U168, R1162_U169, R1162_U17, R1162_U170, R1162_U171, R1162_U172, R1162_U173, R1162_U174, R1162_U175, R1162_U176, R1162_U177, R1162_U178, R1162_U179, R1162_U18, R1162_U180, R1162_U181, R1162_U182, R1162_U183, R1162_U184, R1162_U185, R1162_U186, R1162_U187, R1162_U188, R1162_U189, R1162_U19, R1162_U190, R1162_U191, R1162_U192, R1162_U193, R1162_U194, R1162_U195, R1162_U196, R1162_U197, R1162_U198, R1162_U199, R1162_U20, R1162_U200, R1162_U201, R1162_U202, R1162_U203, R1162_U204, R1162_U205, R1162_U206, R1162_U207, R1162_U208, R1162_U209, R1162_U21, R1162_U210, R1162_U211, R1162_U212, R1162_U213, R1162_U214, R1162_U215, R1162_U216, R1162_U217, R1162_U218, R1162_U219, R1162_U22, R1162_U220, R1162_U221, R1162_U222, R1162_U223, R1162_U224, R1162_U225, R1162_U226, R1162_U227, R1162_U228, R1162_U229, R1162_U23, R1162_U230, R1162_U231, R1162_U232, R1162_U233, R1162_U234, R1162_U235, R1162_U236, R1162_U237, R1162_U238, R1162_U239, R1162_U24, R1162_U240, R1162_U241, R1162_U242, R1162_U243, R1162_U244, R1162_U245, R1162_U246, R1162_U247, R1162_U248, R1162_U249, R1162_U25, R1162_U250, R1162_U251, R1162_U252, R1162_U253, R1162_U254, R1162_U255, R1162_U256, R1162_U257, R1162_U258, R1162_U259, R1162_U26, R1162_U260, R1162_U261, R1162_U262, R1162_U263, R1162_U264, R1162_U265, R1162_U266, R1162_U267, R1162_U268, R1162_U269, R1162_U27, R1162_U270, R1162_U271, R1162_U272, R1162_U273, R1162_U274, R1162_U275, R1162_U276, R1162_U277, R1162_U278, R1162_U279, R1162_U28, R1162_U280, R1162_U281, R1162_U282, R1162_U283, R1162_U284, R1162_U285, R1162_U286, R1162_U287, R1162_U288, R1162_U289, R1162_U29, R1162_U290, R1162_U30, R1162_U31, R1162_U32, R1162_U33, R1162_U34, R1162_U35, R1162_U36, R1162_U37, R1162_U38, R1162_U39, R1162_U4, R1162_U40, R1162_U41, R1162_U42, R1162_U43, R1162_U44, R1162_U45, R1162_U46, R1162_U47, R1162_U48, R1162_U49, R1162_U5, R1162_U50, R1162_U51, R1162_U52, R1162_U53, R1162_U54, R1162_U55, R1162_U56, R1162_U57, R1162_U58, R1162_U59, R1162_U6, R1162_U60, R1162_U61, R1162_U62, R1162_U63, R1162_U64, R1162_U65, R1162_U66, R1162_U67, R1162_U68, R1162_U69, R1162_U7, R1162_U70, R1162_U71, R1162_U72, R1162_U73, R1162_U74, R1162_U75, R1162_U76, R1162_U77, R1162_U78, R1162_U79, R1162_U8, R1162_U80, R1162_U81, R1162_U82, R1162_U83, R1162_U84, R1162_U85, R1162_U86, R1162_U87, R1162_U88, R1162_U89, R1162_U9, R1162_U90, R1162_U91, R1162_U92, R1162_U93, R1162_U94, R1162_U95, R1162_U96, R1162_U97, R1162_U98, R1162_U99, R1165_U10, R1165_U100, R1165_U101, R1165_U102, R1165_U103, R1165_U104, R1165_U105, R1165_U106, R1165_U107, R1165_U108, R1165_U109, R1165_U11, R1165_U110, R1165_U111, R1165_U112, R1165_U113, R1165_U114, R1165_U115, R1165_U116, R1165_U117, R1165_U118, R1165_U119, R1165_U12, R1165_U120, R1165_U121, R1165_U122, R1165_U123, R1165_U124, R1165_U125, R1165_U126, R1165_U127, R1165_U128, R1165_U129, R1165_U13, R1165_U130, R1165_U131, R1165_U132, R1165_U133, R1165_U134, R1165_U135, R1165_U136, R1165_U137, R1165_U138, R1165_U139, R1165_U14, R1165_U140, R1165_U141, R1165_U142, R1165_U143, R1165_U144, R1165_U145, R1165_U146, R1165_U147, R1165_U148, R1165_U149, R1165_U15, R1165_U150, R1165_U151, R1165_U152, R1165_U153, R1165_U154, R1165_U155, R1165_U156, R1165_U157, R1165_U158, R1165_U159, R1165_U16, R1165_U160, R1165_U161, R1165_U162, R1165_U163, R1165_U164, R1165_U165, R1165_U166, R1165_U167, R1165_U168, R1165_U169, R1165_U17, R1165_U170, R1165_U171, R1165_U172, R1165_U173, R1165_U174, R1165_U175, R1165_U176, R1165_U177, R1165_U178, R1165_U179, R1165_U18, R1165_U180, R1165_U181, R1165_U182, R1165_U183, R1165_U184, R1165_U185, R1165_U186, R1165_U187, R1165_U188, R1165_U189, R1165_U19, R1165_U190, R1165_U191, R1165_U192, R1165_U193, R1165_U194, R1165_U195, R1165_U196, R1165_U197, R1165_U198, R1165_U199, R1165_U20, R1165_U200, R1165_U201, R1165_U202, R1165_U203, R1165_U204, R1165_U205, R1165_U206, R1165_U207, R1165_U208, R1165_U209, R1165_U21, R1165_U210, R1165_U211, R1165_U212, R1165_U213, R1165_U214, R1165_U215, R1165_U216, R1165_U217, R1165_U218, R1165_U219, R1165_U22, R1165_U220, R1165_U221, R1165_U222, R1165_U223, R1165_U224, R1165_U225, R1165_U226, R1165_U227, R1165_U228, R1165_U229, R1165_U23, R1165_U230, R1165_U231, R1165_U232, R1165_U233, R1165_U234, R1165_U235, R1165_U236, R1165_U237, R1165_U238, R1165_U239, R1165_U24, R1165_U240, R1165_U241, R1165_U242, R1165_U243, R1165_U244, R1165_U245, R1165_U246, R1165_U247, R1165_U248, R1165_U249, R1165_U25, R1165_U250, R1165_U251, R1165_U252, R1165_U253, R1165_U254, R1165_U255, R1165_U256, R1165_U257, R1165_U258, R1165_U259, R1165_U26, R1165_U260, R1165_U261, R1165_U262, R1165_U263, R1165_U264, R1165_U265, R1165_U266, R1165_U267, R1165_U268, R1165_U269, R1165_U27, R1165_U270, R1165_U271, R1165_U272, R1165_U273, R1165_U274, R1165_U275, R1165_U276, R1165_U277, R1165_U278, R1165_U279, R1165_U28, R1165_U280, R1165_U281, R1165_U282, R1165_U283, R1165_U284, R1165_U285, R1165_U286, R1165_U287, R1165_U288, R1165_U289, R1165_U29, R1165_U290, R1165_U291, R1165_U292, R1165_U293, R1165_U294, R1165_U295, R1165_U296, R1165_U297, R1165_U298, R1165_U299, R1165_U30, R1165_U300, R1165_U301, R1165_U302, R1165_U303, R1165_U304, R1165_U305, R1165_U306, R1165_U307, R1165_U308, R1165_U309, R1165_U31, R1165_U310, R1165_U311, R1165_U312, R1165_U313, R1165_U314, R1165_U315, R1165_U316, R1165_U317, R1165_U318, R1165_U319, R1165_U32, R1165_U320, R1165_U321, R1165_U322, R1165_U323, R1165_U324, R1165_U325, R1165_U326, R1165_U327, R1165_U328, R1165_U329, R1165_U33, R1165_U330, R1165_U331, R1165_U332, R1165_U333, R1165_U334, R1165_U335, R1165_U336, R1165_U337, R1165_U338, R1165_U339, R1165_U34, R1165_U340, R1165_U341, R1165_U342, R1165_U343, R1165_U344, R1165_U345, R1165_U346, R1165_U347, R1165_U348, R1165_U349, R1165_U35, R1165_U350, R1165_U351, R1165_U352, R1165_U353, R1165_U354, R1165_U355, R1165_U356, R1165_U357, R1165_U358, R1165_U359, R1165_U36, R1165_U360, R1165_U361, R1165_U362, R1165_U363, R1165_U364, R1165_U365, R1165_U366, R1165_U367, R1165_U368, R1165_U369, R1165_U37, R1165_U370, R1165_U371, R1165_U372, R1165_U373, R1165_U374, R1165_U375, R1165_U376, R1165_U377, R1165_U378, R1165_U379, R1165_U38, R1165_U380, R1165_U381, R1165_U382, R1165_U383, R1165_U384, R1165_U385, R1165_U386, R1165_U387, R1165_U388, R1165_U389, R1165_U39, R1165_U390, R1165_U391, R1165_U392, R1165_U393, R1165_U394, R1165_U395, R1165_U396, R1165_U397, R1165_U398, R1165_U399, R1165_U4, R1165_U40, R1165_U400, R1165_U401, R1165_U402, R1165_U403, R1165_U404, R1165_U405, R1165_U406, R1165_U407, R1165_U408, R1165_U409, R1165_U41, R1165_U410, R1165_U411, R1165_U412, R1165_U413, R1165_U414, R1165_U415, R1165_U416, R1165_U417, R1165_U418, R1165_U419, R1165_U42, R1165_U420, R1165_U421, R1165_U422, R1165_U423, R1165_U424, R1165_U425, R1165_U426, R1165_U427, R1165_U428, R1165_U429, R1165_U43, R1165_U430, R1165_U431, R1165_U432, R1165_U433, R1165_U434, R1165_U435, R1165_U436, R1165_U437, R1165_U438, R1165_U439, R1165_U44, R1165_U440, R1165_U441, R1165_U442, R1165_U443, R1165_U444, R1165_U445, R1165_U446, R1165_U447, R1165_U448, R1165_U449, R1165_U45, R1165_U450, R1165_U451, R1165_U452, R1165_U453, R1165_U454, R1165_U455, R1165_U456, R1165_U457, R1165_U458, R1165_U459, R1165_U46, R1165_U460, R1165_U461, R1165_U462, R1165_U463, R1165_U464, R1165_U465, R1165_U466, R1165_U467, R1165_U468, R1165_U469, R1165_U47, R1165_U470, R1165_U471, R1165_U472, R1165_U473, R1165_U474, R1165_U475, R1165_U476, R1165_U477, R1165_U478, R1165_U479, R1165_U48, R1165_U480, R1165_U481, R1165_U482, R1165_U483, R1165_U484, R1165_U485, R1165_U486, R1165_U487, R1165_U488, R1165_U489, R1165_U49, R1165_U490, R1165_U491, R1165_U492, R1165_U493, R1165_U494, R1165_U495, R1165_U496, R1165_U497, R1165_U498, R1165_U499, R1165_U5, R1165_U50, R1165_U500, R1165_U501, R1165_U502, R1165_U503, R1165_U504, R1165_U505, R1165_U506, R1165_U507, R1165_U508, R1165_U509, R1165_U51, R1165_U510, R1165_U511, R1165_U512, R1165_U513, R1165_U514, R1165_U515, R1165_U516, R1165_U517, R1165_U518, R1165_U519, R1165_U52, R1165_U520, R1165_U521, R1165_U522, R1165_U523, R1165_U524, R1165_U525, R1165_U526, R1165_U527, R1165_U528, R1165_U529, R1165_U53, R1165_U530, R1165_U531, R1165_U532, R1165_U533, R1165_U534, R1165_U535, R1165_U536, R1165_U537, R1165_U538, R1165_U539, R1165_U54, R1165_U540, R1165_U541, R1165_U542, R1165_U543, R1165_U544, R1165_U545, R1165_U546, R1165_U547, R1165_U548, R1165_U549, R1165_U55, R1165_U550, R1165_U551, R1165_U552, R1165_U553, R1165_U554, R1165_U555, R1165_U556, R1165_U557, R1165_U558, R1165_U559, R1165_U56, R1165_U560, R1165_U561, R1165_U562, R1165_U563, R1165_U564, R1165_U565, R1165_U566, R1165_U567, R1165_U568, R1165_U569, R1165_U57, R1165_U570, R1165_U571, R1165_U572, R1165_U573, R1165_U574, R1165_U575, R1165_U576, R1165_U577, R1165_U578, R1165_U579, R1165_U58, R1165_U580, R1165_U581, R1165_U582, R1165_U583, R1165_U584, R1165_U585, R1165_U586, R1165_U587, R1165_U588, R1165_U589, R1165_U59, R1165_U590, R1165_U591, R1165_U592, R1165_U593, R1165_U594, R1165_U595, R1165_U596, R1165_U597, R1165_U598, R1165_U599, R1165_U6, R1165_U60, R1165_U600, R1165_U601, R1165_U602, R1165_U603, R1165_U604, R1165_U605, R1165_U606, R1165_U607, R1165_U608, R1165_U609, R1165_U61, R1165_U610, R1165_U611, R1165_U612, R1165_U613, R1165_U62, R1165_U63, R1165_U64, R1165_U65, R1165_U66, R1165_U67, R1165_U68, R1165_U69, R1165_U7, R1165_U70, R1165_U71, R1165_U72, R1165_U73, R1165_U74, R1165_U75, R1165_U76, R1165_U77, R1165_U78, R1165_U79, R1165_U8, R1165_U80, R1165_U81, R1165_U82, R1165_U83, R1165_U84, R1165_U85, R1165_U86, R1165_U87, R1165_U88, R1165_U89, R1165_U9, R1165_U90, R1165_U91, R1165_U92, R1165_U93, R1165_U94, R1165_U95, R1165_U96, R1165_U97, R1165_U98, R1165_U99, R1171_U10, R1171_U100, R1171_U101, R1171_U102, R1171_U103, R1171_U104, R1171_U105, R1171_U106, R1171_U107, R1171_U108, R1171_U109, R1171_U11, R1171_U110, R1171_U111, R1171_U112, R1171_U113, R1171_U114, R1171_U115, R1171_U116, R1171_U117, R1171_U118, R1171_U119, R1171_U12, R1171_U120, R1171_U121, R1171_U122, R1171_U123, R1171_U124, R1171_U125, R1171_U126, R1171_U127, R1171_U128, R1171_U129, R1171_U13, R1171_U130, R1171_U131, R1171_U132, R1171_U133, R1171_U134, R1171_U135, R1171_U136, R1171_U137, R1171_U138, R1171_U139, R1171_U14, R1171_U140, R1171_U141, R1171_U142, R1171_U143, R1171_U144, R1171_U145, R1171_U146, R1171_U147, R1171_U148, R1171_U149, R1171_U15, R1171_U150, R1171_U151, R1171_U152, R1171_U153, R1171_U154, R1171_U155, R1171_U156, R1171_U157, R1171_U158, R1171_U159, R1171_U16, R1171_U160, R1171_U161, R1171_U162, R1171_U163, R1171_U164, R1171_U165, R1171_U166, R1171_U167, R1171_U168, R1171_U169, R1171_U17, R1171_U170, R1171_U171, R1171_U172, R1171_U173, R1171_U174, R1171_U175, R1171_U176, R1171_U177, R1171_U178, R1171_U179, R1171_U18, R1171_U180, R1171_U181, R1171_U182, R1171_U183, R1171_U184, R1171_U185, R1171_U186, R1171_U187, R1171_U188, R1171_U189, R1171_U19, R1171_U190, R1171_U191, R1171_U192, R1171_U193, R1171_U194, R1171_U195, R1171_U196, R1171_U197, R1171_U198, R1171_U199, R1171_U20, R1171_U200, R1171_U201, R1171_U202, R1171_U203, R1171_U204, R1171_U205, R1171_U206, R1171_U207, R1171_U208, R1171_U209, R1171_U21, R1171_U210, R1171_U211, R1171_U212, R1171_U213, R1171_U214, R1171_U215, R1171_U216, R1171_U217, R1171_U218, R1171_U219, R1171_U22, R1171_U220, R1171_U221, R1171_U222, R1171_U223, R1171_U224, R1171_U225, R1171_U226, R1171_U227, R1171_U228, R1171_U229, R1171_U23, R1171_U230, R1171_U231, R1171_U232, R1171_U233, R1171_U234, R1171_U235, R1171_U236, R1171_U237, R1171_U238, R1171_U239, R1171_U24, R1171_U240, R1171_U241, R1171_U242, R1171_U243, R1171_U244, R1171_U245, R1171_U246, R1171_U247, R1171_U248, R1171_U249, R1171_U25, R1171_U250, R1171_U251, R1171_U252, R1171_U253, R1171_U254, R1171_U255, R1171_U256, R1171_U257, R1171_U258, R1171_U259, R1171_U26, R1171_U260, R1171_U261, R1171_U262, R1171_U263, R1171_U264, R1171_U265, R1171_U266, R1171_U267, R1171_U268, R1171_U269, R1171_U27, R1171_U270, R1171_U271, R1171_U272, R1171_U273, R1171_U274, R1171_U275, R1171_U276, R1171_U277, R1171_U278, R1171_U279, R1171_U28, R1171_U280, R1171_U281, R1171_U282, R1171_U283, R1171_U284, R1171_U285, R1171_U286, R1171_U287, R1171_U288, R1171_U289, R1171_U29, R1171_U290, R1171_U291, R1171_U292, R1171_U293, R1171_U294, R1171_U295, R1171_U296, R1171_U297, R1171_U298, R1171_U299, R1171_U30, R1171_U300, R1171_U301, R1171_U302, R1171_U303, R1171_U304, R1171_U305, R1171_U306, R1171_U307, R1171_U308, R1171_U309, R1171_U31, R1171_U310, R1171_U311, R1171_U312, R1171_U313, R1171_U314, R1171_U315, R1171_U316, R1171_U317, R1171_U318, R1171_U319, R1171_U32, R1171_U320, R1171_U321, R1171_U322, R1171_U323, R1171_U324, R1171_U325, R1171_U326, R1171_U327, R1171_U328, R1171_U329, R1171_U33, R1171_U330, R1171_U331, R1171_U332, R1171_U333, R1171_U334, R1171_U335, R1171_U336, R1171_U337, R1171_U338, R1171_U339, R1171_U34, R1171_U340, R1171_U341, R1171_U342, R1171_U343, R1171_U344, R1171_U345, R1171_U346, R1171_U347, R1171_U348, R1171_U349, R1171_U35, R1171_U350, R1171_U351, R1171_U352, R1171_U353, R1171_U354, R1171_U355, R1171_U356, R1171_U357, R1171_U358, R1171_U359, R1171_U36, R1171_U360, R1171_U361, R1171_U362, R1171_U363, R1171_U364, R1171_U365, R1171_U366, R1171_U367, R1171_U368, R1171_U369, R1171_U37, R1171_U370, R1171_U371, R1171_U372, R1171_U373, R1171_U374, R1171_U375, R1171_U376, R1171_U377, R1171_U378, R1171_U379, R1171_U38, R1171_U380, R1171_U381, R1171_U382, R1171_U383, R1171_U384, R1171_U385, R1171_U386, R1171_U387, R1171_U388, R1171_U389, R1171_U39, R1171_U390, R1171_U391, R1171_U392, R1171_U393, R1171_U394, R1171_U395, R1171_U396, R1171_U397, R1171_U398, R1171_U399, R1171_U4, R1171_U40, R1171_U400, R1171_U401, R1171_U402, R1171_U403, R1171_U404, R1171_U405, R1171_U406, R1171_U407, R1171_U408, R1171_U409, R1171_U41, R1171_U410, R1171_U411, R1171_U412, R1171_U413, R1171_U414, R1171_U415, R1171_U416, R1171_U417, R1171_U418, R1171_U419, R1171_U42, R1171_U420, R1171_U421, R1171_U422, R1171_U423, R1171_U424, R1171_U425, R1171_U426, R1171_U427, R1171_U428, R1171_U429, R1171_U43, R1171_U430, R1171_U431, R1171_U432, R1171_U433, R1171_U434, R1171_U435, R1171_U436, R1171_U437, R1171_U438, R1171_U439, R1171_U44, R1171_U440, R1171_U441, R1171_U442, R1171_U443, R1171_U444, R1171_U445, R1171_U446, R1171_U447, R1171_U448, R1171_U449, R1171_U45, R1171_U450, R1171_U451, R1171_U452, R1171_U453, R1171_U454, R1171_U455, R1171_U456, R1171_U457, R1171_U458, R1171_U459, R1171_U46, R1171_U460, R1171_U461, R1171_U462, R1171_U463, R1171_U464, R1171_U465, R1171_U466, R1171_U467, R1171_U468, R1171_U469, R1171_U47, R1171_U470, R1171_U471, R1171_U472, R1171_U473, R1171_U474, R1171_U475, R1171_U476, R1171_U477, R1171_U478, R1171_U479, R1171_U48, R1171_U480, R1171_U481, R1171_U482, R1171_U483, R1171_U484, R1171_U485, R1171_U486, R1171_U487, R1171_U488, R1171_U489, R1171_U49, R1171_U490, R1171_U491, R1171_U492, R1171_U493, R1171_U494, R1171_U495, R1171_U496, R1171_U497, R1171_U498, R1171_U499, R1171_U5, R1171_U50, R1171_U500, R1171_U501, R1171_U502, R1171_U503, R1171_U504, R1171_U505, R1171_U506, R1171_U507, R1171_U508, R1171_U509, R1171_U51, R1171_U510, R1171_U511, R1171_U512, R1171_U513, R1171_U514, R1171_U515, R1171_U516, R1171_U517, R1171_U518, R1171_U519, R1171_U52, R1171_U520, R1171_U521, R1171_U522, R1171_U523, R1171_U524, R1171_U525, R1171_U526, R1171_U527, R1171_U528, R1171_U529, R1171_U53, R1171_U530, R1171_U531, R1171_U54, R1171_U55, R1171_U56, R1171_U57, R1171_U58, R1171_U59, R1171_U6, R1171_U60, R1171_U61, R1171_U62, R1171_U63, R1171_U64, R1171_U65, R1171_U66, R1171_U67, R1171_U68, R1171_U69, R1171_U7, R1171_U70, R1171_U71, R1171_U72, R1171_U73, R1171_U74, R1171_U75, R1171_U76, R1171_U77, R1171_U78, R1171_U79, R1171_U8, R1171_U80, R1171_U81, R1171_U82, R1171_U83, R1171_U84, R1171_U85, R1171_U86, R1171_U87, R1171_U88, R1171_U89, R1171_U9, R1171_U90, R1171_U91, R1171_U92, R1171_U93, R1171_U94, R1171_U95, R1171_U96, R1171_U97, R1171_U98, R1171_U99, R1192_U10, R1192_U100, R1192_U101, R1192_U102, R1192_U103, R1192_U104, R1192_U105, R1192_U106, R1192_U107, R1192_U108, R1192_U109, R1192_U11, R1192_U110, R1192_U111, R1192_U112, R1192_U113, R1192_U114, R1192_U115, R1192_U116, R1192_U117, R1192_U118, R1192_U119, R1192_U12, R1192_U120, R1192_U121, R1192_U122, R1192_U123, R1192_U124, R1192_U125, R1192_U126, R1192_U127, R1192_U128, R1192_U129, R1192_U13, R1192_U130, R1192_U131, R1192_U132, R1192_U133, R1192_U134, R1192_U135, R1192_U136, R1192_U137, R1192_U138, R1192_U139, R1192_U14, R1192_U140, R1192_U141, R1192_U142, R1192_U143, R1192_U144, R1192_U145, R1192_U146, R1192_U147, R1192_U148, R1192_U149, R1192_U15, R1192_U150, R1192_U151, R1192_U152, R1192_U153, R1192_U154, R1192_U155, R1192_U156, R1192_U157, R1192_U158, R1192_U159, R1192_U16, R1192_U160, R1192_U161, R1192_U162, R1192_U163, R1192_U164, R1192_U165, R1192_U166, R1192_U167, R1192_U168, R1192_U169, R1192_U17, R1192_U170, R1192_U171, R1192_U172, R1192_U173, R1192_U174, R1192_U175, R1192_U176, R1192_U177, R1192_U178, R1192_U179, R1192_U18, R1192_U180, R1192_U181, R1192_U182, R1192_U183, R1192_U184, R1192_U185, R1192_U186, R1192_U187, R1192_U188, R1192_U189, R1192_U19, R1192_U190, R1192_U191, R1192_U192, R1192_U193, R1192_U194, R1192_U195, R1192_U196, R1192_U197, R1192_U198, R1192_U199, R1192_U20, R1192_U200, R1192_U201, R1192_U202, R1192_U203, R1192_U204, R1192_U205, R1192_U206, R1192_U207, R1192_U208, R1192_U209, R1192_U21, R1192_U210, R1192_U211, R1192_U212, R1192_U213, R1192_U214, R1192_U215, R1192_U216, R1192_U217, R1192_U218, R1192_U219, R1192_U22, R1192_U220, R1192_U221, R1192_U222, R1192_U223, R1192_U224, R1192_U225, R1192_U226, R1192_U227, R1192_U228, R1192_U229, R1192_U23, R1192_U230, R1192_U231, R1192_U232, R1192_U233, R1192_U234, R1192_U235, R1192_U236, R1192_U237, R1192_U238, R1192_U239, R1192_U24, R1192_U240, R1192_U241, R1192_U242, R1192_U243, R1192_U244, R1192_U245, R1192_U246, R1192_U247, R1192_U248, R1192_U249, R1192_U25, R1192_U250, R1192_U251, R1192_U252, R1192_U253, R1192_U254, R1192_U255, R1192_U256, R1192_U257, R1192_U258, R1192_U259, R1192_U26, R1192_U260, R1192_U261, R1192_U262, R1192_U263, R1192_U264, R1192_U265, R1192_U266, R1192_U267, R1192_U268, R1192_U269, R1192_U27, R1192_U270, R1192_U271, R1192_U272, R1192_U273, R1192_U274, R1192_U275, R1192_U276, R1192_U277, R1192_U278, R1192_U279, R1192_U28, R1192_U280, R1192_U281, R1192_U282, R1192_U283, R1192_U284, R1192_U285, R1192_U286, R1192_U287, R1192_U288, R1192_U289, R1192_U29, R1192_U290, R1192_U291, R1192_U292, R1192_U293, R1192_U294, R1192_U295, R1192_U296, R1192_U297, R1192_U298, R1192_U299, R1192_U30, R1192_U300, R1192_U301, R1192_U302, R1192_U303, R1192_U304, R1192_U305, R1192_U306, R1192_U307, R1192_U308, R1192_U309, R1192_U31, R1192_U310, R1192_U311, R1192_U312, R1192_U313, R1192_U314, R1192_U315, R1192_U316, R1192_U317, R1192_U318, R1192_U319, R1192_U32, R1192_U320, R1192_U321, R1192_U322, R1192_U323, R1192_U324, R1192_U325, R1192_U326, R1192_U327, R1192_U328, R1192_U329, R1192_U33, R1192_U330, R1192_U331, R1192_U332, R1192_U333, R1192_U334, R1192_U335, R1192_U336, R1192_U337, R1192_U338, R1192_U339, R1192_U34, R1192_U340, R1192_U341, R1192_U342, R1192_U343, R1192_U344, R1192_U345, R1192_U346, R1192_U347, R1192_U348, R1192_U349, R1192_U35, R1192_U350, R1192_U351, R1192_U352, R1192_U353, R1192_U354, R1192_U355, R1192_U356, R1192_U357, R1192_U358, R1192_U359, R1192_U36, R1192_U360, R1192_U361, R1192_U362, R1192_U363, R1192_U364, R1192_U365, R1192_U366, R1192_U367, R1192_U368, R1192_U369, R1192_U37, R1192_U370, R1192_U371, R1192_U372, R1192_U373, R1192_U374, R1192_U375, R1192_U376, R1192_U377, R1192_U378, R1192_U379, R1192_U38, R1192_U380, R1192_U381, R1192_U382, R1192_U383, R1192_U384, R1192_U385, R1192_U386, R1192_U387, R1192_U388, R1192_U389, R1192_U39, R1192_U390, R1192_U391, R1192_U392, R1192_U393, R1192_U394, R1192_U395, R1192_U396, R1192_U397, R1192_U398, R1192_U399, R1192_U40, R1192_U400, R1192_U401, R1192_U402, R1192_U403, R1192_U404, R1192_U405, R1192_U406, R1192_U407, R1192_U408, R1192_U409, R1192_U41, R1192_U410, R1192_U411, R1192_U412, R1192_U413, R1192_U414, R1192_U415, R1192_U416, R1192_U417, R1192_U418, R1192_U419, R1192_U42, R1192_U420, R1192_U421, R1192_U422, R1192_U423, R1192_U424, R1192_U425, R1192_U426, R1192_U427, R1192_U428, R1192_U429, R1192_U43, R1192_U430, R1192_U431, R1192_U432, R1192_U433, R1192_U434, R1192_U435, R1192_U436, R1192_U437, R1192_U438, R1192_U439, R1192_U44, R1192_U440, R1192_U441, R1192_U442, R1192_U443, R1192_U444, R1192_U445, R1192_U446, R1192_U447, R1192_U448, R1192_U449, R1192_U45, R1192_U450, R1192_U451, R1192_U452, R1192_U453, R1192_U454, R1192_U455, R1192_U456, R1192_U457, R1192_U458, R1192_U459, R1192_U46, R1192_U460, R1192_U461, R1192_U462, R1192_U463, R1192_U464, R1192_U465, R1192_U466, R1192_U467, R1192_U468, R1192_U469, R1192_U47, R1192_U470, R1192_U471, R1192_U472, R1192_U473, R1192_U474, R1192_U475, R1192_U476, R1192_U477, R1192_U478, R1192_U479, R1192_U48, R1192_U480, R1192_U481, R1192_U482, R1192_U483, R1192_U484, R1192_U485, R1192_U486, R1192_U487, R1192_U488, R1192_U489, R1192_U49, R1192_U490, R1192_U491, R1192_U492, R1192_U493, R1192_U494, R1192_U495, R1192_U496, R1192_U497, R1192_U498, R1192_U499, R1192_U50, R1192_U500, R1192_U501, R1192_U502, R1192_U503, R1192_U504, R1192_U505, R1192_U506, R1192_U507, R1192_U508, R1192_U509, R1192_U51, R1192_U510, R1192_U511, R1192_U512, R1192_U513, R1192_U514, R1192_U515, R1192_U516, R1192_U517, R1192_U518, R1192_U519, R1192_U52, R1192_U520, R1192_U53, R1192_U54, R1192_U55, R1192_U56, R1192_U57, R1192_U58, R1192_U59, R1192_U6, R1192_U60, R1192_U61, R1192_U62, R1192_U63, R1192_U64, R1192_U65, R1192_U66, R1192_U67, R1192_U68, R1192_U69, R1192_U7, R1192_U70, R1192_U71, R1192_U72, R1192_U73, R1192_U74, R1192_U75, R1192_U76, R1192_U77, R1192_U78, R1192_U79, R1192_U8, R1192_U80, R1192_U81, R1192_U82, R1192_U83, R1192_U84, R1192_U85, R1192_U86, R1192_U87, R1192_U88, R1192_U89, R1192_U9, R1192_U90, R1192_U91, R1192_U92, R1192_U93, R1192_U94, R1192_U95, R1192_U96, R1192_U97, R1192_U98, R1192_U99, R1207_U10, R1207_U100, R1207_U101, R1207_U102, R1207_U103, R1207_U104, R1207_U105, R1207_U106, R1207_U107, R1207_U108, R1207_U109, R1207_U11, R1207_U110, R1207_U111, R1207_U112, R1207_U113, R1207_U114, R1207_U115, R1207_U116, R1207_U117, R1207_U118, R1207_U119, R1207_U12, R1207_U120, R1207_U121, R1207_U122, R1207_U123, R1207_U124, R1207_U125, R1207_U126, R1207_U127, R1207_U128, R1207_U129, R1207_U13, R1207_U130, R1207_U131, R1207_U132, R1207_U133, R1207_U134, R1207_U135, R1207_U136, R1207_U137, R1207_U138, R1207_U139, R1207_U14, R1207_U140, R1207_U141, R1207_U142, R1207_U143, R1207_U144, R1207_U145, R1207_U146, R1207_U147, R1207_U148, R1207_U149, R1207_U15, R1207_U150, R1207_U151, R1207_U152, R1207_U153, R1207_U154, R1207_U155, R1207_U156, R1207_U157, R1207_U158, R1207_U159, R1207_U16, R1207_U160, R1207_U161, R1207_U162, R1207_U163, R1207_U164, R1207_U165, R1207_U166, R1207_U167, R1207_U168, R1207_U169, R1207_U17, R1207_U170, R1207_U171, R1207_U172, R1207_U173, R1207_U174, R1207_U175, R1207_U176, R1207_U177, R1207_U178, R1207_U179, R1207_U18, R1207_U180, R1207_U181, R1207_U182, R1207_U183, R1207_U184, R1207_U185, R1207_U186, R1207_U187, R1207_U188, R1207_U189, R1207_U19, R1207_U190, R1207_U191, R1207_U192, R1207_U193, R1207_U194, R1207_U195, R1207_U196, R1207_U197, R1207_U198, R1207_U199, R1207_U20, R1207_U200, R1207_U201, R1207_U202, R1207_U203, R1207_U204, R1207_U205, R1207_U206, R1207_U207, R1207_U208, R1207_U209, R1207_U21, R1207_U210, R1207_U211, R1207_U212, R1207_U213, R1207_U214, R1207_U215, R1207_U216, R1207_U217, R1207_U218, R1207_U219, R1207_U22, R1207_U220, R1207_U221, R1207_U222, R1207_U223, R1207_U224, R1207_U225, R1207_U226, R1207_U227, R1207_U228, R1207_U229, R1207_U23, R1207_U230, R1207_U231, R1207_U232, R1207_U233, R1207_U234, R1207_U235, R1207_U236, R1207_U237, R1207_U238, R1207_U239, R1207_U24, R1207_U240, R1207_U241, R1207_U242, R1207_U243, R1207_U244, R1207_U245, R1207_U246, R1207_U247, R1207_U248, R1207_U249, R1207_U25, R1207_U250, R1207_U251, R1207_U252, R1207_U253, R1207_U254, R1207_U255, R1207_U256, R1207_U257, R1207_U258, R1207_U259, R1207_U26, R1207_U260, R1207_U261, R1207_U262, R1207_U263, R1207_U264, R1207_U265, R1207_U266, R1207_U267, R1207_U268, R1207_U269, R1207_U27, R1207_U270, R1207_U271, R1207_U272, R1207_U273, R1207_U274, R1207_U275, R1207_U276, R1207_U277, R1207_U278, R1207_U279, R1207_U28, R1207_U280, R1207_U281, R1207_U282, R1207_U283, R1207_U284, R1207_U285, R1207_U286, R1207_U287, R1207_U288, R1207_U289, R1207_U29, R1207_U290, R1207_U291, R1207_U292, R1207_U293, R1207_U294, R1207_U295, R1207_U296, R1207_U297, R1207_U298, R1207_U299, R1207_U30, R1207_U300, R1207_U301, R1207_U302, R1207_U303, R1207_U304, R1207_U305, R1207_U306, R1207_U307, R1207_U308, R1207_U309, R1207_U31, R1207_U310, R1207_U311, R1207_U312, R1207_U313, R1207_U314, R1207_U315, R1207_U316, R1207_U317, R1207_U318, R1207_U319, R1207_U32, R1207_U320, R1207_U321, R1207_U322, R1207_U323, R1207_U324, R1207_U325, R1207_U326, R1207_U327, R1207_U328, R1207_U329, R1207_U33, R1207_U330, R1207_U331, R1207_U332, R1207_U333, R1207_U334, R1207_U335, R1207_U336, R1207_U337, R1207_U338, R1207_U339, R1207_U34, R1207_U340, R1207_U341, R1207_U342, R1207_U343, R1207_U344, R1207_U345, R1207_U346, R1207_U347, R1207_U348, R1207_U349, R1207_U35, R1207_U350, R1207_U351, R1207_U352, R1207_U353, R1207_U354, R1207_U355, R1207_U356, R1207_U357, R1207_U358, R1207_U359, R1207_U36, R1207_U360, R1207_U361, R1207_U362, R1207_U363, R1207_U364, R1207_U365, R1207_U366, R1207_U367, R1207_U368, R1207_U369, R1207_U37, R1207_U370, R1207_U371, R1207_U372, R1207_U373, R1207_U374, R1207_U375, R1207_U376, R1207_U377, R1207_U378, R1207_U379, R1207_U38, R1207_U380, R1207_U381, R1207_U382, R1207_U383, R1207_U384, R1207_U385, R1207_U386, R1207_U387, R1207_U388, R1207_U389, R1207_U39, R1207_U390, R1207_U391, R1207_U392, R1207_U393, R1207_U394, R1207_U395, R1207_U396, R1207_U397, R1207_U398, R1207_U399, R1207_U40, R1207_U400, R1207_U401, R1207_U402, R1207_U403, R1207_U404, R1207_U405, R1207_U406, R1207_U407, R1207_U408, R1207_U409, R1207_U41, R1207_U410, R1207_U411, R1207_U412, R1207_U413, R1207_U414, R1207_U415, R1207_U416, R1207_U417, R1207_U418, R1207_U419, R1207_U42, R1207_U420, R1207_U421, R1207_U422, R1207_U423, R1207_U424, R1207_U425, R1207_U426, R1207_U427, R1207_U428, R1207_U429, R1207_U43, R1207_U430, R1207_U431, R1207_U432, R1207_U433, R1207_U434, R1207_U435, R1207_U436, R1207_U437, R1207_U438, R1207_U439, R1207_U44, R1207_U440, R1207_U441, R1207_U442, R1207_U443, R1207_U444, R1207_U445, R1207_U446, R1207_U447, R1207_U448, R1207_U449, R1207_U45, R1207_U450, R1207_U451, R1207_U452, R1207_U453, R1207_U454, R1207_U455, R1207_U456, R1207_U457, R1207_U458, R1207_U459, R1207_U46, R1207_U460, R1207_U461, R1207_U462, R1207_U463, R1207_U464, R1207_U465, R1207_U466, R1207_U467, R1207_U468, R1207_U469, R1207_U47, R1207_U470, R1207_U471, R1207_U472, R1207_U473, R1207_U474, R1207_U475, R1207_U476, R1207_U477, R1207_U478, R1207_U479, R1207_U48, R1207_U480, R1207_U481, R1207_U482, R1207_U483, R1207_U484, R1207_U485, R1207_U486, R1207_U487, R1207_U488, R1207_U489, R1207_U49, R1207_U490, R1207_U491, R1207_U492, R1207_U493, R1207_U494, R1207_U495, R1207_U496, R1207_U497, R1207_U498, R1207_U499, R1207_U50, R1207_U500, R1207_U501, R1207_U502, R1207_U503, R1207_U504, R1207_U505, R1207_U506, R1207_U507, R1207_U508, R1207_U509, R1207_U51, R1207_U510, R1207_U511, R1207_U512, R1207_U513, R1207_U514, R1207_U515, R1207_U516, R1207_U517, R1207_U518, R1207_U519, R1207_U52, R1207_U520, R1207_U53, R1207_U54, R1207_U55, R1207_U56, R1207_U57, R1207_U58, R1207_U59, R1207_U6, R1207_U60, R1207_U61, R1207_U62, R1207_U63, R1207_U64, R1207_U65, R1207_U66, R1207_U67, R1207_U68, R1207_U69, R1207_U7, R1207_U70, R1207_U71, R1207_U72, R1207_U73, R1207_U74, R1207_U75, R1207_U76, R1207_U77, R1207_U78, R1207_U79, R1207_U8, R1207_U80, R1207_U81, R1207_U82, R1207_U83, R1207_U84, R1207_U85, R1207_U86, R1207_U87, R1207_U88, R1207_U89, R1207_U9, R1207_U90, R1207_U91, R1207_U92, R1207_U93, R1207_U94, R1207_U95, R1207_U96, R1207_U97, R1207_U98, R1207_U99, R1222_U10, R1222_U100, R1222_U101, R1222_U102, R1222_U103, R1222_U104, R1222_U105, R1222_U106, R1222_U107, R1222_U108, R1222_U109, R1222_U11, R1222_U110, R1222_U111, R1222_U112, R1222_U113, R1222_U114, R1222_U115, R1222_U116, R1222_U117, R1222_U118, R1222_U119, R1222_U12, R1222_U120, R1222_U121, R1222_U122, R1222_U123, R1222_U124, R1222_U125, R1222_U126, R1222_U127, R1222_U128, R1222_U129, R1222_U13, R1222_U130, R1222_U131, R1222_U132, R1222_U133, R1222_U134, R1222_U135, R1222_U136, R1222_U137, R1222_U138, R1222_U139, R1222_U14, R1222_U140, R1222_U141, R1222_U142, R1222_U143, R1222_U144, R1222_U145, R1222_U146, R1222_U147, R1222_U148, R1222_U149, R1222_U15, R1222_U150, R1222_U151, R1222_U152, R1222_U153, R1222_U154, R1222_U155, R1222_U156, R1222_U157, R1222_U158, R1222_U159, R1222_U16, R1222_U160, R1222_U161, R1222_U162, R1222_U163, R1222_U164, R1222_U165, R1222_U166, R1222_U167, R1222_U168, R1222_U169, R1222_U17, R1222_U170, R1222_U171, R1222_U172, R1222_U173, R1222_U174, R1222_U175, R1222_U176, R1222_U177, R1222_U178, R1222_U179, R1222_U18, R1222_U180, R1222_U181, R1222_U182, R1222_U183, R1222_U184, R1222_U185, R1222_U186, R1222_U187, R1222_U188, R1222_U189, R1222_U19, R1222_U190, R1222_U191, R1222_U192, R1222_U193, R1222_U194, R1222_U195, R1222_U196, R1222_U197, R1222_U198, R1222_U199, R1222_U20, R1222_U200, R1222_U201, R1222_U202, R1222_U203, R1222_U204, R1222_U205, R1222_U206, R1222_U207, R1222_U208, R1222_U209, R1222_U21, R1222_U210, R1222_U211, R1222_U212, R1222_U213, R1222_U214, R1222_U215, R1222_U216, R1222_U217, R1222_U218, R1222_U219, R1222_U22, R1222_U220, R1222_U221, R1222_U222, R1222_U223, R1222_U224, R1222_U225, R1222_U226, R1222_U227, R1222_U228, R1222_U229, R1222_U23, R1222_U230, R1222_U231, R1222_U232, R1222_U233, R1222_U234, R1222_U235, R1222_U236, R1222_U237, R1222_U238, R1222_U239, R1222_U24, R1222_U240, R1222_U241, R1222_U242, R1222_U243, R1222_U244, R1222_U245, R1222_U246, R1222_U247, R1222_U248, R1222_U249, R1222_U25, R1222_U250, R1222_U251, R1222_U252, R1222_U253, R1222_U254, R1222_U255, R1222_U256, R1222_U257, R1222_U258, R1222_U259, R1222_U26, R1222_U260, R1222_U261, R1222_U262, R1222_U263, R1222_U264, R1222_U265, R1222_U266, R1222_U267, R1222_U268, R1222_U269, R1222_U27, R1222_U270, R1222_U271, R1222_U272, R1222_U273, R1222_U274, R1222_U275, R1222_U276, R1222_U277, R1222_U278, R1222_U279, R1222_U28, R1222_U280, R1222_U281, R1222_U282, R1222_U283, R1222_U284, R1222_U285, R1222_U286, R1222_U287, R1222_U288, R1222_U289, R1222_U29, R1222_U290, R1222_U291, R1222_U292, R1222_U293, R1222_U294, R1222_U295, R1222_U296, R1222_U297, R1222_U298, R1222_U299, R1222_U30, R1222_U300, R1222_U301, R1222_U302, R1222_U303, R1222_U304, R1222_U305, R1222_U306, R1222_U307, R1222_U308, R1222_U309, R1222_U31, R1222_U310, R1222_U311, R1222_U312, R1222_U313, R1222_U314, R1222_U315, R1222_U316, R1222_U317, R1222_U318, R1222_U319, R1222_U32, R1222_U320, R1222_U321, R1222_U322, R1222_U323, R1222_U324, R1222_U325, R1222_U326, R1222_U327, R1222_U328, R1222_U329, R1222_U33, R1222_U330, R1222_U331, R1222_U332, R1222_U333, R1222_U334, R1222_U335, R1222_U336, R1222_U337, R1222_U338, R1222_U339, R1222_U34, R1222_U340, R1222_U341, R1222_U342, R1222_U343, R1222_U344, R1222_U345, R1222_U346, R1222_U347, R1222_U348, R1222_U349, R1222_U35, R1222_U350, R1222_U351, R1222_U352, R1222_U353, R1222_U354, R1222_U355, R1222_U356, R1222_U357, R1222_U358, R1222_U359, R1222_U36, R1222_U360, R1222_U361, R1222_U362, R1222_U363, R1222_U364, R1222_U365, R1222_U366, R1222_U367, R1222_U368, R1222_U369, R1222_U37, R1222_U370, R1222_U371, R1222_U372, R1222_U373, R1222_U374, R1222_U375, R1222_U376, R1222_U377, R1222_U378, R1222_U379, R1222_U38, R1222_U380, R1222_U381, R1222_U382, R1222_U383, R1222_U384, R1222_U385, R1222_U386, R1222_U387, R1222_U388, R1222_U389, R1222_U39, R1222_U390, R1222_U391, R1222_U392, R1222_U393, R1222_U394, R1222_U395, R1222_U396, R1222_U397, R1222_U398, R1222_U399, R1222_U4, R1222_U40, R1222_U400, R1222_U401, R1222_U402, R1222_U403, R1222_U404, R1222_U405, R1222_U406, R1222_U407, R1222_U408, R1222_U409, R1222_U41, R1222_U410, R1222_U411, R1222_U412, R1222_U413, R1222_U414, R1222_U415, R1222_U416, R1222_U417, R1222_U418, R1222_U419, R1222_U42, R1222_U420, R1222_U421, R1222_U422, R1222_U423, R1222_U424, R1222_U425, R1222_U426, R1222_U427, R1222_U428, R1222_U429, R1222_U43, R1222_U430, R1222_U431, R1222_U432, R1222_U433, R1222_U434, R1222_U435, R1222_U436, R1222_U437, R1222_U438, R1222_U439, R1222_U44, R1222_U440, R1222_U441, R1222_U442, R1222_U443, R1222_U444, R1222_U445, R1222_U446, R1222_U447, R1222_U448, R1222_U449, R1222_U45, R1222_U450, R1222_U451, R1222_U452, R1222_U453, R1222_U454, R1222_U455, R1222_U456, R1222_U457, R1222_U458, R1222_U459, R1222_U46, R1222_U460, R1222_U461, R1222_U462, R1222_U463, R1222_U464, R1222_U465, R1222_U466, R1222_U467, R1222_U468, R1222_U469, R1222_U47, R1222_U470, R1222_U471, R1222_U472, R1222_U473, R1222_U474, R1222_U475, R1222_U476, R1222_U477, R1222_U478, R1222_U479, R1222_U48, R1222_U480, R1222_U481, R1222_U482, R1222_U483, R1222_U484, R1222_U485, R1222_U486, R1222_U487, R1222_U488, R1222_U489, R1222_U49, R1222_U490, R1222_U491, R1222_U492, R1222_U493, R1222_U494, R1222_U495, R1222_U496, R1222_U497, R1222_U498, R1222_U499, R1222_U5, R1222_U50, R1222_U500, R1222_U501, R1222_U502, R1222_U503, R1222_U504, R1222_U505, R1222_U506, R1222_U507, R1222_U508, R1222_U509, R1222_U51, R1222_U510, R1222_U511, R1222_U512, R1222_U513, R1222_U514, R1222_U515, R1222_U516, R1222_U517, R1222_U518, R1222_U519, R1222_U52, R1222_U53, R1222_U54, R1222_U55, R1222_U56, R1222_U57, R1222_U58, R1222_U59, R1222_U6, R1222_U60, R1222_U61, R1222_U62, R1222_U63, R1222_U64, R1222_U65, R1222_U66, R1222_U67, R1222_U68, R1222_U69, R1222_U7, R1222_U70, R1222_U71, R1222_U72, R1222_U73, R1222_U74, R1222_U75, R1222_U76, R1222_U77, R1222_U78, R1222_U79, R1222_U8, R1222_U80, R1222_U81, R1222_U82, R1222_U83, R1222_U84, R1222_U85, R1222_U86, R1222_U87, R1222_U88, R1222_U89, R1222_U9, R1222_U90, R1222_U91, R1222_U92, R1222_U93, R1222_U94, R1222_U95, R1222_U96, R1222_U97, R1222_U98, R1222_U99, R1240_U10, R1240_U100, R1240_U101, R1240_U102, R1240_U103, R1240_U104, R1240_U105, R1240_U106, R1240_U107, R1240_U108, R1240_U109, R1240_U11, R1240_U110, R1240_U111, R1240_U112, R1240_U113, R1240_U114, R1240_U115, R1240_U116, R1240_U117, R1240_U118, R1240_U119, R1240_U12, R1240_U120, R1240_U121, R1240_U122, R1240_U123, R1240_U124, R1240_U125, R1240_U126, R1240_U127, R1240_U128, R1240_U129, R1240_U13, R1240_U130, R1240_U131, R1240_U132, R1240_U133, R1240_U134, R1240_U135, R1240_U136, R1240_U137, R1240_U138, R1240_U139, R1240_U14, R1240_U140, R1240_U141, R1240_U142, R1240_U143, R1240_U144, R1240_U145, R1240_U146, R1240_U147, R1240_U148, R1240_U149, R1240_U15, R1240_U150, R1240_U151, R1240_U152, R1240_U153, R1240_U154, R1240_U155, R1240_U156, R1240_U157, R1240_U158, R1240_U159, R1240_U16, R1240_U160, R1240_U161, R1240_U162, R1240_U163, R1240_U164, R1240_U165, R1240_U166, R1240_U167, R1240_U168, R1240_U169, R1240_U17, R1240_U170, R1240_U171, R1240_U172, R1240_U173, R1240_U174, R1240_U175, R1240_U176, R1240_U177, R1240_U178, R1240_U179, R1240_U18, R1240_U180, R1240_U181, R1240_U182, R1240_U183, R1240_U184, R1240_U185, R1240_U186, R1240_U187, R1240_U188, R1240_U189, R1240_U19, R1240_U190, R1240_U191, R1240_U192, R1240_U193, R1240_U194, R1240_U195, R1240_U196, R1240_U197, R1240_U198, R1240_U199, R1240_U20, R1240_U200, R1240_U201, R1240_U202, R1240_U203, R1240_U204, R1240_U205, R1240_U206, R1240_U207, R1240_U208, R1240_U209, R1240_U21, R1240_U210, R1240_U211, R1240_U212, R1240_U213, R1240_U214, R1240_U215, R1240_U216, R1240_U217, R1240_U218, R1240_U219, R1240_U22, R1240_U220, R1240_U221, R1240_U222, R1240_U223, R1240_U224, R1240_U225, R1240_U226, R1240_U227, R1240_U228, R1240_U229, R1240_U23, R1240_U230, R1240_U231, R1240_U232, R1240_U233, R1240_U234, R1240_U235, R1240_U236, R1240_U237, R1240_U238, R1240_U239, R1240_U24, R1240_U240, R1240_U241, R1240_U242, R1240_U243, R1240_U244, R1240_U245, R1240_U246, R1240_U247, R1240_U248, R1240_U249, R1240_U25, R1240_U250, R1240_U251, R1240_U252, R1240_U253, R1240_U254, R1240_U255, R1240_U256, R1240_U257, R1240_U258, R1240_U259, R1240_U26, R1240_U260, R1240_U261, R1240_U262, R1240_U263, R1240_U264, R1240_U265, R1240_U266, R1240_U267, R1240_U268, R1240_U269, R1240_U27, R1240_U270, R1240_U271, R1240_U272, R1240_U273, R1240_U274, R1240_U275, R1240_U276, R1240_U277, R1240_U278, R1240_U279, R1240_U28, R1240_U280, R1240_U281, R1240_U282, R1240_U283, R1240_U284, R1240_U285, R1240_U286, R1240_U287, R1240_U288, R1240_U289, R1240_U29, R1240_U290, R1240_U291, R1240_U292, R1240_U293, R1240_U294, R1240_U295, R1240_U296, R1240_U297, R1240_U298, R1240_U299, R1240_U30, R1240_U300, R1240_U301, R1240_U302, R1240_U303, R1240_U304, R1240_U305, R1240_U306, R1240_U307, R1240_U308, R1240_U309, R1240_U31, R1240_U310, R1240_U311, R1240_U312, R1240_U313, R1240_U314, R1240_U315, R1240_U316, R1240_U317, R1240_U318, R1240_U319, R1240_U32, R1240_U320, R1240_U321, R1240_U322, R1240_U323, R1240_U324, R1240_U325, R1240_U326, R1240_U327, R1240_U328, R1240_U329, R1240_U33, R1240_U330, R1240_U331, R1240_U332, R1240_U333, R1240_U334, R1240_U335, R1240_U336, R1240_U337, R1240_U338, R1240_U339, R1240_U34, R1240_U340, R1240_U341, R1240_U342, R1240_U343, R1240_U344, R1240_U345, R1240_U346, R1240_U347, R1240_U348, R1240_U349, R1240_U35, R1240_U350, R1240_U351, R1240_U352, R1240_U353, R1240_U354, R1240_U355, R1240_U356, R1240_U357, R1240_U358, R1240_U359, R1240_U36, R1240_U360, R1240_U361, R1240_U362, R1240_U363, R1240_U364, R1240_U365, R1240_U366, R1240_U367, R1240_U368, R1240_U369, R1240_U37, R1240_U370, R1240_U371, R1240_U372, R1240_U373, R1240_U374, R1240_U375, R1240_U376, R1240_U377, R1240_U378, R1240_U379, R1240_U38, R1240_U380, R1240_U381, R1240_U382, R1240_U383, R1240_U384, R1240_U385, R1240_U386, R1240_U387, R1240_U388, R1240_U389, R1240_U39, R1240_U390, R1240_U391, R1240_U392, R1240_U393, R1240_U394, R1240_U395, R1240_U396, R1240_U397, R1240_U398, R1240_U399, R1240_U4, R1240_U40, R1240_U400, R1240_U401, R1240_U402, R1240_U403, R1240_U404, R1240_U405, R1240_U406, R1240_U407, R1240_U408, R1240_U409, R1240_U41, R1240_U410, R1240_U411, R1240_U412, R1240_U413, R1240_U414, R1240_U415, R1240_U416, R1240_U417, R1240_U418, R1240_U419, R1240_U42, R1240_U420, R1240_U421, R1240_U422, R1240_U423, R1240_U424, R1240_U425, R1240_U426, R1240_U427, R1240_U428, R1240_U429, R1240_U43, R1240_U430, R1240_U431, R1240_U432, R1240_U433, R1240_U434, R1240_U435, R1240_U436, R1240_U437, R1240_U438, R1240_U439, R1240_U44, R1240_U440, R1240_U441, R1240_U442, R1240_U443, R1240_U444, R1240_U445, R1240_U446, R1240_U447, R1240_U448, R1240_U449, R1240_U45, R1240_U450, R1240_U451, R1240_U452, R1240_U453, R1240_U454, R1240_U455, R1240_U456, R1240_U457, R1240_U458, R1240_U459, R1240_U46, R1240_U460, R1240_U461, R1240_U462, R1240_U463, R1240_U464, R1240_U465, R1240_U466, R1240_U467, R1240_U468, R1240_U469, R1240_U47, R1240_U470, R1240_U471, R1240_U472, R1240_U473, R1240_U474, R1240_U475, R1240_U476, R1240_U477, R1240_U478, R1240_U479, R1240_U48, R1240_U480, R1240_U481, R1240_U482, R1240_U483, R1240_U484, R1240_U485, R1240_U486, R1240_U487, R1240_U488, R1240_U489, R1240_U49, R1240_U490, R1240_U491, R1240_U492, R1240_U493, R1240_U494, R1240_U495, R1240_U496, R1240_U497, R1240_U498, R1240_U499, R1240_U5, R1240_U50, R1240_U500, R1240_U501, R1240_U502, R1240_U503, R1240_U504, R1240_U505, R1240_U506, R1240_U507, R1240_U508, R1240_U509, R1240_U51, R1240_U510, R1240_U511, R1240_U512, R1240_U513, R1240_U514, R1240_U515, R1240_U516, R1240_U517, R1240_U518, R1240_U519, R1240_U52, R1240_U520, R1240_U521, R1240_U522, R1240_U523, R1240_U524, R1240_U525, R1240_U526, R1240_U527, R1240_U528, R1240_U529, R1240_U53, R1240_U530, R1240_U531, R1240_U54, R1240_U55, R1240_U56, R1240_U57, R1240_U58, R1240_U59, R1240_U6, R1240_U60, R1240_U61, R1240_U62, R1240_U63, R1240_U64, R1240_U65, R1240_U66, R1240_U67, R1240_U68, R1240_U69, R1240_U7, R1240_U70, R1240_U71, R1240_U72, R1240_U73, R1240_U74, R1240_U75, R1240_U76, R1240_U77, R1240_U78, R1240_U79, R1240_U8, R1240_U80, R1240_U81, R1240_U82, R1240_U83, R1240_U84, R1240_U85, R1240_U86, R1240_U87, R1240_U88, R1240_U89, R1240_U9, R1240_U90, R1240_U91, R1240_U92, R1240_U93, R1240_U94, R1240_U95, R1240_U96, R1240_U97, R1240_U98, R1240_U99, R1282_U10, R1282_U100, R1282_U101, R1282_U102, R1282_U103, R1282_U104, R1282_U105, R1282_U106, R1282_U107, R1282_U108, R1282_U109, R1282_U11, R1282_U110, R1282_U111, R1282_U112, R1282_U113, R1282_U114, R1282_U115, R1282_U116, R1282_U117, R1282_U118, R1282_U119, R1282_U12, R1282_U120, R1282_U121, R1282_U122, R1282_U123, R1282_U124, R1282_U125, R1282_U126, R1282_U127, R1282_U128, R1282_U129, R1282_U13, R1282_U130, R1282_U131, R1282_U132, R1282_U133, R1282_U134, R1282_U135, R1282_U136, R1282_U137, R1282_U138, R1282_U139, R1282_U14, R1282_U140, R1282_U141, R1282_U142, R1282_U143, R1282_U144, R1282_U145, R1282_U146, R1282_U147, R1282_U148, R1282_U149, R1282_U15, R1282_U150, R1282_U151, R1282_U152, R1282_U153, R1282_U154, R1282_U155, R1282_U156, R1282_U157, R1282_U158, R1282_U159, R1282_U16, R1282_U160, R1282_U161, R1282_U162, R1282_U163, R1282_U164, R1282_U165, R1282_U166, R1282_U167, R1282_U168, R1282_U169, R1282_U17, R1282_U170, R1282_U171, R1282_U172, R1282_U173, R1282_U174, R1282_U175, R1282_U176, R1282_U177, R1282_U178, R1282_U179, R1282_U18, R1282_U180, R1282_U19, R1282_U20, R1282_U21, R1282_U22, R1282_U23, R1282_U24, R1282_U25, R1282_U26, R1282_U27, R1282_U28, R1282_U29, R1282_U30, R1282_U31, R1282_U32, R1282_U33, R1282_U34, R1282_U35, R1282_U36, R1282_U37, R1282_U38, R1282_U39, R1282_U40, R1282_U41, R1282_U42, R1282_U43, R1282_U44, R1282_U45, R1282_U46, R1282_U47, R1282_U48, R1282_U49, R1282_U50, R1282_U51, R1282_U52, R1282_U53, R1282_U54, R1282_U55, R1282_U56, R1282_U57, R1282_U58, R1282_U59, R1282_U6, R1282_U60, R1282_U61, R1282_U62, R1282_U63, R1282_U64, R1282_U65, R1282_U66, R1282_U67, R1282_U68, R1282_U69, R1282_U7, R1282_U70, R1282_U71, R1282_U72, R1282_U73, R1282_U74, R1282_U75, R1282_U76, R1282_U77, R1282_U78, R1282_U79, R1282_U8, R1282_U80, R1282_U81, R1282_U82, R1282_U83, R1282_U84, R1282_U85, R1282_U86, R1282_U87, R1282_U88, R1282_U89, R1282_U9, R1282_U90, R1282_U91, R1282_U92, R1282_U93, R1282_U94, R1282_U95, R1282_U96, R1282_U97, R1282_U98, R1282_U99, R1309_U10, R1309_U6, R1309_U7, R1309_U8, R1309_U9, R1347_U10, R1347_U100, R1347_U101, R1347_U102, R1347_U103, R1347_U104, R1347_U105, R1347_U106, R1347_U107, R1347_U108, R1347_U109, R1347_U11, R1347_U110, R1347_U111, R1347_U112, R1347_U113, R1347_U114, R1347_U115, R1347_U116, R1347_U117, R1347_U118, R1347_U119, R1347_U12, R1347_U120, R1347_U121, R1347_U122, R1347_U123, R1347_U124, R1347_U125, R1347_U126, R1347_U127, R1347_U128, R1347_U129, R1347_U13, R1347_U130, R1347_U131, R1347_U132, R1347_U133, R1347_U134, R1347_U135, R1347_U136, R1347_U137, R1347_U138, R1347_U139, R1347_U14, R1347_U140, R1347_U141, R1347_U142, R1347_U143, R1347_U144, R1347_U145, R1347_U146, R1347_U147, R1347_U148, R1347_U149, R1347_U15, R1347_U150, R1347_U151, R1347_U152, R1347_U153, R1347_U154, R1347_U155, R1347_U156, R1347_U157, R1347_U158, R1347_U159, R1347_U16, R1347_U160, R1347_U161, R1347_U162, R1347_U163, R1347_U164, R1347_U165, R1347_U166, R1347_U167, R1347_U168, R1347_U169, R1347_U17, R1347_U170, R1347_U171, R1347_U172, R1347_U173, R1347_U174, R1347_U175, R1347_U176, R1347_U177, R1347_U178, R1347_U179, R1347_U18, R1347_U180, R1347_U181, R1347_U182, R1347_U183, R1347_U184, R1347_U185, R1347_U186, R1347_U187, R1347_U188, R1347_U189, R1347_U19, R1347_U190, R1347_U191, R1347_U192, R1347_U193, R1347_U194, R1347_U195, R1347_U196, R1347_U197, R1347_U198, R1347_U199, R1347_U20, R1347_U200, R1347_U201, R1347_U202, R1347_U203, R1347_U204, R1347_U205, R1347_U206, R1347_U207, R1347_U208, R1347_U209, R1347_U21, R1347_U210, R1347_U211, R1347_U212, R1347_U22, R1347_U23, R1347_U24, R1347_U25, R1347_U26, R1347_U27, R1347_U28, R1347_U29, R1347_U30, R1347_U31, R1347_U32, R1347_U33, R1347_U34, R1347_U35, R1347_U36, R1347_U37, R1347_U38, R1347_U39, R1347_U40, R1347_U41, R1347_U42, R1347_U43, R1347_U44, R1347_U45, R1347_U46, R1347_U47, R1347_U48, R1347_U49, R1347_U50, R1347_U51, R1347_U52, R1347_U53, R1347_U54, R1347_U55, R1347_U56, R1347_U57, R1347_U58, R1347_U59, R1347_U6, R1347_U60, R1347_U61, R1347_U62, R1347_U63, R1347_U64, R1347_U65, R1347_U66, R1347_U67, R1347_U68, R1347_U69, R1347_U7, R1347_U70, R1347_U71, R1347_U72, R1347_U73, R1347_U74, R1347_U75, R1347_U76, R1347_U77, R1347_U78, R1347_U79, R1347_U8, R1347_U80, R1347_U81, R1347_U82, R1347_U83, R1347_U84, R1347_U85, R1347_U86, R1347_U87, R1347_U88, R1347_U89, R1347_U9, R1347_U90, R1347_U91, R1347_U92, R1347_U93, R1347_U94, R1347_U95, R1347_U96, R1347_U97, R1347_U98, R1347_U99, R1352_U6, R1352_U7, R1375_U10, R1375_U100, R1375_U101, R1375_U102, R1375_U103, R1375_U104, R1375_U105, R1375_U106, R1375_U107, R1375_U108, R1375_U109, R1375_U11, R1375_U110, R1375_U111, R1375_U112, R1375_U113, R1375_U114, R1375_U115, R1375_U116, R1375_U117, R1375_U118, R1375_U119, R1375_U12, R1375_U120, R1375_U121, R1375_U122, R1375_U123, R1375_U124, R1375_U125, R1375_U126, R1375_U127, R1375_U128, R1375_U129, R1375_U13, R1375_U130, R1375_U131, R1375_U132, R1375_U133, R1375_U134, R1375_U135, R1375_U136, R1375_U137, R1375_U138, R1375_U139, R1375_U14, R1375_U140, R1375_U141, R1375_U142, R1375_U143, R1375_U144, R1375_U145, R1375_U146, R1375_U147, R1375_U148, R1375_U149, R1375_U15, R1375_U150, R1375_U151, R1375_U152, R1375_U153, R1375_U154, R1375_U155, R1375_U156, R1375_U157, R1375_U158, R1375_U159, R1375_U16, R1375_U160, R1375_U161, R1375_U162, R1375_U163, R1375_U164, R1375_U165, R1375_U166, R1375_U167, R1375_U168, R1375_U169, R1375_U17, R1375_U170, R1375_U171, R1375_U172, R1375_U173, R1375_U174, R1375_U175, R1375_U176, R1375_U177, R1375_U178, R1375_U179, R1375_U18, R1375_U180, R1375_U181, R1375_U182, R1375_U183, R1375_U184, R1375_U185, R1375_U186, R1375_U187, R1375_U188, R1375_U189, R1375_U19, R1375_U190, R1375_U191, R1375_U192, R1375_U193, R1375_U194, R1375_U195, R1375_U196, R1375_U197, R1375_U198, R1375_U199, R1375_U20, R1375_U200, R1375_U201, R1375_U202, R1375_U203, R1375_U204, R1375_U205, R1375_U206, R1375_U207, R1375_U208, R1375_U209, R1375_U21, R1375_U210, R1375_U211, R1375_U212, R1375_U213, R1375_U214, R1375_U215, R1375_U216, R1375_U217, R1375_U218, R1375_U219, R1375_U22, R1375_U220, R1375_U221, R1375_U222, R1375_U223, R1375_U224, R1375_U225, R1375_U23, R1375_U24, R1375_U25, R1375_U26, R1375_U27, R1375_U28, R1375_U29, R1375_U30, R1375_U31, R1375_U32, R1375_U33, R1375_U34, R1375_U35, R1375_U36, R1375_U37, R1375_U38, R1375_U39, R1375_U40, R1375_U41, R1375_U42, R1375_U43, R1375_U44, R1375_U45, R1375_U46, R1375_U47, R1375_U48, R1375_U49, R1375_U50, R1375_U51, R1375_U52, R1375_U53, R1375_U54, R1375_U55, R1375_U56, R1375_U57, R1375_U58, R1375_U59, R1375_U6, R1375_U60, R1375_U61, R1375_U62, R1375_U63, R1375_U64, R1375_U65, R1375_U66, R1375_U67, R1375_U68, R1375_U69, R1375_U7, R1375_U70, R1375_U71, R1375_U72, R1375_U73, R1375_U74, R1375_U75, R1375_U76, R1375_U77, R1375_U78, R1375_U79, R1375_U8, R1375_U80, R1375_U81, R1375_U82, R1375_U83, R1375_U84, R1375_U85, R1375_U86, R1375_U87, R1375_U88, R1375_U89, R1375_U9, R1375_U90, R1375_U91, R1375_U92, R1375_U93, R1375_U94, R1375_U95, R1375_U96, R1375_U97, R1375_U98, R1375_U99, R395_U10, R395_U100, R395_U101, R395_U102, R395_U103, R395_U104, R395_U105, R395_U106, R395_U107, R395_U108, R395_U109, R395_U11, R395_U110, R395_U111, R395_U112, R395_U113, R395_U114, R395_U115, R395_U116, R395_U117, R395_U118, R395_U119, R395_U12, R395_U120, R395_U121, R395_U122, R395_U123, R395_U124, R395_U125, R395_U126, R395_U127, R395_U128, R395_U129, R395_U13, R395_U130, R395_U131, R395_U132, R395_U133, R395_U134, R395_U135, R395_U136, R395_U137, R395_U138, R395_U139, R395_U14, R395_U140, R395_U141, R395_U142, R395_U143, R395_U144, R395_U145, R395_U146, R395_U147, R395_U148, R395_U149, R395_U15, R395_U150, R395_U151, R395_U152, R395_U153, R395_U154, R395_U155, R395_U156, R395_U157, R395_U158, R395_U159, R395_U16, R395_U160, R395_U161, R395_U162, R395_U163, R395_U164, R395_U165, R395_U166, R395_U167, R395_U168, R395_U169, R395_U17, R395_U170, R395_U171, R395_U172, R395_U173, R395_U174, R395_U175, R395_U176, R395_U177, R395_U178, R395_U179, R395_U18, R395_U180, R395_U181, R395_U182, R395_U183, R395_U184, R395_U185, R395_U186, R395_U187, R395_U188, R395_U19, R395_U20, R395_U21, R395_U22, R395_U23, R395_U24, R395_U25, R395_U26, R395_U27, R395_U28, R395_U29, R395_U30, R395_U31, R395_U32, R395_U33, R395_U34, R395_U35, R395_U36, R395_U37, R395_U38, R395_U39, R395_U40, R395_U41, R395_U42, R395_U43, R395_U44, R395_U45, R395_U46, R395_U47, R395_U48, R395_U49, R395_U50, R395_U51, R395_U52, R395_U53, R395_U54, R395_U55, R395_U56, R395_U57, R395_U58, R395_U59, R395_U6, R395_U60, R395_U61, R395_U62, R395_U63, R395_U64, R395_U65, R395_U66, R395_U67, R395_U68, R395_U69, R395_U7, R395_U70, R395_U71, R395_U72, R395_U73, R395_U74, R395_U75, R395_U76, R395_U77, R395_U78, R395_U79, R395_U8, R395_U80, R395_U81, R395_U82, R395_U83, R395_U84, R395_U85, R395_U86, R395_U87, R395_U88, R395_U89, R395_U9, R395_U90, R395_U91, R395_U92, R395_U93, R395_U94, R395_U95, R395_U96, R395_U97, R395_U98, R395_U99, SUB_84_U10, SUB_84_U100, SUB_84_U101, SUB_84_U102, SUB_84_U103, SUB_84_U104, SUB_84_U105, SUB_84_U106, SUB_84_U107, SUB_84_U108, SUB_84_U109, SUB_84_U11, SUB_84_U110, SUB_84_U111, SUB_84_U112, SUB_84_U113, SUB_84_U114, SUB_84_U115, SUB_84_U116, SUB_84_U117, SUB_84_U118, SUB_84_U119, SUB_84_U12, SUB_84_U120, SUB_84_U121, SUB_84_U122, SUB_84_U123, SUB_84_U124, SUB_84_U125, SUB_84_U126, SUB_84_U127, SUB_84_U128, SUB_84_U129, SUB_84_U13, SUB_84_U130, SUB_84_U131, SUB_84_U132, SUB_84_U133, SUB_84_U134, SUB_84_U135, SUB_84_U136, SUB_84_U137, SUB_84_U138, SUB_84_U139, SUB_84_U14, SUB_84_U140, SUB_84_U141, SUB_84_U142, SUB_84_U143, SUB_84_U144, SUB_84_U145, SUB_84_U146, SUB_84_U147, SUB_84_U148, SUB_84_U149, SUB_84_U15, SUB_84_U150, SUB_84_U151, SUB_84_U152, SUB_84_U153, SUB_84_U154, SUB_84_U155, SUB_84_U156, SUB_84_U157, SUB_84_U158, SUB_84_U159, SUB_84_U16, SUB_84_U160, SUB_84_U161, SUB_84_U17, SUB_84_U18, SUB_84_U19, SUB_84_U20, SUB_84_U21, SUB_84_U22, SUB_84_U23, SUB_84_U24, SUB_84_U25, SUB_84_U26, SUB_84_U27, SUB_84_U28, SUB_84_U29, SUB_84_U30, SUB_84_U31, SUB_84_U32, SUB_84_U33, SUB_84_U34, SUB_84_U35, SUB_84_U36, SUB_84_U37, SUB_84_U38, SUB_84_U39, SUB_84_U4, SUB_84_U40, SUB_84_U41, SUB_84_U42, SUB_84_U43, SUB_84_U44, SUB_84_U45, SUB_84_U46, SUB_84_U47, SUB_84_U48, SUB_84_U49, SUB_84_U5, SUB_84_U50, SUB_84_U51, SUB_84_U52, SUB_84_U53, SUB_84_U54, SUB_84_U55, SUB_84_U56, SUB_84_U57, SUB_84_U58, SUB_84_U59, SUB_84_U6, SUB_84_U60, SUB_84_U61, SUB_84_U62, SUB_84_U63, SUB_84_U64, SUB_84_U65, SUB_84_U66, SUB_84_U67, SUB_84_U68, SUB_84_U69, SUB_84_U7, SUB_84_U70, SUB_84_U71, SUB_84_U72, SUB_84_U73, SUB_84_U74, SUB_84_U75, SUB_84_U76, SUB_84_U77, SUB_84_U78, SUB_84_U79, SUB_84_U8, SUB_84_U80, SUB_84_U81, SUB_84_U82, SUB_84_U83, SUB_84_U84, SUB_84_U85, SUB_84_U86, SUB_84_U87, SUB_84_U88, SUB_84_U89, SUB_84_U9, SUB_84_U90, SUB_84_U91, SUB_84_U92, SUB_84_U93, SUB_84_U94, SUB_84_U95, SUB_84_U96, SUB_84_U97, SUB_84_U98, SUB_84_U99, U3014, U3015, U3016, U3017, U3018, U3019, U3020, U3021, U3022, U3023, U3024, U3025, U3026, U3027, U3028, U3029, U3030, U3031, U3032, U3033, U3034, U3035, U3036, U3037, U3038, U3039, U3040, U3041, U3042, U3043, U3044, U3045, U3046, U3047, U3048, U3049, U3050, U3051, U3052, U3053, U3054, U3055, U3056, U3057, U3058, U3059, U3060, U3061, U3062, U3063, U3064, U3065, U3066, U3067, U3068, U3069, U3070, U3071, U3072, U3073, U3074, U3075, U3076, U3077, U3078, U3079, U3080, U3081, U3082, U3083, U3084, U3085, U3086, U3087, U3088, U3089, U3090, U3091, U3092, U3093, U3094, U3095, U3096, U3097, U3098, U3099, U3100, U3101, U3102, U3103, U3104, U3105, U3106, U3107, U3108, U3109, U3110, U3111, U3112, U3113, U3114, U3115, U3116, U3117, U3118, U3119, U3120, U3121, U3122, U3123, U3124, U3125, U3126, U3127, U3128, U3129, U3130, U3131, U3132, U3133, U3134, U3135, U3136, U3137, U3138, U3139, U3140, U3141, U3142, U3143, U3144, U3145, U3146, U3147, U3150, U3151, U3152, U3153, U3154, U3155, U3156, U3157, U3158, U3159, U3160, U3161, U3162, U3163, U3164, U3165, U3166, U3167, U3168, U3169, U3170, U3171, U3172, U3173, U3174, U3175, U3176, U3177, U3178, U3179, U3180, U3181, U3182, U3183, U3184, U3185, U3186, U3187, U3188, U3189, U3190, U3191, U3192, U3193, U3194, U3195, U3196, U3197, U3198, U3199, U3200, U3201, U3202, U3203, U3204, U3205, U3206, U3207, U3208, U3209, U3353, U3355, U3356, U3357, U3358, U3359, U3360, U3361, U3362, U3363, U3364, U3365, U3366, U3367, U3368, U3369, U3370, U3371, U3372, U3373, U3374, U3375, U3376, U3377, U3378, U3379, U3380, U3381, U3382, U3383, U3384, U3385, U3386, U3387, U3388, U3389, U3390, U3391, U3392, U3393, U3394, U3395, U3396, U3397, U3398, U3399, U3400, U3401, U3402, U3403, U3404, U3405, U3406, U3407, U3408, U3409, U3410, U3411, U3412, U3413, U3414, U3415, U3416, U3417, U3418, U3419, U3420, U3421, U3422, U3423, U3424, U3425, U3426, U3427, U3428, U3429, U3430, U3431, U3432, U3433, U3434, U3435, U3436, U3437, U3438, U3439, U3440, U3441, U3442, U3443, U3444, U3445, U3446, U3447, U3448, U3449, U3450, U3451, U3452, U3453, U3454, U3455, U3456, U3457, U3460, U3461, U3462, U3463, U3464, U3465, U3466, U3468, U3470, U3472, U3474, U3476, U3478, U3480, U3482, U3484, U3486, U3488, U3490, U3492, U3494, U3496, U3498, U3500, U3502, U3504, U3582, U3583, U3584, U3585, U3586, U3587, U3588, U3589, U3590, U3591, U3592, U3593, U3594, U3595, U3596, U3597, U3598, U3599, U3600, U3601, U3602, U3603, U3604, U3605, U3606, U3607, U3608, U3609, U3610, U3611, U3612, U3613, U3614, U3615, U3616, U3617, U3618, U3619, U3620, U3621, U3622, U3623, U3624, U3625, U3626, U3627, U3628, U3629, U3630, U3631, U3632, U3633, U3634, U3635, U3636, U3637, U3638, U3639, U3640, U3641, U3642, U3643, U3644, U3645, U3646, U3647, U3648, U3649, U3650, U3651, U3652, U3653, U3654, U3655, U3656, U3657, U3658, U3659, U3660, U3661, U3662, U3663, U3664, U3665, U3666, U3667, U3668, U3669, U3670, U3671, U3672, U3673, U3674, U3675, U3676, U3677, U3678, U3679, U3680, U3681, U3682, U3683, U3684, U3685, U3686, U3687, U3688, U3689, U3690, U3691, U3692, U3693, U3694, U3695, U3696, U3697, U3698, U3699, U3700, U3701, U3702, U3703, U3704, U3705, U3706, U3707, U3708, U3709, U3710, U3711, U3712, U3713, U3714, U3715, U3716, U3717, U3718, U3719, U3720, U3721, U3722, U3723, U3724, U3725, U3726, U3727, U3728, U3729, U3730, U3731, U3732, U3733, U3734, U3735, U3736, U3737, U3738, U3739, U3740, U3741, U3742, U3743, U3744, U3745, U3746, U3747, U3748, U3749, U3750, U3751, U3752, U3753, U3754, U3755, U3756, U3757, U3758, U3759, U3760, U3761, U3762, U3763, U3764, U3765, U3766, U3767, U3768, U3769, U3770, U3771, U3772, U3773, U3774, U3775, U3776, U3777, U3778, U3779, U3780, U3781, U3782, U3783, U3784, U3785, U3786, U3787, U3788, U3789, U3790, U3791, U3792, U3793, U3794, U3795, U3796, U3797, U3798, U3799, U3800, U3801, U3802, U3803, U3804, U3805, U3806, U3807, U3808, U3809, U3810, U3811, U3812, U3813, U3814, U3815, U3816, U3817, U3818, U3819, U3820, U3821, U3822, U3823, U3824, U3825, U3826, U3827, U3828, U3829, U3830, U3831, U3832, U3833, U3834, U3835, U3836, U3837, U3838, U3839, U3840, U3841, U3842, U3843, U3844, U3845, U3846, U3847, U3848, U3849, U3850, U3851, U3852, U3853, U3854, U3855, U3856, U3857, U3858, U3859, U3860, U3861, U3862, U3863, U3864, U3865, U3866, U3867, U3868, U3869, U3870, U3871, U3872, U3873, U3874, U3875, U3876, U3877, U3878, U3879, U3880, U3881, U3882, U3883, U3884, U3885, U3886, U3887, U3888, U3889, U3890, U3891, U3892, U3893, U3894, U3895, U3896, U3897, U3898, U3899, U3900, U3901, U3902, U3903, U3904, U3905, U3906, U3907, U3908, U3909, U3910, U3911, U3912, U3913, U3914, U3915, U3916, U3917, U3918, U3919, U3920, U3921, U3922, U3923, U3924, U3925, U3926, U3927, U3928, U3929, U3930, U3931, U3932, U3933, U3934, U3935, U3936, U3937, U3938, U3939, U3940, U3941, U3942, U3943, U3944, U3945, U3946, U3947, U3948, U3949, U3950, U3951, U3952, U3953, U3954, U3955, U3956, U3957, U3958, U3959, U3960, U3961, U3962, U3963, U3964, U3965, U3966, U3967, U3968, U3969, U3970, U3971, U3972, U3973, U3974, U3975, U3976, U3977, U3978, U3979, U3980, U3981, U3982, U3983, U3984, U3985, U3986, U3987, U3988, U3989, U3990, U3991, U3992, U3993, U3994, U3995, U3996, U3997, U3998, U3999, U4000, U4001, U4002, U4003, U4004, U4005, U4006, U4007, U4008, U4009, U4010, U4011, U4012, U4013, U4014, U4015, U4016, U4017, U4018, U4019, U4020, U4021, U4022, U4023, U4024, U4025, U4026, U4027, U4028, U4029, U4030, U4031, U4032, U4033, U4034, U4035, U4036, U4037, U4038, U4039, U4040, U4041, U4042, U4044, U4045, U4046, U4047, U4048, U4049, U4050, U4051, U4052, U4053, U4054, U4055, U4056, U4057, U4058, U4059, U4060, U4061, U4062, U4063, U4064, U4065, U4066, U4067, U4068, U4069, U4070, U4071, U4072, U4073, U4074, U4075, U4076, U4077, U4078, U4079, U4080, U4081, U4082, U4083, U4084, U4085, U4086, U4087, U4088, U4089, U4090, U4091, U4092, U4093, U4094, U4095, U4096, U4097, U4098, U4099, U4100, U4101, U4102, U4103, U4104, U4105, U4106, U4107, U4108, U4109, U4110, U4111, U4112, U4113, U4114, U4115, U4116, U4117, U4118, U4119, U4120, U4121, U4122, U4123, U4124, U4125, U4126, U4127, U4128, U4129, U4130, U4131, U4132, U4133, U4134, U4135, U4136, U4137, U4138, U4139, U4140, U4141, U4142, U4143, U4144, U4145, U4146, U4147, U4148, U4149, U4150, U4151, U4152, U4153, U4154, U4155, U4156, U4157, U4158, U4159, U4160, U4161, U4162, U4163, U4164, U4165, U4166, U4167, U4168, U4169, U4170, U4171, U4172, U4173, U4174, U4175, U4176, U4177, U4178, U4179, U4180, U4181, U4182, U4183, U4184, U4185, U4186, U4187, U4188, U4189, U4190, U4191, U4192, U4193, U4194, U4195, U4196, U4197, U4198, U4199, U4200, U4201, U4202, U4203, U4204, U4205, U4206, U4207, U4208, U4209, U4210, U4211, U4212, U4213, U4214, U4215, U4216, U4217, U4218, U4219, U4220, U4221, U4222, U4223, U4224, U4225, U4226, U4227, U4228, U4229, U4230, U4231, U4232, U4233, U4234, U4235, U4236, U4237, U4238, U4239, U4240, U4241, U4242, U4243, U4244, U4245, U4246, U4247, U4248, U4249, U4250, U4251, U4252, U4253, U4254, U4255, U4256, U4257, U4258, U4259, U4260, U4261, U4262, U4263, U4264, U4265, U4266, U4267, U4268, U4269, U4270, U4271, U4272, U4273, U4274, U4275, U4276, U4277, U4278, U4279, U4280, U4281, U4282, U4283, U4284, U4285, U4286, U4287, U4288, U4289, U4290, U4291, U4292, U4293, U4294, U4295, U4296, U4297, U4298, U4299, U4300, U4301, U4302, U4303, U4304, U4305, U4306, U4307, U4308, U4309, U4310, U4311, U4312, U4313, U4314, U4315, U4316, U4317, U4318, U4319, U4320, U4321, U4322, U4323, U4324, U4325, U4326, U4327, U4328, U4329, U4330, U4331, U4332, U4333, U4334, U4335, U4336, U4337, U4338, U4339, U4340, U4341, U4342, U4343, U4344, U4345, U4346, U4347, U4348, U4349, U4350, U4351, U4352, U4353, U4354, U4355, U4356, U4357, U4358, U4359, U4360, U4361, U4362, U4363, U4364, U4365, U4366, U4367, U4368, U4369, U4370, U4371, U4372, U4373, U4374, U4375, U4376, U4377, U4378, U4379, U4380, U4381, U4382, U4383, U4384, U4385, U4386, U4387, U4388, U4389, U4390, U4391, U4392, U4393, U4394, U4395, U4396, U4397, U4398, U4399, U4400, U4401, U4402, U4403, U4404, U4405, U4406, U4407, U4408, U4409, U4410, U4411, U4412, U4413, U4414, U4415, U4416, U4417, U4418, U4419, U4420, U4421, U4422, U4423, U4424, U4425, U4426, U4427, U4428, U4429, U4430, U4431, U4432, U4433, U4434, U4435, U4436, U4437, U4438, U4439, U4440, U4441, U4442, U4443, U4444, U4445, U4446, U4447, U4448, U4449, U4450, U4451, U4452, U4453, U4454, U4455, U4456, U4457, U4458, U4459, U4460, U4461, U4462, U4463, U4464, U4465, U4466, U4467, U4468, U4469, U4470, U4471, U4472, U4473, U4474, U4475, U4476, U4477, U4478, U4479, U4480, U4481, U4482, U4483, U4484, U4485, U4486, U4487, U4488, U4489, U4490, U4491, U4492, U4493, U4494, U4495, U4496, U4497, U4498, U4499, U4500, U4501, U4502, U4503, U4504, U4505, U4506, U4507, U4508, U4509, U4510, U4511, U4512, U4513, U4514, U4515, U4516, U4517, U4518, U4519, U4520, U4521, U4522, U4523, U4524, U4525, U4526, U4527, U4528, U4529, U4530, U4531, U4532, U4533, U4534, U4535, U4536, U4537, U4538, U4539, U4540, U4541, U4542, U4543, U4544, U4545, U4546, U4547, U4548, U4549, U4550, U4551, U4552, U4553, U4554, U4555, U4556, U4557, U4558, U4559, U4560, U4561, U4562, U4563, U4564, U4565, U4566, U4567, U4568, U4569, U4570, U4571, U4572, U4573, U4574, U4575, U4576, U4577, U4578, U4579, U4580, U4581, U4582, U4583, U4584, U4585, U4586, U4587, U4588, U4589, U4590, U4591, U4592, U4593, U4594, U4595, U4596, U4597, U4598, U4599, U4600, U4601, U4602, U4603, U4604, U4605, U4606, U4607, U4608, U4609, U4610, U4611, U4612, U4613, U4614, U4615, U4616, U4617, U4618, U4619, U4620, U4621, U4622, U4623, U4624, U4625, U4626, U4627, U4628, U4629, U4630, U4631, U4632, U4633, U4634, U4635, U4636, U4637, U4638, U4639, U4640, U4641, U4642, U4643, U4644, U4645, U4646, U4647, U4648, U4649, U4650, U4651, U4652, U4653, U4654, U4655, U4656, U4657, U4658, U4659, U4660, U4661, U4662, U4663, U4664, U4665, U4666, U4667, U4668, U4669, U4670, U4671, U4672, U4673, U4674, U4675, U4676, U4677, U4678, U4679, U4680, U4681, U4682, U4683, U4684, U4685, U4686, U4687, U4688, U4689, U4690, U4691, U4692, U4693, U4694, U4695, U4696, U4697, U4698, U4699, U4700, U4701, U4702, U4703, U4704, U4705, U4706, U4707, U4708, U4709, U4710, U4711, U4712, U4713, U4714, U4715, U4716, U4717, U4718, U4719, U4720, U4721, U4722, U4723, U4724, U4725, U4726, U4727, U4728, U4729, U4730, U4731, U4732, U4733, U4734, U4735, U4736, U4737, U4738, U4739, U4740, U4741, U4742, U4743, U4744, U4745, U4746, U4747, U4748, U4749, U4750, U4751, U4752, U4753, U4754, U4755, U4756, U4757, U4758, U4759, U4760, U4761, U4762, U4763, U4764, U4765, U4766, U4767, U4768, U4769, U4770, U4771, U4772, U4773, U4774, U4775, U4776, U4777, U4778, U4779, U4780, U4781, U4782, U4783, U4784, U4785, U4786, U4787, U4788, U4789, U4790, U4791, U4792, U4793, U4794, U4795, U4796, U4797, U4798, U4799, U4800, U4801, U4802, U4803, U4804, U4805, U4806, U4807, U4808, U4809, U4810, U4811, U4812, U4813, U4814, U4815, U4816, U4817, U4818, U4819, U4820, U4821, U4822, U4823, U4824, U4825, U4826, U4827, U4828, U4829, U4830, U4831, U4832, U4833, U4834, U4835, U4836, U4837, U4838, U4839, U4840, U4841, U4842, U4843, U4844, U4845, U4846, U4847, U4848, U4849, U4850, U4851, U4852, U4853, U4854, U4855, U4856, U4857, U4858, U4859, U4860, U4861, U4862, U4863, U4864, U4865, U4866, U4867, U4868, U4869, U4870, U4871, U4872, U4873, U4874, U4875, U4876, U4877, U4878, U4879, U4880, U4881, U4882, U4883, U4884, U4885, U4886, U4887, U4888, U4889, U4890, U4891, U4892, U4893, U4894, U4895, U4896, U4897, U4898, U4899, U4900, U4901, U4902, U4903, U4904, U4905, U4906, U4907, U4908, U4909, U4910, U4911, U4912, U4913, U4914, U4915, U4916, U4917, U4918, U4919, U4920, U4921, U4922, U4923, U4924, U4925, U4926, U4927, U4928, U4929, U4930, U4931, U4932, U4933, U4934, U4935, U4936, U4937, U4938, U4939, U4940, U4941, U4942, U4943, U4944, U4945, U4946, U4947, U4948, U4949, U4950, U4951, U4952, U4953, U4954, U4955, U4956, U4957, U4958, U4959, U4960, U4961, U4962, U4963, U4964, U4965, U4966, U4967, U4968, U4969, U4970, U4971, U4972, U4973, U4974, U4975, U4976, U4977, U4978, U4979, U4980, U4981, U4982, U4983, U4984, U4985, U4986, U4987, U4988, U4989, U4990, U4991, U4992, U4993, U4994, U4995, U4996, U4997, U4998, U4999, U5000, U5001, U5002, U5003, U5004, U5005, U5006, U5007, U5008, U5009, U5010, U5011, U5012, U5013, U5014, U5015, U5016, U5017, U5018, U5019, U5020, U5021, U5022, U5023, U5024, U5025, U5026, U5027, U5028, U5029, U5030, U5031, U5032, U5033, U5034, U5035, U5036, U5037, U5038, U5039, U5040, U5041, U5042, U5043, U5044, U5045, U5046, U5047, U5048, U5049, U5050, U5051, U5052, U5053, U5054, U5055, U5056, U5057, U5058, U5059, U5060, U5061, U5062, U5063, U5064, U5065, U5066, U5067, U5068, U5069, U5070, U5071, U5072, U5073, U5074, U5075, U5076, U5077, U5078, U5079, U5080, U5081, U5082, U5083, U5084, U5085, U5086, U5087, U5088, U5089, U5090, U5091, U5092, U5093, U5094, U5095, U5096, U5097, U5098, U5099, U5100, U5101, U5102, U5103, U5104, U5105, U5106, U5107, U5108, U5109, U5110, U5111, U5112, U5113, U5114, U5115, U5116, U5117, U5118, U5119, U5120, U5121, U5122, U5123, U5124, U5125, U5126, U5127, U5128, U5129, U5130, U5131, U5132, U5133, U5134, U5135, U5136, U5137, U5138, U5139, U5140, U5141, U5142, U5143, U5144, U5145, U5146, U5147, U5148, U5149, U5150, U5151, U5152, U5153, U5154, U5155, U5156, U5157, U5158, U5159, U5160, U5161, U5162, U5163, U5164, U5165, U5166, U5167, U5168, U5169, U5170, U5171, U5172, U5173, U5174, U5175, U5176, U5177, U5178, U5179, U5180, U5181, U5182, U5183, U5184, U5185, U5186, U5187, U5188, U5189, U5190, U5191, U5192, U5193, U5194, U5195, U5196, U5197, U5198, U5199, U5200, U5201, U5202, U5203, U5204, U5205, U5206, U5207, U5208, U5209, U5210, U5211, U5212, U5213, U5214, U5215, U5216, U5217, U5218, U5219, U5220, U5221, U5222, U5223, U5224, U5225, U5226, U5227, U5228, U5229, U5230, U5231, U5232, U5233, U5234, U5235, U5236, U5237, U5238, U5239, U5240, U5241, U5242, U5243, U5244, U5245, U5246, U5247, U5248, U5249, U5250, U5251, U5252, U5253, U5254, U5255, U5256, U5257, U5258, U5259, U5260, U5261, U5262, U5263, U5264, U5265, U5266, U5267, U5268, U5269, U5270, U5271, U5272, U5273, U5274, U5275, U5276, U5277, U5278, U5279, U5280, U5281, U5282, U5283, U5284, U5285, U5286, U5287, U5288, U5289, U5290, U5291, U5292, U5293, U5294, U5295, U5296, U5297, U5298, U5299, U5300, U5301, U5302, U5303, U5304, U5305, U5306, U5307, U5308, U5309, U5310, U5311, U5312, U5313, U5314, U5315, U5316, U5317, U5318, U5319, U5320, U5321, U5322, U5323, U5324, U5325, U5326, U5327, U5328, U5329, U5330, U5331, U5332, U5333, U5334, U5335, U5336, U5337, U5338, U5339, U5340, U5341, U5342, U5343, U5344, U5345, U5346, U5347, U5348, U5349, U5350, U5351, U5352, U5353, U5354, U5355, U5356, U5357, U5358, U5359, U5360, U5361, U5362, U5363, U5364, U5365, U5366, U5367, U5368, U5369, U5370, U5371, U5372, U5373, U5374, U5375, U5376, U5377, U5378, U5379, U5380, U5381, U5382, U5383, U5384, U5385, U5386, U5387, U5388, U5389, U5390, U5391, U5392, U5393, U5394, U5395, U5396, U5397, U5398, U5399, U5400, U5401, U5402, U5403, U5404, U5405, U5406, U5407, U5408, U5409, U5410, U5411, U5412, U5413, U5414, U5415, U5416, U5417, U5418, U5419, U5420, U5421, U5422, U5423, U5424, U5425, U5426, U5427, U5428, U5429, U5430, U5431, U5432, U5433, U5434, U5435, U5436, U5437, U5438, U5439, U5440, U5441, U5442, U5443, U5444, U5445, U5446, U5447, U5448, U5449, U5450, U5451, U5452, U5453, U5454, U5455, U5456, U5457, U5458, U5459, U5460, U5461, U5462, U5463, U5464, U5465, U5466, U5467, U5468, U5469, U5470, U5471, U5472, U5473, U5474, U5475, U5476, U5477, U5478, U5479, U5480, U5481, U5482, U5483, U5484, U5485, U5486, U5487, U5488, U5489, U5490, U5491, U5492, U5493, U5494, U5495, U5496, U5497, U5498, U5499, U5500, U5501, U5502, U5503, U5504, U5505, U5506, U5507, U5508, U5509, U5510, U5511, U5512, U5513, U5514, U5515, U5516, U5517, U5518, U5519, U5520, U5521, U5522, U5523, U5524, U5525, U5526, U5527, U5528, U5529, U5530, U5531, U5532, U5533, U5534, U5535, U5536, U5537, U5538, U5539, U5540, U5541, U5542, U5543, U5544, U5545, U5546, U5547, U5548, U5549, U5550, U5551, U5552, U5553, U5554, U5555, U5556, U5557, U5558, U5559, U5560, U5561, U5562, U5563, U5564, U5565, U5566, U5567, U5568, U5569, U5570, U5571, U5572, U5573, U5574, U5575, U5576, U5577, U5578, U5579, U5580, U5581, U5582, U5583, U5584, U5585, U5586, U5587, U5588, U5589, U5590, U5591, U5592, U5593, U5594, U5595, U5596, U5597, U5598, U5599, U5600, U5601, U5602, U5603, U5604, U5605, U5606, U5607, U5608, U5609, U5610, U5611, U5612, U5613, U5614, U5615, U5616, U5617, U5618, U5619, U5620, U5621, U5622, U5623, U5624, U5625, U5626, U5627, U5628, U5629, U5630, U5631, U5632, U5633, U5634, U5635, U5636, U5637, U5638, U5639, U5640, U5641, U5642, U5643, U5644, U5645, U5646, U5647, U5648, U5649, U5650, U5651, U5652, U5653, U5654, U5655, U5656, U5657, U5658, U5659, U5660, U5661, U5662, U5663, U5664, U5665, U5666, U5667, U5668, U5669, U5670, U5671, U5672, U5673, U5674, U5675, U5676, U5677, U5678, U5679, U5680, U5681, U5682, U5683, U5684, U5685, U5686, U5687, U5688, U5689, U5690, U5691, U5692, U5693, U5694, U5695, U5696, U5697, U5698, U5699, U5700, U5701, U5702, U5703, U5704, U5705, U5706, U5707, U5708, U5709, U5710, U5711, U5712, U5713, U5714, U5715, U5716, U5717, U5718, U5719, U5720, U5721, U5722, U5723, U5724, U5725, U5726, U5727, U5728, U5729, U5730, U5731, U5732, U5733, U5734, U5735, U5736, U5737, U5738, U5739, U5740, U5741, U5742, U5743, U5744, U5745, U5746, U5747, U5748, U5749, U5750, U5751, U5752, U5753, U5754, U5755, U5756, U5757, U5758, U5759, U5760, U5761, U5762, U5763, U5764, U5765, U5766, U5767, U5768, U5769, U5770, U5771, U5772, U5773, U5774, U5775, U5776, U5777, U5778, U5779, U5780, U5781, U5782, U5783, U5784, U5785, U5786, U5787, U5788, U5789, U5790, U5791, U5792, U5793, U5794, U5795, U5796, U5797, U5798, U5799, U5800, U5801, U5802, U5803, U5804, U5805, U5806, U5807, U5808, U5809, U5810, U5811, U5812, U5813, U5814, U5815, U5816, U5817, U5818, U5819, U5820, U5821, U5822, U5823, U5824, U5825, U5826, U5827, U5828, U5829, U5830, U5831, U5832, U5833, U5834, U5835, U5836, U5837, U5838, U5839, U5840, U5841, U5842, U5843, U5844, U5845, U5846, U5847, U5848, U5849, U5850, U5851, U5852, U5853, U5854, U5855, U5856, U5857, U5858, U5859, U5860, U5861, U5862, U5863, U5864, U5865, U5866, U5867, U5868, U5869, U5870, U5871, U5872, U5873, U5874, U5875, U5876, U5877, U5878, U5879, U5880, U5881, U5882, U5883, U5884, U5885, U5886, U5887, U5888, U5889, U5890, U5891, U5892, U5893, U5894, U5895, U5896, U5897, U5898, U5899, U5900, U5901, U5902, U5903, U5904, U5905, U5906, U5907, U5908, U5909, U5910, U5911, U5912, U5913, U5914, U5915, U5916, U5917, U5918, U5919, U5920, U5921, U5922, U5923, U5924, U5925, U5926, U5927, U5928, U5929, U5930, U5931, U5932, U5933, U5934, U5935, U5936, U5937, U5938, U5939, U5940, U5941, U5942, U5943, U5944, U5945, U5946, U5947, U5948, U5949, U5950, U5951, U5952, U5953, U5954, U5955, U5956, U5957, U5958, U5959, U5960, U5961, U5962, U5963, U5964, U5965, U5966, U5967, U5968, U5969, U5970, U5971, U5972, U5973, U5974, U5975, U5976, U5977, U5978, U5979, U5980, U5981, U5982, U5983, U5984, U5985, U5986, U5987, U5988, U5989, U5990, U5991, U5992, U5993, U5994, U5995, U5996, U5997, U5998, U5999, U6000, U6001, U6002, U6003, U6004, U6005, U6006, U6007, U6008, U6009, U6010, U6011, U6012, U6013, U6014, U6015, U6016, U6017, U6018, U6019, U6020, U6021, U6022, U6023, U6024, U6025, U6026, U6027, U6028, U6029, U6030, U6031, U6032, U6033, U6034, U6035, U6036, U6037, U6038, U6039, U6040, U6041, U6042, U6043, U6044, U6045, U6046, U6047, U6048, U6049, U6050, U6051, U6052, U6053, U6054, U6055, U6056, U6057, U6058, U6059, U6060, U6061, U6062, U6063, U6064, U6065, U6066, U6067, U6068, U6069, U6070, U6071, U6072, U6073, U6074, U6075, U6076, U6077, U6078, U6079, U6080, U6081, U6082, U6083, U6084, U6085, U6086, U6087, U6088, U6089, U6090, U6091, U6092, U6093, U6094, U6095, U6096, U6097, U6098, U6099, U6100, U6101, U6102, U6103, U6104, U6105, U6106, U6107, U6108, U6109, U6110, U6111, U6112, U6113, U6114, U6115, U6116, U6117, U6118, U6119, U6120, U6121, U6122, U6123, U6124, U6125, U6126, U6127, U6128, U6129, U6130, U6131, U6132, U6133, U6134, U6135, U6136, U6137, U6138, U6139, U6140, U6141, U6142, U6143, U6144, U6145, U6146, U6147, U6148, U6149, U6150, U6151, U6152, U6153, U6154, U6155, U6156, U6157, U6158, U6159, U6160, U6161, U6162, U6163, U6164, U6165, U6166, U6167, U6168, U6169, U6170, U6171, U6172, U6173, U6174, U6175, U6176, U6177, U6178, U6179, U6180, U6181, U6182, U6183, U6184, U6185, U6186, U6187, U6188, U6189, U6190, U6191, U6192, U6193, U6194, U6195, U6196, U6197, U6198, U6199, U6200, U6201, U6202, U6203, U6204, U6205, U6206, U6207, U6208, U6209, U6210, U6211, U6212, U6213, U6214, U6215, U6216, U6217, U6218, U6219, U6220, U6221, U6222, U6223, U6224, U6225, U6226, U6227, U6228, U6229, U6230, U6231, U6232, U6233, U6234, U6235, U6236, U6237, U6238, U6239, U6240, U6241, U6242, U6243, U6244, U6245, U6246, U6247, U6248, U6249, U6250, U6251, U6252, U6253, U6254, U6255, U6256, U6257, U6258, U6259, U6260, U6261, U6262, U6263, U6264, U6265, U6266, U6267, U6268, U6269, U6270, U6271, U6272, U6273, U6274, U6275, U6276, U6277, U6278, U6279, U6280, U6281, U6282, U6283, U6284, U6285, U6286, U6287, U6288, U6289, U6290, U6291, U6292, U6293, U6294, U6295, U6296, U6297, U6298, U6299, U6300, U6301, U6302, U6303, U6304, U6305, U6306, U6307, U6308, U6309, U6310, U6311, U6312, U6313, U6314, U6315, U6316, U6317, U6318, U6319, U6320, U6321, U6322, U6323, U3316_in, flip_signal;

  nand ginst1 (ADD_95_U10, REG3_REG_7__SCAN_IN, REG3_REG_3__SCAN_IN, REG3_REG_5__SCAN_IN, REG3_REG_4__SCAN_IN, REG3_REG_6__SCAN_IN);
  not ginst2 (ADD_95_U100, ADD_95_U29);
  not ginst3 (ADD_95_U101, ADD_95_U31);
  not ginst4 (ADD_95_U102, ADD_95_U33);
  not ginst5 (ADD_95_U103, ADD_95_U35);
  not ginst6 (ADD_95_U104, ADD_95_U37);
  not ginst7 (ADD_95_U105, ADD_95_U39);
  not ginst8 (ADD_95_U106, ADD_95_U41);
  not ginst9 (ADD_95_U107, ADD_95_U43);
  not ginst10 (ADD_95_U108, ADD_95_U81);
  not ginst11 (ADD_95_U109, ADD_95_U79);
  not ginst12 (ADD_95_U11, REG3_REG_8__SCAN_IN);
  nand ginst13 (ADD_95_U110, REG3_REG_9__SCAN_IN, ADD_95_U77);
  nand ginst14 (ADD_95_U111, ADD_95_U12, ADD_95_U89);
  nand ginst15 (ADD_95_U112, REG3_REG_8__SCAN_IN, ADD_95_U10);
  nand ginst16 (ADD_95_U113, ADD_95_U11, ADD_95_U88);
  nand ginst17 (ADD_95_U114, REG3_REG_7__SCAN_IN, ADD_95_U78);
  nand ginst18 (ADD_95_U115, ADD_95_U6, ADD_95_U87);
  nand ginst19 (ADD_95_U116, REG3_REG_6__SCAN_IN, ADD_95_U79);
  nand ginst20 (ADD_95_U117, ADD_95_U109, ADD_95_U7);
  nand ginst21 (ADD_95_U118, REG3_REG_5__SCAN_IN, ADD_95_U80);
  nand ginst22 (ADD_95_U119, ADD_95_U8, ADD_95_U86);
  not ginst23 (ADD_95_U12, REG3_REG_9__SCAN_IN);
  nand ginst24 (ADD_95_U120, REG3_REG_4__SCAN_IN, ADD_95_U4);
  nand ginst25 (ADD_95_U121, REG3_REG_3__SCAN_IN, ADD_95_U9);
  nand ginst26 (ADD_95_U122, REG3_REG_28__SCAN_IN, ADD_95_U81);
  nand ginst27 (ADD_95_U123, ADD_95_U108, ADD_95_U44);
  nand ginst28 (ADD_95_U124, REG3_REG_27__SCAN_IN, ADD_95_U43);
  nand ginst29 (ADD_95_U125, ADD_95_U107, ADD_95_U45);
  nand ginst30 (ADD_95_U126, REG3_REG_26__SCAN_IN, ADD_95_U41);
  nand ginst31 (ADD_95_U127, ADD_95_U106, ADD_95_U42);
  nand ginst32 (ADD_95_U128, REG3_REG_25__SCAN_IN, ADD_95_U39);
  nand ginst33 (ADD_95_U129, ADD_95_U105, ADD_95_U40);
  nand ginst34 (ADD_95_U13, ADD_95_U71, ADD_95_U88);
  nand ginst35 (ADD_95_U130, REG3_REG_24__SCAN_IN, ADD_95_U37);
  nand ginst36 (ADD_95_U131, ADD_95_U104, ADD_95_U38);
  nand ginst37 (ADD_95_U132, REG3_REG_23__SCAN_IN, ADD_95_U35);
  nand ginst38 (ADD_95_U133, ADD_95_U103, ADD_95_U36);
  nand ginst39 (ADD_95_U134, REG3_REG_22__SCAN_IN, ADD_95_U33);
  nand ginst40 (ADD_95_U135, ADD_95_U102, ADD_95_U34);
  nand ginst41 (ADD_95_U136, REG3_REG_21__SCAN_IN, ADD_95_U31);
  nand ginst42 (ADD_95_U137, ADD_95_U101, ADD_95_U32);
  nand ginst43 (ADD_95_U138, REG3_REG_20__SCAN_IN, ADD_95_U29);
  nand ginst44 (ADD_95_U139, ADD_95_U100, ADD_95_U30);
  not ginst45 (ADD_95_U14, REG3_REG_11__SCAN_IN);
  nand ginst46 (ADD_95_U140, REG3_REG_19__SCAN_IN, ADD_95_U27);
  nand ginst47 (ADD_95_U141, ADD_95_U28, ADD_95_U99);
  nand ginst48 (ADD_95_U142, REG3_REG_18__SCAN_IN, ADD_95_U25);
  nand ginst49 (ADD_95_U143, ADD_95_U26, ADD_95_U98);
  nand ginst50 (ADD_95_U144, REG3_REG_17__SCAN_IN, ADD_95_U82);
  nand ginst51 (ADD_95_U145, ADD_95_U23, ADD_95_U97);
  nand ginst52 (ADD_95_U146, REG3_REG_16__SCAN_IN, ADD_95_U22);
  nand ginst53 (ADD_95_U147, ADD_95_U24, ADD_95_U96);
  nand ginst54 (ADD_95_U148, REG3_REG_15__SCAN_IN, ADD_95_U83);
  nand ginst55 (ADD_95_U149, ADD_95_U20, ADD_95_U95);
  not ginst56 (ADD_95_U15, REG3_REG_10__SCAN_IN);
  nand ginst57 (ADD_95_U150, REG3_REG_14__SCAN_IN, ADD_95_U19);
  nand ginst58 (ADD_95_U151, ADD_95_U21, ADD_95_U94);
  nand ginst59 (ADD_95_U152, REG3_REG_13__SCAN_IN, ADD_95_U84);
  nand ginst60 (ADD_95_U153, ADD_95_U17, ADD_95_U93);
  nand ginst61 (ADD_95_U154, REG3_REG_12__SCAN_IN, ADD_95_U16);
  nand ginst62 (ADD_95_U155, ADD_95_U18, ADD_95_U92);
  nand ginst63 (ADD_95_U156, REG3_REG_11__SCAN_IN, ADD_95_U85);
  nand ginst64 (ADD_95_U157, ADD_95_U14, ADD_95_U91);
  nand ginst65 (ADD_95_U158, REG3_REG_10__SCAN_IN, ADD_95_U13);
  nand ginst66 (ADD_95_U159, ADD_95_U15, ADD_95_U90);
  nand ginst67 (ADD_95_U16, ADD_95_U72, ADD_95_U90);
  not ginst68 (ADD_95_U17, REG3_REG_13__SCAN_IN);
  not ginst69 (ADD_95_U18, REG3_REG_12__SCAN_IN);
  nand ginst70 (ADD_95_U19, ADD_95_U73, ADD_95_U92);
  not ginst71 (ADD_95_U20, REG3_REG_15__SCAN_IN);
  not ginst72 (ADD_95_U21, REG3_REG_14__SCAN_IN);
  nand ginst73 (ADD_95_U22, ADD_95_U74, ADD_95_U94);
  not ginst74 (ADD_95_U23, REG3_REG_17__SCAN_IN);
  not ginst75 (ADD_95_U24, REG3_REG_16__SCAN_IN);
  nand ginst76 (ADD_95_U25, ADD_95_U75, ADD_95_U96);
  not ginst77 (ADD_95_U26, REG3_REG_18__SCAN_IN);
  nand ginst78 (ADD_95_U27, REG3_REG_18__SCAN_IN, ADD_95_U98);
  not ginst79 (ADD_95_U28, REG3_REG_19__SCAN_IN);
  nand ginst80 (ADD_95_U29, REG3_REG_19__SCAN_IN, ADD_95_U99);
  not ginst81 (ADD_95_U30, REG3_REG_20__SCAN_IN);
  nand ginst82 (ADD_95_U31, REG3_REG_20__SCAN_IN, ADD_95_U100);
  not ginst83 (ADD_95_U32, REG3_REG_21__SCAN_IN);
  nand ginst84 (ADD_95_U33, REG3_REG_21__SCAN_IN, ADD_95_U101);
  not ginst85 (ADD_95_U34, REG3_REG_22__SCAN_IN);
  nand ginst86 (ADD_95_U35, REG3_REG_22__SCAN_IN, ADD_95_U102);
  not ginst87 (ADD_95_U36, REG3_REG_23__SCAN_IN);
  nand ginst88 (ADD_95_U37, REG3_REG_23__SCAN_IN, ADD_95_U103);
  not ginst89 (ADD_95_U38, REG3_REG_24__SCAN_IN);
  nand ginst90 (ADD_95_U39, REG3_REG_24__SCAN_IN, ADD_95_U104);
  not ginst91 (ADD_95_U4, REG3_REG_3__SCAN_IN);
  not ginst92 (ADD_95_U40, REG3_REG_25__SCAN_IN);
  nand ginst93 (ADD_95_U41, REG3_REG_25__SCAN_IN, ADD_95_U105);
  not ginst94 (ADD_95_U42, REG3_REG_26__SCAN_IN);
  nand ginst95 (ADD_95_U43, REG3_REG_26__SCAN_IN, ADD_95_U106);
  not ginst96 (ADD_95_U44, REG3_REG_28__SCAN_IN);
  not ginst97 (ADD_95_U45, REG3_REG_27__SCAN_IN);
  nand ginst98 (ADD_95_U46, ADD_95_U110, ADD_95_U111);
  nand ginst99 (ADD_95_U47, ADD_95_U112, ADD_95_U113);
  nand ginst100 (ADD_95_U48, ADD_95_U114, ADD_95_U115);
  nand ginst101 (ADD_95_U49, ADD_95_U116, ADD_95_U117);
  and ginst102 (ADD_95_U5, ADD_95_U107, ADD_95_U76);
  nand ginst103 (ADD_95_U50, ADD_95_U118, ADD_95_U119);
  nand ginst104 (ADD_95_U51, ADD_95_U120, ADD_95_U121);
  nand ginst105 (ADD_95_U52, ADD_95_U122, ADD_95_U123);
  nand ginst106 (ADD_95_U53, ADD_95_U124, ADD_95_U125);
  nand ginst107 (ADD_95_U54, ADD_95_U126, ADD_95_U127);
  nand ginst108 (ADD_95_U55, ADD_95_U128, ADD_95_U129);
  nand ginst109 (ADD_95_U56, ADD_95_U130, ADD_95_U131);
  nand ginst110 (ADD_95_U57, ADD_95_U132, ADD_95_U133);
  nand ginst111 (ADD_95_U58, ADD_95_U134, ADD_95_U135);
  nand ginst112 (ADD_95_U59, ADD_95_U136, ADD_95_U137);
  not ginst113 (ADD_95_U6, REG3_REG_7__SCAN_IN);
  nand ginst114 (ADD_95_U60, ADD_95_U138, ADD_95_U139);
  nand ginst115 (ADD_95_U61, ADD_95_U140, ADD_95_U141);
  nand ginst116 (ADD_95_U62, ADD_95_U142, ADD_95_U143);
  nand ginst117 (ADD_95_U63, ADD_95_U144, ADD_95_U145);
  nand ginst118 (ADD_95_U64, ADD_95_U146, ADD_95_U147);
  nand ginst119 (ADD_95_U65, ADD_95_U148, ADD_95_U149);
  nand ginst120 (ADD_95_U66, ADD_95_U150, ADD_95_U151);
  nand ginst121 (ADD_95_U67, ADD_95_U152, ADD_95_U153);
  nand ginst122 (ADD_95_U68, ADD_95_U154, ADD_95_U155);
  nand ginst123 (ADD_95_U69, ADD_95_U156, ADD_95_U157);
  not ginst124 (ADD_95_U7, REG3_REG_6__SCAN_IN);
  nand ginst125 (ADD_95_U70, ADD_95_U158, ADD_95_U159);
  and ginst126 (ADD_95_U71, REG3_REG_8__SCAN_IN, REG3_REG_9__SCAN_IN);
  and ginst127 (ADD_95_U72, REG3_REG_10__SCAN_IN, REG3_REG_11__SCAN_IN);
  and ginst128 (ADD_95_U73, REG3_REG_12__SCAN_IN, REG3_REG_13__SCAN_IN);
  and ginst129 (ADD_95_U74, REG3_REG_14__SCAN_IN, REG3_REG_15__SCAN_IN);
  and ginst130 (ADD_95_U75, REG3_REG_16__SCAN_IN, REG3_REG_17__SCAN_IN);
  and ginst131 (ADD_95_U76, REG3_REG_27__SCAN_IN, REG3_REG_28__SCAN_IN);
  nand ginst132 (ADD_95_U77, REG3_REG_8__SCAN_IN, ADD_95_U88);
  nand ginst133 (ADD_95_U78, REG3_REG_3__SCAN_IN, REG3_REG_5__SCAN_IN, REG3_REG_4__SCAN_IN, REG3_REG_6__SCAN_IN);
  nand ginst134 (ADD_95_U79, REG3_REG_3__SCAN_IN, REG3_REG_5__SCAN_IN, REG3_REG_4__SCAN_IN);
  not ginst135 (ADD_95_U8, REG3_REG_5__SCAN_IN);
  nand ginst136 (ADD_95_U80, REG3_REG_3__SCAN_IN, REG3_REG_4__SCAN_IN);
  nand ginst137 (ADD_95_U81, REG3_REG_27__SCAN_IN, ADD_95_U107);
  nand ginst138 (ADD_95_U82, REG3_REG_16__SCAN_IN, ADD_95_U96);
  nand ginst139 (ADD_95_U83, REG3_REG_14__SCAN_IN, ADD_95_U94);
  nand ginst140 (ADD_95_U84, REG3_REG_12__SCAN_IN, ADD_95_U92);
  nand ginst141 (ADD_95_U85, REG3_REG_10__SCAN_IN, ADD_95_U90);
  not ginst142 (ADD_95_U86, ADD_95_U80);
  not ginst143 (ADD_95_U87, ADD_95_U78);
  not ginst144 (ADD_95_U88, ADD_95_U10);
  not ginst145 (ADD_95_U89, ADD_95_U77);
  not ginst146 (ADD_95_U9, REG3_REG_4__SCAN_IN);
  not ginst147 (ADD_95_U90, ADD_95_U13);
  not ginst148 (ADD_95_U91, ADD_95_U85);
  not ginst149 (ADD_95_U92, ADD_95_U16);
  not ginst150 (ADD_95_U93, ADD_95_U84);
  not ginst151 (ADD_95_U94, ADD_95_U19);
  not ginst152 (ADD_95_U95, ADD_95_U83);
  not ginst153 (ADD_95_U96, ADD_95_U22);
  not ginst154 (ADD_95_U97, ADD_95_U82);
  not ginst155 (ADD_95_U98, ADD_95_U25);
  not ginst156 (ADD_95_U99, ADD_95_U27);
  not ginst157 (R1105_U10, U3443);
  nand ginst158 (R1105_U100, R1105_U141, R1105_U142);
  and ginst159 (R1105_U101, R1105_U303, R1105_U304);
  nand ginst160 (R1105_U102, R1105_U137, R1105_U138);
  not ginst161 (R1105_U103, R1105_U82);
  not ginst162 (R1105_U104, R1105_U9);
  nand ginst163 (R1105_U105, R1105_U10, R1105_U9);
  nand ginst164 (R1105_U106, REG2_REG_1__SCAN_IN, R1105_U105);
  not ginst165 (R1105_U107, R1105_U81);
  or ginst166 (R1105_U108, REG2_REG_2__SCAN_IN, U3442);
  nand ginst167 (R1105_U109, R1105_U108, R1105_U81);
  not ginst168 (R1105_U11, REG2_REG_2__SCAN_IN);
  nand ginst169 (R1105_U110, REG2_REG_2__SCAN_IN, U3442);
  not ginst170 (R1105_U111, R1105_U79);
  or ginst171 (R1105_U112, REG2_REG_3__SCAN_IN, U3441);
  nand ginst172 (R1105_U113, R1105_U112, R1105_U79);
  nand ginst173 (R1105_U114, REG2_REG_3__SCAN_IN, U3441);
  not ginst174 (R1105_U115, R1105_U77);
  or ginst175 (R1105_U116, REG2_REG_4__SCAN_IN, U3440);
  nand ginst176 (R1105_U117, R1105_U116, R1105_U77);
  nand ginst177 (R1105_U118, REG2_REG_4__SCAN_IN, U3440);
  not ginst178 (R1105_U119, R1105_U75);
  not ginst179 (R1105_U12, U3442);
  or ginst180 (R1105_U120, REG2_REG_5__SCAN_IN, U3439);
  nand ginst181 (R1105_U121, R1105_U120, R1105_U75);
  nand ginst182 (R1105_U122, REG2_REG_5__SCAN_IN, U3439);
  not ginst183 (R1105_U123, R1105_U73);
  or ginst184 (R1105_U124, REG2_REG_6__SCAN_IN, U3438);
  nand ginst185 (R1105_U125, R1105_U124, R1105_U73);
  nand ginst186 (R1105_U126, REG2_REG_6__SCAN_IN, U3438);
  not ginst187 (R1105_U127, R1105_U71);
  or ginst188 (R1105_U128, REG2_REG_7__SCAN_IN, U3437);
  nand ginst189 (R1105_U129, R1105_U128, R1105_U71);
  not ginst190 (R1105_U13, REG2_REG_3__SCAN_IN);
  nand ginst191 (R1105_U130, REG2_REG_7__SCAN_IN, U3437);
  not ginst192 (R1105_U131, R1105_U69);
  or ginst193 (R1105_U132, REG2_REG_8__SCAN_IN, U3436);
  nand ginst194 (R1105_U133, R1105_U132, R1105_U69);
  nand ginst195 (R1105_U134, REG2_REG_8__SCAN_IN, U3436);
  not ginst196 (R1105_U135, R1105_U67);
  or ginst197 (R1105_U136, REG2_REG_9__SCAN_IN, U3435);
  nand ginst198 (R1105_U137, R1105_U136, R1105_U67);
  nand ginst199 (R1105_U138, REG2_REG_9__SCAN_IN, U3435);
  not ginst200 (R1105_U139, R1105_U102);
  not ginst201 (R1105_U14, U3441);
  or ginst202 (R1105_U140, REG2_REG_10__SCAN_IN, U3452);
  nand ginst203 (R1105_U141, R1105_U102, R1105_U140);
  nand ginst204 (R1105_U142, REG2_REG_10__SCAN_IN, U3452);
  not ginst205 (R1105_U143, R1105_U100);
  or ginst206 (R1105_U144, REG2_REG_11__SCAN_IN, U3451);
  nand ginst207 (R1105_U145, R1105_U100, R1105_U144);
  nand ginst208 (R1105_U146, REG2_REG_11__SCAN_IN, U3451);
  not ginst209 (R1105_U147, R1105_U98);
  or ginst210 (R1105_U148, REG2_REG_12__SCAN_IN, U3450);
  nand ginst211 (R1105_U149, R1105_U148, R1105_U98);
  not ginst212 (R1105_U15, REG2_REG_4__SCAN_IN);
  nand ginst213 (R1105_U150, REG2_REG_12__SCAN_IN, U3450);
  not ginst214 (R1105_U151, R1105_U96);
  or ginst215 (R1105_U152, REG2_REG_13__SCAN_IN, U3449);
  nand ginst216 (R1105_U153, R1105_U152, R1105_U96);
  nand ginst217 (R1105_U154, REG2_REG_13__SCAN_IN, U3449);
  not ginst218 (R1105_U155, R1105_U94);
  or ginst219 (R1105_U156, REG2_REG_14__SCAN_IN, U3448);
  nand ginst220 (R1105_U157, R1105_U156, R1105_U94);
  nand ginst221 (R1105_U158, REG2_REG_14__SCAN_IN, U3448);
  not ginst222 (R1105_U159, R1105_U92);
  not ginst223 (R1105_U16, U3440);
  or ginst224 (R1105_U160, REG2_REG_15__SCAN_IN, U3447);
  nand ginst225 (R1105_U161, R1105_U160, R1105_U92);
  nand ginst226 (R1105_U162, REG2_REG_15__SCAN_IN, U3447);
  not ginst227 (R1105_U163, R1105_U90);
  or ginst228 (R1105_U164, REG2_REG_16__SCAN_IN, U3446);
  nand ginst229 (R1105_U165, R1105_U164, R1105_U90);
  nand ginst230 (R1105_U166, REG2_REG_16__SCAN_IN, U3446);
  not ginst231 (R1105_U167, R1105_U88);
  or ginst232 (R1105_U168, REG2_REG_17__SCAN_IN, U3445);
  nand ginst233 (R1105_U169, R1105_U168, R1105_U88);
  not ginst234 (R1105_U17, REG2_REG_5__SCAN_IN);
  nand ginst235 (R1105_U170, REG2_REG_17__SCAN_IN, U3445);
  not ginst236 (R1105_U171, R1105_U45);
  or ginst237 (R1105_U172, REG2_REG_18__SCAN_IN, U3444);
  nand ginst238 (R1105_U173, R1105_U172, R1105_U45);
  nand ginst239 (R1105_U174, REG2_REG_18__SCAN_IN, U3444);
  nand ginst240 (R1105_U175, R1105_U173, R1105_U64);
  nand ginst241 (R1105_U176, REG2_REG_18__SCAN_IN, U3444);
  nand ginst242 (R1105_U177, R1105_U171, R1105_U176);
  or ginst243 (R1105_U178, REG2_REG_18__SCAN_IN, U3444);
  nand ginst244 (R1105_U179, R1105_U177, R1105_U65);
  not ginst245 (R1105_U18, U3439);
  nand ginst246 (R1105_U180, R1105_U10, R1105_U239);
  nand ginst247 (R1105_U181, R1105_U26, U3435);
  nand ginst248 (R1105_U182, REG2_REG_9__SCAN_IN, R1105_U25);
  nand ginst249 (R1105_U183, R1105_U26, U3435);
  nand ginst250 (R1105_U184, REG2_REG_9__SCAN_IN, R1105_U25);
  nand ginst251 (R1105_U185, R1105_U183, R1105_U184);
  nand ginst252 (R1105_U186, R1105_U66, R1105_U67);
  nand ginst253 (R1105_U187, R1105_U135, R1105_U185);
  nand ginst254 (R1105_U188, R1105_U23, U3436);
  nand ginst255 (R1105_U189, REG2_REG_8__SCAN_IN, R1105_U24);
  not ginst256 (R1105_U19, REG2_REG_6__SCAN_IN);
  nand ginst257 (R1105_U190, R1105_U23, U3436);
  nand ginst258 (R1105_U191, REG2_REG_8__SCAN_IN, R1105_U24);
  nand ginst259 (R1105_U192, R1105_U190, R1105_U191);
  nand ginst260 (R1105_U193, R1105_U68, R1105_U69);
  nand ginst261 (R1105_U194, R1105_U131, R1105_U192);
  nand ginst262 (R1105_U195, R1105_U21, U3437);
  nand ginst263 (R1105_U196, REG2_REG_7__SCAN_IN, R1105_U22);
  nand ginst264 (R1105_U197, R1105_U21, U3437);
  nand ginst265 (R1105_U198, REG2_REG_7__SCAN_IN, R1105_U22);
  nand ginst266 (R1105_U199, R1105_U197, R1105_U198);
  not ginst267 (R1105_U20, U3438);
  nand ginst268 (R1105_U200, R1105_U70, R1105_U71);
  nand ginst269 (R1105_U201, R1105_U127, R1105_U199);
  nand ginst270 (R1105_U202, R1105_U19, U3438);
  nand ginst271 (R1105_U203, REG2_REG_6__SCAN_IN, R1105_U20);
  nand ginst272 (R1105_U204, R1105_U19, U3438);
  nand ginst273 (R1105_U205, REG2_REG_6__SCAN_IN, R1105_U20);
  nand ginst274 (R1105_U206, R1105_U204, R1105_U205);
  nand ginst275 (R1105_U207, R1105_U72, R1105_U73);
  nand ginst276 (R1105_U208, R1105_U123, R1105_U206);
  nand ginst277 (R1105_U209, R1105_U17, U3439);
  not ginst278 (R1105_U21, REG2_REG_7__SCAN_IN);
  nand ginst279 (R1105_U210, REG2_REG_5__SCAN_IN, R1105_U18);
  nand ginst280 (R1105_U211, R1105_U17, U3439);
  nand ginst281 (R1105_U212, REG2_REG_5__SCAN_IN, R1105_U18);
  nand ginst282 (R1105_U213, R1105_U211, R1105_U212);
  nand ginst283 (R1105_U214, R1105_U74, R1105_U75);
  nand ginst284 (R1105_U215, R1105_U119, R1105_U213);
  nand ginst285 (R1105_U216, R1105_U15, U3440);
  nand ginst286 (R1105_U217, REG2_REG_4__SCAN_IN, R1105_U16);
  nand ginst287 (R1105_U218, R1105_U15, U3440);
  nand ginst288 (R1105_U219, REG2_REG_4__SCAN_IN, R1105_U16);
  not ginst289 (R1105_U22, U3437);
  nand ginst290 (R1105_U220, R1105_U218, R1105_U219);
  nand ginst291 (R1105_U221, R1105_U76, R1105_U77);
  nand ginst292 (R1105_U222, R1105_U115, R1105_U220);
  nand ginst293 (R1105_U223, R1105_U13, U3441);
  nand ginst294 (R1105_U224, REG2_REG_3__SCAN_IN, R1105_U14);
  nand ginst295 (R1105_U225, R1105_U13, U3441);
  nand ginst296 (R1105_U226, REG2_REG_3__SCAN_IN, R1105_U14);
  nand ginst297 (R1105_U227, R1105_U225, R1105_U226);
  nand ginst298 (R1105_U228, R1105_U78, R1105_U79);
  nand ginst299 (R1105_U229, R1105_U111, R1105_U227);
  not ginst300 (R1105_U23, REG2_REG_8__SCAN_IN);
  nand ginst301 (R1105_U230, R1105_U11, U3442);
  nand ginst302 (R1105_U231, REG2_REG_2__SCAN_IN, R1105_U12);
  nand ginst303 (R1105_U232, R1105_U11, U3442);
  nand ginst304 (R1105_U233, REG2_REG_2__SCAN_IN, R1105_U12);
  nand ginst305 (R1105_U234, R1105_U232, R1105_U233);
  nand ginst306 (R1105_U235, R1105_U80, R1105_U81);
  nand ginst307 (R1105_U236, R1105_U107, R1105_U234);
  nand ginst308 (R1105_U237, REG2_REG_1__SCAN_IN, R1105_U9);
  nand ginst309 (R1105_U238, R1105_U104, R1105_U8);
  nand ginst310 (R1105_U239, R1105_U237, R1105_U238);
  not ginst311 (R1105_U24, U3436);
  nand ginst312 (R1105_U240, R1105_U8, R1105_U9, U3443);
  nand ginst313 (R1105_U241, REG2_REG_1__SCAN_IN, R1105_U103);
  nand ginst314 (R1105_U242, R1105_U85, U3461);
  nand ginst315 (R1105_U243, REG2_REG_19__SCAN_IN, R1105_U84);
  nand ginst316 (R1105_U244, R1105_U85, U3461);
  nand ginst317 (R1105_U245, REG2_REG_19__SCAN_IN, R1105_U84);
  nand ginst318 (R1105_U246, R1105_U244, R1105_U245);
  nand ginst319 (R1105_U247, R1105_U43, U3444);
  nand ginst320 (R1105_U248, REG2_REG_18__SCAN_IN, R1105_U44);
  nand ginst321 (R1105_U249, R1105_U43, U3444);
  not ginst322 (R1105_U25, U3435);
  nand ginst323 (R1105_U250, REG2_REG_18__SCAN_IN, R1105_U44);
  nand ginst324 (R1105_U251, R1105_U249, R1105_U250);
  nand ginst325 (R1105_U252, R1105_U45, R1105_U86);
  nand ginst326 (R1105_U253, R1105_U171, R1105_U251);
  nand ginst327 (R1105_U254, R1105_U41, U3445);
  nand ginst328 (R1105_U255, REG2_REG_17__SCAN_IN, R1105_U42);
  nand ginst329 (R1105_U256, R1105_U41, U3445);
  nand ginst330 (R1105_U257, REG2_REG_17__SCAN_IN, R1105_U42);
  nand ginst331 (R1105_U258, R1105_U256, R1105_U257);
  nand ginst332 (R1105_U259, R1105_U87, R1105_U88);
  not ginst333 (R1105_U26, REG2_REG_9__SCAN_IN);
  nand ginst334 (R1105_U260, R1105_U167, R1105_U258);
  nand ginst335 (R1105_U261, R1105_U39, U3446);
  nand ginst336 (R1105_U262, REG2_REG_16__SCAN_IN, R1105_U40);
  nand ginst337 (R1105_U263, R1105_U39, U3446);
  nand ginst338 (R1105_U264, REG2_REG_16__SCAN_IN, R1105_U40);
  nand ginst339 (R1105_U265, R1105_U263, R1105_U264);
  nand ginst340 (R1105_U266, R1105_U89, R1105_U90);
  nand ginst341 (R1105_U267, R1105_U163, R1105_U265);
  nand ginst342 (R1105_U268, R1105_U37, U3447);
  nand ginst343 (R1105_U269, REG2_REG_15__SCAN_IN, R1105_U38);
  not ginst344 (R1105_U27, REG2_REG_10__SCAN_IN);
  nand ginst345 (R1105_U270, R1105_U37, U3447);
  nand ginst346 (R1105_U271, REG2_REG_15__SCAN_IN, R1105_U38);
  nand ginst347 (R1105_U272, R1105_U270, R1105_U271);
  nand ginst348 (R1105_U273, R1105_U91, R1105_U92);
  nand ginst349 (R1105_U274, R1105_U159, R1105_U272);
  nand ginst350 (R1105_U275, R1105_U35, U3448);
  nand ginst351 (R1105_U276, REG2_REG_14__SCAN_IN, R1105_U36);
  nand ginst352 (R1105_U277, R1105_U35, U3448);
  nand ginst353 (R1105_U278, REG2_REG_14__SCAN_IN, R1105_U36);
  nand ginst354 (R1105_U279, R1105_U277, R1105_U278);
  not ginst355 (R1105_U28, U3452);
  nand ginst356 (R1105_U280, R1105_U93, R1105_U94);
  nand ginst357 (R1105_U281, R1105_U155, R1105_U279);
  nand ginst358 (R1105_U282, R1105_U33, U3449);
  nand ginst359 (R1105_U283, REG2_REG_13__SCAN_IN, R1105_U34);
  nand ginst360 (R1105_U284, R1105_U33, U3449);
  nand ginst361 (R1105_U285, REG2_REG_13__SCAN_IN, R1105_U34);
  nand ginst362 (R1105_U286, R1105_U284, R1105_U285);
  nand ginst363 (R1105_U287, R1105_U95, R1105_U96);
  nand ginst364 (R1105_U288, R1105_U151, R1105_U286);
  nand ginst365 (R1105_U289, R1105_U31, U3450);
  not ginst366 (R1105_U29, REG2_REG_11__SCAN_IN);
  nand ginst367 (R1105_U290, REG2_REG_12__SCAN_IN, R1105_U32);
  nand ginst368 (R1105_U291, R1105_U31, U3450);
  nand ginst369 (R1105_U292, REG2_REG_12__SCAN_IN, R1105_U32);
  nand ginst370 (R1105_U293, R1105_U291, R1105_U292);
  nand ginst371 (R1105_U294, R1105_U97, R1105_U98);
  nand ginst372 (R1105_U295, R1105_U147, R1105_U293);
  nand ginst373 (R1105_U296, R1105_U29, U3451);
  nand ginst374 (R1105_U297, REG2_REG_11__SCAN_IN, R1105_U30);
  nand ginst375 (R1105_U298, R1105_U29, U3451);
  nand ginst376 (R1105_U299, REG2_REG_11__SCAN_IN, R1105_U30);
  not ginst377 (R1105_U30, U3451);
  nand ginst378 (R1105_U300, R1105_U298, R1105_U299);
  nand ginst379 (R1105_U301, R1105_U100, R1105_U99);
  nand ginst380 (R1105_U302, R1105_U143, R1105_U300);
  nand ginst381 (R1105_U303, R1105_U27, U3452);
  nand ginst382 (R1105_U304, REG2_REG_10__SCAN_IN, R1105_U28);
  nand ginst383 (R1105_U305, R1105_U27, U3452);
  nand ginst384 (R1105_U306, REG2_REG_10__SCAN_IN, R1105_U28);
  nand ginst385 (R1105_U307, R1105_U305, R1105_U306);
  nand ginst386 (R1105_U308, R1105_U101, R1105_U102);
  nand ginst387 (R1105_U309, R1105_U139, R1105_U307);
  not ginst388 (R1105_U31, REG2_REG_12__SCAN_IN);
  nand ginst389 (R1105_U310, R1105_U6, U3453);
  nand ginst390 (R1105_U311, REG2_REG_0__SCAN_IN, R1105_U7);
  not ginst391 (R1105_U32, U3450);
  not ginst392 (R1105_U33, REG2_REG_13__SCAN_IN);
  not ginst393 (R1105_U34, U3449);
  not ginst394 (R1105_U35, REG2_REG_14__SCAN_IN);
  not ginst395 (R1105_U36, U3448);
  not ginst396 (R1105_U37, REG2_REG_15__SCAN_IN);
  not ginst397 (R1105_U38, U3447);
  not ginst398 (R1105_U39, REG2_REG_16__SCAN_IN);
  and ginst399 (R1105_U4, R1105_U175, R1105_U179);
  not ginst400 (R1105_U40, U3446);
  not ginst401 (R1105_U41, REG2_REG_17__SCAN_IN);
  not ginst402 (R1105_U42, U3445);
  not ginst403 (R1105_U43, REG2_REG_18__SCAN_IN);
  not ginst404 (R1105_U44, U3444);
  nand ginst405 (R1105_U45, R1105_U169, R1105_U170);
  nand ginst406 (R1105_U46, R1105_U310, R1105_U311);
  nand ginst407 (R1105_U47, R1105_U186, R1105_U187);
  nand ginst408 (R1105_U48, R1105_U193, R1105_U194);
  nand ginst409 (R1105_U49, R1105_U200, R1105_U201);
  nand ginst410 (R1105_U5, R1105_U180, R1105_U83);
  nand ginst411 (R1105_U50, R1105_U207, R1105_U208);
  nand ginst412 (R1105_U51, R1105_U214, R1105_U215);
  nand ginst413 (R1105_U52, R1105_U221, R1105_U222);
  nand ginst414 (R1105_U53, R1105_U228, R1105_U229);
  nand ginst415 (R1105_U54, R1105_U235, R1105_U236);
  nand ginst416 (R1105_U55, R1105_U252, R1105_U253);
  nand ginst417 (R1105_U56, R1105_U259, R1105_U260);
  nand ginst418 (R1105_U57, R1105_U266, R1105_U267);
  nand ginst419 (R1105_U58, R1105_U273, R1105_U274);
  nand ginst420 (R1105_U59, R1105_U280, R1105_U281);
  not ginst421 (R1105_U6, REG2_REG_0__SCAN_IN);
  nand ginst422 (R1105_U60, R1105_U287, R1105_U288);
  nand ginst423 (R1105_U61, R1105_U294, R1105_U295);
  nand ginst424 (R1105_U62, R1105_U301, R1105_U302);
  nand ginst425 (R1105_U63, R1105_U308, R1105_U309);
  and ginst426 (R1105_U64, R1105_U174, R1105_U242, R1105_U243);
  and ginst427 (R1105_U65, R1105_U178, R1105_U246);
  and ginst428 (R1105_U66, R1105_U181, R1105_U182);
  nand ginst429 (R1105_U67, R1105_U133, R1105_U134);
  and ginst430 (R1105_U68, R1105_U188, R1105_U189);
  nand ginst431 (R1105_U69, R1105_U129, R1105_U130);
  not ginst432 (R1105_U7, U3453);
  and ginst433 (R1105_U70, R1105_U195, R1105_U196);
  nand ginst434 (R1105_U71, R1105_U125, R1105_U126);
  and ginst435 (R1105_U72, R1105_U202, R1105_U203);
  nand ginst436 (R1105_U73, R1105_U121, R1105_U122);
  and ginst437 (R1105_U74, R1105_U209, R1105_U210);
  nand ginst438 (R1105_U75, R1105_U117, R1105_U118);
  and ginst439 (R1105_U76, R1105_U216, R1105_U217);
  nand ginst440 (R1105_U77, R1105_U113, R1105_U114);
  and ginst441 (R1105_U78, R1105_U223, R1105_U224);
  nand ginst442 (R1105_U79, R1105_U109, R1105_U110);
  not ginst443 (R1105_U8, REG2_REG_1__SCAN_IN);
  and ginst444 (R1105_U80, R1105_U230, R1105_U231);
  nand ginst445 (R1105_U81, R1105_U106, R1105_U82);
  nand ginst446 (R1105_U82, R1105_U104, U3443);
  and ginst447 (R1105_U83, R1105_U240, R1105_U241);
  not ginst448 (R1105_U84, U3461);
  not ginst449 (R1105_U85, REG2_REG_19__SCAN_IN);
  and ginst450 (R1105_U86, R1105_U247, R1105_U248);
  and ginst451 (R1105_U87, R1105_U254, R1105_U255);
  nand ginst452 (R1105_U88, R1105_U165, R1105_U166);
  and ginst453 (R1105_U89, R1105_U261, R1105_U262);
  nand ginst454 (R1105_U9, REG2_REG_0__SCAN_IN, U3453);
  nand ginst455 (R1105_U90, R1105_U161, R1105_U162);
  and ginst456 (R1105_U91, R1105_U268, R1105_U269);
  nand ginst457 (R1105_U92, R1105_U157, R1105_U158);
  and ginst458 (R1105_U93, R1105_U275, R1105_U276);
  nand ginst459 (R1105_U94, R1105_U153, R1105_U154);
  and ginst460 (R1105_U95, R1105_U282, R1105_U283);
  nand ginst461 (R1105_U96, R1105_U149, R1105_U150);
  and ginst462 (R1105_U97, R1105_U289, R1105_U290);
  nand ginst463 (R1105_U98, R1105_U145, R1105_U146);
  and ginst464 (R1105_U99, R1105_U296, R1105_U297);
  and ginst465 (R1117_U10, R1117_U273, R1117_U274);
  not ginst466 (R1117_U100, U4030);
  not ginst467 (R1117_U101, U3051);
  nand ginst468 (R1117_U102, R1117_U211, R1117_U431);
  nand ginst469 (R1117_U103, R1117_U297, R1117_U346);
  nand ginst470 (R1117_U104, R1117_U157, R1117_U356);
  nand ginst471 (R1117_U105, R1117_U289, R1117_U344);
  nand ginst472 (R1117_U106, R1117_U315, R1117_U94);
  nand ginst473 (R1117_U107, R1117_U360, R1117_U88);
  not ginst474 (R1117_U108, U3074);
  nand ginst475 (R1117_U109, R1117_U427, R1117_U428);
  and ginst476 (R1117_U11, R1117_U186, R1117_U290);
  nand ginst477 (R1117_U110, R1117_U443, R1117_U444);
  nand ginst478 (R1117_U111, R1117_U448, R1117_U449);
  nand ginst479 (R1117_U112, R1117_U466, R1117_U467);
  nand ginst480 (R1117_U113, R1117_U471, R1117_U472);
  nand ginst481 (R1117_U114, R1117_U476, R1117_U477);
  nand ginst482 (R1117_U115, R1117_U481, R1117_U482);
  nand ginst483 (R1117_U116, R1117_U486, R1117_U487);
  nand ginst484 (R1117_U117, R1117_U502, R1117_U503);
  nand ginst485 (R1117_U118, R1117_U507, R1117_U508);
  nand ginst486 (R1117_U119, R1117_U386, R1117_U387);
  and ginst487 (R1117_U12, R1117_U291, R1117_U292);
  nand ginst488 (R1117_U120, R1117_U395, R1117_U396);
  nand ginst489 (R1117_U121, R1117_U402, R1117_U403);
  nand ginst490 (R1117_U122, R1117_U406, R1117_U407);
  nand ginst491 (R1117_U123, R1117_U415, R1117_U416);
  nand ginst492 (R1117_U124, R1117_U438, R1117_U439);
  nand ginst493 (R1117_U125, R1117_U457, R1117_U458);
  nand ginst494 (R1117_U126, R1117_U461, R1117_U462);
  nand ginst495 (R1117_U127, R1117_U493, R1117_U494);
  nand ginst496 (R1117_U128, R1117_U497, R1117_U498);
  nand ginst497 (R1117_U129, R1117_U514, R1117_U515);
  and ginst498 (R1117_U13, R1117_U211, R1117_U304);
  and ginst499 (R1117_U130, R1117_U212, R1117_U222);
  and ginst500 (R1117_U131, R1117_U224, R1117_U225);
  and ginst501 (R1117_U132, R1117_U14, R1117_U15);
  and ginst502 (R1117_U133, R1117_U238, R1117_U239);
  and ginst503 (R1117_U134, R1117_U133, R1117_U338);
  and ginst504 (R1117_U135, R1117_U33, R1117_U388, R1117_U389);
  and ginst505 (R1117_U136, R1117_U214, R1117_U392);
  and ginst506 (R1117_U137, R1117_U254, R1117_U6);
  and ginst507 (R1117_U138, R1117_U213, R1117_U399);
  and ginst508 (R1117_U139, R1117_U408, R1117_U409, R1117_U41);
  and ginst509 (R1117_U14, R1117_U213, R1117_U226, R1117_U231);
  and ginst510 (R1117_U140, R1117_U212, R1117_U412);
  and ginst511 (R1117_U141, R1117_U19, R1117_U270);
  and ginst512 (R1117_U142, R1117_U17, R1117_U282);
  and ginst513 (R1117_U143, R1117_U283, R1117_U343);
  and ginst514 (R1117_U144, R1117_U21, R1117_U298);
  and ginst515 (R1117_U145, R1117_U299, R1117_U348);
  and ginst516 (R1117_U146, R1117_U306, R1117_U307);
  and ginst517 (R1117_U147, R1117_U308, R1117_U419);
  and ginst518 (R1117_U148, R1117_U22, R1117_U307);
  and ginst519 (R1117_U149, R1117_U148, R1117_U306, R1117_U309);
  and ginst520 (R1117_U15, R1117_U214, R1117_U236);
  and ginst521 (R1117_U150, R1117_U179, R1117_U375);
  nand ginst522 (R1117_U151, R1117_U424, R1117_U425);
  and ginst523 (R1117_U152, R1117_U102, R1117_U211);
  nand ginst524 (R1117_U153, R1117_U440, R1117_U441);
  nand ginst525 (R1117_U154, R1117_U445, R1117_U446);
  and ginst526 (R1117_U155, R1117_U67, U3058);
  and ginst527 (R1117_U156, R1117_U20, R1117_U295);
  and ginst528 (R1117_U157, R1117_U349, R1117_U68);
  and ginst529 (R1117_U158, R1117_U12, R1117_U311);
  nand ginst530 (R1117_U159, R1117_U463, R1117_U464);
  and ginst531 (R1117_U16, R1117_U241, R1117_U7);
  nand ginst532 (R1117_U160, R1117_U468, R1117_U469);
  nand ginst533 (R1117_U161, R1117_U473, R1117_U474);
  nand ginst534 (R1117_U162, R1117_U478, R1117_U479);
  nand ginst535 (R1117_U163, R1117_U483, R1117_U484);
  and ginst536 (R1117_U164, R1117_U10, R1117_U321);
  and ginst537 (R1117_U165, R1117_U209, R1117_U490);
  nand ginst538 (R1117_U166, R1117_U499, R1117_U500);
  nand ginst539 (R1117_U167, R1117_U504, R1117_U505);
  and ginst540 (R1117_U168, R1117_U330, R1117_U8);
  and ginst541 (R1117_U169, R1117_U208, R1117_U511);
  and ginst542 (R1117_U17, R1117_U277, R1117_U9);
  and ginst543 (R1117_U170, R1117_U384, R1117_U385);
  nand ginst544 (R1117_U171, R1117_U134, R1117_U337);
  and ginst545 (R1117_U172, R1117_U393, R1117_U394);
  and ginst546 (R1117_U173, R1117_U400, R1117_U401);
  and ginst547 (R1117_U174, R1117_U404, R1117_U405);
  nand ginst548 (R1117_U175, R1117_U131, R1117_U368);
  and ginst549 (R1117_U176, R1117_U413, R1117_U414);
  not ginst550 (R1117_U177, U4040);
  not ginst551 (R1117_U178, U3052);
  and ginst552 (R1117_U179, R1117_U422, R1117_U423);
  and ginst553 (R1117_U18, R1117_U11, R1117_U295);
  nand ginst554 (R1117_U180, R1117_U146, R1117_U376);
  and ginst555 (R1117_U181, R1117_U434, R1117_U435);
  and ginst556 (R1117_U182, R1117_U436, R1117_U437);
  nand ginst557 (R1117_U183, R1117_U301, R1117_U302);
  nand ginst558 (R1117_U184, R1117_U145, R1117_U358);
  nand ginst559 (R1117_U185, R1117_U347, R1117_U354);
  nand ginst560 (R1117_U186, R1117_U64, U4035);
  and ginst561 (R1117_U187, R1117_U455, R1117_U456);
  and ginst562 (R1117_U188, R1117_U459, R1117_U460);
  nand ginst563 (R1117_U189, R1117_U345, R1117_U352);
  and ginst564 (R1117_U19, R1117_U16, R1117_U268);
  nand ginst565 (R1117_U190, R1117_U350, R1117_U73);
  not ginst566 (R1117_U191, U3468);
  nand ginst567 (R1117_U192, R1117_U108, U3464);
  nand ginst568 (R1117_U193, R1117_U336, R1117_U380);
  nand ginst569 (R1117_U194, R1117_U143, R1117_U342);
  nand ginst570 (R1117_U195, R1117_U279, R1117_U95);
  and ginst571 (R1117_U196, R1117_U491, R1117_U492);
  and ginst572 (R1117_U197, R1117_U495, R1117_U496);
  nand ginst573 (R1117_U198, R1117_U271, R1117_U341, R1117_U366);
  nand ginst574 (R1117_U199, R1117_U364, R1117_U90);
  and ginst575 (R1117_U20, R1117_U286, R1117_U288);
  nand ginst576 (R1117_U200, R1117_U267, R1117_U362);
  and ginst577 (R1117_U201, R1117_U512, R1117_U513);
  not ginst578 (R1117_U202, R1117_U102);
  nand ginst579 (R1117_U203, R1117_U147, R1117_U180);
  nand ginst580 (R1117_U204, R1117_U191, R1117_U192);
  not ginst581 (R1117_U205, R1117_U59);
  not ginst582 (R1117_U206, R1117_U41);
  not ginst583 (R1117_U207, R1117_U33);
  nand ginst584 (R1117_U208, R1117_U85, U3486);
  nand ginst585 (R1117_U209, R1117_U92, U3496);
  and ginst586 (R1117_U21, R1117_U18, R1117_U20);
  not ginst587 (R1117_U210, R1117_U186);
  nand ginst588 (R1117_U211, R1117_U58, U4031);
  nand ginst589 (R1117_U212, R1117_U40, U3470);
  nand ginst590 (R1117_U213, R1117_U48, U3476);
  nand ginst591 (R1117_U214, R1117_U32, U3480);
  not ginst592 (R1117_U215, R1117_U94);
  not ginst593 (R1117_U216, R1117_U68);
  not ginst594 (R1117_U217, R1117_U50);
  not ginst595 (R1117_U218, R1117_U88);
  not ginst596 (R1117_U219, R1117_U192);
  and ginst597 (R1117_U22, R1117_U420, R1117_U421);
  nand ginst598 (R1117_U220, R1117_U192, U3075);
  not ginst599 (R1117_U221, R1117_U56);
  nand ginst600 (R1117_U222, R1117_U42, U3472);
  nand ginst601 (R1117_U223, R1117_U41, R1117_U42);
  nand ginst602 (R1117_U224, R1117_U223, R1117_U46);
  nand ginst603 (R1117_U225, R1117_U206, U3061);
  nand ginst604 (R1117_U226, R1117_U47, U3478);
  nand ginst605 (R1117_U227, R1117_U36, U3068);
  nand ginst606 (R1117_U228, R1117_U35, U3064);
  nand ginst607 (R1117_U229, R1117_U213, R1117_U217);
  nand ginst608 (R1117_U23, R1117_U328, R1117_U331);
  nand ginst609 (R1117_U230, R1117_U229, R1117_U6);
  nand ginst610 (R1117_U231, R1117_U49, U3474);
  nand ginst611 (R1117_U232, R1117_U47, U3478);
  nand ginst612 (R1117_U233, R1117_U14, R1117_U175);
  not ginst613 (R1117_U234, R1117_U51);
  not ginst614 (R1117_U235, R1117_U54);
  nand ginst615 (R1117_U236, R1117_U34, U3482);
  nand ginst616 (R1117_U237, R1117_U33, R1117_U34);
  nand ginst617 (R1117_U238, R1117_U237, R1117_U39);
  nand ginst618 (R1117_U239, R1117_U207, U3081);
  nand ginst619 (R1117_U24, R1117_U319, R1117_U322);
  not ginst620 (R1117_U240, R1117_U171);
  nand ginst621 (R1117_U241, R1117_U53, U3484);
  nand ginst622 (R1117_U242, R1117_U241, R1117_U88);
  nand ginst623 (R1117_U243, R1117_U235, R1117_U33);
  nand ginst624 (R1117_U244, R1117_U136, R1117_U243);
  nand ginst625 (R1117_U245, R1117_U214, R1117_U54);
  nand ginst626 (R1117_U246, R1117_U135, R1117_U245);
  nand ginst627 (R1117_U247, R1117_U214, R1117_U33);
  nand ginst628 (R1117_U248, R1117_U175, R1117_U231);
  not ginst629 (R1117_U249, R1117_U55);
  nand ginst630 (R1117_U25, R1117_U382, R1117_U383, R1117_U453, R1117_U454);
  nand ginst631 (R1117_U250, R1117_U35, U3064);
  nand ginst632 (R1117_U251, R1117_U249, R1117_U250);
  nand ginst633 (R1117_U252, R1117_U138, R1117_U251);
  nand ginst634 (R1117_U253, R1117_U213, R1117_U55);
  nand ginst635 (R1117_U254, R1117_U47, U3478);
  nand ginst636 (R1117_U255, R1117_U137, R1117_U253);
  nand ginst637 (R1117_U256, R1117_U35, U3064);
  nand ginst638 (R1117_U257, R1117_U213, R1117_U256);
  nand ginst639 (R1117_U258, R1117_U231, R1117_U50);
  nand ginst640 (R1117_U259, R1117_U140, R1117_U372);
  nand ginst641 (R1117_U26, R1117_U150, R1117_U203);
  nand ginst642 (R1117_U260, R1117_U212, R1117_U41);
  nand ginst643 (R1117_U261, R1117_U84, U3488);
  nand ginst644 (R1117_U262, R1117_U86, U3060);
  nand ginst645 (R1117_U263, R1117_U87, U3059);
  nand ginst646 (R1117_U264, R1117_U218, R1117_U7);
  nand ginst647 (R1117_U265, R1117_U264, R1117_U8);
  nand ginst648 (R1117_U266, R1117_U84, U3488);
  nand ginst649 (R1117_U267, R1117_U265, R1117_U266);
  nand ginst650 (R1117_U268, R1117_U89, U3490);
  nand ginst651 (R1117_U269, R1117_U83, U3069);
  nand ginst652 (R1117_U27, R1117_U259, R1117_U371);
  nand ginst653 (R1117_U270, R1117_U81, U3492);
  nand ginst654 (R1117_U271, R1117_U82, U3077);
  nand ginst655 (R1117_U272, R1117_U91, U3498);
  nand ginst656 (R1117_U273, R1117_U78, U3070);
  nand ginst657 (R1117_U274, R1117_U79, U3071);
  nand ginst658 (R1117_U275, R1117_U215, R1117_U9);
  nand ginst659 (R1117_U276, R1117_U10, R1117_U275);
  nand ginst660 (R1117_U277, R1117_U93, U3494);
  nand ginst661 (R1117_U278, R1117_U91, U3498);
  nand ginst662 (R1117_U279, R1117_U17, R1117_U198);
  nand ginst663 (R1117_U28, R1117_U252, R1117_U255);
  not ginst664 (R1117_U280, R1117_U95);
  not ginst665 (R1117_U281, R1117_U195);
  nand ginst666 (R1117_U282, R1117_U76, U3500);
  nand ginst667 (R1117_U283, R1117_U77, U3066);
  not ginst668 (R1117_U284, R1117_U194);
  nand ginst669 (R1117_U285, R1117_U75, U3502);
  nand ginst670 (R1117_U286, R1117_U71, U3504);
  not ginst671 (R1117_U287, R1117_U73);
  nand ginst672 (R1117_U288, R1117_U70, U4037);
  nand ginst673 (R1117_U289, R1117_U72, U3073);
  nand ginst674 (R1117_U29, R1117_U244, R1117_U246);
  nand ginst675 (R1117_U290, R1117_U63, U4034);
  nand ginst676 (R1117_U291, R1117_U66, U3063);
  nand ginst677 (R1117_U292, R1117_U67, U3058);
  nand ginst678 (R1117_U293, R1117_U11, R1117_U216);
  nand ginst679 (R1117_U294, R1117_U12, R1117_U293);
  nand ginst680 (R1117_U295, R1117_U65, U4036);
  nand ginst681 (R1117_U296, R1117_U63, U4034);
  nand ginst682 (R1117_U297, R1117_U294, R1117_U296);
  nand ginst683 (R1117_U298, R1117_U61, U4033);
  nand ginst684 (R1117_U299, R1117_U62, U3062);
  nand ginst685 (R1117_U30, R1117_U192, R1117_U334);
  nand ginst686 (R1117_U300, R1117_U98, U4032);
  nand ginst687 (R1117_U301, R1117_U184, R1117_U300);
  nand ginst688 (R1117_U302, R1117_U97, U3055);
  not ginst689 (R1117_U303, R1117_U183);
  nand ginst690 (R1117_U304, R1117_U60, U4030);
  nand ginst691 (R1117_U305, R1117_U59, R1117_U60);
  nand ginst692 (R1117_U306, R1117_U100, R1117_U305);
  nand ginst693 (R1117_U307, R1117_U205, U3050);
  nand ginst694 (R1117_U308, R1117_U101, U4029);
  nand ginst695 (R1117_U309, R1117_U57, U3051);
  and ginst696 (R1117_U31, R1117_U373, R1117_U379);
  nand ginst697 (R1117_U310, R1117_U211, R1117_U59);
  nand ginst698 (R1117_U311, R1117_U63, U4034);
  nand ginst699 (R1117_U312, R1117_U67, U3058);
  nand ginst700 (R1117_U313, R1117_U186, R1117_U312);
  nand ginst701 (R1117_U314, R1117_U295, R1117_U68);
  nand ginst702 (R1117_U315, R1117_U198, R1117_U277);
  not ginst703 (R1117_U316, R1117_U106);
  nand ginst704 (R1117_U317, R1117_U79, U3071);
  nand ginst705 (R1117_U318, R1117_U316, R1117_U317);
  nand ginst706 (R1117_U319, R1117_U165, R1117_U318);
  not ginst707 (R1117_U32, U3067);
  nand ginst708 (R1117_U320, R1117_U106, R1117_U209);
  nand ginst709 (R1117_U321, R1117_U91, U3498);
  nand ginst710 (R1117_U322, R1117_U164, R1117_U320);
  nand ginst711 (R1117_U323, R1117_U79, U3071);
  nand ginst712 (R1117_U324, R1117_U209, R1117_U323);
  nand ginst713 (R1117_U325, R1117_U277, R1117_U94);
  nand ginst714 (R1117_U326, R1117_U87, U3059);
  nand ginst715 (R1117_U327, R1117_U326, R1117_U361);
  nand ginst716 (R1117_U328, R1117_U169, R1117_U327);
  nand ginst717 (R1117_U329, R1117_U107, R1117_U208);
  nand ginst718 (R1117_U33, R1117_U38, U3067);
  nand ginst719 (R1117_U330, R1117_U84, U3488);
  nand ginst720 (R1117_U331, R1117_U168, R1117_U329);
  nand ginst721 (R1117_U332, R1117_U87, U3059);
  nand ginst722 (R1117_U333, R1117_U208, R1117_U332);
  nand ginst723 (R1117_U334, R1117_U44, U3074);
  nand ginst724 (R1117_U335, R1117_U191, U3075);
  nand ginst725 (R1117_U336, R1117_U96, U3079);
  nand ginst726 (R1117_U337, R1117_U132, R1117_U175);
  nand ginst727 (R1117_U338, R1117_U15, R1117_U234);
  nand ginst728 (R1117_U339, R1117_U267, R1117_U269);
  not ginst729 (R1117_U34, U3081);
  not ginst730 (R1117_U340, R1117_U90);
  nand ginst731 (R1117_U341, R1117_U270, R1117_U340);
  nand ginst732 (R1117_U342, R1117_U142, R1117_U198);
  nand ginst733 (R1117_U343, R1117_U280, R1117_U282);
  nand ginst734 (R1117_U344, R1117_U287, R1117_U288);
  not ginst735 (R1117_U345, R1117_U105);
  nand ginst736 (R1117_U346, R1117_U105, R1117_U18);
  not ginst737 (R1117_U347, R1117_U103);
  nand ginst738 (R1117_U348, R1117_U103, R1117_U298);
  nand ginst739 (R1117_U349, R1117_U105, R1117_U295);
  not ginst740 (R1117_U35, U3476);
  nand ginst741 (R1117_U350, R1117_U193, R1117_U286);
  not ginst742 (R1117_U351, R1117_U190);
  nand ginst743 (R1117_U352, R1117_U193, R1117_U20);
  not ginst744 (R1117_U353, R1117_U189);
  nand ginst745 (R1117_U354, R1117_U193, R1117_U21);
  not ginst746 (R1117_U355, R1117_U185);
  nand ginst747 (R1117_U356, R1117_U156, R1117_U193);
  not ginst748 (R1117_U357, R1117_U104);
  nand ginst749 (R1117_U358, R1117_U144, R1117_U193);
  not ginst750 (R1117_U359, R1117_U184);
  not ginst751 (R1117_U36, U3478);
  nand ginst752 (R1117_U360, R1117_U171, R1117_U241);
  not ginst753 (R1117_U361, R1117_U107);
  nand ginst754 (R1117_U362, R1117_U16, R1117_U171);
  not ginst755 (R1117_U363, R1117_U200);
  nand ginst756 (R1117_U364, R1117_U171, R1117_U19);
  not ginst757 (R1117_U365, R1117_U199);
  nand ginst758 (R1117_U366, R1117_U141, R1117_U171);
  not ginst759 (R1117_U367, R1117_U198);
  nand ginst760 (R1117_U368, R1117_U130, R1117_U56);
  not ginst761 (R1117_U369, R1117_U175);
  not ginst762 (R1117_U37, U3474);
  nand ginst763 (R1117_U370, R1117_U212, R1117_U56);
  nand ginst764 (R1117_U371, R1117_U139, R1117_U370);
  nand ginst765 (R1117_U372, R1117_U221, R1117_U41);
  nand ginst766 (R1117_U373, R1117_U152, R1117_U183);
  nand ginst767 (R1117_U374, R1117_U13, R1117_U183);
  nand ginst768 (R1117_U375, R1117_U149, R1117_U374);
  nand ginst769 (R1117_U376, R1117_U13, R1117_U183);
  not ginst770 (R1117_U377, R1117_U180);
  nand ginst771 (R1117_U378, R1117_U183, R1117_U202);
  nand ginst772 (R1117_U379, R1117_U181, R1117_U378);
  not ginst773 (R1117_U38, U3480);
  nand ginst774 (R1117_U380, R1117_U194, R1117_U285);
  not ginst775 (R1117_U381, R1117_U193);
  nand ginst776 (R1117_U382, R1117_U155, R1117_U452);
  nand ginst777 (R1117_U383, R1117_U158, R1117_U357);
  nand ginst778 (R1117_U384, R1117_U53, U3484);
  nand ginst779 (R1117_U385, R1117_U52, U3080);
  nand ginst780 (R1117_U386, R1117_U171, R1117_U242);
  nand ginst781 (R1117_U387, R1117_U170, R1117_U240);
  nand ginst782 (R1117_U388, R1117_U34, U3482);
  nand ginst783 (R1117_U389, R1117_U39, U3081);
  not ginst784 (R1117_U39, U3482);
  nand ginst785 (R1117_U390, R1117_U34, U3482);
  nand ginst786 (R1117_U391, R1117_U39, U3081);
  nand ginst787 (R1117_U392, R1117_U390, R1117_U391);
  nand ginst788 (R1117_U393, R1117_U32, U3480);
  nand ginst789 (R1117_U394, R1117_U38, U3067);
  nand ginst790 (R1117_U395, R1117_U247, R1117_U54);
  nand ginst791 (R1117_U396, R1117_U172, R1117_U235);
  nand ginst792 (R1117_U397, R1117_U47, U3478);
  nand ginst793 (R1117_U398, R1117_U36, U3068);
  nand ginst794 (R1117_U399, R1117_U397, R1117_U398);
  not ginst795 (R1117_U40, U3065);
  nand ginst796 (R1117_U400, R1117_U48, U3476);
  nand ginst797 (R1117_U401, R1117_U35, U3064);
  nand ginst798 (R1117_U402, R1117_U257, R1117_U55);
  nand ginst799 (R1117_U403, R1117_U173, R1117_U249);
  nand ginst800 (R1117_U404, R1117_U49, U3474);
  nand ginst801 (R1117_U405, R1117_U37, U3057);
  nand ginst802 (R1117_U406, R1117_U175, R1117_U258);
  nand ginst803 (R1117_U407, R1117_U174, R1117_U369);
  nand ginst804 (R1117_U408, R1117_U42, U3472);
  nand ginst805 (R1117_U409, R1117_U46, U3061);
  nand ginst806 (R1117_U41, R1117_U43, U3065);
  nand ginst807 (R1117_U410, R1117_U42, U3472);
  nand ginst808 (R1117_U411, R1117_U46, U3061);
  nand ginst809 (R1117_U412, R1117_U410, R1117_U411);
  nand ginst810 (R1117_U413, R1117_U40, U3470);
  nand ginst811 (R1117_U414, R1117_U43, U3065);
  nand ginst812 (R1117_U415, R1117_U260, R1117_U56);
  nand ginst813 (R1117_U416, R1117_U176, R1117_U221);
  nand ginst814 (R1117_U417, R1117_U178, U4040);
  nand ginst815 (R1117_U418, R1117_U177, U3052);
  nand ginst816 (R1117_U419, R1117_U417, R1117_U418);
  not ginst817 (R1117_U42, U3061);
  nand ginst818 (R1117_U420, R1117_U178, U4040);
  nand ginst819 (R1117_U421, R1117_U177, U3052);
  nand ginst820 (R1117_U422, R1117_U419, R1117_U57, U3051);
  nand ginst821 (R1117_U423, R1117_U101, R1117_U22, U4029);
  nand ginst822 (R1117_U424, R1117_U101, U4029);
  nand ginst823 (R1117_U425, R1117_U57, U3051);
  not ginst824 (R1117_U426, R1117_U151);
  nand ginst825 (R1117_U427, R1117_U377, R1117_U426);
  nand ginst826 (R1117_U428, R1117_U151, R1117_U180);
  nand ginst827 (R1117_U429, R1117_U60, U4030);
  not ginst828 (R1117_U43, U3470);
  nand ginst829 (R1117_U430, R1117_U100, U3050);
  nand ginst830 (R1117_U431, R1117_U429, R1117_U430);
  nand ginst831 (R1117_U432, R1117_U60, U4030);
  nand ginst832 (R1117_U433, R1117_U100, U3050);
  nand ginst833 (R1117_U434, R1117_U432, R1117_U433, R1117_U59);
  nand ginst834 (R1117_U435, R1117_U205, R1117_U431);
  nand ginst835 (R1117_U436, R1117_U58, U4031);
  nand ginst836 (R1117_U437, R1117_U99, U3054);
  nand ginst837 (R1117_U438, R1117_U183, R1117_U310);
  nand ginst838 (R1117_U439, R1117_U182, R1117_U303);
  not ginst839 (R1117_U44, U3464);
  nand ginst840 (R1117_U440, R1117_U98, U4032);
  nand ginst841 (R1117_U441, R1117_U97, U3055);
  not ginst842 (R1117_U442, R1117_U153);
  nand ginst843 (R1117_U443, R1117_U359, R1117_U442);
  nand ginst844 (R1117_U444, R1117_U153, R1117_U184);
  nand ginst845 (R1117_U445, R1117_U61, U4033);
  nand ginst846 (R1117_U446, R1117_U62, U3062);
  not ginst847 (R1117_U447, R1117_U154);
  nand ginst848 (R1117_U448, R1117_U355, R1117_U447);
  nand ginst849 (R1117_U449, R1117_U154, R1117_U185);
  not ginst850 (R1117_U45, U3075);
  nand ginst851 (R1117_U450, R1117_U63, U4034);
  nand ginst852 (R1117_U451, R1117_U66, U3063);
  nand ginst853 (R1117_U452, R1117_U450, R1117_U451);
  nand ginst854 (R1117_U453, R1117_U104, R1117_U186, R1117_U452);
  nand ginst855 (R1117_U454, R1117_U12, R1117_U210, R1117_U311);
  nand ginst856 (R1117_U455, R1117_U64, U4035);
  nand ginst857 (R1117_U456, R1117_U67, U3058);
  nand ginst858 (R1117_U457, R1117_U104, R1117_U313);
  nand ginst859 (R1117_U458, R1117_U187, R1117_U357);
  nand ginst860 (R1117_U459, R1117_U65, U4036);
  not ginst861 (R1117_U46, U3472);
  nand ginst862 (R1117_U460, R1117_U69, U3072);
  nand ginst863 (R1117_U461, R1117_U189, R1117_U314);
  nand ginst864 (R1117_U462, R1117_U188, R1117_U353);
  nand ginst865 (R1117_U463, R1117_U70, U4037);
  nand ginst866 (R1117_U464, R1117_U72, U3073);
  not ginst867 (R1117_U465, R1117_U159);
  nand ginst868 (R1117_U466, R1117_U351, R1117_U465);
  nand ginst869 (R1117_U467, R1117_U159, R1117_U190);
  nand ginst870 (R1117_U468, R1117_U45, U3468);
  nand ginst871 (R1117_U469, R1117_U191, U3075);
  not ginst872 (R1117_U47, U3068);
  not ginst873 (R1117_U470, R1117_U160);
  nand ginst874 (R1117_U471, R1117_U219, R1117_U470);
  nand ginst875 (R1117_U472, R1117_U160, R1117_U192);
  nand ginst876 (R1117_U473, R1117_U71, U3504);
  nand ginst877 (R1117_U474, R1117_U74, U3078);
  not ginst878 (R1117_U475, R1117_U161);
  nand ginst879 (R1117_U476, R1117_U381, R1117_U475);
  nand ginst880 (R1117_U477, R1117_U161, R1117_U193);
  nand ginst881 (R1117_U478, R1117_U75, U3502);
  nand ginst882 (R1117_U479, R1117_U96, U3079);
  not ginst883 (R1117_U48, U3064);
  not ginst884 (R1117_U480, R1117_U162);
  nand ginst885 (R1117_U481, R1117_U284, R1117_U480);
  nand ginst886 (R1117_U482, R1117_U162, R1117_U194);
  nand ginst887 (R1117_U483, R1117_U76, U3500);
  nand ginst888 (R1117_U484, R1117_U77, U3066);
  not ginst889 (R1117_U485, R1117_U163);
  nand ginst890 (R1117_U486, R1117_U281, R1117_U485);
  nand ginst891 (R1117_U487, R1117_U163, R1117_U195);
  nand ginst892 (R1117_U488, R1117_U91, U3498);
  nand ginst893 (R1117_U489, R1117_U78, U3070);
  not ginst894 (R1117_U49, U3057);
  nand ginst895 (R1117_U490, R1117_U488, R1117_U489);
  nand ginst896 (R1117_U491, R1117_U92, U3496);
  nand ginst897 (R1117_U492, R1117_U79, U3071);
  nand ginst898 (R1117_U493, R1117_U106, R1117_U324);
  nand ginst899 (R1117_U494, R1117_U196, R1117_U316);
  nand ginst900 (R1117_U495, R1117_U93, U3494);
  nand ginst901 (R1117_U496, R1117_U80, U3076);
  nand ginst902 (R1117_U497, R1117_U198, R1117_U325);
  nand ginst903 (R1117_U498, R1117_U197, R1117_U367);
  nand ginst904 (R1117_U499, R1117_U81, U3492);
  nand ginst905 (R1117_U50, R1117_U37, U3057);
  nand ginst906 (R1117_U500, R1117_U82, U3077);
  not ginst907 (R1117_U501, R1117_U166);
  nand ginst908 (R1117_U502, R1117_U365, R1117_U501);
  nand ginst909 (R1117_U503, R1117_U166, R1117_U199);
  nand ginst910 (R1117_U504, R1117_U89, U3490);
  nand ginst911 (R1117_U505, R1117_U83, U3069);
  not ginst912 (R1117_U506, R1117_U167);
  nand ginst913 (R1117_U507, R1117_U363, R1117_U506);
  nand ginst914 (R1117_U508, R1117_U167, R1117_U200);
  nand ginst915 (R1117_U509, R1117_U84, U3488);
  nand ginst916 (R1117_U51, R1117_U230, R1117_U232);
  nand ginst917 (R1117_U510, R1117_U86, U3060);
  nand ginst918 (R1117_U511, R1117_U509, R1117_U510);
  nand ginst919 (R1117_U512, R1117_U85, U3486);
  nand ginst920 (R1117_U513, R1117_U87, U3059);
  nand ginst921 (R1117_U514, R1117_U107, R1117_U333);
  nand ginst922 (R1117_U515, R1117_U201, R1117_U361);
  not ginst923 (R1117_U52, U3484);
  not ginst924 (R1117_U53, U3080);
  nand ginst925 (R1117_U54, R1117_U233, R1117_U51);
  nand ginst926 (R1117_U55, R1117_U248, R1117_U50);
  nand ginst927 (R1117_U56, R1117_U204, R1117_U220, R1117_U335);
  not ginst928 (R1117_U57, U4029);
  not ginst929 (R1117_U58, U3054);
  nand ginst930 (R1117_U59, R1117_U99, U3054);
  and ginst931 (R1117_U6, R1117_U227, R1117_U228);
  not ginst932 (R1117_U60, U3050);
  not ginst933 (R1117_U61, U3062);
  not ginst934 (R1117_U62, U4033);
  not ginst935 (R1117_U63, U3063);
  not ginst936 (R1117_U64, U3058);
  not ginst937 (R1117_U65, U3072);
  not ginst938 (R1117_U66, U4034);
  not ginst939 (R1117_U67, U4035);
  nand ginst940 (R1117_U68, R1117_U69, U3072);
  not ginst941 (R1117_U69, U4036);
  and ginst942 (R1117_U7, R1117_U208, R1117_U261);
  not ginst943 (R1117_U70, U3073);
  not ginst944 (R1117_U71, U3078);
  not ginst945 (R1117_U72, U4037);
  nand ginst946 (R1117_U73, R1117_U74, U3078);
  not ginst947 (R1117_U74, U3504);
  not ginst948 (R1117_U75, U3079);
  not ginst949 (R1117_U76, U3066);
  not ginst950 (R1117_U77, U3500);
  not ginst951 (R1117_U78, U3498);
  not ginst952 (R1117_U79, U3496);
  and ginst953 (R1117_U8, R1117_U262, R1117_U263);
  not ginst954 (R1117_U80, U3494);
  not ginst955 (R1117_U81, U3077);
  not ginst956 (R1117_U82, U3492);
  not ginst957 (R1117_U83, U3490);
  not ginst958 (R1117_U84, U3060);
  not ginst959 (R1117_U85, U3059);
  not ginst960 (R1117_U86, U3488);
  not ginst961 (R1117_U87, U3486);
  nand ginst962 (R1117_U88, R1117_U52, U3080);
  not ginst963 (R1117_U89, U3069);
  and ginst964 (R1117_U9, R1117_U209, R1117_U272);
  nand ginst965 (R1117_U90, R1117_U268, R1117_U339);
  not ginst966 (R1117_U91, U3070);
  not ginst967 (R1117_U92, U3071);
  not ginst968 (R1117_U93, U3076);
  nand ginst969 (R1117_U94, R1117_U80, U3076);
  nand ginst970 (R1117_U95, R1117_U276, R1117_U278);
  not ginst971 (R1117_U96, U3502);
  not ginst972 (R1117_U97, U4032);
  not ginst973 (R1117_U98, U3055);
  not ginst974 (R1117_U99, U4031);
  and ginst975 (R1138_U10, R1138_U281, R1138_U282);
  nand ginst976 (R1138_U100, R1138_U314, R1138_U60);
  nand ginst977 (R1138_U101, R1138_U294, R1138_U385);
  nand ginst978 (R1138_U102, R1138_U277, R1138_U278);
  not ginst979 (R1138_U103, U3073);
  nand ginst980 (R1138_U104, R1138_U323, R1138_U84);
  nand ginst981 (R1138_U105, R1138_U271, R1138_U382, R1138_U383);
  nand ginst982 (R1138_U106, R1138_U345, R1138_U72);
  nand ginst983 (R1138_U107, R1138_U483, R1138_U484);
  nand ginst984 (R1138_U108, R1138_U530, R1138_U531);
  nand ginst985 (R1138_U109, R1138_U401, R1138_U402);
  and ginst986 (R1138_U11, R1138_U10, R1138_U283);
  nand ginst987 (R1138_U110, R1138_U406, R1138_U407);
  nand ginst988 (R1138_U111, R1138_U413, R1138_U414);
  nand ginst989 (R1138_U112, R1138_U420, R1138_U421);
  nand ginst990 (R1138_U113, R1138_U425, R1138_U426);
  nand ginst991 (R1138_U114, R1138_U434, R1138_U435);
  nand ginst992 (R1138_U115, R1138_U441, R1138_U442);
  nand ginst993 (R1138_U116, R1138_U448, R1138_U449);
  nand ginst994 (R1138_U117, R1138_U455, R1138_U456);
  nand ginst995 (R1138_U118, R1138_U460, R1138_U461);
  nand ginst996 (R1138_U119, R1138_U467, R1138_U468);
  and ginst997 (R1138_U12, R1138_U217, R1138_U7);
  nand ginst998 (R1138_U120, R1138_U474, R1138_U475);
  nand ginst999 (R1138_U121, R1138_U488, R1138_U489);
  nand ginst1000 (R1138_U122, R1138_U493, R1138_U494);
  nand ginst1001 (R1138_U123, R1138_U500, R1138_U501);
  nand ginst1002 (R1138_U124, R1138_U507, R1138_U508);
  nand ginst1003 (R1138_U125, R1138_U514, R1138_U515);
  nand ginst1004 (R1138_U126, R1138_U521, R1138_U522);
  nand ginst1005 (R1138_U127, R1138_U526, R1138_U527);
  and ginst1006 (R1138_U128, R1138_U129, R1138_U197);
  and ginst1007 (R1138_U129, U3065, U3470);
  and ginst1008 (R1138_U13, R1138_U262, R1138_U8);
  and ginst1009 (R1138_U130, U3061, U3472);
  and ginst1010 (R1138_U131, U3074, U3464);
  and ginst1011 (R1138_U132, R1138_U203, R1138_U204, R1138_U206);
  and ginst1012 (R1138_U133, R1138_U207, R1138_U373, R1138_U374);
  and ginst1013 (R1138_U134, R1138_U408, R1138_U409, R1138_U43);
  and ginst1014 (R1138_U135, R1138_U225, R1138_U6);
  and ginst1015 (R1138_U136, R1138_U231, R1138_U233);
  and ginst1016 (R1138_U137, R1138_U34, R1138_U415, R1138_U416);
  and ginst1017 (R1138_U138, R1138_U239, R1138_U4);
  and ginst1018 (R1138_U139, R1138_U198, R1138_U247);
  and ginst1019 (R1138_U14, R1138_U11, R1138_U292);
  and ginst1020 (R1138_U140, R1138_U188, R1138_U252);
  and ginst1021 (R1138_U141, R1138_U12, R1138_U6);
  and ginst1022 (R1138_U142, R1138_U255, R1138_U378);
  and ginst1023 (R1138_U143, R1138_U15, R1138_U270);
  and ginst1024 (R1138_U144, R1138_U189, R1138_U260);
  and ginst1025 (R1138_U145, R1138_U16, R1138_U296);
  and ginst1026 (R1138_U146, R1138_U297, R1138_U389);
  and ginst1027 (R1138_U147, R1138_U185, R1138_U309);
  and ginst1028 (R1138_U148, R1138_U310, R1138_U393, R1138_U395);
  and ginst1029 (R1138_U149, R1138_U17, R1138_U185);
  and ginst1030 (R1138_U15, R1138_U13, R1138_U267);
  and ginst1031 (R1138_U150, R1138_U304, R1138_U97);
  and ginst1032 (R1138_U151, R1138_U190, R1138_U450, R1138_U451);
  and ginst1033 (R1138_U152, R1138_U185, R1138_U320);
  and ginst1034 (R1138_U153, R1138_U176, R1138_U288);
  and ginst1035 (R1138_U154, R1138_U481, R1138_U482, R1138_U80);
  and ginst1036 (R1138_U155, R1138_U10, R1138_U333);
  and ginst1037 (R1138_U156, R1138_U495, R1138_U496, R1138_U90);
  and ginst1038 (R1138_U157, R1138_U342, R1138_U9);
  and ginst1039 (R1138_U158, R1138_U189, R1138_U516, R1138_U517);
  and ginst1040 (R1138_U159, R1138_U351, R1138_U8);
  and ginst1041 (R1138_U16, R1138_U14, R1138_U9);
  and ginst1042 (R1138_U160, R1138_U188, R1138_U528, R1138_U529);
  and ginst1043 (R1138_U161, R1138_U358, R1138_U7);
  nand ginst1044 (R1138_U162, R1138_U215, R1138_U375);
  nand ginst1045 (R1138_U163, R1138_U230, R1138_U242);
  not ginst1046 (R1138_U164, U3052);
  not ginst1047 (R1138_U165, U4040);
  and ginst1048 (R1138_U166, R1138_U429, R1138_U430);
  nand ginst1049 (R1138_U167, R1138_U186, R1138_U312, R1138_U372);
  and ginst1050 (R1138_U168, R1138_U436, R1138_U437);
  nand ginst1051 (R1138_U169, R1138_U148, R1138_U394);
  and ginst1052 (R1138_U17, R1138_U299, R1138_U305);
  and ginst1053 (R1138_U170, R1138_U443, R1138_U444);
  nand ginst1054 (R1138_U171, R1138_U150, R1138_U307);
  nand ginst1055 (R1138_U172, R1138_U300, R1138_U301);
  and ginst1056 (R1138_U173, R1138_U462, R1138_U463);
  and ginst1057 (R1138_U174, R1138_U469, R1138_U470);
  nand ginst1058 (R1138_U175, R1138_U384, R1138_U386);
  and ginst1059 (R1138_U176, R1138_U476, R1138_U477);
  nand ginst1060 (R1138_U177, U3074, U3464);
  nand ginst1061 (R1138_U178, R1138_U335, R1138_U36);
  nand ginst1062 (R1138_U179, R1138_U279, R1138_U376);
  and ginst1063 (R1138_U18, R1138_U356, R1138_U359);
  and ginst1064 (R1138_U180, R1138_U502, R1138_U503);
  nand ginst1065 (R1138_U181, R1138_U379, R1138_U77);
  and ginst1066 (R1138_U182, R1138_U509, R1138_U510);
  nand ginst1067 (R1138_U183, R1138_U264, R1138_U265);
  nand ginst1068 (R1138_U184, R1138_U142, R1138_U377);
  nand ginst1069 (R1138_U185, R1138_U390, R1138_U391);
  nand ginst1070 (R1138_U186, R1138_U169, U3051);
  not ginst1071 (R1138_U187, R1138_U34);
  nand ginst1072 (R1138_U188, U3080, U3484);
  nand ginst1073 (R1138_U189, U3069, U3490);
  and ginst1074 (R1138_U19, R1138_U349, R1138_U352);
  nand ginst1075 (R1138_U190, U3055, U4032);
  not ginst1076 (R1138_U191, R1138_U72);
  not ginst1077 (R1138_U192, R1138_U84);
  not ginst1078 (R1138_U193, R1138_U60);
  not ginst1079 (R1138_U194, R1138_U65);
  or ginst1080 (R1138_U195, U3064, U3476);
  or ginst1081 (R1138_U196, U3057, U3474);
  or ginst1082 (R1138_U197, U3061, U3472);
  or ginst1083 (R1138_U198, U3065, U3470);
  not ginst1084 (R1138_U199, R1138_U177);
  and ginst1085 (R1138_U20, R1138_U340, R1138_U343);
  or ginst1086 (R1138_U200, U3075, U3468);
  not ginst1087 (R1138_U201, R1138_U39);
  not ginst1088 (R1138_U202, R1138_U36);
  nand ginst1089 (R1138_U203, R1138_U128, R1138_U4);
  nand ginst1090 (R1138_U204, R1138_U130, R1138_U4);
  nand ginst1091 (R1138_U205, R1138_U34, R1138_U35);
  nand ginst1092 (R1138_U206, R1138_U205, U3064);
  nand ginst1093 (R1138_U207, R1138_U187, U3476);
  not ginst1094 (R1138_U208, R1138_U51);
  or ginst1095 (R1138_U209, U3067, U3480);
  and ginst1096 (R1138_U21, R1138_U331, R1138_U334);
  or ginst1097 (R1138_U210, U3068, U3478);
  not ginst1098 (R1138_U211, R1138_U43);
  nand ginst1099 (R1138_U212, R1138_U43, R1138_U44);
  nand ginst1100 (R1138_U213, R1138_U212, U3067);
  nand ginst1101 (R1138_U214, R1138_U211, U3480);
  nand ginst1102 (R1138_U215, R1138_U51, R1138_U6);
  not ginst1103 (R1138_U216, R1138_U162);
  or ginst1104 (R1138_U217, U3081, U3482);
  nand ginst1105 (R1138_U218, R1138_U162, R1138_U217);
  not ginst1106 (R1138_U219, R1138_U50);
  and ginst1107 (R1138_U22, R1138_U326, R1138_U328);
  or ginst1108 (R1138_U220, U3080, U3484);
  or ginst1109 (R1138_U221, U3068, U3478);
  nand ginst1110 (R1138_U222, R1138_U221, R1138_U51);
  nand ginst1111 (R1138_U223, R1138_U134, R1138_U222);
  nand ginst1112 (R1138_U224, R1138_U208, R1138_U43);
  nand ginst1113 (R1138_U225, U3067, U3480);
  nand ginst1114 (R1138_U226, R1138_U135, R1138_U224);
  or ginst1115 (R1138_U227, U3068, U3478);
  nand ginst1116 (R1138_U228, R1138_U198, R1138_U202);
  nand ginst1117 (R1138_U229, U3065, U3470);
  and ginst1118 (R1138_U23, R1138_U318, R1138_U321);
  not ginst1119 (R1138_U230, R1138_U53);
  nand ginst1120 (R1138_U231, R1138_U201, R1138_U5);
  nand ginst1121 (R1138_U232, R1138_U197, R1138_U53);
  nand ginst1122 (R1138_U233, U3061, U3472);
  not ginst1123 (R1138_U234, R1138_U52);
  or ginst1124 (R1138_U235, U3057, U3474);
  nand ginst1125 (R1138_U236, R1138_U235, R1138_U52);
  nand ginst1126 (R1138_U237, R1138_U137, R1138_U236);
  nand ginst1127 (R1138_U238, R1138_U234, R1138_U34);
  nand ginst1128 (R1138_U239, U3064, U3476);
  and ginst1129 (R1138_U24, R1138_U245, R1138_U248);
  nand ginst1130 (R1138_U240, R1138_U138, R1138_U238);
  or ginst1131 (R1138_U241, U3057, U3474);
  nand ginst1132 (R1138_U242, R1138_U198, R1138_U201);
  not ginst1133 (R1138_U243, R1138_U163);
  nand ginst1134 (R1138_U244, U3061, U3472);
  nand ginst1135 (R1138_U245, R1138_U36, R1138_U39, R1138_U427, R1138_U428);
  nand ginst1136 (R1138_U246, R1138_U36, R1138_U39);
  nand ginst1137 (R1138_U247, U3065, U3470);
  nand ginst1138 (R1138_U248, R1138_U139, R1138_U246);
  or ginst1139 (R1138_U249, U3080, U3484);
  and ginst1140 (R1138_U25, R1138_U237, R1138_U240);
  or ginst1141 (R1138_U250, U3059, U3486);
  nand ginst1142 (R1138_U251, R1138_U194, R1138_U7);
  nand ginst1143 (R1138_U252, U3059, U3486);
  nand ginst1144 (R1138_U253, R1138_U140, R1138_U251);
  or ginst1145 (R1138_U254, U3059, U3486);
  nand ginst1146 (R1138_U255, R1138_U253, R1138_U254);
  not ginst1147 (R1138_U256, R1138_U184);
  or ginst1148 (R1138_U257, U3077, U3492);
  or ginst1149 (R1138_U258, U3069, U3490);
  nand ginst1150 (R1138_U259, R1138_U191, R1138_U8);
  and ginst1151 (R1138_U26, R1138_U223, R1138_U226);
  nand ginst1152 (R1138_U260, U3077, U3492);
  nand ginst1153 (R1138_U261, R1138_U144, R1138_U259);
  or ginst1154 (R1138_U262, U3060, U3488);
  or ginst1155 (R1138_U263, U3077, U3492);
  nand ginst1156 (R1138_U264, R1138_U13, R1138_U184);
  nand ginst1157 (R1138_U265, R1138_U261, R1138_U263);
  not ginst1158 (R1138_U266, R1138_U183);
  or ginst1159 (R1138_U267, U3076, U3494);
  nand ginst1160 (R1138_U268, U3076, U3494);
  not ginst1161 (R1138_U269, R1138_U181);
  not ginst1162 (R1138_U27, U3470);
  or ginst1163 (R1138_U270, U3071, U3496);
  nand ginst1164 (R1138_U271, U3071, U3496);
  not ginst1165 (R1138_U272, R1138_U105);
  or ginst1166 (R1138_U273, U3066, U3500);
  or ginst1167 (R1138_U274, U3070, U3498);
  not ginst1168 (R1138_U275, R1138_U90);
  nand ginst1169 (R1138_U276, R1138_U90, R1138_U91);
  nand ginst1170 (R1138_U277, R1138_U276, U3066);
  nand ginst1171 (R1138_U278, R1138_U275, U3500);
  nand ginst1172 (R1138_U279, R1138_U105, R1138_U9);
  not ginst1173 (R1138_U28, U3065);
  not ginst1174 (R1138_U280, R1138_U179);
  or ginst1175 (R1138_U281, U3073, U4037);
  or ginst1176 (R1138_U282, U3078, U3504);
  or ginst1177 (R1138_U283, U3072, U4036);
  not ginst1178 (R1138_U284, R1138_U80);
  nand ginst1179 (R1138_U285, R1138_U284, U4037);
  nand ginst1180 (R1138_U286, R1138_U103, R1138_U285);
  nand ginst1181 (R1138_U287, R1138_U80, R1138_U81);
  nand ginst1182 (R1138_U288, R1138_U286, R1138_U287);
  nand ginst1183 (R1138_U289, R1138_U11, R1138_U192);
  not ginst1184 (R1138_U29, U3472);
  nand ginst1185 (R1138_U290, U3072, U4036);
  nand ginst1186 (R1138_U291, R1138_U288, R1138_U289, R1138_U290);
  or ginst1187 (R1138_U292, U3079, U3502);
  or ginst1188 (R1138_U293, U3072, U4036);
  nand ginst1189 (R1138_U294, R1138_U291, R1138_U293);
  not ginst1190 (R1138_U295, R1138_U175);
  or ginst1191 (R1138_U296, U3058, U4035);
  nand ginst1192 (R1138_U297, U3058, U4035);
  not ginst1193 (R1138_U298, R1138_U94);
  or ginst1194 (R1138_U299, U3063, U4034);
  not ginst1195 (R1138_U30, U3061);
  nand ginst1196 (R1138_U300, R1138_U299, R1138_U94);
  nand ginst1197 (R1138_U301, U3063, U4034);
  not ginst1198 (R1138_U302, R1138_U172);
  or ginst1199 (R1138_U303, U3055, U4032);
  nand ginst1200 (R1138_U304, R1138_U185, R1138_U193);
  or ginst1201 (R1138_U305, U3062, U4033);
  or ginst1202 (R1138_U306, U3054, U4031);
  nand ginst1203 (R1138_U307, R1138_U149, R1138_U392);
  not ginst1204 (R1138_U308, R1138_U171);
  or ginst1205 (R1138_U309, U3050, U4030);
  not ginst1206 (R1138_U31, U3474);
  nand ginst1207 (R1138_U310, U3050, U4030);
  not ginst1208 (R1138_U311, R1138_U169);
  nand ginst1209 (R1138_U312, R1138_U169, U4029);
  not ginst1210 (R1138_U313, R1138_U167);
  nand ginst1211 (R1138_U314, R1138_U172, R1138_U305);
  not ginst1212 (R1138_U315, R1138_U100);
  or ginst1213 (R1138_U316, U3055, U4032);
  nand ginst1214 (R1138_U317, R1138_U100, R1138_U316);
  nand ginst1215 (R1138_U318, R1138_U151, R1138_U317);
  nand ginst1216 (R1138_U319, R1138_U190, R1138_U315);
  not ginst1217 (R1138_U32, U3057);
  nand ginst1218 (R1138_U320, U3054, U4031);
  nand ginst1219 (R1138_U321, R1138_U152, R1138_U319);
  or ginst1220 (R1138_U322, U3055, U4032);
  nand ginst1221 (R1138_U323, R1138_U179, R1138_U292);
  not ginst1222 (R1138_U324, R1138_U104);
  nand ginst1223 (R1138_U325, R1138_U10, R1138_U104);
  nand ginst1224 (R1138_U326, R1138_U153, R1138_U325);
  nand ginst1225 (R1138_U327, R1138_U288, R1138_U325);
  nand ginst1226 (R1138_U328, R1138_U327, R1138_U480);
  or ginst1227 (R1138_U329, U3078, U3504);
  not ginst1228 (R1138_U33, U3064);
  nand ginst1229 (R1138_U330, R1138_U104, R1138_U329);
  nand ginst1230 (R1138_U331, R1138_U154, R1138_U330);
  nand ginst1231 (R1138_U332, R1138_U324, R1138_U80);
  nand ginst1232 (R1138_U333, U3073, U4037);
  nand ginst1233 (R1138_U334, R1138_U155, R1138_U332);
  or ginst1234 (R1138_U335, U3075, U3468);
  not ginst1235 (R1138_U336, R1138_U178);
  or ginst1236 (R1138_U337, U3078, U3504);
  or ginst1237 (R1138_U338, U3070, U3498);
  nand ginst1238 (R1138_U339, R1138_U105, R1138_U338);
  nand ginst1239 (R1138_U34, U3057, U3474);
  nand ginst1240 (R1138_U340, R1138_U156, R1138_U339);
  nand ginst1241 (R1138_U341, R1138_U272, R1138_U90);
  nand ginst1242 (R1138_U342, U3066, U3500);
  nand ginst1243 (R1138_U343, R1138_U157, R1138_U341);
  or ginst1244 (R1138_U344, U3070, U3498);
  nand ginst1245 (R1138_U345, R1138_U184, R1138_U262);
  not ginst1246 (R1138_U346, R1138_U106);
  or ginst1247 (R1138_U347, U3069, U3490);
  nand ginst1248 (R1138_U348, R1138_U106, R1138_U347);
  nand ginst1249 (R1138_U349, R1138_U158, R1138_U348);
  not ginst1250 (R1138_U35, U3476);
  nand ginst1251 (R1138_U350, R1138_U189, R1138_U346);
  nand ginst1252 (R1138_U351, U3077, U3492);
  nand ginst1253 (R1138_U352, R1138_U159, R1138_U350);
  or ginst1254 (R1138_U353, U3069, U3490);
  or ginst1255 (R1138_U354, U3080, U3484);
  nand ginst1256 (R1138_U355, R1138_U354, R1138_U50);
  nand ginst1257 (R1138_U356, R1138_U160, R1138_U355);
  nand ginst1258 (R1138_U357, R1138_U188, R1138_U219);
  nand ginst1259 (R1138_U358, U3059, U3486);
  nand ginst1260 (R1138_U359, R1138_U161, R1138_U357);
  nand ginst1261 (R1138_U36, U3075, U3468);
  nand ginst1262 (R1138_U360, R1138_U188, R1138_U220);
  nand ginst1263 (R1138_U361, R1138_U217, R1138_U65);
  nand ginst1264 (R1138_U362, R1138_U227, R1138_U43);
  nand ginst1265 (R1138_U363, R1138_U241, R1138_U34);
  nand ginst1266 (R1138_U364, R1138_U197, R1138_U244);
  nand ginst1267 (R1138_U365, R1138_U190, R1138_U322);
  nand ginst1268 (R1138_U366, R1138_U305, R1138_U60);
  nand ginst1269 (R1138_U367, R1138_U337, R1138_U80);
  nand ginst1270 (R1138_U368, R1138_U292, R1138_U84);
  nand ginst1271 (R1138_U369, R1138_U344, R1138_U90);
  not ginst1272 (R1138_U37, U3464);
  nand ginst1273 (R1138_U370, R1138_U189, R1138_U353);
  nand ginst1274 (R1138_U371, R1138_U262, R1138_U72);
  nand ginst1275 (R1138_U372, U3051, U4029);
  nand ginst1276 (R1138_U373, R1138_U202, R1138_U4, R1138_U5);
  nand ginst1277 (R1138_U374, R1138_U201, R1138_U4, R1138_U5);
  not ginst1278 (R1138_U375, R1138_U45);
  not ginst1279 (R1138_U376, R1138_U102);
  nand ginst1280 (R1138_U377, R1138_U141, R1138_U51);
  nand ginst1281 (R1138_U378, R1138_U12, R1138_U45);
  nand ginst1282 (R1138_U379, R1138_U15, R1138_U184);
  not ginst1283 (R1138_U38, U3074);
  nand ginst1284 (R1138_U380, R1138_U265, R1138_U268);
  not ginst1285 (R1138_U381, R1138_U77);
  nand ginst1286 (R1138_U382, R1138_U143, R1138_U184);
  nand ginst1287 (R1138_U383, R1138_U270, R1138_U381);
  nand ginst1288 (R1138_U384, R1138_U105, R1138_U16);
  nand ginst1289 (R1138_U385, R1138_U102, R1138_U14);
  not ginst1290 (R1138_U386, R1138_U101);
  not ginst1291 (R1138_U387, R1138_U97);
  nand ginst1292 (R1138_U388, R1138_U105, R1138_U145);
  nand ginst1293 (R1138_U389, R1138_U101, R1138_U296);
  nand ginst1294 (R1138_U39, R1138_U131, R1138_U200);
  nand ginst1295 (R1138_U390, R1138_U303, U3054);
  nand ginst1296 (R1138_U391, R1138_U303, U4031);
  nand ginst1297 (R1138_U392, R1138_U298, R1138_U301);
  nand ginst1298 (R1138_U393, R1138_U185, R1138_U193, R1138_U309);
  nand ginst1299 (R1138_U394, R1138_U147, R1138_U17, R1138_U392);
  nand ginst1300 (R1138_U395, R1138_U309, R1138_U387);
  nand ginst1301 (R1138_U396, R1138_U190, R1138_U57);
  nand ginst1302 (R1138_U397, R1138_U190, R1138_U56);
  nand ginst1303 (R1138_U398, R1138_U49, U3080);
  nand ginst1304 (R1138_U399, R1138_U48, U3484);
  and ginst1305 (R1138_U4, R1138_U195, R1138_U196);
  not ginst1306 (R1138_U40, U3478);
  nand ginst1307 (R1138_U400, R1138_U398, R1138_U399);
  nand ginst1308 (R1138_U401, R1138_U360, R1138_U50);
  nand ginst1309 (R1138_U402, R1138_U219, R1138_U400);
  nand ginst1310 (R1138_U403, R1138_U46, U3081);
  nand ginst1311 (R1138_U404, R1138_U47, U3482);
  nand ginst1312 (R1138_U405, R1138_U403, R1138_U404);
  nand ginst1313 (R1138_U406, R1138_U162, R1138_U361);
  nand ginst1314 (R1138_U407, R1138_U216, R1138_U405);
  nand ginst1315 (R1138_U408, R1138_U44, U3067);
  nand ginst1316 (R1138_U409, R1138_U42, U3480);
  not ginst1317 (R1138_U41, U3068);
  nand ginst1318 (R1138_U410, R1138_U40, U3068);
  nand ginst1319 (R1138_U411, R1138_U41, U3478);
  nand ginst1320 (R1138_U412, R1138_U410, R1138_U411);
  nand ginst1321 (R1138_U413, R1138_U362, R1138_U51);
  nand ginst1322 (R1138_U414, R1138_U208, R1138_U412);
  nand ginst1323 (R1138_U415, R1138_U35, U3064);
  nand ginst1324 (R1138_U416, R1138_U33, U3476);
  nand ginst1325 (R1138_U417, R1138_U31, U3057);
  nand ginst1326 (R1138_U418, R1138_U32, U3474);
  nand ginst1327 (R1138_U419, R1138_U417, R1138_U418);
  not ginst1328 (R1138_U42, U3067);
  nand ginst1329 (R1138_U420, R1138_U363, R1138_U52);
  nand ginst1330 (R1138_U421, R1138_U234, R1138_U419);
  nand ginst1331 (R1138_U422, R1138_U29, U3061);
  nand ginst1332 (R1138_U423, R1138_U30, U3472);
  nand ginst1333 (R1138_U424, R1138_U422, R1138_U423);
  nand ginst1334 (R1138_U425, R1138_U163, R1138_U364);
  nand ginst1335 (R1138_U426, R1138_U243, R1138_U424);
  nand ginst1336 (R1138_U427, R1138_U27, U3065);
  nand ginst1337 (R1138_U428, R1138_U28, U3470);
  nand ginst1338 (R1138_U429, R1138_U165, U3052);
  nand ginst1339 (R1138_U43, U3068, U3478);
  nand ginst1340 (R1138_U430, R1138_U164, U4040);
  nand ginst1341 (R1138_U431, R1138_U165, U3052);
  nand ginst1342 (R1138_U432, R1138_U164, U4040);
  nand ginst1343 (R1138_U433, R1138_U431, R1138_U432);
  nand ginst1344 (R1138_U434, R1138_U166, R1138_U167);
  nand ginst1345 (R1138_U435, R1138_U313, R1138_U433);
  nand ginst1346 (R1138_U436, R1138_U99, U3051);
  nand ginst1347 (R1138_U437, R1138_U98, U4029);
  nand ginst1348 (R1138_U438, R1138_U99, U3051);
  nand ginst1349 (R1138_U439, R1138_U98, U4029);
  not ginst1350 (R1138_U44, U3480);
  nand ginst1351 (R1138_U440, R1138_U438, R1138_U439);
  nand ginst1352 (R1138_U441, R1138_U168, R1138_U169);
  nand ginst1353 (R1138_U442, R1138_U311, R1138_U440);
  nand ginst1354 (R1138_U443, R1138_U54, U3050);
  nand ginst1355 (R1138_U444, R1138_U55, U4030);
  nand ginst1356 (R1138_U445, R1138_U54, U3050);
  nand ginst1357 (R1138_U446, R1138_U55, U4030);
  nand ginst1358 (R1138_U447, R1138_U445, R1138_U446);
  nand ginst1359 (R1138_U448, R1138_U170, R1138_U171);
  nand ginst1360 (R1138_U449, R1138_U308, R1138_U447);
  nand ginst1361 (R1138_U45, R1138_U213, R1138_U214);
  nand ginst1362 (R1138_U450, R1138_U57, U3054);
  nand ginst1363 (R1138_U451, R1138_U56, U4031);
  nand ginst1364 (R1138_U452, R1138_U95, U3055);
  nand ginst1365 (R1138_U453, R1138_U96, U4032);
  nand ginst1366 (R1138_U454, R1138_U452, R1138_U453);
  nand ginst1367 (R1138_U455, R1138_U100, R1138_U365);
  nand ginst1368 (R1138_U456, R1138_U315, R1138_U454);
  nand ginst1369 (R1138_U457, R1138_U58, U3062);
  nand ginst1370 (R1138_U458, R1138_U59, U4033);
  nand ginst1371 (R1138_U459, R1138_U457, R1138_U458);
  not ginst1372 (R1138_U46, U3482);
  nand ginst1373 (R1138_U460, R1138_U172, R1138_U366);
  nand ginst1374 (R1138_U461, R1138_U302, R1138_U459);
  nand ginst1375 (R1138_U462, R1138_U92, U3063);
  nand ginst1376 (R1138_U463, R1138_U93, U4034);
  nand ginst1377 (R1138_U464, R1138_U92, U3063);
  nand ginst1378 (R1138_U465, R1138_U93, U4034);
  nand ginst1379 (R1138_U466, R1138_U464, R1138_U465);
  nand ginst1380 (R1138_U467, R1138_U173, R1138_U94);
  nand ginst1381 (R1138_U468, R1138_U298, R1138_U466);
  nand ginst1382 (R1138_U469, R1138_U61, U3058);
  not ginst1383 (R1138_U47, U3081);
  nand ginst1384 (R1138_U470, R1138_U62, U4035);
  nand ginst1385 (R1138_U471, R1138_U61, U3058);
  nand ginst1386 (R1138_U472, R1138_U62, U4035);
  nand ginst1387 (R1138_U473, R1138_U471, R1138_U472);
  nand ginst1388 (R1138_U474, R1138_U174, R1138_U175);
  nand ginst1389 (R1138_U475, R1138_U295, R1138_U473);
  nand ginst1390 (R1138_U476, R1138_U85, U3072);
  nand ginst1391 (R1138_U477, R1138_U86, U4036);
  nand ginst1392 (R1138_U478, R1138_U85, U3072);
  nand ginst1393 (R1138_U479, R1138_U86, U4036);
  not ginst1394 (R1138_U48, U3080);
  nand ginst1395 (R1138_U480, R1138_U478, R1138_U479);
  nand ginst1396 (R1138_U481, R1138_U81, U3073);
  nand ginst1397 (R1138_U482, R1138_U103, U4037);
  nand ginst1398 (R1138_U483, R1138_U178, R1138_U199);
  nand ginst1399 (R1138_U484, R1138_U177, R1138_U336);
  nand ginst1400 (R1138_U485, R1138_U78, U3078);
  nand ginst1401 (R1138_U486, R1138_U79, U3504);
  nand ginst1402 (R1138_U487, R1138_U485, R1138_U486);
  nand ginst1403 (R1138_U488, R1138_U104, R1138_U367);
  nand ginst1404 (R1138_U489, R1138_U324, R1138_U487);
  not ginst1405 (R1138_U49, U3484);
  nand ginst1406 (R1138_U490, R1138_U82, U3079);
  nand ginst1407 (R1138_U491, R1138_U83, U3502);
  nand ginst1408 (R1138_U492, R1138_U490, R1138_U491);
  nand ginst1409 (R1138_U493, R1138_U179, R1138_U368);
  nand ginst1410 (R1138_U494, R1138_U280, R1138_U492);
  nand ginst1411 (R1138_U495, R1138_U91, U3066);
  nand ginst1412 (R1138_U496, R1138_U89, U3500);
  nand ginst1413 (R1138_U497, R1138_U87, U3070);
  nand ginst1414 (R1138_U498, R1138_U88, U3498);
  nand ginst1415 (R1138_U499, R1138_U497, R1138_U498);
  and ginst1416 (R1138_U5, R1138_U197, R1138_U198);
  nand ginst1417 (R1138_U50, R1138_U218, R1138_U65);
  nand ginst1418 (R1138_U500, R1138_U105, R1138_U369);
  nand ginst1419 (R1138_U501, R1138_U272, R1138_U499);
  nand ginst1420 (R1138_U502, R1138_U63, U3071);
  nand ginst1421 (R1138_U503, R1138_U64, U3496);
  nand ginst1422 (R1138_U504, R1138_U63, U3071);
  nand ginst1423 (R1138_U505, R1138_U64, U3496);
  nand ginst1424 (R1138_U506, R1138_U504, R1138_U505);
  nand ginst1425 (R1138_U507, R1138_U180, R1138_U181);
  nand ginst1426 (R1138_U508, R1138_U269, R1138_U506);
  nand ginst1427 (R1138_U509, R1138_U75, U3076);
  nand ginst1428 (R1138_U51, R1138_U132, R1138_U133);
  nand ginst1429 (R1138_U510, R1138_U76, U3494);
  nand ginst1430 (R1138_U511, R1138_U75, U3076);
  nand ginst1431 (R1138_U512, R1138_U76, U3494);
  nand ginst1432 (R1138_U513, R1138_U511, R1138_U512);
  nand ginst1433 (R1138_U514, R1138_U182, R1138_U183);
  nand ginst1434 (R1138_U515, R1138_U266, R1138_U513);
  nand ginst1435 (R1138_U516, R1138_U73, U3077);
  nand ginst1436 (R1138_U517, R1138_U74, U3492);
  nand ginst1437 (R1138_U518, R1138_U68, U3069);
  nand ginst1438 (R1138_U519, R1138_U69, U3490);
  nand ginst1439 (R1138_U52, R1138_U136, R1138_U232);
  nand ginst1440 (R1138_U520, R1138_U518, R1138_U519);
  nand ginst1441 (R1138_U521, R1138_U106, R1138_U370);
  nand ginst1442 (R1138_U522, R1138_U346, R1138_U520);
  nand ginst1443 (R1138_U523, R1138_U70, U3060);
  nand ginst1444 (R1138_U524, R1138_U71, U3488);
  nand ginst1445 (R1138_U525, R1138_U523, R1138_U524);
  nand ginst1446 (R1138_U526, R1138_U184, R1138_U371);
  nand ginst1447 (R1138_U527, R1138_U256, R1138_U525);
  nand ginst1448 (R1138_U528, R1138_U66, U3059);
  nand ginst1449 (R1138_U529, R1138_U67, U3486);
  nand ginst1450 (R1138_U53, R1138_U228, R1138_U229);
  nand ginst1451 (R1138_U530, R1138_U37, U3074);
  nand ginst1452 (R1138_U531, R1138_U38, U3464);
  not ginst1453 (R1138_U54, U4030);
  not ginst1454 (R1138_U55, U3050);
  not ginst1455 (R1138_U56, U3054);
  not ginst1456 (R1138_U57, U4031);
  not ginst1457 (R1138_U58, U4033);
  not ginst1458 (R1138_U59, U3062);
  and ginst1459 (R1138_U6, R1138_U209, R1138_U210);
  nand ginst1460 (R1138_U60, U3062, U4033);
  not ginst1461 (R1138_U61, U4035);
  not ginst1462 (R1138_U62, U3058);
  not ginst1463 (R1138_U63, U3496);
  not ginst1464 (R1138_U64, U3071);
  nand ginst1465 (R1138_U65, U3081, U3482);
  not ginst1466 (R1138_U66, U3486);
  not ginst1467 (R1138_U67, U3059);
  not ginst1468 (R1138_U68, U3490);
  not ginst1469 (R1138_U69, U3069);
  and ginst1470 (R1138_U7, R1138_U249, R1138_U250);
  not ginst1471 (R1138_U70, U3488);
  not ginst1472 (R1138_U71, U3060);
  nand ginst1473 (R1138_U72, U3060, U3488);
  not ginst1474 (R1138_U73, U3492);
  not ginst1475 (R1138_U74, U3077);
  not ginst1476 (R1138_U75, U3494);
  not ginst1477 (R1138_U76, U3076);
  nand ginst1478 (R1138_U77, R1138_U267, R1138_U380);
  not ginst1479 (R1138_U78, U3504);
  not ginst1480 (R1138_U79, U3078);
  and ginst1481 (R1138_U8, R1138_U257, R1138_U258);
  nand ginst1482 (R1138_U80, U3078, U3504);
  not ginst1483 (R1138_U81, U4037);
  not ginst1484 (R1138_U82, U3502);
  not ginst1485 (R1138_U83, U3079);
  nand ginst1486 (R1138_U84, U3079, U3502);
  not ginst1487 (R1138_U85, U4036);
  not ginst1488 (R1138_U86, U3072);
  not ginst1489 (R1138_U87, U3498);
  not ginst1490 (R1138_U88, U3070);
  not ginst1491 (R1138_U89, U3066);
  and ginst1492 (R1138_U9, R1138_U273, R1138_U274);
  nand ginst1493 (R1138_U90, U3070, U3498);
  not ginst1494 (R1138_U91, U3500);
  not ginst1495 (R1138_U92, U4034);
  not ginst1496 (R1138_U93, U3063);
  nand ginst1497 (R1138_U94, R1138_U146, R1138_U388);
  not ginst1498 (R1138_U95, U4032);
  not ginst1499 (R1138_U96, U3055);
  nand ginst1500 (R1138_U97, R1138_U306, R1138_U396, R1138_U397);
  not ginst1501 (R1138_U98, U3051);
  not ginst1502 (R1138_U99, U4029);
  and ginst1503 (R1150_U10, R1150_U269, R1150_U270);
  not ginst1504 (R1150_U100, U4029);
  not ginst1505 (R1150_U101, U3051);
  nand ginst1506 (R1150_U102, R1150_U146, R1150_U367);
  nand ginst1507 (R1150_U103, R1150_U295, R1150_U356);
  nand ginst1508 (R1150_U104, R1150_U293, R1150_U354);
  nand ginst1509 (R1150_U105, R1150_U285, R1150_U352);
  nand ginst1510 (R1150_U106, R1150_U311, R1150_U68);
  nand ginst1511 (R1150_U107, R1150_U322, R1150_U94);
  nand ginst1512 (R1150_U108, R1150_U369, R1150_U88);
  not ginst1513 (R1150_U109, U3074);
  and ginst1514 (R1150_U11, R1150_U206, R1150_U286);
  nand ginst1515 (R1150_U110, R1150_U427, R1150_U428);
  nand ginst1516 (R1150_U111, R1150_U441, R1150_U442);
  nand ginst1517 (R1150_U112, R1150_U446, R1150_U447);
  nand ginst1518 (R1150_U113, R1150_U462, R1150_U463);
  nand ginst1519 (R1150_U114, R1150_U467, R1150_U468);
  nand ginst1520 (R1150_U115, R1150_U472, R1150_U473);
  nand ginst1521 (R1150_U116, R1150_U477, R1150_U478);
  nand ginst1522 (R1150_U117, R1150_U482, R1150_U483);
  nand ginst1523 (R1150_U118, R1150_U498, R1150_U499);
  nand ginst1524 (R1150_U119, R1150_U503, R1150_U504);
  and ginst1525 (R1150_U12, R1150_U287, R1150_U288);
  nand ginst1526 (R1150_U120, R1150_U386, R1150_U387);
  nand ginst1527 (R1150_U121, R1150_U395, R1150_U396);
  nand ginst1528 (R1150_U122, R1150_U402, R1150_U403);
  nand ginst1529 (R1150_U123, R1150_U406, R1150_U407);
  nand ginst1530 (R1150_U124, R1150_U415, R1150_U416);
  nand ginst1531 (R1150_U125, R1150_U436, R1150_U437);
  nand ginst1532 (R1150_U126, R1150_U453, R1150_U454);
  nand ginst1533 (R1150_U127, R1150_U457, R1150_U458);
  nand ginst1534 (R1150_U128, R1150_U489, R1150_U490);
  nand ginst1535 (R1150_U129, R1150_U493, R1150_U494);
  and ginst1536 (R1150_U13, R1150_U209, R1150_U222, R1150_U227);
  nand ginst1537 (R1150_U130, R1150_U510, R1150_U511);
  and ginst1538 (R1150_U131, R1150_U208, R1150_U218);
  and ginst1539 (R1150_U132, R1150_U220, R1150_U221);
  and ginst1540 (R1150_U133, R1150_U13, R1150_U14);
  and ginst1541 (R1150_U134, R1150_U234, R1150_U235);
  and ginst1542 (R1150_U135, R1150_U134, R1150_U346);
  and ginst1543 (R1150_U136, R1150_U33, R1150_U388, R1150_U389);
  and ginst1544 (R1150_U137, R1150_U210, R1150_U392);
  and ginst1545 (R1150_U138, R1150_U250, R1150_U6);
  and ginst1546 (R1150_U139, R1150_U209, R1150_U399);
  and ginst1547 (R1150_U14, R1150_U210, R1150_U232);
  and ginst1548 (R1150_U140, R1150_U408, R1150_U409, R1150_U41);
  and ginst1549 (R1150_U141, R1150_U208, R1150_U412);
  and ginst1550 (R1150_U142, R1150_U18, R1150_U266);
  and ginst1551 (R1150_U143, R1150_U16, R1150_U278);
  and ginst1552 (R1150_U144, R1150_U279, R1150_U351);
  and ginst1553 (R1150_U145, R1150_U21, R1150_U296);
  and ginst1554 (R1150_U146, R1150_U297, R1150_U358);
  and ginst1555 (R1150_U147, R1150_U207, R1150_U298);
  and ginst1556 (R1150_U148, R1150_U301, R1150_U302);
  and ginst1557 (R1150_U149, R1150_U304, R1150_U421);
  and ginst1558 (R1150_U15, R1150_U237, R1150_U7);
  and ginst1559 (R1150_U150, R1150_U301, R1150_U302);
  and ginst1560 (R1150_U151, R1150_U22, R1150_U305);
  nand ginst1561 (R1150_U152, R1150_U424, R1150_U425);
  and ginst1562 (R1150_U153, R1150_U429, R1150_U430, R1150_U98);
  and ginst1563 (R1150_U154, R1150_U207, R1150_U433);
  nand ginst1564 (R1150_U155, R1150_U438, R1150_U439);
  nand ginst1565 (R1150_U156, R1150_U443, R1150_U444);
  and ginst1566 (R1150_U157, R1150_U12, R1150_U317);
  and ginst1567 (R1150_U158, R1150_U206, R1150_U450);
  nand ginst1568 (R1150_U159, R1150_U459, R1150_U460);
  and ginst1569 (R1150_U16, R1150_U273, R1150_U9);
  nand ginst1570 (R1150_U160, R1150_U464, R1150_U465);
  nand ginst1571 (R1150_U161, R1150_U469, R1150_U470);
  nand ginst1572 (R1150_U162, R1150_U474, R1150_U475);
  nand ginst1573 (R1150_U163, R1150_U479, R1150_U480);
  and ginst1574 (R1150_U164, R1150_U10, R1150_U328);
  and ginst1575 (R1150_U165, R1150_U205, R1150_U486);
  nand ginst1576 (R1150_U166, R1150_U495, R1150_U496);
  nand ginst1577 (R1150_U167, R1150_U500, R1150_U501);
  and ginst1578 (R1150_U168, R1150_U337, R1150_U8);
  and ginst1579 (R1150_U169, R1150_U204, R1150_U507);
  and ginst1580 (R1150_U17, R1150_U11, R1150_U291);
  and ginst1581 (R1150_U170, R1150_U384, R1150_U385);
  nand ginst1582 (R1150_U171, R1150_U135, R1150_U345);
  and ginst1583 (R1150_U172, R1150_U393, R1150_U394);
  and ginst1584 (R1150_U173, R1150_U400, R1150_U401);
  and ginst1585 (R1150_U174, R1150_U404, R1150_U405);
  nand ginst1586 (R1150_U175, R1150_U132, R1150_U377);
  and ginst1587 (R1150_U176, R1150_U413, R1150_U414);
  not ginst1588 (R1150_U177, U4040);
  not ginst1589 (R1150_U178, U3052);
  and ginst1590 (R1150_U179, R1150_U422, R1150_U423);
  and ginst1591 (R1150_U18, R1150_U15, R1150_U264);
  nand ginst1592 (R1150_U180, R1150_U148, R1150_U299);
  and ginst1593 (R1150_U181, R1150_U434, R1150_U435);
  nand ginst1594 (R1150_U182, R1150_U357, R1150_U365);
  nand ginst1595 (R1150_U183, R1150_U355, R1150_U363);
  and ginst1596 (R1150_U184, R1150_U451, R1150_U452);
  and ginst1597 (R1150_U185, R1150_U455, R1150_U456);
  nand ginst1598 (R1150_U186, R1150_U353, R1150_U361);
  nand ginst1599 (R1150_U187, R1150_U359, R1150_U73);
  not ginst1600 (R1150_U188, U3468);
  nand ginst1601 (R1150_U189, R1150_U109, U3464);
  and ginst1602 (R1150_U19, R1150_U282, R1150_U284);
  nand ginst1603 (R1150_U190, R1150_U343, R1150_U382);
  nand ginst1604 (R1150_U191, R1150_U144, R1150_U350);
  nand ginst1605 (R1150_U192, R1150_U275, R1150_U95);
  and ginst1606 (R1150_U193, R1150_U487, R1150_U488);
  and ginst1607 (R1150_U194, R1150_U491, R1150_U492);
  nand ginst1608 (R1150_U195, R1150_U267, R1150_U349, R1150_U375);
  nand ginst1609 (R1150_U196, R1150_U373, R1150_U90);
  nand ginst1610 (R1150_U197, R1150_U263, R1150_U371);
  and ginst1611 (R1150_U198, R1150_U508, R1150_U509);
  nand ginst1612 (R1150_U199, R1150_U149, R1150_U180);
  and ginst1613 (R1150_U20, R1150_U17, R1150_U19);
  nand ginst1614 (R1150_U200, R1150_U188, R1150_U189);
  not ginst1615 (R1150_U201, R1150_U98);
  not ginst1616 (R1150_U202, R1150_U41);
  not ginst1617 (R1150_U203, R1150_U33);
  nand ginst1618 (R1150_U204, R1150_U85, U3486);
  nand ginst1619 (R1150_U205, R1150_U92, U3496);
  nand ginst1620 (R1150_U206, R1150_U64, U4035);
  nand ginst1621 (R1150_U207, R1150_U97, U4031);
  nand ginst1622 (R1150_U208, R1150_U40, U3470);
  nand ginst1623 (R1150_U209, R1150_U48, U3476);
  and ginst1624 (R1150_U21, R1150_U20, R1150_U294);
  nand ginst1625 (R1150_U210, R1150_U32, U3480);
  not ginst1626 (R1150_U211, R1150_U94);
  not ginst1627 (R1150_U212, R1150_U68);
  not ginst1628 (R1150_U213, R1150_U50);
  not ginst1629 (R1150_U214, R1150_U88);
  not ginst1630 (R1150_U215, R1150_U189);
  nand ginst1631 (R1150_U216, R1150_U189, U3075);
  not ginst1632 (R1150_U217, R1150_U56);
  nand ginst1633 (R1150_U218, R1150_U42, U3472);
  nand ginst1634 (R1150_U219, R1150_U41, R1150_U42);
  and ginst1635 (R1150_U22, R1150_U417, R1150_U418);
  nand ginst1636 (R1150_U220, R1150_U219, R1150_U46);
  nand ginst1637 (R1150_U221, R1150_U202, U3061);
  nand ginst1638 (R1150_U222, R1150_U47, U3478);
  nand ginst1639 (R1150_U223, R1150_U36, U3068);
  nand ginst1640 (R1150_U224, R1150_U35, U3064);
  nand ginst1641 (R1150_U225, R1150_U209, R1150_U213);
  nand ginst1642 (R1150_U226, R1150_U225, R1150_U6);
  nand ginst1643 (R1150_U227, R1150_U49, U3474);
  nand ginst1644 (R1150_U228, R1150_U47, U3478);
  nand ginst1645 (R1150_U229, R1150_U13, R1150_U175);
  nand ginst1646 (R1150_U23, R1150_U335, R1150_U338);
  not ginst1647 (R1150_U230, R1150_U51);
  not ginst1648 (R1150_U231, R1150_U54);
  nand ginst1649 (R1150_U232, R1150_U34, U3482);
  nand ginst1650 (R1150_U233, R1150_U33, R1150_U34);
  nand ginst1651 (R1150_U234, R1150_U233, R1150_U39);
  nand ginst1652 (R1150_U235, R1150_U203, U3081);
  not ginst1653 (R1150_U236, R1150_U171);
  nand ginst1654 (R1150_U237, R1150_U53, U3484);
  nand ginst1655 (R1150_U238, R1150_U237, R1150_U88);
  nand ginst1656 (R1150_U239, R1150_U231, R1150_U33);
  nand ginst1657 (R1150_U24, R1150_U326, R1150_U329);
  nand ginst1658 (R1150_U240, R1150_U137, R1150_U239);
  nand ginst1659 (R1150_U241, R1150_U210, R1150_U54);
  nand ginst1660 (R1150_U242, R1150_U136, R1150_U241);
  nand ginst1661 (R1150_U243, R1150_U210, R1150_U33);
  nand ginst1662 (R1150_U244, R1150_U175, R1150_U227);
  not ginst1663 (R1150_U245, R1150_U55);
  nand ginst1664 (R1150_U246, R1150_U35, U3064);
  nand ginst1665 (R1150_U247, R1150_U245, R1150_U246);
  nand ginst1666 (R1150_U248, R1150_U139, R1150_U247);
  nand ginst1667 (R1150_U249, R1150_U209, R1150_U55);
  nand ginst1668 (R1150_U25, R1150_U315, R1150_U318);
  nand ginst1669 (R1150_U250, R1150_U47, U3478);
  nand ginst1670 (R1150_U251, R1150_U138, R1150_U249);
  nand ginst1671 (R1150_U252, R1150_U35, U3064);
  nand ginst1672 (R1150_U253, R1150_U209, R1150_U252);
  nand ginst1673 (R1150_U254, R1150_U227, R1150_U50);
  nand ginst1674 (R1150_U255, R1150_U141, R1150_U381);
  nand ginst1675 (R1150_U256, R1150_U208, R1150_U41);
  nand ginst1676 (R1150_U257, R1150_U84, U3488);
  nand ginst1677 (R1150_U258, R1150_U86, U3060);
  nand ginst1678 (R1150_U259, R1150_U87, U3059);
  nand ginst1679 (R1150_U26, R1150_U307, R1150_U309);
  nand ginst1680 (R1150_U260, R1150_U214, R1150_U7);
  nand ginst1681 (R1150_U261, R1150_U260, R1150_U8);
  nand ginst1682 (R1150_U262, R1150_U84, U3488);
  nand ginst1683 (R1150_U263, R1150_U261, R1150_U262);
  nand ginst1684 (R1150_U264, R1150_U89, U3490);
  nand ginst1685 (R1150_U265, R1150_U83, U3069);
  nand ginst1686 (R1150_U266, R1150_U81, U3492);
  nand ginst1687 (R1150_U267, R1150_U82, U3077);
  nand ginst1688 (R1150_U268, R1150_U91, U3498);
  nand ginst1689 (R1150_U269, R1150_U78, U3070);
  nand ginst1690 (R1150_U27, R1150_U179, R1150_U199, R1150_U344);
  nand ginst1691 (R1150_U270, R1150_U79, U3071);
  nand ginst1692 (R1150_U271, R1150_U211, R1150_U9);
  nand ginst1693 (R1150_U272, R1150_U10, R1150_U271);
  nand ginst1694 (R1150_U273, R1150_U93, U3494);
  nand ginst1695 (R1150_U274, R1150_U91, U3498);
  nand ginst1696 (R1150_U275, R1150_U16, R1150_U195);
  not ginst1697 (R1150_U276, R1150_U95);
  not ginst1698 (R1150_U277, R1150_U192);
  nand ginst1699 (R1150_U278, R1150_U76, U3500);
  nand ginst1700 (R1150_U279, R1150_U77, U3066);
  nand ginst1701 (R1150_U28, R1150_U255, R1150_U380);
  not ginst1702 (R1150_U280, R1150_U191);
  nand ginst1703 (R1150_U281, R1150_U75, U3502);
  nand ginst1704 (R1150_U282, R1150_U71, U3504);
  not ginst1705 (R1150_U283, R1150_U73);
  nand ginst1706 (R1150_U284, R1150_U70, U4037);
  nand ginst1707 (R1150_U285, R1150_U72, U3073);
  nand ginst1708 (R1150_U286, R1150_U63, U4034);
  nand ginst1709 (R1150_U287, R1150_U66, U3063);
  nand ginst1710 (R1150_U288, R1150_U67, U3058);
  nand ginst1711 (R1150_U289, R1150_U11, R1150_U212);
  nand ginst1712 (R1150_U29, R1150_U248, R1150_U251);
  nand ginst1713 (R1150_U290, R1150_U12, R1150_U289);
  nand ginst1714 (R1150_U291, R1150_U65, U4036);
  nand ginst1715 (R1150_U292, R1150_U63, U4034);
  nand ginst1716 (R1150_U293, R1150_U290, R1150_U292);
  nand ginst1717 (R1150_U294, R1150_U61, U4033);
  nand ginst1718 (R1150_U295, R1150_U62, U3062);
  nand ginst1719 (R1150_U296, R1150_U59, U4032);
  nand ginst1720 (R1150_U297, R1150_U60, U3055);
  nand ginst1721 (R1150_U298, R1150_U99, U4030);
  nand ginst1722 (R1150_U299, R1150_U102, R1150_U147);
  nand ginst1723 (R1150_U30, R1150_U240, R1150_U242);
  nand ginst1724 (R1150_U300, R1150_U98, R1150_U99);
  nand ginst1725 (R1150_U301, R1150_U300, R1150_U58);
  nand ginst1726 (R1150_U302, R1150_U201, U3050);
  not ginst1727 (R1150_U303, R1150_U180);
  nand ginst1728 (R1150_U304, R1150_U101, U4029);
  nand ginst1729 (R1150_U305, R1150_U100, U3051);
  nand ginst1730 (R1150_U306, R1150_U368, R1150_U98);
  nand ginst1731 (R1150_U307, R1150_U154, R1150_U306);
  nand ginst1732 (R1150_U308, R1150_U102, R1150_U207);
  nand ginst1733 (R1150_U309, R1150_U153, R1150_U308);
  nand ginst1734 (R1150_U31, R1150_U189, R1150_U341);
  nand ginst1735 (R1150_U310, R1150_U207, R1150_U98);
  nand ginst1736 (R1150_U311, R1150_U186, R1150_U291);
  not ginst1737 (R1150_U312, R1150_U106);
  nand ginst1738 (R1150_U313, R1150_U67, U3058);
  nand ginst1739 (R1150_U314, R1150_U312, R1150_U313);
  nand ginst1740 (R1150_U315, R1150_U158, R1150_U314);
  nand ginst1741 (R1150_U316, R1150_U106, R1150_U206);
  nand ginst1742 (R1150_U317, R1150_U63, U4034);
  nand ginst1743 (R1150_U318, R1150_U157, R1150_U316);
  nand ginst1744 (R1150_U319, R1150_U67, U3058);
  not ginst1745 (R1150_U32, U3067);
  nand ginst1746 (R1150_U320, R1150_U206, R1150_U319);
  nand ginst1747 (R1150_U321, R1150_U291, R1150_U68);
  nand ginst1748 (R1150_U322, R1150_U195, R1150_U273);
  not ginst1749 (R1150_U323, R1150_U107);
  nand ginst1750 (R1150_U324, R1150_U79, U3071);
  nand ginst1751 (R1150_U325, R1150_U323, R1150_U324);
  nand ginst1752 (R1150_U326, R1150_U165, R1150_U325);
  nand ginst1753 (R1150_U327, R1150_U107, R1150_U205);
  nand ginst1754 (R1150_U328, R1150_U91, U3498);
  nand ginst1755 (R1150_U329, R1150_U164, R1150_U327);
  nand ginst1756 (R1150_U33, R1150_U38, U3067);
  nand ginst1757 (R1150_U330, R1150_U79, U3071);
  nand ginst1758 (R1150_U331, R1150_U205, R1150_U330);
  nand ginst1759 (R1150_U332, R1150_U273, R1150_U94);
  nand ginst1760 (R1150_U333, R1150_U87, U3059);
  nand ginst1761 (R1150_U334, R1150_U333, R1150_U370);
  nand ginst1762 (R1150_U335, R1150_U169, R1150_U334);
  nand ginst1763 (R1150_U336, R1150_U108, R1150_U204);
  nand ginst1764 (R1150_U337, R1150_U84, U3488);
  nand ginst1765 (R1150_U338, R1150_U168, R1150_U336);
  nand ginst1766 (R1150_U339, R1150_U87, U3059);
  not ginst1767 (R1150_U34, U3081);
  nand ginst1768 (R1150_U340, R1150_U204, R1150_U339);
  nand ginst1769 (R1150_U341, R1150_U44, U3074);
  nand ginst1770 (R1150_U342, R1150_U188, U3075);
  nand ginst1771 (R1150_U343, R1150_U96, U3079);
  nand ginst1772 (R1150_U344, R1150_U150, R1150_U151, R1150_U299);
  nand ginst1773 (R1150_U345, R1150_U133, R1150_U175);
  nand ginst1774 (R1150_U346, R1150_U14, R1150_U230);
  nand ginst1775 (R1150_U347, R1150_U263, R1150_U265);
  not ginst1776 (R1150_U348, R1150_U90);
  nand ginst1777 (R1150_U349, R1150_U266, R1150_U348);
  not ginst1778 (R1150_U35, U3476);
  nand ginst1779 (R1150_U350, R1150_U143, R1150_U195);
  nand ginst1780 (R1150_U351, R1150_U276, R1150_U278);
  nand ginst1781 (R1150_U352, R1150_U283, R1150_U284);
  not ginst1782 (R1150_U353, R1150_U105);
  nand ginst1783 (R1150_U354, R1150_U105, R1150_U17);
  not ginst1784 (R1150_U355, R1150_U104);
  nand ginst1785 (R1150_U356, R1150_U104, R1150_U294);
  not ginst1786 (R1150_U357, R1150_U103);
  nand ginst1787 (R1150_U358, R1150_U103, R1150_U296);
  nand ginst1788 (R1150_U359, R1150_U190, R1150_U282);
  not ginst1789 (R1150_U36, U3478);
  not ginst1790 (R1150_U360, R1150_U187);
  nand ginst1791 (R1150_U361, R1150_U19, R1150_U190);
  not ginst1792 (R1150_U362, R1150_U186);
  nand ginst1793 (R1150_U363, R1150_U190, R1150_U20);
  not ginst1794 (R1150_U364, R1150_U183);
  nand ginst1795 (R1150_U365, R1150_U190, R1150_U21);
  not ginst1796 (R1150_U366, R1150_U182);
  nand ginst1797 (R1150_U367, R1150_U145, R1150_U190);
  not ginst1798 (R1150_U368, R1150_U102);
  nand ginst1799 (R1150_U369, R1150_U171, R1150_U237);
  not ginst1800 (R1150_U37, U3474);
  not ginst1801 (R1150_U370, R1150_U108);
  nand ginst1802 (R1150_U371, R1150_U15, R1150_U171);
  not ginst1803 (R1150_U372, R1150_U197);
  nand ginst1804 (R1150_U373, R1150_U171, R1150_U18);
  not ginst1805 (R1150_U374, R1150_U196);
  nand ginst1806 (R1150_U375, R1150_U142, R1150_U171);
  not ginst1807 (R1150_U376, R1150_U195);
  nand ginst1808 (R1150_U377, R1150_U131, R1150_U56);
  not ginst1809 (R1150_U378, R1150_U175);
  nand ginst1810 (R1150_U379, R1150_U208, R1150_U56);
  not ginst1811 (R1150_U38, U3480);
  nand ginst1812 (R1150_U380, R1150_U140, R1150_U379);
  nand ginst1813 (R1150_U381, R1150_U217, R1150_U41);
  nand ginst1814 (R1150_U382, R1150_U191, R1150_U281);
  not ginst1815 (R1150_U383, R1150_U190);
  nand ginst1816 (R1150_U384, R1150_U53, U3484);
  nand ginst1817 (R1150_U385, R1150_U52, U3080);
  nand ginst1818 (R1150_U386, R1150_U171, R1150_U238);
  nand ginst1819 (R1150_U387, R1150_U170, R1150_U236);
  nand ginst1820 (R1150_U388, R1150_U34, U3482);
  nand ginst1821 (R1150_U389, R1150_U39, U3081);
  not ginst1822 (R1150_U39, U3482);
  nand ginst1823 (R1150_U390, R1150_U34, U3482);
  nand ginst1824 (R1150_U391, R1150_U39, U3081);
  nand ginst1825 (R1150_U392, R1150_U390, R1150_U391);
  nand ginst1826 (R1150_U393, R1150_U32, U3480);
  nand ginst1827 (R1150_U394, R1150_U38, U3067);
  nand ginst1828 (R1150_U395, R1150_U243, R1150_U54);
  nand ginst1829 (R1150_U396, R1150_U172, R1150_U231);
  nand ginst1830 (R1150_U397, R1150_U47, U3478);
  nand ginst1831 (R1150_U398, R1150_U36, U3068);
  nand ginst1832 (R1150_U399, R1150_U397, R1150_U398);
  not ginst1833 (R1150_U40, U3065);
  nand ginst1834 (R1150_U400, R1150_U48, U3476);
  nand ginst1835 (R1150_U401, R1150_U35, U3064);
  nand ginst1836 (R1150_U402, R1150_U253, R1150_U55);
  nand ginst1837 (R1150_U403, R1150_U173, R1150_U245);
  nand ginst1838 (R1150_U404, R1150_U49, U3474);
  nand ginst1839 (R1150_U405, R1150_U37, U3057);
  nand ginst1840 (R1150_U406, R1150_U175, R1150_U254);
  nand ginst1841 (R1150_U407, R1150_U174, R1150_U378);
  nand ginst1842 (R1150_U408, R1150_U42, U3472);
  nand ginst1843 (R1150_U409, R1150_U46, U3061);
  nand ginst1844 (R1150_U41, R1150_U43, U3065);
  nand ginst1845 (R1150_U410, R1150_U42, U3472);
  nand ginst1846 (R1150_U411, R1150_U46, U3061);
  nand ginst1847 (R1150_U412, R1150_U410, R1150_U411);
  nand ginst1848 (R1150_U413, R1150_U40, U3470);
  nand ginst1849 (R1150_U414, R1150_U43, U3065);
  nand ginst1850 (R1150_U415, R1150_U256, R1150_U56);
  nand ginst1851 (R1150_U416, R1150_U176, R1150_U217);
  nand ginst1852 (R1150_U417, R1150_U178, U4040);
  nand ginst1853 (R1150_U418, R1150_U177, U3052);
  nand ginst1854 (R1150_U419, R1150_U178, U4040);
  not ginst1855 (R1150_U42, U3061);
  nand ginst1856 (R1150_U420, R1150_U177, U3052);
  nand ginst1857 (R1150_U421, R1150_U419, R1150_U420);
  nand ginst1858 (R1150_U422, R1150_U100, R1150_U421, U3051);
  nand ginst1859 (R1150_U423, R1150_U101, R1150_U22, U4029);
  nand ginst1860 (R1150_U424, R1150_U101, U4029);
  nand ginst1861 (R1150_U425, R1150_U100, U3051);
  not ginst1862 (R1150_U426, R1150_U152);
  nand ginst1863 (R1150_U427, R1150_U303, R1150_U426);
  nand ginst1864 (R1150_U428, R1150_U152, R1150_U180);
  nand ginst1865 (R1150_U429, R1150_U99, U4030);
  not ginst1866 (R1150_U43, U3470);
  nand ginst1867 (R1150_U430, R1150_U58, U3050);
  nand ginst1868 (R1150_U431, R1150_U99, U4030);
  nand ginst1869 (R1150_U432, R1150_U58, U3050);
  nand ginst1870 (R1150_U433, R1150_U431, R1150_U432);
  nand ginst1871 (R1150_U434, R1150_U97, U4031);
  nand ginst1872 (R1150_U435, R1150_U57, U3054);
  nand ginst1873 (R1150_U436, R1150_U102, R1150_U310);
  nand ginst1874 (R1150_U437, R1150_U181, R1150_U368);
  nand ginst1875 (R1150_U438, R1150_U59, U4032);
  nand ginst1876 (R1150_U439, R1150_U60, U3055);
  not ginst1877 (R1150_U44, U3464);
  not ginst1878 (R1150_U440, R1150_U155);
  nand ginst1879 (R1150_U441, R1150_U366, R1150_U440);
  nand ginst1880 (R1150_U442, R1150_U155, R1150_U182);
  nand ginst1881 (R1150_U443, R1150_U61, U4033);
  nand ginst1882 (R1150_U444, R1150_U62, U3062);
  not ginst1883 (R1150_U445, R1150_U156);
  nand ginst1884 (R1150_U446, R1150_U364, R1150_U445);
  nand ginst1885 (R1150_U447, R1150_U156, R1150_U183);
  nand ginst1886 (R1150_U448, R1150_U63, U4034);
  nand ginst1887 (R1150_U449, R1150_U66, U3063);
  not ginst1888 (R1150_U45, U3075);
  nand ginst1889 (R1150_U450, R1150_U448, R1150_U449);
  nand ginst1890 (R1150_U451, R1150_U64, U4035);
  nand ginst1891 (R1150_U452, R1150_U67, U3058);
  nand ginst1892 (R1150_U453, R1150_U106, R1150_U320);
  nand ginst1893 (R1150_U454, R1150_U184, R1150_U312);
  nand ginst1894 (R1150_U455, R1150_U65, U4036);
  nand ginst1895 (R1150_U456, R1150_U69, U3072);
  nand ginst1896 (R1150_U457, R1150_U186, R1150_U321);
  nand ginst1897 (R1150_U458, R1150_U185, R1150_U362);
  nand ginst1898 (R1150_U459, R1150_U70, U4037);
  not ginst1899 (R1150_U46, U3472);
  nand ginst1900 (R1150_U460, R1150_U72, U3073);
  not ginst1901 (R1150_U461, R1150_U159);
  nand ginst1902 (R1150_U462, R1150_U360, R1150_U461);
  nand ginst1903 (R1150_U463, R1150_U159, R1150_U187);
  nand ginst1904 (R1150_U464, R1150_U45, U3468);
  nand ginst1905 (R1150_U465, R1150_U188, U3075);
  not ginst1906 (R1150_U466, R1150_U160);
  nand ginst1907 (R1150_U467, R1150_U215, R1150_U466);
  nand ginst1908 (R1150_U468, R1150_U160, R1150_U189);
  nand ginst1909 (R1150_U469, R1150_U71, U3504);
  not ginst1910 (R1150_U47, U3068);
  nand ginst1911 (R1150_U470, R1150_U74, U3078);
  not ginst1912 (R1150_U471, R1150_U161);
  nand ginst1913 (R1150_U472, R1150_U383, R1150_U471);
  nand ginst1914 (R1150_U473, R1150_U161, R1150_U190);
  nand ginst1915 (R1150_U474, R1150_U75, U3502);
  nand ginst1916 (R1150_U475, R1150_U96, U3079);
  not ginst1917 (R1150_U476, R1150_U162);
  nand ginst1918 (R1150_U477, R1150_U280, R1150_U476);
  nand ginst1919 (R1150_U478, R1150_U162, R1150_U191);
  nand ginst1920 (R1150_U479, R1150_U76, U3500);
  not ginst1921 (R1150_U48, U3064);
  nand ginst1922 (R1150_U480, R1150_U77, U3066);
  not ginst1923 (R1150_U481, R1150_U163);
  nand ginst1924 (R1150_U482, R1150_U277, R1150_U481);
  nand ginst1925 (R1150_U483, R1150_U163, R1150_U192);
  nand ginst1926 (R1150_U484, R1150_U91, U3498);
  nand ginst1927 (R1150_U485, R1150_U78, U3070);
  nand ginst1928 (R1150_U486, R1150_U484, R1150_U485);
  nand ginst1929 (R1150_U487, R1150_U92, U3496);
  nand ginst1930 (R1150_U488, R1150_U79, U3071);
  nand ginst1931 (R1150_U489, R1150_U107, R1150_U331);
  not ginst1932 (R1150_U49, U3057);
  nand ginst1933 (R1150_U490, R1150_U193, R1150_U323);
  nand ginst1934 (R1150_U491, R1150_U93, U3494);
  nand ginst1935 (R1150_U492, R1150_U80, U3076);
  nand ginst1936 (R1150_U493, R1150_U195, R1150_U332);
  nand ginst1937 (R1150_U494, R1150_U194, R1150_U376);
  nand ginst1938 (R1150_U495, R1150_U81, U3492);
  nand ginst1939 (R1150_U496, R1150_U82, U3077);
  not ginst1940 (R1150_U497, R1150_U166);
  nand ginst1941 (R1150_U498, R1150_U374, R1150_U497);
  nand ginst1942 (R1150_U499, R1150_U166, R1150_U196);
  nand ginst1943 (R1150_U50, R1150_U37, U3057);
  nand ginst1944 (R1150_U500, R1150_U89, U3490);
  nand ginst1945 (R1150_U501, R1150_U83, U3069);
  not ginst1946 (R1150_U502, R1150_U167);
  nand ginst1947 (R1150_U503, R1150_U372, R1150_U502);
  nand ginst1948 (R1150_U504, R1150_U167, R1150_U197);
  nand ginst1949 (R1150_U505, R1150_U84, U3488);
  nand ginst1950 (R1150_U506, R1150_U86, U3060);
  nand ginst1951 (R1150_U507, R1150_U505, R1150_U506);
  nand ginst1952 (R1150_U508, R1150_U85, U3486);
  nand ginst1953 (R1150_U509, R1150_U87, U3059);
  nand ginst1954 (R1150_U51, R1150_U226, R1150_U228);
  nand ginst1955 (R1150_U510, R1150_U108, R1150_U340);
  nand ginst1956 (R1150_U511, R1150_U198, R1150_U370);
  not ginst1957 (R1150_U52, U3484);
  not ginst1958 (R1150_U53, U3080);
  nand ginst1959 (R1150_U54, R1150_U229, R1150_U51);
  nand ginst1960 (R1150_U55, R1150_U244, R1150_U50);
  nand ginst1961 (R1150_U56, R1150_U200, R1150_U216, R1150_U342);
  not ginst1962 (R1150_U57, U4031);
  not ginst1963 (R1150_U58, U4030);
  not ginst1964 (R1150_U59, U3055);
  and ginst1965 (R1150_U6, R1150_U223, R1150_U224);
  not ginst1966 (R1150_U60, U4032);
  not ginst1967 (R1150_U61, U3062);
  not ginst1968 (R1150_U62, U4033);
  not ginst1969 (R1150_U63, U3063);
  not ginst1970 (R1150_U64, U3058);
  not ginst1971 (R1150_U65, U3072);
  not ginst1972 (R1150_U66, U4034);
  not ginst1973 (R1150_U67, U4035);
  nand ginst1974 (R1150_U68, R1150_U69, U3072);
  not ginst1975 (R1150_U69, U4036);
  and ginst1976 (R1150_U7, R1150_U204, R1150_U257);
  not ginst1977 (R1150_U70, U3073);
  not ginst1978 (R1150_U71, U3078);
  not ginst1979 (R1150_U72, U4037);
  nand ginst1980 (R1150_U73, R1150_U74, U3078);
  not ginst1981 (R1150_U74, U3504);
  not ginst1982 (R1150_U75, U3079);
  not ginst1983 (R1150_U76, U3066);
  not ginst1984 (R1150_U77, U3500);
  not ginst1985 (R1150_U78, U3498);
  not ginst1986 (R1150_U79, U3496);
  and ginst1987 (R1150_U8, R1150_U258, R1150_U259);
  not ginst1988 (R1150_U80, U3494);
  not ginst1989 (R1150_U81, U3077);
  not ginst1990 (R1150_U82, U3492);
  not ginst1991 (R1150_U83, U3490);
  not ginst1992 (R1150_U84, U3060);
  not ginst1993 (R1150_U85, U3059);
  not ginst1994 (R1150_U86, U3488);
  not ginst1995 (R1150_U87, U3486);
  nand ginst1996 (R1150_U88, R1150_U52, U3080);
  not ginst1997 (R1150_U89, U3069);
  and ginst1998 (R1150_U9, R1150_U205, R1150_U268);
  nand ginst1999 (R1150_U90, R1150_U264, R1150_U347);
  not ginst2000 (R1150_U91, U3070);
  not ginst2001 (R1150_U92, U3071);
  not ginst2002 (R1150_U93, U3076);
  nand ginst2003 (R1150_U94, R1150_U80, U3076);
  nand ginst2004 (R1150_U95, R1150_U272, R1150_U274);
  not ginst2005 (R1150_U96, U3502);
  not ginst2006 (R1150_U97, U3054);
  nand ginst2007 (R1150_U98, R1150_U57, U3054);
  not ginst2008 (R1150_U99, U3050);
  not ginst2009 (R1162_U10, REG1_REG_1__SCAN_IN);
  not ginst2010 (R1162_U100, R1162_U82);
  or ginst2011 (R1162_U101, REG1_REG_2__SCAN_IN, U3442);
  nand ginst2012 (R1162_U102, R1162_U101, R1162_U82);
  nand ginst2013 (R1162_U103, REG1_REG_2__SCAN_IN, U3442);
  not ginst2014 (R1162_U104, R1162_U13);
  nand ginst2015 (R1162_U105, R1162_U208, U3441);
  nand ginst2016 (R1162_U106, REG1_REG_3__SCAN_IN, R1162_U13);
  not ginst2017 (R1162_U107, R1162_U80);
  or ginst2018 (R1162_U108, REG1_REG_4__SCAN_IN, U3440);
  nand ginst2019 (R1162_U109, R1162_U108, R1162_U80);
  not ginst2020 (R1162_U11, REG1_REG_2__SCAN_IN);
  nand ginst2021 (R1162_U110, REG1_REG_4__SCAN_IN, U3440);
  not ginst2022 (R1162_U111, R1162_U18);
  nand ginst2023 (R1162_U112, R1162_U195, U3439);
  nand ginst2024 (R1162_U113, REG1_REG_5__SCAN_IN, R1162_U18);
  not ginst2025 (R1162_U114, R1162_U78);
  or ginst2026 (R1162_U115, REG1_REG_6__SCAN_IN, U3438);
  nand ginst2027 (R1162_U116, R1162_U115, R1162_U78);
  nand ginst2028 (R1162_U117, REG1_REG_6__SCAN_IN, U3438);
  not ginst2029 (R1162_U118, R1162_U76);
  or ginst2030 (R1162_U119, REG1_REG_7__SCAN_IN, U3437);
  not ginst2031 (R1162_U12, U3442);
  nand ginst2032 (R1162_U120, R1162_U119, R1162_U76);
  nand ginst2033 (R1162_U121, REG1_REG_7__SCAN_IN, U3437);
  not ginst2034 (R1162_U122, R1162_U25);
  nand ginst2035 (R1162_U123, R1162_U175, U3436);
  nand ginst2036 (R1162_U124, REG1_REG_8__SCAN_IN, R1162_U25);
  not ginst2037 (R1162_U125, R1162_U74);
  or ginst2038 (R1162_U126, REG1_REG_9__SCAN_IN, U3435);
  nand ginst2039 (R1162_U127, R1162_U126, R1162_U74);
  nand ginst2040 (R1162_U128, REG1_REG_9__SCAN_IN, U3435);
  not ginst2041 (R1162_U129, R1162_U30);
  nand ginst2042 (R1162_U13, R1162_U102, R1162_U103);
  nand ginst2043 (R1162_U130, R1162_U284, U3452);
  nand ginst2044 (R1162_U131, REG1_REG_10__SCAN_IN, R1162_U30);
  not ginst2045 (R1162_U132, R1162_U95);
  or ginst2046 (R1162_U133, REG1_REG_11__SCAN_IN, U3451);
  nand ginst2047 (R1162_U134, R1162_U133, R1162_U95);
  nand ginst2048 (R1162_U135, REG1_REG_11__SCAN_IN, U3451);
  not ginst2049 (R1162_U136, R1162_U93);
  or ginst2050 (R1162_U137, REG1_REG_12__SCAN_IN, U3450);
  nand ginst2051 (R1162_U138, R1162_U137, R1162_U93);
  nand ginst2052 (R1162_U139, REG1_REG_12__SCAN_IN, U3450);
  not ginst2053 (R1162_U14, U3441);
  not ginst2054 (R1162_U140, R1162_U37);
  nand ginst2055 (R1162_U141, R1162_U264, U3449);
  nand ginst2056 (R1162_U142, REG1_REG_13__SCAN_IN, R1162_U37);
  not ginst2057 (R1162_U143, R1162_U40);
  nand ginst2058 (R1162_U144, R1162_U258, U3448);
  nand ginst2059 (R1162_U145, REG1_REG_14__SCAN_IN, R1162_U40);
  not ginst2060 (R1162_U146, R1162_U43);
  nand ginst2061 (R1162_U147, R1162_U252, U3447);
  nand ginst2062 (R1162_U148, REG1_REG_15__SCAN_IN, R1162_U43);
  not ginst2063 (R1162_U149, R1162_U91);
  not ginst2064 (R1162_U15, REG1_REG_3__SCAN_IN);
  or ginst2065 (R1162_U150, REG1_REG_16__SCAN_IN, U3446);
  nand ginst2066 (R1162_U151, R1162_U150, R1162_U91);
  nand ginst2067 (R1162_U152, REG1_REG_16__SCAN_IN, U3446);
  not ginst2068 (R1162_U153, R1162_U89);
  or ginst2069 (R1162_U154, REG1_REG_17__SCAN_IN, U3445);
  nand ginst2070 (R1162_U155, R1162_U154, R1162_U89);
  nand ginst2071 (R1162_U156, REG1_REG_17__SCAN_IN, U3445);
  not ginst2072 (R1162_U157, R1162_U52);
  or ginst2073 (R1162_U158, REG1_REG_18__SCAN_IN, U3444);
  nand ginst2074 (R1162_U159, R1162_U158, R1162_U52);
  not ginst2075 (R1162_U16, REG1_REG_4__SCAN_IN);
  nand ginst2076 (R1162_U160, REG1_REG_18__SCAN_IN, U3444);
  nand ginst2077 (R1162_U161, R1162_U159, R1162_U71);
  nand ginst2078 (R1162_U162, REG1_REG_18__SCAN_IN, U3444);
  nand ginst2079 (R1162_U163, R1162_U157, R1162_U162);
  or ginst2080 (R1162_U164, REG1_REG_18__SCAN_IN, U3444);
  nand ginst2081 (R1162_U165, R1162_U163, R1162_U72);
  nand ginst2082 (R1162_U166, R1162_U10, R1162_U222);
  nand ginst2083 (R1162_U167, R1162_U29, U3435);
  nand ginst2084 (R1162_U168, REG1_REG_9__SCAN_IN, R1162_U28);
  nand ginst2085 (R1162_U169, R1162_U29, U3435);
  not ginst2086 (R1162_U17, U3440);
  nand ginst2087 (R1162_U170, REG1_REG_9__SCAN_IN, R1162_U28);
  nand ginst2088 (R1162_U171, R1162_U169, R1162_U170);
  nand ginst2089 (R1162_U172, R1162_U73, R1162_U74);
  nand ginst2090 (R1162_U173, R1162_U125, R1162_U171);
  nand ginst2091 (R1162_U174, REG1_REG_8__SCAN_IN, R1162_U25);
  nand ginst2092 (R1162_U175, R1162_U122, R1162_U27);
  nand ginst2093 (R1162_U176, REG1_REG_8__SCAN_IN, R1162_U25);
  nand ginst2094 (R1162_U177, R1162_U175, R1162_U176);
  nand ginst2095 (R1162_U178, R1162_U174, R1162_U175, R1162_U26);
  nand ginst2096 (R1162_U179, R1162_U177, U3436);
  nand ginst2097 (R1162_U18, R1162_U109, R1162_U110);
  nand ginst2098 (R1162_U180, R1162_U23, U3437);
  nand ginst2099 (R1162_U181, REG1_REG_7__SCAN_IN, R1162_U24);
  nand ginst2100 (R1162_U182, R1162_U23, U3437);
  nand ginst2101 (R1162_U183, REG1_REG_7__SCAN_IN, R1162_U24);
  nand ginst2102 (R1162_U184, R1162_U182, R1162_U183);
  nand ginst2103 (R1162_U185, R1162_U75, R1162_U76);
  nand ginst2104 (R1162_U186, R1162_U118, R1162_U184);
  nand ginst2105 (R1162_U187, R1162_U21, U3438);
  nand ginst2106 (R1162_U188, REG1_REG_6__SCAN_IN, R1162_U22);
  nand ginst2107 (R1162_U189, R1162_U21, U3438);
  not ginst2108 (R1162_U19, U3439);
  nand ginst2109 (R1162_U190, REG1_REG_6__SCAN_IN, R1162_U22);
  nand ginst2110 (R1162_U191, R1162_U189, R1162_U190);
  nand ginst2111 (R1162_U192, R1162_U77, R1162_U78);
  nand ginst2112 (R1162_U193, R1162_U114, R1162_U191);
  nand ginst2113 (R1162_U194, REG1_REG_5__SCAN_IN, R1162_U18);
  nand ginst2114 (R1162_U195, R1162_U111, R1162_U20);
  nand ginst2115 (R1162_U196, REG1_REG_5__SCAN_IN, R1162_U18);
  nand ginst2116 (R1162_U197, R1162_U195, R1162_U196);
  nand ginst2117 (R1162_U198, R1162_U19, R1162_U194, R1162_U195);
  nand ginst2118 (R1162_U199, R1162_U197, U3439);
  not ginst2119 (R1162_U20, REG1_REG_5__SCAN_IN);
  nand ginst2120 (R1162_U200, R1162_U16, U3440);
  nand ginst2121 (R1162_U201, REG1_REG_4__SCAN_IN, R1162_U17);
  nand ginst2122 (R1162_U202, R1162_U16, U3440);
  nand ginst2123 (R1162_U203, REG1_REG_4__SCAN_IN, R1162_U17);
  nand ginst2124 (R1162_U204, R1162_U202, R1162_U203);
  nand ginst2125 (R1162_U205, R1162_U79, R1162_U80);
  nand ginst2126 (R1162_U206, R1162_U107, R1162_U204);
  nand ginst2127 (R1162_U207, REG1_REG_3__SCAN_IN, R1162_U13);
  nand ginst2128 (R1162_U208, R1162_U104, R1162_U15);
  nand ginst2129 (R1162_U209, REG1_REG_3__SCAN_IN, R1162_U13);
  not ginst2130 (R1162_U21, REG1_REG_6__SCAN_IN);
  nand ginst2131 (R1162_U210, R1162_U208, R1162_U209);
  nand ginst2132 (R1162_U211, R1162_U14, R1162_U207, R1162_U208);
  nand ginst2133 (R1162_U212, R1162_U210, U3441);
  nand ginst2134 (R1162_U213, R1162_U11, U3442);
  nand ginst2135 (R1162_U214, REG1_REG_2__SCAN_IN, R1162_U12);
  nand ginst2136 (R1162_U215, R1162_U11, U3442);
  nand ginst2137 (R1162_U216, REG1_REG_2__SCAN_IN, R1162_U12);
  nand ginst2138 (R1162_U217, R1162_U215, R1162_U216);
  nand ginst2139 (R1162_U218, R1162_U81, R1162_U82);
  nand ginst2140 (R1162_U219, R1162_U100, R1162_U217);
  not ginst2141 (R1162_U22, U3438);
  nand ginst2142 (R1162_U220, R1162_U9, U3443);
  nand ginst2143 (R1162_U221, R1162_U8, R1162_U97);
  nand ginst2144 (R1162_U222, R1162_U220, R1162_U221);
  nand ginst2145 (R1162_U223, REG1_REG_1__SCAN_IN, R1162_U8, R1162_U9);
  nand ginst2146 (R1162_U224, R1162_U96, U3443);
  nand ginst2147 (R1162_U225, R1162_U86, U3461);
  nand ginst2148 (R1162_U226, REG1_REG_19__SCAN_IN, R1162_U85);
  nand ginst2149 (R1162_U227, R1162_U86, U3461);
  nand ginst2150 (R1162_U228, REG1_REG_19__SCAN_IN, R1162_U85);
  nand ginst2151 (R1162_U229, R1162_U227, R1162_U228);
  not ginst2152 (R1162_U23, REG1_REG_7__SCAN_IN);
  nand ginst2153 (R1162_U230, R1162_U50, U3444);
  nand ginst2154 (R1162_U231, REG1_REG_18__SCAN_IN, R1162_U51);
  nand ginst2155 (R1162_U232, R1162_U50, U3444);
  nand ginst2156 (R1162_U233, REG1_REG_18__SCAN_IN, R1162_U51);
  nand ginst2157 (R1162_U234, R1162_U232, R1162_U233);
  nand ginst2158 (R1162_U235, R1162_U52, R1162_U87);
  nand ginst2159 (R1162_U236, R1162_U157, R1162_U234);
  nand ginst2160 (R1162_U237, R1162_U48, U3445);
  nand ginst2161 (R1162_U238, REG1_REG_17__SCAN_IN, R1162_U49);
  nand ginst2162 (R1162_U239, R1162_U48, U3445);
  not ginst2163 (R1162_U24, U3437);
  nand ginst2164 (R1162_U240, REG1_REG_17__SCAN_IN, R1162_U49);
  nand ginst2165 (R1162_U241, R1162_U239, R1162_U240);
  nand ginst2166 (R1162_U242, R1162_U88, R1162_U89);
  nand ginst2167 (R1162_U243, R1162_U153, R1162_U241);
  nand ginst2168 (R1162_U244, R1162_U46, U3446);
  nand ginst2169 (R1162_U245, REG1_REG_16__SCAN_IN, R1162_U47);
  nand ginst2170 (R1162_U246, R1162_U46, U3446);
  nand ginst2171 (R1162_U247, REG1_REG_16__SCAN_IN, R1162_U47);
  nand ginst2172 (R1162_U248, R1162_U246, R1162_U247);
  nand ginst2173 (R1162_U249, R1162_U90, R1162_U91);
  nand ginst2174 (R1162_U25, R1162_U120, R1162_U121);
  nand ginst2175 (R1162_U250, R1162_U149, R1162_U248);
  nand ginst2176 (R1162_U251, REG1_REG_15__SCAN_IN, R1162_U43);
  nand ginst2177 (R1162_U252, R1162_U146, R1162_U45);
  nand ginst2178 (R1162_U253, REG1_REG_15__SCAN_IN, R1162_U43);
  nand ginst2179 (R1162_U254, R1162_U252, R1162_U253);
  nand ginst2180 (R1162_U255, R1162_U251, R1162_U252, R1162_U44);
  nand ginst2181 (R1162_U256, R1162_U254, U3447);
  nand ginst2182 (R1162_U257, REG1_REG_14__SCAN_IN, R1162_U40);
  nand ginst2183 (R1162_U258, R1162_U143, R1162_U42);
  nand ginst2184 (R1162_U259, REG1_REG_14__SCAN_IN, R1162_U40);
  not ginst2185 (R1162_U26, U3436);
  nand ginst2186 (R1162_U260, R1162_U258, R1162_U259);
  nand ginst2187 (R1162_U261, R1162_U257, R1162_U258, R1162_U41);
  nand ginst2188 (R1162_U262, R1162_U260, U3448);
  nand ginst2189 (R1162_U263, REG1_REG_13__SCAN_IN, R1162_U37);
  nand ginst2190 (R1162_U264, R1162_U140, R1162_U39);
  nand ginst2191 (R1162_U265, REG1_REG_13__SCAN_IN, R1162_U37);
  nand ginst2192 (R1162_U266, R1162_U264, R1162_U265);
  nand ginst2193 (R1162_U267, R1162_U263, R1162_U264, R1162_U38);
  nand ginst2194 (R1162_U268, R1162_U266, U3449);
  nand ginst2195 (R1162_U269, R1162_U35, U3450);
  not ginst2196 (R1162_U27, REG1_REG_8__SCAN_IN);
  nand ginst2197 (R1162_U270, REG1_REG_12__SCAN_IN, R1162_U36);
  nand ginst2198 (R1162_U271, R1162_U35, U3450);
  nand ginst2199 (R1162_U272, REG1_REG_12__SCAN_IN, R1162_U36);
  nand ginst2200 (R1162_U273, R1162_U271, R1162_U272);
  nand ginst2201 (R1162_U274, R1162_U92, R1162_U93);
  nand ginst2202 (R1162_U275, R1162_U136, R1162_U273);
  nand ginst2203 (R1162_U276, R1162_U33, U3451);
  nand ginst2204 (R1162_U277, REG1_REG_11__SCAN_IN, R1162_U34);
  nand ginst2205 (R1162_U278, R1162_U33, U3451);
  nand ginst2206 (R1162_U279, REG1_REG_11__SCAN_IN, R1162_U34);
  not ginst2207 (R1162_U28, U3435);
  nand ginst2208 (R1162_U280, R1162_U278, R1162_U279);
  nand ginst2209 (R1162_U281, R1162_U94, R1162_U95);
  nand ginst2210 (R1162_U282, R1162_U132, R1162_U280);
  nand ginst2211 (R1162_U283, REG1_REG_10__SCAN_IN, R1162_U30);
  nand ginst2212 (R1162_U284, R1162_U129, R1162_U32);
  nand ginst2213 (R1162_U285, REG1_REG_10__SCAN_IN, R1162_U30);
  nand ginst2214 (R1162_U286, R1162_U284, R1162_U285);
  nand ginst2215 (R1162_U287, R1162_U283, R1162_U284, R1162_U31);
  nand ginst2216 (R1162_U288, R1162_U286, U3452);
  nand ginst2217 (R1162_U289, R1162_U6, U3453);
  not ginst2218 (R1162_U29, REG1_REG_9__SCAN_IN);
  nand ginst2219 (R1162_U290, REG1_REG_0__SCAN_IN, R1162_U7);
  nand ginst2220 (R1162_U30, R1162_U127, R1162_U128);
  not ginst2221 (R1162_U31, U3452);
  not ginst2222 (R1162_U32, REG1_REG_10__SCAN_IN);
  not ginst2223 (R1162_U33, REG1_REG_11__SCAN_IN);
  not ginst2224 (R1162_U34, U3451);
  not ginst2225 (R1162_U35, REG1_REG_12__SCAN_IN);
  not ginst2226 (R1162_U36, U3450);
  nand ginst2227 (R1162_U37, R1162_U138, R1162_U139);
  not ginst2228 (R1162_U38, U3449);
  not ginst2229 (R1162_U39, REG1_REG_13__SCAN_IN);
  and ginst2230 (R1162_U4, R1162_U161, R1162_U165);
  nand ginst2231 (R1162_U40, R1162_U141, R1162_U142);
  not ginst2232 (R1162_U41, U3448);
  not ginst2233 (R1162_U42, REG1_REG_14__SCAN_IN);
  nand ginst2234 (R1162_U43, R1162_U144, R1162_U145);
  not ginst2235 (R1162_U44, U3447);
  not ginst2236 (R1162_U45, REG1_REG_15__SCAN_IN);
  not ginst2237 (R1162_U46, REG1_REG_16__SCAN_IN);
  not ginst2238 (R1162_U47, U3446);
  not ginst2239 (R1162_U48, REG1_REG_17__SCAN_IN);
  not ginst2240 (R1162_U49, U3445);
  nand ginst2241 (R1162_U5, R1162_U166, R1162_U84);
  not ginst2242 (R1162_U50, REG1_REG_18__SCAN_IN);
  not ginst2243 (R1162_U51, U3444);
  nand ginst2244 (R1162_U52, R1162_U155, R1162_U156);
  nand ginst2245 (R1162_U53, R1162_U289, R1162_U290);
  nand ginst2246 (R1162_U54, R1162_U172, R1162_U173);
  nand ginst2247 (R1162_U55, R1162_U178, R1162_U179);
  nand ginst2248 (R1162_U56, R1162_U185, R1162_U186);
  nand ginst2249 (R1162_U57, R1162_U192, R1162_U193);
  nand ginst2250 (R1162_U58, R1162_U198, R1162_U199);
  nand ginst2251 (R1162_U59, R1162_U205, R1162_U206);
  not ginst2252 (R1162_U6, REG1_REG_0__SCAN_IN);
  nand ginst2253 (R1162_U60, R1162_U211, R1162_U212);
  nand ginst2254 (R1162_U61, R1162_U218, R1162_U219);
  nand ginst2255 (R1162_U62, R1162_U235, R1162_U236);
  nand ginst2256 (R1162_U63, R1162_U242, R1162_U243);
  nand ginst2257 (R1162_U64, R1162_U249, R1162_U250);
  nand ginst2258 (R1162_U65, R1162_U255, R1162_U256);
  nand ginst2259 (R1162_U66, R1162_U261, R1162_U262);
  nand ginst2260 (R1162_U67, R1162_U267, R1162_U268);
  nand ginst2261 (R1162_U68, R1162_U274, R1162_U275);
  nand ginst2262 (R1162_U69, R1162_U281, R1162_U282);
  not ginst2263 (R1162_U7, U3453);
  nand ginst2264 (R1162_U70, R1162_U287, R1162_U288);
  and ginst2265 (R1162_U71, R1162_U160, R1162_U225, R1162_U226);
  and ginst2266 (R1162_U72, R1162_U164, R1162_U229);
  and ginst2267 (R1162_U73, R1162_U167, R1162_U168);
  nand ginst2268 (R1162_U74, R1162_U123, R1162_U124);
  and ginst2269 (R1162_U75, R1162_U180, R1162_U181);
  nand ginst2270 (R1162_U76, R1162_U116, R1162_U117);
  and ginst2271 (R1162_U77, R1162_U187, R1162_U188);
  nand ginst2272 (R1162_U78, R1162_U112, R1162_U113);
  and ginst2273 (R1162_U79, R1162_U200, R1162_U201);
  not ginst2274 (R1162_U8, U3443);
  nand ginst2275 (R1162_U80, R1162_U105, R1162_U106);
  and ginst2276 (R1162_U81, R1162_U213, R1162_U214);
  nand ginst2277 (R1162_U82, R1162_U83, R1162_U99);
  nand ginst2278 (R1162_U83, REG1_REG_1__SCAN_IN, R1162_U97);
  and ginst2279 (R1162_U84, R1162_U223, R1162_U224);
  not ginst2280 (R1162_U85, U3461);
  not ginst2281 (R1162_U86, REG1_REG_19__SCAN_IN);
  and ginst2282 (R1162_U87, R1162_U230, R1162_U231);
  and ginst2283 (R1162_U88, R1162_U237, R1162_U238);
  nand ginst2284 (R1162_U89, R1162_U151, R1162_U152);
  nand ginst2285 (R1162_U9, REG1_REG_0__SCAN_IN, U3453);
  and ginst2286 (R1162_U90, R1162_U244, R1162_U245);
  nand ginst2287 (R1162_U91, R1162_U147, R1162_U148);
  and ginst2288 (R1162_U92, R1162_U269, R1162_U270);
  nand ginst2289 (R1162_U93, R1162_U134, R1162_U135);
  and ginst2290 (R1162_U94, R1162_U276, R1162_U277);
  nand ginst2291 (R1162_U95, R1162_U130, R1162_U131);
  not ginst2292 (R1162_U96, R1162_U83);
  not ginst2293 (R1162_U97, R1162_U9);
  nand ginst2294 (R1162_U98, R1162_U10, R1162_U9);
  nand ginst2295 (R1162_U99, R1162_U98, U3443);
  and ginst2296 (R1165_U10, R1165_U256, R1165_U6);
  nand ginst2297 (R1165_U100, R1165_U522, R1165_U523);
  nand ginst2298 (R1165_U101, R1165_U527, R1165_U528);
  nand ginst2299 (R1165_U102, R1165_U534, R1165_U535);
  nand ginst2300 (R1165_U103, R1165_U541, R1165_U542);
  nand ginst2301 (R1165_U104, R1165_U548, R1165_U549);
  nand ginst2302 (R1165_U105, R1165_U555, R1165_U556);
  nand ginst2303 (R1165_U106, R1165_U560, R1165_U561);
  nand ginst2304 (R1165_U107, R1165_U567, R1165_U568);
  nand ginst2305 (R1165_U108, R1165_U574, R1165_U575);
  nand ginst2306 (R1165_U109, R1165_U581, R1165_U582);
  and ginst2307 (R1165_U11, R1165_U223, R1165_U5);
  nand ginst2308 (R1165_U110, R1165_U588, R1165_U589);
  nand ginst2309 (R1165_U111, R1165_U595, R1165_U596);
  nand ginst2310 (R1165_U112, R1165_U600, R1165_U601);
  nand ginst2311 (R1165_U113, R1165_U607, R1165_U608);
  and ginst2312 (R1165_U114, R1165_U209, R1165_U71);
  and ginst2313 (R1165_U115, R1165_U218, R1165_U219);
  and ginst2314 (R1165_U116, R1165_U11, R1165_U231);
  and ginst2315 (R1165_U117, R1165_U232, R1165_U362);
  and ginst2316 (R1165_U118, R1165_U21, R1165_U420, R1165_U421);
  and ginst2317 (R1165_U119, R1165_U237, R1165_U5);
  and ginst2318 (R1165_U12, R1165_U340, R1165_U343);
  and ginst2319 (R1165_U120, R1165_U27, R1165_U441, R1165_U442);
  and ginst2320 (R1165_U121, R1165_U244, R1165_U4);
  and ginst2321 (R1165_U122, R1165_U203, R1165_U254);
  and ginst2322 (R1165_U123, R1165_U10, R1165_U249);
  and ginst2323 (R1165_U124, R1165_U258, R1165_U363);
  and ginst2324 (R1165_U125, R1165_U271, R1165_U272);
  and ginst2325 (R1165_U126, R1165_U284, R1165_U8);
  and ginst2326 (R1165_U127, R1165_U204, R1165_U282);
  and ginst2327 (R1165_U128, R1165_U302, R1165_U9);
  and ginst2328 (R1165_U129, R1165_U205, R1165_U300);
  and ginst2329 (R1165_U13, R1165_U331, R1165_U334);
  and ginst2330 (R1165_U130, R1165_U305, R1165_U308);
  nand ginst2331 (R1165_U131, R1165_U502, R1165_U503);
  and ginst2332 (R1165_U132, R1165_U205, R1165_U517, R1165_U518);
  and ginst2333 (R1165_U133, R1165_U205, R1165_U56);
  and ginst2334 (R1165_U134, R1165_U317, R1165_U9);
  and ginst2335 (R1165_U135, R1165_U204, R1165_U543, R1165_U544);
  and ginst2336 (R1165_U136, R1165_U326, R1165_U8);
  and ginst2337 (R1165_U137, R1165_U37, R1165_U569, R1165_U570);
  and ginst2338 (R1165_U138, R1165_U333, R1165_U7);
  and ginst2339 (R1165_U139, R1165_U203, R1165_U590, R1165_U591);
  and ginst2340 (R1165_U14, R1165_U324, R1165_U327);
  and ginst2341 (R1165_U140, R1165_U342, R1165_U6);
  nand ginst2342 (R1165_U141, R1165_U609, R1165_U610);
  not ginst2343 (R1165_U142, U3198);
  and ginst2344 (R1165_U143, R1165_U379, R1165_U380);
  not ginst2345 (R1165_U144, U3203);
  not ginst2346 (R1165_U145, U3206);
  not ginst2347 (R1165_U146, U3207);
  not ginst2348 (R1165_U147, U3204);
  not ginst2349 (R1165_U148, U3205);
  not ginst2350 (R1165_U149, U3199);
  and ginst2351 (R1165_U15, R1165_U315, R1165_U318);
  not ginst2352 (R1165_U150, U3202);
  not ginst2353 (R1165_U151, U3200);
  not ginst2354 (R1165_U152, U3201);
  nand ginst2355 (R1165_U153, R1165_U117, R1165_U368);
  and ginst2356 (R1165_U154, R1165_U413, R1165_U414);
  nand ginst2357 (R1165_U155, R1165_U361, R1165_U366);
  and ginst2358 (R1165_U156, R1165_U427, R1165_U428);
  nand ginst2359 (R1165_U157, R1165_U354, R1165_U370);
  and ginst2360 (R1165_U158, R1165_U434, R1165_U435);
  nand ginst2361 (R1165_U159, R1165_U115, R1165_U220);
  and ginst2362 (R1165_U16, R1165_U242, R1165_U245);
  not ginst2363 (R1165_U160, U3180);
  not ginst2364 (R1165_U161, U3196);
  not ginst2365 (R1165_U162, U3194);
  not ginst2366 (R1165_U163, U3195);
  not ginst2367 (R1165_U164, U3197);
  not ginst2368 (R1165_U165, U3193);
  not ginst2369 (R1165_U166, U3192);
  not ginst2370 (R1165_U167, U3190);
  not ginst2371 (R1165_U168, U3191);
  not ginst2372 (R1165_U169, U3189);
  and ginst2373 (R1165_U17, R1165_U235, R1165_U238);
  not ginst2374 (R1165_U170, U3186);
  not ginst2375 (R1165_U171, U3187);
  not ginst2376 (R1165_U172, U3188);
  not ginst2377 (R1165_U173, U3185);
  not ginst2378 (R1165_U174, U3184);
  not ginst2379 (R1165_U175, U3181);
  not ginst2380 (R1165_U176, U3182);
  not ginst2381 (R1165_U177, U3183);
  not ginst2382 (R1165_U178, U3150);
  not ginst2383 (R1165_U179, U3179);
  not ginst2384 (R1165_U18, U3208);
  and ginst2385 (R1165_U180, R1165_U510, R1165_U511);
  nand ginst2386 (R1165_U181, R1165_U304, R1165_U305);
  nand ginst2387 (R1165_U182, R1165_U311, R1165_U56);
  nand ginst2388 (R1165_U183, R1165_U294, R1165_U295);
  and ginst2389 (R1165_U184, R1165_U529, R1165_U530);
  nand ginst2390 (R1165_U185, R1165_U290, R1165_U291);
  and ginst2391 (R1165_U186, R1165_U536, R1165_U537);
  nand ginst2392 (R1165_U187, R1165_U286, R1165_U287);
  and ginst2393 (R1165_U188, R1165_U550, R1165_U551);
  nand ginst2394 (R1165_U189, R1165_U210, R1165_U31);
  not ginst2395 (R1165_U19, U3170);
  nand ginst2396 (R1165_U190, R1165_U276, R1165_U277);
  and ginst2397 (R1165_U191, R1165_U562, R1165_U563);
  nand ginst2398 (R1165_U192, R1165_U125, R1165_U273);
  and ginst2399 (R1165_U193, R1165_U576, R1165_U577);
  nand ginst2400 (R1165_U194, R1165_U260, R1165_U261);
  and ginst2401 (R1165_U195, R1165_U583, R1165_U584);
  nand ginst2402 (R1165_U196, R1165_U124, R1165_U374);
  nand ginst2403 (R1165_U197, R1165_U372, R1165_U44);
  and ginst2404 (R1165_U198, R1165_U602, R1165_U603);
  nand ginst2405 (R1165_U199, R1165_U201, R1165_U247, R1165_U355);
  not ginst2406 (R1165_U20, U3172);
  nand ginst2407 (R1165_U200, R1165_U181, R1165_U310);
  nand ginst2408 (R1165_U201, R1165_U153, R1165_U62);
  not ginst2409 (R1165_U202, R1165_U27);
  nand ginst2410 (R1165_U203, R1165_U74, U3166);
  nand ginst2411 (R1165_U204, R1165_U83, U3158);
  nand ginst2412 (R1165_U205, R1165_U88, U3153);
  not ginst2413 (R1165_U206, R1165_U41);
  not ginst2414 (R1165_U207, R1165_U50);
  not ginst2415 (R1165_U208, R1165_U56);
  or ginst2416 (R1165_U209, U3178, U3208);
  nand ginst2417 (R1165_U21, R1165_U64, U3172);
  nand ginst2418 (R1165_U210, R1165_U209, R1165_U71);
  not ginst2419 (R1165_U211, R1165_U31);
  not ginst2420 (R1165_U212, R1165_U189);
  nand ginst2421 (R1165_U213, R1165_U70, U3177);
  not ginst2422 (R1165_U214, R1165_U35);
  nand ginst2423 (R1165_U215, R1165_U28, R1165_U395);
  nand ginst2424 (R1165_U216, R1165_U26, R1165_U398);
  nand ginst2425 (R1165_U217, R1165_U27, R1165_U28);
  nand ginst2426 (R1165_U218, R1165_U217, R1165_U69);
  nand ginst2427 (R1165_U219, R1165_U202, U3175);
  not ginst2428 (R1165_U22, U3171);
  nand ginst2429 (R1165_U220, R1165_U35, R1165_U4);
  not ginst2430 (R1165_U221, R1165_U159);
  nand ginst2431 (R1165_U222, R1165_U25, R1165_U386);
  nand ginst2432 (R1165_U223, R1165_U23, R1165_U404);
  not ginst2433 (R1165_U224, R1165_U24);
  nand ginst2434 (R1165_U225, R1165_U22, R1165_U407);
  nand ginst2435 (R1165_U226, R1165_U20, R1165_U410);
  not ginst2436 (R1165_U227, R1165_U21);
  nand ginst2437 (R1165_U228, R1165_U21, R1165_U22);
  nand ginst2438 (R1165_U229, R1165_U228, R1165_U65);
  not ginst2439 (R1165_U23, U3173);
  nand ginst2440 (R1165_U230, R1165_U227, U3171);
  nand ginst2441 (R1165_U231, R1165_U19, R1165_U401);
  nand ginst2442 (R1165_U232, R1165_U63, U3170);
  nand ginst2443 (R1165_U233, R1165_U20, R1165_U410);
  nand ginst2444 (R1165_U234, R1165_U233, R1165_U34);
  nand ginst2445 (R1165_U235, R1165_U118, R1165_U234);
  nand ginst2446 (R1165_U236, R1165_U21, R1165_U365);
  nand ginst2447 (R1165_U237, R1165_U65, U3171);
  nand ginst2448 (R1165_U238, R1165_U119, R1165_U236);
  nand ginst2449 (R1165_U239, R1165_U20, R1165_U410);
  nand ginst2450 (R1165_U24, R1165_U66, U3173);
  nand ginst2451 (R1165_U240, R1165_U26, R1165_U398);
  nand ginst2452 (R1165_U241, R1165_U240, R1165_U35);
  nand ginst2453 (R1165_U242, R1165_U120, R1165_U241);
  nand ginst2454 (R1165_U243, R1165_U214, R1165_U27);
  nand ginst2455 (R1165_U244, R1165_U69, U3175);
  nand ginst2456 (R1165_U245, R1165_U121, R1165_U243);
  nand ginst2457 (R1165_U246, R1165_U26, R1165_U398);
  nand ginst2458 (R1165_U247, R1165_U153, U3169);
  not ginst2459 (R1165_U248, R1165_U199);
  nand ginst2460 (R1165_U249, R1165_U43, R1165_U462);
  not ginst2461 (R1165_U25, U3174);
  not ginst2462 (R1165_U250, R1165_U44);
  nand ginst2463 (R1165_U251, R1165_U42, R1165_U456);
  nand ginst2464 (R1165_U252, R1165_U39, R1165_U459);
  nand ginst2465 (R1165_U253, R1165_U206, R1165_U6);
  nand ginst2466 (R1165_U254, R1165_U75, U3165);
  nand ginst2467 (R1165_U255, R1165_U122, R1165_U253);
  nand ginst2468 (R1165_U256, R1165_U40, R1165_U453);
  nand ginst2469 (R1165_U257, R1165_U42, R1165_U456);
  nand ginst2470 (R1165_U258, R1165_U255, R1165_U257);
  nand ginst2471 (R1165_U259, R1165_U45, R1165_U465);
  not ginst2472 (R1165_U26, U3176);
  nand ginst2473 (R1165_U260, R1165_U196, R1165_U259);
  nand ginst2474 (R1165_U261, R1165_U78, U3164);
  not ginst2475 (R1165_U262, R1165_U194);
  nand ginst2476 (R1165_U263, R1165_U46, R1165_U468);
  nand ginst2477 (R1165_U264, R1165_U194, R1165_U263);
  nand ginst2478 (R1165_U265, R1165_U79, U3163);
  not ginst2479 (R1165_U266, R1165_U60);
  nand ginst2480 (R1165_U267, R1165_U38, R1165_U471);
  nand ginst2481 (R1165_U268, R1165_U36, R1165_U474);
  not ginst2482 (R1165_U269, R1165_U37);
  nand ginst2483 (R1165_U27, R1165_U68, U3176);
  nand ginst2484 (R1165_U270, R1165_U37, R1165_U38);
  nand ginst2485 (R1165_U271, R1165_U270, R1165_U73);
  nand ginst2486 (R1165_U272, R1165_U269, U3161);
  nand ginst2487 (R1165_U273, R1165_U60, R1165_U7);
  not ginst2488 (R1165_U274, R1165_U192);
  nand ginst2489 (R1165_U275, R1165_U47, R1165_U477);
  nand ginst2490 (R1165_U276, R1165_U192, R1165_U275);
  nand ginst2491 (R1165_U277, R1165_U80, U3160);
  not ginst2492 (R1165_U278, R1165_U190);
  nand ginst2493 (R1165_U279, R1165_U480, R1165_U51);
  not ginst2494 (R1165_U28, U3175);
  nand ginst2495 (R1165_U280, R1165_U48, R1165_U483);
  nand ginst2496 (R1165_U281, R1165_U207, R1165_U8);
  nand ginst2497 (R1165_U282, R1165_U82, U3157);
  nand ginst2498 (R1165_U283, R1165_U127, R1165_U281);
  nand ginst2499 (R1165_U284, R1165_U486, R1165_U49);
  nand ginst2500 (R1165_U285, R1165_U480, R1165_U51);
  nand ginst2501 (R1165_U286, R1165_U126, R1165_U190);
  nand ginst2502 (R1165_U287, R1165_U283, R1165_U285);
  not ginst2503 (R1165_U288, R1165_U187);
  nand ginst2504 (R1165_U289, R1165_U489, R1165_U52);
  not ginst2505 (R1165_U29, U3177);
  nand ginst2506 (R1165_U290, R1165_U187, R1165_U289);
  nand ginst2507 (R1165_U291, R1165_U84, U3156);
  not ginst2508 (R1165_U292, R1165_U185);
  nand ginst2509 (R1165_U293, R1165_U492, R1165_U53);
  nand ginst2510 (R1165_U294, R1165_U185, R1165_U293);
  nand ginst2511 (R1165_U295, R1165_U85, U3155);
  not ginst2512 (R1165_U296, R1165_U183);
  nand ginst2513 (R1165_U297, R1165_U495, R1165_U57);
  nand ginst2514 (R1165_U298, R1165_U498, R1165_U54);
  nand ginst2515 (R1165_U299, R1165_U208, R1165_U9);
  not ginst2516 (R1165_U30, U3178);
  nand ginst2517 (R1165_U300, R1165_U87, U3152);
  nand ginst2518 (R1165_U301, R1165_U129, R1165_U299);
  nand ginst2519 (R1165_U302, R1165_U501, R1165_U55);
  nand ginst2520 (R1165_U303, R1165_U495, R1165_U57);
  nand ginst2521 (R1165_U304, R1165_U128, R1165_U183);
  nand ginst2522 (R1165_U305, R1165_U301, R1165_U303);
  not ginst2523 (R1165_U306, R1165_U181);
  nand ginst2524 (R1165_U307, R1165_U450, R1165_U58);
  nand ginst2525 (R1165_U308, R1165_U89, U3151);
  nand ginst2526 (R1165_U309, R1165_U89, U3151);
  nand ginst2527 (R1165_U31, U3178, U3208);
  nand ginst2528 (R1165_U310, R1165_U450, R1165_U58);
  nand ginst2529 (R1165_U311, R1165_U183, R1165_U302);
  not ginst2530 (R1165_U312, R1165_U182);
  nand ginst2531 (R1165_U313, R1165_U498, R1165_U54);
  nand ginst2532 (R1165_U314, R1165_U182, R1165_U313);
  nand ginst2533 (R1165_U315, R1165_U132, R1165_U314);
  nand ginst2534 (R1165_U316, R1165_U133, R1165_U311);
  nand ginst2535 (R1165_U317, R1165_U87, U3152);
  nand ginst2536 (R1165_U318, R1165_U134, R1165_U316);
  nand ginst2537 (R1165_U319, R1165_U498, R1165_U54);
  not ginst2538 (R1165_U32, U3169);
  nand ginst2539 (R1165_U320, R1165_U190, R1165_U284);
  not ginst2540 (R1165_U321, R1165_U59);
  nand ginst2541 (R1165_U322, R1165_U48, R1165_U483);
  nand ginst2542 (R1165_U323, R1165_U322, R1165_U59);
  nand ginst2543 (R1165_U324, R1165_U135, R1165_U323);
  nand ginst2544 (R1165_U325, R1165_U204, R1165_U321);
  nand ginst2545 (R1165_U326, R1165_U82, U3157);
  nand ginst2546 (R1165_U327, R1165_U136, R1165_U325);
  nand ginst2547 (R1165_U328, R1165_U48, R1165_U483);
  nand ginst2548 (R1165_U329, R1165_U36, R1165_U474);
  nand ginst2549 (R1165_U33, R1165_U229, R1165_U230, R1165_U360);
  nand ginst2550 (R1165_U330, R1165_U329, R1165_U60);
  nand ginst2551 (R1165_U331, R1165_U137, R1165_U330);
  nand ginst2552 (R1165_U332, R1165_U266, R1165_U37);
  nand ginst2553 (R1165_U333, R1165_U73, U3161);
  nand ginst2554 (R1165_U334, R1165_U138, R1165_U332);
  nand ginst2555 (R1165_U335, R1165_U36, R1165_U474);
  nand ginst2556 (R1165_U336, R1165_U197, R1165_U256);
  not ginst2557 (R1165_U337, R1165_U61);
  nand ginst2558 (R1165_U338, R1165_U39, R1165_U459);
  nand ginst2559 (R1165_U339, R1165_U338, R1165_U61);
  nand ginst2560 (R1165_U34, R1165_U24, R1165_U364);
  nand ginst2561 (R1165_U340, R1165_U139, R1165_U339);
  nand ginst2562 (R1165_U341, R1165_U203, R1165_U337);
  nand ginst2563 (R1165_U342, R1165_U75, U3165);
  nand ginst2564 (R1165_U343, R1165_U140, R1165_U341);
  nand ginst2565 (R1165_U344, R1165_U39, R1165_U459);
  nand ginst2566 (R1165_U345, R1165_U21, R1165_U239);
  nand ginst2567 (R1165_U346, R1165_U246, R1165_U27);
  nand ginst2568 (R1165_U347, R1165_U205, R1165_U319);
  nand ginst2569 (R1165_U348, R1165_U302, R1165_U56);
  nand ginst2570 (R1165_U349, R1165_U204, R1165_U328);
  nand ginst2571 (R1165_U35, R1165_U213, R1165_U357, R1165_U358);
  nand ginst2572 (R1165_U350, R1165_U284, R1165_U50);
  nand ginst2573 (R1165_U351, R1165_U335, R1165_U37);
  nand ginst2574 (R1165_U352, R1165_U203, R1165_U344);
  nand ginst2575 (R1165_U353, R1165_U256, R1165_U41);
  nand ginst2576 (R1165_U354, R1165_U67, U3174);
  nand ginst2577 (R1165_U355, R1165_U62, U3169);
  nand ginst2578 (R1165_U356, R1165_U130, R1165_U304);
  nand ginst2579 (R1165_U357, R1165_U114, R1165_U359);
  nand ginst2580 (R1165_U358, R1165_U211, R1165_U359);
  nand ginst2581 (R1165_U359, R1165_U29, R1165_U389);
  not ginst2582 (R1165_U36, U3162);
  nand ginst2583 (R1165_U360, R1165_U224, R1165_U5);
  not ginst2584 (R1165_U361, R1165_U33);
  nand ginst2585 (R1165_U362, R1165_U231, R1165_U33);
  nand ginst2586 (R1165_U363, R1165_U10, R1165_U250);
  nand ginst2587 (R1165_U364, R1165_U157, R1165_U223);
  not ginst2588 (R1165_U365, R1165_U34);
  nand ginst2589 (R1165_U366, R1165_U11, R1165_U157);
  not ginst2590 (R1165_U367, R1165_U155);
  nand ginst2591 (R1165_U368, R1165_U116, R1165_U157);
  not ginst2592 (R1165_U369, R1165_U153);
  nand ginst2593 (R1165_U37, R1165_U72, U3162);
  nand ginst2594 (R1165_U370, R1165_U159, R1165_U222);
  not ginst2595 (R1165_U371, R1165_U157);
  nand ginst2596 (R1165_U372, R1165_U199, R1165_U249);
  not ginst2597 (R1165_U373, R1165_U197);
  nand ginst2598 (R1165_U374, R1165_U123, R1165_U199);
  not ginst2599 (R1165_U375, R1165_U196);
  nand ginst2600 (R1165_U376, R1165_U142, U3208);
  nand ginst2601 (R1165_U377, R1165_U18, U3198);
  not ginst2602 (R1165_U378, R1165_U62);
  nand ginst2603 (R1165_U379, R1165_U378, U3169);
  not ginst2604 (R1165_U38, U3161);
  nand ginst2605 (R1165_U380, R1165_U32, R1165_U62);
  nand ginst2606 (R1165_U381, R1165_U378, U3169);
  nand ginst2607 (R1165_U382, R1165_U32, R1165_U62);
  nand ginst2608 (R1165_U383, R1165_U381, R1165_U382);
  nand ginst2609 (R1165_U384, R1165_U144, U3208);
  nand ginst2610 (R1165_U385, R1165_U18, U3203);
  not ginst2611 (R1165_U386, R1165_U67);
  nand ginst2612 (R1165_U387, R1165_U145, U3208);
  nand ginst2613 (R1165_U388, R1165_U18, U3206);
  not ginst2614 (R1165_U389, R1165_U70);
  not ginst2615 (R1165_U39, U3166);
  nand ginst2616 (R1165_U390, R1165_U146, U3208);
  nand ginst2617 (R1165_U391, R1165_U18, U3207);
  not ginst2618 (R1165_U392, R1165_U71);
  nand ginst2619 (R1165_U393, R1165_U147, U3208);
  nand ginst2620 (R1165_U394, R1165_U18, U3204);
  not ginst2621 (R1165_U395, R1165_U69);
  nand ginst2622 (R1165_U396, R1165_U148, U3208);
  nand ginst2623 (R1165_U397, R1165_U18, U3205);
  not ginst2624 (R1165_U398, R1165_U68);
  nand ginst2625 (R1165_U399, R1165_U149, U3208);
  and ginst2626 (R1165_U4, R1165_U215, R1165_U216);
  not ginst2627 (R1165_U40, U3167);
  nand ginst2628 (R1165_U400, R1165_U18, U3199);
  not ginst2629 (R1165_U401, R1165_U63);
  nand ginst2630 (R1165_U402, R1165_U150, U3208);
  nand ginst2631 (R1165_U403, R1165_U18, U3202);
  not ginst2632 (R1165_U404, R1165_U66);
  nand ginst2633 (R1165_U405, R1165_U151, U3208);
  nand ginst2634 (R1165_U406, R1165_U18, U3200);
  not ginst2635 (R1165_U407, R1165_U65);
  nand ginst2636 (R1165_U408, R1165_U152, U3208);
  nand ginst2637 (R1165_U409, R1165_U18, U3201);
  nand ginst2638 (R1165_U41, R1165_U76, U3167);
  not ginst2639 (R1165_U410, R1165_U64);
  nand ginst2640 (R1165_U411, R1165_U143, R1165_U153);
  nand ginst2641 (R1165_U412, R1165_U369, R1165_U383);
  nand ginst2642 (R1165_U413, R1165_U401, U3170);
  nand ginst2643 (R1165_U414, R1165_U19, R1165_U63);
  nand ginst2644 (R1165_U415, R1165_U401, U3170);
  nand ginst2645 (R1165_U416, R1165_U19, R1165_U63);
  nand ginst2646 (R1165_U417, R1165_U415, R1165_U416);
  nand ginst2647 (R1165_U418, R1165_U154, R1165_U155);
  nand ginst2648 (R1165_U419, R1165_U367, R1165_U417);
  not ginst2649 (R1165_U42, U3165);
  nand ginst2650 (R1165_U420, R1165_U407, U3171);
  nand ginst2651 (R1165_U421, R1165_U22, R1165_U65);
  nand ginst2652 (R1165_U422, R1165_U410, U3172);
  nand ginst2653 (R1165_U423, R1165_U20, R1165_U64);
  nand ginst2654 (R1165_U424, R1165_U422, R1165_U423);
  nand ginst2655 (R1165_U425, R1165_U34, R1165_U345);
  nand ginst2656 (R1165_U426, R1165_U365, R1165_U424);
  nand ginst2657 (R1165_U427, R1165_U404, U3173);
  nand ginst2658 (R1165_U428, R1165_U23, R1165_U66);
  nand ginst2659 (R1165_U429, R1165_U404, U3173);
  not ginst2660 (R1165_U43, U3168);
  nand ginst2661 (R1165_U430, R1165_U23, R1165_U66);
  nand ginst2662 (R1165_U431, R1165_U429, R1165_U430);
  nand ginst2663 (R1165_U432, R1165_U156, R1165_U157);
  nand ginst2664 (R1165_U433, R1165_U371, R1165_U431);
  nand ginst2665 (R1165_U434, R1165_U386, U3174);
  nand ginst2666 (R1165_U435, R1165_U25, R1165_U67);
  nand ginst2667 (R1165_U436, R1165_U386, U3174);
  nand ginst2668 (R1165_U437, R1165_U25, R1165_U67);
  nand ginst2669 (R1165_U438, R1165_U436, R1165_U437);
  nand ginst2670 (R1165_U439, R1165_U158, R1165_U159);
  nand ginst2671 (R1165_U44, R1165_U77, U3168);
  nand ginst2672 (R1165_U440, R1165_U221, R1165_U438);
  nand ginst2673 (R1165_U441, R1165_U395, U3175);
  nand ginst2674 (R1165_U442, R1165_U28, R1165_U69);
  nand ginst2675 (R1165_U443, R1165_U398, U3176);
  nand ginst2676 (R1165_U444, R1165_U26, R1165_U68);
  nand ginst2677 (R1165_U445, R1165_U443, R1165_U444);
  nand ginst2678 (R1165_U446, R1165_U346, R1165_U35);
  nand ginst2679 (R1165_U447, R1165_U214, R1165_U445);
  nand ginst2680 (R1165_U448, R1165_U160, U3208);
  nand ginst2681 (R1165_U449, R1165_U18, U3180);
  not ginst2682 (R1165_U45, U3164);
  not ginst2683 (R1165_U450, R1165_U89);
  nand ginst2684 (R1165_U451, R1165_U161, U3208);
  nand ginst2685 (R1165_U452, R1165_U18, U3196);
  not ginst2686 (R1165_U453, R1165_U76);
  nand ginst2687 (R1165_U454, R1165_U162, U3208);
  nand ginst2688 (R1165_U455, R1165_U18, U3194);
  not ginst2689 (R1165_U456, R1165_U75);
  nand ginst2690 (R1165_U457, R1165_U163, U3208);
  nand ginst2691 (R1165_U458, R1165_U18, U3195);
  not ginst2692 (R1165_U459, R1165_U74);
  not ginst2693 (R1165_U46, U3163);
  nand ginst2694 (R1165_U460, R1165_U164, U3208);
  nand ginst2695 (R1165_U461, R1165_U18, U3197);
  not ginst2696 (R1165_U462, R1165_U77);
  nand ginst2697 (R1165_U463, R1165_U165, U3208);
  nand ginst2698 (R1165_U464, R1165_U18, U3193);
  not ginst2699 (R1165_U465, R1165_U78);
  nand ginst2700 (R1165_U466, R1165_U166, U3208);
  nand ginst2701 (R1165_U467, R1165_U18, U3192);
  not ginst2702 (R1165_U468, R1165_U79);
  nand ginst2703 (R1165_U469, R1165_U167, U3208);
  not ginst2704 (R1165_U47, U3160);
  nand ginst2705 (R1165_U470, R1165_U18, U3190);
  not ginst2706 (R1165_U471, R1165_U73);
  nand ginst2707 (R1165_U472, R1165_U168, U3208);
  nand ginst2708 (R1165_U473, R1165_U18, U3191);
  not ginst2709 (R1165_U474, R1165_U72);
  nand ginst2710 (R1165_U475, R1165_U169, U3208);
  nand ginst2711 (R1165_U476, R1165_U18, U3189);
  not ginst2712 (R1165_U477, R1165_U80);
  nand ginst2713 (R1165_U478, R1165_U170, U3208);
  nand ginst2714 (R1165_U479, R1165_U18, U3186);
  not ginst2715 (R1165_U48, U3158);
  not ginst2716 (R1165_U480, R1165_U82);
  nand ginst2717 (R1165_U481, R1165_U171, U3208);
  nand ginst2718 (R1165_U482, R1165_U18, U3187);
  not ginst2719 (R1165_U483, R1165_U83);
  nand ginst2720 (R1165_U484, R1165_U172, U3208);
  nand ginst2721 (R1165_U485, R1165_U18, U3188);
  not ginst2722 (R1165_U486, R1165_U81);
  nand ginst2723 (R1165_U487, R1165_U173, U3208);
  nand ginst2724 (R1165_U488, R1165_U18, U3185);
  not ginst2725 (R1165_U489, R1165_U84);
  not ginst2726 (R1165_U49, U3159);
  nand ginst2727 (R1165_U490, R1165_U174, U3208);
  nand ginst2728 (R1165_U491, R1165_U18, U3184);
  not ginst2729 (R1165_U492, R1165_U85);
  nand ginst2730 (R1165_U493, R1165_U175, U3208);
  nand ginst2731 (R1165_U494, R1165_U18, U3181);
  not ginst2732 (R1165_U495, R1165_U87);
  nand ginst2733 (R1165_U496, R1165_U176, U3208);
  nand ginst2734 (R1165_U497, R1165_U18, U3182);
  not ginst2735 (R1165_U498, R1165_U88);
  nand ginst2736 (R1165_U499, R1165_U177, U3208);
  and ginst2737 (R1165_U5, R1165_U225, R1165_U226);
  nand ginst2738 (R1165_U50, R1165_U81, U3159);
  nand ginst2739 (R1165_U500, R1165_U18, U3183);
  not ginst2740 (R1165_U501, R1165_U86);
  nand ginst2741 (R1165_U502, R1165_U178, U3208);
  nand ginst2742 (R1165_U503, R1165_U18, U3150);
  not ginst2743 (R1165_U504, R1165_U131);
  nand ginst2744 (R1165_U505, R1165_U504, U3179);
  nand ginst2745 (R1165_U506, R1165_U131, R1165_U179);
  not ginst2746 (R1165_U507, R1165_U90);
  nand ginst2747 (R1165_U508, R1165_U307, R1165_U356, R1165_U507);
  nand ginst2748 (R1165_U509, R1165_U200, R1165_U309, R1165_U90);
  not ginst2749 (R1165_U51, U3157);
  nand ginst2750 (R1165_U510, R1165_U450, U3151);
  nand ginst2751 (R1165_U511, R1165_U58, R1165_U89);
  nand ginst2752 (R1165_U512, R1165_U450, U3151);
  nand ginst2753 (R1165_U513, R1165_U58, R1165_U89);
  nand ginst2754 (R1165_U514, R1165_U512, R1165_U513);
  nand ginst2755 (R1165_U515, R1165_U180, R1165_U181);
  nand ginst2756 (R1165_U516, R1165_U306, R1165_U514);
  nand ginst2757 (R1165_U517, R1165_U495, U3152);
  nand ginst2758 (R1165_U518, R1165_U57, R1165_U87);
  nand ginst2759 (R1165_U519, R1165_U498, U3153);
  not ginst2760 (R1165_U52, U3156);
  nand ginst2761 (R1165_U520, R1165_U54, R1165_U88);
  nand ginst2762 (R1165_U521, R1165_U519, R1165_U520);
  nand ginst2763 (R1165_U522, R1165_U182, R1165_U347);
  nand ginst2764 (R1165_U523, R1165_U312, R1165_U521);
  nand ginst2765 (R1165_U524, R1165_U501, U3154);
  nand ginst2766 (R1165_U525, R1165_U55, R1165_U86);
  nand ginst2767 (R1165_U526, R1165_U524, R1165_U525);
  nand ginst2768 (R1165_U527, R1165_U183, R1165_U348);
  nand ginst2769 (R1165_U528, R1165_U296, R1165_U526);
  nand ginst2770 (R1165_U529, R1165_U492, U3155);
  not ginst2771 (R1165_U53, U3155);
  nand ginst2772 (R1165_U530, R1165_U53, R1165_U85);
  nand ginst2773 (R1165_U531, R1165_U492, U3155);
  nand ginst2774 (R1165_U532, R1165_U53, R1165_U85);
  nand ginst2775 (R1165_U533, R1165_U531, R1165_U532);
  nand ginst2776 (R1165_U534, R1165_U184, R1165_U185);
  nand ginst2777 (R1165_U535, R1165_U292, R1165_U533);
  nand ginst2778 (R1165_U536, R1165_U489, U3156);
  nand ginst2779 (R1165_U537, R1165_U52, R1165_U84);
  nand ginst2780 (R1165_U538, R1165_U489, U3156);
  nand ginst2781 (R1165_U539, R1165_U52, R1165_U84);
  not ginst2782 (R1165_U54, U3153);
  nand ginst2783 (R1165_U540, R1165_U538, R1165_U539);
  nand ginst2784 (R1165_U541, R1165_U186, R1165_U187);
  nand ginst2785 (R1165_U542, R1165_U288, R1165_U540);
  nand ginst2786 (R1165_U543, R1165_U480, U3157);
  nand ginst2787 (R1165_U544, R1165_U51, R1165_U82);
  nand ginst2788 (R1165_U545, R1165_U483, U3158);
  nand ginst2789 (R1165_U546, R1165_U48, R1165_U83);
  nand ginst2790 (R1165_U547, R1165_U545, R1165_U546);
  nand ginst2791 (R1165_U548, R1165_U349, R1165_U59);
  nand ginst2792 (R1165_U549, R1165_U321, R1165_U547);
  not ginst2793 (R1165_U55, U3154);
  nand ginst2794 (R1165_U550, R1165_U389, U3177);
  nand ginst2795 (R1165_U551, R1165_U29, R1165_U70);
  nand ginst2796 (R1165_U552, R1165_U389, U3177);
  nand ginst2797 (R1165_U553, R1165_U29, R1165_U70);
  nand ginst2798 (R1165_U554, R1165_U552, R1165_U553);
  nand ginst2799 (R1165_U555, R1165_U188, R1165_U189);
  nand ginst2800 (R1165_U556, R1165_U212, R1165_U554);
  nand ginst2801 (R1165_U557, R1165_U486, U3159);
  nand ginst2802 (R1165_U558, R1165_U49, R1165_U81);
  nand ginst2803 (R1165_U559, R1165_U557, R1165_U558);
  nand ginst2804 (R1165_U56, R1165_U86, U3154);
  nand ginst2805 (R1165_U560, R1165_U190, R1165_U350);
  nand ginst2806 (R1165_U561, R1165_U278, R1165_U559);
  nand ginst2807 (R1165_U562, R1165_U477, U3160);
  nand ginst2808 (R1165_U563, R1165_U47, R1165_U80);
  nand ginst2809 (R1165_U564, R1165_U477, U3160);
  nand ginst2810 (R1165_U565, R1165_U47, R1165_U80);
  nand ginst2811 (R1165_U566, R1165_U564, R1165_U565);
  nand ginst2812 (R1165_U567, R1165_U191, R1165_U192);
  nand ginst2813 (R1165_U568, R1165_U274, R1165_U566);
  nand ginst2814 (R1165_U569, R1165_U471, U3161);
  not ginst2815 (R1165_U57, U3152);
  nand ginst2816 (R1165_U570, R1165_U38, R1165_U73);
  nand ginst2817 (R1165_U571, R1165_U474, U3162);
  nand ginst2818 (R1165_U572, R1165_U36, R1165_U72);
  nand ginst2819 (R1165_U573, R1165_U571, R1165_U572);
  nand ginst2820 (R1165_U574, R1165_U351, R1165_U60);
  nand ginst2821 (R1165_U575, R1165_U266, R1165_U573);
  nand ginst2822 (R1165_U576, R1165_U468, U3163);
  nand ginst2823 (R1165_U577, R1165_U46, R1165_U79);
  nand ginst2824 (R1165_U578, R1165_U468, U3163);
  nand ginst2825 (R1165_U579, R1165_U46, R1165_U79);
  not ginst2826 (R1165_U58, U3151);
  nand ginst2827 (R1165_U580, R1165_U578, R1165_U579);
  nand ginst2828 (R1165_U581, R1165_U193, R1165_U194);
  nand ginst2829 (R1165_U582, R1165_U262, R1165_U580);
  nand ginst2830 (R1165_U583, R1165_U465, U3164);
  nand ginst2831 (R1165_U584, R1165_U45, R1165_U78);
  nand ginst2832 (R1165_U585, R1165_U465, U3164);
  nand ginst2833 (R1165_U586, R1165_U45, R1165_U78);
  nand ginst2834 (R1165_U587, R1165_U585, R1165_U586);
  nand ginst2835 (R1165_U588, R1165_U195, R1165_U196);
  nand ginst2836 (R1165_U589, R1165_U375, R1165_U587);
  nand ginst2837 (R1165_U59, R1165_U320, R1165_U50);
  nand ginst2838 (R1165_U590, R1165_U456, U3165);
  nand ginst2839 (R1165_U591, R1165_U42, R1165_U75);
  nand ginst2840 (R1165_U592, R1165_U459, U3166);
  nand ginst2841 (R1165_U593, R1165_U39, R1165_U74);
  nand ginst2842 (R1165_U594, R1165_U592, R1165_U593);
  nand ginst2843 (R1165_U595, R1165_U352, R1165_U61);
  nand ginst2844 (R1165_U596, R1165_U337, R1165_U594);
  nand ginst2845 (R1165_U597, R1165_U453, U3167);
  nand ginst2846 (R1165_U598, R1165_U40, R1165_U76);
  nand ginst2847 (R1165_U599, R1165_U597, R1165_U598);
  and ginst2848 (R1165_U6, R1165_U251, R1165_U252);
  nand ginst2849 (R1165_U60, R1165_U264, R1165_U265);
  nand ginst2850 (R1165_U600, R1165_U197, R1165_U353);
  nand ginst2851 (R1165_U601, R1165_U373, R1165_U599);
  nand ginst2852 (R1165_U602, R1165_U462, U3168);
  nand ginst2853 (R1165_U603, R1165_U43, R1165_U77);
  nand ginst2854 (R1165_U604, R1165_U462, U3168);
  nand ginst2855 (R1165_U605, R1165_U43, R1165_U77);
  nand ginst2856 (R1165_U606, R1165_U604, R1165_U605);
  nand ginst2857 (R1165_U607, R1165_U198, R1165_U199);
  nand ginst2858 (R1165_U608, R1165_U248, R1165_U606);
  nand ginst2859 (R1165_U609, R1165_U18, U3178);
  nand ginst2860 (R1165_U61, R1165_U336, R1165_U41);
  nand ginst2861 (R1165_U610, R1165_U30, U3208);
  not ginst2862 (R1165_U611, R1165_U141);
  nand ginst2863 (R1165_U612, R1165_U611, R1165_U71);
  nand ginst2864 (R1165_U613, R1165_U141, R1165_U392);
  nand ginst2865 (R1165_U62, R1165_U376, R1165_U377);
  nand ginst2866 (R1165_U63, R1165_U399, R1165_U400);
  nand ginst2867 (R1165_U64, R1165_U408, R1165_U409);
  nand ginst2868 (R1165_U65, R1165_U405, R1165_U406);
  nand ginst2869 (R1165_U66, R1165_U402, R1165_U403);
  nand ginst2870 (R1165_U67, R1165_U384, R1165_U385);
  nand ginst2871 (R1165_U68, R1165_U396, R1165_U397);
  nand ginst2872 (R1165_U69, R1165_U393, R1165_U394);
  and ginst2873 (R1165_U7, R1165_U267, R1165_U268);
  nand ginst2874 (R1165_U70, R1165_U387, R1165_U388);
  nand ginst2875 (R1165_U71, R1165_U390, R1165_U391);
  nand ginst2876 (R1165_U72, R1165_U472, R1165_U473);
  nand ginst2877 (R1165_U73, R1165_U469, R1165_U470);
  nand ginst2878 (R1165_U74, R1165_U457, R1165_U458);
  nand ginst2879 (R1165_U75, R1165_U454, R1165_U455);
  nand ginst2880 (R1165_U76, R1165_U451, R1165_U452);
  nand ginst2881 (R1165_U77, R1165_U460, R1165_U461);
  nand ginst2882 (R1165_U78, R1165_U463, R1165_U464);
  nand ginst2883 (R1165_U79, R1165_U466, R1165_U467);
  and ginst2884 (R1165_U8, R1165_U279, R1165_U280);
  nand ginst2885 (R1165_U80, R1165_U475, R1165_U476);
  nand ginst2886 (R1165_U81, R1165_U484, R1165_U485);
  nand ginst2887 (R1165_U82, R1165_U478, R1165_U479);
  nand ginst2888 (R1165_U83, R1165_U481, R1165_U482);
  nand ginst2889 (R1165_U84, R1165_U487, R1165_U488);
  nand ginst2890 (R1165_U85, R1165_U490, R1165_U491);
  nand ginst2891 (R1165_U86, R1165_U499, R1165_U500);
  nand ginst2892 (R1165_U87, R1165_U493, R1165_U494);
  nand ginst2893 (R1165_U88, R1165_U496, R1165_U497);
  nand ginst2894 (R1165_U89, R1165_U448, R1165_U449);
  and ginst2895 (R1165_U9, R1165_U297, R1165_U298);
  nand ginst2896 (R1165_U90, R1165_U505, R1165_U506);
  nand ginst2897 (R1165_U91, R1165_U612, R1165_U613);
  nand ginst2898 (R1165_U92, R1165_U411, R1165_U412);
  nand ginst2899 (R1165_U93, R1165_U418, R1165_U419);
  nand ginst2900 (R1165_U94, R1165_U425, R1165_U426);
  nand ginst2901 (R1165_U95, R1165_U432, R1165_U433);
  nand ginst2902 (R1165_U96, R1165_U439, R1165_U440);
  nand ginst2903 (R1165_U97, R1165_U446, R1165_U447);
  nand ginst2904 (R1165_U98, R1165_U508, R1165_U509);
  nand ginst2905 (R1165_U99, R1165_U515, R1165_U516);
  and ginst2906 (R1171_U10, R1171_U281, R1171_U282);
  nand ginst2907 (R1171_U100, R1171_U314, R1171_U60);
  nand ginst2908 (R1171_U101, R1171_U294, R1171_U385);
  nand ginst2909 (R1171_U102, R1171_U277, R1171_U278);
  not ginst2910 (R1171_U103, U3073);
  nand ginst2911 (R1171_U104, R1171_U323, R1171_U84);
  nand ginst2912 (R1171_U105, R1171_U271, R1171_U382, R1171_U383);
  nand ginst2913 (R1171_U106, R1171_U345, R1171_U72);
  nand ginst2914 (R1171_U107, R1171_U483, R1171_U484);
  nand ginst2915 (R1171_U108, R1171_U530, R1171_U531);
  nand ginst2916 (R1171_U109, R1171_U401, R1171_U402);
  and ginst2917 (R1171_U11, R1171_U10, R1171_U283);
  nand ginst2918 (R1171_U110, R1171_U406, R1171_U407);
  nand ginst2919 (R1171_U111, R1171_U413, R1171_U414);
  nand ginst2920 (R1171_U112, R1171_U420, R1171_U421);
  nand ginst2921 (R1171_U113, R1171_U425, R1171_U426);
  nand ginst2922 (R1171_U114, R1171_U434, R1171_U435);
  nand ginst2923 (R1171_U115, R1171_U441, R1171_U442);
  nand ginst2924 (R1171_U116, R1171_U448, R1171_U449);
  nand ginst2925 (R1171_U117, R1171_U455, R1171_U456);
  nand ginst2926 (R1171_U118, R1171_U460, R1171_U461);
  nand ginst2927 (R1171_U119, R1171_U467, R1171_U468);
  and ginst2928 (R1171_U12, R1171_U217, R1171_U7);
  nand ginst2929 (R1171_U120, R1171_U474, R1171_U475);
  nand ginst2930 (R1171_U121, R1171_U488, R1171_U489);
  nand ginst2931 (R1171_U122, R1171_U493, R1171_U494);
  nand ginst2932 (R1171_U123, R1171_U500, R1171_U501);
  nand ginst2933 (R1171_U124, R1171_U507, R1171_U508);
  nand ginst2934 (R1171_U125, R1171_U514, R1171_U515);
  nand ginst2935 (R1171_U126, R1171_U521, R1171_U522);
  nand ginst2936 (R1171_U127, R1171_U526, R1171_U527);
  and ginst2937 (R1171_U128, R1171_U129, R1171_U197);
  and ginst2938 (R1171_U129, U3065, U3470);
  and ginst2939 (R1171_U13, R1171_U262, R1171_U8);
  and ginst2940 (R1171_U130, U3061, U3472);
  and ginst2941 (R1171_U131, U3074, U3464);
  and ginst2942 (R1171_U132, R1171_U203, R1171_U204, R1171_U206);
  and ginst2943 (R1171_U133, R1171_U207, R1171_U373, R1171_U374);
  and ginst2944 (R1171_U134, R1171_U408, R1171_U409, R1171_U43);
  and ginst2945 (R1171_U135, R1171_U225, R1171_U6);
  and ginst2946 (R1171_U136, R1171_U231, R1171_U233);
  and ginst2947 (R1171_U137, R1171_U34, R1171_U415, R1171_U416);
  and ginst2948 (R1171_U138, R1171_U239, R1171_U4);
  and ginst2949 (R1171_U139, R1171_U198, R1171_U247);
  and ginst2950 (R1171_U14, R1171_U11, R1171_U292);
  and ginst2951 (R1171_U140, R1171_U188, R1171_U252);
  and ginst2952 (R1171_U141, R1171_U12, R1171_U6);
  and ginst2953 (R1171_U142, R1171_U255, R1171_U378);
  and ginst2954 (R1171_U143, R1171_U15, R1171_U270);
  and ginst2955 (R1171_U144, R1171_U189, R1171_U260);
  and ginst2956 (R1171_U145, R1171_U16, R1171_U296);
  and ginst2957 (R1171_U146, R1171_U297, R1171_U389);
  and ginst2958 (R1171_U147, R1171_U185, R1171_U309);
  and ginst2959 (R1171_U148, R1171_U310, R1171_U393, R1171_U395);
  and ginst2960 (R1171_U149, R1171_U17, R1171_U185);
  and ginst2961 (R1171_U15, R1171_U13, R1171_U267);
  and ginst2962 (R1171_U150, R1171_U304, R1171_U97);
  and ginst2963 (R1171_U151, R1171_U190, R1171_U450, R1171_U451);
  and ginst2964 (R1171_U152, R1171_U185, R1171_U320);
  and ginst2965 (R1171_U153, R1171_U176, R1171_U288);
  and ginst2966 (R1171_U154, R1171_U481, R1171_U482, R1171_U80);
  and ginst2967 (R1171_U155, R1171_U10, R1171_U333);
  and ginst2968 (R1171_U156, R1171_U495, R1171_U496, R1171_U90);
  and ginst2969 (R1171_U157, R1171_U342, R1171_U9);
  and ginst2970 (R1171_U158, R1171_U189, R1171_U516, R1171_U517);
  and ginst2971 (R1171_U159, R1171_U351, R1171_U8);
  and ginst2972 (R1171_U16, R1171_U14, R1171_U9);
  and ginst2973 (R1171_U160, R1171_U188, R1171_U528, R1171_U529);
  and ginst2974 (R1171_U161, R1171_U358, R1171_U7);
  nand ginst2975 (R1171_U162, R1171_U215, R1171_U375);
  nand ginst2976 (R1171_U163, R1171_U230, R1171_U242);
  not ginst2977 (R1171_U164, U3052);
  not ginst2978 (R1171_U165, U4040);
  and ginst2979 (R1171_U166, R1171_U429, R1171_U430);
  nand ginst2980 (R1171_U167, R1171_U186, R1171_U312, R1171_U372);
  and ginst2981 (R1171_U168, R1171_U436, R1171_U437);
  nand ginst2982 (R1171_U169, R1171_U148, R1171_U394);
  and ginst2983 (R1171_U17, R1171_U299, R1171_U305);
  and ginst2984 (R1171_U170, R1171_U443, R1171_U444);
  nand ginst2985 (R1171_U171, R1171_U150, R1171_U307);
  nand ginst2986 (R1171_U172, R1171_U300, R1171_U301);
  and ginst2987 (R1171_U173, R1171_U462, R1171_U463);
  and ginst2988 (R1171_U174, R1171_U469, R1171_U470);
  nand ginst2989 (R1171_U175, R1171_U384, R1171_U386);
  and ginst2990 (R1171_U176, R1171_U476, R1171_U477);
  nand ginst2991 (R1171_U177, U3074, U3464);
  nand ginst2992 (R1171_U178, R1171_U335, R1171_U36);
  nand ginst2993 (R1171_U179, R1171_U279, R1171_U376);
  and ginst2994 (R1171_U18, R1171_U356, R1171_U359);
  and ginst2995 (R1171_U180, R1171_U502, R1171_U503);
  nand ginst2996 (R1171_U181, R1171_U379, R1171_U77);
  and ginst2997 (R1171_U182, R1171_U509, R1171_U510);
  nand ginst2998 (R1171_U183, R1171_U264, R1171_U265);
  nand ginst2999 (R1171_U184, R1171_U142, R1171_U377);
  nand ginst3000 (R1171_U185, R1171_U390, R1171_U391);
  nand ginst3001 (R1171_U186, R1171_U169, U3051);
  not ginst3002 (R1171_U187, R1171_U34);
  nand ginst3003 (R1171_U188, U3080, U3484);
  nand ginst3004 (R1171_U189, U3069, U3490);
  and ginst3005 (R1171_U19, R1171_U349, R1171_U352);
  nand ginst3006 (R1171_U190, U3055, U4032);
  not ginst3007 (R1171_U191, R1171_U72);
  not ginst3008 (R1171_U192, R1171_U84);
  not ginst3009 (R1171_U193, R1171_U60);
  not ginst3010 (R1171_U194, R1171_U65);
  or ginst3011 (R1171_U195, U3064, U3476);
  or ginst3012 (R1171_U196, U3057, U3474);
  or ginst3013 (R1171_U197, U3061, U3472);
  or ginst3014 (R1171_U198, U3065, U3470);
  not ginst3015 (R1171_U199, R1171_U177);
  and ginst3016 (R1171_U20, R1171_U340, R1171_U343);
  or ginst3017 (R1171_U200, U3075, U3468);
  not ginst3018 (R1171_U201, R1171_U39);
  not ginst3019 (R1171_U202, R1171_U36);
  nand ginst3020 (R1171_U203, R1171_U128, R1171_U4);
  nand ginst3021 (R1171_U204, R1171_U130, R1171_U4);
  nand ginst3022 (R1171_U205, R1171_U34, R1171_U35);
  nand ginst3023 (R1171_U206, R1171_U205, U3064);
  nand ginst3024 (R1171_U207, R1171_U187, U3476);
  not ginst3025 (R1171_U208, R1171_U51);
  or ginst3026 (R1171_U209, U3067, U3480);
  and ginst3027 (R1171_U21, R1171_U331, R1171_U334);
  or ginst3028 (R1171_U210, U3068, U3478);
  not ginst3029 (R1171_U211, R1171_U43);
  nand ginst3030 (R1171_U212, R1171_U43, R1171_U44);
  nand ginst3031 (R1171_U213, R1171_U212, U3067);
  nand ginst3032 (R1171_U214, R1171_U211, U3480);
  nand ginst3033 (R1171_U215, R1171_U51, R1171_U6);
  not ginst3034 (R1171_U216, R1171_U162);
  or ginst3035 (R1171_U217, U3081, U3482);
  nand ginst3036 (R1171_U218, R1171_U162, R1171_U217);
  not ginst3037 (R1171_U219, R1171_U50);
  and ginst3038 (R1171_U22, R1171_U326, R1171_U328);
  or ginst3039 (R1171_U220, U3080, U3484);
  or ginst3040 (R1171_U221, U3068, U3478);
  nand ginst3041 (R1171_U222, R1171_U221, R1171_U51);
  nand ginst3042 (R1171_U223, R1171_U134, R1171_U222);
  nand ginst3043 (R1171_U224, R1171_U208, R1171_U43);
  nand ginst3044 (R1171_U225, U3067, U3480);
  nand ginst3045 (R1171_U226, R1171_U135, R1171_U224);
  or ginst3046 (R1171_U227, U3068, U3478);
  nand ginst3047 (R1171_U228, R1171_U198, R1171_U202);
  nand ginst3048 (R1171_U229, U3065, U3470);
  and ginst3049 (R1171_U23, R1171_U318, R1171_U321);
  not ginst3050 (R1171_U230, R1171_U53);
  nand ginst3051 (R1171_U231, R1171_U201, R1171_U5);
  nand ginst3052 (R1171_U232, R1171_U197, R1171_U53);
  nand ginst3053 (R1171_U233, U3061, U3472);
  not ginst3054 (R1171_U234, R1171_U52);
  or ginst3055 (R1171_U235, U3057, U3474);
  nand ginst3056 (R1171_U236, R1171_U235, R1171_U52);
  nand ginst3057 (R1171_U237, R1171_U137, R1171_U236);
  nand ginst3058 (R1171_U238, R1171_U234, R1171_U34);
  nand ginst3059 (R1171_U239, U3064, U3476);
  and ginst3060 (R1171_U24, R1171_U245, R1171_U248);
  nand ginst3061 (R1171_U240, R1171_U138, R1171_U238);
  or ginst3062 (R1171_U241, U3057, U3474);
  nand ginst3063 (R1171_U242, R1171_U198, R1171_U201);
  not ginst3064 (R1171_U243, R1171_U163);
  nand ginst3065 (R1171_U244, U3061, U3472);
  nand ginst3066 (R1171_U245, R1171_U36, R1171_U39, R1171_U427, R1171_U428);
  nand ginst3067 (R1171_U246, R1171_U36, R1171_U39);
  nand ginst3068 (R1171_U247, U3065, U3470);
  nand ginst3069 (R1171_U248, R1171_U139, R1171_U246);
  or ginst3070 (R1171_U249, U3080, U3484);
  and ginst3071 (R1171_U25, R1171_U237, R1171_U240);
  or ginst3072 (R1171_U250, U3059, U3486);
  nand ginst3073 (R1171_U251, R1171_U194, R1171_U7);
  nand ginst3074 (R1171_U252, U3059, U3486);
  nand ginst3075 (R1171_U253, R1171_U140, R1171_U251);
  or ginst3076 (R1171_U254, U3059, U3486);
  nand ginst3077 (R1171_U255, R1171_U253, R1171_U254);
  not ginst3078 (R1171_U256, R1171_U184);
  or ginst3079 (R1171_U257, U3077, U3492);
  or ginst3080 (R1171_U258, U3069, U3490);
  nand ginst3081 (R1171_U259, R1171_U191, R1171_U8);
  and ginst3082 (R1171_U26, R1171_U223, R1171_U226);
  nand ginst3083 (R1171_U260, U3077, U3492);
  nand ginst3084 (R1171_U261, R1171_U144, R1171_U259);
  or ginst3085 (R1171_U262, U3060, U3488);
  or ginst3086 (R1171_U263, U3077, U3492);
  nand ginst3087 (R1171_U264, R1171_U13, R1171_U184);
  nand ginst3088 (R1171_U265, R1171_U261, R1171_U263);
  not ginst3089 (R1171_U266, R1171_U183);
  or ginst3090 (R1171_U267, U3076, U3494);
  nand ginst3091 (R1171_U268, U3076, U3494);
  not ginst3092 (R1171_U269, R1171_U181);
  not ginst3093 (R1171_U27, U3470);
  or ginst3094 (R1171_U270, U3071, U3496);
  nand ginst3095 (R1171_U271, U3071, U3496);
  not ginst3096 (R1171_U272, R1171_U105);
  or ginst3097 (R1171_U273, U3066, U3500);
  or ginst3098 (R1171_U274, U3070, U3498);
  not ginst3099 (R1171_U275, R1171_U90);
  nand ginst3100 (R1171_U276, R1171_U90, R1171_U91);
  nand ginst3101 (R1171_U277, R1171_U276, U3066);
  nand ginst3102 (R1171_U278, R1171_U275, U3500);
  nand ginst3103 (R1171_U279, R1171_U105, R1171_U9);
  not ginst3104 (R1171_U28, U3065);
  not ginst3105 (R1171_U280, R1171_U179);
  or ginst3106 (R1171_U281, U3073, U4037);
  or ginst3107 (R1171_U282, U3078, U3504);
  or ginst3108 (R1171_U283, U3072, U4036);
  not ginst3109 (R1171_U284, R1171_U80);
  nand ginst3110 (R1171_U285, R1171_U284, U4037);
  nand ginst3111 (R1171_U286, R1171_U103, R1171_U285);
  nand ginst3112 (R1171_U287, R1171_U80, R1171_U81);
  nand ginst3113 (R1171_U288, R1171_U286, R1171_U287);
  nand ginst3114 (R1171_U289, R1171_U11, R1171_U192);
  not ginst3115 (R1171_U29, U3472);
  nand ginst3116 (R1171_U290, U3072, U4036);
  nand ginst3117 (R1171_U291, R1171_U288, R1171_U289, R1171_U290);
  or ginst3118 (R1171_U292, U3079, U3502);
  or ginst3119 (R1171_U293, U3072, U4036);
  nand ginst3120 (R1171_U294, R1171_U291, R1171_U293);
  not ginst3121 (R1171_U295, R1171_U175);
  or ginst3122 (R1171_U296, U3058, U4035);
  nand ginst3123 (R1171_U297, U3058, U4035);
  not ginst3124 (R1171_U298, R1171_U94);
  or ginst3125 (R1171_U299, U3063, U4034);
  not ginst3126 (R1171_U30, U3061);
  nand ginst3127 (R1171_U300, R1171_U299, R1171_U94);
  nand ginst3128 (R1171_U301, U3063, U4034);
  not ginst3129 (R1171_U302, R1171_U172);
  or ginst3130 (R1171_U303, U3055, U4032);
  nand ginst3131 (R1171_U304, R1171_U185, R1171_U193);
  or ginst3132 (R1171_U305, U3062, U4033);
  or ginst3133 (R1171_U306, U3054, U4031);
  nand ginst3134 (R1171_U307, R1171_U149, R1171_U392);
  not ginst3135 (R1171_U308, R1171_U171);
  or ginst3136 (R1171_U309, U3050, U4030);
  not ginst3137 (R1171_U31, U3474);
  nand ginst3138 (R1171_U310, U3050, U4030);
  not ginst3139 (R1171_U311, R1171_U169);
  nand ginst3140 (R1171_U312, R1171_U169, U4029);
  not ginst3141 (R1171_U313, R1171_U167);
  nand ginst3142 (R1171_U314, R1171_U172, R1171_U305);
  not ginst3143 (R1171_U315, R1171_U100);
  or ginst3144 (R1171_U316, U3055, U4032);
  nand ginst3145 (R1171_U317, R1171_U100, R1171_U316);
  nand ginst3146 (R1171_U318, R1171_U151, R1171_U317);
  nand ginst3147 (R1171_U319, R1171_U190, R1171_U315);
  not ginst3148 (R1171_U32, U3057);
  nand ginst3149 (R1171_U320, U3054, U4031);
  nand ginst3150 (R1171_U321, R1171_U152, R1171_U319);
  or ginst3151 (R1171_U322, U3055, U4032);
  nand ginst3152 (R1171_U323, R1171_U179, R1171_U292);
  not ginst3153 (R1171_U324, R1171_U104);
  nand ginst3154 (R1171_U325, R1171_U10, R1171_U104);
  nand ginst3155 (R1171_U326, R1171_U153, R1171_U325);
  nand ginst3156 (R1171_U327, R1171_U288, R1171_U325);
  nand ginst3157 (R1171_U328, R1171_U327, R1171_U480);
  or ginst3158 (R1171_U329, U3078, U3504);
  not ginst3159 (R1171_U33, U3064);
  nand ginst3160 (R1171_U330, R1171_U104, R1171_U329);
  nand ginst3161 (R1171_U331, R1171_U154, R1171_U330);
  nand ginst3162 (R1171_U332, R1171_U324, R1171_U80);
  nand ginst3163 (R1171_U333, U3073, U4037);
  nand ginst3164 (R1171_U334, R1171_U155, R1171_U332);
  or ginst3165 (R1171_U335, U3075, U3468);
  not ginst3166 (R1171_U336, R1171_U178);
  or ginst3167 (R1171_U337, U3078, U3504);
  or ginst3168 (R1171_U338, U3070, U3498);
  nand ginst3169 (R1171_U339, R1171_U105, R1171_U338);
  nand ginst3170 (R1171_U34, U3057, U3474);
  nand ginst3171 (R1171_U340, R1171_U156, R1171_U339);
  nand ginst3172 (R1171_U341, R1171_U272, R1171_U90);
  nand ginst3173 (R1171_U342, U3066, U3500);
  nand ginst3174 (R1171_U343, R1171_U157, R1171_U341);
  or ginst3175 (R1171_U344, U3070, U3498);
  nand ginst3176 (R1171_U345, R1171_U184, R1171_U262);
  not ginst3177 (R1171_U346, R1171_U106);
  or ginst3178 (R1171_U347, U3069, U3490);
  nand ginst3179 (R1171_U348, R1171_U106, R1171_U347);
  nand ginst3180 (R1171_U349, R1171_U158, R1171_U348);
  not ginst3181 (R1171_U35, U3476);
  nand ginst3182 (R1171_U350, R1171_U189, R1171_U346);
  nand ginst3183 (R1171_U351, U3077, U3492);
  nand ginst3184 (R1171_U352, R1171_U159, R1171_U350);
  or ginst3185 (R1171_U353, U3069, U3490);
  or ginst3186 (R1171_U354, U3080, U3484);
  nand ginst3187 (R1171_U355, R1171_U354, R1171_U50);
  nand ginst3188 (R1171_U356, R1171_U160, R1171_U355);
  nand ginst3189 (R1171_U357, R1171_U188, R1171_U219);
  nand ginst3190 (R1171_U358, U3059, U3486);
  nand ginst3191 (R1171_U359, R1171_U161, R1171_U357);
  nand ginst3192 (R1171_U36, U3075, U3468);
  nand ginst3193 (R1171_U360, R1171_U188, R1171_U220);
  nand ginst3194 (R1171_U361, R1171_U217, R1171_U65);
  nand ginst3195 (R1171_U362, R1171_U227, R1171_U43);
  nand ginst3196 (R1171_U363, R1171_U241, R1171_U34);
  nand ginst3197 (R1171_U364, R1171_U197, R1171_U244);
  nand ginst3198 (R1171_U365, R1171_U190, R1171_U322);
  nand ginst3199 (R1171_U366, R1171_U305, R1171_U60);
  nand ginst3200 (R1171_U367, R1171_U337, R1171_U80);
  nand ginst3201 (R1171_U368, R1171_U292, R1171_U84);
  nand ginst3202 (R1171_U369, R1171_U344, R1171_U90);
  not ginst3203 (R1171_U37, U3464);
  nand ginst3204 (R1171_U370, R1171_U189, R1171_U353);
  nand ginst3205 (R1171_U371, R1171_U262, R1171_U72);
  nand ginst3206 (R1171_U372, U3051, U4029);
  nand ginst3207 (R1171_U373, R1171_U202, R1171_U4, R1171_U5);
  nand ginst3208 (R1171_U374, R1171_U201, R1171_U4, R1171_U5);
  not ginst3209 (R1171_U375, R1171_U45);
  not ginst3210 (R1171_U376, R1171_U102);
  nand ginst3211 (R1171_U377, R1171_U141, R1171_U51);
  nand ginst3212 (R1171_U378, R1171_U12, R1171_U45);
  nand ginst3213 (R1171_U379, R1171_U15, R1171_U184);
  not ginst3214 (R1171_U38, U3074);
  nand ginst3215 (R1171_U380, R1171_U265, R1171_U268);
  not ginst3216 (R1171_U381, R1171_U77);
  nand ginst3217 (R1171_U382, R1171_U143, R1171_U184);
  nand ginst3218 (R1171_U383, R1171_U270, R1171_U381);
  nand ginst3219 (R1171_U384, R1171_U105, R1171_U16);
  nand ginst3220 (R1171_U385, R1171_U102, R1171_U14);
  not ginst3221 (R1171_U386, R1171_U101);
  not ginst3222 (R1171_U387, R1171_U97);
  nand ginst3223 (R1171_U388, R1171_U105, R1171_U145);
  nand ginst3224 (R1171_U389, R1171_U101, R1171_U296);
  nand ginst3225 (R1171_U39, R1171_U131, R1171_U200);
  nand ginst3226 (R1171_U390, R1171_U303, U3054);
  nand ginst3227 (R1171_U391, R1171_U303, U4031);
  nand ginst3228 (R1171_U392, R1171_U298, R1171_U301);
  nand ginst3229 (R1171_U393, R1171_U185, R1171_U193, R1171_U309);
  nand ginst3230 (R1171_U394, R1171_U147, R1171_U17, R1171_U392);
  nand ginst3231 (R1171_U395, R1171_U309, R1171_U387);
  nand ginst3232 (R1171_U396, R1171_U190, R1171_U57);
  nand ginst3233 (R1171_U397, R1171_U190, R1171_U56);
  nand ginst3234 (R1171_U398, R1171_U49, U3080);
  nand ginst3235 (R1171_U399, R1171_U48, U3484);
  and ginst3236 (R1171_U4, R1171_U195, R1171_U196);
  not ginst3237 (R1171_U40, U3478);
  nand ginst3238 (R1171_U400, R1171_U398, R1171_U399);
  nand ginst3239 (R1171_U401, R1171_U360, R1171_U50);
  nand ginst3240 (R1171_U402, R1171_U219, R1171_U400);
  nand ginst3241 (R1171_U403, R1171_U46, U3081);
  nand ginst3242 (R1171_U404, R1171_U47, U3482);
  nand ginst3243 (R1171_U405, R1171_U403, R1171_U404);
  nand ginst3244 (R1171_U406, R1171_U162, R1171_U361);
  nand ginst3245 (R1171_U407, R1171_U216, R1171_U405);
  nand ginst3246 (R1171_U408, R1171_U44, U3067);
  nand ginst3247 (R1171_U409, R1171_U42, U3480);
  not ginst3248 (R1171_U41, U3068);
  nand ginst3249 (R1171_U410, R1171_U40, U3068);
  nand ginst3250 (R1171_U411, R1171_U41, U3478);
  nand ginst3251 (R1171_U412, R1171_U410, R1171_U411);
  nand ginst3252 (R1171_U413, R1171_U362, R1171_U51);
  nand ginst3253 (R1171_U414, R1171_U208, R1171_U412);
  nand ginst3254 (R1171_U415, R1171_U35, U3064);
  nand ginst3255 (R1171_U416, R1171_U33, U3476);
  nand ginst3256 (R1171_U417, R1171_U31, U3057);
  nand ginst3257 (R1171_U418, R1171_U32, U3474);
  nand ginst3258 (R1171_U419, R1171_U417, R1171_U418);
  not ginst3259 (R1171_U42, U3067);
  nand ginst3260 (R1171_U420, R1171_U363, R1171_U52);
  nand ginst3261 (R1171_U421, R1171_U234, R1171_U419);
  nand ginst3262 (R1171_U422, R1171_U29, U3061);
  nand ginst3263 (R1171_U423, R1171_U30, U3472);
  nand ginst3264 (R1171_U424, R1171_U422, R1171_U423);
  nand ginst3265 (R1171_U425, R1171_U163, R1171_U364);
  nand ginst3266 (R1171_U426, R1171_U243, R1171_U424);
  nand ginst3267 (R1171_U427, R1171_U27, U3065);
  nand ginst3268 (R1171_U428, R1171_U28, U3470);
  nand ginst3269 (R1171_U429, R1171_U165, U3052);
  nand ginst3270 (R1171_U43, U3068, U3478);
  nand ginst3271 (R1171_U430, R1171_U164, U4040);
  nand ginst3272 (R1171_U431, R1171_U165, U3052);
  nand ginst3273 (R1171_U432, R1171_U164, U4040);
  nand ginst3274 (R1171_U433, R1171_U431, R1171_U432);
  nand ginst3275 (R1171_U434, R1171_U166, R1171_U167);
  nand ginst3276 (R1171_U435, R1171_U313, R1171_U433);
  nand ginst3277 (R1171_U436, R1171_U99, U3051);
  nand ginst3278 (R1171_U437, R1171_U98, U4029);
  nand ginst3279 (R1171_U438, R1171_U99, U3051);
  nand ginst3280 (R1171_U439, R1171_U98, U4029);
  not ginst3281 (R1171_U44, U3480);
  nand ginst3282 (R1171_U440, R1171_U438, R1171_U439);
  nand ginst3283 (R1171_U441, R1171_U168, R1171_U169);
  nand ginst3284 (R1171_U442, R1171_U311, R1171_U440);
  nand ginst3285 (R1171_U443, R1171_U54, U3050);
  nand ginst3286 (R1171_U444, R1171_U55, U4030);
  nand ginst3287 (R1171_U445, R1171_U54, U3050);
  nand ginst3288 (R1171_U446, R1171_U55, U4030);
  nand ginst3289 (R1171_U447, R1171_U445, R1171_U446);
  nand ginst3290 (R1171_U448, R1171_U170, R1171_U171);
  nand ginst3291 (R1171_U449, R1171_U308, R1171_U447);
  nand ginst3292 (R1171_U45, R1171_U213, R1171_U214);
  nand ginst3293 (R1171_U450, R1171_U57, U3054);
  nand ginst3294 (R1171_U451, R1171_U56, U4031);
  nand ginst3295 (R1171_U452, R1171_U95, U3055);
  nand ginst3296 (R1171_U453, R1171_U96, U4032);
  nand ginst3297 (R1171_U454, R1171_U452, R1171_U453);
  nand ginst3298 (R1171_U455, R1171_U100, R1171_U365);
  nand ginst3299 (R1171_U456, R1171_U315, R1171_U454);
  nand ginst3300 (R1171_U457, R1171_U58, U3062);
  nand ginst3301 (R1171_U458, R1171_U59, U4033);
  nand ginst3302 (R1171_U459, R1171_U457, R1171_U458);
  not ginst3303 (R1171_U46, U3482);
  nand ginst3304 (R1171_U460, R1171_U172, R1171_U366);
  nand ginst3305 (R1171_U461, R1171_U302, R1171_U459);
  nand ginst3306 (R1171_U462, R1171_U92, U3063);
  nand ginst3307 (R1171_U463, R1171_U93, U4034);
  nand ginst3308 (R1171_U464, R1171_U92, U3063);
  nand ginst3309 (R1171_U465, R1171_U93, U4034);
  nand ginst3310 (R1171_U466, R1171_U464, R1171_U465);
  nand ginst3311 (R1171_U467, R1171_U173, R1171_U94);
  nand ginst3312 (R1171_U468, R1171_U298, R1171_U466);
  nand ginst3313 (R1171_U469, R1171_U61, U3058);
  not ginst3314 (R1171_U47, U3081);
  nand ginst3315 (R1171_U470, R1171_U62, U4035);
  nand ginst3316 (R1171_U471, R1171_U61, U3058);
  nand ginst3317 (R1171_U472, R1171_U62, U4035);
  nand ginst3318 (R1171_U473, R1171_U471, R1171_U472);
  nand ginst3319 (R1171_U474, R1171_U174, R1171_U175);
  nand ginst3320 (R1171_U475, R1171_U295, R1171_U473);
  nand ginst3321 (R1171_U476, R1171_U85, U3072);
  nand ginst3322 (R1171_U477, R1171_U86, U4036);
  nand ginst3323 (R1171_U478, R1171_U85, U3072);
  nand ginst3324 (R1171_U479, R1171_U86, U4036);
  not ginst3325 (R1171_U48, U3080);
  nand ginst3326 (R1171_U480, R1171_U478, R1171_U479);
  nand ginst3327 (R1171_U481, R1171_U81, U3073);
  nand ginst3328 (R1171_U482, R1171_U103, U4037);
  nand ginst3329 (R1171_U483, R1171_U178, R1171_U199);
  nand ginst3330 (R1171_U484, R1171_U177, R1171_U336);
  nand ginst3331 (R1171_U485, R1171_U78, U3078);
  nand ginst3332 (R1171_U486, R1171_U79, U3504);
  nand ginst3333 (R1171_U487, R1171_U485, R1171_U486);
  nand ginst3334 (R1171_U488, R1171_U104, R1171_U367);
  nand ginst3335 (R1171_U489, R1171_U324, R1171_U487);
  not ginst3336 (R1171_U49, U3484);
  nand ginst3337 (R1171_U490, R1171_U82, U3079);
  nand ginst3338 (R1171_U491, R1171_U83, U3502);
  nand ginst3339 (R1171_U492, R1171_U490, R1171_U491);
  nand ginst3340 (R1171_U493, R1171_U179, R1171_U368);
  nand ginst3341 (R1171_U494, R1171_U280, R1171_U492);
  nand ginst3342 (R1171_U495, R1171_U91, U3066);
  nand ginst3343 (R1171_U496, R1171_U89, U3500);
  nand ginst3344 (R1171_U497, R1171_U87, U3070);
  nand ginst3345 (R1171_U498, R1171_U88, U3498);
  nand ginst3346 (R1171_U499, R1171_U497, R1171_U498);
  and ginst3347 (R1171_U5, R1171_U197, R1171_U198);
  nand ginst3348 (R1171_U50, R1171_U218, R1171_U65);
  nand ginst3349 (R1171_U500, R1171_U105, R1171_U369);
  nand ginst3350 (R1171_U501, R1171_U272, R1171_U499);
  nand ginst3351 (R1171_U502, R1171_U63, U3071);
  nand ginst3352 (R1171_U503, R1171_U64, U3496);
  nand ginst3353 (R1171_U504, R1171_U63, U3071);
  nand ginst3354 (R1171_U505, R1171_U64, U3496);
  nand ginst3355 (R1171_U506, R1171_U504, R1171_U505);
  nand ginst3356 (R1171_U507, R1171_U180, R1171_U181);
  nand ginst3357 (R1171_U508, R1171_U269, R1171_U506);
  nand ginst3358 (R1171_U509, R1171_U75, U3076);
  nand ginst3359 (R1171_U51, R1171_U132, R1171_U133);
  nand ginst3360 (R1171_U510, R1171_U76, U3494);
  nand ginst3361 (R1171_U511, R1171_U75, U3076);
  nand ginst3362 (R1171_U512, R1171_U76, U3494);
  nand ginst3363 (R1171_U513, R1171_U511, R1171_U512);
  nand ginst3364 (R1171_U514, R1171_U182, R1171_U183);
  nand ginst3365 (R1171_U515, R1171_U266, R1171_U513);
  nand ginst3366 (R1171_U516, R1171_U73, U3077);
  nand ginst3367 (R1171_U517, R1171_U74, U3492);
  nand ginst3368 (R1171_U518, R1171_U68, U3069);
  nand ginst3369 (R1171_U519, R1171_U69, U3490);
  nand ginst3370 (R1171_U52, R1171_U136, R1171_U232);
  nand ginst3371 (R1171_U520, R1171_U518, R1171_U519);
  nand ginst3372 (R1171_U521, R1171_U106, R1171_U370);
  nand ginst3373 (R1171_U522, R1171_U346, R1171_U520);
  nand ginst3374 (R1171_U523, R1171_U70, U3060);
  nand ginst3375 (R1171_U524, R1171_U71, U3488);
  nand ginst3376 (R1171_U525, R1171_U523, R1171_U524);
  nand ginst3377 (R1171_U526, R1171_U184, R1171_U371);
  nand ginst3378 (R1171_U527, R1171_U256, R1171_U525);
  nand ginst3379 (R1171_U528, R1171_U66, U3059);
  nand ginst3380 (R1171_U529, R1171_U67, U3486);
  nand ginst3381 (R1171_U53, R1171_U228, R1171_U229);
  nand ginst3382 (R1171_U530, R1171_U37, U3074);
  nand ginst3383 (R1171_U531, R1171_U38, U3464);
  not ginst3384 (R1171_U54, U4030);
  not ginst3385 (R1171_U55, U3050);
  not ginst3386 (R1171_U56, U3054);
  not ginst3387 (R1171_U57, U4031);
  not ginst3388 (R1171_U58, U4033);
  not ginst3389 (R1171_U59, U3062);
  and ginst3390 (R1171_U6, R1171_U209, R1171_U210);
  nand ginst3391 (R1171_U60, U3062, U4033);
  not ginst3392 (R1171_U61, U4035);
  not ginst3393 (R1171_U62, U3058);
  not ginst3394 (R1171_U63, U3496);
  not ginst3395 (R1171_U64, U3071);
  nand ginst3396 (R1171_U65, U3081, U3482);
  not ginst3397 (R1171_U66, U3486);
  not ginst3398 (R1171_U67, U3059);
  not ginst3399 (R1171_U68, U3490);
  not ginst3400 (R1171_U69, U3069);
  and ginst3401 (R1171_U7, R1171_U249, R1171_U250);
  not ginst3402 (R1171_U70, U3488);
  not ginst3403 (R1171_U71, U3060);
  nand ginst3404 (R1171_U72, U3060, U3488);
  not ginst3405 (R1171_U73, U3492);
  not ginst3406 (R1171_U74, U3077);
  not ginst3407 (R1171_U75, U3494);
  not ginst3408 (R1171_U76, U3076);
  nand ginst3409 (R1171_U77, R1171_U267, R1171_U380);
  not ginst3410 (R1171_U78, U3504);
  not ginst3411 (R1171_U79, U3078);
  and ginst3412 (R1171_U8, R1171_U257, R1171_U258);
  nand ginst3413 (R1171_U80, U3078, U3504);
  not ginst3414 (R1171_U81, U4037);
  not ginst3415 (R1171_U82, U3502);
  not ginst3416 (R1171_U83, U3079);
  nand ginst3417 (R1171_U84, U3079, U3502);
  not ginst3418 (R1171_U85, U4036);
  not ginst3419 (R1171_U86, U3072);
  not ginst3420 (R1171_U87, U3498);
  not ginst3421 (R1171_U88, U3070);
  not ginst3422 (R1171_U89, U3066);
  and ginst3423 (R1171_U9, R1171_U273, R1171_U274);
  nand ginst3424 (R1171_U90, U3070, U3498);
  not ginst3425 (R1171_U91, U3500);
  not ginst3426 (R1171_U92, U4034);
  not ginst3427 (R1171_U93, U3063);
  nand ginst3428 (R1171_U94, R1171_U146, R1171_U388);
  not ginst3429 (R1171_U95, U4032);
  not ginst3430 (R1171_U96, U3055);
  nand ginst3431 (R1171_U97, R1171_U306, R1171_U396, R1171_U397);
  not ginst3432 (R1171_U98, U3051);
  not ginst3433 (R1171_U99, U4029);
  and ginst3434 (R1192_U10, R1192_U276, R1192_U277);
  not ginst3435 (R1192_U100, U3050);
  not ginst3436 (R1192_U101, U4029);
  not ginst3437 (R1192_U102, U3051);
  nand ginst3438 (R1192_U103, R1192_U302, R1192_U356);
  nand ginst3439 (R1192_U104, R1192_U300, R1192_U354);
  nand ginst3440 (R1192_U105, R1192_U292, R1192_U352);
  nand ginst3441 (R1192_U106, R1192_U65, U4035);
  nand ginst3442 (R1192_U107, R1192_U321, R1192_U95);
  nand ginst3443 (R1192_U108, R1192_U372, R1192_U89);
  not ginst3444 (R1192_U109, U3074);
  and ginst3445 (R1192_U11, R1192_U106, R1192_U293);
  nand ginst3446 (R1192_U110, R1192_U432, R1192_U433);
  nand ginst3447 (R1192_U111, R1192_U448, R1192_U449);
  nand ginst3448 (R1192_U112, R1192_U453, R1192_U454);
  nand ginst3449 (R1192_U113, R1192_U471, R1192_U472);
  nand ginst3450 (R1192_U114, R1192_U476, R1192_U477);
  nand ginst3451 (R1192_U115, R1192_U481, R1192_U482);
  nand ginst3452 (R1192_U116, R1192_U486, R1192_U487);
  nand ginst3453 (R1192_U117, R1192_U491, R1192_U492);
  nand ginst3454 (R1192_U118, R1192_U507, R1192_U508);
  nand ginst3455 (R1192_U119, R1192_U512, R1192_U513);
  and ginst3456 (R1192_U12, R1192_U294, R1192_U295);
  nand ginst3457 (R1192_U120, R1192_U391, R1192_U392);
  nand ginst3458 (R1192_U121, R1192_U400, R1192_U401);
  nand ginst3459 (R1192_U122, R1192_U407, R1192_U408);
  nand ginst3460 (R1192_U123, R1192_U411, R1192_U412);
  nand ginst3461 (R1192_U124, R1192_U420, R1192_U421);
  nand ginst3462 (R1192_U125, R1192_U443, R1192_U444);
  nand ginst3463 (R1192_U126, R1192_U462, R1192_U463);
  nand ginst3464 (R1192_U127, R1192_U466, R1192_U467);
  nand ginst3465 (R1192_U128, R1192_U498, R1192_U499);
  nand ginst3466 (R1192_U129, R1192_U502, R1192_U503);
  and ginst3467 (R1192_U13, R1192_U216, R1192_U229, R1192_U234);
  nand ginst3468 (R1192_U130, R1192_U519, R1192_U520);
  and ginst3469 (R1192_U131, R1192_U215, R1192_U225);
  and ginst3470 (R1192_U132, R1192_U227, R1192_U228);
  and ginst3471 (R1192_U133, R1192_U13, R1192_U14);
  and ginst3472 (R1192_U134, R1192_U241, R1192_U242);
  and ginst3473 (R1192_U135, R1192_U134, R1192_U346);
  and ginst3474 (R1192_U136, R1192_U34, R1192_U393, R1192_U394);
  and ginst3475 (R1192_U137, R1192_U217, R1192_U397);
  and ginst3476 (R1192_U138, R1192_U257, R1192_U6);
  and ginst3477 (R1192_U139, R1192_U216, R1192_U404);
  and ginst3478 (R1192_U14, R1192_U217, R1192_U239);
  and ginst3479 (R1192_U140, R1192_U413, R1192_U414, R1192_U42);
  and ginst3480 (R1192_U141, R1192_U215, R1192_U417);
  and ginst3481 (R1192_U142, R1192_U18, R1192_U273);
  and ginst3482 (R1192_U143, R1192_U16, R1192_U285);
  and ginst3483 (R1192_U144, R1192_U286, R1192_U351);
  and ginst3484 (R1192_U145, R1192_U21, R1192_U303);
  and ginst3485 (R1192_U146, R1192_U304, R1192_U358);
  and ginst3486 (R1192_U147, R1192_U214, R1192_U305);
  and ginst3487 (R1192_U148, R1192_U308, R1192_U309);
  and ginst3488 (R1192_U149, R1192_U311, R1192_U426);
  and ginst3489 (R1192_U15, R1192_U244, R1192_U7);
  and ginst3490 (R1192_U150, R1192_U308, R1192_U309);
  and ginst3491 (R1192_U151, R1192_U23, R1192_U312);
  nand ginst3492 (R1192_U152, R1192_U429, R1192_U430);
  and ginst3493 (R1192_U153, R1192_U214, R1192_U436);
  and ginst3494 (R1192_U154, R1192_U186, R1192_U214);
  nand ginst3495 (R1192_U155, R1192_U445, R1192_U446);
  nand ginst3496 (R1192_U156, R1192_U450, R1192_U451);
  and ginst3497 (R1192_U157, R1192_U22, R1192_U298);
  and ginst3498 (R1192_U158, R1192_U213, R1192_U317);
  and ginst3499 (R1192_U159, R1192_U68, U3058);
  and ginst3500 (R1192_U16, R1192_U280, R1192_U9);
  and ginst3501 (R1192_U160, R1192_U19, R1192_U298);
  and ginst3502 (R1192_U161, R1192_U12, R1192_U317, R1192_U360);
  nand ginst3503 (R1192_U162, R1192_U468, R1192_U469);
  nand ginst3504 (R1192_U163, R1192_U473, R1192_U474);
  nand ginst3505 (R1192_U164, R1192_U478, R1192_U479);
  nand ginst3506 (R1192_U165, R1192_U483, R1192_U484);
  nand ginst3507 (R1192_U166, R1192_U488, R1192_U489);
  and ginst3508 (R1192_U167, R1192_U10, R1192_U327);
  and ginst3509 (R1192_U168, R1192_U212, R1192_U495);
  nand ginst3510 (R1192_U169, R1192_U504, R1192_U505);
  and ginst3511 (R1192_U17, R1192_U11, R1192_U298);
  nand ginst3512 (R1192_U170, R1192_U509, R1192_U510);
  and ginst3513 (R1192_U171, R1192_U336, R1192_U8);
  and ginst3514 (R1192_U172, R1192_U211, R1192_U516);
  and ginst3515 (R1192_U173, R1192_U389, R1192_U390);
  nand ginst3516 (R1192_U174, R1192_U135, R1192_U345);
  and ginst3517 (R1192_U175, R1192_U398, R1192_U399);
  and ginst3518 (R1192_U176, R1192_U405, R1192_U406);
  and ginst3519 (R1192_U177, R1192_U409, R1192_U410);
  nand ginst3520 (R1192_U178, R1192_U132, R1192_U380);
  and ginst3521 (R1192_U179, R1192_U418, R1192_U419);
  and ginst3522 (R1192_U18, R1192_U15, R1192_U271);
  not ginst3523 (R1192_U180, U4040);
  not ginst3524 (R1192_U181, U3052);
  and ginst3525 (R1192_U182, R1192_U427, R1192_U428);
  nand ginst3526 (R1192_U183, R1192_U148, R1192_U306);
  and ginst3527 (R1192_U184, R1192_U439, R1192_U440);
  and ginst3528 (R1192_U185, R1192_U441, R1192_U442);
  nand ginst3529 (R1192_U186, R1192_U146, R1192_U370);
  nand ginst3530 (R1192_U187, R1192_U357, R1192_U367);
  nand ginst3531 (R1192_U188, R1192_U355, R1192_U365);
  and ginst3532 (R1192_U189, R1192_U460, R1192_U461);
  and ginst3533 (R1192_U19, R1192_U289, R1192_U291);
  nand ginst3534 (R1192_U190, R1192_U315, R1192_U69);
  and ginst3535 (R1192_U191, R1192_U464, R1192_U465);
  nand ginst3536 (R1192_U192, R1192_U353, R1192_U363);
  nand ginst3537 (R1192_U193, R1192_U361, R1192_U74);
  not ginst3538 (R1192_U194, U3468);
  nand ginst3539 (R1192_U195, R1192_U109, U3464);
  nand ginst3540 (R1192_U196, R1192_U342, R1192_U385);
  nand ginst3541 (R1192_U197, R1192_U144, R1192_U350);
  nand ginst3542 (R1192_U198, R1192_U282, R1192_U96);
  and ginst3543 (R1192_U199, R1192_U496, R1192_U497);
  and ginst3544 (R1192_U20, R1192_U17, R1192_U19);
  and ginst3545 (R1192_U200, R1192_U500, R1192_U501);
  nand ginst3546 (R1192_U201, R1192_U274, R1192_U349, R1192_U378);
  nand ginst3547 (R1192_U202, R1192_U376, R1192_U91);
  nand ginst3548 (R1192_U203, R1192_U270, R1192_U374);
  and ginst3549 (R1192_U204, R1192_U517, R1192_U518);
  nand ginst3550 (R1192_U205, R1192_U153, R1192_U186);
  nand ginst3551 (R1192_U206, R1192_U149, R1192_U183);
  nand ginst3552 (R1192_U207, R1192_U194, R1192_U195);
  not ginst3553 (R1192_U208, R1192_U99);
  not ginst3554 (R1192_U209, R1192_U42);
  and ginst3555 (R1192_U21, R1192_U20, R1192_U301);
  not ginst3556 (R1192_U210, R1192_U34);
  nand ginst3557 (R1192_U211, R1192_U86, U3486);
  nand ginst3558 (R1192_U212, R1192_U93, U3496);
  not ginst3559 (R1192_U213, R1192_U106);
  nand ginst3560 (R1192_U214, R1192_U98, U4031);
  nand ginst3561 (R1192_U215, R1192_U41, U3470);
  nand ginst3562 (R1192_U216, R1192_U49, U3476);
  nand ginst3563 (R1192_U217, R1192_U33, U3480);
  not ginst3564 (R1192_U218, R1192_U95);
  not ginst3565 (R1192_U219, R1192_U69);
  and ginst3566 (R1192_U22, R1192_U106, R1192_U457);
  not ginst3567 (R1192_U220, R1192_U51);
  not ginst3568 (R1192_U221, R1192_U89);
  not ginst3569 (R1192_U222, R1192_U195);
  nand ginst3570 (R1192_U223, R1192_U195, U3075);
  not ginst3571 (R1192_U224, R1192_U57);
  nand ginst3572 (R1192_U225, R1192_U43, U3472);
  nand ginst3573 (R1192_U226, R1192_U42, R1192_U43);
  nand ginst3574 (R1192_U227, R1192_U226, R1192_U47);
  nand ginst3575 (R1192_U228, R1192_U209, U3061);
  nand ginst3576 (R1192_U229, R1192_U48, U3478);
  and ginst3577 (R1192_U23, R1192_U422, R1192_U423);
  nand ginst3578 (R1192_U230, R1192_U37, U3068);
  nand ginst3579 (R1192_U231, R1192_U36, U3064);
  nand ginst3580 (R1192_U232, R1192_U216, R1192_U220);
  nand ginst3581 (R1192_U233, R1192_U232, R1192_U6);
  nand ginst3582 (R1192_U234, R1192_U50, U3474);
  nand ginst3583 (R1192_U235, R1192_U48, U3478);
  nand ginst3584 (R1192_U236, R1192_U13, R1192_U178);
  not ginst3585 (R1192_U237, R1192_U52);
  not ginst3586 (R1192_U238, R1192_U55);
  nand ginst3587 (R1192_U239, R1192_U35, U3482);
  nand ginst3588 (R1192_U24, R1192_U334, R1192_U337);
  nand ginst3589 (R1192_U240, R1192_U34, R1192_U35);
  nand ginst3590 (R1192_U241, R1192_U240, R1192_U40);
  nand ginst3591 (R1192_U242, R1192_U210, U3081);
  not ginst3592 (R1192_U243, R1192_U174);
  nand ginst3593 (R1192_U244, R1192_U54, U3484);
  nand ginst3594 (R1192_U245, R1192_U244, R1192_U89);
  nand ginst3595 (R1192_U246, R1192_U238, R1192_U34);
  nand ginst3596 (R1192_U247, R1192_U137, R1192_U246);
  nand ginst3597 (R1192_U248, R1192_U217, R1192_U55);
  nand ginst3598 (R1192_U249, R1192_U136, R1192_U248);
  nand ginst3599 (R1192_U25, R1192_U325, R1192_U328);
  nand ginst3600 (R1192_U250, R1192_U217, R1192_U34);
  nand ginst3601 (R1192_U251, R1192_U178, R1192_U234);
  not ginst3602 (R1192_U252, R1192_U56);
  nand ginst3603 (R1192_U253, R1192_U36, U3064);
  nand ginst3604 (R1192_U254, R1192_U252, R1192_U253);
  nand ginst3605 (R1192_U255, R1192_U139, R1192_U254);
  nand ginst3606 (R1192_U256, R1192_U216, R1192_U56);
  nand ginst3607 (R1192_U257, R1192_U48, U3478);
  nand ginst3608 (R1192_U258, R1192_U138, R1192_U256);
  nand ginst3609 (R1192_U259, R1192_U36, U3064);
  nand ginst3610 (R1192_U26, R1192_U359, R1192_U387, R1192_U388, R1192_U458, R1192_U459);
  nand ginst3611 (R1192_U260, R1192_U216, R1192_U259);
  nand ginst3612 (R1192_U261, R1192_U234, R1192_U51);
  nand ginst3613 (R1192_U262, R1192_U141, R1192_U384);
  nand ginst3614 (R1192_U263, R1192_U215, R1192_U42);
  nand ginst3615 (R1192_U264, R1192_U85, U3488);
  nand ginst3616 (R1192_U265, R1192_U87, U3060);
  nand ginst3617 (R1192_U266, R1192_U88, U3059);
  nand ginst3618 (R1192_U267, R1192_U221, R1192_U7);
  nand ginst3619 (R1192_U268, R1192_U267, R1192_U8);
  nand ginst3620 (R1192_U269, R1192_U85, U3488);
  and ginst3621 (R1192_U27, R1192_U313, R1192_U344);
  nand ginst3622 (R1192_U270, R1192_U268, R1192_U269);
  nand ginst3623 (R1192_U271, R1192_U90, U3490);
  nand ginst3624 (R1192_U272, R1192_U84, U3069);
  nand ginst3625 (R1192_U273, R1192_U82, U3492);
  nand ginst3626 (R1192_U274, R1192_U83, U3077);
  nand ginst3627 (R1192_U275, R1192_U92, U3498);
  nand ginst3628 (R1192_U276, R1192_U79, U3070);
  nand ginst3629 (R1192_U277, R1192_U80, U3071);
  nand ginst3630 (R1192_U278, R1192_U218, R1192_U9);
  nand ginst3631 (R1192_U279, R1192_U10, R1192_U278);
  nand ginst3632 (R1192_U28, R1192_U182, R1192_U206, R1192_U343);
  nand ginst3633 (R1192_U280, R1192_U94, U3494);
  nand ginst3634 (R1192_U281, R1192_U92, U3498);
  nand ginst3635 (R1192_U282, R1192_U16, R1192_U201);
  not ginst3636 (R1192_U283, R1192_U96);
  not ginst3637 (R1192_U284, R1192_U198);
  nand ginst3638 (R1192_U285, R1192_U77, U3500);
  nand ginst3639 (R1192_U286, R1192_U78, U3066);
  not ginst3640 (R1192_U287, R1192_U197);
  nand ginst3641 (R1192_U288, R1192_U76, U3502);
  nand ginst3642 (R1192_U289, R1192_U72, U3504);
  nand ginst3643 (R1192_U29, R1192_U262, R1192_U383);
  not ginst3644 (R1192_U290, R1192_U74);
  nand ginst3645 (R1192_U291, R1192_U71, U4037);
  nand ginst3646 (R1192_U292, R1192_U73, U3073);
  nand ginst3647 (R1192_U293, R1192_U64, U4034);
  nand ginst3648 (R1192_U294, R1192_U67, U3063);
  nand ginst3649 (R1192_U295, R1192_U68, U3058);
  nand ginst3650 (R1192_U296, R1192_U11, R1192_U219);
  nand ginst3651 (R1192_U297, R1192_U12, R1192_U296);
  nand ginst3652 (R1192_U298, R1192_U66, U4036);
  nand ginst3653 (R1192_U299, R1192_U64, U4034);
  nand ginst3654 (R1192_U30, R1192_U255, R1192_U258);
  nand ginst3655 (R1192_U300, R1192_U297, R1192_U299);
  nand ginst3656 (R1192_U301, R1192_U62, U4033);
  nand ginst3657 (R1192_U302, R1192_U63, U3062);
  nand ginst3658 (R1192_U303, R1192_U60, U4032);
  nand ginst3659 (R1192_U304, R1192_U61, U3055);
  nand ginst3660 (R1192_U305, R1192_U100, U4030);
  nand ginst3661 (R1192_U306, R1192_U147, R1192_U186);
  nand ginst3662 (R1192_U307, R1192_U100, R1192_U99);
  nand ginst3663 (R1192_U308, R1192_U307, R1192_U59);
  nand ginst3664 (R1192_U309, R1192_U208, U3050);
  nand ginst3665 (R1192_U31, R1192_U247, R1192_U249);
  not ginst3666 (R1192_U310, R1192_U183);
  nand ginst3667 (R1192_U311, R1192_U102, U4029);
  nand ginst3668 (R1192_U312, R1192_U101, U3051);
  nand ginst3669 (R1192_U313, R1192_U154, R1192_U205);
  nand ginst3670 (R1192_U314, R1192_U214, R1192_U99);
  nand ginst3671 (R1192_U315, R1192_U192, R1192_U298);
  not ginst3672 (R1192_U316, R1192_U190);
  nand ginst3673 (R1192_U317, R1192_U64, U4034);
  nand ginst3674 (R1192_U318, R1192_U68, U3058);
  nand ginst3675 (R1192_U319, R1192_U106, R1192_U318);
  nand ginst3676 (R1192_U32, R1192_U195, R1192_U340);
  nand ginst3677 (R1192_U320, R1192_U298, R1192_U69);
  nand ginst3678 (R1192_U321, R1192_U201, R1192_U280);
  not ginst3679 (R1192_U322, R1192_U107);
  nand ginst3680 (R1192_U323, R1192_U80, U3071);
  nand ginst3681 (R1192_U324, R1192_U322, R1192_U323);
  nand ginst3682 (R1192_U325, R1192_U168, R1192_U324);
  nand ginst3683 (R1192_U326, R1192_U107, R1192_U212);
  nand ginst3684 (R1192_U327, R1192_U92, U3498);
  nand ginst3685 (R1192_U328, R1192_U167, R1192_U326);
  nand ginst3686 (R1192_U329, R1192_U80, U3071);
  not ginst3687 (R1192_U33, U3067);
  nand ginst3688 (R1192_U330, R1192_U212, R1192_U329);
  nand ginst3689 (R1192_U331, R1192_U280, R1192_U95);
  nand ginst3690 (R1192_U332, R1192_U88, U3059);
  nand ginst3691 (R1192_U333, R1192_U332, R1192_U373);
  nand ginst3692 (R1192_U334, R1192_U172, R1192_U333);
  nand ginst3693 (R1192_U335, R1192_U108, R1192_U211);
  nand ginst3694 (R1192_U336, R1192_U85, U3488);
  nand ginst3695 (R1192_U337, R1192_U171, R1192_U335);
  nand ginst3696 (R1192_U338, R1192_U88, U3059);
  nand ginst3697 (R1192_U339, R1192_U211, R1192_U338);
  nand ginst3698 (R1192_U34, R1192_U39, U3067);
  nand ginst3699 (R1192_U340, R1192_U45, U3074);
  nand ginst3700 (R1192_U341, R1192_U194, U3075);
  nand ginst3701 (R1192_U342, R1192_U97, U3079);
  nand ginst3702 (R1192_U343, R1192_U150, R1192_U151, R1192_U306);
  nand ginst3703 (R1192_U344, R1192_U184, R1192_U205);
  nand ginst3704 (R1192_U345, R1192_U133, R1192_U178);
  nand ginst3705 (R1192_U346, R1192_U14, R1192_U237);
  nand ginst3706 (R1192_U347, R1192_U270, R1192_U272);
  not ginst3707 (R1192_U348, R1192_U91);
  nand ginst3708 (R1192_U349, R1192_U273, R1192_U348);
  not ginst3709 (R1192_U35, U3081);
  nand ginst3710 (R1192_U350, R1192_U143, R1192_U201);
  nand ginst3711 (R1192_U351, R1192_U283, R1192_U285);
  nand ginst3712 (R1192_U352, R1192_U290, R1192_U291);
  not ginst3713 (R1192_U353, R1192_U105);
  nand ginst3714 (R1192_U354, R1192_U105, R1192_U17);
  not ginst3715 (R1192_U355, R1192_U104);
  nand ginst3716 (R1192_U356, R1192_U104, R1192_U301);
  not ginst3717 (R1192_U357, R1192_U103);
  nand ginst3718 (R1192_U358, R1192_U103, R1192_U303);
  nand ginst3719 (R1192_U359, R1192_U157, R1192_U192);
  not ginst3720 (R1192_U36, U3476);
  nand ginst3721 (R1192_U360, R1192_U105, R1192_U298);
  nand ginst3722 (R1192_U361, R1192_U196, R1192_U289);
  not ginst3723 (R1192_U362, R1192_U193);
  nand ginst3724 (R1192_U363, R1192_U19, R1192_U196);
  not ginst3725 (R1192_U364, R1192_U192);
  nand ginst3726 (R1192_U365, R1192_U196, R1192_U20);
  not ginst3727 (R1192_U366, R1192_U188);
  nand ginst3728 (R1192_U367, R1192_U196, R1192_U21);
  not ginst3729 (R1192_U368, R1192_U187);
  nand ginst3730 (R1192_U369, R1192_U160, R1192_U196);
  not ginst3731 (R1192_U37, U3478);
  nand ginst3732 (R1192_U370, R1192_U145, R1192_U196);
  not ginst3733 (R1192_U371, R1192_U186);
  nand ginst3734 (R1192_U372, R1192_U174, R1192_U244);
  not ginst3735 (R1192_U373, R1192_U108);
  nand ginst3736 (R1192_U374, R1192_U15, R1192_U174);
  not ginst3737 (R1192_U375, R1192_U203);
  nand ginst3738 (R1192_U376, R1192_U174, R1192_U18);
  not ginst3739 (R1192_U377, R1192_U202);
  nand ginst3740 (R1192_U378, R1192_U142, R1192_U174);
  not ginst3741 (R1192_U379, R1192_U201);
  not ginst3742 (R1192_U38, U3474);
  nand ginst3743 (R1192_U380, R1192_U131, R1192_U57);
  not ginst3744 (R1192_U381, R1192_U178);
  nand ginst3745 (R1192_U382, R1192_U215, R1192_U57);
  nand ginst3746 (R1192_U383, R1192_U140, R1192_U382);
  nand ginst3747 (R1192_U384, R1192_U224, R1192_U42);
  nand ginst3748 (R1192_U385, R1192_U197, R1192_U288);
  not ginst3749 (R1192_U386, R1192_U196);
  nand ginst3750 (R1192_U387, R1192_U12, R1192_U158);
  nand ginst3751 (R1192_U388, R1192_U159, R1192_U457);
  nand ginst3752 (R1192_U389, R1192_U54, U3484);
  not ginst3753 (R1192_U39, U3480);
  nand ginst3754 (R1192_U390, R1192_U53, U3080);
  nand ginst3755 (R1192_U391, R1192_U174, R1192_U245);
  nand ginst3756 (R1192_U392, R1192_U173, R1192_U243);
  nand ginst3757 (R1192_U393, R1192_U35, U3482);
  nand ginst3758 (R1192_U394, R1192_U40, U3081);
  nand ginst3759 (R1192_U395, R1192_U35, U3482);
  nand ginst3760 (R1192_U396, R1192_U40, U3081);
  nand ginst3761 (R1192_U397, R1192_U395, R1192_U396);
  nand ginst3762 (R1192_U398, R1192_U33, U3480);
  nand ginst3763 (R1192_U399, R1192_U39, U3067);
  not ginst3764 (R1192_U40, U3482);
  nand ginst3765 (R1192_U400, R1192_U250, R1192_U55);
  nand ginst3766 (R1192_U401, R1192_U175, R1192_U238);
  nand ginst3767 (R1192_U402, R1192_U48, U3478);
  nand ginst3768 (R1192_U403, R1192_U37, U3068);
  nand ginst3769 (R1192_U404, R1192_U402, R1192_U403);
  nand ginst3770 (R1192_U405, R1192_U49, U3476);
  nand ginst3771 (R1192_U406, R1192_U36, U3064);
  nand ginst3772 (R1192_U407, R1192_U260, R1192_U56);
  nand ginst3773 (R1192_U408, R1192_U176, R1192_U252);
  nand ginst3774 (R1192_U409, R1192_U50, U3474);
  not ginst3775 (R1192_U41, U3065);
  nand ginst3776 (R1192_U410, R1192_U38, U3057);
  nand ginst3777 (R1192_U411, R1192_U178, R1192_U261);
  nand ginst3778 (R1192_U412, R1192_U177, R1192_U381);
  nand ginst3779 (R1192_U413, R1192_U43, U3472);
  nand ginst3780 (R1192_U414, R1192_U47, U3061);
  nand ginst3781 (R1192_U415, R1192_U43, U3472);
  nand ginst3782 (R1192_U416, R1192_U47, U3061);
  nand ginst3783 (R1192_U417, R1192_U415, R1192_U416);
  nand ginst3784 (R1192_U418, R1192_U41, U3470);
  nand ginst3785 (R1192_U419, R1192_U44, U3065);
  nand ginst3786 (R1192_U42, R1192_U44, U3065);
  nand ginst3787 (R1192_U420, R1192_U263, R1192_U57);
  nand ginst3788 (R1192_U421, R1192_U179, R1192_U224);
  nand ginst3789 (R1192_U422, R1192_U181, U4040);
  nand ginst3790 (R1192_U423, R1192_U180, U3052);
  nand ginst3791 (R1192_U424, R1192_U181, U4040);
  nand ginst3792 (R1192_U425, R1192_U180, U3052);
  nand ginst3793 (R1192_U426, R1192_U424, R1192_U425);
  nand ginst3794 (R1192_U427, R1192_U102, R1192_U23, U4029);
  nand ginst3795 (R1192_U428, R1192_U101, R1192_U426, U3051);
  nand ginst3796 (R1192_U429, R1192_U102, U4029);
  not ginst3797 (R1192_U43, U3061);
  nand ginst3798 (R1192_U430, R1192_U101, U3051);
  not ginst3799 (R1192_U431, R1192_U152);
  nand ginst3800 (R1192_U432, R1192_U310, R1192_U431);
  nand ginst3801 (R1192_U433, R1192_U152, R1192_U183);
  nand ginst3802 (R1192_U434, R1192_U100, U4030);
  nand ginst3803 (R1192_U435, R1192_U59, U3050);
  nand ginst3804 (R1192_U436, R1192_U434, R1192_U435);
  nand ginst3805 (R1192_U437, R1192_U100, U4030);
  nand ginst3806 (R1192_U438, R1192_U59, U3050);
  nand ginst3807 (R1192_U439, R1192_U437, R1192_U438, R1192_U99);
  not ginst3808 (R1192_U44, U3470);
  nand ginst3809 (R1192_U440, R1192_U208, R1192_U436);
  nand ginst3810 (R1192_U441, R1192_U98, U4031);
  nand ginst3811 (R1192_U442, R1192_U58, U3054);
  nand ginst3812 (R1192_U443, R1192_U186, R1192_U314);
  nand ginst3813 (R1192_U444, R1192_U185, R1192_U371);
  nand ginst3814 (R1192_U445, R1192_U60, U4032);
  nand ginst3815 (R1192_U446, R1192_U61, U3055);
  not ginst3816 (R1192_U447, R1192_U155);
  nand ginst3817 (R1192_U448, R1192_U368, R1192_U447);
  nand ginst3818 (R1192_U449, R1192_U155, R1192_U187);
  not ginst3819 (R1192_U45, U3464);
  nand ginst3820 (R1192_U450, R1192_U62, U4033);
  nand ginst3821 (R1192_U451, R1192_U63, U3062);
  not ginst3822 (R1192_U452, R1192_U156);
  nand ginst3823 (R1192_U453, R1192_U366, R1192_U452);
  nand ginst3824 (R1192_U454, R1192_U156, R1192_U188);
  nand ginst3825 (R1192_U455, R1192_U64, U4034);
  nand ginst3826 (R1192_U456, R1192_U67, U3063);
  nand ginst3827 (R1192_U457, R1192_U455, R1192_U456);
  nand ginst3828 (R1192_U458, R1192_U161, R1192_U369, R1192_U69);
  nand ginst3829 (R1192_U459, R1192_U219, R1192_U22);
  not ginst3830 (R1192_U46, U3075);
  nand ginst3831 (R1192_U460, R1192_U65, U4035);
  nand ginst3832 (R1192_U461, R1192_U68, U3058);
  nand ginst3833 (R1192_U462, R1192_U190, R1192_U319);
  nand ginst3834 (R1192_U463, R1192_U189, R1192_U316);
  nand ginst3835 (R1192_U464, R1192_U66, U4036);
  nand ginst3836 (R1192_U465, R1192_U70, U3072);
  nand ginst3837 (R1192_U466, R1192_U192, R1192_U320);
  nand ginst3838 (R1192_U467, R1192_U191, R1192_U364);
  nand ginst3839 (R1192_U468, R1192_U71, U4037);
  nand ginst3840 (R1192_U469, R1192_U73, U3073);
  not ginst3841 (R1192_U47, U3472);
  not ginst3842 (R1192_U470, R1192_U162);
  nand ginst3843 (R1192_U471, R1192_U362, R1192_U470);
  nand ginst3844 (R1192_U472, R1192_U162, R1192_U193);
  nand ginst3845 (R1192_U473, R1192_U46, U3468);
  nand ginst3846 (R1192_U474, R1192_U194, U3075);
  not ginst3847 (R1192_U475, R1192_U163);
  nand ginst3848 (R1192_U476, R1192_U222, R1192_U475);
  nand ginst3849 (R1192_U477, R1192_U163, R1192_U195);
  nand ginst3850 (R1192_U478, R1192_U72, U3504);
  nand ginst3851 (R1192_U479, R1192_U75, U3078);
  not ginst3852 (R1192_U48, U3068);
  not ginst3853 (R1192_U480, R1192_U164);
  nand ginst3854 (R1192_U481, R1192_U386, R1192_U480);
  nand ginst3855 (R1192_U482, R1192_U164, R1192_U196);
  nand ginst3856 (R1192_U483, R1192_U76, U3502);
  nand ginst3857 (R1192_U484, R1192_U97, U3079);
  not ginst3858 (R1192_U485, R1192_U165);
  nand ginst3859 (R1192_U486, R1192_U287, R1192_U485);
  nand ginst3860 (R1192_U487, R1192_U165, R1192_U197);
  nand ginst3861 (R1192_U488, R1192_U77, U3500);
  nand ginst3862 (R1192_U489, R1192_U78, U3066);
  not ginst3863 (R1192_U49, U3064);
  not ginst3864 (R1192_U490, R1192_U166);
  nand ginst3865 (R1192_U491, R1192_U284, R1192_U490);
  nand ginst3866 (R1192_U492, R1192_U166, R1192_U198);
  nand ginst3867 (R1192_U493, R1192_U92, U3498);
  nand ginst3868 (R1192_U494, R1192_U79, U3070);
  nand ginst3869 (R1192_U495, R1192_U493, R1192_U494);
  nand ginst3870 (R1192_U496, R1192_U93, U3496);
  nand ginst3871 (R1192_U497, R1192_U80, U3071);
  nand ginst3872 (R1192_U498, R1192_U107, R1192_U330);
  nand ginst3873 (R1192_U499, R1192_U199, R1192_U322);
  not ginst3874 (R1192_U50, U3057);
  nand ginst3875 (R1192_U500, R1192_U94, U3494);
  nand ginst3876 (R1192_U501, R1192_U81, U3076);
  nand ginst3877 (R1192_U502, R1192_U201, R1192_U331);
  nand ginst3878 (R1192_U503, R1192_U200, R1192_U379);
  nand ginst3879 (R1192_U504, R1192_U82, U3492);
  nand ginst3880 (R1192_U505, R1192_U83, U3077);
  not ginst3881 (R1192_U506, R1192_U169);
  nand ginst3882 (R1192_U507, R1192_U377, R1192_U506);
  nand ginst3883 (R1192_U508, R1192_U169, R1192_U202);
  nand ginst3884 (R1192_U509, R1192_U90, U3490);
  nand ginst3885 (R1192_U51, R1192_U38, U3057);
  nand ginst3886 (R1192_U510, R1192_U84, U3069);
  not ginst3887 (R1192_U511, R1192_U170);
  nand ginst3888 (R1192_U512, R1192_U375, R1192_U511);
  nand ginst3889 (R1192_U513, R1192_U170, R1192_U203);
  nand ginst3890 (R1192_U514, R1192_U85, U3488);
  nand ginst3891 (R1192_U515, R1192_U87, U3060);
  nand ginst3892 (R1192_U516, R1192_U514, R1192_U515);
  nand ginst3893 (R1192_U517, R1192_U86, U3486);
  nand ginst3894 (R1192_U518, R1192_U88, U3059);
  nand ginst3895 (R1192_U519, R1192_U108, R1192_U339);
  nand ginst3896 (R1192_U52, R1192_U233, R1192_U235);
  nand ginst3897 (R1192_U520, R1192_U204, R1192_U373);
  not ginst3898 (R1192_U53, U3484);
  not ginst3899 (R1192_U54, U3080);
  nand ginst3900 (R1192_U55, R1192_U236, R1192_U52);
  nand ginst3901 (R1192_U56, R1192_U251, R1192_U51);
  nand ginst3902 (R1192_U57, R1192_U207, R1192_U223, R1192_U341);
  not ginst3903 (R1192_U58, U4031);
  not ginst3904 (R1192_U59, U4030);
  and ginst3905 (R1192_U6, R1192_U230, R1192_U231);
  not ginst3906 (R1192_U60, U3055);
  not ginst3907 (R1192_U61, U4032);
  not ginst3908 (R1192_U62, U3062);
  not ginst3909 (R1192_U63, U4033);
  not ginst3910 (R1192_U64, U3063);
  not ginst3911 (R1192_U65, U3058);
  not ginst3912 (R1192_U66, U3072);
  not ginst3913 (R1192_U67, U4034);
  not ginst3914 (R1192_U68, U4035);
  nand ginst3915 (R1192_U69, R1192_U70, U3072);
  and ginst3916 (R1192_U7, R1192_U211, R1192_U264);
  not ginst3917 (R1192_U70, U4036);
  not ginst3918 (R1192_U71, U3073);
  not ginst3919 (R1192_U72, U3078);
  not ginst3920 (R1192_U73, U4037);
  nand ginst3921 (R1192_U74, R1192_U75, U3078);
  not ginst3922 (R1192_U75, U3504);
  not ginst3923 (R1192_U76, U3079);
  not ginst3924 (R1192_U77, U3066);
  not ginst3925 (R1192_U78, U3500);
  not ginst3926 (R1192_U79, U3498);
  and ginst3927 (R1192_U8, R1192_U265, R1192_U266);
  not ginst3928 (R1192_U80, U3496);
  not ginst3929 (R1192_U81, U3494);
  not ginst3930 (R1192_U82, U3077);
  not ginst3931 (R1192_U83, U3492);
  not ginst3932 (R1192_U84, U3490);
  not ginst3933 (R1192_U85, U3060);
  not ginst3934 (R1192_U86, U3059);
  not ginst3935 (R1192_U87, U3488);
  not ginst3936 (R1192_U88, U3486);
  nand ginst3937 (R1192_U89, R1192_U53, U3080);
  and ginst3938 (R1192_U9, R1192_U212, R1192_U275);
  not ginst3939 (R1192_U90, U3069);
  nand ginst3940 (R1192_U91, R1192_U271, R1192_U347);
  not ginst3941 (R1192_U92, U3070);
  not ginst3942 (R1192_U93, U3071);
  not ginst3943 (R1192_U94, U3076);
  nand ginst3944 (R1192_U95, R1192_U81, U3076);
  nand ginst3945 (R1192_U96, R1192_U279, R1192_U281);
  not ginst3946 (R1192_U97, U3502);
  not ginst3947 (R1192_U98, U3054);
  nand ginst3948 (R1192_U99, R1192_U58, U3054);
  and ginst3949 (R1207_U10, R1207_U276, R1207_U277);
  not ginst3950 (R1207_U100, U3050);
  not ginst3951 (R1207_U101, U4029);
  not ginst3952 (R1207_U102, U3051);
  nand ginst3953 (R1207_U103, R1207_U302, R1207_U356);
  nand ginst3954 (R1207_U104, R1207_U300, R1207_U354);
  nand ginst3955 (R1207_U105, R1207_U292, R1207_U352);
  nand ginst3956 (R1207_U106, R1207_U65, U4035);
  nand ginst3957 (R1207_U107, R1207_U321, R1207_U95);
  nand ginst3958 (R1207_U108, R1207_U372, R1207_U89);
  not ginst3959 (R1207_U109, U3074);
  and ginst3960 (R1207_U11, R1207_U106, R1207_U293);
  nand ginst3961 (R1207_U110, R1207_U432, R1207_U433);
  nand ginst3962 (R1207_U111, R1207_U448, R1207_U449);
  nand ginst3963 (R1207_U112, R1207_U453, R1207_U454);
  nand ginst3964 (R1207_U113, R1207_U471, R1207_U472);
  nand ginst3965 (R1207_U114, R1207_U476, R1207_U477);
  nand ginst3966 (R1207_U115, R1207_U481, R1207_U482);
  nand ginst3967 (R1207_U116, R1207_U486, R1207_U487);
  nand ginst3968 (R1207_U117, R1207_U491, R1207_U492);
  nand ginst3969 (R1207_U118, R1207_U507, R1207_U508);
  nand ginst3970 (R1207_U119, R1207_U512, R1207_U513);
  and ginst3971 (R1207_U12, R1207_U294, R1207_U295);
  nand ginst3972 (R1207_U120, R1207_U391, R1207_U392);
  nand ginst3973 (R1207_U121, R1207_U400, R1207_U401);
  nand ginst3974 (R1207_U122, R1207_U407, R1207_U408);
  nand ginst3975 (R1207_U123, R1207_U411, R1207_U412);
  nand ginst3976 (R1207_U124, R1207_U420, R1207_U421);
  nand ginst3977 (R1207_U125, R1207_U443, R1207_U444);
  nand ginst3978 (R1207_U126, R1207_U462, R1207_U463);
  nand ginst3979 (R1207_U127, R1207_U466, R1207_U467);
  nand ginst3980 (R1207_U128, R1207_U498, R1207_U499);
  nand ginst3981 (R1207_U129, R1207_U502, R1207_U503);
  and ginst3982 (R1207_U13, R1207_U216, R1207_U229, R1207_U234);
  nand ginst3983 (R1207_U130, R1207_U519, R1207_U520);
  and ginst3984 (R1207_U131, R1207_U215, R1207_U225);
  and ginst3985 (R1207_U132, R1207_U227, R1207_U228);
  and ginst3986 (R1207_U133, R1207_U13, R1207_U14);
  and ginst3987 (R1207_U134, R1207_U241, R1207_U242);
  and ginst3988 (R1207_U135, R1207_U134, R1207_U346);
  and ginst3989 (R1207_U136, R1207_U34, R1207_U393, R1207_U394);
  and ginst3990 (R1207_U137, R1207_U217, R1207_U397);
  and ginst3991 (R1207_U138, R1207_U257, R1207_U6);
  and ginst3992 (R1207_U139, R1207_U216, R1207_U404);
  and ginst3993 (R1207_U14, R1207_U217, R1207_U239);
  and ginst3994 (R1207_U140, R1207_U413, R1207_U414, R1207_U42);
  and ginst3995 (R1207_U141, R1207_U215, R1207_U417);
  and ginst3996 (R1207_U142, R1207_U18, R1207_U273);
  and ginst3997 (R1207_U143, R1207_U16, R1207_U285);
  and ginst3998 (R1207_U144, R1207_U286, R1207_U351);
  and ginst3999 (R1207_U145, R1207_U21, R1207_U303);
  and ginst4000 (R1207_U146, R1207_U304, R1207_U358);
  and ginst4001 (R1207_U147, R1207_U214, R1207_U305);
  and ginst4002 (R1207_U148, R1207_U308, R1207_U309);
  and ginst4003 (R1207_U149, R1207_U311, R1207_U426);
  and ginst4004 (R1207_U15, R1207_U244, R1207_U7);
  and ginst4005 (R1207_U150, R1207_U308, R1207_U309);
  and ginst4006 (R1207_U151, R1207_U23, R1207_U312);
  nand ginst4007 (R1207_U152, R1207_U429, R1207_U430);
  and ginst4008 (R1207_U153, R1207_U214, R1207_U436);
  and ginst4009 (R1207_U154, R1207_U186, R1207_U214);
  nand ginst4010 (R1207_U155, R1207_U445, R1207_U446);
  nand ginst4011 (R1207_U156, R1207_U450, R1207_U451);
  and ginst4012 (R1207_U157, R1207_U22, R1207_U298);
  and ginst4013 (R1207_U158, R1207_U213, R1207_U317);
  and ginst4014 (R1207_U159, R1207_U68, U3058);
  and ginst4015 (R1207_U16, R1207_U280, R1207_U9);
  and ginst4016 (R1207_U160, R1207_U19, R1207_U298);
  and ginst4017 (R1207_U161, R1207_U12, R1207_U317, R1207_U360);
  nand ginst4018 (R1207_U162, R1207_U468, R1207_U469);
  nand ginst4019 (R1207_U163, R1207_U473, R1207_U474);
  nand ginst4020 (R1207_U164, R1207_U478, R1207_U479);
  nand ginst4021 (R1207_U165, R1207_U483, R1207_U484);
  nand ginst4022 (R1207_U166, R1207_U488, R1207_U489);
  and ginst4023 (R1207_U167, R1207_U10, R1207_U327);
  and ginst4024 (R1207_U168, R1207_U212, R1207_U495);
  nand ginst4025 (R1207_U169, R1207_U504, R1207_U505);
  and ginst4026 (R1207_U17, R1207_U11, R1207_U298);
  nand ginst4027 (R1207_U170, R1207_U509, R1207_U510);
  and ginst4028 (R1207_U171, R1207_U336, R1207_U8);
  and ginst4029 (R1207_U172, R1207_U211, R1207_U516);
  and ginst4030 (R1207_U173, R1207_U389, R1207_U390);
  nand ginst4031 (R1207_U174, R1207_U135, R1207_U345);
  and ginst4032 (R1207_U175, R1207_U398, R1207_U399);
  and ginst4033 (R1207_U176, R1207_U405, R1207_U406);
  and ginst4034 (R1207_U177, R1207_U409, R1207_U410);
  nand ginst4035 (R1207_U178, R1207_U132, R1207_U380);
  and ginst4036 (R1207_U179, R1207_U418, R1207_U419);
  and ginst4037 (R1207_U18, R1207_U15, R1207_U271);
  not ginst4038 (R1207_U180, U4040);
  not ginst4039 (R1207_U181, U3052);
  and ginst4040 (R1207_U182, R1207_U427, R1207_U428);
  nand ginst4041 (R1207_U183, R1207_U148, R1207_U306);
  and ginst4042 (R1207_U184, R1207_U439, R1207_U440);
  and ginst4043 (R1207_U185, R1207_U441, R1207_U442);
  nand ginst4044 (R1207_U186, R1207_U146, R1207_U370);
  nand ginst4045 (R1207_U187, R1207_U357, R1207_U367);
  nand ginst4046 (R1207_U188, R1207_U355, R1207_U365);
  and ginst4047 (R1207_U189, R1207_U460, R1207_U461);
  and ginst4048 (R1207_U19, R1207_U289, R1207_U291);
  nand ginst4049 (R1207_U190, R1207_U315, R1207_U69);
  and ginst4050 (R1207_U191, R1207_U464, R1207_U465);
  nand ginst4051 (R1207_U192, R1207_U353, R1207_U363);
  nand ginst4052 (R1207_U193, R1207_U361, R1207_U74);
  not ginst4053 (R1207_U194, U3468);
  nand ginst4054 (R1207_U195, R1207_U109, U3464);
  nand ginst4055 (R1207_U196, R1207_U342, R1207_U385);
  nand ginst4056 (R1207_U197, R1207_U144, R1207_U350);
  nand ginst4057 (R1207_U198, R1207_U282, R1207_U96);
  and ginst4058 (R1207_U199, R1207_U496, R1207_U497);
  and ginst4059 (R1207_U20, R1207_U17, R1207_U19);
  and ginst4060 (R1207_U200, R1207_U500, R1207_U501);
  nand ginst4061 (R1207_U201, R1207_U274, R1207_U349, R1207_U378);
  nand ginst4062 (R1207_U202, R1207_U376, R1207_U91);
  nand ginst4063 (R1207_U203, R1207_U270, R1207_U374);
  and ginst4064 (R1207_U204, R1207_U517, R1207_U518);
  nand ginst4065 (R1207_U205, R1207_U153, R1207_U186);
  nand ginst4066 (R1207_U206, R1207_U149, R1207_U183);
  nand ginst4067 (R1207_U207, R1207_U194, R1207_U195);
  not ginst4068 (R1207_U208, R1207_U99);
  not ginst4069 (R1207_U209, R1207_U42);
  and ginst4070 (R1207_U21, R1207_U20, R1207_U301);
  not ginst4071 (R1207_U210, R1207_U34);
  nand ginst4072 (R1207_U211, R1207_U86, U3486);
  nand ginst4073 (R1207_U212, R1207_U93, U3496);
  not ginst4074 (R1207_U213, R1207_U106);
  nand ginst4075 (R1207_U214, R1207_U98, U4031);
  nand ginst4076 (R1207_U215, R1207_U41, U3470);
  nand ginst4077 (R1207_U216, R1207_U49, U3476);
  nand ginst4078 (R1207_U217, R1207_U33, U3480);
  not ginst4079 (R1207_U218, R1207_U95);
  not ginst4080 (R1207_U219, R1207_U69);
  and ginst4081 (R1207_U22, R1207_U106, R1207_U457);
  not ginst4082 (R1207_U220, R1207_U51);
  not ginst4083 (R1207_U221, R1207_U89);
  not ginst4084 (R1207_U222, R1207_U195);
  nand ginst4085 (R1207_U223, R1207_U195, U3075);
  not ginst4086 (R1207_U224, R1207_U57);
  nand ginst4087 (R1207_U225, R1207_U43, U3472);
  nand ginst4088 (R1207_U226, R1207_U42, R1207_U43);
  nand ginst4089 (R1207_U227, R1207_U226, R1207_U47);
  nand ginst4090 (R1207_U228, R1207_U209, U3061);
  nand ginst4091 (R1207_U229, R1207_U48, U3478);
  and ginst4092 (R1207_U23, R1207_U422, R1207_U423);
  nand ginst4093 (R1207_U230, R1207_U37, U3068);
  nand ginst4094 (R1207_U231, R1207_U36, U3064);
  nand ginst4095 (R1207_U232, R1207_U216, R1207_U220);
  nand ginst4096 (R1207_U233, R1207_U232, R1207_U6);
  nand ginst4097 (R1207_U234, R1207_U50, U3474);
  nand ginst4098 (R1207_U235, R1207_U48, U3478);
  nand ginst4099 (R1207_U236, R1207_U13, R1207_U178);
  not ginst4100 (R1207_U237, R1207_U52);
  not ginst4101 (R1207_U238, R1207_U55);
  nand ginst4102 (R1207_U239, R1207_U35, U3482);
  nand ginst4103 (R1207_U24, R1207_U334, R1207_U337);
  nand ginst4104 (R1207_U240, R1207_U34, R1207_U35);
  nand ginst4105 (R1207_U241, R1207_U240, R1207_U40);
  nand ginst4106 (R1207_U242, R1207_U210, U3081);
  not ginst4107 (R1207_U243, R1207_U174);
  nand ginst4108 (R1207_U244, R1207_U54, U3484);
  nand ginst4109 (R1207_U245, R1207_U244, R1207_U89);
  nand ginst4110 (R1207_U246, R1207_U238, R1207_U34);
  nand ginst4111 (R1207_U247, R1207_U137, R1207_U246);
  nand ginst4112 (R1207_U248, R1207_U217, R1207_U55);
  nand ginst4113 (R1207_U249, R1207_U136, R1207_U248);
  nand ginst4114 (R1207_U25, R1207_U325, R1207_U328);
  nand ginst4115 (R1207_U250, R1207_U217, R1207_U34);
  nand ginst4116 (R1207_U251, R1207_U178, R1207_U234);
  not ginst4117 (R1207_U252, R1207_U56);
  nand ginst4118 (R1207_U253, R1207_U36, U3064);
  nand ginst4119 (R1207_U254, R1207_U252, R1207_U253);
  nand ginst4120 (R1207_U255, R1207_U139, R1207_U254);
  nand ginst4121 (R1207_U256, R1207_U216, R1207_U56);
  nand ginst4122 (R1207_U257, R1207_U48, U3478);
  nand ginst4123 (R1207_U258, R1207_U138, R1207_U256);
  nand ginst4124 (R1207_U259, R1207_U36, U3064);
  nand ginst4125 (R1207_U26, R1207_U359, R1207_U387, R1207_U388, R1207_U458, R1207_U459);
  nand ginst4126 (R1207_U260, R1207_U216, R1207_U259);
  nand ginst4127 (R1207_U261, R1207_U234, R1207_U51);
  nand ginst4128 (R1207_U262, R1207_U141, R1207_U384);
  nand ginst4129 (R1207_U263, R1207_U215, R1207_U42);
  nand ginst4130 (R1207_U264, R1207_U85, U3488);
  nand ginst4131 (R1207_U265, R1207_U87, U3060);
  nand ginst4132 (R1207_U266, R1207_U88, U3059);
  nand ginst4133 (R1207_U267, R1207_U221, R1207_U7);
  nand ginst4134 (R1207_U268, R1207_U267, R1207_U8);
  nand ginst4135 (R1207_U269, R1207_U85, U3488);
  and ginst4136 (R1207_U27, R1207_U313, R1207_U344);
  nand ginst4137 (R1207_U270, R1207_U268, R1207_U269);
  nand ginst4138 (R1207_U271, R1207_U90, U3490);
  nand ginst4139 (R1207_U272, R1207_U84, U3069);
  nand ginst4140 (R1207_U273, R1207_U82, U3492);
  nand ginst4141 (R1207_U274, R1207_U83, U3077);
  nand ginst4142 (R1207_U275, R1207_U92, U3498);
  nand ginst4143 (R1207_U276, R1207_U79, U3070);
  nand ginst4144 (R1207_U277, R1207_U80, U3071);
  nand ginst4145 (R1207_U278, R1207_U218, R1207_U9);
  nand ginst4146 (R1207_U279, R1207_U10, R1207_U278);
  nand ginst4147 (R1207_U28, R1207_U182, R1207_U206, R1207_U343);
  nand ginst4148 (R1207_U280, R1207_U94, U3494);
  nand ginst4149 (R1207_U281, R1207_U92, U3498);
  nand ginst4150 (R1207_U282, R1207_U16, R1207_U201);
  not ginst4151 (R1207_U283, R1207_U96);
  not ginst4152 (R1207_U284, R1207_U198);
  nand ginst4153 (R1207_U285, R1207_U77, U3500);
  nand ginst4154 (R1207_U286, R1207_U78, U3066);
  not ginst4155 (R1207_U287, R1207_U197);
  nand ginst4156 (R1207_U288, R1207_U76, U3502);
  nand ginst4157 (R1207_U289, R1207_U72, U3504);
  nand ginst4158 (R1207_U29, R1207_U262, R1207_U383);
  not ginst4159 (R1207_U290, R1207_U74);
  nand ginst4160 (R1207_U291, R1207_U71, U4037);
  nand ginst4161 (R1207_U292, R1207_U73, U3073);
  nand ginst4162 (R1207_U293, R1207_U64, U4034);
  nand ginst4163 (R1207_U294, R1207_U67, U3063);
  nand ginst4164 (R1207_U295, R1207_U68, U3058);
  nand ginst4165 (R1207_U296, R1207_U11, R1207_U219);
  nand ginst4166 (R1207_U297, R1207_U12, R1207_U296);
  nand ginst4167 (R1207_U298, R1207_U66, U4036);
  nand ginst4168 (R1207_U299, R1207_U64, U4034);
  nand ginst4169 (R1207_U30, R1207_U255, R1207_U258);
  nand ginst4170 (R1207_U300, R1207_U297, R1207_U299);
  nand ginst4171 (R1207_U301, R1207_U62, U4033);
  nand ginst4172 (R1207_U302, R1207_U63, U3062);
  nand ginst4173 (R1207_U303, R1207_U60, U4032);
  nand ginst4174 (R1207_U304, R1207_U61, U3055);
  nand ginst4175 (R1207_U305, R1207_U100, U4030);
  nand ginst4176 (R1207_U306, R1207_U147, R1207_U186);
  nand ginst4177 (R1207_U307, R1207_U100, R1207_U99);
  nand ginst4178 (R1207_U308, R1207_U307, R1207_U59);
  nand ginst4179 (R1207_U309, R1207_U208, U3050);
  nand ginst4180 (R1207_U31, R1207_U247, R1207_U249);
  not ginst4181 (R1207_U310, R1207_U183);
  nand ginst4182 (R1207_U311, R1207_U102, U4029);
  nand ginst4183 (R1207_U312, R1207_U101, U3051);
  nand ginst4184 (R1207_U313, R1207_U154, R1207_U205);
  nand ginst4185 (R1207_U314, R1207_U214, R1207_U99);
  nand ginst4186 (R1207_U315, R1207_U192, R1207_U298);
  not ginst4187 (R1207_U316, R1207_U190);
  nand ginst4188 (R1207_U317, R1207_U64, U4034);
  nand ginst4189 (R1207_U318, R1207_U68, U3058);
  nand ginst4190 (R1207_U319, R1207_U106, R1207_U318);
  nand ginst4191 (R1207_U32, R1207_U195, R1207_U340);
  nand ginst4192 (R1207_U320, R1207_U298, R1207_U69);
  nand ginst4193 (R1207_U321, R1207_U201, R1207_U280);
  not ginst4194 (R1207_U322, R1207_U107);
  nand ginst4195 (R1207_U323, R1207_U80, U3071);
  nand ginst4196 (R1207_U324, R1207_U322, R1207_U323);
  nand ginst4197 (R1207_U325, R1207_U168, R1207_U324);
  nand ginst4198 (R1207_U326, R1207_U107, R1207_U212);
  nand ginst4199 (R1207_U327, R1207_U92, U3498);
  nand ginst4200 (R1207_U328, R1207_U167, R1207_U326);
  nand ginst4201 (R1207_U329, R1207_U80, U3071);
  not ginst4202 (R1207_U33, U3067);
  nand ginst4203 (R1207_U330, R1207_U212, R1207_U329);
  nand ginst4204 (R1207_U331, R1207_U280, R1207_U95);
  nand ginst4205 (R1207_U332, R1207_U88, U3059);
  nand ginst4206 (R1207_U333, R1207_U332, R1207_U373);
  nand ginst4207 (R1207_U334, R1207_U172, R1207_U333);
  nand ginst4208 (R1207_U335, R1207_U108, R1207_U211);
  nand ginst4209 (R1207_U336, R1207_U85, U3488);
  nand ginst4210 (R1207_U337, R1207_U171, R1207_U335);
  nand ginst4211 (R1207_U338, R1207_U88, U3059);
  nand ginst4212 (R1207_U339, R1207_U211, R1207_U338);
  nand ginst4213 (R1207_U34, R1207_U39, U3067);
  nand ginst4214 (R1207_U340, R1207_U45, U3074);
  nand ginst4215 (R1207_U341, R1207_U194, U3075);
  nand ginst4216 (R1207_U342, R1207_U97, U3079);
  nand ginst4217 (R1207_U343, R1207_U150, R1207_U151, R1207_U306);
  nand ginst4218 (R1207_U344, R1207_U184, R1207_U205);
  nand ginst4219 (R1207_U345, R1207_U133, R1207_U178);
  nand ginst4220 (R1207_U346, R1207_U14, R1207_U237);
  nand ginst4221 (R1207_U347, R1207_U270, R1207_U272);
  not ginst4222 (R1207_U348, R1207_U91);
  nand ginst4223 (R1207_U349, R1207_U273, R1207_U348);
  not ginst4224 (R1207_U35, U3081);
  nand ginst4225 (R1207_U350, R1207_U143, R1207_U201);
  nand ginst4226 (R1207_U351, R1207_U283, R1207_U285);
  nand ginst4227 (R1207_U352, R1207_U290, R1207_U291);
  not ginst4228 (R1207_U353, R1207_U105);
  nand ginst4229 (R1207_U354, R1207_U105, R1207_U17);
  not ginst4230 (R1207_U355, R1207_U104);
  nand ginst4231 (R1207_U356, R1207_U104, R1207_U301);
  not ginst4232 (R1207_U357, R1207_U103);
  nand ginst4233 (R1207_U358, R1207_U103, R1207_U303);
  nand ginst4234 (R1207_U359, R1207_U157, R1207_U192);
  not ginst4235 (R1207_U36, U3476);
  nand ginst4236 (R1207_U360, R1207_U105, R1207_U298);
  nand ginst4237 (R1207_U361, R1207_U196, R1207_U289);
  not ginst4238 (R1207_U362, R1207_U193);
  nand ginst4239 (R1207_U363, R1207_U19, R1207_U196);
  not ginst4240 (R1207_U364, R1207_U192);
  nand ginst4241 (R1207_U365, R1207_U196, R1207_U20);
  not ginst4242 (R1207_U366, R1207_U188);
  nand ginst4243 (R1207_U367, R1207_U196, R1207_U21);
  not ginst4244 (R1207_U368, R1207_U187);
  nand ginst4245 (R1207_U369, R1207_U160, R1207_U196);
  not ginst4246 (R1207_U37, U3478);
  nand ginst4247 (R1207_U370, R1207_U145, R1207_U196);
  not ginst4248 (R1207_U371, R1207_U186);
  nand ginst4249 (R1207_U372, R1207_U174, R1207_U244);
  not ginst4250 (R1207_U373, R1207_U108);
  nand ginst4251 (R1207_U374, R1207_U15, R1207_U174);
  not ginst4252 (R1207_U375, R1207_U203);
  nand ginst4253 (R1207_U376, R1207_U174, R1207_U18);
  not ginst4254 (R1207_U377, R1207_U202);
  nand ginst4255 (R1207_U378, R1207_U142, R1207_U174);
  not ginst4256 (R1207_U379, R1207_U201);
  not ginst4257 (R1207_U38, U3474);
  nand ginst4258 (R1207_U380, R1207_U131, R1207_U57);
  not ginst4259 (R1207_U381, R1207_U178);
  nand ginst4260 (R1207_U382, R1207_U215, R1207_U57);
  nand ginst4261 (R1207_U383, R1207_U140, R1207_U382);
  nand ginst4262 (R1207_U384, R1207_U224, R1207_U42);
  nand ginst4263 (R1207_U385, R1207_U197, R1207_U288);
  not ginst4264 (R1207_U386, R1207_U196);
  nand ginst4265 (R1207_U387, R1207_U12, R1207_U158);
  nand ginst4266 (R1207_U388, R1207_U159, R1207_U457);
  nand ginst4267 (R1207_U389, R1207_U54, U3484);
  not ginst4268 (R1207_U39, U3480);
  nand ginst4269 (R1207_U390, R1207_U53, U3080);
  nand ginst4270 (R1207_U391, R1207_U174, R1207_U245);
  nand ginst4271 (R1207_U392, R1207_U173, R1207_U243);
  nand ginst4272 (R1207_U393, R1207_U35, U3482);
  nand ginst4273 (R1207_U394, R1207_U40, U3081);
  nand ginst4274 (R1207_U395, R1207_U35, U3482);
  nand ginst4275 (R1207_U396, R1207_U40, U3081);
  nand ginst4276 (R1207_U397, R1207_U395, R1207_U396);
  nand ginst4277 (R1207_U398, R1207_U33, U3480);
  nand ginst4278 (R1207_U399, R1207_U39, U3067);
  not ginst4279 (R1207_U40, U3482);
  nand ginst4280 (R1207_U400, R1207_U250, R1207_U55);
  nand ginst4281 (R1207_U401, R1207_U175, R1207_U238);
  nand ginst4282 (R1207_U402, R1207_U48, U3478);
  nand ginst4283 (R1207_U403, R1207_U37, U3068);
  nand ginst4284 (R1207_U404, R1207_U402, R1207_U403);
  nand ginst4285 (R1207_U405, R1207_U49, U3476);
  nand ginst4286 (R1207_U406, R1207_U36, U3064);
  nand ginst4287 (R1207_U407, R1207_U260, R1207_U56);
  nand ginst4288 (R1207_U408, R1207_U176, R1207_U252);
  nand ginst4289 (R1207_U409, R1207_U50, U3474);
  not ginst4290 (R1207_U41, U3065);
  nand ginst4291 (R1207_U410, R1207_U38, U3057);
  nand ginst4292 (R1207_U411, R1207_U178, R1207_U261);
  nand ginst4293 (R1207_U412, R1207_U177, R1207_U381);
  nand ginst4294 (R1207_U413, R1207_U43, U3472);
  nand ginst4295 (R1207_U414, R1207_U47, U3061);
  nand ginst4296 (R1207_U415, R1207_U43, U3472);
  nand ginst4297 (R1207_U416, R1207_U47, U3061);
  nand ginst4298 (R1207_U417, R1207_U415, R1207_U416);
  nand ginst4299 (R1207_U418, R1207_U41, U3470);
  nand ginst4300 (R1207_U419, R1207_U44, U3065);
  nand ginst4301 (R1207_U42, R1207_U44, U3065);
  nand ginst4302 (R1207_U420, R1207_U263, R1207_U57);
  nand ginst4303 (R1207_U421, R1207_U179, R1207_U224);
  nand ginst4304 (R1207_U422, R1207_U181, U4040);
  nand ginst4305 (R1207_U423, R1207_U180, U3052);
  nand ginst4306 (R1207_U424, R1207_U181, U4040);
  nand ginst4307 (R1207_U425, R1207_U180, U3052);
  nand ginst4308 (R1207_U426, R1207_U424, R1207_U425);
  nand ginst4309 (R1207_U427, R1207_U102, R1207_U23, U4029);
  nand ginst4310 (R1207_U428, R1207_U101, R1207_U426, U3051);
  nand ginst4311 (R1207_U429, R1207_U102, U4029);
  not ginst4312 (R1207_U43, U3061);
  nand ginst4313 (R1207_U430, R1207_U101, U3051);
  not ginst4314 (R1207_U431, R1207_U152);
  nand ginst4315 (R1207_U432, R1207_U310, R1207_U431);
  nand ginst4316 (R1207_U433, R1207_U152, R1207_U183);
  nand ginst4317 (R1207_U434, R1207_U100, U4030);
  nand ginst4318 (R1207_U435, R1207_U59, U3050);
  nand ginst4319 (R1207_U436, R1207_U434, R1207_U435);
  nand ginst4320 (R1207_U437, R1207_U100, U4030);
  nand ginst4321 (R1207_U438, R1207_U59, U3050);
  nand ginst4322 (R1207_U439, R1207_U437, R1207_U438, R1207_U99);
  not ginst4323 (R1207_U44, U3470);
  nand ginst4324 (R1207_U440, R1207_U208, R1207_U436);
  nand ginst4325 (R1207_U441, R1207_U98, U4031);
  nand ginst4326 (R1207_U442, R1207_U58, U3054);
  nand ginst4327 (R1207_U443, R1207_U186, R1207_U314);
  nand ginst4328 (R1207_U444, R1207_U185, R1207_U371);
  nand ginst4329 (R1207_U445, R1207_U60, U4032);
  nand ginst4330 (R1207_U446, R1207_U61, U3055);
  not ginst4331 (R1207_U447, R1207_U155);
  nand ginst4332 (R1207_U448, R1207_U368, R1207_U447);
  nand ginst4333 (R1207_U449, R1207_U155, R1207_U187);
  not ginst4334 (R1207_U45, U3464);
  nand ginst4335 (R1207_U450, R1207_U62, U4033);
  nand ginst4336 (R1207_U451, R1207_U63, U3062);
  not ginst4337 (R1207_U452, R1207_U156);
  nand ginst4338 (R1207_U453, R1207_U366, R1207_U452);
  nand ginst4339 (R1207_U454, R1207_U156, R1207_U188);
  nand ginst4340 (R1207_U455, R1207_U64, U4034);
  nand ginst4341 (R1207_U456, R1207_U67, U3063);
  nand ginst4342 (R1207_U457, R1207_U455, R1207_U456);
  nand ginst4343 (R1207_U458, R1207_U161, R1207_U369, R1207_U69);
  nand ginst4344 (R1207_U459, R1207_U219, R1207_U22);
  not ginst4345 (R1207_U46, U3075);
  nand ginst4346 (R1207_U460, R1207_U65, U4035);
  nand ginst4347 (R1207_U461, R1207_U68, U3058);
  nand ginst4348 (R1207_U462, R1207_U190, R1207_U319);
  nand ginst4349 (R1207_U463, R1207_U189, R1207_U316);
  nand ginst4350 (R1207_U464, R1207_U66, U4036);
  nand ginst4351 (R1207_U465, R1207_U70, U3072);
  nand ginst4352 (R1207_U466, R1207_U192, R1207_U320);
  nand ginst4353 (R1207_U467, R1207_U191, R1207_U364);
  nand ginst4354 (R1207_U468, R1207_U71, U4037);
  nand ginst4355 (R1207_U469, R1207_U73, U3073);
  not ginst4356 (R1207_U47, U3472);
  not ginst4357 (R1207_U470, R1207_U162);
  nand ginst4358 (R1207_U471, R1207_U362, R1207_U470);
  nand ginst4359 (R1207_U472, R1207_U162, R1207_U193);
  nand ginst4360 (R1207_U473, R1207_U46, U3468);
  nand ginst4361 (R1207_U474, R1207_U194, U3075);
  not ginst4362 (R1207_U475, R1207_U163);
  nand ginst4363 (R1207_U476, R1207_U222, R1207_U475);
  nand ginst4364 (R1207_U477, R1207_U163, R1207_U195);
  nand ginst4365 (R1207_U478, R1207_U72, U3504);
  nand ginst4366 (R1207_U479, R1207_U75, U3078);
  not ginst4367 (R1207_U48, U3068);
  not ginst4368 (R1207_U480, R1207_U164);
  nand ginst4369 (R1207_U481, R1207_U386, R1207_U480);
  nand ginst4370 (R1207_U482, R1207_U164, R1207_U196);
  nand ginst4371 (R1207_U483, R1207_U76, U3502);
  nand ginst4372 (R1207_U484, R1207_U97, U3079);
  not ginst4373 (R1207_U485, R1207_U165);
  nand ginst4374 (R1207_U486, R1207_U287, R1207_U485);
  nand ginst4375 (R1207_U487, R1207_U165, R1207_U197);
  nand ginst4376 (R1207_U488, R1207_U77, U3500);
  nand ginst4377 (R1207_U489, R1207_U78, U3066);
  not ginst4378 (R1207_U49, U3064);
  not ginst4379 (R1207_U490, R1207_U166);
  nand ginst4380 (R1207_U491, R1207_U284, R1207_U490);
  nand ginst4381 (R1207_U492, R1207_U166, R1207_U198);
  nand ginst4382 (R1207_U493, R1207_U92, U3498);
  nand ginst4383 (R1207_U494, R1207_U79, U3070);
  nand ginst4384 (R1207_U495, R1207_U493, R1207_U494);
  nand ginst4385 (R1207_U496, R1207_U93, U3496);
  nand ginst4386 (R1207_U497, R1207_U80, U3071);
  nand ginst4387 (R1207_U498, R1207_U107, R1207_U330);
  nand ginst4388 (R1207_U499, R1207_U199, R1207_U322);
  not ginst4389 (R1207_U50, U3057);
  nand ginst4390 (R1207_U500, R1207_U94, U3494);
  nand ginst4391 (R1207_U501, R1207_U81, U3076);
  nand ginst4392 (R1207_U502, R1207_U201, R1207_U331);
  nand ginst4393 (R1207_U503, R1207_U200, R1207_U379);
  nand ginst4394 (R1207_U504, R1207_U82, U3492);
  nand ginst4395 (R1207_U505, R1207_U83, U3077);
  not ginst4396 (R1207_U506, R1207_U169);
  nand ginst4397 (R1207_U507, R1207_U377, R1207_U506);
  nand ginst4398 (R1207_U508, R1207_U169, R1207_U202);
  nand ginst4399 (R1207_U509, R1207_U90, U3490);
  nand ginst4400 (R1207_U51, R1207_U38, U3057);
  nand ginst4401 (R1207_U510, R1207_U84, U3069);
  not ginst4402 (R1207_U511, R1207_U170);
  nand ginst4403 (R1207_U512, R1207_U375, R1207_U511);
  nand ginst4404 (R1207_U513, R1207_U170, R1207_U203);
  nand ginst4405 (R1207_U514, R1207_U85, U3488);
  nand ginst4406 (R1207_U515, R1207_U87, U3060);
  nand ginst4407 (R1207_U516, R1207_U514, R1207_U515);
  nand ginst4408 (R1207_U517, R1207_U86, U3486);
  nand ginst4409 (R1207_U518, R1207_U88, U3059);
  nand ginst4410 (R1207_U519, R1207_U108, R1207_U339);
  nand ginst4411 (R1207_U52, R1207_U233, R1207_U235);
  nand ginst4412 (R1207_U520, R1207_U204, R1207_U373);
  not ginst4413 (R1207_U53, U3484);
  not ginst4414 (R1207_U54, U3080);
  nand ginst4415 (R1207_U55, R1207_U236, R1207_U52);
  nand ginst4416 (R1207_U56, R1207_U251, R1207_U51);
  nand ginst4417 (R1207_U57, R1207_U207, R1207_U223, R1207_U341);
  not ginst4418 (R1207_U58, U4031);
  not ginst4419 (R1207_U59, U4030);
  and ginst4420 (R1207_U6, R1207_U230, R1207_U231);
  not ginst4421 (R1207_U60, U3055);
  not ginst4422 (R1207_U61, U4032);
  not ginst4423 (R1207_U62, U3062);
  not ginst4424 (R1207_U63, U4033);
  not ginst4425 (R1207_U64, U3063);
  not ginst4426 (R1207_U65, U3058);
  not ginst4427 (R1207_U66, U3072);
  not ginst4428 (R1207_U67, U4034);
  not ginst4429 (R1207_U68, U4035);
  nand ginst4430 (R1207_U69, R1207_U70, U3072);
  and ginst4431 (R1207_U7, R1207_U211, R1207_U264);
  not ginst4432 (R1207_U70, U4036);
  not ginst4433 (R1207_U71, U3073);
  not ginst4434 (R1207_U72, U3078);
  not ginst4435 (R1207_U73, U4037);
  nand ginst4436 (R1207_U74, R1207_U75, U3078);
  not ginst4437 (R1207_U75, U3504);
  not ginst4438 (R1207_U76, U3079);
  not ginst4439 (R1207_U77, U3066);
  not ginst4440 (R1207_U78, U3500);
  not ginst4441 (R1207_U79, U3498);
  and ginst4442 (R1207_U8, R1207_U265, R1207_U266);
  not ginst4443 (R1207_U80, U3496);
  not ginst4444 (R1207_U81, U3494);
  not ginst4445 (R1207_U82, U3077);
  not ginst4446 (R1207_U83, U3492);
  not ginst4447 (R1207_U84, U3490);
  not ginst4448 (R1207_U85, U3060);
  not ginst4449 (R1207_U86, U3059);
  not ginst4450 (R1207_U87, U3488);
  not ginst4451 (R1207_U88, U3486);
  nand ginst4452 (R1207_U89, R1207_U53, U3080);
  and ginst4453 (R1207_U9, R1207_U212, R1207_U275);
  not ginst4454 (R1207_U90, U3069);
  nand ginst4455 (R1207_U91, R1207_U271, R1207_U347);
  not ginst4456 (R1207_U92, U3070);
  not ginst4457 (R1207_U93, U3071);
  not ginst4458 (R1207_U94, U3076);
  nand ginst4459 (R1207_U95, R1207_U81, U3076);
  nand ginst4460 (R1207_U96, R1207_U279, R1207_U281);
  not ginst4461 (R1207_U97, U3502);
  not ginst4462 (R1207_U98, U3054);
  nand ginst4463 (R1207_U99, R1207_U58, U3054);
  and ginst4464 (R1222_U10, R1222_U267, R1222_U268);
  nand ginst4465 (R1222_U100, R1222_U314, R1222_U59);
  nand ginst4466 (R1222_U101, R1222_U259, R1222_U369, R1222_U370);
  nand ginst4467 (R1222_U102, R1222_U333, R1222_U76);
  nand ginst4468 (R1222_U103, R1222_U471, R1222_U472);
  nand ginst4469 (R1222_U104, R1222_U518, R1222_U519);
  nand ginst4470 (R1222_U105, R1222_U389, R1222_U390);
  nand ginst4471 (R1222_U106, R1222_U394, R1222_U395);
  nand ginst4472 (R1222_U107, R1222_U401, R1222_U402);
  nand ginst4473 (R1222_U108, R1222_U408, R1222_U409);
  nand ginst4474 (R1222_U109, R1222_U413, R1222_U414);
  and ginst4475 (R1222_U11, R1222_U10, R1222_U269);
  nand ginst4476 (R1222_U110, R1222_U422, R1222_U423);
  nand ginst4477 (R1222_U111, R1222_U429, R1222_U430);
  nand ginst4478 (R1222_U112, R1222_U436, R1222_U437);
  nand ginst4479 (R1222_U113, R1222_U443, R1222_U444);
  nand ginst4480 (R1222_U114, R1222_U448, R1222_U449);
  nand ginst4481 (R1222_U115, R1222_U455, R1222_U456);
  nand ginst4482 (R1222_U116, R1222_U462, R1222_U463);
  nand ginst4483 (R1222_U117, R1222_U476, R1222_U477);
  nand ginst4484 (R1222_U118, R1222_U481, R1222_U482);
  nand ginst4485 (R1222_U119, R1222_U488, R1222_U489);
  and ginst4486 (R1222_U12, R1222_U289, R1222_U290);
  nand ginst4487 (R1222_U120, R1222_U495, R1222_U496);
  nand ginst4488 (R1222_U121, R1222_U502, R1222_U503);
  nand ginst4489 (R1222_U122, R1222_U509, R1222_U510);
  nand ginst4490 (R1222_U123, R1222_U514, R1222_U515);
  and ginst4491 (R1222_U124, R1222_U125, R1222_U191);
  and ginst4492 (R1222_U125, U3065, U3470);
  and ginst4493 (R1222_U126, U3061, U3472);
  and ginst4494 (R1222_U127, U3074, U3464);
  and ginst4495 (R1222_U128, R1222_U197, R1222_U198, R1222_U200);
  and ginst4496 (R1222_U129, R1222_U201, R1222_U361, R1222_U362);
  and ginst4497 (R1222_U13, R1222_U209, R1222_U7);
  and ginst4498 (R1222_U130, R1222_U29, R1222_U396, R1222_U397);
  and ginst4499 (R1222_U131, R1222_U214, R1222_U6);
  and ginst4500 (R1222_U132, R1222_U220, R1222_U222);
  and ginst4501 (R1222_U133, R1222_U38, R1222_U403, R1222_U404);
  and ginst4502 (R1222_U134, R1222_U228, R1222_U4);
  and ginst4503 (R1222_U135, R1222_U192, R1222_U236);
  and ginst4504 (R1222_U136, R1222_U182, R1222_U241);
  and ginst4505 (R1222_U137, R1222_U13, R1222_U6);
  and ginst4506 (R1222_U138, R1222_U244, R1222_U365);
  and ginst4507 (R1222_U139, R1222_U16, R1222_U258);
  and ginst4508 (R1222_U14, R1222_U250, R1222_U8);
  and ginst4509 (R1222_U140, R1222_U183, R1222_U248);
  and ginst4510 (R1222_U141, R1222_U15, R1222_U9);
  and ginst4511 (R1222_U142, R1222_U280, R1222_U371);
  and ginst4512 (R1222_U143, R1222_U12, R1222_U294);
  and ginst4513 (R1222_U144, R1222_U184, R1222_U292);
  and ginst4514 (R1222_U145, R1222_U184, R1222_U438, R1222_U439);
  and ginst4515 (R1222_U146, R1222_U12, R1222_U311);
  and ginst4516 (R1222_U147, R1222_U171, R1222_U274);
  and ginst4517 (R1222_U148, R1222_U469, R1222_U470, R1222_U55);
  and ginst4518 (R1222_U149, R1222_U10, R1222_U324);
  and ginst4519 (R1222_U15, R1222_U11, R1222_U278);
  and ginst4520 (R1222_U150, R1222_U483, R1222_U484, R1222_U65);
  and ginst4521 (R1222_U151, R1222_U330, R1222_U9);
  and ginst4522 (R1222_U152, R1222_U183, R1222_U504, R1222_U505);
  and ginst4523 (R1222_U153, R1222_U339, R1222_U8);
  and ginst4524 (R1222_U154, R1222_U182, R1222_U516, R1222_U517);
  and ginst4525 (R1222_U155, R1222_U346, R1222_U7);
  nand ginst4526 (R1222_U156, R1222_U363, R1222_U373);
  nand ginst4527 (R1222_U157, R1222_U219, R1222_U231);
  not ginst4528 (R1222_U158, U3052);
  not ginst4529 (R1222_U159, U4040);
  and ginst4530 (R1222_U16, R1222_U14, R1222_U255);
  and ginst4531 (R1222_U160, R1222_U417, R1222_U418);
  nand ginst4532 (R1222_U161, R1222_U180, R1222_U303, R1222_U360);
  and ginst4533 (R1222_U162, R1222_U424, R1222_U425);
  nand ginst4534 (R1222_U163, R1222_U300, R1222_U301);
  and ginst4535 (R1222_U164, R1222_U431, R1222_U432);
  nand ginst4536 (R1222_U165, R1222_U296, R1222_U297);
  nand ginst4537 (R1222_U166, R1222_U286, R1222_U287);
  and ginst4538 (R1222_U167, R1222_U450, R1222_U451);
  nand ginst4539 (R1222_U168, R1222_U282, R1222_U283);
  and ginst4540 (R1222_U169, R1222_U457, R1222_U458);
  and ginst4541 (R1222_U17, R1222_U344, R1222_U347);
  nand ginst4542 (R1222_U170, R1222_U142, R1222_U384);
  and ginst4543 (R1222_U171, R1222_U464, R1222_U465);
  nand ginst4544 (R1222_U172, U3074, U3464);
  nand ginst4545 (R1222_U173, R1222_U326, R1222_U40);
  nand ginst4546 (R1222_U174, R1222_U364, R1222_U380);
  and ginst4547 (R1222_U175, R1222_U490, R1222_U491);
  nand ginst4548 (R1222_U176, R1222_U366, R1222_U81);
  and ginst4549 (R1222_U177, R1222_U497, R1222_U498);
  nand ginst4550 (R1222_U178, R1222_U252, R1222_U253);
  nand ginst4551 (R1222_U179, R1222_U138, R1222_U377);
  and ginst4552 (R1222_U18, R1222_U337, R1222_U340);
  nand ginst4553 (R1222_U180, R1222_U163, U3051);
  not ginst4554 (R1222_U181, R1222_U38);
  nand ginst4555 (R1222_U182, U3080, U3484);
  nand ginst4556 (R1222_U183, U3069, U3490);
  nand ginst4557 (R1222_U184, U3055, U4032);
  not ginst4558 (R1222_U185, R1222_U76);
  not ginst4559 (R1222_U186, R1222_U59);
  not ginst4560 (R1222_U187, R1222_U90);
  not ginst4561 (R1222_U188, R1222_U69);
  or ginst4562 (R1222_U189, U3064, U3476);
  and ginst4563 (R1222_U19, R1222_U331, R1222_U383);
  or ginst4564 (R1222_U190, U3057, U3474);
  or ginst4565 (R1222_U191, U3061, U3472);
  or ginst4566 (R1222_U192, U3065, U3470);
  not ginst4567 (R1222_U193, R1222_U172);
  or ginst4568 (R1222_U194, U3075, U3468);
  not ginst4569 (R1222_U195, R1222_U43);
  not ginst4570 (R1222_U196, R1222_U40);
  nand ginst4571 (R1222_U197, R1222_U124, R1222_U4);
  nand ginst4572 (R1222_U198, R1222_U126, R1222_U4);
  nand ginst4573 (R1222_U199, R1222_U38, R1222_U39);
  and ginst4574 (R1222_U20, R1222_U322, R1222_U325);
  nand ginst4575 (R1222_U200, R1222_U199, U3064);
  nand ginst4576 (R1222_U201, R1222_U181, U3476);
  not ginst4577 (R1222_U202, R1222_U50);
  or ginst4578 (R1222_U203, U3067, U3480);
  or ginst4579 (R1222_U204, U3068, U3478);
  not ginst4580 (R1222_U205, R1222_U29);
  nand ginst4581 (R1222_U206, R1222_U29, R1222_U30);
  nand ginst4582 (R1222_U207, R1222_U206, U3067);
  nand ginst4583 (R1222_U208, R1222_U205, U3480);
  or ginst4584 (R1222_U209, U3081, U3482);
  and ginst4585 (R1222_U21, R1222_U317, R1222_U319);
  nand ginst4586 (R1222_U210, R1222_U156, R1222_U209);
  not ginst4587 (R1222_U211, R1222_U49);
  or ginst4588 (R1222_U212, U3080, U3484);
  or ginst4589 (R1222_U213, U3068, U3478);
  nand ginst4590 (R1222_U214, U3067, U3480);
  nand ginst4591 (R1222_U215, R1222_U131, R1222_U372);
  or ginst4592 (R1222_U216, U3068, U3478);
  nand ginst4593 (R1222_U217, R1222_U192, R1222_U196);
  nand ginst4594 (R1222_U218, U3065, U3470);
  not ginst4595 (R1222_U219, R1222_U52);
  and ginst4596 (R1222_U22, R1222_U309, R1222_U312);
  nand ginst4597 (R1222_U220, R1222_U195, R1222_U5);
  nand ginst4598 (R1222_U221, R1222_U191, R1222_U52);
  nand ginst4599 (R1222_U222, U3061, U3472);
  not ginst4600 (R1222_U223, R1222_U51);
  or ginst4601 (R1222_U224, U3057, U3474);
  nand ginst4602 (R1222_U225, R1222_U224, R1222_U51);
  nand ginst4603 (R1222_U226, R1222_U133, R1222_U225);
  nand ginst4604 (R1222_U227, R1222_U223, R1222_U38);
  nand ginst4605 (R1222_U228, U3064, U3476);
  nand ginst4606 (R1222_U229, R1222_U134, R1222_U227);
  and ginst4607 (R1222_U23, R1222_U234, R1222_U237);
  or ginst4608 (R1222_U230, U3057, U3474);
  nand ginst4609 (R1222_U231, R1222_U192, R1222_U195);
  not ginst4610 (R1222_U232, R1222_U157);
  nand ginst4611 (R1222_U233, U3061, U3472);
  nand ginst4612 (R1222_U234, R1222_U40, R1222_U415, R1222_U416, R1222_U43);
  nand ginst4613 (R1222_U235, R1222_U40, R1222_U43);
  nand ginst4614 (R1222_U236, U3065, U3470);
  nand ginst4615 (R1222_U237, R1222_U135, R1222_U235);
  or ginst4616 (R1222_U238, U3080, U3484);
  or ginst4617 (R1222_U239, U3059, U3486);
  and ginst4618 (R1222_U24, R1222_U226, R1222_U229);
  nand ginst4619 (R1222_U240, R1222_U188, R1222_U7);
  nand ginst4620 (R1222_U241, U3059, U3486);
  nand ginst4621 (R1222_U242, R1222_U136, R1222_U240);
  or ginst4622 (R1222_U243, U3059, U3486);
  nand ginst4623 (R1222_U244, R1222_U242, R1222_U243);
  or ginst4624 (R1222_U245, U3077, U3492);
  or ginst4625 (R1222_U246, U3069, U3490);
  nand ginst4626 (R1222_U247, R1222_U185, R1222_U8);
  nand ginst4627 (R1222_U248, U3077, U3492);
  nand ginst4628 (R1222_U249, R1222_U140, R1222_U247);
  and ginst4629 (R1222_U25, R1222_U215, R1222_U376);
  or ginst4630 (R1222_U250, U3060, U3488);
  or ginst4631 (R1222_U251, U3077, U3492);
  nand ginst4632 (R1222_U252, R1222_U14, R1222_U179);
  nand ginst4633 (R1222_U253, R1222_U249, R1222_U251);
  not ginst4634 (R1222_U254, R1222_U178);
  or ginst4635 (R1222_U255, U3076, U3494);
  nand ginst4636 (R1222_U256, U3076, U3494);
  not ginst4637 (R1222_U257, R1222_U176);
  or ginst4638 (R1222_U258, U3071, U3496);
  nand ginst4639 (R1222_U259, U3071, U3496);
  not ginst4640 (R1222_U26, U3478);
  not ginst4641 (R1222_U260, R1222_U101);
  or ginst4642 (R1222_U261, U3066, U3500);
  or ginst4643 (R1222_U262, U3070, U3498);
  not ginst4644 (R1222_U263, R1222_U65);
  nand ginst4645 (R1222_U264, R1222_U65, R1222_U66);
  nand ginst4646 (R1222_U265, R1222_U264, U3066);
  nand ginst4647 (R1222_U266, R1222_U263, U3500);
  or ginst4648 (R1222_U267, U3073, U4037);
  or ginst4649 (R1222_U268, U3078, U3504);
  or ginst4650 (R1222_U269, U3072, U4036);
  not ginst4651 (R1222_U27, U3068);
  not ginst4652 (R1222_U270, R1222_U55);
  nand ginst4653 (R1222_U271, R1222_U270, U4037);
  nand ginst4654 (R1222_U272, R1222_U271, R1222_U99);
  nand ginst4655 (R1222_U273, R1222_U55, R1222_U56);
  nand ginst4656 (R1222_U274, R1222_U272, R1222_U273);
  nand ginst4657 (R1222_U275, R1222_U11, R1222_U186);
  nand ginst4658 (R1222_U276, U3072, U4036);
  nand ginst4659 (R1222_U277, R1222_U274, R1222_U275, R1222_U276);
  or ginst4660 (R1222_U278, U3079, U3502);
  or ginst4661 (R1222_U279, U3072, U4036);
  not ginst4662 (R1222_U28, U3067);
  nand ginst4663 (R1222_U280, R1222_U277, R1222_U279);
  or ginst4664 (R1222_U281, U3058, U4035);
  nand ginst4665 (R1222_U282, R1222_U170, R1222_U281);
  nand ginst4666 (R1222_U283, U3058, U4035);
  not ginst4667 (R1222_U284, R1222_U168);
  or ginst4668 (R1222_U285, U3063, U4034);
  nand ginst4669 (R1222_U286, R1222_U168, R1222_U285);
  nand ginst4670 (R1222_U287, U3063, U4034);
  not ginst4671 (R1222_U288, R1222_U166);
  or ginst4672 (R1222_U289, U3054, U4031);
  nand ginst4673 (R1222_U29, U3068, U3478);
  or ginst4674 (R1222_U290, U3055, U4032);
  nand ginst4675 (R1222_U291, R1222_U12, R1222_U187);
  nand ginst4676 (R1222_U292, U3054, U4031);
  nand ginst4677 (R1222_U293, R1222_U144, R1222_U291);
  or ginst4678 (R1222_U294, U3062, U4033);
  or ginst4679 (R1222_U295, U3054, U4031);
  nand ginst4680 (R1222_U296, R1222_U143, R1222_U166);
  nand ginst4681 (R1222_U297, R1222_U293, R1222_U295);
  not ginst4682 (R1222_U298, R1222_U165);
  or ginst4683 (R1222_U299, U3050, U4030);
  not ginst4684 (R1222_U30, U3480);
  nand ginst4685 (R1222_U300, R1222_U165, R1222_U299);
  nand ginst4686 (R1222_U301, U3050, U4030);
  not ginst4687 (R1222_U302, R1222_U163);
  nand ginst4688 (R1222_U303, R1222_U163, U4029);
  not ginst4689 (R1222_U304, R1222_U161);
  nand ginst4690 (R1222_U305, R1222_U166, R1222_U294);
  not ginst4691 (R1222_U306, R1222_U97);
  or ginst4692 (R1222_U307, U3055, U4032);
  nand ginst4693 (R1222_U308, R1222_U307, R1222_U97);
  nand ginst4694 (R1222_U309, R1222_U145, R1222_U308);
  not ginst4695 (R1222_U31, U3470);
  nand ginst4696 (R1222_U310, R1222_U184, R1222_U306);
  nand ginst4697 (R1222_U311, U3054, U4031);
  nand ginst4698 (R1222_U312, R1222_U146, R1222_U310);
  or ginst4699 (R1222_U313, U3055, U4032);
  nand ginst4700 (R1222_U314, R1222_U174, R1222_U278);
  not ginst4701 (R1222_U315, R1222_U100);
  nand ginst4702 (R1222_U316, R1222_U10, R1222_U100);
  nand ginst4703 (R1222_U317, R1222_U147, R1222_U316);
  nand ginst4704 (R1222_U318, R1222_U274, R1222_U316);
  nand ginst4705 (R1222_U319, R1222_U318, R1222_U468);
  not ginst4706 (R1222_U32, U3065);
  or ginst4707 (R1222_U320, U3078, U3504);
  nand ginst4708 (R1222_U321, R1222_U100, R1222_U320);
  nand ginst4709 (R1222_U322, R1222_U148, R1222_U321);
  nand ginst4710 (R1222_U323, R1222_U315, R1222_U55);
  nand ginst4711 (R1222_U324, U3073, U4037);
  nand ginst4712 (R1222_U325, R1222_U149, R1222_U323);
  or ginst4713 (R1222_U326, U3075, U3468);
  not ginst4714 (R1222_U327, R1222_U173);
  or ginst4715 (R1222_U328, U3078, U3504);
  or ginst4716 (R1222_U329, U3070, U3498);
  not ginst4717 (R1222_U33, U3472);
  nand ginst4718 (R1222_U330, U3066, U3500);
  nand ginst4719 (R1222_U331, R1222_U151, R1222_U379);
  or ginst4720 (R1222_U332, U3070, U3498);
  nand ginst4721 (R1222_U333, R1222_U179, R1222_U250);
  not ginst4722 (R1222_U334, R1222_U102);
  or ginst4723 (R1222_U335, U3069, U3490);
  nand ginst4724 (R1222_U336, R1222_U102, R1222_U335);
  nand ginst4725 (R1222_U337, R1222_U152, R1222_U336);
  nand ginst4726 (R1222_U338, R1222_U183, R1222_U334);
  nand ginst4727 (R1222_U339, U3077, U3492);
  not ginst4728 (R1222_U34, U3061);
  nand ginst4729 (R1222_U340, R1222_U153, R1222_U338);
  or ginst4730 (R1222_U341, U3069, U3490);
  or ginst4731 (R1222_U342, U3080, U3484);
  nand ginst4732 (R1222_U343, R1222_U342, R1222_U49);
  nand ginst4733 (R1222_U344, R1222_U154, R1222_U343);
  nand ginst4734 (R1222_U345, R1222_U182, R1222_U211);
  nand ginst4735 (R1222_U346, U3059, U3486);
  nand ginst4736 (R1222_U347, R1222_U155, R1222_U345);
  nand ginst4737 (R1222_U348, R1222_U182, R1222_U212);
  nand ginst4738 (R1222_U349, R1222_U209, R1222_U69);
  not ginst4739 (R1222_U35, U3474);
  nand ginst4740 (R1222_U350, R1222_U216, R1222_U29);
  nand ginst4741 (R1222_U351, R1222_U230, R1222_U38);
  nand ginst4742 (R1222_U352, R1222_U191, R1222_U233);
  nand ginst4743 (R1222_U353, R1222_U184, R1222_U313);
  nand ginst4744 (R1222_U354, R1222_U294, R1222_U90);
  nand ginst4745 (R1222_U355, R1222_U328, R1222_U55);
  nand ginst4746 (R1222_U356, R1222_U278, R1222_U59);
  nand ginst4747 (R1222_U357, R1222_U332, R1222_U65);
  nand ginst4748 (R1222_U358, R1222_U183, R1222_U341);
  nand ginst4749 (R1222_U359, R1222_U250, R1222_U76);
  not ginst4750 (R1222_U36, U3057);
  nand ginst4751 (R1222_U360, U3051, U4029);
  nand ginst4752 (R1222_U361, R1222_U196, R1222_U4, R1222_U5);
  nand ginst4753 (R1222_U362, R1222_U195, R1222_U4, R1222_U5);
  not ginst4754 (R1222_U363, R1222_U44);
  not ginst4755 (R1222_U364, R1222_U98);
  nand ginst4756 (R1222_U365, R1222_U13, R1222_U44);
  nand ginst4757 (R1222_U366, R1222_U16, R1222_U179);
  nand ginst4758 (R1222_U367, R1222_U253, R1222_U256);
  not ginst4759 (R1222_U368, R1222_U81);
  nand ginst4760 (R1222_U369, R1222_U139, R1222_U179);
  not ginst4761 (R1222_U37, U3064);
  nand ginst4762 (R1222_U370, R1222_U258, R1222_U368);
  nand ginst4763 (R1222_U371, R1222_U15, R1222_U98);
  nand ginst4764 (R1222_U372, R1222_U202, R1222_U29);
  nand ginst4765 (R1222_U373, R1222_U50, R1222_U6);
  not ginst4766 (R1222_U374, R1222_U156);
  nand ginst4767 (R1222_U375, R1222_U213, R1222_U50);
  nand ginst4768 (R1222_U376, R1222_U130, R1222_U375);
  nand ginst4769 (R1222_U377, R1222_U137, R1222_U50);
  not ginst4770 (R1222_U378, R1222_U179);
  nand ginst4771 (R1222_U379, R1222_U260, R1222_U65);
  nand ginst4772 (R1222_U38, U3057, U3474);
  nand ginst4773 (R1222_U380, R1222_U101, R1222_U9);
  not ginst4774 (R1222_U381, R1222_U174);
  nand ginst4775 (R1222_U382, R1222_U101, R1222_U329);
  nand ginst4776 (R1222_U383, R1222_U150, R1222_U382);
  nand ginst4777 (R1222_U384, R1222_U101, R1222_U141);
  not ginst4778 (R1222_U385, R1222_U170);
  nand ginst4779 (R1222_U386, R1222_U48, U3080);
  nand ginst4780 (R1222_U387, R1222_U47, U3484);
  nand ginst4781 (R1222_U388, R1222_U386, R1222_U387);
  nand ginst4782 (R1222_U389, R1222_U348, R1222_U49);
  not ginst4783 (R1222_U39, U3476);
  nand ginst4784 (R1222_U390, R1222_U211, R1222_U388);
  nand ginst4785 (R1222_U391, R1222_U45, U3081);
  nand ginst4786 (R1222_U392, R1222_U46, U3482);
  nand ginst4787 (R1222_U393, R1222_U391, R1222_U392);
  nand ginst4788 (R1222_U394, R1222_U156, R1222_U349);
  nand ginst4789 (R1222_U395, R1222_U374, R1222_U393);
  nand ginst4790 (R1222_U396, R1222_U30, U3067);
  nand ginst4791 (R1222_U397, R1222_U28, U3480);
  nand ginst4792 (R1222_U398, R1222_U26, U3068);
  nand ginst4793 (R1222_U399, R1222_U27, U3478);
  and ginst4794 (R1222_U4, R1222_U189, R1222_U190);
  nand ginst4795 (R1222_U40, U3075, U3468);
  nand ginst4796 (R1222_U400, R1222_U398, R1222_U399);
  nand ginst4797 (R1222_U401, R1222_U350, R1222_U50);
  nand ginst4798 (R1222_U402, R1222_U202, R1222_U400);
  nand ginst4799 (R1222_U403, R1222_U39, U3064);
  nand ginst4800 (R1222_U404, R1222_U37, U3476);
  nand ginst4801 (R1222_U405, R1222_U35, U3057);
  nand ginst4802 (R1222_U406, R1222_U36, U3474);
  nand ginst4803 (R1222_U407, R1222_U405, R1222_U406);
  nand ginst4804 (R1222_U408, R1222_U351, R1222_U51);
  nand ginst4805 (R1222_U409, R1222_U223, R1222_U407);
  not ginst4806 (R1222_U41, U3464);
  nand ginst4807 (R1222_U410, R1222_U33, U3061);
  nand ginst4808 (R1222_U411, R1222_U34, U3472);
  nand ginst4809 (R1222_U412, R1222_U410, R1222_U411);
  nand ginst4810 (R1222_U413, R1222_U157, R1222_U352);
  nand ginst4811 (R1222_U414, R1222_U232, R1222_U412);
  nand ginst4812 (R1222_U415, R1222_U31, U3065);
  nand ginst4813 (R1222_U416, R1222_U32, U3470);
  nand ginst4814 (R1222_U417, R1222_U159, U3052);
  nand ginst4815 (R1222_U418, R1222_U158, U4040);
  nand ginst4816 (R1222_U419, R1222_U159, U3052);
  not ginst4817 (R1222_U42, U3074);
  nand ginst4818 (R1222_U420, R1222_U158, U4040);
  nand ginst4819 (R1222_U421, R1222_U419, R1222_U420);
  nand ginst4820 (R1222_U422, R1222_U160, R1222_U161);
  nand ginst4821 (R1222_U423, R1222_U304, R1222_U421);
  nand ginst4822 (R1222_U424, R1222_U96, U3051);
  nand ginst4823 (R1222_U425, R1222_U95, U4029);
  nand ginst4824 (R1222_U426, R1222_U96, U3051);
  nand ginst4825 (R1222_U427, R1222_U95, U4029);
  nand ginst4826 (R1222_U428, R1222_U426, R1222_U427);
  nand ginst4827 (R1222_U429, R1222_U162, R1222_U163);
  nand ginst4828 (R1222_U43, R1222_U127, R1222_U194);
  nand ginst4829 (R1222_U430, R1222_U302, R1222_U428);
  nand ginst4830 (R1222_U431, R1222_U93, U3050);
  nand ginst4831 (R1222_U432, R1222_U94, U4030);
  nand ginst4832 (R1222_U433, R1222_U93, U3050);
  nand ginst4833 (R1222_U434, R1222_U94, U4030);
  nand ginst4834 (R1222_U435, R1222_U433, R1222_U434);
  nand ginst4835 (R1222_U436, R1222_U164, R1222_U165);
  nand ginst4836 (R1222_U437, R1222_U298, R1222_U435);
  nand ginst4837 (R1222_U438, R1222_U91, U3054);
  nand ginst4838 (R1222_U439, R1222_U92, U4031);
  nand ginst4839 (R1222_U44, R1222_U207, R1222_U208);
  nand ginst4840 (R1222_U440, R1222_U86, U3055);
  nand ginst4841 (R1222_U441, R1222_U87, U4032);
  nand ginst4842 (R1222_U442, R1222_U440, R1222_U441);
  nand ginst4843 (R1222_U443, R1222_U353, R1222_U97);
  nand ginst4844 (R1222_U444, R1222_U306, R1222_U442);
  nand ginst4845 (R1222_U445, R1222_U88, U3062);
  nand ginst4846 (R1222_U446, R1222_U89, U4033);
  nand ginst4847 (R1222_U447, R1222_U445, R1222_U446);
  nand ginst4848 (R1222_U448, R1222_U166, R1222_U354);
  nand ginst4849 (R1222_U449, R1222_U288, R1222_U447);
  not ginst4850 (R1222_U45, U3482);
  nand ginst4851 (R1222_U450, R1222_U84, U3063);
  nand ginst4852 (R1222_U451, R1222_U85, U4034);
  nand ginst4853 (R1222_U452, R1222_U84, U3063);
  nand ginst4854 (R1222_U453, R1222_U85, U4034);
  nand ginst4855 (R1222_U454, R1222_U452, R1222_U453);
  nand ginst4856 (R1222_U455, R1222_U167, R1222_U168);
  nand ginst4857 (R1222_U456, R1222_U284, R1222_U454);
  nand ginst4858 (R1222_U457, R1222_U82, U3058);
  nand ginst4859 (R1222_U458, R1222_U83, U4035);
  nand ginst4860 (R1222_U459, R1222_U82, U3058);
  not ginst4861 (R1222_U46, U3081);
  nand ginst4862 (R1222_U460, R1222_U83, U4035);
  nand ginst4863 (R1222_U461, R1222_U459, R1222_U460);
  nand ginst4864 (R1222_U462, R1222_U169, R1222_U170);
  nand ginst4865 (R1222_U463, R1222_U385, R1222_U461);
  nand ginst4866 (R1222_U464, R1222_U60, U3072);
  nand ginst4867 (R1222_U465, R1222_U61, U4036);
  nand ginst4868 (R1222_U466, R1222_U60, U3072);
  nand ginst4869 (R1222_U467, R1222_U61, U4036);
  nand ginst4870 (R1222_U468, R1222_U466, R1222_U467);
  nand ginst4871 (R1222_U469, R1222_U56, U3073);
  not ginst4872 (R1222_U47, U3080);
  nand ginst4873 (R1222_U470, R1222_U99, U4037);
  nand ginst4874 (R1222_U471, R1222_U173, R1222_U193);
  nand ginst4875 (R1222_U472, R1222_U172, R1222_U327);
  nand ginst4876 (R1222_U473, R1222_U53, U3078);
  nand ginst4877 (R1222_U474, R1222_U54, U3504);
  nand ginst4878 (R1222_U475, R1222_U473, R1222_U474);
  nand ginst4879 (R1222_U476, R1222_U100, R1222_U355);
  nand ginst4880 (R1222_U477, R1222_U315, R1222_U475);
  nand ginst4881 (R1222_U478, R1222_U57, U3079);
  nand ginst4882 (R1222_U479, R1222_U58, U3502);
  not ginst4883 (R1222_U48, U3484);
  nand ginst4884 (R1222_U480, R1222_U478, R1222_U479);
  nand ginst4885 (R1222_U481, R1222_U174, R1222_U356);
  nand ginst4886 (R1222_U482, R1222_U381, R1222_U480);
  nand ginst4887 (R1222_U483, R1222_U66, U3066);
  nand ginst4888 (R1222_U484, R1222_U64, U3500);
  nand ginst4889 (R1222_U485, R1222_U62, U3070);
  nand ginst4890 (R1222_U486, R1222_U63, U3498);
  nand ginst4891 (R1222_U487, R1222_U485, R1222_U486);
  nand ginst4892 (R1222_U488, R1222_U101, R1222_U357);
  nand ginst4893 (R1222_U489, R1222_U260, R1222_U487);
  nand ginst4894 (R1222_U49, R1222_U210, R1222_U69);
  nand ginst4895 (R1222_U490, R1222_U67, U3071);
  nand ginst4896 (R1222_U491, R1222_U68, U3496);
  nand ginst4897 (R1222_U492, R1222_U67, U3071);
  nand ginst4898 (R1222_U493, R1222_U68, U3496);
  nand ginst4899 (R1222_U494, R1222_U492, R1222_U493);
  nand ginst4900 (R1222_U495, R1222_U175, R1222_U176);
  nand ginst4901 (R1222_U496, R1222_U257, R1222_U494);
  nand ginst4902 (R1222_U497, R1222_U79, U3076);
  nand ginst4903 (R1222_U498, R1222_U80, U3494);
  nand ginst4904 (R1222_U499, R1222_U79, U3076);
  and ginst4905 (R1222_U5, R1222_U191, R1222_U192);
  nand ginst4906 (R1222_U50, R1222_U128, R1222_U129);
  nand ginst4907 (R1222_U500, R1222_U80, U3494);
  nand ginst4908 (R1222_U501, R1222_U499, R1222_U500);
  nand ginst4909 (R1222_U502, R1222_U177, R1222_U178);
  nand ginst4910 (R1222_U503, R1222_U254, R1222_U501);
  nand ginst4911 (R1222_U504, R1222_U77, U3077);
  nand ginst4912 (R1222_U505, R1222_U78, U3492);
  nand ginst4913 (R1222_U506, R1222_U72, U3069);
  nand ginst4914 (R1222_U507, R1222_U73, U3490);
  nand ginst4915 (R1222_U508, R1222_U506, R1222_U507);
  nand ginst4916 (R1222_U509, R1222_U102, R1222_U358);
  nand ginst4917 (R1222_U51, R1222_U132, R1222_U221);
  nand ginst4918 (R1222_U510, R1222_U334, R1222_U508);
  nand ginst4919 (R1222_U511, R1222_U74, U3060);
  nand ginst4920 (R1222_U512, R1222_U75, U3488);
  nand ginst4921 (R1222_U513, R1222_U511, R1222_U512);
  nand ginst4922 (R1222_U514, R1222_U179, R1222_U359);
  nand ginst4923 (R1222_U515, R1222_U378, R1222_U513);
  nand ginst4924 (R1222_U516, R1222_U70, U3059);
  nand ginst4925 (R1222_U517, R1222_U71, U3486);
  nand ginst4926 (R1222_U518, R1222_U41, U3074);
  nand ginst4927 (R1222_U519, R1222_U42, U3464);
  nand ginst4928 (R1222_U52, R1222_U217, R1222_U218);
  not ginst4929 (R1222_U53, U3504);
  not ginst4930 (R1222_U54, U3078);
  nand ginst4931 (R1222_U55, U3078, U3504);
  not ginst4932 (R1222_U56, U4037);
  not ginst4933 (R1222_U57, U3502);
  not ginst4934 (R1222_U58, U3079);
  nand ginst4935 (R1222_U59, U3079, U3502);
  and ginst4936 (R1222_U6, R1222_U203, R1222_U204);
  not ginst4937 (R1222_U60, U4036);
  not ginst4938 (R1222_U61, U3072);
  not ginst4939 (R1222_U62, U3498);
  not ginst4940 (R1222_U63, U3070);
  not ginst4941 (R1222_U64, U3066);
  nand ginst4942 (R1222_U65, U3070, U3498);
  not ginst4943 (R1222_U66, U3500);
  not ginst4944 (R1222_U67, U3496);
  not ginst4945 (R1222_U68, U3071);
  nand ginst4946 (R1222_U69, U3081, U3482);
  and ginst4947 (R1222_U7, R1222_U238, R1222_U239);
  not ginst4948 (R1222_U70, U3486);
  not ginst4949 (R1222_U71, U3059);
  not ginst4950 (R1222_U72, U3490);
  not ginst4951 (R1222_U73, U3069);
  not ginst4952 (R1222_U74, U3488);
  not ginst4953 (R1222_U75, U3060);
  nand ginst4954 (R1222_U76, U3060, U3488);
  not ginst4955 (R1222_U77, U3492);
  not ginst4956 (R1222_U78, U3077);
  not ginst4957 (R1222_U79, U3494);
  and ginst4958 (R1222_U8, R1222_U245, R1222_U246);
  not ginst4959 (R1222_U80, U3076);
  nand ginst4960 (R1222_U81, R1222_U255, R1222_U367);
  not ginst4961 (R1222_U82, U4035);
  not ginst4962 (R1222_U83, U3058);
  not ginst4963 (R1222_U84, U4034);
  not ginst4964 (R1222_U85, U3063);
  not ginst4965 (R1222_U86, U4032);
  not ginst4966 (R1222_U87, U3055);
  not ginst4967 (R1222_U88, U4033);
  not ginst4968 (R1222_U89, U3062);
  and ginst4969 (R1222_U9, R1222_U261, R1222_U262);
  nand ginst4970 (R1222_U90, U3062, U4033);
  not ginst4971 (R1222_U91, U4031);
  not ginst4972 (R1222_U92, U3054);
  not ginst4973 (R1222_U93, U4030);
  not ginst4974 (R1222_U94, U3050);
  not ginst4975 (R1222_U95, U3051);
  not ginst4976 (R1222_U96, U4029);
  nand ginst4977 (R1222_U97, R1222_U305, R1222_U90);
  nand ginst4978 (R1222_U98, R1222_U265, R1222_U266);
  not ginst4979 (R1222_U99, U3073);
  and ginst4980 (R1240_U10, R1240_U281, R1240_U282);
  nand ginst4981 (R1240_U100, R1240_U314, R1240_U60);
  nand ginst4982 (R1240_U101, R1240_U294, R1240_U385);
  nand ginst4983 (R1240_U102, R1240_U277, R1240_U278);
  not ginst4984 (R1240_U103, U3073);
  nand ginst4985 (R1240_U104, R1240_U323, R1240_U84);
  nand ginst4986 (R1240_U105, R1240_U271, R1240_U382, R1240_U383);
  nand ginst4987 (R1240_U106, R1240_U345, R1240_U72);
  nand ginst4988 (R1240_U107, R1240_U483, R1240_U484);
  nand ginst4989 (R1240_U108, R1240_U530, R1240_U531);
  nand ginst4990 (R1240_U109, R1240_U401, R1240_U402);
  and ginst4991 (R1240_U11, R1240_U10, R1240_U283);
  nand ginst4992 (R1240_U110, R1240_U406, R1240_U407);
  nand ginst4993 (R1240_U111, R1240_U413, R1240_U414);
  nand ginst4994 (R1240_U112, R1240_U420, R1240_U421);
  nand ginst4995 (R1240_U113, R1240_U425, R1240_U426);
  nand ginst4996 (R1240_U114, R1240_U434, R1240_U435);
  nand ginst4997 (R1240_U115, R1240_U441, R1240_U442);
  nand ginst4998 (R1240_U116, R1240_U448, R1240_U449);
  nand ginst4999 (R1240_U117, R1240_U455, R1240_U456);
  nand ginst5000 (R1240_U118, R1240_U460, R1240_U461);
  nand ginst5001 (R1240_U119, R1240_U467, R1240_U468);
  and ginst5002 (R1240_U12, R1240_U217, R1240_U7);
  nand ginst5003 (R1240_U120, R1240_U474, R1240_U475);
  nand ginst5004 (R1240_U121, R1240_U488, R1240_U489);
  nand ginst5005 (R1240_U122, R1240_U493, R1240_U494);
  nand ginst5006 (R1240_U123, R1240_U500, R1240_U501);
  nand ginst5007 (R1240_U124, R1240_U507, R1240_U508);
  nand ginst5008 (R1240_U125, R1240_U514, R1240_U515);
  nand ginst5009 (R1240_U126, R1240_U521, R1240_U522);
  nand ginst5010 (R1240_U127, R1240_U526, R1240_U527);
  and ginst5011 (R1240_U128, R1240_U129, R1240_U197);
  and ginst5012 (R1240_U129, U3065, U3470);
  and ginst5013 (R1240_U13, R1240_U262, R1240_U8);
  and ginst5014 (R1240_U130, U3061, U3472);
  and ginst5015 (R1240_U131, U3074, U3464);
  and ginst5016 (R1240_U132, R1240_U203, R1240_U204, R1240_U206);
  and ginst5017 (R1240_U133, R1240_U207, R1240_U373, R1240_U374);
  and ginst5018 (R1240_U134, R1240_U408, R1240_U409, R1240_U43);
  and ginst5019 (R1240_U135, R1240_U225, R1240_U6);
  and ginst5020 (R1240_U136, R1240_U231, R1240_U233);
  and ginst5021 (R1240_U137, R1240_U34, R1240_U415, R1240_U416);
  and ginst5022 (R1240_U138, R1240_U239, R1240_U4);
  and ginst5023 (R1240_U139, R1240_U198, R1240_U247);
  and ginst5024 (R1240_U14, R1240_U11, R1240_U292);
  and ginst5025 (R1240_U140, R1240_U188, R1240_U252);
  and ginst5026 (R1240_U141, R1240_U12, R1240_U6);
  and ginst5027 (R1240_U142, R1240_U255, R1240_U378);
  and ginst5028 (R1240_U143, R1240_U15, R1240_U270);
  and ginst5029 (R1240_U144, R1240_U189, R1240_U260);
  and ginst5030 (R1240_U145, R1240_U16, R1240_U296);
  and ginst5031 (R1240_U146, R1240_U297, R1240_U389);
  and ginst5032 (R1240_U147, R1240_U185, R1240_U309);
  and ginst5033 (R1240_U148, R1240_U310, R1240_U393, R1240_U395);
  and ginst5034 (R1240_U149, R1240_U17, R1240_U185);
  and ginst5035 (R1240_U15, R1240_U13, R1240_U267);
  and ginst5036 (R1240_U150, R1240_U304, R1240_U97);
  and ginst5037 (R1240_U151, R1240_U190, R1240_U450, R1240_U451);
  and ginst5038 (R1240_U152, R1240_U185, R1240_U320);
  and ginst5039 (R1240_U153, R1240_U176, R1240_U288);
  and ginst5040 (R1240_U154, R1240_U481, R1240_U482, R1240_U80);
  and ginst5041 (R1240_U155, R1240_U10, R1240_U333);
  and ginst5042 (R1240_U156, R1240_U495, R1240_U496, R1240_U90);
  and ginst5043 (R1240_U157, R1240_U342, R1240_U9);
  and ginst5044 (R1240_U158, R1240_U189, R1240_U516, R1240_U517);
  and ginst5045 (R1240_U159, R1240_U351, R1240_U8);
  and ginst5046 (R1240_U16, R1240_U14, R1240_U9);
  and ginst5047 (R1240_U160, R1240_U188, R1240_U528, R1240_U529);
  and ginst5048 (R1240_U161, R1240_U358, R1240_U7);
  nand ginst5049 (R1240_U162, R1240_U215, R1240_U375);
  nand ginst5050 (R1240_U163, R1240_U230, R1240_U242);
  not ginst5051 (R1240_U164, U3052);
  not ginst5052 (R1240_U165, U4040);
  and ginst5053 (R1240_U166, R1240_U429, R1240_U430);
  nand ginst5054 (R1240_U167, R1240_U186, R1240_U312, R1240_U372);
  and ginst5055 (R1240_U168, R1240_U436, R1240_U437);
  nand ginst5056 (R1240_U169, R1240_U148, R1240_U394);
  and ginst5057 (R1240_U17, R1240_U299, R1240_U305);
  and ginst5058 (R1240_U170, R1240_U443, R1240_U444);
  nand ginst5059 (R1240_U171, R1240_U150, R1240_U307);
  nand ginst5060 (R1240_U172, R1240_U300, R1240_U301);
  and ginst5061 (R1240_U173, R1240_U462, R1240_U463);
  and ginst5062 (R1240_U174, R1240_U469, R1240_U470);
  nand ginst5063 (R1240_U175, R1240_U384, R1240_U386);
  and ginst5064 (R1240_U176, R1240_U476, R1240_U477);
  nand ginst5065 (R1240_U177, U3074, U3464);
  nand ginst5066 (R1240_U178, R1240_U335, R1240_U36);
  nand ginst5067 (R1240_U179, R1240_U279, R1240_U376);
  and ginst5068 (R1240_U18, R1240_U356, R1240_U359);
  and ginst5069 (R1240_U180, R1240_U502, R1240_U503);
  nand ginst5070 (R1240_U181, R1240_U379, R1240_U77);
  and ginst5071 (R1240_U182, R1240_U509, R1240_U510);
  nand ginst5072 (R1240_U183, R1240_U264, R1240_U265);
  nand ginst5073 (R1240_U184, R1240_U142, R1240_U377);
  nand ginst5074 (R1240_U185, R1240_U390, R1240_U391);
  nand ginst5075 (R1240_U186, R1240_U169, U3051);
  not ginst5076 (R1240_U187, R1240_U34);
  nand ginst5077 (R1240_U188, U3080, U3484);
  nand ginst5078 (R1240_U189, U3069, U3490);
  and ginst5079 (R1240_U19, R1240_U349, R1240_U352);
  nand ginst5080 (R1240_U190, U3055, U4032);
  not ginst5081 (R1240_U191, R1240_U72);
  not ginst5082 (R1240_U192, R1240_U84);
  not ginst5083 (R1240_U193, R1240_U60);
  not ginst5084 (R1240_U194, R1240_U65);
  or ginst5085 (R1240_U195, U3064, U3476);
  or ginst5086 (R1240_U196, U3057, U3474);
  or ginst5087 (R1240_U197, U3061, U3472);
  or ginst5088 (R1240_U198, U3065, U3470);
  not ginst5089 (R1240_U199, R1240_U177);
  and ginst5090 (R1240_U20, R1240_U340, R1240_U343);
  or ginst5091 (R1240_U200, U3075, U3468);
  not ginst5092 (R1240_U201, R1240_U39);
  not ginst5093 (R1240_U202, R1240_U36);
  nand ginst5094 (R1240_U203, R1240_U128, R1240_U4);
  nand ginst5095 (R1240_U204, R1240_U130, R1240_U4);
  nand ginst5096 (R1240_U205, R1240_U34, R1240_U35);
  nand ginst5097 (R1240_U206, R1240_U205, U3064);
  nand ginst5098 (R1240_U207, R1240_U187, U3476);
  not ginst5099 (R1240_U208, R1240_U51);
  or ginst5100 (R1240_U209, U3067, U3480);
  and ginst5101 (R1240_U21, R1240_U331, R1240_U334);
  or ginst5102 (R1240_U210, U3068, U3478);
  not ginst5103 (R1240_U211, R1240_U43);
  nand ginst5104 (R1240_U212, R1240_U43, R1240_U44);
  nand ginst5105 (R1240_U213, R1240_U212, U3067);
  nand ginst5106 (R1240_U214, R1240_U211, U3480);
  nand ginst5107 (R1240_U215, R1240_U51, R1240_U6);
  not ginst5108 (R1240_U216, R1240_U162);
  or ginst5109 (R1240_U217, U3081, U3482);
  nand ginst5110 (R1240_U218, R1240_U162, R1240_U217);
  not ginst5111 (R1240_U219, R1240_U50);
  and ginst5112 (R1240_U22, R1240_U326, R1240_U328);
  or ginst5113 (R1240_U220, U3080, U3484);
  or ginst5114 (R1240_U221, U3068, U3478);
  nand ginst5115 (R1240_U222, R1240_U221, R1240_U51);
  nand ginst5116 (R1240_U223, R1240_U134, R1240_U222);
  nand ginst5117 (R1240_U224, R1240_U208, R1240_U43);
  nand ginst5118 (R1240_U225, U3067, U3480);
  nand ginst5119 (R1240_U226, R1240_U135, R1240_U224);
  or ginst5120 (R1240_U227, U3068, U3478);
  nand ginst5121 (R1240_U228, R1240_U198, R1240_U202);
  nand ginst5122 (R1240_U229, U3065, U3470);
  and ginst5123 (R1240_U23, R1240_U318, R1240_U321);
  not ginst5124 (R1240_U230, R1240_U53);
  nand ginst5125 (R1240_U231, R1240_U201, R1240_U5);
  nand ginst5126 (R1240_U232, R1240_U197, R1240_U53);
  nand ginst5127 (R1240_U233, U3061, U3472);
  not ginst5128 (R1240_U234, R1240_U52);
  or ginst5129 (R1240_U235, U3057, U3474);
  nand ginst5130 (R1240_U236, R1240_U235, R1240_U52);
  nand ginst5131 (R1240_U237, R1240_U137, R1240_U236);
  nand ginst5132 (R1240_U238, R1240_U234, R1240_U34);
  nand ginst5133 (R1240_U239, U3064, U3476);
  and ginst5134 (R1240_U24, R1240_U245, R1240_U248);
  nand ginst5135 (R1240_U240, R1240_U138, R1240_U238);
  or ginst5136 (R1240_U241, U3057, U3474);
  nand ginst5137 (R1240_U242, R1240_U198, R1240_U201);
  not ginst5138 (R1240_U243, R1240_U163);
  nand ginst5139 (R1240_U244, U3061, U3472);
  nand ginst5140 (R1240_U245, R1240_U36, R1240_U39, R1240_U427, R1240_U428);
  nand ginst5141 (R1240_U246, R1240_U36, R1240_U39);
  nand ginst5142 (R1240_U247, U3065, U3470);
  nand ginst5143 (R1240_U248, R1240_U139, R1240_U246);
  or ginst5144 (R1240_U249, U3080, U3484);
  and ginst5145 (R1240_U25, R1240_U237, R1240_U240);
  or ginst5146 (R1240_U250, U3059, U3486);
  nand ginst5147 (R1240_U251, R1240_U194, R1240_U7);
  nand ginst5148 (R1240_U252, U3059, U3486);
  nand ginst5149 (R1240_U253, R1240_U140, R1240_U251);
  or ginst5150 (R1240_U254, U3059, U3486);
  nand ginst5151 (R1240_U255, R1240_U253, R1240_U254);
  not ginst5152 (R1240_U256, R1240_U184);
  or ginst5153 (R1240_U257, U3077, U3492);
  or ginst5154 (R1240_U258, U3069, U3490);
  nand ginst5155 (R1240_U259, R1240_U191, R1240_U8);
  and ginst5156 (R1240_U26, R1240_U223, R1240_U226);
  nand ginst5157 (R1240_U260, U3077, U3492);
  nand ginst5158 (R1240_U261, R1240_U144, R1240_U259);
  or ginst5159 (R1240_U262, U3060, U3488);
  or ginst5160 (R1240_U263, U3077, U3492);
  nand ginst5161 (R1240_U264, R1240_U13, R1240_U184);
  nand ginst5162 (R1240_U265, R1240_U261, R1240_U263);
  not ginst5163 (R1240_U266, R1240_U183);
  or ginst5164 (R1240_U267, U3076, U3494);
  nand ginst5165 (R1240_U268, U3076, U3494);
  not ginst5166 (R1240_U269, R1240_U181);
  not ginst5167 (R1240_U27, U3470);
  or ginst5168 (R1240_U270, U3071, U3496);
  nand ginst5169 (R1240_U271, U3071, U3496);
  not ginst5170 (R1240_U272, R1240_U105);
  or ginst5171 (R1240_U273, U3066, U3500);
  or ginst5172 (R1240_U274, U3070, U3498);
  not ginst5173 (R1240_U275, R1240_U90);
  nand ginst5174 (R1240_U276, R1240_U90, R1240_U91);
  nand ginst5175 (R1240_U277, R1240_U276, U3066);
  nand ginst5176 (R1240_U278, R1240_U275, U3500);
  nand ginst5177 (R1240_U279, R1240_U105, R1240_U9);
  not ginst5178 (R1240_U28, U3065);
  not ginst5179 (R1240_U280, R1240_U179);
  or ginst5180 (R1240_U281, U3073, U4037);
  or ginst5181 (R1240_U282, U3078, U3504);
  or ginst5182 (R1240_U283, U3072, U4036);
  not ginst5183 (R1240_U284, R1240_U80);
  nand ginst5184 (R1240_U285, R1240_U284, U4037);
  nand ginst5185 (R1240_U286, R1240_U103, R1240_U285);
  nand ginst5186 (R1240_U287, R1240_U80, R1240_U81);
  nand ginst5187 (R1240_U288, R1240_U286, R1240_U287);
  nand ginst5188 (R1240_U289, R1240_U11, R1240_U192);
  not ginst5189 (R1240_U29, U3472);
  nand ginst5190 (R1240_U290, U3072, U4036);
  nand ginst5191 (R1240_U291, R1240_U288, R1240_U289, R1240_U290);
  or ginst5192 (R1240_U292, U3079, U3502);
  or ginst5193 (R1240_U293, U3072, U4036);
  nand ginst5194 (R1240_U294, R1240_U291, R1240_U293);
  not ginst5195 (R1240_U295, R1240_U175);
  or ginst5196 (R1240_U296, U3058, U4035);
  nand ginst5197 (R1240_U297, U3058, U4035);
  not ginst5198 (R1240_U298, R1240_U94);
  or ginst5199 (R1240_U299, U3063, U4034);
  not ginst5200 (R1240_U30, U3061);
  nand ginst5201 (R1240_U300, R1240_U299, R1240_U94);
  nand ginst5202 (R1240_U301, U3063, U4034);
  not ginst5203 (R1240_U302, R1240_U172);
  or ginst5204 (R1240_U303, U3055, U4032);
  nand ginst5205 (R1240_U304, R1240_U185, R1240_U193);
  or ginst5206 (R1240_U305, U3062, U4033);
  or ginst5207 (R1240_U306, U3054, U4031);
  nand ginst5208 (R1240_U307, R1240_U149, R1240_U392);
  not ginst5209 (R1240_U308, R1240_U171);
  or ginst5210 (R1240_U309, U3050, U4030);
  not ginst5211 (R1240_U31, U3474);
  nand ginst5212 (R1240_U310, U3050, U4030);
  not ginst5213 (R1240_U311, R1240_U169);
  nand ginst5214 (R1240_U312, R1240_U169, U4029);
  not ginst5215 (R1240_U313, R1240_U167);
  nand ginst5216 (R1240_U314, R1240_U172, R1240_U305);
  not ginst5217 (R1240_U315, R1240_U100);
  or ginst5218 (R1240_U316, U3055, U4032);
  nand ginst5219 (R1240_U317, R1240_U100, R1240_U316);
  nand ginst5220 (R1240_U318, R1240_U151, R1240_U317);
  nand ginst5221 (R1240_U319, R1240_U190, R1240_U315);
  not ginst5222 (R1240_U32, U3057);
  nand ginst5223 (R1240_U320, U3054, U4031);
  nand ginst5224 (R1240_U321, R1240_U152, R1240_U319);
  or ginst5225 (R1240_U322, U3055, U4032);
  nand ginst5226 (R1240_U323, R1240_U179, R1240_U292);
  not ginst5227 (R1240_U324, R1240_U104);
  nand ginst5228 (R1240_U325, R1240_U10, R1240_U104);
  nand ginst5229 (R1240_U326, R1240_U153, R1240_U325);
  nand ginst5230 (R1240_U327, R1240_U288, R1240_U325);
  nand ginst5231 (R1240_U328, R1240_U327, R1240_U480);
  or ginst5232 (R1240_U329, U3078, U3504);
  not ginst5233 (R1240_U33, U3064);
  nand ginst5234 (R1240_U330, R1240_U104, R1240_U329);
  nand ginst5235 (R1240_U331, R1240_U154, R1240_U330);
  nand ginst5236 (R1240_U332, R1240_U324, R1240_U80);
  nand ginst5237 (R1240_U333, U3073, U4037);
  nand ginst5238 (R1240_U334, R1240_U155, R1240_U332);
  or ginst5239 (R1240_U335, U3075, U3468);
  not ginst5240 (R1240_U336, R1240_U178);
  or ginst5241 (R1240_U337, U3078, U3504);
  or ginst5242 (R1240_U338, U3070, U3498);
  nand ginst5243 (R1240_U339, R1240_U105, R1240_U338);
  nand ginst5244 (R1240_U34, U3057, U3474);
  nand ginst5245 (R1240_U340, R1240_U156, R1240_U339);
  nand ginst5246 (R1240_U341, R1240_U272, R1240_U90);
  nand ginst5247 (R1240_U342, U3066, U3500);
  nand ginst5248 (R1240_U343, R1240_U157, R1240_U341);
  or ginst5249 (R1240_U344, U3070, U3498);
  nand ginst5250 (R1240_U345, R1240_U184, R1240_U262);
  not ginst5251 (R1240_U346, R1240_U106);
  or ginst5252 (R1240_U347, U3069, U3490);
  nand ginst5253 (R1240_U348, R1240_U106, R1240_U347);
  nand ginst5254 (R1240_U349, R1240_U158, R1240_U348);
  not ginst5255 (R1240_U35, U3476);
  nand ginst5256 (R1240_U350, R1240_U189, R1240_U346);
  nand ginst5257 (R1240_U351, U3077, U3492);
  nand ginst5258 (R1240_U352, R1240_U159, R1240_U350);
  or ginst5259 (R1240_U353, U3069, U3490);
  or ginst5260 (R1240_U354, U3080, U3484);
  nand ginst5261 (R1240_U355, R1240_U354, R1240_U50);
  nand ginst5262 (R1240_U356, R1240_U160, R1240_U355);
  nand ginst5263 (R1240_U357, R1240_U188, R1240_U219);
  nand ginst5264 (R1240_U358, U3059, U3486);
  nand ginst5265 (R1240_U359, R1240_U161, R1240_U357);
  nand ginst5266 (R1240_U36, U3075, U3468);
  nand ginst5267 (R1240_U360, R1240_U188, R1240_U220);
  nand ginst5268 (R1240_U361, R1240_U217, R1240_U65);
  nand ginst5269 (R1240_U362, R1240_U227, R1240_U43);
  nand ginst5270 (R1240_U363, R1240_U241, R1240_U34);
  nand ginst5271 (R1240_U364, R1240_U197, R1240_U244);
  nand ginst5272 (R1240_U365, R1240_U190, R1240_U322);
  nand ginst5273 (R1240_U366, R1240_U305, R1240_U60);
  nand ginst5274 (R1240_U367, R1240_U337, R1240_U80);
  nand ginst5275 (R1240_U368, R1240_U292, R1240_U84);
  nand ginst5276 (R1240_U369, R1240_U344, R1240_U90);
  not ginst5277 (R1240_U37, U3464);
  nand ginst5278 (R1240_U370, R1240_U189, R1240_U353);
  nand ginst5279 (R1240_U371, R1240_U262, R1240_U72);
  nand ginst5280 (R1240_U372, U3051, U4029);
  nand ginst5281 (R1240_U373, R1240_U202, R1240_U4, R1240_U5);
  nand ginst5282 (R1240_U374, R1240_U201, R1240_U4, R1240_U5);
  not ginst5283 (R1240_U375, R1240_U45);
  not ginst5284 (R1240_U376, R1240_U102);
  nand ginst5285 (R1240_U377, R1240_U141, R1240_U51);
  nand ginst5286 (R1240_U378, R1240_U12, R1240_U45);
  nand ginst5287 (R1240_U379, R1240_U15, R1240_U184);
  not ginst5288 (R1240_U38, U3074);
  nand ginst5289 (R1240_U380, R1240_U265, R1240_U268);
  not ginst5290 (R1240_U381, R1240_U77);
  nand ginst5291 (R1240_U382, R1240_U143, R1240_U184);
  nand ginst5292 (R1240_U383, R1240_U270, R1240_U381);
  nand ginst5293 (R1240_U384, R1240_U105, R1240_U16);
  nand ginst5294 (R1240_U385, R1240_U102, R1240_U14);
  not ginst5295 (R1240_U386, R1240_U101);
  not ginst5296 (R1240_U387, R1240_U97);
  nand ginst5297 (R1240_U388, R1240_U105, R1240_U145);
  nand ginst5298 (R1240_U389, R1240_U101, R1240_U296);
  nand ginst5299 (R1240_U39, R1240_U131, R1240_U200);
  nand ginst5300 (R1240_U390, R1240_U303, U3054);
  nand ginst5301 (R1240_U391, R1240_U303, U4031);
  nand ginst5302 (R1240_U392, R1240_U298, R1240_U301);
  nand ginst5303 (R1240_U393, R1240_U185, R1240_U193, R1240_U309);
  nand ginst5304 (R1240_U394, R1240_U147, R1240_U17, R1240_U392);
  nand ginst5305 (R1240_U395, R1240_U309, R1240_U387);
  nand ginst5306 (R1240_U396, R1240_U190, R1240_U57);
  nand ginst5307 (R1240_U397, R1240_U190, R1240_U56);
  nand ginst5308 (R1240_U398, R1240_U49, U3080);
  nand ginst5309 (R1240_U399, R1240_U48, U3484);
  and ginst5310 (R1240_U4, R1240_U195, R1240_U196);
  not ginst5311 (R1240_U40, U3478);
  nand ginst5312 (R1240_U400, R1240_U398, R1240_U399);
  nand ginst5313 (R1240_U401, R1240_U360, R1240_U50);
  nand ginst5314 (R1240_U402, R1240_U219, R1240_U400);
  nand ginst5315 (R1240_U403, R1240_U46, U3081);
  nand ginst5316 (R1240_U404, R1240_U47, U3482);
  nand ginst5317 (R1240_U405, R1240_U403, R1240_U404);
  nand ginst5318 (R1240_U406, R1240_U162, R1240_U361);
  nand ginst5319 (R1240_U407, R1240_U216, R1240_U405);
  nand ginst5320 (R1240_U408, R1240_U44, U3067);
  nand ginst5321 (R1240_U409, R1240_U42, U3480);
  not ginst5322 (R1240_U41, U3068);
  nand ginst5323 (R1240_U410, R1240_U40, U3068);
  nand ginst5324 (R1240_U411, R1240_U41, U3478);
  nand ginst5325 (R1240_U412, R1240_U410, R1240_U411);
  nand ginst5326 (R1240_U413, R1240_U362, R1240_U51);
  nand ginst5327 (R1240_U414, R1240_U208, R1240_U412);
  nand ginst5328 (R1240_U415, R1240_U35, U3064);
  nand ginst5329 (R1240_U416, R1240_U33, U3476);
  nand ginst5330 (R1240_U417, R1240_U31, U3057);
  nand ginst5331 (R1240_U418, R1240_U32, U3474);
  nand ginst5332 (R1240_U419, R1240_U417, R1240_U418);
  not ginst5333 (R1240_U42, U3067);
  nand ginst5334 (R1240_U420, R1240_U363, R1240_U52);
  nand ginst5335 (R1240_U421, R1240_U234, R1240_U419);
  nand ginst5336 (R1240_U422, R1240_U29, U3061);
  nand ginst5337 (R1240_U423, R1240_U30, U3472);
  nand ginst5338 (R1240_U424, R1240_U422, R1240_U423);
  nand ginst5339 (R1240_U425, R1240_U163, R1240_U364);
  nand ginst5340 (R1240_U426, R1240_U243, R1240_U424);
  nand ginst5341 (R1240_U427, R1240_U27, U3065);
  nand ginst5342 (R1240_U428, R1240_U28, U3470);
  nand ginst5343 (R1240_U429, R1240_U165, U3052);
  nand ginst5344 (R1240_U43, U3068, U3478);
  nand ginst5345 (R1240_U430, R1240_U164, U4040);
  nand ginst5346 (R1240_U431, R1240_U165, U3052);
  nand ginst5347 (R1240_U432, R1240_U164, U4040);
  nand ginst5348 (R1240_U433, R1240_U431, R1240_U432);
  nand ginst5349 (R1240_U434, R1240_U166, R1240_U167);
  nand ginst5350 (R1240_U435, R1240_U313, R1240_U433);
  nand ginst5351 (R1240_U436, R1240_U99, U3051);
  nand ginst5352 (R1240_U437, R1240_U98, U4029);
  nand ginst5353 (R1240_U438, R1240_U99, U3051);
  nand ginst5354 (R1240_U439, R1240_U98, U4029);
  not ginst5355 (R1240_U44, U3480);
  nand ginst5356 (R1240_U440, R1240_U438, R1240_U439);
  nand ginst5357 (R1240_U441, R1240_U168, R1240_U169);
  nand ginst5358 (R1240_U442, R1240_U311, R1240_U440);
  nand ginst5359 (R1240_U443, R1240_U54, U3050);
  nand ginst5360 (R1240_U444, R1240_U55, U4030);
  nand ginst5361 (R1240_U445, R1240_U54, U3050);
  nand ginst5362 (R1240_U446, R1240_U55, U4030);
  nand ginst5363 (R1240_U447, R1240_U445, R1240_U446);
  nand ginst5364 (R1240_U448, R1240_U170, R1240_U171);
  nand ginst5365 (R1240_U449, R1240_U308, R1240_U447);
  nand ginst5366 (R1240_U45, R1240_U213, R1240_U214);
  nand ginst5367 (R1240_U450, R1240_U57, U3054);
  nand ginst5368 (R1240_U451, R1240_U56, U4031);
  nand ginst5369 (R1240_U452, R1240_U95, U3055);
  nand ginst5370 (R1240_U453, R1240_U96, U4032);
  nand ginst5371 (R1240_U454, R1240_U452, R1240_U453);
  nand ginst5372 (R1240_U455, R1240_U100, R1240_U365);
  nand ginst5373 (R1240_U456, R1240_U315, R1240_U454);
  nand ginst5374 (R1240_U457, R1240_U58, U3062);
  nand ginst5375 (R1240_U458, R1240_U59, U4033);
  nand ginst5376 (R1240_U459, R1240_U457, R1240_U458);
  not ginst5377 (R1240_U46, U3482);
  nand ginst5378 (R1240_U460, R1240_U172, R1240_U366);
  nand ginst5379 (R1240_U461, R1240_U302, R1240_U459);
  nand ginst5380 (R1240_U462, R1240_U92, U3063);
  nand ginst5381 (R1240_U463, R1240_U93, U4034);
  nand ginst5382 (R1240_U464, R1240_U92, U3063);
  nand ginst5383 (R1240_U465, R1240_U93, U4034);
  nand ginst5384 (R1240_U466, R1240_U464, R1240_U465);
  nand ginst5385 (R1240_U467, R1240_U173, R1240_U94);
  nand ginst5386 (R1240_U468, R1240_U298, R1240_U466);
  nand ginst5387 (R1240_U469, R1240_U61, U3058);
  not ginst5388 (R1240_U47, U3081);
  nand ginst5389 (R1240_U470, R1240_U62, U4035);
  nand ginst5390 (R1240_U471, R1240_U61, U3058);
  nand ginst5391 (R1240_U472, R1240_U62, U4035);
  nand ginst5392 (R1240_U473, R1240_U471, R1240_U472);
  nand ginst5393 (R1240_U474, R1240_U174, R1240_U175);
  nand ginst5394 (R1240_U475, R1240_U295, R1240_U473);
  nand ginst5395 (R1240_U476, R1240_U85, U3072);
  nand ginst5396 (R1240_U477, R1240_U86, U4036);
  nand ginst5397 (R1240_U478, R1240_U85, U3072);
  nand ginst5398 (R1240_U479, R1240_U86, U4036);
  not ginst5399 (R1240_U48, U3080);
  nand ginst5400 (R1240_U480, R1240_U478, R1240_U479);
  nand ginst5401 (R1240_U481, R1240_U81, U3073);
  nand ginst5402 (R1240_U482, R1240_U103, U4037);
  nand ginst5403 (R1240_U483, R1240_U178, R1240_U199);
  nand ginst5404 (R1240_U484, R1240_U177, R1240_U336);
  nand ginst5405 (R1240_U485, R1240_U78, U3078);
  nand ginst5406 (R1240_U486, R1240_U79, U3504);
  nand ginst5407 (R1240_U487, R1240_U485, R1240_U486);
  nand ginst5408 (R1240_U488, R1240_U104, R1240_U367);
  nand ginst5409 (R1240_U489, R1240_U324, R1240_U487);
  not ginst5410 (R1240_U49, U3484);
  nand ginst5411 (R1240_U490, R1240_U82, U3079);
  nand ginst5412 (R1240_U491, R1240_U83, U3502);
  nand ginst5413 (R1240_U492, R1240_U490, R1240_U491);
  nand ginst5414 (R1240_U493, R1240_U179, R1240_U368);
  nand ginst5415 (R1240_U494, R1240_U280, R1240_U492);
  nand ginst5416 (R1240_U495, R1240_U91, U3066);
  nand ginst5417 (R1240_U496, R1240_U89, U3500);
  nand ginst5418 (R1240_U497, R1240_U87, U3070);
  nand ginst5419 (R1240_U498, R1240_U88, U3498);
  nand ginst5420 (R1240_U499, R1240_U497, R1240_U498);
  and ginst5421 (R1240_U5, R1240_U197, R1240_U198);
  nand ginst5422 (R1240_U50, R1240_U218, R1240_U65);
  nand ginst5423 (R1240_U500, R1240_U105, R1240_U369);
  nand ginst5424 (R1240_U501, R1240_U272, R1240_U499);
  nand ginst5425 (R1240_U502, R1240_U63, U3071);
  nand ginst5426 (R1240_U503, R1240_U64, U3496);
  nand ginst5427 (R1240_U504, R1240_U63, U3071);
  nand ginst5428 (R1240_U505, R1240_U64, U3496);
  nand ginst5429 (R1240_U506, R1240_U504, R1240_U505);
  nand ginst5430 (R1240_U507, R1240_U180, R1240_U181);
  nand ginst5431 (R1240_U508, R1240_U269, R1240_U506);
  nand ginst5432 (R1240_U509, R1240_U75, U3076);
  nand ginst5433 (R1240_U51, R1240_U132, R1240_U133);
  nand ginst5434 (R1240_U510, R1240_U76, U3494);
  nand ginst5435 (R1240_U511, R1240_U75, U3076);
  nand ginst5436 (R1240_U512, R1240_U76, U3494);
  nand ginst5437 (R1240_U513, R1240_U511, R1240_U512);
  nand ginst5438 (R1240_U514, R1240_U182, R1240_U183);
  nand ginst5439 (R1240_U515, R1240_U266, R1240_U513);
  nand ginst5440 (R1240_U516, R1240_U73, U3077);
  nand ginst5441 (R1240_U517, R1240_U74, U3492);
  nand ginst5442 (R1240_U518, R1240_U68, U3069);
  nand ginst5443 (R1240_U519, R1240_U69, U3490);
  nand ginst5444 (R1240_U52, R1240_U136, R1240_U232);
  nand ginst5445 (R1240_U520, R1240_U518, R1240_U519);
  nand ginst5446 (R1240_U521, R1240_U106, R1240_U370);
  nand ginst5447 (R1240_U522, R1240_U346, R1240_U520);
  nand ginst5448 (R1240_U523, R1240_U70, U3060);
  nand ginst5449 (R1240_U524, R1240_U71, U3488);
  nand ginst5450 (R1240_U525, R1240_U523, R1240_U524);
  nand ginst5451 (R1240_U526, R1240_U184, R1240_U371);
  nand ginst5452 (R1240_U527, R1240_U256, R1240_U525);
  nand ginst5453 (R1240_U528, R1240_U66, U3059);
  nand ginst5454 (R1240_U529, R1240_U67, U3486);
  nand ginst5455 (R1240_U53, R1240_U228, R1240_U229);
  nand ginst5456 (R1240_U530, R1240_U37, U3074);
  nand ginst5457 (R1240_U531, R1240_U38, U3464);
  not ginst5458 (R1240_U54, U4030);
  not ginst5459 (R1240_U55, U3050);
  not ginst5460 (R1240_U56, U3054);
  not ginst5461 (R1240_U57, U4031);
  not ginst5462 (R1240_U58, U4033);
  not ginst5463 (R1240_U59, U3062);
  and ginst5464 (R1240_U6, R1240_U209, R1240_U210);
  nand ginst5465 (R1240_U60, U3062, U4033);
  not ginst5466 (R1240_U61, U4035);
  not ginst5467 (R1240_U62, U3058);
  not ginst5468 (R1240_U63, U3496);
  not ginst5469 (R1240_U64, U3071);
  nand ginst5470 (R1240_U65, U3081, U3482);
  not ginst5471 (R1240_U66, U3486);
  not ginst5472 (R1240_U67, U3059);
  not ginst5473 (R1240_U68, U3490);
  not ginst5474 (R1240_U69, U3069);
  and ginst5475 (R1240_U7, R1240_U249, R1240_U250);
  not ginst5476 (R1240_U70, U3488);
  not ginst5477 (R1240_U71, U3060);
  nand ginst5478 (R1240_U72, U3060, U3488);
  not ginst5479 (R1240_U73, U3492);
  not ginst5480 (R1240_U74, U3077);
  not ginst5481 (R1240_U75, U3494);
  not ginst5482 (R1240_U76, U3076);
  nand ginst5483 (R1240_U77, R1240_U267, R1240_U380);
  not ginst5484 (R1240_U78, U3504);
  not ginst5485 (R1240_U79, U3078);
  and ginst5486 (R1240_U8, R1240_U257, R1240_U258);
  nand ginst5487 (R1240_U80, U3078, U3504);
  not ginst5488 (R1240_U81, U4037);
  not ginst5489 (R1240_U82, U3502);
  not ginst5490 (R1240_U83, U3079);
  nand ginst5491 (R1240_U84, U3079, U3502);
  not ginst5492 (R1240_U85, U4036);
  not ginst5493 (R1240_U86, U3072);
  not ginst5494 (R1240_U87, U3498);
  not ginst5495 (R1240_U88, U3070);
  not ginst5496 (R1240_U89, U3066);
  and ginst5497 (R1240_U9, R1240_U273, R1240_U274);
  nand ginst5498 (R1240_U90, U3070, U3498);
  not ginst5499 (R1240_U91, U3500);
  not ginst5500 (R1240_U92, U4034);
  not ginst5501 (R1240_U93, U3063);
  nand ginst5502 (R1240_U94, R1240_U146, R1240_U388);
  not ginst5503 (R1240_U95, U4032);
  not ginst5504 (R1240_U96, U3055);
  nand ginst5505 (R1240_U97, R1240_U306, R1240_U396, R1240_U397);
  not ginst5506 (R1240_U98, U3051);
  not ginst5507 (R1240_U99, U4029);
  and ginst5508 (R1282_U10, R1282_U103, R1282_U14);
  not ginst5509 (R1282_U100, R1282_U35);
  not ginst5510 (R1282_U101, R1282_U15);
  nand ginst5511 (R1282_U102, R1282_U14, U3480);
  nand ginst5512 (R1282_U103, R1282_U98, U3478);
  nand ginst5513 (R1282_U104, R1282_U13, U3476);
  nand ginst5514 (R1282_U105, R1282_U96, U3474);
  nand ginst5515 (R1282_U106, R1282_U12, U3472);
  not ginst5516 (R1282_U107, R1282_U93);
  not ginst5517 (R1282_U108, R1282_U21);
  not ginst5518 (R1282_U109, R1282_U88);
  and ginst5519 (R1282_U11, R1282_U102, R1282_U35);
  not ginst5520 (R1282_U110, R1282_U22);
  not ginst5521 (R1282_U111, R1282_U83);
  not ginst5522 (R1282_U112, R1282_U23);
  not ginst5523 (R1282_U113, R1282_U78);
  not ginst5524 (R1282_U114, R1282_U24);
  not ginst5525 (R1282_U115, R1282_U73);
  not ginst5526 (R1282_U116, R1282_U25);
  not ginst5527 (R1282_U117, R1282_U66);
  not ginst5528 (R1282_U118, R1282_U26);
  not ginst5529 (R1282_U119, R1282_U61);
  or ginst5530 (R1282_U12, U3464, U3468, U3470);
  not ginst5531 (R1282_U120, R1282_U27);
  not ginst5532 (R1282_U121, R1282_U56);
  not ginst5533 (R1282_U122, R1282_U28);
  not ginst5534 (R1282_U123, R1282_U51);
  not ginst5535 (R1282_U124, R1282_U29);
  not ginst5536 (R1282_U125, R1282_U46);
  not ginst5537 (R1282_U126, R1282_U30);
  not ginst5538 (R1282_U127, R1282_U41);
  not ginst5539 (R1282_U128, R1282_U38);
  or ginst5540 (R1282_U129, U3464, U3468);
  nand ginst5541 (R1282_U13, R1282_U19, R1282_U20, R1282_U95);
  nand ginst5542 (R1282_U130, R1282_U129, U3470);
  nand ginst5543 (R1282_U131, R1282_U15, U3484);
  nand ginst5544 (R1282_U132, R1282_U101, R1282_U32);
  nand ginst5545 (R1282_U133, R1282_U35, U3482);
  nand ginst5546 (R1282_U134, R1282_U100, R1282_U34);
  nand ginst5547 (R1282_U135, R1282_U38, U4038);
  nand ginst5548 (R1282_U136, R1282_U128, R1282_U37);
  nand ginst5549 (R1282_U137, R1282_U41, U4039);
  nand ginst5550 (R1282_U138, R1282_U127, R1282_U40);
  nand ginst5551 (R1282_U139, R1282_U30, U4040);
  nand ginst5552 (R1282_U14, R1282_U17, R1282_U18, R1282_U97);
  nand ginst5553 (R1282_U140, R1282_U126, R1282_U43);
  nand ginst5554 (R1282_U141, R1282_U46, U4029);
  nand ginst5555 (R1282_U142, R1282_U125, R1282_U45);
  nand ginst5556 (R1282_U143, R1282_U29, U4030);
  nand ginst5557 (R1282_U144, R1282_U124, R1282_U48);
  nand ginst5558 (R1282_U145, R1282_U51, U4031);
  nand ginst5559 (R1282_U146, R1282_U123, R1282_U50);
  nand ginst5560 (R1282_U147, R1282_U28, U4032);
  nand ginst5561 (R1282_U148, R1282_U122, R1282_U53);
  nand ginst5562 (R1282_U149, R1282_U56, U4033);
  nand ginst5563 (R1282_U15, R1282_U16, R1282_U34, R1282_U99);
  nand ginst5564 (R1282_U150, R1282_U121, R1282_U55);
  nand ginst5565 (R1282_U151, R1282_U27, U4034);
  nand ginst5566 (R1282_U152, R1282_U120, R1282_U58);
  nand ginst5567 (R1282_U153, R1282_U61, U4035);
  nand ginst5568 (R1282_U154, R1282_U119, R1282_U60);
  nand ginst5569 (R1282_U155, R1282_U26, U4036);
  nand ginst5570 (R1282_U156, R1282_U118, R1282_U63);
  nand ginst5571 (R1282_U157, R1282_U66, U4037);
  nand ginst5572 (R1282_U158, R1282_U117, R1282_U65);
  nand ginst5573 (R1282_U159, R1282_U69, U3468);
  not ginst5574 (R1282_U16, U3480);
  nand ginst5575 (R1282_U160, R1282_U68, U3464);
  nand ginst5576 (R1282_U161, R1282_U25, U3504);
  nand ginst5577 (R1282_U162, R1282_U116, R1282_U70);
  nand ginst5578 (R1282_U163, R1282_U73, U3502);
  nand ginst5579 (R1282_U164, R1282_U115, R1282_U72);
  nand ginst5580 (R1282_U165, R1282_U24, U3500);
  nand ginst5581 (R1282_U166, R1282_U114, R1282_U75);
  nand ginst5582 (R1282_U167, R1282_U78, U3498);
  nand ginst5583 (R1282_U168, R1282_U113, R1282_U77);
  nand ginst5584 (R1282_U169, R1282_U23, U3496);
  not ginst5585 (R1282_U17, U3478);
  nand ginst5586 (R1282_U170, R1282_U112, R1282_U80);
  nand ginst5587 (R1282_U171, R1282_U83, U3494);
  nand ginst5588 (R1282_U172, R1282_U111, R1282_U82);
  nand ginst5589 (R1282_U173, R1282_U22, U3492);
  nand ginst5590 (R1282_U174, R1282_U110, R1282_U85);
  nand ginst5591 (R1282_U175, R1282_U88, U3490);
  nand ginst5592 (R1282_U176, R1282_U109, R1282_U87);
  nand ginst5593 (R1282_U177, R1282_U21, U3488);
  nand ginst5594 (R1282_U178, R1282_U108, R1282_U90);
  nand ginst5595 (R1282_U179, R1282_U93, U3486);
  not ginst5596 (R1282_U18, U3476);
  nand ginst5597 (R1282_U180, R1282_U107, R1282_U92);
  not ginst5598 (R1282_U19, U3474);
  not ginst5599 (R1282_U20, U3472);
  nand ginst5600 (R1282_U21, R1282_U101, R1282_U32, R1282_U92);
  nand ginst5601 (R1282_U22, R1282_U108, R1282_U87, R1282_U90);
  nand ginst5602 (R1282_U23, R1282_U110, R1282_U82, R1282_U85);
  nand ginst5603 (R1282_U24, R1282_U112, R1282_U77, R1282_U80);
  nand ginst5604 (R1282_U25, R1282_U114, R1282_U72, R1282_U75);
  nand ginst5605 (R1282_U26, R1282_U116, R1282_U65, R1282_U70);
  nand ginst5606 (R1282_U27, R1282_U118, R1282_U60, R1282_U63);
  nand ginst5607 (R1282_U28, R1282_U120, R1282_U55, R1282_U58);
  nand ginst5608 (R1282_U29, R1282_U122, R1282_U50, R1282_U53);
  nand ginst5609 (R1282_U30, R1282_U124, R1282_U45, R1282_U48);
  nand ginst5610 (R1282_U31, R1282_U159, R1282_U160);
  not ginst5611 (R1282_U32, U3484);
  and ginst5612 (R1282_U33, R1282_U131, R1282_U132);
  not ginst5613 (R1282_U34, U3482);
  nand ginst5614 (R1282_U35, R1282_U16, R1282_U99);
  and ginst5615 (R1282_U36, R1282_U133, R1282_U134);
  not ginst5616 (R1282_U37, U4038);
  nand ginst5617 (R1282_U38, R1282_U126, R1282_U40, R1282_U43);
  and ginst5618 (R1282_U39, R1282_U135, R1282_U136);
  not ginst5619 (R1282_U40, U4039);
  nand ginst5620 (R1282_U41, R1282_U126, R1282_U43);
  and ginst5621 (R1282_U42, R1282_U137, R1282_U138);
  not ginst5622 (R1282_U43, U4040);
  and ginst5623 (R1282_U44, R1282_U139, R1282_U140);
  not ginst5624 (R1282_U45, U4029);
  nand ginst5625 (R1282_U46, R1282_U124, R1282_U48);
  and ginst5626 (R1282_U47, R1282_U141, R1282_U142);
  not ginst5627 (R1282_U48, U4030);
  and ginst5628 (R1282_U49, R1282_U143, R1282_U144);
  not ginst5629 (R1282_U50, U4031);
  nand ginst5630 (R1282_U51, R1282_U122, R1282_U53);
  and ginst5631 (R1282_U52, R1282_U145, R1282_U146);
  not ginst5632 (R1282_U53, U4032);
  and ginst5633 (R1282_U54, R1282_U147, R1282_U148);
  not ginst5634 (R1282_U55, U4033);
  nand ginst5635 (R1282_U56, R1282_U120, R1282_U58);
  and ginst5636 (R1282_U57, R1282_U149, R1282_U150);
  not ginst5637 (R1282_U58, U4034);
  and ginst5638 (R1282_U59, R1282_U151, R1282_U152);
  and ginst5639 (R1282_U6, R1282_U12, R1282_U130);
  not ginst5640 (R1282_U60, U4035);
  nand ginst5641 (R1282_U61, R1282_U118, R1282_U63);
  and ginst5642 (R1282_U62, R1282_U153, R1282_U154);
  not ginst5643 (R1282_U63, U4036);
  and ginst5644 (R1282_U64, R1282_U155, R1282_U156);
  not ginst5645 (R1282_U65, U4037);
  nand ginst5646 (R1282_U66, R1282_U116, R1282_U70);
  and ginst5647 (R1282_U67, R1282_U157, R1282_U158);
  not ginst5648 (R1282_U68, U3468);
  not ginst5649 (R1282_U69, U3464);
  and ginst5650 (R1282_U7, R1282_U106, R1282_U96);
  not ginst5651 (R1282_U70, U3504);
  and ginst5652 (R1282_U71, R1282_U161, R1282_U162);
  not ginst5653 (R1282_U72, U3502);
  nand ginst5654 (R1282_U73, R1282_U114, R1282_U75);
  and ginst5655 (R1282_U74, R1282_U163, R1282_U164);
  not ginst5656 (R1282_U75, U3500);
  and ginst5657 (R1282_U76, R1282_U165, R1282_U166);
  not ginst5658 (R1282_U77, U3498);
  nand ginst5659 (R1282_U78, R1282_U112, R1282_U80);
  and ginst5660 (R1282_U79, R1282_U167, R1282_U168);
  and ginst5661 (R1282_U8, R1282_U105, R1282_U13);
  not ginst5662 (R1282_U80, U3496);
  and ginst5663 (R1282_U81, R1282_U169, R1282_U170);
  not ginst5664 (R1282_U82, U3494);
  nand ginst5665 (R1282_U83, R1282_U110, R1282_U85);
  and ginst5666 (R1282_U84, R1282_U171, R1282_U172);
  not ginst5667 (R1282_U85, U3492);
  and ginst5668 (R1282_U86, R1282_U173, R1282_U174);
  not ginst5669 (R1282_U87, U3490);
  nand ginst5670 (R1282_U88, R1282_U108, R1282_U90);
  and ginst5671 (R1282_U89, R1282_U175, R1282_U176);
  and ginst5672 (R1282_U9, R1282_U104, R1282_U98);
  not ginst5673 (R1282_U90, U3488);
  and ginst5674 (R1282_U91, R1282_U177, R1282_U178);
  not ginst5675 (R1282_U92, U3486);
  nand ginst5676 (R1282_U93, R1282_U101, R1282_U32);
  and ginst5677 (R1282_U94, R1282_U179, R1282_U180);
  not ginst5678 (R1282_U95, R1282_U12);
  nand ginst5679 (R1282_U96, R1282_U20, R1282_U95);
  not ginst5680 (R1282_U97, R1282_U13);
  nand ginst5681 (R1282_U98, R1282_U18, R1282_U97);
  not ginst5682 (R1282_U99, R1282_U14);
  nand ginst5683 (R1309_U10, R1309_U7, U3056);
  not ginst5684 (R1309_U6, U3056);
  not ginst5685 (R1309_U7, U3053);
  and ginst5686 (R1309_U8, R1309_U10, R1309_U9);
  nand ginst5687 (R1309_U9, R1309_U6, U3053);
  and ginst5688 (R1347_U10, R1347_U11, R1347_U83);
  and ginst5689 (R1347_U100, R1347_U41, U3604);
  and ginst5690 (R1347_U101, R1347_U43, U3600);
  and ginst5691 (R1347_U102, R1347_U35, U3599);
  and ginst5692 (R1347_U103, R1347_U133, R1347_U151, R1347_U165);
  and ginst5693 (R1347_U104, R1347_U166, R1347_U167);
  and ginst5694 (R1347_U105, R1347_U168, R1347_U169, R1347_U170, R1347_U176);
  and ginst5695 (R1347_U106, R1347_U177, R1347_U178);
  and ginst5696 (R1347_U107, R1347_U108, R1347_U179);
  and ginst5697 (R1347_U108, R1347_U186, R1347_U188);
  and ginst5698 (R1347_U109, R1347_U189, R1347_U190);
  and ginst5699 (R1347_U11, R1347_U183, R1347_U78, R1347_U79);
  and ginst5700 (R1347_U110, R1347_U109, R1347_U206);
  and ginst5701 (R1347_U111, R1347_U106, R1347_U107, R1347_U110, R1347_U207);
  and ginst5702 (R1347_U112, R1347_U61, U4034);
  and ginst5703 (R1347_U113, R1347_U192, R1347_U193);
  and ginst5704 (R1347_U114, R1347_U123, R1347_U132);
  and ginst5705 (R1347_U115, R1347_U12, R1347_U197);
  and ginst5706 (R1347_U116, R1347_U115, R1347_U210);
  and ginst5707 (R1347_U117, R1347_U67, U3589);
  and ginst5708 (R1347_U118, R1347_U120, R1347_U212);
  and ginst5709 (R1347_U119, R1347_U199, R1347_U201, R1347_U204);
  and ginst5710 (R1347_U12, R1347_U132, R1347_U209);
  and ginst5711 (R1347_U120, R1347_U119, R1347_U205);
  not ginst5712 (R1347_U121, U3613);
  not ginst5713 (R1347_U122, U4040);
  not ginst5714 (R1347_U123, U4029);
  not ginst5715 (R1347_U124, U3595);
  nand ginst5716 (R1347_U125, R1347_U202, R1347_U203);
  nand ginst5717 (R1347_U126, R1347_U131, R1347_U208);
  nand ginst5718 (R1347_U127, R1347_U194, U4032);
  nand ginst5719 (R1347_U128, R1347_U69, U3588);
  nand ginst5720 (R1347_U129, R1347_U122, R1347_U128, R1347_U130);
  and ginst5721 (R1347_U13, R1347_U118, R1347_U198);
  nand ginst5722 (R1347_U130, R1347_U68, U4039);
  nand ginst5723 (R1347_U131, R1347_U114, R1347_U209);
  nand ginst5724 (R1347_U132, R1347_U71, U4030);
  nand ginst5725 (R1347_U133, R1347_U63, U3596);
  nand ginst5726 (R1347_U134, R1347_U56, U3498);
  nand ginst5727 (R1347_U135, R1347_U42, U3602);
  nand ginst5728 (R1347_U136, R1347_U38, U3603);
  not ginst5729 (R1347_U137, R1347_U40);
  nand ginst5730 (R1347_U138, R1347_U55, U3496);
  nand ginst5731 (R1347_U139, R1347_U52, U3486);
  not ginst5732 (R1347_U14, U3596);
  nand ginst5733 (R1347_U140, R1347_U25, U3612);
  nand ginst5734 (R1347_U141, R1347_U51, U3484);
  nand ginst5735 (R1347_U142, R1347_U49, U3480);
  nand ginst5736 (R1347_U143, R1347_U50, U3482);
  nand ginst5737 (R1347_U144, R1347_U48, U3478);
  nand ginst5738 (R1347_U145, R1347_U47, U3476);
  nand ginst5739 (R1347_U146, R1347_U46, U3474);
  nand ginst5740 (R1347_U147, R1347_U45, U3472);
  nand ginst5741 (R1347_U148, R1347_U140, R1347_U73);
  nand ginst5742 (R1347_U149, R1347_U44, U3470);
  not ginst5743 (R1347_U15, U3486);
  nand ginst5744 (R1347_U150, R1347_U23, U3468);
  nand ginst5745 (R1347_U151, R1347_U10, R1347_U8, R1347_U86);
  nand ginst5746 (R1347_U152, R1347_U29, U3609);
  nand ginst5747 (R1347_U153, R1347_U33, U3608);
  not ginst5748 (R1347_U154, R1347_U31);
  nand ginst5749 (R1347_U155, R1347_U18, U3583);
  nand ginst5750 (R1347_U156, R1347_U16, U3582);
  nand ginst5751 (R1347_U157, R1347_U155, R1347_U156);
  nand ginst5752 (R1347_U158, R1347_U21, U3587);
  nand ginst5753 (R1347_U159, R1347_U20, U3586);
  not ginst5754 (R1347_U16, U3484);
  nand ginst5755 (R1347_U160, R1347_U158, R1347_U159);
  nand ginst5756 (R1347_U161, R1347_U160, R1347_U89);
  nand ginst5757 (R1347_U162, R1347_U19, U3585);
  nand ginst5758 (R1347_U163, R1347_U17, U3584);
  nand ginst5759 (R1347_U164, R1347_U161, R1347_U90);
  nand ginst5760 (R1347_U165, R1347_U10, R1347_U24, R1347_U8, U3601);
  nand ginst5761 (R1347_U166, R1347_U10, R1347_U88);
  nand ginst5762 (R1347_U167, R1347_U10, R1347_U91);
  nand ginst5763 (R1347_U168, R1347_U10, R1347_U93);
  nand ginst5764 (R1347_U169, R1347_U10, R1347_U94);
  not ginst5765 (R1347_U17, U3480);
  nand ginst5766 (R1347_U170, R1347_U10, R1347_U95);
  nand ginst5767 (R1347_U171, R1347_U33, U3608);
  nand ginst5768 (R1347_U172, R1347_U171, R1347_U74);
  nand ginst5769 (R1347_U173, R1347_U154, R1347_U75);
  nand ginst5770 (R1347_U174, R1347_U28, U3492);
  nand ginst5771 (R1347_U175, R1347_U54, U3494);
  nand ginst5772 (R1347_U176, R1347_U11, R1347_U96);
  nand ginst5773 (R1347_U177, R1347_U11, R1347_U98);
  nand ginst5774 (R1347_U178, R1347_U11, R1347_U99);
  nand ginst5775 (R1347_U179, R1347_U100, R1347_U11);
  not ginst5776 (R1347_U18, U3482);
  nand ginst5777 (R1347_U180, R1347_U59, U4036);
  nand ginst5778 (R1347_U181, R1347_U60, U4035);
  nand ginst5779 (R1347_U182, R1347_U135, R1347_U76);
  nand ginst5780 (R1347_U183, R1347_U137, R1347_U77);
  nand ginst5781 (R1347_U184, R1347_U37, U3504);
  nand ginst5782 (R1347_U185, R1347_U58, U4037);
  nand ginst5783 (R1347_U186, R1347_U101, R1347_U9);
  nand ginst5784 (R1347_U187, R1347_U60, U4035);
  nand ginst5785 (R1347_U188, R1347_U102, R1347_U187);
  nand ginst5786 (R1347_U189, R1347_U36, U3598);
  not ginst5787 (R1347_U19, U3478);
  nand ginst5788 (R1347_U190, R1347_U62, U3597);
  nand ginst5789 (R1347_U191, R1347_U103, R1347_U104, R1347_U105, R1347_U111);
  nand ginst5790 (R1347_U192, R1347_U112, R1347_U133);
  nand ginst5791 (R1347_U193, R1347_U14, U4033);
  nand ginst5792 (R1347_U194, R1347_U113, R1347_U191);
  nand ginst5793 (R1347_U195, R1347_U124, U4032);
  nand ginst5794 (R1347_U196, R1347_U124, R1347_U194);
  nand ginst5795 (R1347_U197, R1347_U72, U4031);
  nand ginst5796 (R1347_U198, R1347_U116, R1347_U127, R1347_U195, R1347_U196);
  nand ginst5797 (R1347_U199, R1347_U117, R1347_U128);
  not ginst5798 (R1347_U20, U3476);
  nand ginst5799 (R1347_U200, R1347_U68, U4039);
  nand ginst5800 (R1347_U201, R1347_U122, R1347_U128, R1347_U200, U3591);
  nand ginst5801 (R1347_U202, R1347_U65, U3593);
  nand ginst5802 (R1347_U203, R1347_U64, U3594);
  nand ginst5803 (R1347_U204, R1347_U66, U4038);
  nand ginst5804 (R1347_U205, R1347_U123, R1347_U209, U3592);
  nand ginst5805 (R1347_U206, R1347_U11, R1347_U40);
  nand ginst5806 (R1347_U207, R1347_U10, R1347_U31);
  nand ginst5807 (R1347_U208, R1347_U12, U3592);
  nand ginst5808 (R1347_U209, R1347_U129, R1347_U211);
  not ginst5809 (R1347_U21, U3474);
  nand ginst5810 (R1347_U210, R1347_U131, R1347_U70);
  nand ginst5811 (R1347_U211, R1347_U128, R1347_U130, U3591);
  nand ginst5812 (R1347_U212, R1347_U125, R1347_U126);
  not ginst5813 (R1347_U22, U3472);
  not ginst5814 (R1347_U23, U3612);
  not ginst5815 (R1347_U24, U3470);
  not ginst5816 (R1347_U25, U3468);
  not ginst5817 (R1347_U26, U3498);
  not ginst5818 (R1347_U27, U3496);
  not ginst5819 (R1347_U28, U3608);
  not ginst5820 (R1347_U29, U3490);
  not ginst5821 (R1347_U30, U3609);
  nand ginst5822 (R1347_U31, R1347_U152, R1347_U153);
  not ginst5823 (R1347_U32, U3488);
  not ginst5824 (R1347_U33, U3492);
  not ginst5825 (R1347_U34, U3494);
  not ginst5826 (R1347_U35, U4036);
  not ginst5827 (R1347_U36, U4035);
  not ginst5828 (R1347_U37, U3602);
  not ginst5829 (R1347_U38, U3502);
  not ginst5830 (R1347_U39, U3603);
  nand ginst5831 (R1347_U40, R1347_U135, R1347_U136);
  not ginst5832 (R1347_U41, U3500);
  not ginst5833 (R1347_U42, U3504);
  not ginst5834 (R1347_U43, U4037);
  not ginst5835 (R1347_U44, U3601);
  not ginst5836 (R1347_U45, U3590);
  not ginst5837 (R1347_U46, U3587);
  not ginst5838 (R1347_U47, U3586);
  not ginst5839 (R1347_U48, U3585);
  not ginst5840 (R1347_U49, U3584);
  not ginst5841 (R1347_U50, U3583);
  not ginst5842 (R1347_U51, U3582);
  not ginst5843 (R1347_U52, U3611);
  not ginst5844 (R1347_U53, U3610);
  not ginst5845 (R1347_U54, U3607);
  not ginst5846 (R1347_U55, U3606);
  not ginst5847 (R1347_U56, U3605);
  not ginst5848 (R1347_U57, U3604);
  not ginst5849 (R1347_U58, U3600);
  not ginst5850 (R1347_U59, U3599);
  and ginst5851 (R1347_U6, R1347_U139, R1347_U141, R1347_U142, R1347_U143);
  not ginst5852 (R1347_U60, U3598);
  not ginst5853 (R1347_U61, U3597);
  not ginst5854 (R1347_U62, U4034);
  not ginst5855 (R1347_U63, U4033);
  not ginst5856 (R1347_U64, U4031);
  not ginst5857 (R1347_U65, U4030);
  not ginst5858 (R1347_U66, U3588);
  not ginst5859 (R1347_U67, U4039);
  not ginst5860 (R1347_U68, U3589);
  not ginst5861 (R1347_U69, U4038);
  and ginst5862 (R1347_U7, R1347_U6, R1347_U84);
  not ginst5863 (R1347_U70, U3592);
  not ginst5864 (R1347_U71, U3593);
  not ginst5865 (R1347_U72, U3594);
  and ginst5866 (R1347_U73, R1347_U121, U3464);
  and ginst5867 (R1347_U74, R1347_U30, U3490);
  and ginst5868 (R1347_U75, R1347_U53, U3488);
  and ginst5869 (R1347_U76, R1347_U39, U3502);
  and ginst5870 (R1347_U77, R1347_U57, U3500);
  and ginst5871 (R1347_U78, R1347_U182, R1347_U184);
  and ginst5872 (R1347_U79, R1347_U185, R1347_U9);
  and ginst5873 (R1347_U8, R1347_U147, R1347_U7);
  and ginst5874 (R1347_U80, R1347_U134, R1347_U138);
  and ginst5875 (R1347_U81, R1347_U172, R1347_U80);
  and ginst5876 (R1347_U82, R1347_U174, R1347_U175);
  and ginst5877 (R1347_U83, R1347_U173, R1347_U81, R1347_U82);
  and ginst5878 (R1347_U84, R1347_U144, R1347_U145, R1347_U146);
  and ginst5879 (R1347_U85, R1347_U149, R1347_U150);
  and ginst5880 (R1347_U86, R1347_U148, R1347_U85);
  and ginst5881 (R1347_U87, R1347_U22, U3590);
  and ginst5882 (R1347_U88, R1347_U7, R1347_U87);
  and ginst5883 (R1347_U89, R1347_U144, R1347_U145);
  and ginst5884 (R1347_U9, R1347_U180, R1347_U181);
  and ginst5885 (R1347_U90, R1347_U162, R1347_U163);
  and ginst5886 (R1347_U91, R1347_U164, R1347_U6);
  and ginst5887 (R1347_U92, R1347_U139, R1347_U141);
  and ginst5888 (R1347_U93, R1347_U157, R1347_U92);
  and ginst5889 (R1347_U94, R1347_U15, U3611);
  and ginst5890 (R1347_U95, R1347_U32, U3610);
  and ginst5891 (R1347_U96, R1347_U134, R1347_U138, R1347_U34, U3607);
  and ginst5892 (R1347_U97, R1347_U27, U3606);
  and ginst5893 (R1347_U98, R1347_U134, R1347_U97);
  and ginst5894 (R1347_U99, R1347_U26, U3605);
  and ginst5895 (R1352_U6, R1352_U7, U3056);
  not ginst5896 (R1352_U7, U3053);
  and ginst5897 (R1375_U10, R1375_U9, R1375_U98);
  and ginst5898 (R1375_U100, R1375_U158, R1375_U24);
  and ginst5899 (R1375_U101, R1375_U15, R1375_U65);
  and ginst5900 (R1375_U102, R1375_U13, U3468);
  and ginst5901 (R1375_U103, R1375_U189, R1375_U190);
  and ginst5902 (R1375_U104, R1375_U156, R1375_U192);
  and ginst5903 (R1375_U105, R1375_U10, R1375_U100, R1375_U12, R1375_U14, R1375_U15);
  and ginst5904 (R1375_U106, R1375_U156, R1375_U53);
  and ginst5905 (R1375_U107, R1375_U15, R1375_U166);
  and ginst5906 (R1375_U108, R1375_U15, R1375_U56);
  and ginst5907 (R1375_U109, R1375_U158, R1375_U165, R1375_U178);
  and ginst5908 (R1375_U11, R1375_U181, R1375_U182);
  and ginst5909 (R1375_U110, R1375_U15, R1375_U60);
  and ginst5910 (R1375_U111, R1375_U15, R1375_U44);
  and ginst5911 (R1375_U112, R1375_U8, U3496);
  and ginst5912 (R1375_U113, R1375_U156, R1375_U54);
  and ginst5913 (R1375_U114, R1375_U15, U3478);
  and ginst5914 (R1375_U115, R1375_U156, R1375_U39);
  and ginst5915 (R1375_U116, R1375_U100, R1375_U12, R1375_U15, R1375_U19, U3476);
  and ginst5916 (R1375_U117, R1375_U156, R1375_U184, R1375_U36);
  and ginst5917 (R1375_U118, R1375_U15, R1375_U50);
  and ginst5918 (R1375_U119, R1375_U15, R1375_U43);
  and ginst5919 (R1375_U12, R1375_U183, R1375_U23);
  and ginst5920 (R1375_U120, R1375_U15, R1375_U58);
  and ginst5921 (R1375_U121, R1375_U11, U3480);
  and ginst5922 (R1375_U122, R1375_U156, R1375_U169, R1375_U45);
  and ginst5923 (R1375_U123, R1375_U156, R1375_U51);
  and ginst5924 (R1375_U124, R1375_U15, R1375_U171);
  and ginst5925 (R1375_U125, R1375_U7, U3498);
  and ginst5926 (R1375_U126, R1375_U156, R1375_U52);
  and ginst5927 (R1375_U127, R1375_U15, R1375_U167);
  and ginst5928 (R1375_U128, R1375_U8, U3494);
  and ginst5929 (R1375_U129, R1375_U156, R1375_U57);
  and ginst5930 (R1375_U13, R1375_U184, R1375_U185, R1375_U186);
  and ginst5931 (R1375_U130, R1375_U100, R1375_U15, R1375_U178, R1375_U19, U3486);
  and ginst5932 (R1375_U131, R1375_U156, R1375_U181, R1375_U59);
  and ginst5933 (R1375_U132, R1375_U15, R1375_U35);
  and ginst5934 (R1375_U133, R1375_U156, R1375_U184, R1375_U185, R1375_U37);
  and ginst5935 (R1375_U134, R1375_U217, R1375_U218);
  and ginst5936 (R1375_U135, R1375_U156, R1375_U219);
  and ginst5937 (R1375_U136, R1375_U156, R1375_U172, R1375_U49);
  and ginst5938 (R1375_U137, R1375_U15, R1375_U48);
  and ginst5939 (R1375_U138, R1375_U7, U3500);
  and ginst5940 (R1375_U139, R1375_U193, R1375_U199);
  and ginst5941 (R1375_U14, R1375_U103, R1375_U13, R1375_U152, R1375_U191);
  and ginst5942 (R1375_U140, R1375_U200, R1375_U201, R1375_U202);
  and ginst5943 (R1375_U141, R1375_U139, R1375_U140, R1375_U150, R1375_U187);
  and ginst5944 (R1375_U142, R1375_U203, R1375_U204);
  and ginst5945 (R1375_U143, R1375_U207, R1375_U208);
  and ginst5946 (R1375_U144, R1375_U142, R1375_U143, R1375_U205, R1375_U206, R1375_U209);
  and ginst5947 (R1375_U145, R1375_U210, R1375_U211);
  and ginst5948 (R1375_U146, R1375_U145, R1375_U212, R1375_U213);
  and ginst5949 (R1375_U147, R1375_U214, R1375_U215, R1375_U216);
  and ginst5950 (R1375_U148, R1375_U223, R1375_U224, R1375_U225);
  and ginst5951 (R1375_U149, R1375_U148, R1375_U220, R1375_U221, R1375_U222);
  and ginst5952 (R1375_U15, R1375_U153, R1375_U154, R1375_U155, R1375_U157);
  nand ginst5953 (R1375_U150, R1375_U15, R1375_U156, R1375_U196);
  nand ginst5954 (R1375_U151, R1375_U54, U3478);
  nand ginst5955 (R1375_U152, R1375_U151, R1375_U92);
  nand ginst5956 (R1375_U153, R1375_U66, U4038);
  nand ginst5957 (R1375_U154, R1375_U88, U3056);
  nand ginst5958 (R1375_U155, R1375_U87, U3052);
  nand ginst5959 (R1375_U156, R1375_U86, U3051);
  nand ginst5960 (R1375_U157, R1375_U85, U3050);
  nand ginst5961 (R1375_U158, R1375_U30, U3054);
  nand ginst5962 (R1375_U159, R1375_U63, U4033);
  and ginst5963 (R1375_U16, R1375_U158, R1375_U165, R1375_U168, R1375_U169, R1375_U24);
  nand ginst5964 (R1375_U160, R1375_U159, R1375_U91);
  nand ginst5965 (R1375_U161, R1375_U29, U3055);
  nand ginst5966 (R1375_U162, R1375_U41, U3062);
  nand ginst5967 (R1375_U163, R1375_U61, U4034);
  nand ginst5968 (R1375_U164, R1375_U63, U4033);
  nand ginst5969 (R1375_U165, R1375_U6, R1375_U93);
  nand ginst5970 (R1375_U166, R1375_U73, U3077);
  nand ginst5971 (R1375_U167, R1375_U69, U3071);
  nand ginst5972 (R1375_U168, R1375_U75, U3073);
  nand ginst5973 (R1375_U169, R1375_U82, U3072);
  and ginst5974 (R1375_U17, R1375_U10, R1375_U109, R1375_U179, R1375_U24);
  nand ginst5975 (R1375_U170, R1375_U49, U3502);
  nand ginst5976 (R1375_U171, R1375_U170, R1375_U95);
  nand ginst5977 (R1375_U172, R1375_U72, U3078);
  nand ginst5978 (R1375_U173, R1375_U47, U3079);
  nand ginst5979 (R1375_U174, R1375_U76, U3070);
  nand ginst5980 (R1375_U175, R1375_U77, U3076);
  nand ginst5981 (R1375_U176, R1375_U55, U3069);
  nand ginst5982 (R1375_U177, R1375_U53, U3490);
  nand ginst5983 (R1375_U178, R1375_U177, R1375_U94);
  nand ginst5984 (R1375_U179, R1375_U78, U3059);
  and ginst5985 (R1375_U18, R1375_U100, R1375_U22);
  nand ginst5986 (R1375_U180, R1375_U74, U3067);
  nand ginst5987 (R1375_U181, R1375_U68, U3080);
  nand ginst5988 (R1375_U182, R1375_U79, U3081);
  nand ginst5989 (R1375_U183, R1375_U38, U3068);
  nand ginst5990 (R1375_U184, R1375_U80, U3057);
  nand ginst5991 (R1375_U185, R1375_U71, U3061);
  nand ginst5992 (R1375_U186, R1375_U81, U3065);
  nand ginst5993 (R1375_U187, R1375_U101, R1375_U102, R1375_U156, R1375_U18);
  nand ginst5994 (R1375_U188, U3147, U3464);
  nand ginst5995 (R1375_U189, R1375_U188, U3074);
  and ginst5996 (R1375_U19, R1375_U10, R1375_U165);
  nand ginst5997 (R1375_U190, R1375_U64, U3075);
  or ginst5998 (R1375_U191, U3147, U3464);
  nand ginst5999 (R1375_U192, R1375_U83, U3058);
  nand ginst6000 (R1375_U193, R1375_U104, R1375_U105);
  nand ginst6001 (R1375_U194, R1375_U158, R1375_U90);
  nand ginst6002 (R1375_U195, R1375_U28, U4031);
  nand ginst6003 (R1375_U196, R1375_U194, R1375_U195);
  nand ginst6004 (R1375_U197, R1375_U154, R1375_U33, U4040);
  nand ginst6005 (R1375_U198, R1375_U32, U4039);
  nand ginst6006 (R1375_U199, R1375_U31, U3053);
  and ginst6007 (R1375_U20, R1375_U154, R1375_U155, R1375_U34, U4030);
  nand ginst6008 (R1375_U200, R1375_U106, R1375_U107, R1375_U25, R1375_U9, U3490);
  nand ginst6009 (R1375_U201, R1375_U100, R1375_U108, R1375_U156, R1375_U19, U3488);
  nand ginst6010 (R1375_U202, R1375_U110, R1375_U156, R1375_U17, U3484);
  nand ginst6011 (R1375_U203, R1375_U111, R1375_U112, R1375_U156, R1375_U25);
  nand ginst6012 (R1375_U204, R1375_U10, R1375_U113, R1375_U114, R1375_U23, R1375_U25);
  nand ginst6013 (R1375_U205, R1375_U115, R1375_U116);
  nand ginst6014 (R1375_U206, R1375_U117, R1375_U15, R1375_U18, U3472);
  nand ginst6015 (R1375_U207, R1375_U118, R1375_U156, R1375_U16, U3504);
  nand ginst6016 (R1375_U208, R1375_U119, R1375_U156, R1375_U25, R1375_U9, U3492);
  nand ginst6017 (R1375_U209, R1375_U120, R1375_U121, R1375_U156, R1375_U17);
  and ginst6018 (R1375_U21, R1375_U154, R1375_U155, R1375_U27, U4029);
  nand ginst6019 (R1375_U210, R1375_U122, R1375_U15, R1375_U25, U4037);
  nand ginst6020 (R1375_U211, R1375_U123, R1375_U124, R1375_U125, R1375_U16);
  nand ginst6021 (R1375_U212, R1375_U126, R1375_U127, R1375_U128, R1375_U25);
  nand ginst6022 (R1375_U213, R1375_U129, R1375_U130);
  nand ginst6023 (R1375_U214, R1375_U131, R1375_U15, R1375_U17, U3482);
  nand ginst6024 (R1375_U215, R1375_U132, R1375_U156, R1375_U18, U3474);
  nand ginst6025 (R1375_U216, R1375_U100, R1375_U133, R1375_U15, R1375_U22, U3470);
  nand ginst6026 (R1375_U217, R1375_U46, U4036);
  nand ginst6027 (R1375_U218, R1375_U42, U4035);
  nand ginst6028 (R1375_U219, R1375_U134, R1375_U6);
  and ginst6029 (R1375_U22, R1375_U10, R1375_U12, R1375_U99);
  nand ginst6030 (R1375_U220, R1375_U135, R1375_U15, R1375_U25);
  nand ginst6031 (R1375_U221, R1375_U136, R1375_U15, R1375_U16, U3502);
  nand ginst6032 (R1375_U222, R1375_U137, R1375_U138, R1375_U156, R1375_U16);
  nand ginst6033 (R1375_U223, R1375_U153, R1375_U156, R1375_U20);
  nand ginst6034 (R1375_U224, R1375_U153, R1375_U21);
  nand ginst6035 (R1375_U225, R1375_U153, R1375_U89);
  and ginst6036 (R1375_U23, R1375_U11, R1375_U178, R1375_U179, R1375_U180);
  and ginst6037 (R1375_U24, R1375_U160, R1375_U161, R1375_U162);
  and ginst6038 (R1375_U25, R1375_U100, R1375_U165);
  nand ginst6039 (R1375_U26, R1375_U141, R1375_U144, R1375_U146, R1375_U147, R1375_U149);
  not ginst6040 (R1375_U27, U3051);
  not ginst6041 (R1375_U28, U3054);
  not ginst6042 (R1375_U29, U4032);
  not ginst6043 (R1375_U30, U4031);
  not ginst6044 (R1375_U31, U4038);
  not ginst6045 (R1375_U32, U3056);
  not ginst6046 (R1375_U33, U3052);
  not ginst6047 (R1375_U34, U3050);
  not ginst6048 (R1375_U35, U3057);
  not ginst6049 (R1375_U36, U3061);
  not ginst6050 (R1375_U37, U3065);
  not ginst6051 (R1375_U38, U3478);
  not ginst6052 (R1375_U39, U3064);
  not ginst6053 (R1375_U40, U4034);
  not ginst6054 (R1375_U41, U4033);
  not ginst6055 (R1375_U42, U3058);
  not ginst6056 (R1375_U43, U3077);
  not ginst6057 (R1375_U44, U3071);
  not ginst6058 (R1375_U45, U3073);
  not ginst6059 (R1375_U46, U3072);
  not ginst6060 (R1375_U47, U3502);
  not ginst6061 (R1375_U48, U3066);
  not ginst6062 (R1375_U49, U3079);
  not ginst6063 (R1375_U50, U3078);
  not ginst6064 (R1375_U51, U3070);
  not ginst6065 (R1375_U52, U3076);
  not ginst6066 (R1375_U53, U3069);
  not ginst6067 (R1375_U54, U3068);
  not ginst6068 (R1375_U55, U3490);
  not ginst6069 (R1375_U56, U3060);
  not ginst6070 (R1375_U57, U3059);
  not ginst6071 (R1375_U58, U3067);
  not ginst6072 (R1375_U59, U3081);
  and ginst6073 (R1375_U6, R1375_U163, R1375_U164);
  not ginst6074 (R1375_U60, U3080);
  not ginst6075 (R1375_U61, U3063);
  not ginst6076 (R1375_U62, U3055);
  not ginst6077 (R1375_U63, U3062);
  not ginst6078 (R1375_U64, U3468);
  not ginst6079 (R1375_U65, U3075);
  not ginst6080 (R1375_U66, U3053);
  not ginst6081 (R1375_U67, U3488);
  not ginst6082 (R1375_U68, U3484);
  not ginst6083 (R1375_U69, U3496);
  and ginst6084 (R1375_U7, R1375_U172, R1375_U173);
  not ginst6085 (R1375_U70, U3476);
  not ginst6086 (R1375_U71, U3472);
  not ginst6087 (R1375_U72, U3504);
  not ginst6088 (R1375_U73, U3492);
  not ginst6089 (R1375_U74, U3480);
  not ginst6090 (R1375_U75, U4037);
  not ginst6091 (R1375_U76, U3498);
  not ginst6092 (R1375_U77, U3494);
  not ginst6093 (R1375_U78, U3486);
  not ginst6094 (R1375_U79, U3482);
  and ginst6095 (R1375_U8, R1375_U171, R1375_U174, R1375_U7, R1375_U96);
  not ginst6096 (R1375_U80, U3474);
  not ginst6097 (R1375_U81, U3470);
  not ginst6098 (R1375_U82, U4036);
  not ginst6099 (R1375_U83, U4035);
  not ginst6100 (R1375_U84, U3500);
  not ginst6101 (R1375_U85, U4030);
  not ginst6102 (R1375_U86, U4029);
  not ginst6103 (R1375_U87, U4040);
  not ginst6104 (R1375_U88, U4039);
  nand ginst6105 (R1375_U89, R1375_U197, R1375_U198);
  and ginst6106 (R1375_U9, R1375_U8, R1375_U97);
  and ginst6107 (R1375_U90, R1375_U62, U4032);
  and ginst6108 (R1375_U91, R1375_U40, U3063);
  and ginst6109 (R1375_U92, R1375_U70, U3064);
  and ginst6110 (R1375_U93, R1375_U83, U3058);
  and ginst6111 (R1375_U94, R1375_U67, U3060);
  and ginst6112 (R1375_U95, R1375_U84, U3066);
  and ginst6113 (R1375_U96, R1375_U168, R1375_U169);
  and ginst6114 (R1375_U97, R1375_U167, R1375_U175);
  and ginst6115 (R1375_U98, R1375_U166, R1375_U176);
  and ginst6116 (R1375_U99, R1375_U152, R1375_U165);
  not ginst6117 (R395_U10, U3143);
  not ginst6118 (R395_U100, U3144);
  not ginst6119 (R395_U101, U3145);
  nand ginst6120 (R395_U102, R395_U100, R395_U101, U3113);
  nand ginst6121 (R395_U103, R395_U100, U3112);
  nand ginst6122 (R395_U104, R395_U10, U3111);
  nand ginst6123 (R395_U105, R395_U67, R395_U68);
  nand ginst6124 (R395_U106, R395_U108, R395_U109, R395_U7, U3143);
  nand ginst6125 (R395_U107, R395_U109, R395_U69);
  nand ginst6126 (R395_U108, R395_U11, U3110);
  nand ginst6127 (R395_U109, R395_U12, U3109);
  not ginst6128 (R395_U11, U3142);
  nand ginst6129 (R395_U110, R395_U9, U3141);
  nand ginst6130 (R395_U111, R395_U16, U3140);
  nand ginst6131 (R395_U112, R395_U105, R395_U70, R395_U71);
  nand ginst6132 (R395_U113, R395_U115, R395_U116, R395_U13, U3108);
  nand ginst6133 (R395_U114, R395_U116, R395_U72);
  nand ginst6134 (R395_U115, R395_U17, U3139);
  nand ginst6135 (R395_U116, R395_U18, U3138);
  nand ginst6136 (R395_U117, R395_U15, U3106);
  nand ginst6137 (R395_U118, R395_U22, U3105);
  nand ginst6138 (R395_U119, R395_U112, R395_U73);
  not ginst6139 (R395_U12, U3141);
  nand ginst6140 (R395_U120, R395_U122, R395_U123, R395_U19, U3137);
  nand ginst6141 (R395_U121, R395_U123, R395_U75);
  nand ginst6142 (R395_U122, R395_U23, U3104);
  nand ginst6143 (R395_U123, R395_U24, U3103);
  nand ginst6144 (R395_U124, R395_U21, U3135);
  nand ginst6145 (R395_U125, R395_U28, U3134);
  nand ginst6146 (R395_U126, R395_U119, R395_U76);
  nand ginst6147 (R395_U127, R395_U129, R395_U130, R395_U25, U3102);
  nand ginst6148 (R395_U128, R395_U130, R395_U78);
  nand ginst6149 (R395_U129, R395_U29, U3133);
  not ginst6150 (R395_U13, U3140);
  nand ginst6151 (R395_U130, R395_U30, U3132);
  nand ginst6152 (R395_U131, R395_U27, U3100);
  nand ginst6153 (R395_U132, R395_U32, U3099);
  nand ginst6154 (R395_U133, R395_U126, R395_U79);
  nand ginst6155 (R395_U134, R395_U31, U3131);
  nand ginst6156 (R395_U135, R395_U34, U3130);
  nand ginst6157 (R395_U136, R395_U133, R395_U81);
  nand ginst6158 (R395_U137, R395_U33, U3098);
  nand ginst6159 (R395_U138, R395_U36, U3097);
  nand ginst6160 (R395_U139, R395_U136, R395_U82);
  not ginst6161 (R395_U14, U3139);
  nand ginst6162 (R395_U140, R395_U35, U3129);
  nand ginst6163 (R395_U141, R395_U38, U3128);
  nand ginst6164 (R395_U142, R395_U139, R395_U83);
  nand ginst6165 (R395_U143, R395_U37, U3096);
  nand ginst6166 (R395_U144, R395_U40, U3095);
  nand ginst6167 (R395_U145, R395_U142, R395_U84);
  nand ginst6168 (R395_U146, R395_U39, U3127);
  nand ginst6169 (R395_U147, R395_U42, U3126);
  nand ginst6170 (R395_U148, R395_U145, R395_U85);
  nand ginst6171 (R395_U149, R395_U41, U3094);
  not ginst6172 (R395_U15, U3138);
  nand ginst6173 (R395_U150, R395_U44, U3093);
  nand ginst6174 (R395_U151, R395_U148, R395_U86);
  nand ginst6175 (R395_U152, R395_U43, U3125);
  nand ginst6176 (R395_U153, R395_U46, U3124);
  nand ginst6177 (R395_U154, R395_U151, R395_U87);
  nand ginst6178 (R395_U155, R395_U45, U3092);
  nand ginst6179 (R395_U156, R395_U48, U3091);
  nand ginst6180 (R395_U157, R395_U154, R395_U88);
  nand ginst6181 (R395_U158, R395_U47, U3123);
  nand ginst6182 (R395_U159, R395_U50, U3122);
  not ginst6183 (R395_U16, U3108);
  nand ginst6184 (R395_U160, R395_U157, R395_U89);
  nand ginst6185 (R395_U161, R395_U49, U3090);
  nand ginst6186 (R395_U162, R395_U52, U3089);
  nand ginst6187 (R395_U163, R395_U160, R395_U90);
  nand ginst6188 (R395_U164, R395_U51, U3121);
  nand ginst6189 (R395_U165, R395_U54, U3120);
  nand ginst6190 (R395_U166, R395_U163, R395_U91);
  nand ginst6191 (R395_U167, R395_U53, U3088);
  nand ginst6192 (R395_U168, R395_U56, U3087);
  nand ginst6193 (R395_U169, R395_U166, R395_U92);
  not ginst6194 (R395_U17, U3107);
  nand ginst6195 (R395_U170, R395_U55, U3119);
  nand ginst6196 (R395_U171, R395_U58, U3118);
  nand ginst6197 (R395_U172, R395_U169, R395_U93);
  nand ginst6198 (R395_U173, R395_U57, U3086);
  nand ginst6199 (R395_U174, R395_U60, U3085);
  nand ginst6200 (R395_U175, R395_U172, R395_U94);
  nand ginst6201 (R395_U176, R395_U59, U3117);
  nand ginst6202 (R395_U177, R395_U62, U3116);
  nand ginst6203 (R395_U178, R395_U175, R395_U95);
  nand ginst6204 (R395_U179, R395_U61, U3084);
  not ginst6205 (R395_U18, U3106);
  nand ginst6206 (R395_U180, R395_U64, U3083);
  nand ginst6207 (R395_U181, R395_U178, R395_U96);
  nand ginst6208 (R395_U182, R395_U63, U3115);
  nand ginst6209 (R395_U183, R395_U181, R395_U97);
  nand ginst6210 (R395_U184, R395_U101, U3112, U3113);
  nand ginst6211 (R395_U185, R395_U98, U3114);
  nand ginst6212 (R395_U186, R395_U65, U3082);
  nand ginst6213 (R395_U187, R395_U98, U3114, U3146);
  nand ginst6214 (R395_U188, R395_U65, R395_U66, U3082);
  not ginst6215 (R395_U19, U3105);
  not ginst6216 (R395_U20, U3104);
  not ginst6217 (R395_U21, U3103);
  not ginst6218 (R395_U22, U3137);
  not ginst6219 (R395_U23, U3136);
  not ginst6220 (R395_U24, U3135);
  not ginst6221 (R395_U25, U3134);
  not ginst6222 (R395_U26, U3133);
  not ginst6223 (R395_U27, U3132);
  not ginst6224 (R395_U28, U3102);
  not ginst6225 (R395_U29, U3101);
  not ginst6226 (R395_U30, U3100);
  not ginst6227 (R395_U31, U3099);
  not ginst6228 (R395_U32, U3131);
  not ginst6229 (R395_U33, U3130);
  not ginst6230 (R395_U34, U3098);
  not ginst6231 (R395_U35, U3097);
  not ginst6232 (R395_U36, U3129);
  not ginst6233 (R395_U37, U3128);
  not ginst6234 (R395_U38, U3096);
  not ginst6235 (R395_U39, U3095);
  not ginst6236 (R395_U40, U3127);
  not ginst6237 (R395_U41, U3126);
  not ginst6238 (R395_U42, U3094);
  not ginst6239 (R395_U43, U3093);
  not ginst6240 (R395_U44, U3125);
  not ginst6241 (R395_U45, U3124);
  not ginst6242 (R395_U46, U3092);
  not ginst6243 (R395_U47, U3091);
  not ginst6244 (R395_U48, U3123);
  not ginst6245 (R395_U49, U3122);
  not ginst6246 (R395_U50, U3090);
  not ginst6247 (R395_U51, U3089);
  not ginst6248 (R395_U52, U3121);
  not ginst6249 (R395_U53, U3120);
  not ginst6250 (R395_U54, U3088);
  not ginst6251 (R395_U55, U3087);
  not ginst6252 (R395_U56, U3119);
  not ginst6253 (R395_U57, U3118);
  not ginst6254 (R395_U58, U3086);
  not ginst6255 (R395_U59, U3085);
  nand ginst6256 (R395_U6, R395_U183, R395_U99);
  not ginst6257 (R395_U60, U3117);
  not ginst6258 (R395_U61, U3116);
  not ginst6259 (R395_U62, U3084);
  not ginst6260 (R395_U63, U3083);
  not ginst6261 (R395_U64, U3115);
  not ginst6262 (R395_U65, U3114);
  not ginst6263 (R395_U66, U3146);
  and ginst6264 (R395_U67, R395_U102, R395_U103, R395_U104);
  and ginst6265 (R395_U68, R395_U108, R395_U109, R395_U184);
  and ginst6266 (R395_U69, R395_U8, U3142);
  not ginst6267 (R395_U7, U3111);
  and ginst6268 (R395_U70, R395_U106, R395_U107, R395_U110);
  and ginst6269 (R395_U71, R395_U111, R395_U115, R395_U116);
  and ginst6270 (R395_U72, R395_U14, U3107);
  and ginst6271 (R395_U73, R395_U113, R395_U114, R395_U117, R395_U74);
  and ginst6272 (R395_U74, R395_U118, R395_U122, R395_U123);
  and ginst6273 (R395_U75, R395_U20, U3136);
  and ginst6274 (R395_U76, R395_U120, R395_U121, R395_U124, R395_U77);
  and ginst6275 (R395_U77, R395_U125, R395_U129, R395_U130);
  and ginst6276 (R395_U78, R395_U26, U3101);
  and ginst6277 (R395_U79, R395_U127, R395_U128, R395_U80);
  not ginst6278 (R395_U8, U3110);
  and ginst6279 (R395_U80, R395_U131, R395_U132);
  and ginst6280 (R395_U81, R395_U134, R395_U135);
  and ginst6281 (R395_U82, R395_U137, R395_U138);
  and ginst6282 (R395_U83, R395_U140, R395_U141);
  and ginst6283 (R395_U84, R395_U143, R395_U144);
  and ginst6284 (R395_U85, R395_U146, R395_U147);
  and ginst6285 (R395_U86, R395_U149, R395_U150);
  and ginst6286 (R395_U87, R395_U152, R395_U153);
  and ginst6287 (R395_U88, R395_U155, R395_U156);
  and ginst6288 (R395_U89, R395_U158, R395_U159);
  not ginst6289 (R395_U9, U3109);
  and ginst6290 (R395_U90, R395_U161, R395_U162);
  and ginst6291 (R395_U91, R395_U164, R395_U165);
  and ginst6292 (R395_U92, R395_U167, R395_U168);
  and ginst6293 (R395_U93, R395_U170, R395_U171);
  and ginst6294 (R395_U94, R395_U173, R395_U174);
  and ginst6295 (R395_U95, R395_U176, R395_U177);
  and ginst6296 (R395_U96, R395_U179, R395_U180);
  and ginst6297 (R395_U97, R395_U182, R395_U185, R395_U186);
  not ginst6298 (R395_U98, U3082);
  and ginst6299 (R395_U99, R395_U187, R395_U188);
  and ginst6300 (SUB_84_U10, SUB_84_U133, SUB_84_U43);
  nand ginst6301 (SUB_84_U100, SUB_84_U69, SUB_84_U91);
  nand ginst6302 (SUB_84_U101, IR_REG_5__SCAN_IN, SUB_84_U100);
  nand ginst6303 (SUB_84_U102, IR_REG_3__SCAN_IN, SUB_84_U29);
  nand ginst6304 (SUB_84_U103, SUB_84_U47, SUB_84_U95);
  not ginst6305 (SUB_84_U104, SUB_84_U46);
  not ginst6306 (SUB_84_U105, SUB_84_U32);
  nand ginst6307 (SUB_84_U106, SUB_84_U105, SUB_84_U44);
  not ginst6308 (SUB_84_U107, SUB_84_U43);
  not ginst6309 (SUB_84_U108, SUB_84_U34);
  nand ginst6310 (SUB_84_U109, SUB_84_U105, SUB_84_U35, SUB_84_U4, SUB_84_U5);
  and ginst6311 (SUB_84_U11, SUB_84_U132, SUB_84_U38);
  not ginst6312 (SUB_84_U110, SUB_84_U33);
  or ginst6313 (SUB_84_U111, IR_REG_0__SCAN_IN, IR_REG_1__SCAN_IN);
  nand ginst6314 (SUB_84_U112, IR_REG_2__SCAN_IN, SUB_84_U111);
  nand ginst6315 (SUB_84_U113, IR_REG_29__SCAN_IN, SUB_84_U109);
  nand ginst6316 (SUB_84_U114, SUB_84_U108, SUB_84_U4);
  nand ginst6317 (SUB_84_U115, IR_REG_28__SCAN_IN, SUB_84_U114);
  not ginst6318 (SUB_84_U116, SUB_84_U36);
  not ginst6319 (SUB_84_U117, SUB_84_U75);
  nand ginst6320 (SUB_84_U118, IR_REG_26__SCAN_IN, SUB_84_U36);
  nand ginst6321 (SUB_84_U119, SUB_84_U108, SUB_84_U77);
  and ginst6322 (SUB_84_U12, SUB_84_U122, SUB_84_U130);
  nand ginst6323 (SUB_84_U120, IR_REG_25__SCAN_IN, SUB_84_U119);
  not ginst6324 (SUB_84_U121, SUB_84_U38);
  nand ginst6325 (SUB_84_U122, SUB_84_U121, SUB_84_U42);
  not ginst6326 (SUB_84_U123, SUB_84_U39);
  not ginst6327 (SUB_84_U124, SUB_84_U40);
  not ginst6328 (SUB_84_U125, SUB_84_U80);
  nand ginst6329 (SUB_84_U126, IR_REG_22__SCAN_IN, SUB_84_U40);
  nand ginst6330 (SUB_84_U127, SUB_84_U123, SUB_84_U82);
  nand ginst6331 (SUB_84_U128, IR_REG_21__SCAN_IN, SUB_84_U127);
  nand ginst6332 (SUB_84_U129, IR_REG_19__SCAN_IN, SUB_84_U122);
  and ginst6333 (SUB_84_U13, SUB_84_U129, SUB_84_U39);
  nand ginst6334 (SUB_84_U130, IR_REG_18__SCAN_IN, SUB_84_U38);
  nand ginst6335 (SUB_84_U131, SUB_84_U107, SUB_84_U86);
  nand ginst6336 (SUB_84_U132, IR_REG_17__SCAN_IN, SUB_84_U131);
  nand ginst6337 (SUB_84_U133, IR_REG_15__SCAN_IN, SUB_84_U106);
  nand ginst6338 (SUB_84_U134, IR_REG_14__SCAN_IN, SUB_84_U32);
  nand ginst6339 (SUB_84_U135, SUB_84_U104, SUB_84_U88);
  nand ginst6340 (SUB_84_U136, IR_REG_13__SCAN_IN, SUB_84_U135);
  nand ginst6341 (SUB_84_U137, IR_REG_11__SCAN_IN, SUB_84_U103);
  nand ginst6342 (SUB_84_U138, IR_REG_10__SCAN_IN, SUB_84_U45);
  nand ginst6343 (SUB_84_U139, SUB_84_U110, SUB_84_U72);
  and ginst6344 (SUB_84_U14, SUB_84_U128, SUB_84_U40);
  nand ginst6345 (SUB_84_U140, IR_REG_8__SCAN_IN, SUB_84_U27);
  nand ginst6346 (SUB_84_U141, SUB_84_U67, SUB_84_U94);
  nand ginst6347 (SUB_84_U142, IR_REG_4__SCAN_IN, SUB_84_U30);
  nand ginst6348 (SUB_84_U143, SUB_84_U69, SUB_84_U91);
  nand ginst6349 (SUB_84_U144, SUB_84_U139, SUB_84_U71);
  nand ginst6350 (SUB_84_U145, IR_REG_31__SCAN_IN, SUB_84_U110, SUB_84_U72);
  nand ginst6351 (SUB_84_U146, IR_REG_30__SCAN_IN, SUB_84_U33);
  nand ginst6352 (SUB_84_U147, SUB_84_U110, SUB_84_U72);
  nand ginst6353 (SUB_84_U148, IR_REG_27__SCAN_IN, SUB_84_U75);
  nand ginst6354 (SUB_84_U149, SUB_84_U117, SUB_84_U74);
  and ginst6355 (SUB_84_U15, SUB_84_U126, SUB_84_U80);
  nand ginst6356 (SUB_84_U150, IR_REG_24__SCAN_IN, SUB_84_U34);
  nand ginst6357 (SUB_84_U151, SUB_84_U108, SUB_84_U77);
  nand ginst6358 (SUB_84_U152, IR_REG_23__SCAN_IN, SUB_84_U80);
  nand ginst6359 (SUB_84_U153, SUB_84_U125, SUB_84_U79);
  nand ginst6360 (SUB_84_U154, IR_REG_20__SCAN_IN, SUB_84_U39);
  nand ginst6361 (SUB_84_U155, SUB_84_U123, SUB_84_U82);
  nand ginst6362 (SUB_84_U156, IR_REG_1__SCAN_IN, SUB_84_U85);
  nand ginst6363 (SUB_84_U157, IR_REG_0__SCAN_IN, SUB_84_U84);
  nand ginst6364 (SUB_84_U158, IR_REG_16__SCAN_IN, SUB_84_U43);
  nand ginst6365 (SUB_84_U159, SUB_84_U107, SUB_84_U86);
  and ginst6366 (SUB_84_U16, SUB_84_U120, SUB_84_U36);
  nand ginst6367 (SUB_84_U160, IR_REG_12__SCAN_IN, SUB_84_U46);
  nand ginst6368 (SUB_84_U161, SUB_84_U104, SUB_84_U88);
  and ginst6369 (SUB_84_U17, SUB_84_U118, SUB_84_U75);
  and ginst6370 (SUB_84_U18, SUB_84_U109, SUB_84_U115);
  and ginst6371 (SUB_84_U19, SUB_84_U113, SUB_84_U33);
  and ginst6372 (SUB_84_U20, SUB_84_U112, SUB_84_U29);
  and ginst6373 (SUB_84_U21, SUB_84_U102, SUB_84_U30);
  and ginst6374 (SUB_84_U22, SUB_84_U101, SUB_84_U26);
  and ginst6375 (SUB_84_U23, SUB_84_U93, SUB_84_U99);
  and ginst6376 (SUB_84_U24, SUB_84_U27, SUB_84_U98);
  and ginst6377 (SUB_84_U25, SUB_84_U45, SUB_84_U97);
  nand ginst6378 (SUB_84_U26, SUB_84_U50, SUB_84_U51);
  nand ginst6379 (SUB_84_U27, SUB_84_U53, SUB_84_U92);
  not ginst6380 (SUB_84_U28, IR_REG_6__SCAN_IN);
  or ginst6381 (SUB_84_U29, IR_REG_0__SCAN_IN, IR_REG_1__SCAN_IN, IR_REG_2__SCAN_IN);
  nand ginst6382 (SUB_84_U30, SUB_84_U31, SUB_84_U90);
  not ginst6383 (SUB_84_U31, IR_REG_3__SCAN_IN);
  nand ginst6384 (SUB_84_U32, SUB_84_U56, SUB_84_U57, SUB_84_U58, SUB_84_U59);
  nand ginst6385 (SUB_84_U33, SUB_84_U105, SUB_84_U4, SUB_84_U5, SUB_84_U60);
  nand ginst6386 (SUB_84_U34, SUB_84_U105, SUB_84_U5);
  not ginst6387 (SUB_84_U35, IR_REG_28__SCAN_IN);
  nand ginst6388 (SUB_84_U36, SUB_84_U108, SUB_84_U61);
  not ginst6389 (SUB_84_U37, IR_REG_26__SCAN_IN);
  nand ginst6390 (SUB_84_U38, SUB_84_U105, SUB_84_U62);
  nand ginst6391 (SUB_84_U39, SUB_84_U121, SUB_84_U63);
  nor ginst6392 (SUB_84_U4, IR_REG_24__SCAN_IN, IR_REG_25__SCAN_IN, IR_REG_26__SCAN_IN, IR_REG_27__SCAN_IN);
  nand ginst6393 (SUB_84_U40, SUB_84_U123, SUB_84_U64);
  not ginst6394 (SUB_84_U41, IR_REG_22__SCAN_IN);
  not ginst6395 (SUB_84_U42, IR_REG_18__SCAN_IN);
  nand ginst6396 (SUB_84_U43, SUB_84_U105, SUB_84_U65);
  not ginst6397 (SUB_84_U44, IR_REG_14__SCAN_IN);
  nand ginst6398 (SUB_84_U45, SUB_84_U52, SUB_84_U92);
  nand ginst6399 (SUB_84_U46, SUB_84_U66, SUB_84_U95);
  not ginst6400 (SUB_84_U47, IR_REG_10__SCAN_IN);
  nand ginst6401 (SUB_84_U48, SUB_84_U156, SUB_84_U157);
  nand ginst6402 (SUB_84_U49, SUB_84_U144, SUB_84_U145);
  and ginst6403 (SUB_84_U5, SUB_84_U54, SUB_84_U55);
  nor ginst6404 (SUB_84_U50, IR_REG_0__SCAN_IN, IR_REG_1__SCAN_IN, IR_REG_2__SCAN_IN);
  nor ginst6405 (SUB_84_U51, IR_REG_3__SCAN_IN, IR_REG_4__SCAN_IN, IR_REG_5__SCAN_IN);
  nor ginst6406 (SUB_84_U52, IR_REG_6__SCAN_IN, IR_REG_7__SCAN_IN, IR_REG_8__SCAN_IN, IR_REG_9__SCAN_IN);
  nor ginst6407 (SUB_84_U53, IR_REG_6__SCAN_IN, IR_REG_7__SCAN_IN);
  nor ginst6408 (SUB_84_U54, IR_REG_14__SCAN_IN, IR_REG_15__SCAN_IN, IR_REG_16__SCAN_IN, IR_REG_17__SCAN_IN, IR_REG_18__SCAN_IN);
  nor ginst6409 (SUB_84_U55, IR_REG_19__SCAN_IN, IR_REG_20__SCAN_IN, IR_REG_21__SCAN_IN, IR_REG_22__SCAN_IN, IR_REG_23__SCAN_IN);
  nor ginst6410 (SUB_84_U56, IR_REG_10__SCAN_IN, IR_REG_11__SCAN_IN, IR_REG_12__SCAN_IN, IR_REG_13__SCAN_IN);
  nor ginst6411 (SUB_84_U57, IR_REG_0__SCAN_IN, IR_REG_1__SCAN_IN, IR_REG_2__SCAN_IN);
  nor ginst6412 (SUB_84_U58, IR_REG_3__SCAN_IN, IR_REG_4__SCAN_IN, IR_REG_5__SCAN_IN, IR_REG_6__SCAN_IN);
  nor ginst6413 (SUB_84_U59, IR_REG_7__SCAN_IN, IR_REG_8__SCAN_IN, IR_REG_9__SCAN_IN);
  and ginst6414 (SUB_84_U6, SUB_84_U103, SUB_84_U138);
  nor ginst6415 (SUB_84_U60, IR_REG_28__SCAN_IN, IR_REG_29__SCAN_IN);
  nor ginst6416 (SUB_84_U61, IR_REG_24__SCAN_IN, IR_REG_25__SCAN_IN);
  nor ginst6417 (SUB_84_U62, IR_REG_14__SCAN_IN, IR_REG_15__SCAN_IN, IR_REG_16__SCAN_IN, IR_REG_17__SCAN_IN);
  nor ginst6418 (SUB_84_U63, IR_REG_18__SCAN_IN, IR_REG_19__SCAN_IN);
  nor ginst6419 (SUB_84_U64, IR_REG_20__SCAN_IN, IR_REG_21__SCAN_IN);
  nor ginst6420 (SUB_84_U65, IR_REG_14__SCAN_IN, IR_REG_15__SCAN_IN);
  nor ginst6421 (SUB_84_U66, IR_REG_10__SCAN_IN, IR_REG_11__SCAN_IN);
  not ginst6422 (SUB_84_U67, IR_REG_8__SCAN_IN);
  and ginst6423 (SUB_84_U68, SUB_84_U140, SUB_84_U141);
  not ginst6424 (SUB_84_U69, IR_REG_4__SCAN_IN);
  and ginst6425 (SUB_84_U7, SUB_84_U137, SUB_84_U46);
  and ginst6426 (SUB_84_U70, SUB_84_U142, SUB_84_U143);
  not ginst6427 (SUB_84_U71, IR_REG_31__SCAN_IN);
  not ginst6428 (SUB_84_U72, IR_REG_30__SCAN_IN);
  and ginst6429 (SUB_84_U73, SUB_84_U146, SUB_84_U147);
  not ginst6430 (SUB_84_U74, IR_REG_27__SCAN_IN);
  nand ginst6431 (SUB_84_U75, SUB_84_U116, SUB_84_U37);
  and ginst6432 (SUB_84_U76, SUB_84_U148, SUB_84_U149);
  not ginst6433 (SUB_84_U77, IR_REG_24__SCAN_IN);
  and ginst6434 (SUB_84_U78, SUB_84_U150, SUB_84_U151);
  not ginst6435 (SUB_84_U79, IR_REG_23__SCAN_IN);
  and ginst6436 (SUB_84_U8, SUB_84_U136, SUB_84_U32);
  nand ginst6437 (SUB_84_U80, SUB_84_U124, SUB_84_U41);
  and ginst6438 (SUB_84_U81, SUB_84_U152, SUB_84_U153);
  not ginst6439 (SUB_84_U82, IR_REG_20__SCAN_IN);
  and ginst6440 (SUB_84_U83, SUB_84_U154, SUB_84_U155);
  not ginst6441 (SUB_84_U84, IR_REG_1__SCAN_IN);
  not ginst6442 (SUB_84_U85, IR_REG_0__SCAN_IN);
  not ginst6443 (SUB_84_U86, IR_REG_16__SCAN_IN);
  and ginst6444 (SUB_84_U87, SUB_84_U158, SUB_84_U159);
  not ginst6445 (SUB_84_U88, IR_REG_12__SCAN_IN);
  and ginst6446 (SUB_84_U89, SUB_84_U160, SUB_84_U161);
  and ginst6447 (SUB_84_U9, SUB_84_U106, SUB_84_U134);
  not ginst6448 (SUB_84_U90, SUB_84_U29);
  not ginst6449 (SUB_84_U91, SUB_84_U30);
  not ginst6450 (SUB_84_U92, SUB_84_U26);
  nand ginst6451 (SUB_84_U93, SUB_84_U28, SUB_84_U92);
  not ginst6452 (SUB_84_U94, SUB_84_U27);
  not ginst6453 (SUB_84_U95, SUB_84_U45);
  nand ginst6454 (SUB_84_U96, SUB_84_U67, SUB_84_U94);
  nand ginst6455 (SUB_84_U97, IR_REG_9__SCAN_IN, SUB_84_U96);
  nand ginst6456 (SUB_84_U98, IR_REG_7__SCAN_IN, SUB_84_U93);
  nand ginst6457 (SUB_84_U99, IR_REG_6__SCAN_IN, SUB_84_U26);
  and ginst6458 (U3014, U3431, U4201);
  and ginst6459 (U3015, U3456, U4011);
  and ginst6460 (U3016, U3454, U3455);
  and ginst6461 (U3017, U3654, U3659);
  and ginst6462 (U3018, U3462, U3463);
  and ginst6463 (U3019, U3462, U5826);
  and ginst6464 (U3020, U3463, U5823);
  and ginst6465 (U3021, U5823, U5826);
  and ginst6466 (U3022, U3355, U5613);
  and ginst6467 (U3023, STATE_REG_SCAN_IN, U3047);
  and ginst6468 (U3024, U5805, U5808, U5820);
  and ginst6469 (U3025, U3421, U3845);
  and ginst6470 (U3026, U4042, U5799);
  and ginst6471 (U3027, U4010, U5820);
  and ginst6472 (U3028, U3908, U4028);
  and ginst6473 (U3029, STATE_REG_SCAN_IN, U3357);
  and ginst6474 (U3030, U4019, U4044);
  and ginst6475 (U3031, U4021, U4044);
  and ginst6476 (U3032, U4012, U4044);
  and ginst6477 (U3033, U4020, U4044);
  and ginst6478 (U3034, U3454, U4042);
  and ginst6479 (U3035, U4028, U5799);
  and ginst6480 (U3036, U3026, U4044);
  and ginst6481 (U3037, U3454, U4028);
  and ginst6482 (U3038, U4938, U5802);
  and ginst6483 (U3039, U3025, U5802);
  and ginst6484 (U3040, U4938, U5799);
  and ginst6485 (U3041, U3025, U5799);
  and ginst6486 (U3042, U3016, U4938);
  and ginst6487 (U3043, U3016, U3025);
  and ginst6488 (U3044, U3023, U3421);
  and ginst6489 (U3045, STATE_REG_SCAN_IN, U5170);
  and ginst6490 (U3046, U3023, U5172);
  and ginst6491 (U3047, U3355, U5748);
  and ginst6492 (U3048, U3017, U3660);
  and ginst6493 (U3049, U4758, U4759, U4762, U4765, U4766);
  nand ginst6494 (U3050, U4695, U4696, U4697, U4698);
  nand ginst6495 (U3051, U4714, U4715, U4716, U4717);
  nand ginst6496 (U3052, U4733, U4734, U4735, U4736);
  nand ginst6497 (U3053, U4772, U4773, U4774);
  nand ginst6498 (U3054, U4676, U4677, U4678, U4679);
  nand ginst6499 (U3055, U4657, U4658, U4659, U4660);
  nand ginst6500 (U3056, U4752, U4753, U4754);
  nand ginst6501 (U3057, U4258, U4259, U4260, U4261);
  nand ginst6502 (U3058, U4600, U4601, U4602, U4603);
  nand ginst6503 (U3059, U4372, U4373, U4374, U4375);
  nand ginst6504 (U3060, U4391, U4392, U4393, U4394);
  nand ginst6505 (U3061, U4239, U4240, U4241, U4242);
  nand ginst6506 (U3062, U4638, U4639, U4640, U4641);
  nand ginst6507 (U3063, U4619, U4620, U4621, U4622);
  nand ginst6508 (U3064, U4277, U4278, U4279, U4280);
  nand ginst6509 (U3065, U4215, U4216, U4217, U4218);
  nand ginst6510 (U3066, U4505, U4506, U4507, U4508);
  nand ginst6511 (U3067, U4315, U4316, U4317, U4318);
  nand ginst6512 (U3068, U4296, U4297, U4298, U4299);
  nand ginst6513 (U3069, U4410, U4411, U4412, U4413);
  nand ginst6514 (U3070, U4486, U4487, U4488, U4489);
  nand ginst6515 (U3071, U4467, U4468, U4469, U4470);
  nand ginst6516 (U3072, U4581, U4582, U4583, U4584);
  nand ginst6517 (U3073, U4562, U4563, U4564, U4565);
  nand ginst6518 (U3074, U4220, U4221, U4222, U4223);
  nand ginst6519 (U3075, U4196, U4197, U4198, U4199);
  nand ginst6520 (U3076, U4448, U4449, U4450, U4451);
  nand ginst6521 (U3077, U4429, U4430, U4431, U4432);
  nand ginst6522 (U3078, U4543, U4544, U4545, U4546);
  nand ginst6523 (U3079, U4524, U4525, U4526, U4527);
  nand ginst6524 (U3080, U4353, U4354, U4355, U4356);
  nand ginst6525 (U3081, U4334, U4335, U4336, U4337);
  nand ginst6526 (U3082, U5537, U5538);
  nand ginst6527 (U3083, U5539, U5540);
  nand ginst6528 (U3084, U5544, U5545, U5546);
  nand ginst6529 (U3085, U5547, U5548, U5549);
  nand ginst6530 (U3086, U5550, U5551, U5552);
  nand ginst6531 (U3087, U5553, U5554, U5555);
  nand ginst6532 (U3088, U5556, U5557, U5558);
  nand ginst6533 (U3089, U5559, U5560, U5561);
  nand ginst6534 (U3090, U5562, U5563, U5564);
  nand ginst6535 (U3091, U5565, U5566, U5567);
  nand ginst6536 (U3092, U5568, U5569, U5570);
  nand ginst6537 (U3093, U5571, U5572, U5573);
  nand ginst6538 (U3094, U5577, U5578, U5579);
  nand ginst6539 (U3095, U5580, U5581, U5582);
  nand ginst6540 (U3096, U5583, U5584, U5585);
  nand ginst6541 (U3097, U5586, U5587, U5588);
  nand ginst6542 (U3098, U5589, U5590, U5591);
  nand ginst6543 (U3099, U5592, U5593, U5594);
  nand ginst6544 (U3100, U5595, U5596, U5597);
  nand ginst6545 (U3101, U5598, U5599, U5600);
  nand ginst6546 (U3102, U5601, U5602, U5603);
  nand ginst6547 (U3103, U5604, U5605, U5606);
  nand ginst6548 (U3104, U5519, U5520, U5521);
  nand ginst6549 (U3105, U5522, U5523, U5524);
  nand ginst6550 (U3106, U5525, U5526, U5527);
  nand ginst6551 (U3107, U5528, U5529, U5530);
  nand ginst6552 (U3108, U5531, U5532, U5533);
  nand ginst6553 (U3109, U5534, U5535, U5536);
  nand ginst6554 (U3110, U5541, U5542, U5543);
  nand ginst6555 (U3111, U5574, U5575, U5576);
  nand ginst6556 (U3112, U5607, U5608, U5609);
  nand ginst6557 (U3113, U5610, U5611);
  nand ginst6558 (U3114, U3926, U5441);
  nand ginst6559 (U3115, U3927, U5444);
  nand ginst6560 (U3116, U3929, U5450);
  nand ginst6561 (U3117, U3931, U5453);
  nand ginst6562 (U3118, U3933, U5456);
  nand ginst6563 (U3119, U3935, U5459);
  nand ginst6564 (U3120, U3937, U5462);
  nand ginst6565 (U3121, U3939, U5465);
  nand ginst6566 (U3122, U3941, U5468);
  nand ginst6567 (U3123, U3943, U5471);
  nand ginst6568 (U3124, U3945, U5474);
  nand ginst6569 (U3125, U3947, U5477);
  nand ginst6570 (U3126, U3950, U5484);
  nand ginst6571 (U3127, U3951, U5487);
  nand ginst6572 (U3128, U3952, U5490);
  nand ginst6573 (U3129, U3953, U5493);
  nand ginst6574 (U3130, U3954, U5496);
  nand ginst6575 (U3131, U3955, U5499);
  nand ginst6576 (U3132, U3956, U5502);
  nand ginst6577 (U3133, U3957, U5505);
  nand ginst6578 (U3134, U3958, U5508);
  nand ginst6579 (U3135, U3959, U5511);
  nand ginst6580 (U3136, U3920, U5424);
  nand ginst6581 (U3137, U3921, U5427);
  nand ginst6582 (U3138, U3922, U5430);
  nand ginst6583 (U3139, U3923, U5433);
  nand ginst6584 (U3140, U3924, U5436);
  nand ginst6585 (U3141, U3925, U5439);
  nand ginst6586 (U3142, U3928, U5448);
  nand ginst6587 (U3143, U3949, U5481);
  nand ginst6588 (U3144, U3960, U5514);
  nand ginst6589 (U3145, U3961, U5517);
  nand ginst6590 (U3146, U4201, U5748);
  nand ginst6591 (U3147, U3372, U5808);
  nand ginst6592 (U3148, STATE_REG_SCAN_IN, U4062);
  not ginst6593 (U3149, STATE_REG_SCAN_IN);
  nand ginst6594 (U3150, U5692, U5693);
  nand ginst6595 (U3151, U5694, U5695);
  nand ginst6596 (U3152, U5696, U5697);
  nand ginst6597 (U3153, U5698, U5699);
  nand ginst6598 (U3154, U5700, U5701);
  nand ginst6599 (U3155, U5702, U5703);
  nand ginst6600 (U3156, U5704, U5705);
  nand ginst6601 (U3157, U5706, U5707);
  nand ginst6602 (U3158, U5708, U5709);
  nand ginst6603 (U3159, U5712, U5713);
  nand ginst6604 (U3160, U5714, U5715);
  nand ginst6605 (U3161, U5716, U5717);
  nand ginst6606 (U3162, U5718, U5719);
  nand ginst6607 (U3163, U5720, U5721);
  nand ginst6608 (U3164, U5722, U5723);
  nand ginst6609 (U3165, U5724, U5725);
  nand ginst6610 (U3166, U5726, U5727);
  nand ginst6611 (U3167, U5728, U5729);
  nand ginst6612 (U3168, U5730, U5731);
  nand ginst6613 (U3169, U5678, U5679);
  nand ginst6614 (U3170, U5680, U5681);
  nand ginst6615 (U3171, U5682, U5683);
  nand ginst6616 (U3172, U5684, U5685);
  nand ginst6617 (U3173, U5686, U5687);
  nand ginst6618 (U3174, U5688, U5689);
  nand ginst6619 (U3175, U5690, U5691);
  nand ginst6620 (U3176, U5710, U5711);
  nand ginst6621 (U3177, U5732, U5733);
  nand ginst6622 (U3178, U3966, U5735);
  nand ginst6623 (U3179, U5633, U5634);
  nand ginst6624 (U3180, U5635, U5636);
  nand ginst6625 (U3181, U5637, U5638);
  nand ginst6626 (U3182, U5639, U5640);
  nand ginst6627 (U3183, U5641, U5642);
  nand ginst6628 (U3184, U5643, U5644);
  nand ginst6629 (U3185, U5645, U5646);
  nand ginst6630 (U3186, U5647, U5648);
  nand ginst6631 (U3187, U5649, U5650);
  nand ginst6632 (U3188, U5653, U5654);
  nand ginst6633 (U3189, U5655, U5656);
  nand ginst6634 (U3190, U5657, U5658);
  nand ginst6635 (U3191, U5659, U5660);
  nand ginst6636 (U3192, U5661, U5662);
  nand ginst6637 (U3193, U5663, U5664);
  nand ginst6638 (U3194, U5665, U5666);
  nand ginst6639 (U3195, U5667, U5668);
  nand ginst6640 (U3196, U5669, U5670);
  nand ginst6641 (U3197, U5671, U5672);
  nand ginst6642 (U3198, U5619, U5620);
  nand ginst6643 (U3199, U5621, U5622);
  nand ginst6644 (U3200, U5623, U5624);
  nand ginst6645 (U3201, U5625, U5626);
  nand ginst6646 (U3202, U5627, U5628);
  nand ginst6647 (U3203, U5629, U5630);
  nand ginst6648 (U3204, U5631, U5632);
  nand ginst6649 (U3205, U5651, U5652);
  nand ginst6650 (U3206, U5673, U5674);
  nand ginst6651 (U3207, U3965, U5675);
  and ginst6652 (U3208, U3355, U5612);
  nand ginst6653 (U3209, U5422, U6258, U6259);
  nand ginst6654 (U3210, U5415, U5416, U5417, U5418, U5419);
  nand ginst6655 (U3211, U5406, U5407, U5408, U5409, U5410);
  nand ginst6656 (U3212, U5397, U5398, U5399, U5400, U5401);
  nand ginst6657 (U3213, U5388, U5389, U5390, U5391, U5392);
  nand ginst6658 (U3214, U5379, U5380, U5381, U5382, U5383);
  nand ginst6659 (U3215, U3918, U5371, U5372);
  nand ginst6660 (U3216, U5361, U5362, U5363, U5364, U5365);
  nand ginst6661 (U3217, U5352, U5353, U5354, U5355, U5356);
  nand ginst6662 (U3218, U5343, U5344, U5345, U5346, U5347);
  nand ginst6663 (U3219, U3916, U5335, U5336);
  nand ginst6664 (U3220, U5325, U5326, U5327, U5328, U5329);
  nand ginst6665 (U3221, U5316, U5317, U5318, U5319, U5320);
  nand ginst6666 (U3222, U5307, U5308, U5309, U5310, U5311);
  nand ginst6667 (U3223, U5298, U5299, U5300, U5301, U5302);
  nand ginst6668 (U3224, U3915, U5289, U5290, U5291);
  nand ginst6669 (U3225, U5280, U5281, U5282, U5283, U5284);
  nand ginst6670 (U3226, U5271, U5272, U5273, U5274, U5275);
  nand ginst6671 (U3227, U3914, U5262, U5263, U5264);
  nand ginst6672 (U3228, U5253, U5254, U5255, U5256, U5257);
  nand ginst6673 (U3229, U3912, U3913, U5246);
  nand ginst6674 (U3230, U5236, U5237, U5238, U5239, U5240);
  nand ginst6675 (U3231, U5227, U5228, U5229, U5230, U5231);
  nand ginst6676 (U3232, U5218, U5219, U5220, U5221, U5222);
  nand ginst6677 (U3233, U5209, U5210, U5211, U5212, U5213);
  nand ginst6678 (U3234, U3909, U5201, U5202);
  nand ginst6679 (U3235, U5191, U5192, U5193, U5194, U5195);
  nand ginst6680 (U3236, U5182, U5183, U5184, U5185, U5186);
  nand ginst6681 (U3237, U5173, U5174, U5175, U5176, U5177);
  nand ginst6682 (U3238, U5160, U5161, U5162, U5163, U5164);
  nand ginst6683 (U3239, U3904, U5147);
  nand ginst6684 (U3240, U3889, U3890);
  nand ginst6685 (U3241, U3887, U3888);
  nand ginst6686 (U3242, U3885, U3886);
  nand ginst6687 (U3243, U3882, U3883);
  nand ginst6688 (U3244, U3880, U3881);
  nand ginst6689 (U3245, U3877, U3878);
  nand ginst6690 (U3246, U3875, U3876);
  nand ginst6691 (U3247, U3873, U3874);
  nand ginst6692 (U3248, U3871, U3872, U5050, U5054);
  nand ginst6693 (U3249, U3869, U3870, U5040, U5044);
  nand ginst6694 (U3250, U3867, U3868, U5030, U5034);
  nand ginst6695 (U3251, U3865, U3866, U5020, U5024);
  nand ginst6696 (U3252, U3863, U3864, U5010, U5014);
  nand ginst6697 (U3253, U3861, U3862, U5000, U5004);
  nand ginst6698 (U3254, U3859, U3860, U4990, U4994);
  nand ginst6699 (U3255, U3857, U3858, U4980, U4984);
  nand ginst6700 (U3256, U3855, U3856, U4970, U4974);
  nand ginst6701 (U3257, U3853, U3854, U4960, U4964);
  nand ginst6702 (U3258, U3850, U3852);
  nand ginst6703 (U3259, U3846, U3848);
  nand ginst6704 (U3260, U4004, U4936, U4937);
  nand ginst6705 (U3261, U4003, U4934, U4935);
  nand ginst6706 (U3262, U3836, U3837, U4000, U4927);
  nand ginst6707 (U3263, U3834, U3835, U3999, U4922);
  nand ginst6708 (U3264, U3832, U3833, U3998, U4917);
  nand ginst6709 (U3265, U3830, U3831, U3997, U4912);
  nand ginst6710 (U3266, U3828, U3829, U3996, U4907);
  nand ginst6711 (U3267, U3826, U3827, U3995, U4902);
  nand ginst6712 (U3268, U3824, U3825, U3994, U4897);
  nand ginst6713 (U3269, U3822, U3823, U3993, U4892);
  nand ginst6714 (U3270, U3820, U3821, U3992, U4887);
  nand ginst6715 (U3271, U3818, U3819, U3991, U4882);
  nand ginst6716 (U3272, U3816, U3817, U3990, U4877);
  nand ginst6717 (U3273, U3814, U3815, U3989, U4872);
  nand ginst6718 (U3274, U3812, U3813, U3988, U4867);
  nand ginst6719 (U3275, U3810, U3811, U3987, U4862);
  nand ginst6720 (U3276, U3808, U3809, U3986);
  nand ginst6721 (U3277, U3806, U3807, U3985, U4852);
  nand ginst6722 (U3278, U3804, U3805, U3984);
  nand ginst6723 (U3279, U3802, U3803, U3983);
  nand ginst6724 (U3280, U3800, U3801, U3982);
  nand ginst6725 (U3281, U3798, U3799, U3981);
  nand ginst6726 (U3282, U3796, U3797, U3980);
  nand ginst6727 (U3283, U3794, U3795, U3979);
  nand ginst6728 (U3284, U3792, U3793, U3978);
  nand ginst6729 (U3285, U3790, U3791, U3977);
  nand ginst6730 (U3286, U3788, U3789);
  nand ginst6731 (U3287, U3786, U3787);
  nand ginst6732 (U3288, U3784, U3785);
  nand ginst6733 (U3289, U3782, U3783);
  nand ginst6734 (U3290, U3780, U3781);
  and ginst6735 (U3291, D_REG_31__SCAN_IN, U3968);
  and ginst6736 (U3292, D_REG_30__SCAN_IN, U3968);
  and ginst6737 (U3293, D_REG_29__SCAN_IN, U3968);
  and ginst6738 (U3294, D_REG_28__SCAN_IN, U3968);
  and ginst6739 (U3295, D_REG_27__SCAN_IN, U3968);
  and ginst6740 (U3296, D_REG_26__SCAN_IN, U3968);
  and ginst6741 (U3297, D_REG_25__SCAN_IN, U3968);
  and ginst6742 (U3298, D_REG_24__SCAN_IN, U3968);
  and ginst6743 (U3299, D_REG_23__SCAN_IN, U3968);
  and ginst6744 (U3300, D_REG_22__SCAN_IN, U3968);
  and ginst6745 (U3301, D_REG_21__SCAN_IN, U3968);
  and ginst6746 (U3302, D_REG_20__SCAN_IN, U3968);
  and ginst6747 (U3303, D_REG_19__SCAN_IN, U3968);
  and ginst6748 (U3304, D_REG_18__SCAN_IN, U3968);
  and ginst6749 (U3305, D_REG_17__SCAN_IN, U3968);
  and ginst6750 (U3306, D_REG_16__SCAN_IN, U3968);
  and ginst6751 (U3307, D_REG_15__SCAN_IN, U3968);
  and ginst6752 (U3308, D_REG_14__SCAN_IN, U3968);
  and ginst6753 (U3309, D_REG_13__SCAN_IN, U3968);
  and ginst6754 (U3310, D_REG_12__SCAN_IN, U3968);
  and ginst6755 (U3311, D_REG_11__SCAN_IN, U3968);
  and ginst6756 (U3312, D_REG_10__SCAN_IN, U3968);
  and ginst6757 (U3313, D_REG_9__SCAN_IN, U3968);
  and ginst6758 (U3314, D_REG_8__SCAN_IN, U3968);
  and ginst6759 (U3315, D_REG_7__SCAN_IN, U3968);
  xor ginst6760 (U3316, U3316_in, flip_signal);
  and ginst6761 (U3316_in, D_REG_6__SCAN_IN, U3968);
  and ginst6762 (U3317, D_REG_5__SCAN_IN, U3968);
  and ginst6763 (U3318, D_REG_4__SCAN_IN, U3968);
  and ginst6764 (U3319, D_REG_3__SCAN_IN, U3968);
  and ginst6765 (U3320, D_REG_2__SCAN_IN, U3968);
  nand ginst6766 (U3321, U3645, U4159);
  nand ginst6767 (U3322, U3644, U4156);
  nand ginst6768 (U3323, U3643, U4153);
  nand ginst6769 (U3324, U3642, U4150);
  nand ginst6770 (U3325, U3641, U4147);
  nand ginst6771 (U3326, U3640, U4144);
  nand ginst6772 (U3327, U3639, U4141);
  nand ginst6773 (U3328, U3638, U4138);
  nand ginst6774 (U3329, U3637, U4135);
  nand ginst6775 (U3330, U3636, U4132);
  nand ginst6776 (U3331, U3635, U4129);
  nand ginst6777 (U3332, U3634, U4126);
  nand ginst6778 (U3333, U3633, U4123);
  nand ginst6779 (U3334, U3632, U4120);
  nand ginst6780 (U3335, U3631, U4117);
  nand ginst6781 (U3336, U3630, U4114);
  nand ginst6782 (U3337, U3629, U4111);
  nand ginst6783 (U3338, U3628, U4108);
  nand ginst6784 (U3339, U3627, U4105);
  nand ginst6785 (U3340, U3626, U4102);
  nand ginst6786 (U3341, U3625, U4099);
  nand ginst6787 (U3342, U3624, U4096);
  nand ginst6788 (U3343, U3623, U4093);
  nand ginst6789 (U3344, U3622, U4090);
  nand ginst6790 (U3345, U3621, U4087);
  nand ginst6791 (U3346, U3620, U4084);
  nand ginst6792 (U3347, U3619, U4081);
  nand ginst6793 (U3348, U3618, U4078);
  nand ginst6794 (U3349, U3617, U4075);
  nand ginst6795 (U3350, U3616, U4072);
  nand ginst6796 (U3351, U3615, U4069);
  nand ginst6797 (U3352, U3614, U4066);
  nand ginst6798 (U3353, U4055, U5805);
  nand ginst6799 (U3354, U4001, U4930, U4931, U4932, U4933);
  nand ginst6800 (U3355, U3432, U3433, U3434);
  nand ginst6801 (U3356, U4059, U5748);
  nand ginst6802 (U3357, STATE_REG_SCAN_IN, U3967);
  nand ginst6803 (U3358, U3432, U5757);
  not ginst6804 (U3359, B_REG_SCAN_IN);
  nand ginst6805 (U3360, U3432, U5809, U5810);
  nand ginst6806 (U3361, U3456, U5820);
  nand ginst6807 (U3362, U3461, U4201);
  nand ginst6808 (U3363, U3456, U3460, U3461);
  nand ginst6809 (U3364, U3456, U3460, U5817);
  nand ginst6810 (U3365, U3457, U3460);
  nand ginst6811 (U3366, U3461, U4056);
  nand ginst6812 (U3367, U4056, U5817);
  nand ginst6813 (U3368, U4201, U5817);
  nand ginst6814 (U3369, U4015, U5808);
  nand ginst6815 (U3370, U3457, U5817, U5820);
  nand ginst6816 (U3371, U4011, U5805);
  nand ginst6817 (U3372, U3461, U5805);
  nand ginst6818 (U3373, U3456, U3457);
  nand ginst6819 (U3374, U3460, U5808);
  nand ginst6820 (U3375, U3646, U3647, U4206, U4207, U4208);
  not ginst6821 (U3376, REG2_REG_0__SCAN_IN);
  nand ginst6822 (U3377, U3662, U3664, U4225, U4226);
  nand ginst6823 (U3378, U3666, U3668, U4244, U4245);
  nand ginst6824 (U3379, U3670, U3672, U4263, U4264);
  nand ginst6825 (U3380, U3674, U3676, U4282, U4283);
  nand ginst6826 (U3381, U3678, U3680, U4301, U4302);
  nand ginst6827 (U3382, U3682, U3684, U4320, U4321);
  nand ginst6828 (U3383, U3686, U3688, U4339, U4340);
  nand ginst6829 (U3384, U3690, U3692, U4358, U4359);
  nand ginst6830 (U3385, U3694, U3696, U4377, U4378);
  nand ginst6831 (U3386, U3698, U3700, U4396, U4397);
  nand ginst6832 (U3387, U3702, U3704, U4415, U4416);
  nand ginst6833 (U3388, U3706, U3708, U4434, U4435);
  nand ginst6834 (U3389, U3710, U3712, U4453, U4454);
  nand ginst6835 (U3390, U3714, U3716, U4472, U4473);
  nand ginst6836 (U3391, U3718, U3720, U4491, U4492);
  nand ginst6837 (U3392, U3722, U3724, U4510, U4511);
  nand ginst6838 (U3393, U3726, U3728, U4529, U4530);
  nand ginst6839 (U3394, U3730, U3732, U4548, U4549);
  nand ginst6840 (U3395, U3734, U3736, U4567, U4568);
  nand ginst6841 (U3396, DATAI_20_, U3969);
  nand ginst6842 (U3397, U3738, U3740, U4586, U4587);
  nand ginst6843 (U3398, DATAI_21_, U3969);
  nand ginst6844 (U3399, U3742, U3744, U4605, U4606);
  nand ginst6845 (U3400, DATAI_22_, U3969);
  nand ginst6846 (U3401, U3746, U3748, U4624, U4625);
  nand ginst6847 (U3402, DATAI_23_, U3969);
  nand ginst6848 (U3403, U3750, U3752, U4643, U4644);
  nand ginst6849 (U3404, DATAI_24_, U3969);
  nand ginst6850 (U3405, U3754, U3756, U4662, U4663);
  nand ginst6851 (U3406, DATAI_25_, U3969);
  nand ginst6852 (U3407, U3758, U3760, U4681, U4682);
  nand ginst6853 (U3408, DATAI_26_, U3969);
  nand ginst6854 (U3409, U3762, U3764, U4700, U4701);
  nand ginst6855 (U3410, DATAI_27_, U3969);
  nand ginst6856 (U3411, U3766, U3768, U4719, U4720);
  nand ginst6857 (U3412, DATAI_28_, U3969);
  nand ginst6858 (U3413, U3770, U3772, U4738, U4739);
  nand ginst6859 (U3414, DATAI_29_, U3969);
  nand ginst6860 (U3415, DATAI_30_, U3969);
  nand ginst6861 (U3416, DATAI_31_, U3969);
  nand ginst6862 (U3417, U3023, U4784);
  nand ginst6863 (U3418, U4010, U5808, U5820);
  nand ginst6864 (U3419, U3457, U3461, U5820);
  nand ginst6865 (U3420, U3024, U5817);
  nand ginst6866 (U3421, U3356, U4063);
  nand ginst6867 (U3422, STATE_REG_SCAN_IN, U4054);
  nand ginst6868 (U3423, U3015, U3016);
  not ginst6869 (U3424, R395_U6);
  nand ginst6870 (U3425, U3900, U3901);
  nand ginst6871 (U3426, U3023, U4021);
  nand ginst6872 (U3427, U3017, U3905);
  nand ginst6873 (U3428, U3015, U3023);
  nand ginst6874 (U3429, U3907, U5158);
  nand ginst6875 (U3430, U3461, U5808);
  nand ginst6876 (U3431, U5746, U5747);
  nand ginst6877 (U3432, U5752, U5753);
  nand ginst6878 (U3433, U5755, U5756);
  nand ginst6879 (U3434, U5749, U5750);
  nand ginst6880 (U3435, U5758, U5759);
  nand ginst6881 (U3436, U5760, U5761);
  nand ginst6882 (U3437, U5762, U5763);
  nand ginst6883 (U3438, U5764, U5765);
  nand ginst6884 (U3439, U5766, U5767);
  nand ginst6885 (U3440, U5768, U5769);
  nand ginst6886 (U3441, U5770, U5771);
  nand ginst6887 (U3442, U5772, U5773);
  nand ginst6888 (U3443, U5774, U5775);
  nand ginst6889 (U3444, U5776, U5777);
  nand ginst6890 (U3445, U5778, U5779);
  nand ginst6891 (U3446, U5780, U5781);
  nand ginst6892 (U3447, U5782, U5783);
  nand ginst6893 (U3448, U5784, U5785);
  nand ginst6894 (U3449, U5786, U5787);
  nand ginst6895 (U3450, U5788, U5789);
  nand ginst6896 (U3451, U5790, U5791);
  nand ginst6897 (U3452, U5792, U5793);
  nand ginst6898 (U3453, U5794, U5795);
  nand ginst6899 (U3454, U5797, U5798);
  nand ginst6900 (U3455, U5800, U5801);
  nand ginst6901 (U3456, U5803, U5804);
  nand ginst6902 (U3457, U5806, U5807);
  nand ginst6903 (U3458, U5811, U5812);
  nand ginst6904 (U3459, U5813, U5814);
  nand ginst6905 (U3460, U5818, U5819);
  nand ginst6906 (U3461, U5815, U5816);
  nand ginst6907 (U3462, U5821, U5822);
  nand ginst6908 (U3463, U5824, U5825);
  nand ginst6909 (U3464, U5827, U5828);
  nand ginst6910 (U3465, U5835, U5836);
  nand ginst6911 (U3466, U5832, U5833);
  nand ginst6912 (U3467, U5838, U5839);
  nand ginst6913 (U3468, U5840, U5841);
  nand ginst6914 (U3469, U5843, U5844);
  nand ginst6915 (U3470, U5845, U5846);
  nand ginst6916 (U3471, U5848, U5849);
  nand ginst6917 (U3472, U5850, U5851);
  nand ginst6918 (U3473, U5853, U5854);
  nand ginst6919 (U3474, U5855, U5856);
  nand ginst6920 (U3475, U5858, U5859);
  nand ginst6921 (U3476, U5860, U5861);
  nand ginst6922 (U3477, U5863, U5864);
  nand ginst6923 (U3478, U5865, U5866);
  nand ginst6924 (U3479, U5868, U5869);
  nand ginst6925 (U3480, U5870, U5871);
  nand ginst6926 (U3481, U5873, U5874);
  nand ginst6927 (U3482, U5875, U5876);
  nand ginst6928 (U3483, U5878, U5879);
  nand ginst6929 (U3484, U5880, U5881);
  nand ginst6930 (U3485, U5883, U5884);
  nand ginst6931 (U3486, U5885, U5886);
  nand ginst6932 (U3487, U5888, U5889);
  nand ginst6933 (U3488, U5890, U5891);
  nand ginst6934 (U3489, U5893, U5894);
  nand ginst6935 (U3490, U5895, U5896);
  nand ginst6936 (U3491, U5898, U5899);
  nand ginst6937 (U3492, U5900, U5901);
  nand ginst6938 (U3493, U5903, U5904);
  nand ginst6939 (U3494, U5905, U5906);
  nand ginst6940 (U3495, U5908, U5909);
  nand ginst6941 (U3496, U5910, U5911);
  nand ginst6942 (U3497, U5913, U5914);
  nand ginst6943 (U3498, U5915, U5916);
  nand ginst6944 (U3499, U5918, U5919);
  nand ginst6945 (U3500, U5920, U5921);
  nand ginst6946 (U3501, U5923, U5924);
  nand ginst6947 (U3502, U5925, U5926);
  nand ginst6948 (U3503, U5928, U5929);
  nand ginst6949 (U3504, U5930, U5931);
  nand ginst6950 (U3505, U5933, U5934);
  nand ginst6951 (U3506, U5935, U5936);
  nand ginst6952 (U3507, U5937, U5938);
  nand ginst6953 (U3508, U5939, U5940);
  nand ginst6954 (U3509, U5941, U5942);
  nand ginst6955 (U3510, U5943, U5944);
  nand ginst6956 (U3511, U5945, U5946);
  nand ginst6957 (U3512, U5947, U5948);
  nand ginst6958 (U3513, U5949, U5950);
  nand ginst6959 (U3514, U5951, U5952);
  nand ginst6960 (U3515, U5953, U5954);
  nand ginst6961 (U3516, U5955, U5956);
  nand ginst6962 (U3517, U5957, U5958);
  nand ginst6963 (U3518, U5959, U5960);
  nand ginst6964 (U3519, U5961, U5962);
  nand ginst6965 (U3520, U5963, U5964);
  nand ginst6966 (U3521, U5965, U5966);
  nand ginst6967 (U3522, U5967, U5968);
  nand ginst6968 (U3523, U5969, U5970);
  nand ginst6969 (U3524, U5971, U5972);
  nand ginst6970 (U3525, U5973, U5974);
  nand ginst6971 (U3526, U5975, U5976);
  nand ginst6972 (U3527, U5977, U5978);
  nand ginst6973 (U3528, U5979, U5980);
  nand ginst6974 (U3529, U5981, U5982);
  nand ginst6975 (U3530, U5983, U5984);
  nand ginst6976 (U3531, U5985, U5986);
  nand ginst6977 (U3532, U5987, U5988);
  nand ginst6978 (U3533, U5989, U5990);
  nand ginst6979 (U3534, U5991, U5992);
  nand ginst6980 (U3535, U5993, U5994);
  nand ginst6981 (U3536, U5995, U5996);
  nand ginst6982 (U3537, U5997, U5998);
  nand ginst6983 (U3538, U5999, U6000);
  nand ginst6984 (U3539, U6001, U6002);
  nand ginst6985 (U3540, U6003, U6004);
  nand ginst6986 (U3541, U6005, U6006);
  nand ginst6987 (U3542, U6007, U6008);
  nand ginst6988 (U3543, U6009, U6010);
  nand ginst6989 (U3544, U6011, U6012);
  nand ginst6990 (U3545, U6013, U6014);
  nand ginst6991 (U3546, U6015, U6016);
  nand ginst6992 (U3547, U6017, U6018);
  nand ginst6993 (U3548, U6019, U6020);
  nand ginst6994 (U3549, U6021, U6022);
  nand ginst6995 (U3550, U6087, U6088);
  nand ginst6996 (U3551, U6089, U6090);
  nand ginst6997 (U3552, U6091, U6092);
  nand ginst6998 (U3553, U6093, U6094);
  nand ginst6999 (U3554, U6095, U6096);
  nand ginst7000 (U3555, U6097, U6098);
  nand ginst7001 (U3556, U6099, U6100);
  nand ginst7002 (U3557, U6101, U6102);
  nand ginst7003 (U3558, U6103, U6104);
  nand ginst7004 (U3559, U6105, U6106);
  nand ginst7005 (U3560, U6107, U6108);
  nand ginst7006 (U3561, U6109, U6110);
  nand ginst7007 (U3562, U6111, U6112);
  nand ginst7008 (U3563, U6113, U6114);
  nand ginst7009 (U3564, U6115, U6116);
  nand ginst7010 (U3565, U6117, U6118);
  nand ginst7011 (U3566, U6119, U6120);
  nand ginst7012 (U3567, U6121, U6122);
  nand ginst7013 (U3568, U6123, U6124);
  nand ginst7014 (U3569, U6125, U6126);
  nand ginst7015 (U3570, U6127, U6128);
  nand ginst7016 (U3571, U6129, U6130);
  nand ginst7017 (U3572, U6131, U6132);
  nand ginst7018 (U3573, U6133, U6134);
  nand ginst7019 (U3574, U6135, U6136);
  nand ginst7020 (U3575, U6137, U6138);
  nand ginst7021 (U3576, U6139, U6140);
  nand ginst7022 (U3577, U6141, U6142);
  nand ginst7023 (U3578, U6143, U6144);
  nand ginst7024 (U3579, U6145, U6146);
  nand ginst7025 (U3580, U6147, U6148);
  nand ginst7026 (U3581, U6149, U6150);
  nand ginst7027 (U3582, U6260, U6261);
  nand ginst7028 (U3583, U6262, U6263);
  nand ginst7029 (U3584, U6264, U6265);
  nand ginst7030 (U3585, U6266, U6267);
  nand ginst7031 (U3586, U6268, U6269);
  nand ginst7032 (U3587, U6270, U6271);
  nand ginst7033 (U3588, U6272, U6273);
  nand ginst7034 (U3589, U6274, U6275);
  nand ginst7035 (U3590, U6276, U6277);
  nand ginst7036 (U3591, U6278, U6279);
  nand ginst7037 (U3592, U6280, U6281);
  nand ginst7038 (U3593, U6282, U6283);
  nand ginst7039 (U3594, U6284, U6285);
  nand ginst7040 (U3595, U6286, U6287);
  nand ginst7041 (U3596, U6288, U6289);
  nand ginst7042 (U3597, U6290, U6291);
  nand ginst7043 (U3598, U6292, U6293);
  nand ginst7044 (U3599, U6294, U6295);
  nand ginst7045 (U3600, U6296, U6297);
  nand ginst7046 (U3601, U6298, U6299);
  nand ginst7047 (U3602, U6300, U6301);
  nand ginst7048 (U3603, U6302, U6303);
  nand ginst7049 (U3604, U6304, U6305);
  nand ginst7050 (U3605, U6306, U6307);
  nand ginst7051 (U3606, U6308, U6309);
  nand ginst7052 (U3607, U6310, U6311);
  nand ginst7053 (U3608, U6312, U6313);
  nand ginst7054 (U3609, U6314, U6315);
  nand ginst7055 (U3610, U6316, U6317);
  nand ginst7056 (U3611, U6318, U6319);
  nand ginst7057 (U3612, U6320, U6321);
  nand ginst7058 (U3613, U6322, U6323);
  and ginst7059 (U3614, U4065, U4067);
  and ginst7060 (U3615, U4068, U4070);
  and ginst7061 (U3616, U4071, U4073);
  and ginst7062 (U3617, U4074, U4076);
  and ginst7063 (U3618, U4077, U4079);
  and ginst7064 (U3619, U4080, U4082);
  and ginst7065 (U3620, U4083, U4085);
  and ginst7066 (U3621, U4086, U4088);
  and ginst7067 (U3622, U4089, U4091);
  and ginst7068 (U3623, U4092, U4094);
  and ginst7069 (U3624, U4095, U4097);
  and ginst7070 (U3625, U4098, U4100);
  and ginst7071 (U3626, U4101, U4103);
  and ginst7072 (U3627, U4104, U4106);
  and ginst7073 (U3628, U4107, U4109);
  and ginst7074 (U3629, U4110, U4112);
  and ginst7075 (U3630, U4113, U4115);
  and ginst7076 (U3631, U4116, U4118);
  and ginst7077 (U3632, U4119, U4121);
  and ginst7078 (U3633, U4122, U4124);
  and ginst7079 (U3634, U4125, U4127);
  and ginst7080 (U3635, U4128, U4130);
  and ginst7081 (U3636, U4131, U4133);
  and ginst7082 (U3637, U4134, U4136);
  and ginst7083 (U3638, U4137, U4139);
  and ginst7084 (U3639, U4140, U4142);
  and ginst7085 (U3640, U4143, U4145);
  and ginst7086 (U3641, U4146, U4148);
  and ginst7087 (U3642, U4149, U4151);
  and ginst7088 (U3643, U4152, U4154);
  and ginst7089 (U3644, U4155, U4157);
  and ginst7090 (U3645, U4158, U4160);
  and ginst7091 (U3646, U4202, U4203);
  and ginst7092 (U3647, U4204, U4205);
  and ginst7093 (U3648, U4210, U4212);
  and ginst7094 (U3649, U3648, U4211, U4213);
  and ginst7095 (U3650, U4164, U4165, U4166, U4167);
  and ginst7096 (U3651, U4168, U4169, U4170, U4171);
  and ginst7097 (U3652, U4172, U4173, U4174, U4175);
  and ginst7098 (U3653, U4176, U4177, U4178);
  and ginst7099 (U3654, U3650, U3651, U3652, U3653);
  and ginst7100 (U3655, U4179, U4180, U4181, U4182);
  and ginst7101 (U3656, U4183, U4184, U4185, U4186);
  and ginst7102 (U3657, U4187, U4188, U4189, U4190);
  and ginst7103 (U3658, U4191, U4192, U4193);
  and ginst7104 (U3659, U3655, U3656, U3657, U3658);
  and ginst7105 (U3660, U4195, U5834);
  and ginst7106 (U3661, U3023, U5837);
  and ginst7107 (U3662, U4227, U4228);
  and ginst7108 (U3663, U4229, U4230);
  and ginst7109 (U3664, U3663, U4231, U4232);
  and ginst7110 (U3665, U4234, U4235, U4236, U4237);
  and ginst7111 (U3666, U4246, U4247);
  and ginst7112 (U3667, U4248, U4249);
  and ginst7113 (U3668, U3667, U4250, U4251);
  and ginst7114 (U3669, U4253, U4254, U4255, U4256);
  and ginst7115 (U3670, U4265, U4266);
  and ginst7116 (U3671, U4267, U4268);
  and ginst7117 (U3672, U3671, U4269, U4270);
  and ginst7118 (U3673, U4272, U4273, U4274, U4275);
  and ginst7119 (U3674, U4284, U4285);
  and ginst7120 (U3675, U4286, U4287);
  and ginst7121 (U3676, U3675, U4288, U4289);
  and ginst7122 (U3677, U4291, U4292, U4293, U4294);
  and ginst7123 (U3678, U4303, U4304);
  and ginst7124 (U3679, U4305, U4306);
  and ginst7125 (U3680, U3679, U4307, U4308);
  and ginst7126 (U3681, U4310, U4311, U4312, U4313);
  and ginst7127 (U3682, U4322, U4323);
  and ginst7128 (U3683, U4324, U4325);
  and ginst7129 (U3684, U3683, U4326, U4327);
  and ginst7130 (U3685, U4329, U4330, U4331, U4332);
  and ginst7131 (U3686, U4341, U4342);
  and ginst7132 (U3687, U4343, U4344);
  and ginst7133 (U3688, U3687, U4345, U4346);
  and ginst7134 (U3689, U4348, U4349, U4350, U4351);
  and ginst7135 (U3690, U4360, U4361);
  and ginst7136 (U3691, U4362, U4363);
  and ginst7137 (U3692, U3691, U4364, U4365);
  and ginst7138 (U3693, U4367, U4368, U4369, U4370);
  and ginst7139 (U3694, U4379, U4380);
  and ginst7140 (U3695, U4381, U4382);
  and ginst7141 (U3696, U3695, U4383, U4384);
  and ginst7142 (U3697, U4386, U4387, U4388, U4389);
  and ginst7143 (U3698, U4398, U4399);
  and ginst7144 (U3699, U4400, U4401);
  and ginst7145 (U3700, U3699, U4402, U4403);
  and ginst7146 (U3701, U4405, U4406, U4407, U4408);
  and ginst7147 (U3702, U4417, U4418);
  and ginst7148 (U3703, U4419, U4420);
  and ginst7149 (U3704, U3703, U4421, U4422);
  and ginst7150 (U3705, U4424, U4425, U4426, U4427);
  and ginst7151 (U3706, U4436, U4437);
  and ginst7152 (U3707, U4438, U4439);
  and ginst7153 (U3708, U3707, U4440, U4441);
  and ginst7154 (U3709, U4443, U4444, U4445, U4446);
  and ginst7155 (U3710, U4455, U4456);
  and ginst7156 (U3711, U4457, U4458);
  and ginst7157 (U3712, U3711, U4459, U4460);
  and ginst7158 (U3713, U4462, U4463, U4464, U4465);
  and ginst7159 (U3714, U4474, U4475);
  and ginst7160 (U3715, U4476, U4477);
  and ginst7161 (U3716, U3715, U4478, U4479);
  and ginst7162 (U3717, U4481, U4482, U4483, U4484);
  and ginst7163 (U3718, U4493, U4494);
  and ginst7164 (U3719, U4495, U4496);
  and ginst7165 (U3720, U3719, U4497, U4498);
  and ginst7166 (U3721, U4500, U4501, U4502, U4503);
  and ginst7167 (U3722, U4512, U4513);
  and ginst7168 (U3723, U4514, U4515);
  and ginst7169 (U3724, U3723, U4516, U4517);
  and ginst7170 (U3725, U4519, U4520, U4521, U4522);
  and ginst7171 (U3726, U4531, U4532);
  and ginst7172 (U3727, U4533, U4534);
  and ginst7173 (U3728, U3727, U4535, U4536);
  and ginst7174 (U3729, U4538, U4539, U4540, U4541);
  and ginst7175 (U3730, U4550, U4551);
  and ginst7176 (U3731, U4552, U4553);
  and ginst7177 (U3732, U3731, U4554, U4555);
  and ginst7178 (U3733, U4557, U4558, U4559, U4560);
  and ginst7179 (U3734, U4569, U4570);
  and ginst7180 (U3735, U4571, U4572);
  and ginst7181 (U3736, U3735, U4573, U4574);
  and ginst7182 (U3737, U4576, U4577, U4578, U4579);
  and ginst7183 (U3738, U4588, U4589);
  and ginst7184 (U3739, U4590, U4591);
  and ginst7185 (U3740, U3739, U4592, U4593);
  and ginst7186 (U3741, U4595, U4596, U4597, U4598);
  and ginst7187 (U3742, U4607, U4608);
  and ginst7188 (U3743, U4609, U4610);
  and ginst7189 (U3744, U3743, U4611, U4612);
  and ginst7190 (U3745, U4614, U4615, U4616, U4617);
  and ginst7191 (U3746, U4626, U4627);
  and ginst7192 (U3747, U4628, U4629);
  and ginst7193 (U3748, U3747, U4630, U4631);
  and ginst7194 (U3749, U4633, U4634, U4635, U4636);
  and ginst7195 (U3750, U4645, U4646);
  and ginst7196 (U3751, U4647, U4648);
  and ginst7197 (U3752, U3751, U4649, U4650);
  and ginst7198 (U3753, U4652, U4653, U4654, U4655);
  and ginst7199 (U3754, U4664, U4665);
  and ginst7200 (U3755, U4666, U4667);
  and ginst7201 (U3756, U3755, U4668, U4669);
  and ginst7202 (U3757, U4671, U4672, U4673, U4674);
  and ginst7203 (U3758, U4683, U4684);
  and ginst7204 (U3759, U4685, U4686);
  and ginst7205 (U3760, U3759, U4687, U4688);
  and ginst7206 (U3761, U4690, U4691, U4692, U4693);
  and ginst7207 (U3762, U4702, U4703);
  and ginst7208 (U3763, U4704, U4705);
  and ginst7209 (U3764, U3763, U4706, U4707);
  and ginst7210 (U3765, U4709, U4710, U4711, U4712);
  and ginst7211 (U3766, U4721, U4722);
  and ginst7212 (U3767, U4723, U4724);
  and ginst7213 (U3768, U3767, U4725, U4726);
  and ginst7214 (U3769, U4728, U4729, U4730, U4731);
  and ginst7215 (U3770, U4740, U4741);
  and ginst7216 (U3771, U4742, U4743);
  and ginst7217 (U3772, U3771, U4744, U4745);
  and ginst7218 (U3773, U4747, U4748, U4749, U4750);
  and ginst7219 (U3774, U4042, U4757);
  and ginst7220 (U3775, U4760, U4761, U4763, U4764);
  and ginst7221 (U3776, U4768, U4769, U4770);
  and ginst7222 (U3777, U4042, U4757);
  and ginst7223 (U3778, U3023, U3465);
  and ginst7224 (U3779, U3466, U4025, U5837);
  and ginst7225 (U3780, U4785, U4786, U4787);
  and ginst7226 (U3781, U3972, U4788, U4789);
  and ginst7227 (U3782, U4790, U4791, U4792);
  and ginst7228 (U3783, U3973, U4793, U4794);
  and ginst7229 (U3784, U4795, U4796, U4797);
  and ginst7230 (U3785, U3974, U4798, U4799);
  and ginst7231 (U3786, U4800, U4801, U4802);
  and ginst7232 (U3787, U3975, U4803, U4804);
  and ginst7233 (U3788, U4805, U4806, U4807);
  and ginst7234 (U3789, U3976, U4808, U4809);
  and ginst7235 (U3790, U4810, U4811, U4812);
  and ginst7236 (U3791, U4813, U4814);
  and ginst7237 (U3792, U4815, U4816, U4817);
  and ginst7238 (U3793, U4818, U4819);
  and ginst7239 (U3794, U4820, U4821, U4822);
  and ginst7240 (U3795, U4823, U4824);
  and ginst7241 (U3796, U4825, U4826, U4827);
  and ginst7242 (U3797, U4828, U4829);
  and ginst7243 (U3798, U4830, U4831, U4832);
  and ginst7244 (U3799, U4833, U4834);
  and ginst7245 (U3800, U4835, U4836, U4837);
  and ginst7246 (U3801, U4838, U4839);
  and ginst7247 (U3802, U4840, U4841, U4842);
  and ginst7248 (U3803, U4843, U4844);
  and ginst7249 (U3804, U4845, U4846, U4847);
  and ginst7250 (U3805, U4848, U4849);
  and ginst7251 (U3806, U4850, U4851);
  and ginst7252 (U3807, U4853, U4854);
  and ginst7253 (U3808, U4855, U4856, U4857);
  and ginst7254 (U3809, U4858, U4859);
  and ginst7255 (U3810, U4860, U4861);
  and ginst7256 (U3811, U4863, U4864);
  and ginst7257 (U3812, U4865, U4866);
  and ginst7258 (U3813, U4868, U4869);
  and ginst7259 (U3814, U4870, U4871);
  and ginst7260 (U3815, U4873, U4874);
  and ginst7261 (U3816, U4875, U4876);
  and ginst7262 (U3817, U4878, U4879);
  and ginst7263 (U3818, U4880, U4881);
  and ginst7264 (U3819, U4883, U4884);
  and ginst7265 (U3820, U4885, U4886);
  and ginst7266 (U3821, U4888, U4889);
  and ginst7267 (U3822, U4890, U4891);
  and ginst7268 (U3823, U4893, U4894);
  and ginst7269 (U3824, U4895, U4896);
  and ginst7270 (U3825, U4898, U4899);
  and ginst7271 (U3826, U4900, U4901);
  and ginst7272 (U3827, U4903, U4904);
  and ginst7273 (U3828, U4905, U4906);
  and ginst7274 (U3829, U4908, U4909);
  and ginst7275 (U3830, U4910, U4911);
  and ginst7276 (U3831, U4913, U4914);
  and ginst7277 (U3832, U4915, U4916);
  and ginst7278 (U3833, U4918, U4919);
  and ginst7279 (U3834, U4920, U4921);
  and ginst7280 (U3835, U4923, U4924);
  and ginst7281 (U3836, U4925, U4926);
  and ginst7282 (U3837, U4928, U4929);
  and ginst7283 (U3838, U5737, U5738, U5739);
  and ginst7284 (U3839, U3367, U3370, U3419);
  and ginst7285 (U3840, U3362, U3366, U3368);
  and ginst7286 (U3841, U3363, U3364);
  and ginst7287 (U3842, U3420, U3841);
  and ginst7288 (U3843, U3353, U3418);
  and ginst7289 (U3844, U3040, U3461);
  and ginst7290 (U3845, STATE_REG_SCAN_IN, U3431);
  and ginst7291 (U3846, U4939, U4940, U4941, U4943);
  and ginst7292 (U3847, U4944, U4947);
  and ginst7293 (U3848, U3847, U4945, U4946);
  and ginst7294 (U3849, U3040, U3444);
  and ginst7295 (U3850, U4948, U4949, U4950, U4951);
  and ginst7296 (U3851, U4952, U4955);
  and ginst7297 (U3852, U3851, U4953, U4954);
  and ginst7298 (U3853, U4961, U4962);
  and ginst7299 (U3854, U4963, U4965);
  and ginst7300 (U3855, U4971, U4972);
  and ginst7301 (U3856, U4973, U4975);
  and ginst7302 (U3857, U4981, U4982);
  and ginst7303 (U3858, U4983, U4985);
  and ginst7304 (U3859, U4991, U4992);
  and ginst7305 (U3860, U4993, U4995);
  and ginst7306 (U3861, U5001, U5002);
  and ginst7307 (U3862, U5003, U5005);
  and ginst7308 (U3863, U5011, U5012);
  and ginst7309 (U3864, U5013, U5015);
  and ginst7310 (U3865, U5021, U5022);
  and ginst7311 (U3866, U5023, U5025);
  and ginst7312 (U3867, U5031, U5032);
  and ginst7313 (U3868, U5033, U5035);
  and ginst7314 (U3869, U5041, U5042);
  and ginst7315 (U3870, U5043, U5045);
  and ginst7316 (U3871, U5051, U5052);
  and ginst7317 (U3872, U5053, U5055);
  and ginst7318 (U3873, U5060, U5061, U5062);
  and ginst7319 (U3874, U5063, U5064, U5065);
  and ginst7320 (U3875, U5070, U5071, U5072);
  and ginst7321 (U3876, U5073, U5074, U5075);
  and ginst7322 (U3877, U5080, U5081, U5082);
  and ginst7323 (U3878, U5083, U5084, U5085);
  and ginst7324 (U3879, U4053, U5090);
  and ginst7325 (U3880, U3879, U5091, U5092);
  and ginst7326 (U3881, U5093, U5094, U5095);
  and ginst7327 (U3882, U5100, U5101, U5102);
  and ginst7328 (U3883, U5103, U5104, U5105);
  and ginst7329 (U3884, U4053, U5110);
  and ginst7330 (U3885, U3884, U5111, U5112);
  and ginst7331 (U3886, U5113, U5114, U5115);
  and ginst7332 (U3887, U5120, U5121, U5122);
  and ginst7333 (U3888, U5123, U5124, U5125);
  and ginst7334 (U3889, U5130, U5131, U5132);
  and ginst7335 (U3890, U5133, U5134, U5135);
  and ginst7336 (U3891, U6201, U6204, U6207, U6210);
  and ginst7337 (U3892, U6213, U6216, U6219, U6222);
  and ginst7338 (U3893, U6225, U6228, U6231, U6234);
  and ginst7339 (U3894, U6237, U6240, U6243, U6246);
  and ginst7340 (U3895, U6165, U6168, U6171, U6174);
  and ginst7341 (U3896, U6156, U6159, U6162);
  and ginst7342 (U3897, U6183, U6186, U6189, U6192);
  and ginst7343 (U3898, U6177, U6180);
  and ginst7344 (U3899, U6195, U6198);
  and ginst7345 (U3900, U3895, U3896, U3897, U3898, U6153);
  and ginst7346 (U3901, U3891, U3892, U3893, U3894, U3899);
  and ginst7347 (U3902, U5140, U5141, U6254, U6255);
  and ginst7348 (U3903, STATE_REG_SCAN_IN, U3356);
  and ginst7349 (U3904, U5146, U5148);
  and ginst7350 (U3905, U3465, U3466);
  and ginst7351 (U3906, U3371, U3420, U4008);
  and ginst7352 (U3907, U3356, U4025, U5748);
  and ginst7353 (U3908, U3023, U5157);
  and ginst7354 (U3909, U3910, U5200);
  and ginst7355 (U3910, U5203, U5204);
  and ginst7356 (U3911, U3075, U4049);
  and ginst7357 (U3912, U5244, U5245);
  and ginst7358 (U3913, U5247, U5248);
  and ginst7359 (U3914, U5265, U5266);
  and ginst7360 (U3915, U5292, U5293);
  and ginst7361 (U3916, U3917, U5334);
  and ginst7362 (U3917, U5337, U5338);
  and ginst7363 (U3918, U3919, U5370);
  and ginst7364 (U3919, U5373, U5374);
  and ginst7365 (U3920, U3431, U5423, U5425);
  and ginst7366 (U3921, U3431, U5426, U5428);
  and ginst7367 (U3922, U3431, U5429, U5431);
  and ginst7368 (U3923, U3431, U5432, U5434);
  and ginst7369 (U3924, U3431, U5435, U5437);
  and ginst7370 (U3925, U3431, U5438, U5440);
  and ginst7371 (U3926, U5442, U5443);
  and ginst7372 (U3927, U5445, U5446);
  and ginst7373 (U3928, U3431, U5447, U5449);
  and ginst7374 (U3929, U3930, U5452);
  and ginst7375 (U3930, U3431, U5451);
  and ginst7376 (U3931, U3932, U5455);
  and ginst7377 (U3932, U3431, U5454);
  and ginst7378 (U3933, U3934, U5458);
  and ginst7379 (U3934, U3431, U5457);
  and ginst7380 (U3935, U3936, U5461);
  and ginst7381 (U3936, U3431, U5460);
  and ginst7382 (U3937, U3938, U5464);
  and ginst7383 (U3938, U3431, U5463);
  and ginst7384 (U3939, U3940, U5467);
  and ginst7385 (U3940, U3431, U5466);
  and ginst7386 (U3941, U3942, U5470);
  and ginst7387 (U3942, U3431, U5469);
  and ginst7388 (U3943, U3944, U5473);
  and ginst7389 (U3944, U3431, U5472);
  and ginst7390 (U3945, U3946, U5476);
  and ginst7391 (U3946, U3431, U5475);
  and ginst7392 (U3947, U3948, U5479);
  and ginst7393 (U3948, U3431, U5478);
  and ginst7394 (U3949, U3431, U5480, U5482);
  and ginst7395 (U3950, U3431, U5483, U5485);
  and ginst7396 (U3951, U3431, U5486, U5488);
  and ginst7397 (U3952, U3431, U5489, U5491);
  and ginst7398 (U3953, U3431, U5492, U5494);
  and ginst7399 (U3954, U3431, U5495, U5497);
  and ginst7400 (U3955, U3431, U5498, U5500);
  and ginst7401 (U3956, U3431, U5501, U5503);
  and ginst7402 (U3957, U3431, U5504, U5506);
  and ginst7403 (U3958, U3431, U5507, U5509);
  and ginst7404 (U3959, U3431, U5510, U5512);
  and ginst7405 (U3960, U3431, U5513, U5515);
  and ginst7406 (U3961, U3431, U5516, U5518);
  and ginst7407 (U3962, U5805, U5808);
  and ginst7408 (U3963, U3365, U3430);
  and ginst7409 (U3964, U4026, U5616);
  and ginst7410 (U3965, U5676, U5677);
  and ginst7411 (U3966, U5734, U5736);
  not ginst7412 (U3967, IR_REG_31__SCAN_IN);
  nand ginst7413 (U3968, U3023, U3360);
  nand ginst7414 (U3969, U5799, U5802);
  nand ginst7415 (U3970, U3048, U3661);
  nand ginst7416 (U3971, U3048, U3778);
  and ginst7417 (U3972, U6023, U6024);
  and ginst7418 (U3973, U6025, U6026);
  and ginst7419 (U3974, U6027, U6028);
  and ginst7420 (U3975, U6029, U6030);
  and ginst7421 (U3976, U6031, U6032);
  and ginst7422 (U3977, U6033, U6034);
  and ginst7423 (U3978, U6035, U6036);
  and ginst7424 (U3979, U6037, U6038);
  and ginst7425 (U3980, U6039, U6040);
  and ginst7426 (U3981, U6041, U6042);
  and ginst7427 (U3982, U6043, U6044);
  and ginst7428 (U3983, U6045, U6046);
  and ginst7429 (U3984, U6047, U6048);
  and ginst7430 (U3985, U6049, U6050);
  and ginst7431 (U3986, U6051, U6052);
  and ginst7432 (U3987, U6053, U6054);
  and ginst7433 (U3988, U6055, U6056);
  and ginst7434 (U3989, U6057, U6058);
  and ginst7435 (U3990, U6059, U6060);
  and ginst7436 (U3991, U6061, U6062);
  and ginst7437 (U3992, U6063, U6064);
  and ginst7438 (U3993, U6065, U6066);
  and ginst7439 (U3994, U6067, U6068);
  and ginst7440 (U3995, U6069, U6070);
  and ginst7441 (U3996, U6071, U6072);
  and ginst7442 (U3997, U6073, U6074);
  and ginst7443 (U3998, U6075, U6076);
  and ginst7444 (U3999, U6077, U6078);
  and ginst7445 (U4000, U6079, U6080);
  and ginst7446 (U4001, U6081, U6082);
  nand ginst7447 (U4002, U3053, U3777);
  and ginst7448 (U4003, U6083, U6084);
  and ginst7449 (U4004, U6085, U6086);
  not ginst7450 (U4005, R1375_U26);
  and ginst7451 (U4006, U6250, U6251);
  not ginst7452 (U4007, R1347_U13);
  nand ginst7453 (U4008, U4013, U5805);
  not ginst7454 (U4009, R1352_U6);
  not ginst7455 (U4010, U3372);
  not ginst7456 (U4011, U3370);
  not ginst7457 (U4012, U3419);
  not ginst7458 (U4013, U3367);
  not ginst7459 (U4014, U3366);
  not ginst7460 (U4015, U3368);
  not ginst7461 (U4016, U3362);
  not ginst7462 (U4017, U3364);
  not ginst7463 (U4018, U3363);
  not ginst7464 (U4019, U3420);
  not ginst7465 (U4020, U3418);
  not ginst7466 (U4021, U3353);
  not ginst7467 (U4022, U3371);
  not ginst7468 (U4023, U4008);
  not ginst7469 (U4024, U3369);
  nand ginst7470 (U4025, U4042, U4782);
  nand ginst7471 (U4026, U3355, U3962);
  not ginst7472 (U4027, U3969);
  not ginst7473 (U4028, U3427);
  not ginst7474 (U4029, U3412);
  not ginst7475 (U4030, U3410);
  not ginst7476 (U4031, U3408);
  not ginst7477 (U4032, U3406);
  not ginst7478 (U4033, U3404);
  not ginst7479 (U4034, U3402);
  not ginst7480 (U4035, U3400);
  not ginst7481 (U4036, U3398);
  not ginst7482 (U4037, U3396);
  not ginst7483 (U4038, U3416);
  not ginst7484 (U4039, U3415);
  not ginst7485 (U4040, U3414);
  not ginst7486 (U4041, U3423);
  not ginst7487 (U4042, U3373);
  not ginst7488 (U4043, U3422);
  not ginst7489 (U4044, U3417);
  not ginst7490 (U4045, U3971);
  not ginst7491 (U4046, U3970);
  not ginst7492 (U4047, U3968);
  not ginst7493 (U4048, U4002);
  not ginst7494 (U4049, U3428);
  nand ginst7495 (U4050, STATE_REG_SCAN_IN, U3429);
  nand ginst7496 (U4051, U3023, U4020);
  not ginst7497 (U4052, U3426);
  nand ginst7498 (U4053, U3209, U4043);
  not ginst7499 (U4054, U3356);
  not ginst7500 (U4055, U3374);
  not ginst7501 (U4056, U3365);
  not ginst7502 (U4057, U3430);
  not ginst7503 (U4058, U3358);
  not ginst7504 (U4059, U3355);
  nand ginst7505 (U4060, U3047, U3373);
  nand ginst7506 (U4061, U4060, U5748);
  nand ginst7507 (U4062, U3969, U4061);
  not ginst7508 (U4063, U3148);
  not ginst7509 (U4064, U3357);
  nand ginst7510 (U4065, DATAI_0_, U3149);
  nand ginst7511 (U4066, IR_REG_0__SCAN_IN, U3029);
  nand ginst7512 (U4067, IR_REG_0__SCAN_IN, U4064);
  nand ginst7513 (U4068, DATAI_1_, U3149);
  nand ginst7514 (U4069, SUB_84_U48, U3029);
  nand ginst7515 (U4070, IR_REG_1__SCAN_IN, U4064);
  nand ginst7516 (U4071, DATAI_2_, U3149);
  nand ginst7517 (U4072, SUB_84_U20, U3029);
  nand ginst7518 (U4073, IR_REG_2__SCAN_IN, U4064);
  nand ginst7519 (U4074, DATAI_3_, U3149);
  nand ginst7520 (U4075, SUB_84_U21, U3029);
  nand ginst7521 (U4076, IR_REG_3__SCAN_IN, U4064);
  nand ginst7522 (U4077, DATAI_4_, U3149);
  nand ginst7523 (U4078, SUB_84_U70, U3029);
  nand ginst7524 (U4079, IR_REG_4__SCAN_IN, U4064);
  nand ginst7525 (U4080, DATAI_5_, U3149);
  nand ginst7526 (U4081, SUB_84_U22, U3029);
  nand ginst7527 (U4082, IR_REG_5__SCAN_IN, U4064);
  nand ginst7528 (U4083, DATAI_6_, U3149);
  nand ginst7529 (U4084, SUB_84_U23, U3029);
  nand ginst7530 (U4085, IR_REG_6__SCAN_IN, U4064);
  nand ginst7531 (U4086, DATAI_7_, U3149);
  nand ginst7532 (U4087, SUB_84_U24, U3029);
  nand ginst7533 (U4088, IR_REG_7__SCAN_IN, U4064);
  nand ginst7534 (U4089, DATAI_8_, U3149);
  nand ginst7535 (U4090, SUB_84_U68, U3029);
  nand ginst7536 (U4091, IR_REG_8__SCAN_IN, U4064);
  nand ginst7537 (U4092, DATAI_9_, U3149);
  nand ginst7538 (U4093, SUB_84_U25, U3029);
  nand ginst7539 (U4094, IR_REG_9__SCAN_IN, U4064);
  nand ginst7540 (U4095, DATAI_10_, U3149);
  nand ginst7541 (U4096, SUB_84_U6, U3029);
  nand ginst7542 (U4097, IR_REG_10__SCAN_IN, U4064);
  nand ginst7543 (U4098, DATAI_11_, U3149);
  nand ginst7544 (U4099, SUB_84_U7, U3029);
  nand ginst7545 (U4100, IR_REG_11__SCAN_IN, U4064);
  nand ginst7546 (U4101, DATAI_12_, U3149);
  nand ginst7547 (U4102, SUB_84_U89, U3029);
  nand ginst7548 (U4103, IR_REG_12__SCAN_IN, U4064);
  nand ginst7549 (U4104, DATAI_13_, U3149);
  nand ginst7550 (U4105, SUB_84_U8, U3029);
  nand ginst7551 (U4106, IR_REG_13__SCAN_IN, U4064);
  nand ginst7552 (U4107, DATAI_14_, U3149);
  nand ginst7553 (U4108, SUB_84_U9, U3029);
  nand ginst7554 (U4109, IR_REG_14__SCAN_IN, U4064);
  nand ginst7555 (U4110, DATAI_15_, U3149);
  nand ginst7556 (U4111, SUB_84_U10, U3029);
  nand ginst7557 (U4112, IR_REG_15__SCAN_IN, U4064);
  nand ginst7558 (U4113, DATAI_16_, U3149);
  nand ginst7559 (U4114, SUB_84_U87, U3029);
  nand ginst7560 (U4115, IR_REG_16__SCAN_IN, U4064);
  nand ginst7561 (U4116, DATAI_17_, U3149);
  nand ginst7562 (U4117, SUB_84_U11, U3029);
  nand ginst7563 (U4118, IR_REG_17__SCAN_IN, U4064);
  nand ginst7564 (U4119, DATAI_18_, U3149);
  nand ginst7565 (U4120, SUB_84_U12, U3029);
  nand ginst7566 (U4121, IR_REG_18__SCAN_IN, U4064);
  nand ginst7567 (U4122, DATAI_19_, U3149);
  nand ginst7568 (U4123, SUB_84_U13, U3029);
  nand ginst7569 (U4124, IR_REG_19__SCAN_IN, U4064);
  nand ginst7570 (U4125, DATAI_20_, U3149);
  nand ginst7571 (U4126, SUB_84_U83, U3029);
  nand ginst7572 (U4127, IR_REG_20__SCAN_IN, U4064);
  nand ginst7573 (U4128, DATAI_21_, U3149);
  nand ginst7574 (U4129, SUB_84_U14, U3029);
  nand ginst7575 (U4130, IR_REG_21__SCAN_IN, U4064);
  nand ginst7576 (U4131, DATAI_22_, U3149);
  nand ginst7577 (U4132, SUB_84_U15, U3029);
  nand ginst7578 (U4133, IR_REG_22__SCAN_IN, U4064);
  nand ginst7579 (U4134, DATAI_23_, U3149);
  nand ginst7580 (U4135, SUB_84_U81, U3029);
  nand ginst7581 (U4136, IR_REG_23__SCAN_IN, U4064);
  nand ginst7582 (U4137, DATAI_24_, U3149);
  nand ginst7583 (U4138, SUB_84_U78, U3029);
  nand ginst7584 (U4139, IR_REG_24__SCAN_IN, U4064);
  nand ginst7585 (U4140, DATAI_25_, U3149);
  nand ginst7586 (U4141, SUB_84_U16, U3029);
  nand ginst7587 (U4142, IR_REG_25__SCAN_IN, U4064);
  nand ginst7588 (U4143, DATAI_26_, U3149);
  nand ginst7589 (U4144, SUB_84_U17, U3029);
  nand ginst7590 (U4145, IR_REG_26__SCAN_IN, U4064);
  nand ginst7591 (U4146, DATAI_27_, U3149);
  nand ginst7592 (U4147, SUB_84_U76, U3029);
  nand ginst7593 (U4148, IR_REG_27__SCAN_IN, U4064);
  nand ginst7594 (U4149, DATAI_28_, U3149);
  nand ginst7595 (U4150, SUB_84_U18, U3029);
  nand ginst7596 (U4151, IR_REG_28__SCAN_IN, U4064);
  nand ginst7597 (U4152, DATAI_29_, U3149);
  nand ginst7598 (U4153, SUB_84_U19, U3029);
  nand ginst7599 (U4154, IR_REG_29__SCAN_IN, U4064);
  nand ginst7600 (U4155, DATAI_30_, U3149);
  nand ginst7601 (U4156, SUB_84_U73, U3029);
  nand ginst7602 (U4157, IR_REG_30__SCAN_IN, U4064);
  nand ginst7603 (U4158, DATAI_31_, U3149);
  nand ginst7604 (U4159, SUB_84_U49, U3029);
  nand ginst7605 (U4160, IR_REG_31__SCAN_IN, U4064);
  not ginst7606 (U4161, U3360);
  nand ginst7607 (U4162, U3358, U5751);
  nand ginst7608 (U4163, U3358, U5757);
  nand ginst7609 (U4164, D_REG_10__SCAN_IN, U4161);
  nand ginst7610 (U4165, D_REG_11__SCAN_IN, U4161);
  nand ginst7611 (U4166, D_REG_12__SCAN_IN, U4161);
  nand ginst7612 (U4167, D_REG_13__SCAN_IN, U4161);
  nand ginst7613 (U4168, D_REG_14__SCAN_IN, U4161);
  nand ginst7614 (U4169, D_REG_15__SCAN_IN, U4161);
  nand ginst7615 (U4170, D_REG_16__SCAN_IN, U4161);
  nand ginst7616 (U4171, D_REG_17__SCAN_IN, U4161);
  nand ginst7617 (U4172, D_REG_18__SCAN_IN, U4161);
  nand ginst7618 (U4173, D_REG_19__SCAN_IN, U4161);
  nand ginst7619 (U4174, D_REG_20__SCAN_IN, U4161);
  nand ginst7620 (U4175, D_REG_21__SCAN_IN, U4161);
  nand ginst7621 (U4176, D_REG_22__SCAN_IN, U4161);
  nand ginst7622 (U4177, D_REG_23__SCAN_IN, U4161);
  nand ginst7623 (U4178, D_REG_24__SCAN_IN, U4161);
  nand ginst7624 (U4179, D_REG_25__SCAN_IN, U4161);
  nand ginst7625 (U4180, D_REG_26__SCAN_IN, U4161);
  nand ginst7626 (U4181, D_REG_27__SCAN_IN, U4161);
  nand ginst7627 (U4182, D_REG_28__SCAN_IN, U4161);
  nand ginst7628 (U4183, D_REG_29__SCAN_IN, U4161);
  nand ginst7629 (U4184, D_REG_2__SCAN_IN, U4161);
  nand ginst7630 (U4185, D_REG_30__SCAN_IN, U4161);
  nand ginst7631 (U4186, D_REG_31__SCAN_IN, U4161);
  nand ginst7632 (U4187, D_REG_3__SCAN_IN, U4161);
  nand ginst7633 (U4188, D_REG_4__SCAN_IN, U4161);
  nand ginst7634 (U4189, D_REG_5__SCAN_IN, U4161);
  nand ginst7635 (U4190, D_REG_6__SCAN_IN, U4161);
  nand ginst7636 (U4191, D_REG_7__SCAN_IN, U4161);
  nand ginst7637 (U4192, D_REG_8__SCAN_IN, U4161);
  nand ginst7638 (U4193, D_REG_9__SCAN_IN, U4161);
  nand ginst7639 (U4194, U5817, U5820);
  nand ginst7640 (U4195, U3374, U4194, U5830, U5831);
  nand ginst7641 (U4196, REG2_REG_1__SCAN_IN, U3019);
  nand ginst7642 (U4197, REG1_REG_1__SCAN_IN, U3020);
  nand ginst7643 (U4198, REG0_REG_1__SCAN_IN, U3021);
  nand ginst7644 (U4199, REG3_REG_1__SCAN_IN, U3018);
  not ginst7645 (U4200, U3075);
  not ginst7646 (U4201, U3361);
  nand ginst7647 (U4202, R1150_U31, U4016);
  nand ginst7648 (U4203, R1117_U30, U4018);
  nand ginst7649 (U4204, R1138_U108, U4017);
  nand ginst7650 (U4205, R1192_U32, U4014);
  nand ginst7651 (U4206, R1207_U32, U4013);
  nand ginst7652 (U4207, R1171_U108, U4024);
  nand ginst7653 (U4208, R1240_U108, U4022);
  not ginst7654 (U4209, U3375);
  nand ginst7655 (U4210, R1222_U104, U3027);
  nand ginst7656 (U4211, U3026, U3075);
  nand ginst7657 (U4212, U3024, U3464);
  nand ginst7658 (U4213, U3464, U4021);
  nand ginst7659 (U4214, U3649, U4209);
  nand ginst7660 (U4215, REG2_REG_2__SCAN_IN, U3019);
  nand ginst7661 (U4216, REG1_REG_2__SCAN_IN, U3020);
  nand ginst7662 (U4217, REG0_REG_2__SCAN_IN, U3021);
  nand ginst7663 (U4218, REG3_REG_2__SCAN_IN, U3018);
  not ginst7664 (U4219, U3065);
  nand ginst7665 (U4220, REG0_REG_0__SCAN_IN, U3021);
  nand ginst7666 (U4221, REG1_REG_0__SCAN_IN, U3020);
  nand ginst7667 (U4222, REG2_REG_0__SCAN_IN, U3019);
  nand ginst7668 (U4223, REG3_REG_0__SCAN_IN, U3018);
  not ginst7669 (U4224, U3074);
  nand ginst7670 (U4225, U3034, U3074);
  nand ginst7671 (U4226, R1150_U114, U4016);
  nand ginst7672 (U4227, R1117_U113, U4018);
  nand ginst7673 (U4228, R1138_U107, U4017);
  nand ginst7674 (U4229, R1192_U114, U4014);
  nand ginst7675 (U4230, R1207_U114, U4013);
  nand ginst7676 (U4231, R1171_U107, U4024);
  nand ginst7677 (U4232, R1240_U107, U4022);
  not ginst7678 (U4233, U3377);
  nand ginst7679 (U4234, R1222_U103, U3027);
  nand ginst7680 (U4235, U3026, U3065);
  nand ginst7681 (U4236, R1282_U31, U3024);
  nand ginst7682 (U4237, U3468, U4021);
  nand ginst7683 (U4238, U3665, U4233);
  nand ginst7684 (U4239, REG2_REG_3__SCAN_IN, U3019);
  nand ginst7685 (U4240, REG1_REG_3__SCAN_IN, U3020);
  nand ginst7686 (U4241, REG0_REG_3__SCAN_IN, U3021);
  nand ginst7687 (U4242, ADD_95_U4, U3018);
  not ginst7688 (U4243, U3061);
  nand ginst7689 (U4244, U3034, U3075);
  nand ginst7690 (U4245, R1150_U124, U4016);
  nand ginst7691 (U4246, R1117_U123, U4018);
  nand ginst7692 (U4247, R1138_U24, U4017);
  nand ginst7693 (U4248, R1192_U124, U4014);
  nand ginst7694 (U4249, R1207_U124, U4013);
  nand ginst7695 (U4250, R1171_U24, U4024);
  nand ginst7696 (U4251, R1240_U24, U4022);
  not ginst7697 (U4252, U3378);
  nand ginst7698 (U4253, R1222_U23, U3027);
  nand ginst7699 (U4254, U3026, U3061);
  nand ginst7700 (U4255, R1282_U6, U3024);
  nand ginst7701 (U4256, U3470, U4021);
  nand ginst7702 (U4257, U3669, U4252);
  nand ginst7703 (U4258, REG2_REG_4__SCAN_IN, U3019);
  nand ginst7704 (U4259, REG1_REG_4__SCAN_IN, U3020);
  nand ginst7705 (U4260, REG0_REG_4__SCAN_IN, U3021);
  nand ginst7706 (U4261, ADD_95_U51, U3018);
  not ginst7707 (U4262, U3057);
  nand ginst7708 (U4263, U3034, U3065);
  nand ginst7709 (U4264, R1150_U28, U4016);
  nand ginst7710 (U4265, R1117_U27, U4018);
  nand ginst7711 (U4266, R1138_U113, U4017);
  nand ginst7712 (U4267, R1192_U29, U4014);
  nand ginst7713 (U4268, R1207_U29, U4013);
  nand ginst7714 (U4269, R1171_U113, U4024);
  nand ginst7715 (U4270, R1240_U113, U4022);
  not ginst7716 (U4271, U3379);
  nand ginst7717 (U4272, R1222_U109, U3027);
  nand ginst7718 (U4273, U3026, U3057);
  nand ginst7719 (U4274, R1282_U7, U3024);
  nand ginst7720 (U4275, U3472, U4021);
  nand ginst7721 (U4276, U3673, U4271);
  nand ginst7722 (U4277, REG2_REG_5__SCAN_IN, U3019);
  nand ginst7723 (U4278, REG1_REG_5__SCAN_IN, U3020);
  nand ginst7724 (U4279, REG0_REG_5__SCAN_IN, U3021);
  nand ginst7725 (U4280, ADD_95_U50, U3018);
  not ginst7726 (U4281, U3064);
  nand ginst7727 (U4282, U3034, U3061);
  nand ginst7728 (U4283, R1150_U123, U4016);
  nand ginst7729 (U4284, R1117_U122, U4018);
  nand ginst7730 (U4285, R1138_U112, U4017);
  nand ginst7731 (U4286, R1192_U123, U4014);
  nand ginst7732 (U4287, R1207_U123, U4013);
  nand ginst7733 (U4288, R1171_U112, U4024);
  nand ginst7734 (U4289, R1240_U112, U4022);
  not ginst7735 (U4290, U3380);
  nand ginst7736 (U4291, R1222_U108, U3027);
  nand ginst7737 (U4292, U3026, U3064);
  nand ginst7738 (U4293, R1282_U8, U3024);
  nand ginst7739 (U4294, U3474, U4021);
  nand ginst7740 (U4295, U3677, U4290);
  nand ginst7741 (U4296, REG2_REG_6__SCAN_IN, U3019);
  nand ginst7742 (U4297, REG1_REG_6__SCAN_IN, U3020);
  nand ginst7743 (U4298, REG0_REG_6__SCAN_IN, U3021);
  nand ginst7744 (U4299, ADD_95_U49, U3018);
  not ginst7745 (U4300, U3068);
  nand ginst7746 (U4301, U3034, U3057);
  nand ginst7747 (U4302, R1150_U122, U4016);
  nand ginst7748 (U4303, R1117_U121, U4018);
  nand ginst7749 (U4304, R1138_U25, U4017);
  nand ginst7750 (U4305, R1192_U122, U4014);
  nand ginst7751 (U4306, R1207_U122, U4013);
  nand ginst7752 (U4307, R1171_U25, U4024);
  nand ginst7753 (U4308, R1240_U25, U4022);
  not ginst7754 (U4309, U3381);
  nand ginst7755 (U4310, R1222_U24, U3027);
  nand ginst7756 (U4311, U3026, U3068);
  nand ginst7757 (U4312, R1282_U9, U3024);
  nand ginst7758 (U4313, U3476, U4021);
  nand ginst7759 (U4314, U3681, U4309);
  nand ginst7760 (U4315, REG2_REG_7__SCAN_IN, U3019);
  nand ginst7761 (U4316, REG1_REG_7__SCAN_IN, U3020);
  nand ginst7762 (U4317, REG0_REG_7__SCAN_IN, U3021);
  nand ginst7763 (U4318, ADD_95_U48, U3018);
  not ginst7764 (U4319, U3067);
  nand ginst7765 (U4320, U3034, U3064);
  nand ginst7766 (U4321, R1150_U29, U4016);
  nand ginst7767 (U4322, R1117_U28, U4018);
  nand ginst7768 (U4323, R1138_U111, U4017);
  nand ginst7769 (U4324, R1192_U30, U4014);
  nand ginst7770 (U4325, R1207_U30, U4013);
  nand ginst7771 (U4326, R1171_U111, U4024);
  nand ginst7772 (U4327, R1240_U111, U4022);
  not ginst7773 (U4328, U3382);
  nand ginst7774 (U4329, R1222_U107, U3027);
  nand ginst7775 (U4330, U3026, U3067);
  nand ginst7776 (U4331, R1282_U10, U3024);
  nand ginst7777 (U4332, U3478, U4021);
  nand ginst7778 (U4333, U3685, U4328);
  nand ginst7779 (U4334, REG2_REG_8__SCAN_IN, U3019);
  nand ginst7780 (U4335, REG1_REG_8__SCAN_IN, U3020);
  nand ginst7781 (U4336, REG0_REG_8__SCAN_IN, U3021);
  nand ginst7782 (U4337, ADD_95_U47, U3018);
  not ginst7783 (U4338, U3081);
  nand ginst7784 (U4339, U3034, U3068);
  nand ginst7785 (U4340, R1150_U121, U4016);
  nand ginst7786 (U4341, R1117_U120, U4018);
  nand ginst7787 (U4342, R1138_U26, U4017);
  nand ginst7788 (U4343, R1192_U121, U4014);
  nand ginst7789 (U4344, R1207_U121, U4013);
  nand ginst7790 (U4345, R1171_U26, U4024);
  nand ginst7791 (U4346, R1240_U26, U4022);
  not ginst7792 (U4347, U3383);
  nand ginst7793 (U4348, R1222_U25, U3027);
  nand ginst7794 (U4349, U3026, U3081);
  nand ginst7795 (U4350, R1282_U11, U3024);
  nand ginst7796 (U4351, U3480, U4021);
  nand ginst7797 (U4352, U3689, U4347);
  nand ginst7798 (U4353, REG2_REG_9__SCAN_IN, U3019);
  nand ginst7799 (U4354, REG1_REG_9__SCAN_IN, U3020);
  nand ginst7800 (U4355, REG0_REG_9__SCAN_IN, U3021);
  nand ginst7801 (U4356, ADD_95_U46, U3018);
  not ginst7802 (U4357, U3080);
  nand ginst7803 (U4358, U3034, U3067);
  nand ginst7804 (U4359, R1150_U30, U4016);
  nand ginst7805 (U4360, R1117_U29, U4018);
  nand ginst7806 (U4361, R1138_U110, U4017);
  nand ginst7807 (U4362, R1192_U31, U4014);
  nand ginst7808 (U4363, R1207_U31, U4013);
  nand ginst7809 (U4364, R1171_U110, U4024);
  nand ginst7810 (U4365, R1240_U110, U4022);
  not ginst7811 (U4366, U3384);
  nand ginst7812 (U4367, R1222_U106, U3027);
  nand ginst7813 (U4368, U3026, U3080);
  nand ginst7814 (U4369, R1282_U36, U3024);
  nand ginst7815 (U4370, U3482, U4021);
  nand ginst7816 (U4371, U3693, U4366);
  nand ginst7817 (U4372, REG2_REG_10__SCAN_IN, U3019);
  nand ginst7818 (U4373, REG1_REG_10__SCAN_IN, U3020);
  nand ginst7819 (U4374, REG0_REG_10__SCAN_IN, U3021);
  nand ginst7820 (U4375, ADD_95_U70, U3018);
  not ginst7821 (U4376, U3059);
  nand ginst7822 (U4377, U3034, U3081);
  nand ginst7823 (U4378, R1150_U120, U4016);
  nand ginst7824 (U4379, R1117_U119, U4018);
  nand ginst7825 (U4380, R1138_U109, U4017);
  nand ginst7826 (U4381, R1192_U120, U4014);
  nand ginst7827 (U4382, R1207_U120, U4013);
  nand ginst7828 (U4383, R1171_U109, U4024);
  nand ginst7829 (U4384, R1240_U109, U4022);
  not ginst7830 (U4385, U3385);
  nand ginst7831 (U4386, R1222_U105, U3027);
  nand ginst7832 (U4387, U3026, U3059);
  nand ginst7833 (U4388, R1282_U33, U3024);
  nand ginst7834 (U4389, U3484, U4021);
  nand ginst7835 (U4390, U3697, U4385);
  nand ginst7836 (U4391, REG2_REG_11__SCAN_IN, U3019);
  nand ginst7837 (U4392, REG1_REG_11__SCAN_IN, U3020);
  nand ginst7838 (U4393, REG0_REG_11__SCAN_IN, U3021);
  nand ginst7839 (U4394, ADD_95_U69, U3018);
  not ginst7840 (U4395, U3060);
  nand ginst7841 (U4396, U3034, U3080);
  nand ginst7842 (U4397, R1150_U130, U4016);
  nand ginst7843 (U4398, R1117_U129, U4018);
  nand ginst7844 (U4399, R1138_U18, U4017);
  nand ginst7845 (U4400, R1192_U130, U4014);
  nand ginst7846 (U4401, R1207_U130, U4013);
  nand ginst7847 (U4402, R1171_U18, U4024);
  nand ginst7848 (U4403, R1240_U18, U4022);
  not ginst7849 (U4404, U3386);
  nand ginst7850 (U4405, R1222_U17, U3027);
  nand ginst7851 (U4406, U3026, U3060);
  nand ginst7852 (U4407, R1282_U94, U3024);
  nand ginst7853 (U4408, U3486, U4021);
  nand ginst7854 (U4409, U3701, U4404);
  nand ginst7855 (U4410, REG2_REG_12__SCAN_IN, U3019);
  nand ginst7856 (U4411, REG1_REG_12__SCAN_IN, U3020);
  nand ginst7857 (U4412, REG0_REG_12__SCAN_IN, U3021);
  nand ginst7858 (U4413, ADD_95_U68, U3018);
  not ginst7859 (U4414, U3069);
  nand ginst7860 (U4415, U3034, U3059);
  nand ginst7861 (U4416, R1150_U23, U4016);
  nand ginst7862 (U4417, R1117_U23, U4018);
  nand ginst7863 (U4418, R1138_U127, U4017);
  nand ginst7864 (U4419, R1192_U24, U4014);
  nand ginst7865 (U4420, R1207_U24, U4013);
  nand ginst7866 (U4421, R1171_U127, U4024);
  nand ginst7867 (U4422, R1240_U127, U4022);
  not ginst7868 (U4423, U3387);
  nand ginst7869 (U4424, R1222_U123, U3027);
  nand ginst7870 (U4425, U3026, U3069);
  nand ginst7871 (U4426, R1282_U91, U3024);
  nand ginst7872 (U4427, U3488, U4021);
  nand ginst7873 (U4428, U3705, U4423);
  nand ginst7874 (U4429, REG2_REG_13__SCAN_IN, U3019);
  nand ginst7875 (U4430, REG1_REG_13__SCAN_IN, U3020);
  nand ginst7876 (U4431, REG0_REG_13__SCAN_IN, U3021);
  nand ginst7877 (U4432, ADD_95_U67, U3018);
  not ginst7878 (U4433, U3077);
  nand ginst7879 (U4434, U3034, U3060);
  nand ginst7880 (U4435, R1150_U119, U4016);
  nand ginst7881 (U4436, R1117_U118, U4018);
  nand ginst7882 (U4437, R1138_U126, U4017);
  nand ginst7883 (U4438, R1192_U119, U4014);
  nand ginst7884 (U4439, R1207_U119, U4013);
  nand ginst7885 (U4440, R1171_U126, U4024);
  nand ginst7886 (U4441, R1240_U126, U4022);
  not ginst7887 (U4442, U3388);
  nand ginst7888 (U4443, R1222_U122, U3027);
  nand ginst7889 (U4444, U3026, U3077);
  nand ginst7890 (U4445, R1282_U89, U3024);
  nand ginst7891 (U4446, U3490, U4021);
  nand ginst7892 (U4447, U3709, U4442);
  nand ginst7893 (U4448, REG2_REG_14__SCAN_IN, U3019);
  nand ginst7894 (U4449, REG1_REG_14__SCAN_IN, U3020);
  nand ginst7895 (U4450, REG0_REG_14__SCAN_IN, U3021);
  nand ginst7896 (U4451, ADD_95_U66, U3018);
  not ginst7897 (U4452, U3076);
  nand ginst7898 (U4453, U3034, U3069);
  nand ginst7899 (U4454, R1150_U118, U4016);
  nand ginst7900 (U4455, R1117_U117, U4018);
  nand ginst7901 (U4456, R1138_U19, U4017);
  nand ginst7902 (U4457, R1192_U118, U4014);
  nand ginst7903 (U4458, R1207_U118, U4013);
  nand ginst7904 (U4459, R1171_U19, U4024);
  nand ginst7905 (U4460, R1240_U19, U4022);
  not ginst7906 (U4461, U3389);
  nand ginst7907 (U4462, R1222_U18, U3027);
  nand ginst7908 (U4463, U3026, U3076);
  nand ginst7909 (U4464, R1282_U86, U3024);
  nand ginst7910 (U4465, U3492, U4021);
  nand ginst7911 (U4466, U3713, U4461);
  nand ginst7912 (U4467, REG2_REG_15__SCAN_IN, U3019);
  nand ginst7913 (U4468, REG1_REG_15__SCAN_IN, U3020);
  nand ginst7914 (U4469, REG0_REG_15__SCAN_IN, U3021);
  nand ginst7915 (U4470, ADD_95_U65, U3018);
  not ginst7916 (U4471, U3071);
  nand ginst7917 (U4472, U3034, U3077);
  nand ginst7918 (U4473, R1150_U129, U4016);
  nand ginst7919 (U4474, R1117_U128, U4018);
  nand ginst7920 (U4475, R1138_U125, U4017);
  nand ginst7921 (U4476, R1192_U129, U4014);
  nand ginst7922 (U4477, R1207_U129, U4013);
  nand ginst7923 (U4478, R1171_U125, U4024);
  nand ginst7924 (U4479, R1240_U125, U4022);
  not ginst7925 (U4480, U3390);
  nand ginst7926 (U4481, R1222_U121, U3027);
  nand ginst7927 (U4482, U3026, U3071);
  nand ginst7928 (U4483, R1282_U84, U3024);
  nand ginst7929 (U4484, U3494, U4021);
  nand ginst7930 (U4485, U3717, U4480);
  nand ginst7931 (U4486, REG2_REG_16__SCAN_IN, U3019);
  nand ginst7932 (U4487, REG1_REG_16__SCAN_IN, U3020);
  nand ginst7933 (U4488, REG0_REG_16__SCAN_IN, U3021);
  nand ginst7934 (U4489, ADD_95_U64, U3018);
  not ginst7935 (U4490, U3070);
  nand ginst7936 (U4491, U3034, U3076);
  nand ginst7937 (U4492, R1150_U128, U4016);
  nand ginst7938 (U4493, R1117_U127, U4018);
  nand ginst7939 (U4494, R1138_U124, U4017);
  nand ginst7940 (U4495, R1192_U128, U4014);
  nand ginst7941 (U4496, R1207_U128, U4013);
  nand ginst7942 (U4497, R1171_U124, U4024);
  nand ginst7943 (U4498, R1240_U124, U4022);
  not ginst7944 (U4499, U3391);
  nand ginst7945 (U4500, R1222_U120, U3027);
  nand ginst7946 (U4501, U3026, U3070);
  nand ginst7947 (U4502, R1282_U81, U3024);
  nand ginst7948 (U4503, U3496, U4021);
  nand ginst7949 (U4504, U3721, U4499);
  nand ginst7950 (U4505, REG2_REG_17__SCAN_IN, U3019);
  nand ginst7951 (U4506, REG1_REG_17__SCAN_IN, U3020);
  nand ginst7952 (U4507, REG0_REG_17__SCAN_IN, U3021);
  nand ginst7953 (U4508, ADD_95_U63, U3018);
  not ginst7954 (U4509, U3066);
  nand ginst7955 (U4510, U3034, U3071);
  nand ginst7956 (U4511, R1150_U24, U4016);
  nand ginst7957 (U4512, R1117_U24, U4018);
  nand ginst7958 (U4513, R1138_U123, U4017);
  nand ginst7959 (U4514, R1192_U25, U4014);
  nand ginst7960 (U4515, R1207_U25, U4013);
  nand ginst7961 (U4516, R1171_U123, U4024);
  nand ginst7962 (U4517, R1240_U123, U4022);
  not ginst7963 (U4518, U3392);
  nand ginst7964 (U4519, R1222_U119, U3027);
  nand ginst7965 (U4520, U3026, U3066);
  nand ginst7966 (U4521, R1282_U79, U3024);
  nand ginst7967 (U4522, U3498, U4021);
  nand ginst7968 (U4523, U3725, U4518);
  nand ginst7969 (U4524, REG2_REG_18__SCAN_IN, U3019);
  nand ginst7970 (U4525, REG1_REG_18__SCAN_IN, U3020);
  nand ginst7971 (U4526, REG0_REG_18__SCAN_IN, U3021);
  nand ginst7972 (U4527, ADD_95_U62, U3018);
  not ginst7973 (U4528, U3079);
  nand ginst7974 (U4529, U3034, U3070);
  nand ginst7975 (U4530, R1150_U117, U4016);
  nand ginst7976 (U4531, R1117_U116, U4018);
  nand ginst7977 (U4532, R1138_U20, U4017);
  nand ginst7978 (U4533, R1192_U117, U4014);
  nand ginst7979 (U4534, R1207_U117, U4013);
  nand ginst7980 (U4535, R1171_U20, U4024);
  nand ginst7981 (U4536, R1240_U20, U4022);
  not ginst7982 (U4537, U3393);
  nand ginst7983 (U4538, R1222_U19, U3027);
  nand ginst7984 (U4539, U3026, U3079);
  nand ginst7985 (U4540, R1282_U76, U3024);
  nand ginst7986 (U4541, U3500, U4021);
  nand ginst7987 (U4542, U3729, U4537);
  nand ginst7988 (U4543, REG2_REG_19__SCAN_IN, U3019);
  nand ginst7989 (U4544, REG1_REG_19__SCAN_IN, U3020);
  nand ginst7990 (U4545, REG0_REG_19__SCAN_IN, U3021);
  nand ginst7991 (U4546, ADD_95_U61, U3018);
  not ginst7992 (U4547, U3078);
  nand ginst7993 (U4548, U3034, U3066);
  nand ginst7994 (U4549, R1150_U116, U4016);
  nand ginst7995 (U4550, R1117_U115, U4018);
  nand ginst7996 (U4551, R1138_U122, U4017);
  nand ginst7997 (U4552, R1192_U116, U4014);
  nand ginst7998 (U4553, R1207_U116, U4013);
  nand ginst7999 (U4554, R1171_U122, U4024);
  nand ginst8000 (U4555, R1240_U122, U4022);
  not ginst8001 (U4556, U3394);
  nand ginst8002 (U4557, R1222_U118, U3027);
  nand ginst8003 (U4558, U3026, U3078);
  nand ginst8004 (U4559, R1282_U74, U3024);
  nand ginst8005 (U4560, U3502, U4021);
  nand ginst8006 (U4561, U3733, U4556);
  nand ginst8007 (U4562, REG2_REG_20__SCAN_IN, U3019);
  nand ginst8008 (U4563, REG1_REG_20__SCAN_IN, U3020);
  nand ginst8009 (U4564, REG0_REG_20__SCAN_IN, U3021);
  nand ginst8010 (U4565, ADD_95_U60, U3018);
  not ginst8011 (U4566, U3073);
  nand ginst8012 (U4567, U3034, U3079);
  nand ginst8013 (U4568, R1150_U115, U4016);
  nand ginst8014 (U4569, R1117_U114, U4018);
  nand ginst8015 (U4570, R1138_U121, U4017);
  nand ginst8016 (U4571, R1192_U115, U4014);
  nand ginst8017 (U4572, R1207_U115, U4013);
  nand ginst8018 (U4573, R1171_U121, U4024);
  nand ginst8019 (U4574, R1240_U121, U4022);
  not ginst8020 (U4575, U3395);
  nand ginst8021 (U4576, R1222_U117, U3027);
  nand ginst8022 (U4577, U3026, U3073);
  nand ginst8023 (U4578, R1282_U71, U3024);
  nand ginst8024 (U4579, U3504, U4021);
  nand ginst8025 (U4580, U3737, U4575);
  nand ginst8026 (U4581, REG2_REG_21__SCAN_IN, U3019);
  nand ginst8027 (U4582, REG1_REG_21__SCAN_IN, U3020);
  nand ginst8028 (U4583, REG0_REG_21__SCAN_IN, U3021);
  nand ginst8029 (U4584, ADD_95_U59, U3018);
  not ginst8030 (U4585, U3072);
  nand ginst8031 (U4586, U3034, U3078);
  nand ginst8032 (U4587, R1150_U113, U4016);
  nand ginst8033 (U4588, R1117_U112, U4018);
  nand ginst8034 (U4589, R1138_U21, U4017);
  nand ginst8035 (U4590, R1192_U113, U4014);
  nand ginst8036 (U4591, R1207_U113, U4013);
  nand ginst8037 (U4592, R1171_U21, U4024);
  nand ginst8038 (U4593, R1240_U21, U4022);
  not ginst8039 (U4594, U3397);
  nand ginst8040 (U4595, R1222_U20, U3027);
  nand ginst8041 (U4596, U3026, U3072);
  nand ginst8042 (U4597, R1282_U67, U3024);
  nand ginst8043 (U4598, U4021, U4037);
  nand ginst8044 (U4599, U3741, U4594);
  nand ginst8045 (U4600, REG2_REG_22__SCAN_IN, U3019);
  nand ginst8046 (U4601, REG1_REG_22__SCAN_IN, U3020);
  nand ginst8047 (U4602, REG0_REG_22__SCAN_IN, U3021);
  nand ginst8048 (U4603, ADD_95_U58, U3018);
  not ginst8049 (U4604, U3058);
  nand ginst8050 (U4605, U3034, U3073);
  nand ginst8051 (U4606, R1150_U127, U4016);
  nand ginst8052 (U4607, R1117_U126, U4018);
  nand ginst8053 (U4608, R1138_U22, U4017);
  nand ginst8054 (U4609, R1192_U127, U4014);
  nand ginst8055 (U4610, R1207_U127, U4013);
  nand ginst8056 (U4611, R1171_U22, U4024);
  nand ginst8057 (U4612, R1240_U22, U4022);
  not ginst8058 (U4613, U3399);
  nand ginst8059 (U4614, R1222_U21, U3027);
  nand ginst8060 (U4615, U3026, U3058);
  nand ginst8061 (U4616, R1282_U64, U3024);
  nand ginst8062 (U4617, U4021, U4036);
  nand ginst8063 (U4618, U3745, U4613);
  nand ginst8064 (U4619, REG2_REG_23__SCAN_IN, U3019);
  nand ginst8065 (U4620, REG1_REG_23__SCAN_IN, U3020);
  nand ginst8066 (U4621, REG0_REG_23__SCAN_IN, U3021);
  nand ginst8067 (U4622, ADD_95_U57, U3018);
  not ginst8068 (U4623, U3063);
  nand ginst8069 (U4624, U3034, U3072);
  nand ginst8070 (U4625, R1150_U126, U4016);
  nand ginst8071 (U4626, R1117_U125, U4018);
  nand ginst8072 (U4627, R1138_U120, U4017);
  nand ginst8073 (U4628, R1192_U126, U4014);
  nand ginst8074 (U4629, R1207_U126, U4013);
  nand ginst8075 (U4630, R1171_U120, U4024);
  nand ginst8076 (U4631, R1240_U120, U4022);
  not ginst8077 (U4632, U3401);
  nand ginst8078 (U4633, R1222_U116, U3027);
  nand ginst8079 (U4634, U3026, U3063);
  nand ginst8080 (U4635, R1282_U62, U3024);
  nand ginst8081 (U4636, U4021, U4035);
  nand ginst8082 (U4637, U3749, U4632);
  nand ginst8083 (U4638, REG2_REG_24__SCAN_IN, U3019);
  nand ginst8084 (U4639, REG1_REG_24__SCAN_IN, U3020);
  nand ginst8085 (U4640, REG0_REG_24__SCAN_IN, U3021);
  nand ginst8086 (U4641, ADD_95_U56, U3018);
  not ginst8087 (U4642, U3062);
  nand ginst8088 (U4643, U3034, U3058);
  nand ginst8089 (U4644, R1150_U25, U4016);
  nand ginst8090 (U4645, R1117_U25, U4018);
  nand ginst8091 (U4646, R1138_U119, U4017);
  nand ginst8092 (U4647, R1192_U26, U4014);
  nand ginst8093 (U4648, R1207_U26, U4013);
  nand ginst8094 (U4649, R1171_U119, U4024);
  nand ginst8095 (U4650, R1240_U119, U4022);
  not ginst8096 (U4651, U3403);
  nand ginst8097 (U4652, R1222_U115, U3027);
  nand ginst8098 (U4653, U3026, U3062);
  nand ginst8099 (U4654, R1282_U59, U3024);
  nand ginst8100 (U4655, U4021, U4034);
  nand ginst8101 (U4656, U3753, U4651);
  nand ginst8102 (U4657, REG2_REG_25__SCAN_IN, U3019);
  nand ginst8103 (U4658, REG1_REG_25__SCAN_IN, U3020);
  nand ginst8104 (U4659, REG0_REG_25__SCAN_IN, U3021);
  nand ginst8105 (U4660, ADD_95_U55, U3018);
  not ginst8106 (U4661, U3055);
  nand ginst8107 (U4662, U3034, U3063);
  nand ginst8108 (U4663, R1150_U112, U4016);
  nand ginst8109 (U4664, R1117_U111, U4018);
  nand ginst8110 (U4665, R1138_U118, U4017);
  nand ginst8111 (U4666, R1192_U112, U4014);
  nand ginst8112 (U4667, R1207_U112, U4013);
  nand ginst8113 (U4668, R1171_U118, U4024);
  nand ginst8114 (U4669, R1240_U118, U4022);
  not ginst8115 (U4670, U3405);
  nand ginst8116 (U4671, R1222_U114, U3027);
  nand ginst8117 (U4672, U3026, U3055);
  nand ginst8118 (U4673, R1282_U57, U3024);
  nand ginst8119 (U4674, U4021, U4033);
  nand ginst8120 (U4675, U3757, U4670);
  nand ginst8121 (U4676, REG2_REG_26__SCAN_IN, U3019);
  nand ginst8122 (U4677, REG1_REG_26__SCAN_IN, U3020);
  nand ginst8123 (U4678, REG0_REG_26__SCAN_IN, U3021);
  nand ginst8124 (U4679, ADD_95_U54, U3018);
  not ginst8125 (U4680, U3054);
  nand ginst8126 (U4681, U3034, U3062);
  nand ginst8127 (U4682, R1150_U111, U4016);
  nand ginst8128 (U4683, R1117_U110, U4018);
  nand ginst8129 (U4684, R1138_U117, U4017);
  nand ginst8130 (U4685, R1192_U111, U4014);
  nand ginst8131 (U4686, R1207_U111, U4013);
  nand ginst8132 (U4687, R1171_U117, U4024);
  nand ginst8133 (U4688, R1240_U117, U4022);
  not ginst8134 (U4689, U3407);
  nand ginst8135 (U4690, R1222_U113, U3027);
  nand ginst8136 (U4691, U3026, U3054);
  nand ginst8137 (U4692, R1282_U54, U3024);
  nand ginst8138 (U4693, U4021, U4032);
  nand ginst8139 (U4694, U3761, U4689);
  nand ginst8140 (U4695, REG2_REG_27__SCAN_IN, U3019);
  nand ginst8141 (U4696, REG1_REG_27__SCAN_IN, U3020);
  nand ginst8142 (U4697, REG0_REG_27__SCAN_IN, U3021);
  nand ginst8143 (U4698, ADD_95_U53, U3018);
  not ginst8144 (U4699, U3050);
  nand ginst8145 (U4700, U3034, U3055);
  nand ginst8146 (U4701, R1150_U125, U4016);
  nand ginst8147 (U4702, R1117_U124, U4018);
  nand ginst8148 (U4703, R1138_U23, U4017);
  nand ginst8149 (U4704, R1192_U125, U4014);
  nand ginst8150 (U4705, R1207_U125, U4013);
  nand ginst8151 (U4706, R1171_U23, U4024);
  nand ginst8152 (U4707, R1240_U23, U4022);
  not ginst8153 (U4708, U3409);
  nand ginst8154 (U4709, R1222_U22, U3027);
  nand ginst8155 (U4710, U3026, U3050);
  nand ginst8156 (U4711, R1282_U52, U3024);
  nand ginst8157 (U4712, U4021, U4031);
  nand ginst8158 (U4713, U3765, U4708);
  nand ginst8159 (U4714, REG2_REG_28__SCAN_IN, U3019);
  nand ginst8160 (U4715, REG1_REG_28__SCAN_IN, U3020);
  nand ginst8161 (U4716, REG0_REG_28__SCAN_IN, U3021);
  nand ginst8162 (U4717, ADD_95_U52, U3018);
  not ginst8163 (U4718, U3051);
  nand ginst8164 (U4719, U3034, U3054);
  nand ginst8165 (U4720, R1150_U26, U4016);
  nand ginst8166 (U4721, R1117_U31, U4018);
  nand ginst8167 (U4722, R1138_U116, U4017);
  nand ginst8168 (U4723, R1192_U27, U4014);
  nand ginst8169 (U4724, R1207_U27, U4013);
  nand ginst8170 (U4725, R1171_U116, U4024);
  nand ginst8171 (U4726, R1240_U116, U4022);
  not ginst8172 (U4727, U3411);
  nand ginst8173 (U4728, R1222_U112, U3027);
  nand ginst8174 (U4729, U3026, U3051);
  nand ginst8175 (U4730, R1282_U49, U3024);
  nand ginst8176 (U4731, U4021, U4030);
  nand ginst8177 (U4732, U3769, U4727);
  nand ginst8178 (U4733, ADD_95_U5, U3018);
  nand ginst8179 (U4734, REG2_REG_29__SCAN_IN, U3019);
  nand ginst8180 (U4735, REG1_REG_29__SCAN_IN, U3020);
  nand ginst8181 (U4736, REG0_REG_29__SCAN_IN, U3021);
  not ginst8182 (U4737, U3052);
  nand ginst8183 (U4738, U3034, U3050);
  nand ginst8184 (U4739, R1150_U110, U4016);
  nand ginst8185 (U4740, R1117_U109, U4018);
  nand ginst8186 (U4741, R1138_U115, U4017);
  nand ginst8187 (U4742, R1192_U110, U4014);
  nand ginst8188 (U4743, R1207_U110, U4013);
  nand ginst8189 (U4744, R1171_U115, U4024);
  nand ginst8190 (U4745, R1240_U115, U4022);
  not ginst8191 (U4746, U3413);
  nand ginst8192 (U4747, R1222_U111, U3027);
  nand ginst8193 (U4748, U3026, U3052);
  nand ginst8194 (U4749, R1282_U47, U3024);
  nand ginst8195 (U4750, U4021, U4029);
  nand ginst8196 (U4751, U3773, U4746);
  nand ginst8197 (U4752, REG2_REG_30__SCAN_IN, U3019);
  nand ginst8198 (U4753, REG1_REG_30__SCAN_IN, U3020);
  nand ginst8199 (U4754, REG0_REG_30__SCAN_IN, U3021);
  not ginst8200 (U4755, U3056);
  nand ginst8201 (U4756, U3359, U5799);
  nand ginst8202 (U4757, U3969, U4756);
  nand ginst8203 (U4758, U3056, U3774);
  nand ginst8204 (U4759, U3034, U3051);
  nand ginst8205 (U4760, R1150_U27, U4016);
  nand ginst8206 (U4761, R1117_U26, U4018);
  nand ginst8207 (U4762, R1138_U114, U4017);
  nand ginst8208 (U4763, R1192_U28, U4014);
  nand ginst8209 (U4764, R1207_U28, U4013);
  nand ginst8210 (U4765, R1171_U114, U4024);
  nand ginst8211 (U4766, R1240_U114, U4022);
  nand ginst8212 (U4767, U3049, U3838, U5740);
  nand ginst8213 (U4768, R1222_U110, U3027);
  nand ginst8214 (U4769, R1282_U44, U3024);
  nand ginst8215 (U4770, U4021, U4040);
  nand ginst8216 (U4771, U3049, U3775, U3776);
  nand ginst8217 (U4772, REG2_REG_31__SCAN_IN, U3019);
  nand ginst8218 (U4773, REG1_REG_31__SCAN_IN, U3020);
  nand ginst8219 (U4774, REG0_REG_31__SCAN_IN, U3021);
  not ginst8220 (U4775, U3053);
  nand ginst8221 (U4776, R1282_U42, U3024);
  nand ginst8222 (U4777, U4021, U4039);
  nand ginst8223 (U4778, U4002, U4776, U4777);
  nand ginst8224 (U4779, R1282_U39, U3024);
  nand ginst8225 (U4780, U4021, U4038);
  nand ginst8226 (U4781, U4002, U4779, U4780);
  nand ginst8227 (U4782, U5817, U5820);
  nand ginst8228 (U4783, U3017, U3779);
  nand ginst8229 (U4784, U3418, U4783);
  nand ginst8230 (U4785, U3036, U3075);
  nand ginst8231 (U4786, REG3_REG_0__SCAN_IN, U3033);
  nand ginst8232 (U4787, R1222_U104, U3032);
  nand ginst8233 (U4788, U3031, U3464);
  nand ginst8234 (U4789, U3030, U3464);
  nand ginst8235 (U4790, U3036, U3065);
  nand ginst8236 (U4791, REG3_REG_1__SCAN_IN, U3033);
  nand ginst8237 (U4792, R1222_U103, U3032);
  nand ginst8238 (U4793, U3031, U3468);
  nand ginst8239 (U4794, R1282_U31, U3030);
  nand ginst8240 (U4795, U3036, U3061);
  nand ginst8241 (U4796, REG3_REG_2__SCAN_IN, U3033);
  nand ginst8242 (U4797, R1222_U23, U3032);
  nand ginst8243 (U4798, U3031, U3470);
  nand ginst8244 (U4799, R1282_U6, U3030);
  nand ginst8245 (U4800, U3036, U3057);
  nand ginst8246 (U4801, ADD_95_U4, U3033);
  nand ginst8247 (U4802, R1222_U109, U3032);
  nand ginst8248 (U4803, U3031, U3472);
  nand ginst8249 (U4804, R1282_U7, U3030);
  nand ginst8250 (U4805, U3036, U3064);
  nand ginst8251 (U4806, ADD_95_U51, U3033);
  nand ginst8252 (U4807, R1222_U108, U3032);
  nand ginst8253 (U4808, U3031, U3474);
  nand ginst8254 (U4809, R1282_U8, U3030);
  nand ginst8255 (U4810, U3036, U3068);
  nand ginst8256 (U4811, ADD_95_U50, U3033);
  nand ginst8257 (U4812, R1222_U24, U3032);
  nand ginst8258 (U4813, U3031, U3476);
  nand ginst8259 (U4814, R1282_U9, U3030);
  nand ginst8260 (U4815, U3036, U3067);
  nand ginst8261 (U4816, ADD_95_U49, U3033);
  nand ginst8262 (U4817, R1222_U107, U3032);
  nand ginst8263 (U4818, U3031, U3478);
  nand ginst8264 (U4819, R1282_U10, U3030);
  nand ginst8265 (U4820, U3036, U3081);
  nand ginst8266 (U4821, ADD_95_U48, U3033);
  nand ginst8267 (U4822, R1222_U25, U3032);
  nand ginst8268 (U4823, U3031, U3480);
  nand ginst8269 (U4824, R1282_U11, U3030);
  nand ginst8270 (U4825, U3036, U3080);
  nand ginst8271 (U4826, ADD_95_U47, U3033);
  nand ginst8272 (U4827, R1222_U106, U3032);
  nand ginst8273 (U4828, U3031, U3482);
  nand ginst8274 (U4829, R1282_U36, U3030);
  nand ginst8275 (U4830, U3036, U3059);
  nand ginst8276 (U4831, ADD_95_U46, U3033);
  nand ginst8277 (U4832, R1222_U105, U3032);
  nand ginst8278 (U4833, U3031, U3484);
  nand ginst8279 (U4834, R1282_U33, U3030);
  nand ginst8280 (U4835, U3036, U3060);
  nand ginst8281 (U4836, ADD_95_U70, U3033);
  nand ginst8282 (U4837, R1222_U17, U3032);
  nand ginst8283 (U4838, U3031, U3486);
  nand ginst8284 (U4839, R1282_U94, U3030);
  nand ginst8285 (U4840, U3036, U3069);
  nand ginst8286 (U4841, ADD_95_U69, U3033);
  nand ginst8287 (U4842, R1222_U123, U3032);
  nand ginst8288 (U4843, U3031, U3488);
  nand ginst8289 (U4844, R1282_U91, U3030);
  nand ginst8290 (U4845, U3036, U3077);
  nand ginst8291 (U4846, ADD_95_U68, U3033);
  nand ginst8292 (U4847, R1222_U122, U3032);
  nand ginst8293 (U4848, U3031, U3490);
  nand ginst8294 (U4849, R1282_U89, U3030);
  nand ginst8295 (U4850, U3036, U3076);
  nand ginst8296 (U4851, ADD_95_U67, U3033);
  nand ginst8297 (U4852, R1222_U18, U3032);
  nand ginst8298 (U4853, U3031, U3492);
  nand ginst8299 (U4854, R1282_U86, U3030);
  nand ginst8300 (U4855, U3036, U3071);
  nand ginst8301 (U4856, ADD_95_U66, U3033);
  nand ginst8302 (U4857, R1222_U121, U3032);
  nand ginst8303 (U4858, U3031, U3494);
  nand ginst8304 (U4859, R1282_U84, U3030);
  nand ginst8305 (U4860, U3036, U3070);
  nand ginst8306 (U4861, ADD_95_U65, U3033);
  nand ginst8307 (U4862, R1222_U120, U3032);
  nand ginst8308 (U4863, U3031, U3496);
  nand ginst8309 (U4864, R1282_U81, U3030);
  nand ginst8310 (U4865, U3036, U3066);
  nand ginst8311 (U4866, ADD_95_U64, U3033);
  nand ginst8312 (U4867, R1222_U119, U3032);
  nand ginst8313 (U4868, U3031, U3498);
  nand ginst8314 (U4869, R1282_U79, U3030);
  nand ginst8315 (U4870, U3036, U3079);
  nand ginst8316 (U4871, ADD_95_U63, U3033);
  nand ginst8317 (U4872, R1222_U19, U3032);
  nand ginst8318 (U4873, U3031, U3500);
  nand ginst8319 (U4874, R1282_U76, U3030);
  nand ginst8320 (U4875, U3036, U3078);
  nand ginst8321 (U4876, ADD_95_U62, U3033);
  nand ginst8322 (U4877, R1222_U118, U3032);
  nand ginst8323 (U4878, U3031, U3502);
  nand ginst8324 (U4879, R1282_U74, U3030);
  nand ginst8325 (U4880, U3036, U3073);
  nand ginst8326 (U4881, ADD_95_U61, U3033);
  nand ginst8327 (U4882, R1222_U117, U3032);
  nand ginst8328 (U4883, U3031, U3504);
  nand ginst8329 (U4884, R1282_U71, U3030);
  nand ginst8330 (U4885, U3036, U3072);
  nand ginst8331 (U4886, ADD_95_U60, U3033);
  nand ginst8332 (U4887, R1222_U20, U3032);
  nand ginst8333 (U4888, U3031, U4037);
  nand ginst8334 (U4889, R1282_U67, U3030);
  nand ginst8335 (U4890, U3036, U3058);
  nand ginst8336 (U4891, ADD_95_U59, U3033);
  nand ginst8337 (U4892, R1222_U21, U3032);
  nand ginst8338 (U4893, U3031, U4036);
  nand ginst8339 (U4894, R1282_U64, U3030);
  nand ginst8340 (U4895, U3036, U3063);
  nand ginst8341 (U4896, ADD_95_U58, U3033);
  nand ginst8342 (U4897, R1222_U116, U3032);
  nand ginst8343 (U4898, U3031, U4035);
  nand ginst8344 (U4899, R1282_U62, U3030);
  nand ginst8345 (U4900, U3036, U3062);
  nand ginst8346 (U4901, ADD_95_U57, U3033);
  nand ginst8347 (U4902, R1222_U115, U3032);
  nand ginst8348 (U4903, U3031, U4034);
  nand ginst8349 (U4904, R1282_U59, U3030);
  nand ginst8350 (U4905, U3036, U3055);
  nand ginst8351 (U4906, ADD_95_U56, U3033);
  nand ginst8352 (U4907, R1222_U114, U3032);
  nand ginst8353 (U4908, U3031, U4033);
  nand ginst8354 (U4909, R1282_U57, U3030);
  nand ginst8355 (U4910, U3036, U3054);
  nand ginst8356 (U4911, ADD_95_U55, U3033);
  nand ginst8357 (U4912, R1222_U113, U3032);
  nand ginst8358 (U4913, U3031, U4032);
  nand ginst8359 (U4914, R1282_U54, U3030);
  nand ginst8360 (U4915, U3036, U3050);
  nand ginst8361 (U4916, ADD_95_U54, U3033);
  nand ginst8362 (U4917, R1222_U22, U3032);
  nand ginst8363 (U4918, U3031, U4031);
  nand ginst8364 (U4919, R1282_U52, U3030);
  nand ginst8365 (U4920, U3036, U3051);
  nand ginst8366 (U4921, ADD_95_U53, U3033);
  nand ginst8367 (U4922, R1222_U112, U3032);
  nand ginst8368 (U4923, U3031, U4030);
  nand ginst8369 (U4924, R1282_U49, U3030);
  nand ginst8370 (U4925, U3036, U3052);
  nand ginst8371 (U4926, ADD_95_U52, U3033);
  nand ginst8372 (U4927, R1222_U111, U3032);
  nand ginst8373 (U4928, U3031, U4029);
  nand ginst8374 (U4929, R1282_U47, U3030);
  nand ginst8375 (U4930, ADD_95_U5, U3033);
  nand ginst8376 (U4931, R1222_U110, U3032);
  nand ginst8377 (U4932, U3031, U4040);
  nand ginst8378 (U4933, R1282_U44, U3030);
  nand ginst8379 (U4934, U3031, U4039);
  nand ginst8380 (U4935, R1282_U42, U3030);
  nand ginst8381 (U4936, U3031, U4038);
  nand ginst8382 (U4937, R1282_U39, U3030);
  nand ginst8383 (U4938, U3839, U3840, U3842, U3843);
  nand ginst8384 (U4939, R1105_U4, U3042, U3044);
  nand ginst8385 (U4940, U3044, U3844);
  nand ginst8386 (U4941, R1162_U4, U3038, U3044);
  not ginst8387 (U4942, U3421);
  nand ginst8388 (U4943, R1105_U4, U3043);
  nand ginst8389 (U4944, REG3_REG_19__SCAN_IN, U3149);
  nand ginst8390 (U4945, U3041, U3461);
  nand ginst8391 (U4946, R1162_U4, U3039);
  nand ginst8392 (U4947, ADDR_REG_19__SCAN_IN, U4942);
  nand ginst8393 (U4948, R1105_U55, U3042, U3044);
  nand ginst8394 (U4949, U3044, U3849);
  nand ginst8395 (U4950, R1162_U62, U3038, U3044);
  nand ginst8396 (U4951, R1105_U55, U3043);
  nand ginst8397 (U4952, REG3_REG_18__SCAN_IN, U3149);
  nand ginst8398 (U4953, U3041, U3444);
  nand ginst8399 (U4954, R1162_U62, U3039);
  nand ginst8400 (U4955, ADDR_REG_18__SCAN_IN, U4942);
  nand ginst8401 (U4956, R1105_U56, U3042);
  nand ginst8402 (U4957, U3040, U3445);
  nand ginst8403 (U4958, R1162_U63, U3038);
  nand ginst8404 (U4959, U4956, U4957, U4958);
  nand ginst8405 (U4960, U3044, U4959);
  nand ginst8406 (U4961, R1105_U56, U3043);
  nand ginst8407 (U4962, REG3_REG_17__SCAN_IN, U3149);
  nand ginst8408 (U4963, U3041, U3445);
  nand ginst8409 (U4964, R1162_U63, U3039);
  nand ginst8410 (U4965, ADDR_REG_17__SCAN_IN, U4942);
  nand ginst8411 (U4966, R1105_U57, U3042);
  nand ginst8412 (U4967, U3040, U3446);
  nand ginst8413 (U4968, R1162_U64, U3038);
  nand ginst8414 (U4969, U4966, U4967, U4968);
  nand ginst8415 (U4970, U3044, U4969);
  nand ginst8416 (U4971, R1105_U57, U3043);
  nand ginst8417 (U4972, REG3_REG_16__SCAN_IN, U3149);
  nand ginst8418 (U4973, U3041, U3446);
  nand ginst8419 (U4974, R1162_U64, U3039);
  nand ginst8420 (U4975, ADDR_REG_16__SCAN_IN, U4942);
  nand ginst8421 (U4976, R1105_U58, U3042);
  nand ginst8422 (U4977, U3040, U3447);
  nand ginst8423 (U4978, R1162_U65, U3038);
  nand ginst8424 (U4979, U4976, U4977, U4978);
  nand ginst8425 (U4980, U3044, U4979);
  nand ginst8426 (U4981, R1105_U58, U3043);
  nand ginst8427 (U4982, REG3_REG_15__SCAN_IN, U3149);
  nand ginst8428 (U4983, U3041, U3447);
  nand ginst8429 (U4984, R1162_U65, U3039);
  nand ginst8430 (U4985, ADDR_REG_15__SCAN_IN, U4942);
  nand ginst8431 (U4986, R1105_U59, U3042);
  nand ginst8432 (U4987, U3040, U3448);
  nand ginst8433 (U4988, R1162_U66, U3038);
  nand ginst8434 (U4989, U4986, U4987, U4988);
  nand ginst8435 (U4990, U3044, U4989);
  nand ginst8436 (U4991, R1105_U59, U3043);
  nand ginst8437 (U4992, REG3_REG_14__SCAN_IN, U3149);
  nand ginst8438 (U4993, U3041, U3448);
  nand ginst8439 (U4994, R1162_U66, U3039);
  nand ginst8440 (U4995, ADDR_REG_14__SCAN_IN, U4942);
  nand ginst8441 (U4996, R1105_U60, U3042);
  nand ginst8442 (U4997, U3040, U3449);
  nand ginst8443 (U4998, R1162_U67, U3038);
  nand ginst8444 (U4999, U4996, U4997, U4998);
  nand ginst8445 (U5000, U3044, U4999);
  nand ginst8446 (U5001, R1105_U60, U3043);
  nand ginst8447 (U5002, REG3_REG_13__SCAN_IN, U3149);
  nand ginst8448 (U5003, U3041, U3449);
  nand ginst8449 (U5004, R1162_U67, U3039);
  nand ginst8450 (U5005, ADDR_REG_13__SCAN_IN, U4942);
  nand ginst8451 (U5006, R1105_U61, U3042);
  nand ginst8452 (U5007, U3040, U3450);
  nand ginst8453 (U5008, R1162_U68, U3038);
  nand ginst8454 (U5009, U5006, U5007, U5008);
  nand ginst8455 (U5010, U3044, U5009);
  nand ginst8456 (U5011, R1105_U61, U3043);
  nand ginst8457 (U5012, REG3_REG_12__SCAN_IN, U3149);
  nand ginst8458 (U5013, U3041, U3450);
  nand ginst8459 (U5014, R1162_U68, U3039);
  nand ginst8460 (U5015, ADDR_REG_12__SCAN_IN, U4942);
  nand ginst8461 (U5016, R1105_U62, U3042);
  nand ginst8462 (U5017, U3040, U3451);
  nand ginst8463 (U5018, R1162_U69, U3038);
  nand ginst8464 (U5019, U5016, U5017, U5018);
  nand ginst8465 (U5020, U3044, U5019);
  nand ginst8466 (U5021, R1105_U62, U3043);
  nand ginst8467 (U5022, REG3_REG_11__SCAN_IN, U3149);
  nand ginst8468 (U5023, U3041, U3451);
  nand ginst8469 (U5024, R1162_U69, U3039);
  nand ginst8470 (U5025, ADDR_REG_11__SCAN_IN, U4942);
  nand ginst8471 (U5026, R1105_U63, U3042);
  nand ginst8472 (U5027, U3040, U3452);
  nand ginst8473 (U5028, R1162_U70, U3038);
  nand ginst8474 (U5029, U5026, U5027, U5028);
  nand ginst8475 (U5030, U3044, U5029);
  nand ginst8476 (U5031, R1105_U63, U3043);
  nand ginst8477 (U5032, REG3_REG_10__SCAN_IN, U3149);
  nand ginst8478 (U5033, U3041, U3452);
  nand ginst8479 (U5034, R1162_U70, U3039);
  nand ginst8480 (U5035, ADDR_REG_10__SCAN_IN, U4942);
  nand ginst8481 (U5036, R1105_U47, U3042);
  nand ginst8482 (U5037, U3040, U3435);
  nand ginst8483 (U5038, R1162_U54, U3038);
  nand ginst8484 (U5039, U5036, U5037, U5038);
  nand ginst8485 (U5040, U3044, U5039);
  nand ginst8486 (U5041, R1105_U47, U3043);
  nand ginst8487 (U5042, REG3_REG_9__SCAN_IN, U3149);
  nand ginst8488 (U5043, U3041, U3435);
  nand ginst8489 (U5044, R1162_U54, U3039);
  nand ginst8490 (U5045, ADDR_REG_9__SCAN_IN, U4942);
  nand ginst8491 (U5046, R1105_U48, U3042);
  nand ginst8492 (U5047, U3040, U3436);
  nand ginst8493 (U5048, R1162_U55, U3038);
  nand ginst8494 (U5049, U5046, U5047, U5048);
  nand ginst8495 (U5050, U3044, U5049);
  nand ginst8496 (U5051, R1105_U48, U3043);
  nand ginst8497 (U5052, REG3_REG_8__SCAN_IN, U3149);
  nand ginst8498 (U5053, U3041, U3436);
  nand ginst8499 (U5054, R1162_U55, U3039);
  nand ginst8500 (U5055, ADDR_REG_8__SCAN_IN, U4942);
  nand ginst8501 (U5056, R1105_U49, U3042);
  nand ginst8502 (U5057, U3040, U3437);
  nand ginst8503 (U5058, R1162_U56, U3038);
  nand ginst8504 (U5059, U5056, U5057, U5058);
  nand ginst8505 (U5060, U3044, U5059);
  nand ginst8506 (U5061, R1105_U49, U3043);
  nand ginst8507 (U5062, REG3_REG_7__SCAN_IN, U3149);
  nand ginst8508 (U5063, U3041, U3437);
  nand ginst8509 (U5064, R1162_U56, U3039);
  nand ginst8510 (U5065, ADDR_REG_7__SCAN_IN, U4942);
  nand ginst8511 (U5066, R1105_U50, U3042);
  nand ginst8512 (U5067, U3040, U3438);
  nand ginst8513 (U5068, R1162_U57, U3038);
  nand ginst8514 (U5069, U5066, U5067, U5068);
  nand ginst8515 (U5070, U3044, U5069);
  nand ginst8516 (U5071, R1105_U50, U3043);
  nand ginst8517 (U5072, REG3_REG_6__SCAN_IN, U3149);
  nand ginst8518 (U5073, U3041, U3438);
  nand ginst8519 (U5074, R1162_U57, U3039);
  nand ginst8520 (U5075, ADDR_REG_6__SCAN_IN, U4942);
  nand ginst8521 (U5076, R1105_U51, U3042);
  nand ginst8522 (U5077, U3040, U3439);
  nand ginst8523 (U5078, R1162_U58, U3038);
  nand ginst8524 (U5079, U5076, U5077, U5078);
  nand ginst8525 (U5080, U3044, U5079);
  nand ginst8526 (U5081, R1105_U51, U3043);
  nand ginst8527 (U5082, REG3_REG_5__SCAN_IN, U3149);
  nand ginst8528 (U5083, U3041, U3439);
  nand ginst8529 (U5084, R1162_U58, U3039);
  nand ginst8530 (U5085, ADDR_REG_5__SCAN_IN, U4942);
  nand ginst8531 (U5086, R1105_U52, U3042);
  nand ginst8532 (U5087, U3040, U3440);
  nand ginst8533 (U5088, R1162_U59, U3038);
  nand ginst8534 (U5089, U5086, U5087, U5088);
  nand ginst8535 (U5090, U3044, U5089);
  nand ginst8536 (U5091, R1105_U52, U3043);
  nand ginst8537 (U5092, REG3_REG_4__SCAN_IN, U3149);
  nand ginst8538 (U5093, U3041, U3440);
  nand ginst8539 (U5094, R1162_U59, U3039);
  nand ginst8540 (U5095, ADDR_REG_4__SCAN_IN, U4942);
  nand ginst8541 (U5096, R1105_U53, U3042);
  nand ginst8542 (U5097, U3040, U3441);
  nand ginst8543 (U5098, R1162_U60, U3038);
  nand ginst8544 (U5099, U5096, U5097, U5098);
  nand ginst8545 (U5100, U3044, U5099);
  nand ginst8546 (U5101, R1105_U53, U3043);
  nand ginst8547 (U5102, REG3_REG_3__SCAN_IN, U3149);
  nand ginst8548 (U5103, U3041, U3441);
  nand ginst8549 (U5104, R1162_U60, U3039);
  nand ginst8550 (U5105, ADDR_REG_3__SCAN_IN, U4942);
  nand ginst8551 (U5106, R1105_U54, U3042);
  nand ginst8552 (U5107, U3040, U3442);
  nand ginst8553 (U5108, R1162_U61, U3038);
  nand ginst8554 (U5109, U5106, U5107, U5108);
  nand ginst8555 (U5110, U3044, U5109);
  nand ginst8556 (U5111, R1105_U54, U3043);
  nand ginst8557 (U5112, REG3_REG_2__SCAN_IN, U3149);
  nand ginst8558 (U5113, U3041, U3442);
  nand ginst8559 (U5114, R1162_U61, U3039);
  nand ginst8560 (U5115, ADDR_REG_2__SCAN_IN, U4942);
  nand ginst8561 (U5116, R1105_U5, U3042);
  nand ginst8562 (U5117, U3040, U3443);
  nand ginst8563 (U5118, R1162_U5, U3038);
  nand ginst8564 (U5119, U5116, U5117, U5118);
  nand ginst8565 (U5120, U3044, U5119);
  nand ginst8566 (U5121, R1105_U5, U3043);
  nand ginst8567 (U5122, REG3_REG_1__SCAN_IN, U3149);
  nand ginst8568 (U5123, U3041, U3443);
  nand ginst8569 (U5124, R1162_U5, U3039);
  nand ginst8570 (U5125, ADDR_REG_1__SCAN_IN, U4942);
  nand ginst8571 (U5126, R1105_U46, U3042);
  nand ginst8572 (U5127, U3040, U3453);
  nand ginst8573 (U5128, R1162_U53, U3038);
  nand ginst8574 (U5129, U5126, U5127, U5128);
  nand ginst8575 (U5130, U3044, U5129);
  nand ginst8576 (U5131, R1105_U46, U3043);
  nand ginst8577 (U5132, REG3_REG_0__SCAN_IN, U3149);
  nand ginst8578 (U5133, U3041, U3453);
  nand ginst8579 (U5134, R1162_U53, U3039);
  nand ginst8580 (U5135, ADDR_REG_0__SCAN_IN, U4942);
  nand ginst8581 (U5136, U3903, U6256, U6257);
  not ginst8582 (U5137, U3425);
  nand ginst8583 (U5138, U4055, U5137);
  nand ginst8584 (U5139, U4006, U5138);
  nand ginst8585 (U5140, U3424, U4020);
  nand ginst8586 (U5141, U4005, U4012);
  nand ginst8587 (U5142, U3902, U6252, U6253);
  nand ginst8588 (U5143, U3014, U3461, U4005);
  nand ginst8589 (U5144, U3431, U5142);
  nand ginst8590 (U5145, U5143, U5144);
  nand ginst8591 (U5146, R395_U6, U3023, U4041);
  nand ginst8592 (U5147, STATE_REG_SCAN_IN, U5145);
  nand ginst8593 (U5148, B_REG_SCAN_IN, U5136);
  nand ginst8594 (U5149, U3037, U3076);
  nand ginst8595 (U5150, U3035, U3070);
  nand ginst8596 (U5151, ADD_95_U65, U3427);
  nand ginst8597 (U5152, U5149, U5150, U5151);
  nand ginst8598 (U5153, U3362, U3363, U3364);
  nand ginst8599 (U5154, U3366, U3419);
  nand ginst8600 (U5155, U5154, U5805);
  nand ginst8601 (U5156, U5153, U5808);
  nand ginst8602 (U5157, U3369, U3906, U5155, U5156);
  nand ginst8603 (U5158, U3427, U5157);
  not ginst8604 (U5159, U3429);
  nand ginst8605 (U5160, U3496, U5744);
  nand ginst8606 (U5161, ADD_95_U65, U5743);
  nand ginst8607 (U5162, U4049, U5152);
  nand ginst8608 (U5163, R1165_U109, U3028);
  nand ginst8609 (U5164, REG3_REG_15__SCAN_IN, U3149);
  nand ginst8610 (U5165, U3037, U3055);
  nand ginst8611 (U5166, U3035, U3050);
  nand ginst8612 (U5167, ADD_95_U54, U3427);
  nand ginst8613 (U5168, U5165, U5166, U5167);
  nand ginst8614 (U5169, U3427, U4021);
  nand ginst8615 (U5170, U5159, U5169);
  nand ginst8616 (U5171, U4021, U4028);
  nand ginst8617 (U5172, U3418, U5171);
  nand ginst8618 (U5173, U3046, U4031);
  nand ginst8619 (U5174, ADD_95_U54, U3045);
  nand ginst8620 (U5175, U4049, U5168);
  nand ginst8621 (U5176, R1165_U15, U3028);
  nand ginst8622 (U5177, REG3_REG_26__SCAN_IN, U3149);
  nand ginst8623 (U5178, U3037, U3064);
  nand ginst8624 (U5179, U3035, U3067);
  nand ginst8625 (U5180, ADD_95_U49, U3427);
  nand ginst8626 (U5181, U5178, U5179, U5180);
  nand ginst8627 (U5182, U3478, U5744);
  nand ginst8628 (U5183, ADD_95_U49, U5743);
  nand ginst8629 (U5184, U4049, U5181);
  nand ginst8630 (U5185, R1165_U94, U3028);
  nand ginst8631 (U5186, REG3_REG_6__SCAN_IN, U3149);
  nand ginst8632 (U5187, U3037, U3066);
  nand ginst8633 (U5188, U3035, U3078);
  nand ginst8634 (U5189, ADD_95_U62, U3427);
  nand ginst8635 (U5190, U5187, U5188, U5189);
  nand ginst8636 (U5191, U3502, U5744);
  nand ginst8637 (U5192, ADD_95_U62, U5743);
  nand ginst8638 (U5193, U4049, U5190);
  nand ginst8639 (U5194, R1165_U107, U3028);
  nand ginst8640 (U5195, REG3_REG_18__SCAN_IN, U3149);
  nand ginst8641 (U5196, U3037, U3075);
  nand ginst8642 (U5197, U3035, U3061);
  nand ginst8643 (U5198, REG3_REG_2__SCAN_IN, U3427);
  nand ginst8644 (U5199, U5196, U5197, U5198);
  nand ginst8645 (U5200, U3470, U5744);
  nand ginst8646 (U5201, REG3_REG_2__SCAN_IN, U5743);
  nand ginst8647 (U5202, U4049, U5199);
  nand ginst8648 (U5203, R1165_U97, U3028);
  nand ginst8649 (U5204, REG3_REG_2__SCAN_IN, U3149);
  nand ginst8650 (U5205, U3037, U3059);
  nand ginst8651 (U5206, U3035, U3069);
  nand ginst8652 (U5207, ADD_95_U69, U3427);
  nand ginst8653 (U5208, U5205, U5206, U5207);
  nand ginst8654 (U5209, U3488, U5744);
  nand ginst8655 (U5210, ADD_95_U69, U5743);
  nand ginst8656 (U5211, U4049, U5208);
  nand ginst8657 (U5212, R1165_U112, U3028);
  nand ginst8658 (U5213, REG3_REG_11__SCAN_IN, U3149);
  nand ginst8659 (U5214, U3037, U3072);
  nand ginst8660 (U5215, U3035, U3063);
  nand ginst8661 (U5216, ADD_95_U58, U3427);
  nand ginst8662 (U5217, U5214, U5215, U5216);
  nand ginst8663 (U5218, U3046, U4035);
  nand ginst8664 (U5219, ADD_95_U58, U3045);
  nand ginst8665 (U5220, U4049, U5217);
  nand ginst8666 (U5221, R1165_U103, U3028);
  nand ginst8667 (U5222, REG3_REG_22__SCAN_IN, U3149);
  nand ginst8668 (U5223, U3037, U3069);
  nand ginst8669 (U5224, U3035, U3076);
  nand ginst8670 (U5225, ADD_95_U67, U3427);
  nand ginst8671 (U5226, U5223, U5224, U5225);
  nand ginst8672 (U5227, U3492, U5744);
  nand ginst8673 (U5228, ADD_95_U67, U5743);
  nand ginst8674 (U5229, U4049, U5226);
  nand ginst8675 (U5230, R1165_U12, U3028);
  nand ginst8676 (U5231, REG3_REG_13__SCAN_IN, U3149);
  nand ginst8677 (U5232, U3037, U3078);
  nand ginst8678 (U5233, U3035, U3072);
  nand ginst8679 (U5234, ADD_95_U60, U3427);
  nand ginst8680 (U5235, U5232, U5233, U5234);
  nand ginst8681 (U5236, U3046, U4037);
  nand ginst8682 (U5237, ADD_95_U60, U3045);
  nand ginst8683 (U5238, U4049, U5235);
  nand ginst8684 (U5239, R1165_U104, U3028);
  nand ginst8685 (U5240, REG3_REG_20__SCAN_IN, U3149);
  nand ginst8686 (U5241, U3426, U3428);
  nand ginst8687 (U5242, U3427, U5241);
  nand ginst8688 (U5243, U4050, U5242);
  nand ginst8689 (U5244, U3035, U3911);
  nand ginst8690 (U5245, U3464, U5744);
  nand ginst8691 (U5246, REG3_REG_0__SCAN_IN, U5243);
  nand ginst8692 (U5247, R1165_U91, U3028);
  nand ginst8693 (U5248, REG3_REG_0__SCAN_IN, U3149);
  nand ginst8694 (U5249, U3037, U3081);
  nand ginst8695 (U5250, U3035, U3059);
  nand ginst8696 (U5251, ADD_95_U46, U3427);
  nand ginst8697 (U5252, U5249, U5250, U5251);
  nand ginst8698 (U5253, U3484, U5744);
  nand ginst8699 (U5254, ADD_95_U46, U5743);
  nand ginst8700 (U5255, U4049, U5252);
  nand ginst8701 (U5256, R1165_U92, U3028);
  nand ginst8702 (U5257, REG3_REG_9__SCAN_IN, U3149);
  nand ginst8703 (U5258, U3037, U3061);
  nand ginst8704 (U5259, U3035, U3064);
  nand ginst8705 (U5260, ADD_95_U51, U3427);
  nand ginst8706 (U5261, U5258, U5259, U5260);
  nand ginst8707 (U5262, U3474, U5744);
  nand ginst8708 (U5263, ADD_95_U51, U5743);
  nand ginst8709 (U5264, U4049, U5261);
  nand ginst8710 (U5265, R1165_U96, U3028);
  nand ginst8711 (U5266, REG3_REG_4__SCAN_IN, U3149);
  nand ginst8712 (U5267, U3037, U3063);
  nand ginst8713 (U5268, U3035, U3055);
  nand ginst8714 (U5269, ADD_95_U56, U3427);
  nand ginst8715 (U5270, U5267, U5268, U5269);
  nand ginst8716 (U5271, U3046, U4033);
  nand ginst8717 (U5272, ADD_95_U56, U3045);
  nand ginst8718 (U5273, U4049, U5270);
  nand ginst8719 (U5274, R1165_U101, U3028);
  nand ginst8720 (U5275, REG3_REG_24__SCAN_IN, U3149);
  nand ginst8721 (U5276, U3037, U3070);
  nand ginst8722 (U5277, U3035, U3079);
  nand ginst8723 (U5278, ADD_95_U63, U3427);
  nand ginst8724 (U5279, U5276, U5277, U5278);
  nand ginst8725 (U5280, U3500, U5744);
  nand ginst8726 (U5281, ADD_95_U63, U5743);
  nand ginst8727 (U5282, U4049, U5279);
  nand ginst8728 (U5283, R1165_U13, U3028);
  nand ginst8729 (U5284, REG3_REG_17__SCAN_IN, U3149);
  nand ginst8730 (U5285, U3037, U3057);
  nand ginst8731 (U5286, U3035, U3068);
  nand ginst8732 (U5287, ADD_95_U50, U3427);
  nand ginst8733 (U5288, U5285, U5286, U5287);
  nand ginst8734 (U5289, U3476, U5744);
  nand ginst8735 (U5290, ADD_95_U50, U5743);
  nand ginst8736 (U5291, U4049, U5288);
  nand ginst8737 (U5292, R1165_U95, U3028);
  nand ginst8738 (U5293, REG3_REG_5__SCAN_IN, U3149);
  nand ginst8739 (U5294, U3037, U3071);
  nand ginst8740 (U5295, U3035, U3066);
  nand ginst8741 (U5296, ADD_95_U64, U3427);
  nand ginst8742 (U5297, U5294, U5295, U5296);
  nand ginst8743 (U5298, U3498, U5744);
  nand ginst8744 (U5299, ADD_95_U64, U5743);
  nand ginst8745 (U5300, U4049, U5297);
  nand ginst8746 (U5301, R1165_U108, U3028);
  nand ginst8747 (U5302, REG3_REG_16__SCAN_IN, U3149);
  nand ginst8748 (U5303, U3037, U3062);
  nand ginst8749 (U5304, U3035, U3054);
  nand ginst8750 (U5305, ADD_95_U55, U3427);
  nand ginst8751 (U5306, U5303, U5304, U5305);
  nand ginst8752 (U5307, U3046, U4032);
  nand ginst8753 (U5308, ADD_95_U55, U3045);
  nand ginst8754 (U5309, U4049, U5306);
  nand ginst8755 (U5310, R1165_U100, U3028);
  nand ginst8756 (U5311, REG3_REG_25__SCAN_IN, U3149);
  nand ginst8757 (U5312, U3037, U3060);
  nand ginst8758 (U5313, U3035, U3077);
  nand ginst8759 (U5314, ADD_95_U68, U3427);
  nand ginst8760 (U5315, U5312, U5313, U5314);
  nand ginst8761 (U5316, U3490, U5744);
  nand ginst8762 (U5317, ADD_95_U68, U5743);
  nand ginst8763 (U5318, U4049, U5315);
  nand ginst8764 (U5319, R1165_U111, U3028);
  nand ginst8765 (U5320, REG3_REG_12__SCAN_IN, U3149);
  nand ginst8766 (U5321, U3037, U3073);
  nand ginst8767 (U5322, U3035, U3058);
  nand ginst8768 (U5323, ADD_95_U59, U3427);
  nand ginst8769 (U5324, U5321, U5322, U5323);
  nand ginst8770 (U5325, U3046, U4036);
  nand ginst8771 (U5326, ADD_95_U59, U3045);
  nand ginst8772 (U5327, U4049, U5324);
  nand ginst8773 (U5328, R1165_U14, U3028);
  nand ginst8774 (U5329, REG3_REG_21__SCAN_IN, U3149);
  nand ginst8775 (U5330, U3037, U3074);
  nand ginst8776 (U5331, U3035, U3065);
  nand ginst8777 (U5332, REG3_REG_1__SCAN_IN, U3427);
  nand ginst8778 (U5333, U5330, U5331, U5332);
  nand ginst8779 (U5334, U3468, U5744);
  nand ginst8780 (U5335, REG3_REG_1__SCAN_IN, U5743);
  nand ginst8781 (U5336, U4049, U5333);
  nand ginst8782 (U5337, R1165_U105, U3028);
  nand ginst8783 (U5338, REG3_REG_1__SCAN_IN, U3149);
  nand ginst8784 (U5339, U3037, U3067);
  nand ginst8785 (U5340, U3035, U3080);
  nand ginst8786 (U5341, ADD_95_U47, U3427);
  nand ginst8787 (U5342, U5339, U5340, U5341);
  nand ginst8788 (U5343, U3482, U5744);
  nand ginst8789 (U5344, ADD_95_U47, U5743);
  nand ginst8790 (U5345, U4049, U5342);
  nand ginst8791 (U5346, R1165_U93, U3028);
  nand ginst8792 (U5347, REG3_REG_8__SCAN_IN, U3149);
  nand ginst8793 (U5348, U3037, U3050);
  nand ginst8794 (U5349, U3035, U3052);
  nand ginst8795 (U5350, ADD_95_U52, U3427);
  nand ginst8796 (U5351, U5348, U5349, U5350);
  nand ginst8797 (U5352, U3046, U4029);
  nand ginst8798 (U5353, ADD_95_U52, U3045);
  nand ginst8799 (U5354, U4049, U5351);
  nand ginst8800 (U5355, R1165_U98, U3028);
  nand ginst8801 (U5356, REG3_REG_28__SCAN_IN, U3149);
  nand ginst8802 (U5357, U3037, U3079);
  nand ginst8803 (U5358, U3035, U3073);
  nand ginst8804 (U5359, ADD_95_U61, U3427);
  nand ginst8805 (U5360, U5357, U5358, U5359);
  nand ginst8806 (U5361, U3504, U5744);
  nand ginst8807 (U5362, ADD_95_U61, U5743);
  nand ginst8808 (U5363, U4049, U5360);
  nand ginst8809 (U5364, R1165_U106, U3028);
  nand ginst8810 (U5365, REG3_REG_19__SCAN_IN, U3149);
  nand ginst8811 (U5366, U3037, U3065);
  nand ginst8812 (U5367, U3035, U3057);
  nand ginst8813 (U5368, ADD_95_U4, U3427);
  nand ginst8814 (U5369, U5366, U5367, U5368);
  nand ginst8815 (U5370, U3472, U5744);
  nand ginst8816 (U5371, ADD_95_U4, U5743);
  nand ginst8817 (U5372, U4049, U5369);
  nand ginst8818 (U5373, R1165_U16, U3028);
  nand ginst8819 (U5374, REG3_REG_3__SCAN_IN, U3149);
  nand ginst8820 (U5375, U3037, U3080);
  nand ginst8821 (U5376, U3035, U3060);
  nand ginst8822 (U5377, ADD_95_U70, U3427);
  nand ginst8823 (U5378, U5375, U5376, U5377);
  nand ginst8824 (U5379, U3486, U5744);
  nand ginst8825 (U5380, ADD_95_U70, U5743);
  nand ginst8826 (U5381, U4049, U5378);
  nand ginst8827 (U5382, R1165_U113, U3028);
  nand ginst8828 (U5383, REG3_REG_10__SCAN_IN, U3149);
  nand ginst8829 (U5384, U3037, U3058);
  nand ginst8830 (U5385, U3035, U3062);
  nand ginst8831 (U5386, ADD_95_U57, U3427);
  nand ginst8832 (U5387, U5384, U5385, U5386);
  nand ginst8833 (U5388, U3046, U4034);
  nand ginst8834 (U5389, ADD_95_U57, U3045);
  nand ginst8835 (U5390, U4049, U5387);
  nand ginst8836 (U5391, R1165_U102, U3028);
  nand ginst8837 (U5392, REG3_REG_23__SCAN_IN, U3149);
  nand ginst8838 (U5393, U3037, U3077);
  nand ginst8839 (U5394, U3035, U3071);
  nand ginst8840 (U5395, ADD_95_U66, U3427);
  nand ginst8841 (U5396, U5393, U5394, U5395);
  nand ginst8842 (U5397, U3494, U5744);
  nand ginst8843 (U5398, ADD_95_U66, U5743);
  nand ginst8844 (U5399, U4049, U5396);
  nand ginst8845 (U5400, R1165_U110, U3028);
  nand ginst8846 (U5401, REG3_REG_14__SCAN_IN, U3149);
  nand ginst8847 (U5402, U3037, U3054);
  nand ginst8848 (U5403, U3035, U3051);
  nand ginst8849 (U5404, ADD_95_U53, U3427);
  nand ginst8850 (U5405, U5402, U5403, U5404);
  nand ginst8851 (U5406, U3046, U4030);
  nand ginst8852 (U5407, ADD_95_U53, U3045);
  nand ginst8853 (U5408, U4049, U5405);
  nand ginst8854 (U5409, R1165_U99, U3028);
  nand ginst8855 (U5410, REG3_REG_27__SCAN_IN, U3149);
  nand ginst8856 (U5411, U3037, U3068);
  nand ginst8857 (U5412, U3035, U3081);
  nand ginst8858 (U5413, ADD_95_U48, U3427);
  nand ginst8859 (U5414, U5411, U5412, U5413);
  nand ginst8860 (U5415, U3480, U5744);
  nand ginst8861 (U5416, ADD_95_U48, U5743);
  nand ginst8862 (U5417, U4049, U5414);
  nand ginst8863 (U5418, R1165_U17, U3028);
  nand ginst8864 (U5419, REG3_REG_7__SCAN_IN, U3149);
  nand ginst8865 (U5420, U3376, U3455);
  nand ginst8866 (U5421, U3454, U5420);
  nand ginst8867 (U5422, R1165_U91, U3454, U5802);
  nand ginst8868 (U5423, U3014, U3484);
  nand ginst8869 (U5424, U3460, U3582);
  nand ginst8870 (U5425, U3080, U5805);
  nand ginst8871 (U5426, U3014, U3482);
  nand ginst8872 (U5427, U3460, U3583);
  nand ginst8873 (U5428, U3081, U5805);
  nand ginst8874 (U5429, U3014, U3480);
  nand ginst8875 (U5430, U3460, U3584);
  nand ginst8876 (U5431, U3067, U5805);
  nand ginst8877 (U5432, U3014, U3478);
  nand ginst8878 (U5433, U3460, U3585);
  nand ginst8879 (U5434, U3068, U5805);
  nand ginst8880 (U5435, U3014, U3476);
  nand ginst8881 (U5436, U3460, U3586);
  nand ginst8882 (U5437, U3064, U5805);
  nand ginst8883 (U5438, U3014, U3474);
  nand ginst8884 (U5439, U3460, U3587);
  nand ginst8885 (U5440, U3057, U5805);
  nand ginst8886 (U5441, U3460, U3588);
  nand ginst8887 (U5442, U3014, U4038);
  nand ginst8888 (U5443, U3053, U5805);
  nand ginst8889 (U5444, U3460, U3589);
  nand ginst8890 (U5445, U3014, U4039);
  nand ginst8891 (U5446, U3056, U5805);
  nand ginst8892 (U5447, U3014, U3472);
  nand ginst8893 (U5448, U3460, U3590);
  nand ginst8894 (U5449, U3061, U5805);
  nand ginst8895 (U5450, U3460, U3591);
  nand ginst8896 (U5451, U3014, U4040);
  nand ginst8897 (U5452, U3052, U5805);
  nand ginst8898 (U5453, U3460, U3592);
  nand ginst8899 (U5454, U3014, U4029);
  nand ginst8900 (U5455, U3051, U5805);
  nand ginst8901 (U5456, U3460, U3593);
  nand ginst8902 (U5457, U3014, U4030);
  nand ginst8903 (U5458, U3050, U5805);
  nand ginst8904 (U5459, U3460, U3594);
  nand ginst8905 (U5460, U3014, U4031);
  nand ginst8906 (U5461, U3054, U5805);
  nand ginst8907 (U5462, U3460, U3595);
  nand ginst8908 (U5463, U3014, U4032);
  nand ginst8909 (U5464, U3055, U5805);
  nand ginst8910 (U5465, U3460, U3596);
  nand ginst8911 (U5466, U3014, U4033);
  nand ginst8912 (U5467, U3062, U5805);
  nand ginst8913 (U5468, U3460, U3597);
  nand ginst8914 (U5469, U3014, U4034);
  nand ginst8915 (U5470, U3063, U5805);
  nand ginst8916 (U5471, U3460, U3598);
  nand ginst8917 (U5472, U3014, U4035);
  nand ginst8918 (U5473, U3058, U5805);
  nand ginst8919 (U5474, U3460, U3599);
  nand ginst8920 (U5475, U3014, U4036);
  nand ginst8921 (U5476, U3072, U5805);
  nand ginst8922 (U5477, U3460, U3600);
  nand ginst8923 (U5478, U3014, U4037);
  nand ginst8924 (U5479, U3073, U5805);
  nand ginst8925 (U5480, U3014, U3470);
  nand ginst8926 (U5481, U3460, U3601);
  nand ginst8927 (U5482, U3065, U5805);
  nand ginst8928 (U5483, U3014, U3504);
  nand ginst8929 (U5484, U3460, U3602);
  nand ginst8930 (U5485, U3078, U5805);
  nand ginst8931 (U5486, U3014, U3502);
  nand ginst8932 (U5487, U3460, U3603);
  nand ginst8933 (U5488, U3079, U5805);
  nand ginst8934 (U5489, U3014, U3500);
  nand ginst8935 (U5490, U3460, U3604);
  nand ginst8936 (U5491, U3066, U5805);
  nand ginst8937 (U5492, U3014, U3498);
  nand ginst8938 (U5493, U3460, U3605);
  nand ginst8939 (U5494, U3070, U5805);
  nand ginst8940 (U5495, U3014, U3496);
  nand ginst8941 (U5496, U3460, U3606);
  nand ginst8942 (U5497, U3071, U5805);
  nand ginst8943 (U5498, U3014, U3494);
  nand ginst8944 (U5499, U3460, U3607);
  nand ginst8945 (U5500, U3076, U5805);
  nand ginst8946 (U5501, U3014, U3492);
  nand ginst8947 (U5502, U3460, U3608);
  nand ginst8948 (U5503, U3077, U5805);
  nand ginst8949 (U5504, U3014, U3490);
  nand ginst8950 (U5505, U3460, U3609);
  nand ginst8951 (U5506, U3069, U5805);
  nand ginst8952 (U5507, U3014, U3488);
  nand ginst8953 (U5508, U3460, U3610);
  nand ginst8954 (U5509, U3060, U5805);
  nand ginst8955 (U5510, U3014, U3486);
  nand ginst8956 (U5511, U3460, U3611);
  nand ginst8957 (U5512, U3059, U5805);
  nand ginst8958 (U5513, U3014, U3468);
  nand ginst8959 (U5514, U3460, U3612);
  nand ginst8960 (U5515, U3075, U5805);
  nand ginst8961 (U5516, U3014, U3464);
  nand ginst8962 (U5517, U3460, U3613);
  nand ginst8963 (U5518, U3074, U5805);
  nand ginst8964 (U5519, U3361, U3484);
  nand ginst8965 (U5520, U3014, U3080);
  nand ginst8966 (U5521, U3081, U5748);
  nand ginst8967 (U5522, U3361, U3482);
  nand ginst8968 (U5523, U3014, U3081);
  nand ginst8969 (U5524, U3067, U5748);
  nand ginst8970 (U5525, U3361, U3480);
  nand ginst8971 (U5526, U3014, U3067);
  nand ginst8972 (U5527, U3068, U5748);
  nand ginst8973 (U5528, U3361, U3478);
  nand ginst8974 (U5529, U3014, U3068);
  nand ginst8975 (U5530, U3064, U5748);
  nand ginst8976 (U5531, U3361, U3476);
  nand ginst8977 (U5532, U3014, U3064);
  nand ginst8978 (U5533, U3057, U5748);
  nand ginst8979 (U5534, U3361, U3474);
  nand ginst8980 (U5535, U3014, U3057);
  nand ginst8981 (U5536, U3061, U5748);
  nand ginst8982 (U5537, U3361, U4038);
  nand ginst8983 (U5538, U3014, U3053);
  nand ginst8984 (U5539, U3361, U4039);
  nand ginst8985 (U5540, U3014, U3056);
  nand ginst8986 (U5541, U3361, U3472);
  nand ginst8987 (U5542, U3014, U3061);
  nand ginst8988 (U5543, U3065, U5748);
  nand ginst8989 (U5544, U3361, U4040);
  nand ginst8990 (U5545, U3014, U3052);
  nand ginst8991 (U5546, U3051, U5748);
  nand ginst8992 (U5547, U3361, U4029);
  nand ginst8993 (U5548, U3014, U3051);
  nand ginst8994 (U5549, U3050, U5748);
  nand ginst8995 (U5550, U3361, U4030);
  nand ginst8996 (U5551, U3014, U3050);
  nand ginst8997 (U5552, U3054, U5748);
  nand ginst8998 (U5553, U3361, U4031);
  nand ginst8999 (U5554, U3014, U3054);
  nand ginst9000 (U5555, U3055, U5748);
  nand ginst9001 (U5556, U3361, U4032);
  nand ginst9002 (U5557, U3014, U3055);
  nand ginst9003 (U5558, U3062, U5748);
  nand ginst9004 (U5559, U3361, U4033);
  nand ginst9005 (U5560, U3014, U3062);
  nand ginst9006 (U5561, U3063, U5748);
  nand ginst9007 (U5562, U3361, U4034);
  nand ginst9008 (U5563, U3014, U3063);
  nand ginst9009 (U5564, U3058, U5748);
  nand ginst9010 (U5565, U3361, U4035);
  nand ginst9011 (U5566, U3014, U3058);
  nand ginst9012 (U5567, U3072, U5748);
  nand ginst9013 (U5568, U3361, U4036);
  nand ginst9014 (U5569, U3014, U3072);
  nand ginst9015 (U5570, U3073, U5748);
  nand ginst9016 (U5571, U3361, U4037);
  nand ginst9017 (U5572, U3014, U3073);
  nand ginst9018 (U5573, U3078, U5748);
  nand ginst9019 (U5574, U3361, U3470);
  nand ginst9020 (U5575, U3014, U3065);
  nand ginst9021 (U5576, U3075, U5748);
  nand ginst9022 (U5577, U3361, U3504);
  nand ginst9023 (U5578, U3014, U3078);
  nand ginst9024 (U5579, U3079, U5748);
  nand ginst9025 (U5580, U3361, U3502);
  nand ginst9026 (U5581, U3014, U3079);
  nand ginst9027 (U5582, U3066, U5748);
  nand ginst9028 (U5583, U3361, U3500);
  nand ginst9029 (U5584, U3014, U3066);
  nand ginst9030 (U5585, U3070, U5748);
  nand ginst9031 (U5586, U3361, U3498);
  nand ginst9032 (U5587, U3014, U3070);
  nand ginst9033 (U5588, U3071, U5748);
  nand ginst9034 (U5589, U3361, U3496);
  nand ginst9035 (U5590, U3014, U3071);
  nand ginst9036 (U5591, U3076, U5748);
  nand ginst9037 (U5592, U3361, U3494);
  nand ginst9038 (U5593, U3014, U3076);
  nand ginst9039 (U5594, U3077, U5748);
  nand ginst9040 (U5595, U3361, U3492);
  nand ginst9041 (U5596, U3014, U3077);
  nand ginst9042 (U5597, U3069, U5748);
  nand ginst9043 (U5598, U3361, U3490);
  nand ginst9044 (U5599, U3014, U3069);
  nand ginst9045 (U5600, U3060, U5748);
  nand ginst9046 (U5601, U3361, U3488);
  nand ginst9047 (U5602, U3014, U3060);
  nand ginst9048 (U5603, U3059, U5748);
  nand ginst9049 (U5604, U3361, U3486);
  nand ginst9050 (U5605, U3014, U3059);
  nand ginst9051 (U5606, U3080, U5748);
  nand ginst9052 (U5607, U3361, U3468);
  nand ginst9053 (U5608, U3014, U3075);
  nand ginst9054 (U5609, U3074, U5748);
  nand ginst9055 (U5610, U3361, U3464);
  nand ginst9056 (U5611, U3014, U3074);
  nand ginst9057 (U5612, U3963, U4026);
  nand ginst9058 (U5613, U3370, U3419);
  nand ginst9059 (U5614, U3366, U3367, U3368, U3374);
  nand ginst9060 (U5615, U3355, U5614);
  nand ginst9061 (U5616, U3355, U4057);
  nand ginst9062 (U5617, U5615, U5616);
  nand ginst9063 (U5618, U3964, U5615);
  nand ginst9064 (U5619, U3484, U5618);
  nand ginst9065 (U5620, U3022, U3080);
  nand ginst9066 (U5621, U3482, U5618);
  nand ginst9067 (U5622, U3022, U3081);
  nand ginst9068 (U5623, U3480, U5618);
  nand ginst9069 (U5624, U3022, U3067);
  nand ginst9070 (U5625, U3478, U5618);
  nand ginst9071 (U5626, U3022, U3068);
  nand ginst9072 (U5627, U3476, U5618);
  nand ginst9073 (U5628, U3022, U3064);
  nand ginst9074 (U5629, U3474, U5618);
  nand ginst9075 (U5630, U3022, U3057);
  nand ginst9076 (U5631, U3472, U5618);
  nand ginst9077 (U5632, U3022, U3061);
  nand ginst9078 (U5633, U4029, U5618);
  nand ginst9079 (U5634, U3022, U3051);
  nand ginst9080 (U5635, U4030, U5618);
  nand ginst9081 (U5636, U3022, U3050);
  nand ginst9082 (U5637, U4031, U5618);
  nand ginst9083 (U5638, U3022, U3054);
  nand ginst9084 (U5639, U4032, U5618);
  nand ginst9085 (U5640, U3022, U3055);
  nand ginst9086 (U5641, U4033, U5618);
  nand ginst9087 (U5642, U3022, U3062);
  nand ginst9088 (U5643, U4034, U5618);
  nand ginst9089 (U5644, U3022, U3063);
  nand ginst9090 (U5645, U4035, U5618);
  nand ginst9091 (U5646, U3022, U3058);
  nand ginst9092 (U5647, U4036, U5618);
  nand ginst9093 (U5648, U3022, U3072);
  nand ginst9094 (U5649, U4037, U5618);
  nand ginst9095 (U5650, U3022, U3073);
  nand ginst9096 (U5651, U3470, U5618);
  nand ginst9097 (U5652, U3022, U3065);
  nand ginst9098 (U5653, U3504, U5618);
  nand ginst9099 (U5654, U3022, U3078);
  nand ginst9100 (U5655, U3502, U5618);
  nand ginst9101 (U5656, U3022, U3079);
  nand ginst9102 (U5657, U3500, U5618);
  nand ginst9103 (U5658, U3022, U3066);
  nand ginst9104 (U5659, U3498, U5618);
  nand ginst9105 (U5660, U3022, U3070);
  nand ginst9106 (U5661, U3496, U5618);
  nand ginst9107 (U5662, U3022, U3071);
  nand ginst9108 (U5663, U3494, U5618);
  nand ginst9109 (U5664, U3022, U3076);
  nand ginst9110 (U5665, U3492, U5618);
  nand ginst9111 (U5666, U3022, U3077);
  nand ginst9112 (U5667, U3490, U5618);
  nand ginst9113 (U5668, U3022, U3069);
  nand ginst9114 (U5669, U3488, U5618);
  nand ginst9115 (U5670, U3022, U3060);
  nand ginst9116 (U5671, U3486, U5618);
  nand ginst9117 (U5672, U3022, U3059);
  nand ginst9118 (U5673, U3468, U5618);
  nand ginst9119 (U5674, U3022, U3075);
  nand ginst9120 (U5675, U3464, U5618);
  nand ginst9121 (U5676, U3022, U3074);
  nand ginst9122 (U5677, REG1_REG_0__SCAN_IN, U4059);
  nand ginst9123 (U5678, U3022, U3484);
  nand ginst9124 (U5679, U3080, U5617);
  nand ginst9125 (U5680, U3022, U3482);
  nand ginst9126 (U5681, U3081, U5617);
  nand ginst9127 (U5682, U3022, U3480);
  nand ginst9128 (U5683, U3067, U5617);
  nand ginst9129 (U5684, U3022, U3478);
  nand ginst9130 (U5685, U3068, U5617);
  nand ginst9131 (U5686, U3022, U3476);
  nand ginst9132 (U5687, U3064, U5617);
  nand ginst9133 (U5688, U3022, U3474);
  nand ginst9134 (U5689, U3057, U5617);
  nand ginst9135 (U5690, U3022, U3472);
  nand ginst9136 (U5691, U3061, U5617);
  nand ginst9137 (U5692, U3022, U4029);
  nand ginst9138 (U5693, U3051, U5617);
  nand ginst9139 (U5694, U3022, U4030);
  nand ginst9140 (U5695, U3050, U5617);
  nand ginst9141 (U5696, U3022, U4031);
  nand ginst9142 (U5697, U3054, U5617);
  nand ginst9143 (U5698, U3022, U4032);
  nand ginst9144 (U5699, U3055, U5617);
  nand ginst9145 (U5700, U3022, U4033);
  nand ginst9146 (U5701, U3062, U5617);
  nand ginst9147 (U5702, U3022, U4034);
  nand ginst9148 (U5703, U3063, U5617);
  nand ginst9149 (U5704, U3022, U4035);
  nand ginst9150 (U5705, U3058, U5617);
  nand ginst9151 (U5706, U3022, U4036);
  nand ginst9152 (U5707, U3072, U5617);
  nand ginst9153 (U5708, U3022, U4037);
  nand ginst9154 (U5709, U3073, U5617);
  nand ginst9155 (U5710, U3022, U3470);
  nand ginst9156 (U5711, U3065, U5617);
  nand ginst9157 (U5712, U3022, U3504);
  nand ginst9158 (U5713, U3078, U5617);
  nand ginst9159 (U5714, U3022, U3502);
  nand ginst9160 (U5715, U3079, U5617);
  nand ginst9161 (U5716, U3022, U3500);
  nand ginst9162 (U5717, U3066, U5617);
  nand ginst9163 (U5718, U3022, U3498);
  nand ginst9164 (U5719, U3070, U5617);
  nand ginst9165 (U5720, U3022, U3496);
  nand ginst9166 (U5721, U3071, U5617);
  nand ginst9167 (U5722, U3022, U3494);
  nand ginst9168 (U5723, U3076, U5617);
  nand ginst9169 (U5724, U3022, U3492);
  nand ginst9170 (U5725, U3077, U5617);
  nand ginst9171 (U5726, U3022, U3490);
  nand ginst9172 (U5727, U3069, U5617);
  nand ginst9173 (U5728, U3022, U3488);
  nand ginst9174 (U5729, U3060, U5617);
  nand ginst9175 (U5730, U3022, U3486);
  nand ginst9176 (U5731, U3059, U5617);
  nand ginst9177 (U5732, U3022, U3468);
  nand ginst9178 (U5733, U3075, U5617);
  nand ginst9179 (U5734, U3022, U3464);
  nand ginst9180 (U5735, U3074, U5617);
  nand ginst9181 (U5736, U3453, U4059);
  nand ginst9182 (U5737, R1207_U28, U4013);
  nand ginst9183 (U5738, R1192_U28, U4014);
  nand ginst9184 (U5739, R1150_U27, U4016);
  nand ginst9185 (U5740, R1117_U26, U4018);
  nand ginst9186 (U5741, U3427, U4052);
  nand ginst9187 (U5742, U4028, U4052);
  nand ginst9188 (U5743, U4050, U5741);
  nand ginst9189 (U5744, U4051, U5742);
  nand ginst9190 (U5745, U5751, U5754);
  nand ginst9191 (U5746, IR_REG_23__SCAN_IN, U3967);
  nand ginst9192 (U5747, IR_REG_31__SCAN_IN, SUB_84_U81);
  not ginst9193 (U5748, U3431);
  nand ginst9194 (U5749, IR_REG_24__SCAN_IN, U3967);
  nand ginst9195 (U5750, IR_REG_31__SCAN_IN, SUB_84_U78);
  not ginst9196 (U5751, U3434);
  nand ginst9197 (U5752, IR_REG_26__SCAN_IN, U3967);
  nand ginst9198 (U5753, IR_REG_31__SCAN_IN, SUB_84_U17);
  not ginst9199 (U5754, U3432);
  nand ginst9200 (U5755, IR_REG_25__SCAN_IN, U3967);
  nand ginst9201 (U5756, IR_REG_31__SCAN_IN, SUB_84_U16);
  not ginst9202 (U5757, U3433);
  nand ginst9203 (U5758, IR_REG_9__SCAN_IN, U3967);
  nand ginst9204 (U5759, IR_REG_31__SCAN_IN, SUB_84_U25);
  nand ginst9205 (U5760, IR_REG_8__SCAN_IN, U3967);
  nand ginst9206 (U5761, IR_REG_31__SCAN_IN, SUB_84_U68);
  nand ginst9207 (U5762, IR_REG_7__SCAN_IN, U3967);
  nand ginst9208 (U5763, IR_REG_31__SCAN_IN, SUB_84_U24);
  nand ginst9209 (U5764, IR_REG_6__SCAN_IN, U3967);
  nand ginst9210 (U5765, IR_REG_31__SCAN_IN, SUB_84_U23);
  nand ginst9211 (U5766, IR_REG_5__SCAN_IN, U3967);
  nand ginst9212 (U5767, IR_REG_31__SCAN_IN, SUB_84_U22);
  nand ginst9213 (U5768, IR_REG_4__SCAN_IN, U3967);
  nand ginst9214 (U5769, IR_REG_31__SCAN_IN, SUB_84_U70);
  nand ginst9215 (U5770, IR_REG_3__SCAN_IN, U3967);
  nand ginst9216 (U5771, IR_REG_31__SCAN_IN, SUB_84_U21);
  nand ginst9217 (U5772, IR_REG_2__SCAN_IN, U3967);
  nand ginst9218 (U5773, IR_REG_31__SCAN_IN, SUB_84_U20);
  nand ginst9219 (U5774, IR_REG_1__SCAN_IN, U3967);
  nand ginst9220 (U5775, IR_REG_31__SCAN_IN, SUB_84_U48);
  nand ginst9221 (U5776, IR_REG_18__SCAN_IN, U3967);
  nand ginst9222 (U5777, IR_REG_31__SCAN_IN, SUB_84_U12);
  nand ginst9223 (U5778, IR_REG_17__SCAN_IN, U3967);
  nand ginst9224 (U5779, IR_REG_31__SCAN_IN, SUB_84_U11);
  nand ginst9225 (U5780, IR_REG_16__SCAN_IN, U3967);
  nand ginst9226 (U5781, IR_REG_31__SCAN_IN, SUB_84_U87);
  nand ginst9227 (U5782, IR_REG_15__SCAN_IN, U3967);
  nand ginst9228 (U5783, IR_REG_31__SCAN_IN, SUB_84_U10);
  nand ginst9229 (U5784, IR_REG_14__SCAN_IN, U3967);
  nand ginst9230 (U5785, IR_REG_31__SCAN_IN, SUB_84_U9);
  nand ginst9231 (U5786, IR_REG_13__SCAN_IN, U3967);
  nand ginst9232 (U5787, IR_REG_31__SCAN_IN, SUB_84_U8);
  nand ginst9233 (U5788, IR_REG_12__SCAN_IN, U3967);
  nand ginst9234 (U5789, IR_REG_31__SCAN_IN, SUB_84_U89);
  nand ginst9235 (U5790, IR_REG_11__SCAN_IN, U3967);
  nand ginst9236 (U5791, IR_REG_31__SCAN_IN, SUB_84_U7);
  nand ginst9237 (U5792, IR_REG_10__SCAN_IN, U3967);
  nand ginst9238 (U5793, IR_REG_31__SCAN_IN, SUB_84_U6);
  nand ginst9239 (U5794, IR_REG_0__SCAN_IN, U3967);
  nand ginst9240 (U5795, IR_REG_0__SCAN_IN, IR_REG_31__SCAN_IN);
  not ginst9241 (U5796, U3453);
  nand ginst9242 (U5797, IR_REG_28__SCAN_IN, U3967);
  nand ginst9243 (U5798, IR_REG_31__SCAN_IN, SUB_84_U18);
  not ginst9244 (U5799, U3454);
  nand ginst9245 (U5800, IR_REG_27__SCAN_IN, U3967);
  nand ginst9246 (U5801, IR_REG_31__SCAN_IN, SUB_84_U76);
  not ginst9247 (U5802, U3455);
  nand ginst9248 (U5803, IR_REG_22__SCAN_IN, U3967);
  nand ginst9249 (U5804, IR_REG_31__SCAN_IN, SUB_84_U15);
  not ginst9250 (U5805, U3456);
  nand ginst9251 (U5806, IR_REG_21__SCAN_IN, U3967);
  nand ginst9252 (U5807, IR_REG_31__SCAN_IN, SUB_84_U14);
  not ginst9253 (U5808, U3457);
  nand ginst9254 (U5809, U3359, U3434);
  nand ginst9255 (U5810, B_REG_SCAN_IN, U4058, U5751);
  nand ginst9256 (U5811, D_REG_0__SCAN_IN, U3968);
  nand ginst9257 (U5812, U4047, U4162);
  nand ginst9258 (U5813, D_REG_1__SCAN_IN, U3968);
  nand ginst9259 (U5814, U4047, U4163);
  nand ginst9260 (U5815, IR_REG_19__SCAN_IN, U3967);
  nand ginst9261 (U5816, IR_REG_31__SCAN_IN, SUB_84_U13);
  not ginst9262 (U5817, U3461);
  nand ginst9263 (U5818, IR_REG_20__SCAN_IN, U3967);
  nand ginst9264 (U5819, IR_REG_31__SCAN_IN, SUB_84_U83);
  not ginst9265 (U5820, U3460);
  nand ginst9266 (U5821, IR_REG_30__SCAN_IN, U3967);
  nand ginst9267 (U5822, IR_REG_31__SCAN_IN, SUB_84_U73);
  not ginst9268 (U5823, U3462);
  nand ginst9269 (U5824, IR_REG_29__SCAN_IN, U3967);
  nand ginst9270 (U5825, IR_REG_31__SCAN_IN, SUB_84_U19);
  not ginst9271 (U5826, U3463);
  nand ginst9272 (U5827, DATAI_0_, U3969);
  nand ginst9273 (U5828, U3453, U4027);
  not ginst9274 (U5829, U3464);
  nand ginst9275 (U5830, U3456, U5808);
  nand ginst9276 (U5831, U3457, U5805);
  nand ginst9277 (U5832, D_REG_1__SCAN_IN, U4161);
  nand ginst9278 (U5833, U3360, U4163);
  not ginst9279 (U5834, U3466);
  nand ginst9280 (U5835, U3360, U5745);
  nand ginst9281 (U5836, D_REG_0__SCAN_IN, U4161);
  not ginst9282 (U5837, U3465);
  nand ginst9283 (U5838, REG0_REG_0__SCAN_IN, U3970);
  nand ginst9284 (U5839, U4046, U4214);
  nand ginst9285 (U5840, DATAI_1_, U3969);
  nand ginst9286 (U5841, U3443, U4027);
  not ginst9287 (U5842, U3468);
  nand ginst9288 (U5843, REG0_REG_1__SCAN_IN, U3970);
  nand ginst9289 (U5844, U4046, U4238);
  nand ginst9290 (U5845, DATAI_2_, U3969);
  nand ginst9291 (U5846, U3442, U4027);
  not ginst9292 (U5847, U3470);
  nand ginst9293 (U5848, REG0_REG_2__SCAN_IN, U3970);
  nand ginst9294 (U5849, U4046, U4257);
  nand ginst9295 (U5850, DATAI_3_, U3969);
  nand ginst9296 (U5851, U3441, U4027);
  not ginst9297 (U5852, U3472);
  nand ginst9298 (U5853, REG0_REG_3__SCAN_IN, U3970);
  nand ginst9299 (U5854, U4046, U4276);
  nand ginst9300 (U5855, DATAI_4_, U3969);
  nand ginst9301 (U5856, U3440, U4027);
  not ginst9302 (U5857, U3474);
  nand ginst9303 (U5858, REG0_REG_4__SCAN_IN, U3970);
  nand ginst9304 (U5859, U4046, U4295);
  nand ginst9305 (U5860, DATAI_5_, U3969);
  nand ginst9306 (U5861, U3439, U4027);
  not ginst9307 (U5862, U3476);
  nand ginst9308 (U5863, REG0_REG_5__SCAN_IN, U3970);
  nand ginst9309 (U5864, U4046, U4314);
  nand ginst9310 (U5865, DATAI_6_, U3969);
  nand ginst9311 (U5866, U3438, U4027);
  not ginst9312 (U5867, U3478);
  nand ginst9313 (U5868, REG0_REG_6__SCAN_IN, U3970);
  nand ginst9314 (U5869, U4046, U4333);
  nand ginst9315 (U5870, DATAI_7_, U3969);
  nand ginst9316 (U5871, U3437, U4027);
  not ginst9317 (U5872, U3480);
  nand ginst9318 (U5873, REG0_REG_7__SCAN_IN, U3970);
  nand ginst9319 (U5874, U4046, U4352);
  nand ginst9320 (U5875, DATAI_8_, U3969);
  nand ginst9321 (U5876, U3436, U4027);
  not ginst9322 (U5877, U3482);
  nand ginst9323 (U5878, REG0_REG_8__SCAN_IN, U3970);
  nand ginst9324 (U5879, U4046, U4371);
  nand ginst9325 (U5880, DATAI_9_, U3969);
  nand ginst9326 (U5881, U3435, U4027);
  not ginst9327 (U5882, U3484);
  nand ginst9328 (U5883, REG0_REG_9__SCAN_IN, U3970);
  nand ginst9329 (U5884, U4046, U4390);
  nand ginst9330 (U5885, DATAI_10_, U3969);
  nand ginst9331 (U5886, U3452, U4027);
  not ginst9332 (U5887, U3486);
  nand ginst9333 (U5888, REG0_REG_10__SCAN_IN, U3970);
  nand ginst9334 (U5889, U4046, U4409);
  nand ginst9335 (U5890, DATAI_11_, U3969);
  nand ginst9336 (U5891, U3451, U4027);
  not ginst9337 (U5892, U3488);
  nand ginst9338 (U5893, REG0_REG_11__SCAN_IN, U3970);
  nand ginst9339 (U5894, U4046, U4428);
  nand ginst9340 (U5895, DATAI_12_, U3969);
  nand ginst9341 (U5896, U3450, U4027);
  not ginst9342 (U5897, U3490);
  nand ginst9343 (U5898, REG0_REG_12__SCAN_IN, U3970);
  nand ginst9344 (U5899, U4046, U4447);
  nand ginst9345 (U5900, DATAI_13_, U3969);
  nand ginst9346 (U5901, U3449, U4027);
  not ginst9347 (U5902, U3492);
  nand ginst9348 (U5903, REG0_REG_13__SCAN_IN, U3970);
  nand ginst9349 (U5904, U4046, U4466);
  nand ginst9350 (U5905, DATAI_14_, U3969);
  nand ginst9351 (U5906, U3448, U4027);
  not ginst9352 (U5907, U3494);
  nand ginst9353 (U5908, REG0_REG_14__SCAN_IN, U3970);
  nand ginst9354 (U5909, U4046, U4485);
  nand ginst9355 (U5910, DATAI_15_, U3969);
  nand ginst9356 (U5911, U3447, U4027);
  not ginst9357 (U5912, U3496);
  nand ginst9358 (U5913, REG0_REG_15__SCAN_IN, U3970);
  nand ginst9359 (U5914, U4046, U4504);
  nand ginst9360 (U5915, DATAI_16_, U3969);
  nand ginst9361 (U5916, U3446, U4027);
  not ginst9362 (U5917, U3498);
  nand ginst9363 (U5918, REG0_REG_16__SCAN_IN, U3970);
  nand ginst9364 (U5919, U4046, U4523);
  nand ginst9365 (U5920, DATAI_17_, U3969);
  nand ginst9366 (U5921, U3445, U4027);
  not ginst9367 (U5922, U3500);
  nand ginst9368 (U5923, REG0_REG_17__SCAN_IN, U3970);
  nand ginst9369 (U5924, U4046, U4542);
  nand ginst9370 (U5925, DATAI_18_, U3969);
  nand ginst9371 (U5926, U3444, U4027);
  not ginst9372 (U5927, U3502);
  nand ginst9373 (U5928, REG0_REG_18__SCAN_IN, U3970);
  nand ginst9374 (U5929, U4046, U4561);
  nand ginst9375 (U5930, DATAI_19_, U3969);
  nand ginst9376 (U5931, U3461, U4027);
  not ginst9377 (U5932, U3504);
  nand ginst9378 (U5933, REG0_REG_19__SCAN_IN, U3970);
  nand ginst9379 (U5934, U4046, U4580);
  nand ginst9380 (U5935, REG0_REG_20__SCAN_IN, U3970);
  nand ginst9381 (U5936, U4046, U4599);
  nand ginst9382 (U5937, REG0_REG_21__SCAN_IN, U3970);
  nand ginst9383 (U5938, U4046, U4618);
  nand ginst9384 (U5939, REG0_REG_22__SCAN_IN, U3970);
  nand ginst9385 (U5940, U4046, U4637);
  nand ginst9386 (U5941, REG0_REG_23__SCAN_IN, U3970);
  nand ginst9387 (U5942, U4046, U4656);
  nand ginst9388 (U5943, REG0_REG_24__SCAN_IN, U3970);
  nand ginst9389 (U5944, U4046, U4675);
  nand ginst9390 (U5945, REG0_REG_25__SCAN_IN, U3970);
  nand ginst9391 (U5946, U4046, U4694);
  nand ginst9392 (U5947, REG0_REG_26__SCAN_IN, U3970);
  nand ginst9393 (U5948, U4046, U4713);
  nand ginst9394 (U5949, REG0_REG_27__SCAN_IN, U3970);
  nand ginst9395 (U5950, U4046, U4732);
  nand ginst9396 (U5951, REG0_REG_28__SCAN_IN, U3970);
  nand ginst9397 (U5952, U4046, U4751);
  nand ginst9398 (U5953, REG0_REG_29__SCAN_IN, U3970);
  nand ginst9399 (U5954, U4046, U4771);
  nand ginst9400 (U5955, REG0_REG_30__SCAN_IN, U3970);
  nand ginst9401 (U5956, U4046, U4778);
  nand ginst9402 (U5957, REG0_REG_31__SCAN_IN, U3970);
  nand ginst9403 (U5958, U4046, U4781);
  nand ginst9404 (U5959, REG1_REG_0__SCAN_IN, U3971);
  nand ginst9405 (U5960, U4045, U4214);
  nand ginst9406 (U5961, REG1_REG_1__SCAN_IN, U3971);
  nand ginst9407 (U5962, U4045, U4238);
  nand ginst9408 (U5963, REG1_REG_2__SCAN_IN, U3971);
  nand ginst9409 (U5964, U4045, U4257);
  nand ginst9410 (U5965, REG1_REG_3__SCAN_IN, U3971);
  nand ginst9411 (U5966, U4045, U4276);
  nand ginst9412 (U5967, REG1_REG_4__SCAN_IN, U3971);
  nand ginst9413 (U5968, U4045, U4295);
  nand ginst9414 (U5969, REG1_REG_5__SCAN_IN, U3971);
  nand ginst9415 (U5970, U4045, U4314);
  nand ginst9416 (U5971, REG1_REG_6__SCAN_IN, U3971);
  nand ginst9417 (U5972, U4045, U4333);
  nand ginst9418 (U5973, REG1_REG_7__SCAN_IN, U3971);
  nand ginst9419 (U5974, U4045, U4352);
  nand ginst9420 (U5975, REG1_REG_8__SCAN_IN, U3971);
  nand ginst9421 (U5976, U4045, U4371);
  nand ginst9422 (U5977, REG1_REG_9__SCAN_IN, U3971);
  nand ginst9423 (U5978, U4045, U4390);
  nand ginst9424 (U5979, REG1_REG_10__SCAN_IN, U3971);
  nand ginst9425 (U5980, U4045, U4409);
  nand ginst9426 (U5981, REG1_REG_11__SCAN_IN, U3971);
  nand ginst9427 (U5982, U4045, U4428);
  nand ginst9428 (U5983, REG1_REG_12__SCAN_IN, U3971);
  nand ginst9429 (U5984, U4045, U4447);
  nand ginst9430 (U5985, REG1_REG_13__SCAN_IN, U3971);
  nand ginst9431 (U5986, U4045, U4466);
  nand ginst9432 (U5987, REG1_REG_14__SCAN_IN, U3971);
  nand ginst9433 (U5988, U4045, U4485);
  nand ginst9434 (U5989, REG1_REG_15__SCAN_IN, U3971);
  nand ginst9435 (U5990, U4045, U4504);
  nand ginst9436 (U5991, REG1_REG_16__SCAN_IN, U3971);
  nand ginst9437 (U5992, U4045, U4523);
  nand ginst9438 (U5993, REG1_REG_17__SCAN_IN, U3971);
  nand ginst9439 (U5994, U4045, U4542);
  nand ginst9440 (U5995, REG1_REG_18__SCAN_IN, U3971);
  nand ginst9441 (U5996, U4045, U4561);
  nand ginst9442 (U5997, REG1_REG_19__SCAN_IN, U3971);
  nand ginst9443 (U5998, U4045, U4580);
  nand ginst9444 (U5999, REG1_REG_20__SCAN_IN, U3971);
  nand ginst9445 (U6000, U4045, U4599);
  nand ginst9446 (U6001, REG1_REG_21__SCAN_IN, U3971);
  nand ginst9447 (U6002, U4045, U4618);
  nand ginst9448 (U6003, REG1_REG_22__SCAN_IN, U3971);
  nand ginst9449 (U6004, U4045, U4637);
  nand ginst9450 (U6005, REG1_REG_23__SCAN_IN, U3971);
  nand ginst9451 (U6006, U4045, U4656);
  nand ginst9452 (U6007, REG1_REG_24__SCAN_IN, U3971);
  nand ginst9453 (U6008, U4045, U4675);
  nand ginst9454 (U6009, REG1_REG_25__SCAN_IN, U3971);
  nand ginst9455 (U6010, U4045, U4694);
  nand ginst9456 (U6011, REG1_REG_26__SCAN_IN, U3971);
  nand ginst9457 (U6012, U4045, U4713);
  nand ginst9458 (U6013, REG1_REG_27__SCAN_IN, U3971);
  nand ginst9459 (U6014, U4045, U4732);
  nand ginst9460 (U6015, REG1_REG_28__SCAN_IN, U3971);
  nand ginst9461 (U6016, U4045, U4751);
  nand ginst9462 (U6017, REG1_REG_29__SCAN_IN, U3971);
  nand ginst9463 (U6018, U4045, U4771);
  nand ginst9464 (U6019, REG1_REG_30__SCAN_IN, U3971);
  nand ginst9465 (U6020, U4045, U4778);
  nand ginst9466 (U6021, REG1_REG_31__SCAN_IN, U3971);
  nand ginst9467 (U6022, U4045, U4781);
  nand ginst9468 (U6023, REG2_REG_0__SCAN_IN, U3417);
  nand ginst9469 (U6024, U3375, U4044);
  nand ginst9470 (U6025, REG2_REG_1__SCAN_IN, U3417);
  nand ginst9471 (U6026, U3377, U4044);
  nand ginst9472 (U6027, REG2_REG_2__SCAN_IN, U3417);
  nand ginst9473 (U6028, U3378, U4044);
  nand ginst9474 (U6029, REG2_REG_3__SCAN_IN, U3417);
  nand ginst9475 (U6030, U3379, U4044);
  nand ginst9476 (U6031, REG2_REG_4__SCAN_IN, U3417);
  nand ginst9477 (U6032, U3380, U4044);
  nand ginst9478 (U6033, REG2_REG_5__SCAN_IN, U3417);
  nand ginst9479 (U6034, U3381, U4044);
  nand ginst9480 (U6035, REG2_REG_6__SCAN_IN, U3417);
  nand ginst9481 (U6036, U3382, U4044);
  nand ginst9482 (U6037, REG2_REG_7__SCAN_IN, U3417);
  nand ginst9483 (U6038, U3383, U4044);
  nand ginst9484 (U6039, REG2_REG_8__SCAN_IN, U3417);
  nand ginst9485 (U6040, U3384, U4044);
  nand ginst9486 (U6041, REG2_REG_9__SCAN_IN, U3417);
  nand ginst9487 (U6042, U3385, U4044);
  nand ginst9488 (U6043, REG2_REG_10__SCAN_IN, U3417);
  nand ginst9489 (U6044, U3386, U4044);
  nand ginst9490 (U6045, REG2_REG_11__SCAN_IN, U3417);
  nand ginst9491 (U6046, U3387, U4044);
  nand ginst9492 (U6047, REG2_REG_12__SCAN_IN, U3417);
  nand ginst9493 (U6048, U3388, U4044);
  nand ginst9494 (U6049, REG2_REG_13__SCAN_IN, U3417);
  nand ginst9495 (U6050, U3389, U4044);
  nand ginst9496 (U6051, REG2_REG_14__SCAN_IN, U3417);
  nand ginst9497 (U6052, U3390, U4044);
  nand ginst9498 (U6053, REG2_REG_15__SCAN_IN, U3417);
  nand ginst9499 (U6054, U3391, U4044);
  nand ginst9500 (U6055, REG2_REG_16__SCAN_IN, U3417);
  nand ginst9501 (U6056, U3392, U4044);
  nand ginst9502 (U6057, REG2_REG_17__SCAN_IN, U3417);
  nand ginst9503 (U6058, U3393, U4044);
  nand ginst9504 (U6059, REG2_REG_18__SCAN_IN, U3417);
  nand ginst9505 (U6060, U3394, U4044);
  nand ginst9506 (U6061, REG2_REG_19__SCAN_IN, U3417);
  nand ginst9507 (U6062, U3395, U4044);
  nand ginst9508 (U6063, REG2_REG_20__SCAN_IN, U3417);
  nand ginst9509 (U6064, U3397, U4044);
  nand ginst9510 (U6065, REG2_REG_21__SCAN_IN, U3417);
  nand ginst9511 (U6066, U3399, U4044);
  nand ginst9512 (U6067, REG2_REG_22__SCAN_IN, U3417);
  nand ginst9513 (U6068, U3401, U4044);
  nand ginst9514 (U6069, REG2_REG_23__SCAN_IN, U3417);
  nand ginst9515 (U6070, U3403, U4044);
  nand ginst9516 (U6071, REG2_REG_24__SCAN_IN, U3417);
  nand ginst9517 (U6072, U3405, U4044);
  nand ginst9518 (U6073, REG2_REG_25__SCAN_IN, U3417);
  nand ginst9519 (U6074, U3407, U4044);
  nand ginst9520 (U6075, REG2_REG_26__SCAN_IN, U3417);
  nand ginst9521 (U6076, U3409, U4044);
  nand ginst9522 (U6077, REG2_REG_27__SCAN_IN, U3417);
  nand ginst9523 (U6078, U3411, U4044);
  nand ginst9524 (U6079, REG2_REG_28__SCAN_IN, U3417);
  nand ginst9525 (U6080, U3413, U4044);
  nand ginst9526 (U6081, REG2_REG_29__SCAN_IN, U3417);
  nand ginst9527 (U6082, U4044, U4767);
  nand ginst9528 (U6083, REG2_REG_30__SCAN_IN, U3417);
  nand ginst9529 (U6084, U4044, U4048);
  nand ginst9530 (U6085, REG2_REG_31__SCAN_IN, U3417);
  nand ginst9531 (U6086, U4044, U4048);
  nand ginst9532 (U6087, DATAO_REG_0__SCAN_IN, U3422);
  nand ginst9533 (U6088, U3074, U4043);
  nand ginst9534 (U6089, DATAO_REG_1__SCAN_IN, U3422);
  nand ginst9535 (U6090, U3075, U4043);
  nand ginst9536 (U6091, DATAO_REG_2__SCAN_IN, U3422);
  nand ginst9537 (U6092, U3065, U4043);
  nand ginst9538 (U6093, DATAO_REG_3__SCAN_IN, U3422);
  nand ginst9539 (U6094, U3061, U4043);
  nand ginst9540 (U6095, DATAO_REG_4__SCAN_IN, U3422);
  nand ginst9541 (U6096, U3057, U4043);
  nand ginst9542 (U6097, DATAO_REG_5__SCAN_IN, U3422);
  nand ginst9543 (U6098, U3064, U4043);
  nand ginst9544 (U6099, DATAO_REG_6__SCAN_IN, U3422);
  nand ginst9545 (U6100, U3068, U4043);
  nand ginst9546 (U6101, DATAO_REG_7__SCAN_IN, U3422);
  nand ginst9547 (U6102, U3067, U4043);
  nand ginst9548 (U6103, DATAO_REG_8__SCAN_IN, U3422);
  nand ginst9549 (U6104, U3081, U4043);
  nand ginst9550 (U6105, DATAO_REG_9__SCAN_IN, U3422);
  nand ginst9551 (U6106, U3080, U4043);
  nand ginst9552 (U6107, DATAO_REG_10__SCAN_IN, U3422);
  nand ginst9553 (U6108, U3059, U4043);
  nand ginst9554 (U6109, DATAO_REG_11__SCAN_IN, U3422);
  nand ginst9555 (U6110, U3060, U4043);
  nand ginst9556 (U6111, DATAO_REG_12__SCAN_IN, U3422);
  nand ginst9557 (U6112, U3069, U4043);
  nand ginst9558 (U6113, DATAO_REG_13__SCAN_IN, U3422);
  nand ginst9559 (U6114, U3077, U4043);
  nand ginst9560 (U6115, DATAO_REG_14__SCAN_IN, U3422);
  nand ginst9561 (U6116, U3076, U4043);
  nand ginst9562 (U6117, DATAO_REG_15__SCAN_IN, U3422);
  nand ginst9563 (U6118, U3071, U4043);
  nand ginst9564 (U6119, DATAO_REG_16__SCAN_IN, U3422);
  nand ginst9565 (U6120, U3070, U4043);
  nand ginst9566 (U6121, DATAO_REG_17__SCAN_IN, U3422);
  nand ginst9567 (U6122, U3066, U4043);
  nand ginst9568 (U6123, DATAO_REG_18__SCAN_IN, U3422);
  nand ginst9569 (U6124, U3079, U4043);
  nand ginst9570 (U6125, DATAO_REG_19__SCAN_IN, U3422);
  nand ginst9571 (U6126, U3078, U4043);
  nand ginst9572 (U6127, DATAO_REG_20__SCAN_IN, U3422);
  nand ginst9573 (U6128, U3073, U4043);
  nand ginst9574 (U6129, DATAO_REG_21__SCAN_IN, U3422);
  nand ginst9575 (U6130, U3072, U4043);
  nand ginst9576 (U6131, DATAO_REG_22__SCAN_IN, U3422);
  nand ginst9577 (U6132, U3058, U4043);
  nand ginst9578 (U6133, DATAO_REG_23__SCAN_IN, U3422);
  nand ginst9579 (U6134, U3063, U4043);
  nand ginst9580 (U6135, DATAO_REG_24__SCAN_IN, U3422);
  nand ginst9581 (U6136, U3062, U4043);
  nand ginst9582 (U6137, DATAO_REG_25__SCAN_IN, U3422);
  nand ginst9583 (U6138, U3055, U4043);
  nand ginst9584 (U6139, DATAO_REG_26__SCAN_IN, U3422);
  nand ginst9585 (U6140, U3054, U4043);
  nand ginst9586 (U6141, DATAO_REG_27__SCAN_IN, U3422);
  nand ginst9587 (U6142, U3050, U4043);
  nand ginst9588 (U6143, DATAO_REG_28__SCAN_IN, U3422);
  nand ginst9589 (U6144, U3051, U4043);
  nand ginst9590 (U6145, DATAO_REG_29__SCAN_IN, U3422);
  nand ginst9591 (U6146, U3052, U4043);
  nand ginst9592 (U6147, DATAO_REG_30__SCAN_IN, U3422);
  nand ginst9593 (U6148, U3056, U4043);
  nand ginst9594 (U6149, DATAO_REG_31__SCAN_IN, U3422);
  nand ginst9595 (U6150, U3053, U4043);
  nand ginst9596 (U6151, U3052, U4040);
  nand ginst9597 (U6152, U3414, U4737);
  nand ginst9598 (U6153, U6151, U6152);
  nand ginst9599 (U6154, U3053, U4038);
  nand ginst9600 (U6155, U3416, U4775);
  nand ginst9601 (U6156, U6154, U6155);
  nand ginst9602 (U6157, U3056, U4039);
  nand ginst9603 (U6158, U3415, U4755);
  nand ginst9604 (U6159, U6157, U6158);
  nand ginst9605 (U6160, U3073, U4037);
  nand ginst9606 (U6161, U3396, U4566);
  nand ginst9607 (U6162, U6160, U6161);
  nand ginst9608 (U6163, U4395, U5892);
  nand ginst9609 (U6164, U3060, U3488);
  nand ginst9610 (U6165, U6163, U6164);
  nand ginst9611 (U6166, U4376, U5887);
  nand ginst9612 (U6167, U3059, U3486);
  nand ginst9613 (U6168, U6166, U6167);
  nand ginst9614 (U6169, U4262, U5857);
  nand ginst9615 (U6170, U3057, U3474);
  nand ginst9616 (U6171, U6169, U6170);
  nand ginst9617 (U6172, U4547, U5932);
  nand ginst9618 (U6173, U3078, U3504);
  nand ginst9619 (U6174, U6172, U6173);
  nand ginst9620 (U6175, U3055, U4032);
  nand ginst9621 (U6176, U3406, U4661);
  nand ginst9622 (U6177, U6175, U6176);
  nand ginst9623 (U6178, U3054, U4031);
  nand ginst9624 (U6179, U3408, U4680);
  nand ginst9625 (U6180, U6178, U6179);
  nand ginst9626 (U6181, U3072, U4036);
  nand ginst9627 (U6182, U3398, U4585);
  nand ginst9628 (U6183, U6181, U6182);
  nand ginst9629 (U6184, U3058, U4035);
  nand ginst9630 (U6185, U3400, U4604);
  nand ginst9631 (U6186, U6184, U6185);
  nand ginst9632 (U6187, U3063, U4034);
  nand ginst9633 (U6188, U3402, U4623);
  nand ginst9634 (U6189, U6187, U6188);
  nand ginst9635 (U6190, U3062, U4033);
  nand ginst9636 (U6191, U3404, U4642);
  nand ginst9637 (U6192, U6190, U6191);
  nand ginst9638 (U6193, U3050, U4030);
  nand ginst9639 (U6194, U3410, U4699);
  nand ginst9640 (U6195, U6193, U6194);
  nand ginst9641 (U6196, U3051, U4029);
  nand ginst9642 (U6197, U3412, U4718);
  nand ginst9643 (U6198, U6196, U6197);
  nand ginst9644 (U6199, U4338, U5877);
  nand ginst9645 (U6200, U3081, U3482);
  nand ginst9646 (U6201, U6199, U6200);
  nand ginst9647 (U6202, U4357, U5882);
  nand ginst9648 (U6203, U3080, U3484);
  nand ginst9649 (U6204, U6202, U6203);
  nand ginst9650 (U6205, U4528, U5927);
  nand ginst9651 (U6206, U3079, U3502);
  nand ginst9652 (U6207, U6205, U6206);
  nand ginst9653 (U6208, U4433, U5902);
  nand ginst9654 (U6209, U3077, U3492);
  nand ginst9655 (U6210, U6208, U6209);
  nand ginst9656 (U6211, U4452, U5907);
  nand ginst9657 (U6212, U3076, U3494);
  nand ginst9658 (U6213, U6211, U6212);
  nand ginst9659 (U6214, U4200, U5842);
  nand ginst9660 (U6215, U3075, U3468);
  nand ginst9661 (U6216, U6214, U6215);
  nand ginst9662 (U6217, U4224, U5829);
  nand ginst9663 (U6218, U3074, U3464);
  nand ginst9664 (U6219, U6217, U6218);
  nand ginst9665 (U6220, U4471, U5912);
  nand ginst9666 (U6221, U3071, U3496);
  nand ginst9667 (U6222, U6220, U6221);
  nand ginst9668 (U6223, U4490, U5917);
  nand ginst9669 (U6224, U3070, U3498);
  nand ginst9670 (U6225, U6223, U6224);
  nand ginst9671 (U6226, U4414, U5897);
  nand ginst9672 (U6227, U3069, U3490);
  nand ginst9673 (U6228, U6226, U6227);
  nand ginst9674 (U6229, U4300, U5867);
  nand ginst9675 (U6230, U3068, U3478);
  nand ginst9676 (U6231, U6229, U6230);
  nand ginst9677 (U6232, U4319, U5872);
  nand ginst9678 (U6233, U3067, U3480);
  nand ginst9679 (U6234, U6232, U6233);
  nand ginst9680 (U6235, U4509, U5922);
  nand ginst9681 (U6236, U3066, U3500);
  nand ginst9682 (U6237, U6235, U6236);
  nand ginst9683 (U6238, U4219, U5847);
  nand ginst9684 (U6239, U3065, U3470);
  nand ginst9685 (U6240, U6238, U6239);
  nand ginst9686 (U6241, U4281, U5862);
  nand ginst9687 (U6242, U3064, U3476);
  nand ginst9688 (U6243, U6241, U6242);
  nand ginst9689 (U6244, U4243, U5852);
  nand ginst9690 (U6245, U3061, U3472);
  nand ginst9691 (U6246, U6244, U6245);
  nand ginst9692 (U6247, U3424, U4042);
  nand ginst9693 (U6248, R1375_U26, U3373);
  nand ginst9694 (U6249, U6247, U6248);
  nand ginst9695 (U6250, U5820, U6249);
  nand ginst9696 (U6251, R395_U6, U3460, U4042);
  nand ginst9697 (U6252, U5139, U5817);
  nand ginst9698 (U6253, U3425, U3461, U4055);
  nand ginst9699 (U6254, U4007, U4014);
  nand ginst9700 (U6255, R1347_U13, U4023);
  nand ginst9701 (U6256, U3423, U5748);
  nand ginst9702 (U6257, U3431, U3456);
  nand ginst9703 (U6258, U3453, U5421);
  nand ginst9704 (U6259, REG2_REG_0__SCAN_IN, U3016, U5796);
  nand ginst9705 (U6260, R1352_U6, U3080);
  nand ginst9706 (U6261, U3080, U4009);
  nand ginst9707 (U6262, R1352_U6, U3081);
  nand ginst9708 (U6263, U3081, U4009);
  nand ginst9709 (U6264, R1352_U6, U3067);
  nand ginst9710 (U6265, U3067, U4009);
  nand ginst9711 (U6266, R1352_U6, U3068);
  nand ginst9712 (U6267, U3068, U4009);
  nand ginst9713 (U6268, R1352_U6, U3064);
  nand ginst9714 (U6269, U3064, U4009);
  nand ginst9715 (U6270, R1352_U6, U3057);
  nand ginst9716 (U6271, U3057, U4009);
  nand ginst9717 (U6272, R1309_U8, R1352_U6);
  nand ginst9718 (U6273, U3053, U4009);
  nand ginst9719 (U6274, R1309_U6, R1352_U6);
  nand ginst9720 (U6275, U3056, U4009);
  nand ginst9721 (U6276, R1352_U6, U3061);
  nand ginst9722 (U6277, U3061, U4009);
  nand ginst9723 (U6278, R1352_U6, U3052);
  nand ginst9724 (U6279, U3052, U4009);
  nand ginst9725 (U6280, R1352_U6, U3051);
  nand ginst9726 (U6281, U3051, U4009);
  nand ginst9727 (U6282, R1352_U6, U3050);
  nand ginst9728 (U6283, U3050, U4009);
  nand ginst9729 (U6284, R1352_U6, U3054);
  nand ginst9730 (U6285, U3054, U4009);
  nand ginst9731 (U6286, R1352_U6, U3055);
  nand ginst9732 (U6287, U3055, U4009);
  nand ginst9733 (U6288, R1352_U6, U3062);
  nand ginst9734 (U6289, U3062, U4009);
  nand ginst9735 (U6290, R1352_U6, U3063);
  nand ginst9736 (U6291, U3063, U4009);
  nand ginst9737 (U6292, R1352_U6, U3058);
  nand ginst9738 (U6293, U3058, U4009);
  nand ginst9739 (U6294, R1352_U6, U3072);
  nand ginst9740 (U6295, U3072, U4009);
  nand ginst9741 (U6296, R1352_U6, U3073);
  nand ginst9742 (U6297, U3073, U4009);
  nand ginst9743 (U6298, R1352_U6, U3065);
  nand ginst9744 (U6299, U3065, U4009);
  nand ginst9745 (U6300, R1352_U6, U3078);
  nand ginst9746 (U6301, U3078, U4009);
  nand ginst9747 (U6302, R1352_U6, U3079);
  nand ginst9748 (U6303, U3079, U4009);
  nand ginst9749 (U6304, R1352_U6, U3066);
  nand ginst9750 (U6305, U3066, U4009);
  nand ginst9751 (U6306, R1352_U6, U3070);
  nand ginst9752 (U6307, U3070, U4009);
  nand ginst9753 (U6308, R1352_U6, U3071);
  nand ginst9754 (U6309, U3071, U4009);
  nand ginst9755 (U6310, R1352_U6, U3076);
  nand ginst9756 (U6311, U3076, U4009);
  nand ginst9757 (U6312, R1352_U6, U3077);
  nand ginst9758 (U6313, U3077, U4009);
  nand ginst9759 (U6314, R1352_U6, U3069);
  nand ginst9760 (U6315, U3069, U4009);
  nand ginst9761 (U6316, R1352_U6, U3060);
  nand ginst9762 (U6317, U3060, U4009);
  nand ginst9763 (U6318, R1352_U6, U3059);
  nand ginst9764 (U6319, U3059, U4009);
  nand ginst9765 (U6320, R1352_U6, U3075);
  nand ginst9766 (U6321, U3075, U4009);
  nand ginst9767 (U6322, R1352_U6, U3074);
  nand ginst9768 (U6323, U3074, U4009);

SatHard block1 (flip_signal, SUB_84_U63, SUB_84_U80, SUB_84_U64, SUB_84_U150, IR_REG_5__SCAN_IN, U5750, U5753, SUB_84_U125, SUB_84_U78, IR_REG_17__SCAN_IN, D_REG_6__SCAN_IN, SUB_84_U36, SUB_84_U38, SUB_84_U5, U5756, IR_REG_25__SCAN_IN, IR_REG_3__SCAN_IN, SUB_84_U124, U5749, SUB_84_U59, U3968, IR_REG_24__SCAN_IN, SUB_84_U16, IR_REG_1__SCAN_IN, IR_REG_4__SCAN_IN, IR_REG_7__SCAN_IN, U3967, IR_REG_12__SCAN_IN, SUB_84_U81, IR_REG_10__SCAN_IN, IR_REG_21__SCAN_IN, B_REG_SCAN_IN, keyinput0, keyinput1, keyinput2, keyinput3, keyinput4, keyinput5, keyinput6, keyinput7, keyinput8, keyinput9, keyinput10, keyinput11, keyinput12, keyinput13, keyinput14, keyinput15, keyinput16, keyinput17, keyinput18, keyinput19, keyinput20, keyinput21, keyinput22, keyinput23, keyinput24, keyinput25, keyinput26, keyinput27, keyinput28, keyinput29, keyinput30, keyinput31, keyinput32, keyinput33, keyinput34, keyinput35, keyinput36, keyinput37, keyinput38, keyinput39, keyinput40, keyinput41, keyinput42, keyinput43, keyinput44, keyinput45, keyinput46, keyinput47, keyinput48, keyinput49, keyinput50, keyinput51, keyinput52, keyinput53, keyinput54, keyinput55, keyinput56, keyinput57, keyinput58, keyinput59, keyinput60, keyinput61, keyinput62, keyinput63);

endmodule
/*************** SatHard block ***************/
module SatHard (flip_signal, SUB_84_U63, SUB_84_U80, SUB_84_U64, SUB_84_U150, IR_REG_5__SCAN_IN, U5750, U5753, SUB_84_U125, SUB_84_U78, IR_REG_17__SCAN_IN, D_REG_6__SCAN_IN, SUB_84_U36, SUB_84_U38, SUB_84_U5, U5756, IR_REG_25__SCAN_IN, IR_REG_3__SCAN_IN, SUB_84_U124, U5749, SUB_84_U59, U3968, IR_REG_24__SCAN_IN, SUB_84_U16, IR_REG_1__SCAN_IN, IR_REG_4__SCAN_IN, IR_REG_7__SCAN_IN, U3967, IR_REG_12__SCAN_IN, SUB_84_U81, IR_REG_10__SCAN_IN, IR_REG_21__SCAN_IN, B_REG_SCAN_IN, keyinput0, keyinput1, keyinput2, keyinput3, keyinput4, keyinput5, keyinput6, keyinput7, keyinput8, keyinput9, keyinput10, keyinput11, keyinput12, keyinput13, keyinput14, keyinput15, keyinput16, keyinput17, keyinput18, keyinput19, keyinput20, keyinput21, keyinput22, keyinput23, keyinput24, keyinput25, keyinput26, keyinput27, keyinput28, keyinput29, keyinput30, keyinput31, keyinput32, keyinput33, keyinput34, keyinput35, keyinput36, keyinput37, keyinput38, keyinput39, keyinput40, keyinput41, keyinput42, keyinput43, keyinput44, keyinput45, keyinput46, keyinput47, keyinput48, keyinput49, keyinput50, keyinput51, keyinput52, keyinput53, keyinput54, keyinput55, keyinput56, keyinput57, keyinput58, keyinput59, keyinput60, keyinput61, keyinput62, keyinput63);

  input SUB_84_U63, SUB_84_U80, SUB_84_U64, SUB_84_U150, IR_REG_5__SCAN_IN, U5750, U5753, SUB_84_U125, SUB_84_U78, IR_REG_17__SCAN_IN, D_REG_6__SCAN_IN, SUB_84_U36, SUB_84_U38, SUB_84_U5, U5756, IR_REG_25__SCAN_IN, IR_REG_3__SCAN_IN, SUB_84_U124, U5749, SUB_84_U59, U3968, IR_REG_24__SCAN_IN, SUB_84_U16, IR_REG_1__SCAN_IN, IR_REG_4__SCAN_IN, IR_REG_7__SCAN_IN, U3967, IR_REG_12__SCAN_IN, SUB_84_U81, IR_REG_10__SCAN_IN, IR_REG_21__SCAN_IN, B_REG_SCAN_IN, keyinput0, keyinput1, keyinput2, keyinput3, keyinput4, keyinput5, keyinput6, keyinput7, keyinput8, keyinput9, keyinput10, keyinput11, keyinput12, keyinput13, keyinput14, keyinput15, keyinput16, keyinput17, keyinput18, keyinput19, keyinput20, keyinput21, keyinput22, keyinput23, keyinput24, keyinput25, keyinput26, keyinput27, keyinput28, keyinput29, keyinput30, keyinput31, keyinput32, keyinput33, keyinput34, keyinput35, keyinput36, keyinput37, keyinput38, keyinput39, keyinput40, keyinput41, keyinput42, keyinput43, keyinput44, keyinput45, keyinput46, keyinput47, keyinput48, keyinput49, keyinput50, keyinput51, keyinput52, keyinput53, keyinput54, keyinput55, keyinput56, keyinput57, keyinput58, keyinput59, keyinput60, keyinput61, keyinput62, keyinput63;
  output flip_signal;
  //SatHard key=0011110010011111110011011101100011100110100000110010100100111110
  wire [31:0] sat_res_inputs;
  assign sat_res_inputs[31:0] = {SUB_84_U63, SUB_84_U80, SUB_84_U64, SUB_84_U150, IR_REG_5__SCAN_IN, U5750, U5753, SUB_84_U125, SUB_84_U78, IR_REG_17__SCAN_IN, D_REG_6__SCAN_IN, SUB_84_U36, SUB_84_U38, SUB_84_U5, U5756, IR_REG_25__SCAN_IN, IR_REG_3__SCAN_IN, SUB_84_U124, U5749, SUB_84_U59, U3968, IR_REG_24__SCAN_IN, SUB_84_U16, IR_REG_1__SCAN_IN, IR_REG_4__SCAN_IN, IR_REG_7__SCAN_IN, U3967, IR_REG_12__SCAN_IN, SUB_84_U81, IR_REG_10__SCAN_IN, IR_REG_21__SCAN_IN, B_REG_SCAN_IN};
  wire [63:0] keyinputs, keyvalue;
  assign keyinputs[63:0] = {keyinput0, keyinput1, keyinput2, keyinput3, keyinput4, keyinput5, keyinput6, keyinput7, keyinput8, keyinput9, keyinput10, keyinput11, keyinput12, keyinput13, keyinput14, keyinput15, keyinput16, keyinput17, keyinput18, keyinput19, keyinput20, keyinput21, keyinput22, keyinput23, keyinput24, keyinput25, keyinput26, keyinput27, keyinput28, keyinput29, keyinput30, keyinput31, keyinput32, keyinput33, keyinput34, keyinput35, keyinput36, keyinput37, keyinput38, keyinput39, keyinput40, keyinput41, keyinput42, keyinput43, keyinput44, keyinput45, keyinput46, keyinput47, keyinput48, keyinput49, keyinput50, keyinput51, keyinput52, keyinput53, keyinput54, keyinput55, keyinput56, keyinput57, keyinput58, keyinput59, keyinput60, keyinput61, keyinput62, keyinput63};
  assign keyvalue[63:0] = 64'b0011110010011111110011011101100011100110100000110010100100111110;

  wire g, g_bar;
  assign g = &(keyinputs[31:0] ^ sat_res_inputs ^ keyvalue[31:0]);
  assign g_bar = ~&(keyinputs[63:32] ^ sat_res_inputs ^ keyvalue[63:32]);
  assign flip_signal = g & g_bar;

endmodule
/*************** SatHard block ***************/
