/*************** Top Level ***************/
module b22_C_AntiSAT_128_1_top (P3_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, SI_28_, SI_27_, SI_26_, SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, SI_19_, SI_18_, SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, SI_10_, SI_9_, SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, SI_0_, P3_RD_REG_SCAN_IN, P3_STATE_REG_SCAN_IN, P3_REG3_REG_7__SCAN_IN, P3_REG3_REG_27__SCAN_IN, P3_REG3_REG_14__SCAN_IN, P3_REG3_REG_23__SCAN_IN, P3_REG3_REG_10__SCAN_IN, P3_REG3_REG_3__SCAN_IN, P3_REG3_REG_19__SCAN_IN, P3_REG3_REG_28__SCAN_IN, P3_REG3_REG_8__SCAN_IN, P3_REG3_REG_1__SCAN_IN, P3_REG3_REG_21__SCAN_IN, P3_REG3_REG_12__SCAN_IN, P3_REG3_REG_25__SCAN_IN, P3_REG3_REG_16__SCAN_IN, P3_REG3_REG_5__SCAN_IN, P3_REG3_REG_17__SCAN_IN, P3_REG3_REG_24__SCAN_IN, P3_REG3_REG_4__SCAN_IN, P3_REG3_REG_9__SCAN_IN, P3_REG3_REG_0__SCAN_IN, P3_REG3_REG_20__SCAN_IN, P3_REG3_REG_13__SCAN_IN, P3_REG3_REG_22__SCAN_IN, P3_REG3_REG_11__SCAN_IN, P3_REG3_REG_2__SCAN_IN, P3_REG3_REG_18__SCAN_IN, P3_REG3_REG_6__SCAN_IN, P3_REG3_REG_26__SCAN_IN, P3_REG3_REG_15__SCAN_IN, P3_B_REG_SCAN_IN, P3_DATAO_REG_31__SCAN_IN, P3_DATAO_REG_30__SCAN_IN, P3_DATAO_REG_29__SCAN_IN, P3_DATAO_REG_28__SCAN_IN, P3_DATAO_REG_27__SCAN_IN, P3_DATAO_REG_26__SCAN_IN, P3_DATAO_REG_25__SCAN_IN, P3_DATAO_REG_24__SCAN_IN, P3_DATAO_REG_23__SCAN_IN, P3_DATAO_REG_22__SCAN_IN, P3_DATAO_REG_21__SCAN_IN, P3_DATAO_REG_20__SCAN_IN, P3_DATAO_REG_19__SCAN_IN, P3_DATAO_REG_18__SCAN_IN, P3_DATAO_REG_17__SCAN_IN, P3_DATAO_REG_16__SCAN_IN, P3_DATAO_REG_15__SCAN_IN, P3_DATAO_REG_14__SCAN_IN, P3_DATAO_REG_13__SCAN_IN, P3_DATAO_REG_12__SCAN_IN, P3_DATAO_REG_11__SCAN_IN, P3_DATAO_REG_10__SCAN_IN, P3_DATAO_REG_9__SCAN_IN, P3_DATAO_REG_8__SCAN_IN, P3_DATAO_REG_7__SCAN_IN, P3_DATAO_REG_6__SCAN_IN, P3_DATAO_REG_5__SCAN_IN, P3_DATAO_REG_4__SCAN_IN, P3_DATAO_REG_3__SCAN_IN, P3_DATAO_REG_2__SCAN_IN, P3_DATAO_REG_1__SCAN_IN, P3_DATAO_REG_0__SCAN_IN, P3_ADDR_REG_0__SCAN_IN, P3_ADDR_REG_1__SCAN_IN, P3_ADDR_REG_2__SCAN_IN, P3_ADDR_REG_3__SCAN_IN, P3_ADDR_REG_4__SCAN_IN, P3_ADDR_REG_5__SCAN_IN, P3_ADDR_REG_6__SCAN_IN, P3_ADDR_REG_7__SCAN_IN, P3_ADDR_REG_8__SCAN_IN, P3_ADDR_REG_9__SCAN_IN, P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN, P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN, P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN, P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN, P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN, P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN, P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN, P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN, P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN, P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN, P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN, P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN, P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN, P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN, P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN, P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN, P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN, P1_REG1_REG_3__SCAN_IN, P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN, P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN, P1_REG1_REG_9__SCAN_IN, P1_REG1_REG_10__SCAN_IN, P1_REG1_REG_11__SCAN_IN, P1_REG1_REG_12__SCAN_IN, P1_REG1_REG_13__SCAN_IN, P1_REG1_REG_14__SCAN_IN, P1_REG1_REG_15__SCAN_IN, P1_REG1_REG_16__SCAN_IN, P1_REG1_REG_17__SCAN_IN, P1_REG1_REG_18__SCAN_IN, P1_REG1_REG_19__SCAN_IN, P1_REG1_REG_20__SCAN_IN, P1_REG1_REG_21__SCAN_IN, P1_REG1_REG_22__SCAN_IN, P1_REG1_REG_23__SCAN_IN, P1_REG1_REG_24__SCAN_IN, P1_REG1_REG_25__SCAN_IN, P1_REG1_REG_26__SCAN_IN, P1_REG1_REG_27__SCAN_IN, P1_REG1_REG_28__SCAN_IN, P1_REG1_REG_29__SCAN_IN, P1_REG1_REG_30__SCAN_IN, P1_REG1_REG_31__SCAN_IN, P1_REG2_REG_0__SCAN_IN, P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN, P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN, P1_REG2_REG_6__SCAN_IN, P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN, P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN, P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN, P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN, P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN, P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN, P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN, P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN, P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN, P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN, P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN, P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN, P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN, P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN, P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN, P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN, P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN, P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN, P1_ADDR_REG_6__SCAN_IN, P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN, P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN, P1_ADDR_REG_0__SCAN_IN, P1_DATAO_REG_0__SCAN_IN, P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, P1_REG3_REG_15__SCAN_IN, P1_REG3_REG_26__SCAN_IN, P1_REG3_REG_6__SCAN_IN, P1_REG3_REG_18__SCAN_IN, P1_REG3_REG_2__SCAN_IN, P1_REG3_REG_11__SCAN_IN, P1_REG3_REG_22__SCAN_IN, P1_REG3_REG_13__SCAN_IN, P1_REG3_REG_20__SCAN_IN, P1_REG3_REG_0__SCAN_IN, P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN, P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN, P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN, P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN, P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN, P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN, P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN, P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN, P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN, P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN, P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN, P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN, P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN, P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN, P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN, P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN, P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN, P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN, P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN, P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN, P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN, P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN, P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN, P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN, P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN, P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN, P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN, P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN, P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN, P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN, P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN, P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN, P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN, P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN, P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN, P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN, P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN, P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN, P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN, P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN, P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN, P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN, P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN, P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN, P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN, P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN, P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN, P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN, P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN, P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN, P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN, P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN, P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN, P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN, P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN, P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN, P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN, P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN, P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN, P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN, P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN, P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN, P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN, P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN, P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN, P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN, P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN, P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN, P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN, P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN, P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN, P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN, P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN, P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN, P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN, P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN, P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN, P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN, P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN, P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN, P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN, P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN, P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN, P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN, P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN, P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN, P2_DATAO_REG_5__SCAN_IN, P2_DATAO_REG_6__SCAN_IN, P2_DATAO_REG_7__SCAN_IN, P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_9__SCAN_IN, P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_11__SCAN_IN, P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_13__SCAN_IN, P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_15__SCAN_IN, P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_17__SCAN_IN, P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_19__SCAN_IN, P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_21__SCAN_IN, P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_23__SCAN_IN, P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_25__SCAN_IN, P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_27__SCAN_IN, P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_29__SCAN_IN, P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_31__SCAN_IN, P2_B_REG_SCAN_IN, P2_REG3_REG_15__SCAN_IN, P2_REG3_REG_26__SCAN_IN, P2_REG3_REG_6__SCAN_IN, P2_REG3_REG_18__SCAN_IN, P2_REG3_REG_2__SCAN_IN, P2_REG3_REG_11__SCAN_IN, P2_REG3_REG_22__SCAN_IN, P2_REG3_REG_13__SCAN_IN, P2_REG3_REG_20__SCAN_IN, P2_REG3_REG_0__SCAN_IN, P2_REG3_REG_9__SCAN_IN, P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_24__SCAN_IN, P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_5__SCAN_IN, P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_25__SCAN_IN, P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_21__SCAN_IN, P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_8__SCAN_IN, P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_19__SCAN_IN, P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_10__SCAN_IN, P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_14__SCAN_IN, P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_7__SCAN_IN, P2_STATE_REG_SCAN_IN, P2_RD_REG_SCAN_IN, P2_WR_REG_SCAN_IN, P3_IR_REG_0__SCAN_IN, P3_IR_REG_1__SCAN_IN, P3_IR_REG_2__SCAN_IN, P3_IR_REG_3__SCAN_IN, P3_IR_REG_4__SCAN_IN, P3_IR_REG_5__SCAN_IN, P3_IR_REG_6__SCAN_IN, P3_IR_REG_7__SCAN_IN, P3_IR_REG_8__SCAN_IN, P3_IR_REG_9__SCAN_IN, P3_IR_REG_10__SCAN_IN, P3_IR_REG_11__SCAN_IN, P3_IR_REG_12__SCAN_IN, P3_IR_REG_13__SCAN_IN, P3_IR_REG_14__SCAN_IN, P3_IR_REG_15__SCAN_IN, P3_IR_REG_16__SCAN_IN, P3_IR_REG_17__SCAN_IN, P3_IR_REG_18__SCAN_IN, P3_IR_REG_19__SCAN_IN, P3_IR_REG_20__SCAN_IN, P3_IR_REG_21__SCAN_IN, P3_IR_REG_22__SCAN_IN, P3_IR_REG_23__SCAN_IN, P3_IR_REG_24__SCAN_IN, P3_IR_REG_25__SCAN_IN, P3_IR_REG_26__SCAN_IN, P3_IR_REG_27__SCAN_IN, P3_IR_REG_28__SCAN_IN, P3_IR_REG_29__SCAN_IN, P3_IR_REG_30__SCAN_IN, P3_IR_REG_31__SCAN_IN, P3_D_REG_0__SCAN_IN, P3_D_REG_1__SCAN_IN, P3_D_REG_2__SCAN_IN, P3_D_REG_3__SCAN_IN, P3_D_REG_4__SCAN_IN, P3_D_REG_5__SCAN_IN, P3_D_REG_6__SCAN_IN, P3_D_REG_7__SCAN_IN, P3_D_REG_8__SCAN_IN, P3_D_REG_9__SCAN_IN, P3_D_REG_10__SCAN_IN, P3_D_REG_11__SCAN_IN, P3_D_REG_12__SCAN_IN, P3_D_REG_13__SCAN_IN, P3_D_REG_14__SCAN_IN, P3_D_REG_15__SCAN_IN, P3_D_REG_16__SCAN_IN, P3_D_REG_17__SCAN_IN, P3_D_REG_18__SCAN_IN, P3_D_REG_19__SCAN_IN, P3_D_REG_20__SCAN_IN, P3_D_REG_21__SCAN_IN, P3_D_REG_22__SCAN_IN, P3_D_REG_23__SCAN_IN, P3_D_REG_24__SCAN_IN, P3_D_REG_25__SCAN_IN, P3_D_REG_26__SCAN_IN, P3_D_REG_27__SCAN_IN, P3_D_REG_28__SCAN_IN, P3_D_REG_29__SCAN_IN, P3_D_REG_30__SCAN_IN, P3_D_REG_31__SCAN_IN, P3_REG0_REG_0__SCAN_IN, P3_REG0_REG_1__SCAN_IN, P3_REG0_REG_2__SCAN_IN, P3_REG0_REG_3__SCAN_IN, P3_REG0_REG_4__SCAN_IN, P3_REG0_REG_5__SCAN_IN, P3_REG0_REG_6__SCAN_IN, P3_REG0_REG_7__SCAN_IN, P3_REG0_REG_8__SCAN_IN, P3_REG0_REG_9__SCAN_IN, P3_REG0_REG_10__SCAN_IN, P3_REG0_REG_11__SCAN_IN, P3_REG0_REG_12__SCAN_IN, P3_REG0_REG_13__SCAN_IN, P3_REG0_REG_14__SCAN_IN, P3_REG0_REG_15__SCAN_IN, P3_REG0_REG_16__SCAN_IN, P3_REG0_REG_17__SCAN_IN, P3_REG0_REG_18__SCAN_IN, P3_REG0_REG_19__SCAN_IN, P3_REG0_REG_20__SCAN_IN, P3_REG0_REG_21__SCAN_IN, P3_REG0_REG_22__SCAN_IN, P3_REG0_REG_23__SCAN_IN, P3_REG0_REG_24__SCAN_IN, P3_REG0_REG_25__SCAN_IN, P3_REG0_REG_26__SCAN_IN, P3_REG0_REG_27__SCAN_IN, P3_REG0_REG_28__SCAN_IN, P3_REG0_REG_29__SCAN_IN, P3_REG0_REG_30__SCAN_IN, P3_REG0_REG_31__SCAN_IN, P3_REG1_REG_0__SCAN_IN, P3_REG1_REG_1__SCAN_IN, P3_REG1_REG_2__SCAN_IN, P3_REG1_REG_3__SCAN_IN, P3_REG1_REG_4__SCAN_IN, P3_REG1_REG_5__SCAN_IN, P3_REG1_REG_6__SCAN_IN, P3_REG1_REG_7__SCAN_IN, P3_REG1_REG_8__SCAN_IN, P3_REG1_REG_9__SCAN_IN, P3_REG1_REG_10__SCAN_IN, P3_REG1_REG_11__SCAN_IN, P3_REG1_REG_12__SCAN_IN, P3_REG1_REG_13__SCAN_IN, P3_REG1_REG_14__SCAN_IN, P3_REG1_REG_15__SCAN_IN, P3_REG1_REG_16__SCAN_IN, P3_REG1_REG_17__SCAN_IN, P3_REG1_REG_18__SCAN_IN, P3_REG1_REG_19__SCAN_IN, P3_REG1_REG_20__SCAN_IN, P3_REG1_REG_21__SCAN_IN, P3_REG1_REG_22__SCAN_IN, P3_REG1_REG_23__SCAN_IN, P3_REG1_REG_24__SCAN_IN, P3_REG1_REG_25__SCAN_IN, P3_REG1_REG_26__SCAN_IN, P3_REG1_REG_27__SCAN_IN, P3_REG1_REG_28__SCAN_IN, P3_REG1_REG_29__SCAN_IN, P3_REG1_REG_30__SCAN_IN, P3_REG1_REG_31__SCAN_IN, P3_REG2_REG_0__SCAN_IN, P3_REG2_REG_1__SCAN_IN, P3_REG2_REG_2__SCAN_IN, P3_REG2_REG_3__SCAN_IN, P3_REG2_REG_4__SCAN_IN, P3_REG2_REG_5__SCAN_IN, P3_REG2_REG_6__SCAN_IN, P3_REG2_REG_7__SCAN_IN, P3_REG2_REG_8__SCAN_IN, P3_REG2_REG_9__SCAN_IN, P3_REG2_REG_10__SCAN_IN, P3_REG2_REG_11__SCAN_IN, P3_REG2_REG_12__SCAN_IN, P3_REG2_REG_13__SCAN_IN, P3_REG2_REG_14__SCAN_IN, P3_REG2_REG_15__SCAN_IN, P3_REG2_REG_16__SCAN_IN, P3_REG2_REG_17__SCAN_IN, P3_REG2_REG_18__SCAN_IN, P3_REG2_REG_19__SCAN_IN, P3_REG2_REG_20__SCAN_IN, P3_REG2_REG_21__SCAN_IN, P3_REG2_REG_22__SCAN_IN, P3_REG2_REG_23__SCAN_IN, P3_REG2_REG_24__SCAN_IN, P3_REG2_REG_25__SCAN_IN, P3_REG2_REG_26__SCAN_IN, P3_REG2_REG_27__SCAN_IN, P3_REG2_REG_28__SCAN_IN, P3_REG2_REG_29__SCAN_IN, P3_REG2_REG_30__SCAN_IN, P3_REG2_REG_31__SCAN_IN, P3_ADDR_REG_19__SCAN_IN, P3_ADDR_REG_18__SCAN_IN, P3_ADDR_REG_17__SCAN_IN, P3_ADDR_REG_16__SCAN_IN, P3_ADDR_REG_15__SCAN_IN, P3_ADDR_REG_14__SCAN_IN, P3_ADDR_REG_13__SCAN_IN, P3_ADDR_REG_12__SCAN_IN, P3_ADDR_REG_11__SCAN_IN, P3_ADDR_REG_10__SCAN_IN, keyinput0, keyinput1, keyinput2, keyinput3, keyinput4, keyinput5, keyinput6, keyinput7, keyinput8, keyinput9, keyinput10, keyinput11, keyinput12, keyinput13, keyinput14, keyinput15, keyinput16, keyinput17, keyinput18, keyinput19, keyinput20, keyinput21, keyinput22, keyinput23, keyinput24, keyinput25, keyinput26, keyinput27, keyinput28, keyinput29, keyinput30, keyinput31, keyinput32, keyinput33, keyinput34, keyinput35, keyinput36, keyinput37, keyinput38, keyinput39, keyinput40, keyinput41, keyinput42, keyinput43, keyinput44, keyinput45, keyinput46, keyinput47, keyinput48, keyinput49, keyinput50, keyinput51, keyinput52, keyinput53, keyinput54, keyinput55, keyinput56, keyinput57, keyinput58, keyinput59, keyinput60, keyinput61, keyinput62, keyinput63, keyinput64, keyinput65, keyinput66, keyinput67, keyinput68, keyinput69, keyinput70, keyinput71, keyinput72, keyinput73, keyinput74, keyinput75, keyinput76, keyinput77, keyinput78, keyinput79, keyinput80, keyinput81, keyinput82, keyinput83, keyinput84, keyinput85, keyinput86, keyinput87, keyinput88, keyinput89, keyinput90, keyinput91, keyinput92, keyinput93, keyinput94, keyinput95, keyinput96, keyinput97, keyinput98, keyinput99, keyinput100, keyinput101, keyinput102, keyinput103, keyinput104, keyinput105, keyinput106, keyinput107, keyinput108, keyinput109, keyinput110, keyinput111, keyinput112, keyinput113, keyinput114, keyinput115, keyinput116, keyinput117, keyinput118, keyinput119, keyinput120, keyinput121, keyinput122, keyinput123, keyinput124, keyinput125, keyinput126, keyinput127, P3_U3243, P1_U3572, P1_U3356, SUB_1596_U58, P3_U3471, P2_U3278, P2_U3188, P1_U3250, P2_U3316, P3_U3399, P3_U3170, P2_U3251, P1_U3336, P2_U3324, P3_U3272, P1_U3261, P2_U3525, P1_U3278, P1_U3233, P2_U3257, P3_U3483, P2_U3524, P2_U3466, P1_U3578, P3_U3178, P3_U3155, P3_U3520, P1_U3229, P3_U3242, P1_U3241, P2_U3205, P3_U3184, P3_U3268, P1_U3495, P3_U3247, P3_U3246, P1_U3234, P3_U3519, P2_U3275, P2_U3555, SUB_1596_U67, P3_U3450, P1_U3527, P1_U3523, P2_U3488, P3_U3222, P3_U3492, P3_U3252, P2_U3454, P2_U3279, P3_U3491, P2_U3250, P2_U3548, P1_U3515, P3_U3158, P1_U3232, P2_U3185, P1_U3245, P3_U3165, P2_U3294, P2_U3216, P3_U3175, P3_U3208, P2_U3234, P2_U3551, P3_U3181, P2_U3325, P1_U3520, P3_U3396, P3_U3198, P1_U3223, P1_U3086, P3_U3446, P2_U3416, P3_U3461, P3_U3493, P2_U3520, P2_U3535, P2_U3265, P3_U3267, P1_U3537, P1_U3292, P3_U3429, P3_U3460, P3_U3477, P3_U3522, P2_U3498, P1_U3545, P1_U3586, P1_U3272, P2_U3285, P2_U3206, P2_U3228, P3_U3251, P1_U3573, P3_U3263, P3_U3452, P2_U3207, P2_U3512, P3_U3502, P3_U3509, P3_U3196, P1_U3341, P3_U3377, P1_U3550, P3_U3458, P1_U3517, P1_U3280, P2_U3499, P1_U4016, P2_U3269, P2_U3292, P2_U3255, P3_U3188, P2_U3291, P1_U3275, P1_U3235, P1_U3216, P2_U3502, SUB_1596_U65, P2_U3244, P3_U3497, P3_U3441, P1_U3222, P1_U3290, P2_U3282, P1_U3293, P3_U3214, P1_U3590, P2_U3212, P3_U3463, P1_U3347, P3_U3462, P3_U3224, P1_U3282, P2_U3519, P2_U3254, P2_U3513, P2_U3239, P1_U3536, P1_U3581, P2_U3274, P1_U3519, P3_U3221, P1_U3238, P1_U3269, P1_U3344, P3_U3456, P3_U3248, P1_U3333, P3_U3473, P3_U3229, P1_U3308, P2_U3296, P1_U3571, P3_U3289, P3_U3250, P2_U3493, P2_U3211, P1_U3587, P2_U3195, P1_U3543, P3_U3288, P3_U3273, P2_U3544, P3_U3197, U28, P3_U3211, P3_U3187, P1_U3541, P3_U3518, P2_U3270, P1_U3244, P2_U3442, P3_U3226, P1_U3513, P3_U3205, P2_U3503, P1_U3565, P2_U3494, P1_U3215, P1_U3535, SUB_1596_U57, P3_U3185, P3_U3183, P2_U3276, P3_U3438, SUB_1596_U69, P1_U3324, P3_U3506, P1_U3560, P2_U3256, P1_U3558, P2_U3500, P2_U3530, P3_U3163, P1_U3553, P1_U3568, P2_U3214, P1_U3228, P3_U3494, P1_U3291, P1_U3240, P1_U3483, P3_U3154, P3_U3284, P1_U3313, P2_U3264, P2_U3510, P3_U3517, P3_U3513, P3_U3156, P2_U3268, P2_U3259, P3_U3232, P2_U3284, P1_U3263, P2_U3225, P1_U3507, P3_U3166, P2_U3300, P3_U3466, P3_U3164, P3_U3269, P2_U3295, P3_U3233, P2_U3252, P3_U3390, P2_U3550, P3_U3469, P2_U3263, P2_U3310, P3_U3478, P2_U3433, P1_U3338, P2_U3457, P1_U3343, P2_U3193, P1_U3524, P2_U3475, P2_U3280, P1_U3462, P3_U3482, U29, P3_U3227, P3_U3278, P2_U3290, P3_U3508, P3_U3228, P2_U3478, P2_U3490, P1_U3273, P2_U3196, P3_U3168, P2_U3417, P1_U3304, P3_U3271, P1_U3248, P3_U3253, P2_U3491, P2_U3186, P1_U3345, P1_U3346, P3_U3193, P3_U3210, P1_U3510, P3_U3201, P1_U3352, P1_U3221, P2_U3536, P3_U3153, P1_U3085, P3_U3191, SUB_1596_U62, P1_U3249, P2_U3201, P1_U3265, P1_U3486, P3_U3264, P1_U3277, P2_U3463, P3_U3292, P3_U3514, P3_U3296, P2_U3192, SUB_1596_U63, P2_U3299, P2_U3261, P1_U3257, P3_U3236, P2_U3543, P1_U3332, P2_U3309, P2_U3529, P1_U3252, P3_U3215, P1_U3474, P3_U3286, P2_U3227, P1_U3285, P1_U3327, P1_U3504, P3_U3500, P2_U3307, P3_U3280, P1_U3566, P3_U3151, P3_U3487, P1_U3220, P3_U3172, P3_U3167, P1_U3579, P2_U3304, P1_U3294, P2_U3507, P3_U3270, P3_U3432, P1_U3219, P1_U3302, P2_U3549, P3_U3455, P1_U3582, P3_U3467, P3_U3202, P2_U3537, SUB_1596_U53, P2_U3320, P1_U3279, P3_U3294, P1_U3575, P1_U3259, P2_U3240, P1_U3266, P2_U3306, P3_U3501, P1_U3528, P2_U3517, P1_U3534, P1_U3243, P2_U3522, P1_U3226, P1_U3330, P1_U3339, P1_U3547, P1_U3574, P1_U3588, P2_U3293, P1_U3303, P2_U3248, P3_U3414, P3_U3470, P3_U3160, P2_U3489, P3_U3411, P3_U3503, P3_U3449, P1_U3315, P2_U3213, P1_U3555, P1_U3585, P2_U3552, P1_U3549, P2_U3297, P1_U3532, P3_U3453, P3_U3206, P2_U3220, SUB_1596_U4, SUB_1596_U70, P1_U3556, P2_U3508, P3_U3515, P2_U3087, P1_U3349, P1_U3316, P1_U3548, P1_U3271, P3_U3204, P1_U3296, P1_U3237, P2_U3538, P2_U3511, SUB_1596_U60, P1_U3298, P1_U3246, P1_U3218, P1_U3477, P1_U3312, P2_U3301, P2_U3554, P3_U3402, P1_U3459, P1_U3533, P2_U3288, P2_U3222, P1_U3544, P2_U3247, P1_U3583, P2_U3194, P1_U3538, P2_U3258, P2_U3305, P1_U3253, P1_U3284, P2_U3287, P2_U3472, P3_U3516, P1_U3531, P3_U3451, P1_U3564, P3_U3200, SUB_1596_U54, P2_U3226, P2_U3556, P2_U3315, P1_U3224, P1_U3445, P1_U3492, P2_U3545, P2_U3200, P2_U3523, P3_U3510, P2_U3451, P3_U3230, P3_U3176, P3_U3512, P2_U3224, P3_U3207, P3_U3182, P1_U3322, P3_U3474, P2_U3445, P2_U3303, P3_U3157, P3_U3220, P3_U3521, P2_U3547, P3_U3447, P2_U3230, P3_U3257, P3_U3173, P2_U3199, P2_U3273, P3_U3496, P3_U3277, P3_U3507, P1_U3340, P3_U3475, P1_U3307, P2_U3481, P1_U3561, P2_U3436, P3_U3283, P2_U3516, P1_U3334, P1_U3270, P3_U3260, P2_U3232, P1_U3323, P3_U3179, P1_U3231, P3_U3408, P3_U3190, P2_U3558, P1_U3262, P3_U3180, P1_U3213, P1_U3539, P2_U3191, P3_U3499, P2_U3231, P1_U3318, P1_U3354, P1_U3268, P2_U3531, P3_U3171, P3_U3291, P2_U3235, P1_U3569, P1_U3570, P3_U3405, P3_U3465, P1_U3227, P3_U3295, P3_U3199, P1_U3465, P1_U3281, P2_U3439, P1_U3521, P3_U3897, P1_U3299, P2_U3509, P3_U3218, P2_U3198, P3_U3161, P2_U3546, P1_U3255, P2_U3245, P3_U3464, P3_U3484, P2_U3506, P1_U3526, P3_U3249, P1_U3540, P3_U3213, P3_U3489, P3_U3174, P1_U3260, P2_U3208, P1_U3516, P1_U3217, P1_U3551, P3_U3505, P1_U3576, P3_U3235, P1_U3276, SUB_1596_U5, P3_U3225, P1_U3306, P1_U3314, P2_U3237, P3_U3454, P1_U3321, P2_U3533, P3_U3238, P1_U3310, SUB_1596_U56, P2_U3286, P1_U3287, P1_U3264, P2_U3496, P1_U3319, P2_U3262, P3_U3237, P2_U3312, P2_U3528, P3_U3265, P1_U3542, P1_U3242, P2_U3448, P3_U3258, P3_U3498, P1_U3297, P3_U3186, P2_U3318, P3_U3217, P1_U3355, P3_U3485, P1_U3320, P1_U3446, P1_U3489, P2_U3319, P2_U3527, P2_U3553, P3_U3417, P3_U3239, P1_U3557, P2_U3298, P1_U3480, P2_U3223, P1_U3288, P2_U3233, P3_U3216, SUB_1596_U66, SUB_1596_U61, P3_U3472, P2_U3327, P3_U3212, P3_U3511, P1_U3214, P3_U3468, P1_U3239, P3_U3495, P3_U3256, P1_U3529, P1_U3546, P1_U3337, P1_U3522, P2_U3242, P1_U3335, P2_U3532, P2_U3215, P2_U3302, P2_U3277, P2_U3197, P2_U3281, P2_U3560, SUB_1596_U59, P2_U3203, P3_U3423, P2_U3518, P3_U3259, P2_U3088, P2_U3534, P1_U3258, P2_U3484, P1_U3589, P2_U3526, P1_U3328, P2_U3267, SUB_1596_U55, P3_U3241, P1_U3342, P2_U3314, P1_U3309, P1_U3518, P2_U3947, P3_U3245, P1_U3348, SUB_1596_U64, P2_U3317, P2_U3218, P2_U3539, P2_U3542, P2_U3321, P2_U3557, P2_U3210, P2_U3271, P3_U3209, P1_U3552, P2_U3469, P2_U3504, P3_U3262, P3_U3189, P1_U3286, P2_U3322, P3_U3234, P1_U3353, P3_U3159, P1_U3498, P3_U3162, P1_U3350, P3_U3435, P1_U3554, P2_U3492, P2_U3204, P2_U3238, P3_U3490, P3_U3177, P1_U3254, P2_U3311, P3_U3255, P2_U3241, P3_U3444, P1_U3251, P1_U3305, P2_U3501, P2_U3283, P1_U3289, P2_U3430, P2_U3515, P2_U3521, P3_U3203, P1_U3317, P2_U3289, P2_U3260, P2_U3219, P2_U3562, P1_U3563, P3_U3266, P3_U3448, P2_U3514, P1_U3225, P3_U3457, P3_U3282, P1_U3329, SUB_1596_U68, P3_U3195, P2_U3266, P3_U3393, P3_U3275, P2_U3209, P2_U3505, P3_U3244, P3_U3192, P2_U3313, P3_U3376, P3_U3293, P2_U3202, P3_U3479, P3_U3276, P3_U3486, P3_U3290, P2_U3253, P1_U3256, P2_U3308, P3_U3274, P1_U3530, P3_U3254, P1_U3525, P2_U3187, P3_U3480, P2_U3229, P2_U3190, P1_U3267, P3_U3240, P1_U3230, P3_U3285, P3_U3261, P1_U3300, P1_U3325, P2_U3323, P2_U3487, P1_U3274, P2_U3561, P1_U3283, P1_U3236, P3_U3231, P1_U3562, P3_U3287, P2_U3221, P2_U3217, P1_U3311, P3_U3488, P1_U3326, P3_U3194, P1_U3295, P2_U3495, P3_U3219, P1_U3301, P1_U3468, P1_U3580, P1_U3331, P2_U3272, P1_U3501, P3_U3169, P2_U3246, P3_U3426, P3_U3420, P1_U3584, P3_U3223, P2_U3249, P2_U3236, P1_U3559, P1_U3351, P1_U3567, P3_U3481, P2_U3326, P2_U3541, P2_U3559, P3_U3281, P2_U3243, P3_U3150, P3_U3476, P3_U3279, P2_U3540, P1_U3471, P1_U3577, P3_U3459, P2_U3328, P2_U3486, P2_U3497, P3_U3504, P2_U3189, P2_U3460, P1_U3247, P1_U3591);

  input P3_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, SI_28_, SI_27_, SI_26_, SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, SI_19_, SI_18_, SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, SI_10_, SI_9_, SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, SI_0_, P3_RD_REG_SCAN_IN, P3_STATE_REG_SCAN_IN, P3_REG3_REG_7__SCAN_IN, P3_REG3_REG_27__SCAN_IN, P3_REG3_REG_14__SCAN_IN, P3_REG3_REG_23__SCAN_IN, P3_REG3_REG_10__SCAN_IN, P3_REG3_REG_3__SCAN_IN, P3_REG3_REG_19__SCAN_IN, P3_REG3_REG_28__SCAN_IN, P3_REG3_REG_8__SCAN_IN, P3_REG3_REG_1__SCAN_IN, P3_REG3_REG_21__SCAN_IN, P3_REG3_REG_12__SCAN_IN, P3_REG3_REG_25__SCAN_IN, P3_REG3_REG_16__SCAN_IN, P3_REG3_REG_5__SCAN_IN, P3_REG3_REG_17__SCAN_IN, P3_REG3_REG_24__SCAN_IN, P3_REG3_REG_4__SCAN_IN, P3_REG3_REG_9__SCAN_IN, P3_REG3_REG_0__SCAN_IN, P3_REG3_REG_20__SCAN_IN, P3_REG3_REG_13__SCAN_IN, P3_REG3_REG_22__SCAN_IN, P3_REG3_REG_11__SCAN_IN, P3_REG3_REG_2__SCAN_IN, P3_REG3_REG_18__SCAN_IN, P3_REG3_REG_6__SCAN_IN, P3_REG3_REG_26__SCAN_IN, P3_REG3_REG_15__SCAN_IN, P3_B_REG_SCAN_IN, P3_DATAO_REG_31__SCAN_IN, P3_DATAO_REG_30__SCAN_IN, P3_DATAO_REG_29__SCAN_IN, P3_DATAO_REG_28__SCAN_IN, P3_DATAO_REG_27__SCAN_IN, P3_DATAO_REG_26__SCAN_IN, P3_DATAO_REG_25__SCAN_IN, P3_DATAO_REG_24__SCAN_IN, P3_DATAO_REG_23__SCAN_IN, P3_DATAO_REG_22__SCAN_IN, P3_DATAO_REG_21__SCAN_IN, P3_DATAO_REG_20__SCAN_IN, P3_DATAO_REG_19__SCAN_IN, P3_DATAO_REG_18__SCAN_IN, P3_DATAO_REG_17__SCAN_IN, P3_DATAO_REG_16__SCAN_IN, P3_DATAO_REG_15__SCAN_IN, P3_DATAO_REG_14__SCAN_IN, P3_DATAO_REG_13__SCAN_IN, P3_DATAO_REG_12__SCAN_IN, P3_DATAO_REG_11__SCAN_IN, P3_DATAO_REG_10__SCAN_IN, P3_DATAO_REG_9__SCAN_IN, P3_DATAO_REG_8__SCAN_IN, P3_DATAO_REG_7__SCAN_IN, P3_DATAO_REG_6__SCAN_IN, P3_DATAO_REG_5__SCAN_IN, P3_DATAO_REG_4__SCAN_IN, P3_DATAO_REG_3__SCAN_IN, P3_DATAO_REG_2__SCAN_IN, P3_DATAO_REG_1__SCAN_IN, P3_DATAO_REG_0__SCAN_IN, P3_ADDR_REG_0__SCAN_IN, P3_ADDR_REG_1__SCAN_IN, P3_ADDR_REG_2__SCAN_IN, P3_ADDR_REG_3__SCAN_IN, P3_ADDR_REG_4__SCAN_IN, P3_ADDR_REG_5__SCAN_IN, P3_ADDR_REG_6__SCAN_IN, P3_ADDR_REG_7__SCAN_IN, P3_ADDR_REG_8__SCAN_IN, P3_ADDR_REG_9__SCAN_IN, P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN, P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN, P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN, P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN, P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN, P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN, P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN, P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN, P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN, P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN, P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN, P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN, P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN, P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN, P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN, P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN, P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN, P1_REG1_REG_3__SCAN_IN, P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN, P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN, P1_REG1_REG_9__SCAN_IN, P1_REG1_REG_10__SCAN_IN, P1_REG1_REG_11__SCAN_IN, P1_REG1_REG_12__SCAN_IN, P1_REG1_REG_13__SCAN_IN, P1_REG1_REG_14__SCAN_IN, P1_REG1_REG_15__SCAN_IN, P1_REG1_REG_16__SCAN_IN, P1_REG1_REG_17__SCAN_IN, P1_REG1_REG_18__SCAN_IN, P1_REG1_REG_19__SCAN_IN, P1_REG1_REG_20__SCAN_IN, P1_REG1_REG_21__SCAN_IN, P1_REG1_REG_22__SCAN_IN, P1_REG1_REG_23__SCAN_IN, P1_REG1_REG_24__SCAN_IN, P1_REG1_REG_25__SCAN_IN, P1_REG1_REG_26__SCAN_IN, P1_REG1_REG_27__SCAN_IN, P1_REG1_REG_28__SCAN_IN, P1_REG1_REG_29__SCAN_IN, P1_REG1_REG_30__SCAN_IN, P1_REG1_REG_31__SCAN_IN, P1_REG2_REG_0__SCAN_IN, P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN, P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN, P1_REG2_REG_6__SCAN_IN, P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN, P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN, P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN, P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN, P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN, P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN, P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN, P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN, P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN, P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN, P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN, P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN, P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN, P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN, P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN, P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN, P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN, P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN, P1_ADDR_REG_6__SCAN_IN, P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN, P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN, P1_ADDR_REG_0__SCAN_IN, P1_DATAO_REG_0__SCAN_IN, P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, P1_REG3_REG_15__SCAN_IN, P1_REG3_REG_26__SCAN_IN, P1_REG3_REG_6__SCAN_IN, P1_REG3_REG_18__SCAN_IN, P1_REG3_REG_2__SCAN_IN, P1_REG3_REG_11__SCAN_IN, P1_REG3_REG_22__SCAN_IN, P1_REG3_REG_13__SCAN_IN, P1_REG3_REG_20__SCAN_IN, P1_REG3_REG_0__SCAN_IN, P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN, P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN, P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN, P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN, P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN, P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN, P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN, P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN, P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN, P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN, P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN, P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN, P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN, P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN, P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN, P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN, P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN, P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN, P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN, P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN, P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN, P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN, P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN, P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN, P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN, P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN, P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN, P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN, P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN, P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN, P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN, P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN, P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN, P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN, P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN, P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN, P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN, P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN, P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN, P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN, P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN, P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN, P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN, P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN, P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN, P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN, P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN, P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN, P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN, P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN, P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN, P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN, P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN, P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN, P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN, P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN, P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN, P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN, P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN, P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN, P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN, P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN, P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN, P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN, P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN, P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN, P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN, P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN, P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN, P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN, P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN, P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN, P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN, P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN, P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN, P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN, P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN, P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN, P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN, P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN, P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN, P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN, P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN, P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN, P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN, P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN, P2_DATAO_REG_5__SCAN_IN, P2_DATAO_REG_6__SCAN_IN, P2_DATAO_REG_7__SCAN_IN, P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_9__SCAN_IN, P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_11__SCAN_IN, P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_13__SCAN_IN, P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_15__SCAN_IN, P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_17__SCAN_IN, P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_19__SCAN_IN, P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_21__SCAN_IN, P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_23__SCAN_IN, P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_25__SCAN_IN, P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_27__SCAN_IN, P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_29__SCAN_IN, P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_31__SCAN_IN, P2_B_REG_SCAN_IN, P2_REG3_REG_15__SCAN_IN, P2_REG3_REG_26__SCAN_IN, P2_REG3_REG_6__SCAN_IN, P2_REG3_REG_18__SCAN_IN, P2_REG3_REG_2__SCAN_IN, P2_REG3_REG_11__SCAN_IN, P2_REG3_REG_22__SCAN_IN, P2_REG3_REG_13__SCAN_IN, P2_REG3_REG_20__SCAN_IN, P2_REG3_REG_0__SCAN_IN, P2_REG3_REG_9__SCAN_IN, P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_24__SCAN_IN, P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_5__SCAN_IN, P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_25__SCAN_IN, P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_21__SCAN_IN, P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_8__SCAN_IN, P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_19__SCAN_IN, P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_10__SCAN_IN, P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_14__SCAN_IN, P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_7__SCAN_IN, P2_STATE_REG_SCAN_IN, P2_RD_REG_SCAN_IN, P2_WR_REG_SCAN_IN, P3_IR_REG_0__SCAN_IN, P3_IR_REG_1__SCAN_IN, P3_IR_REG_2__SCAN_IN, P3_IR_REG_3__SCAN_IN, P3_IR_REG_4__SCAN_IN, P3_IR_REG_5__SCAN_IN, P3_IR_REG_6__SCAN_IN, P3_IR_REG_7__SCAN_IN, P3_IR_REG_8__SCAN_IN, P3_IR_REG_9__SCAN_IN, P3_IR_REG_10__SCAN_IN, P3_IR_REG_11__SCAN_IN, P3_IR_REG_12__SCAN_IN, P3_IR_REG_13__SCAN_IN, P3_IR_REG_14__SCAN_IN, P3_IR_REG_15__SCAN_IN, P3_IR_REG_16__SCAN_IN, P3_IR_REG_17__SCAN_IN, P3_IR_REG_18__SCAN_IN, P3_IR_REG_19__SCAN_IN, P3_IR_REG_20__SCAN_IN, P3_IR_REG_21__SCAN_IN, P3_IR_REG_22__SCAN_IN, P3_IR_REG_23__SCAN_IN, P3_IR_REG_24__SCAN_IN, P3_IR_REG_25__SCAN_IN, P3_IR_REG_26__SCAN_IN, P3_IR_REG_27__SCAN_IN, P3_IR_REG_28__SCAN_IN, P3_IR_REG_29__SCAN_IN, P3_IR_REG_30__SCAN_IN, P3_IR_REG_31__SCAN_IN, P3_D_REG_0__SCAN_IN, P3_D_REG_1__SCAN_IN, P3_D_REG_2__SCAN_IN, P3_D_REG_3__SCAN_IN, P3_D_REG_4__SCAN_IN, P3_D_REG_5__SCAN_IN, P3_D_REG_6__SCAN_IN, P3_D_REG_7__SCAN_IN, P3_D_REG_8__SCAN_IN, P3_D_REG_9__SCAN_IN, P3_D_REG_10__SCAN_IN, P3_D_REG_11__SCAN_IN, P3_D_REG_12__SCAN_IN, P3_D_REG_13__SCAN_IN, P3_D_REG_14__SCAN_IN, P3_D_REG_15__SCAN_IN, P3_D_REG_16__SCAN_IN, P3_D_REG_17__SCAN_IN, P3_D_REG_18__SCAN_IN, P3_D_REG_19__SCAN_IN, P3_D_REG_20__SCAN_IN, P3_D_REG_21__SCAN_IN, P3_D_REG_22__SCAN_IN, P3_D_REG_23__SCAN_IN, P3_D_REG_24__SCAN_IN, P3_D_REG_25__SCAN_IN, P3_D_REG_26__SCAN_IN, P3_D_REG_27__SCAN_IN, P3_D_REG_28__SCAN_IN, P3_D_REG_29__SCAN_IN, P3_D_REG_30__SCAN_IN, P3_D_REG_31__SCAN_IN, P3_REG0_REG_0__SCAN_IN, P3_REG0_REG_1__SCAN_IN, P3_REG0_REG_2__SCAN_IN, P3_REG0_REG_3__SCAN_IN, P3_REG0_REG_4__SCAN_IN, P3_REG0_REG_5__SCAN_IN, P3_REG0_REG_6__SCAN_IN, P3_REG0_REG_7__SCAN_IN, P3_REG0_REG_8__SCAN_IN, P3_REG0_REG_9__SCAN_IN, P3_REG0_REG_10__SCAN_IN, P3_REG0_REG_11__SCAN_IN, P3_REG0_REG_12__SCAN_IN, P3_REG0_REG_13__SCAN_IN, P3_REG0_REG_14__SCAN_IN, P3_REG0_REG_15__SCAN_IN, P3_REG0_REG_16__SCAN_IN, P3_REG0_REG_17__SCAN_IN, P3_REG0_REG_18__SCAN_IN, P3_REG0_REG_19__SCAN_IN, P3_REG0_REG_20__SCAN_IN, P3_REG0_REG_21__SCAN_IN, P3_REG0_REG_22__SCAN_IN, P3_REG0_REG_23__SCAN_IN, P3_REG0_REG_24__SCAN_IN, P3_REG0_REG_25__SCAN_IN, P3_REG0_REG_26__SCAN_IN, P3_REG0_REG_27__SCAN_IN, P3_REG0_REG_28__SCAN_IN, P3_REG0_REG_29__SCAN_IN, P3_REG0_REG_30__SCAN_IN, P3_REG0_REG_31__SCAN_IN, P3_REG1_REG_0__SCAN_IN, P3_REG1_REG_1__SCAN_IN, P3_REG1_REG_2__SCAN_IN, P3_REG1_REG_3__SCAN_IN, P3_REG1_REG_4__SCAN_IN, P3_REG1_REG_5__SCAN_IN, P3_REG1_REG_6__SCAN_IN, P3_REG1_REG_7__SCAN_IN, P3_REG1_REG_8__SCAN_IN, P3_REG1_REG_9__SCAN_IN, P3_REG1_REG_10__SCAN_IN, P3_REG1_REG_11__SCAN_IN, P3_REG1_REG_12__SCAN_IN, P3_REG1_REG_13__SCAN_IN, P3_REG1_REG_14__SCAN_IN, P3_REG1_REG_15__SCAN_IN, P3_REG1_REG_16__SCAN_IN, P3_REG1_REG_17__SCAN_IN, P3_REG1_REG_18__SCAN_IN, P3_REG1_REG_19__SCAN_IN, P3_REG1_REG_20__SCAN_IN, P3_REG1_REG_21__SCAN_IN, P3_REG1_REG_22__SCAN_IN, P3_REG1_REG_23__SCAN_IN, P3_REG1_REG_24__SCAN_IN, P3_REG1_REG_25__SCAN_IN, P3_REG1_REG_26__SCAN_IN, P3_REG1_REG_27__SCAN_IN, P3_REG1_REG_28__SCAN_IN, P3_REG1_REG_29__SCAN_IN, P3_REG1_REG_30__SCAN_IN, P3_REG1_REG_31__SCAN_IN, P3_REG2_REG_0__SCAN_IN, P3_REG2_REG_1__SCAN_IN, P3_REG2_REG_2__SCAN_IN, P3_REG2_REG_3__SCAN_IN, P3_REG2_REG_4__SCAN_IN, P3_REG2_REG_5__SCAN_IN, P3_REG2_REG_6__SCAN_IN, P3_REG2_REG_7__SCAN_IN, P3_REG2_REG_8__SCAN_IN, P3_REG2_REG_9__SCAN_IN, P3_REG2_REG_10__SCAN_IN, P3_REG2_REG_11__SCAN_IN, P3_REG2_REG_12__SCAN_IN, P3_REG2_REG_13__SCAN_IN, P3_REG2_REG_14__SCAN_IN, P3_REG2_REG_15__SCAN_IN, P3_REG2_REG_16__SCAN_IN, P3_REG2_REG_17__SCAN_IN, P3_REG2_REG_18__SCAN_IN, P3_REG2_REG_19__SCAN_IN, P3_REG2_REG_20__SCAN_IN, P3_REG2_REG_21__SCAN_IN, P3_REG2_REG_22__SCAN_IN, P3_REG2_REG_23__SCAN_IN, P3_REG2_REG_24__SCAN_IN, P3_REG2_REG_25__SCAN_IN, P3_REG2_REG_26__SCAN_IN, P3_REG2_REG_27__SCAN_IN, P3_REG2_REG_28__SCAN_IN, P3_REG2_REG_29__SCAN_IN, P3_REG2_REG_30__SCAN_IN, P3_REG2_REG_31__SCAN_IN, P3_ADDR_REG_19__SCAN_IN, P3_ADDR_REG_18__SCAN_IN, P3_ADDR_REG_17__SCAN_IN, P3_ADDR_REG_16__SCAN_IN, P3_ADDR_REG_15__SCAN_IN, P3_ADDR_REG_14__SCAN_IN, P3_ADDR_REG_13__SCAN_IN, P3_ADDR_REG_12__SCAN_IN, P3_ADDR_REG_11__SCAN_IN, P3_ADDR_REG_10__SCAN_IN, keyinput0, keyinput1, keyinput2, keyinput3, keyinput4, keyinput5, keyinput6, keyinput7, keyinput8, keyinput9, keyinput10, keyinput11, keyinput12, keyinput13, keyinput14, keyinput15, keyinput16, keyinput17, keyinput18, keyinput19, keyinput20, keyinput21, keyinput22, keyinput23, keyinput24, keyinput25, keyinput26, keyinput27, keyinput28, keyinput29, keyinput30, keyinput31, keyinput32, keyinput33, keyinput34, keyinput35, keyinput36, keyinput37, keyinput38, keyinput39, keyinput40, keyinput41, keyinput42, keyinput43, keyinput44, keyinput45, keyinput46, keyinput47, keyinput48, keyinput49, keyinput50, keyinput51, keyinput52, keyinput53, keyinput54, keyinput55, keyinput56, keyinput57, keyinput58, keyinput59, keyinput60, keyinput61, keyinput62, keyinput63, keyinput64, keyinput65, keyinput66, keyinput67, keyinput68, keyinput69, keyinput70, keyinput71, keyinput72, keyinput73, keyinput74, keyinput75, keyinput76, keyinput77, keyinput78, keyinput79, keyinput80, keyinput81, keyinput82, keyinput83, keyinput84, keyinput85, keyinput86, keyinput87, keyinput88, keyinput89, keyinput90, keyinput91, keyinput92, keyinput93, keyinput94, keyinput95, keyinput96, keyinput97, keyinput98, keyinput99, keyinput100, keyinput101, keyinput102, keyinput103, keyinput104, keyinput105, keyinput106, keyinput107, keyinput108, keyinput109, keyinput110, keyinput111, keyinput112, keyinput113, keyinput114, keyinput115, keyinput116, keyinput117, keyinput118, keyinput119, keyinput120, keyinput121, keyinput122, keyinput123, keyinput124, keyinput125, keyinput126, keyinput127;
  output P3_U3243, P1_U3572, P1_U3356, SUB_1596_U58, P3_U3471, P2_U3278, P2_U3188, P1_U3250, P2_U3316, P3_U3399, P3_U3170, P2_U3251, P1_U3336, P2_U3324, P3_U3272, P1_U3261, P2_U3525, P1_U3278, P1_U3233, P2_U3257, P3_U3483, P2_U3524, P2_U3466, P1_U3578, P3_U3178, P3_U3155, P3_U3520, P1_U3229, P3_U3242, P1_U3241, P2_U3205, P3_U3184, P3_U3268, P1_U3495, P3_U3247, P3_U3246, P1_U3234, P3_U3519, P2_U3275, P2_U3555, SUB_1596_U67, P3_U3450, P1_U3527, P1_U3523, P2_U3488, P3_U3222, P3_U3492, P3_U3252, P2_U3454, P2_U3279, P3_U3491, P2_U3250, P2_U3548, P1_U3515, P3_U3158, P1_U3232, P2_U3185, P1_U3245, P3_U3165, P2_U3294, P2_U3216, P3_U3175, P3_U3208, P2_U3234, P2_U3551, P3_U3181, P2_U3325, P1_U3520, P3_U3396, P3_U3198, P1_U3223, P1_U3086, P3_U3446, P2_U3416, P3_U3461, P3_U3493, P2_U3520, P2_U3535, P2_U3265, P3_U3267, P1_U3537, P1_U3292, P3_U3429, P3_U3460, P3_U3477, P3_U3522, P2_U3498, P1_U3545, P1_U3586, P1_U3272, P2_U3285, P2_U3206, P2_U3228, P3_U3251, P1_U3573, P3_U3263, P3_U3452, P2_U3207, P2_U3512, P3_U3502, P3_U3509, P3_U3196, P1_U3341, P3_U3377, P1_U3550, P3_U3458, P1_U3517, P1_U3280, P2_U3499, P1_U4016, P2_U3269, P2_U3292, P2_U3255, P3_U3188, P2_U3291, P1_U3275, P1_U3235, P1_U3216, P2_U3502, SUB_1596_U65, P2_U3244, P3_U3497, P3_U3441, P1_U3222, P1_U3290, P2_U3282, P1_U3293, P3_U3214, P1_U3590, P2_U3212, P3_U3463, P1_U3347, P3_U3462, P3_U3224, P1_U3282, P2_U3519, P2_U3254, P2_U3513, P2_U3239, P1_U3536, P1_U3581, P2_U3274, P1_U3519, P3_U3221, P1_U3238, P1_U3269, P1_U3344, P3_U3456, P3_U3248, P1_U3333, P3_U3473, P3_U3229, P1_U3308, P2_U3296, P1_U3571, P3_U3289, P3_U3250, P2_U3493, P2_U3211, P1_U3587, P2_U3195, P1_U3543, P3_U3288, P3_U3273, P2_U3544, P3_U3197, U28, P3_U3211, P3_U3187, P1_U3541, P3_U3518, P2_U3270, P1_U3244, P2_U3442, P3_U3226, P1_U3513, P3_U3205, P2_U3503, P1_U3565, P2_U3494, P1_U3215, P1_U3535, SUB_1596_U57, P3_U3185, P3_U3183, P2_U3276, P3_U3438, SUB_1596_U69, P1_U3324, P3_U3506, P1_U3560, P2_U3256, P1_U3558, P2_U3500, P2_U3530, P3_U3163, P1_U3553, P1_U3568, P2_U3214, P1_U3228, P3_U3494, P1_U3291, P1_U3240, P1_U3483, P3_U3154, P3_U3284, P1_U3313, P2_U3264, P2_U3510, P3_U3517, P3_U3513, P3_U3156, P2_U3268, P2_U3259, P3_U3232, P2_U3284, P1_U3263, P2_U3225, P1_U3507, P3_U3166, P2_U3300, P3_U3466, P3_U3164, P3_U3269, P2_U3295, P3_U3233, P2_U3252, P3_U3390, P2_U3550, P3_U3469, P2_U3263, P2_U3310, P3_U3478, P2_U3433, P1_U3338, P2_U3457, P1_U3343, P2_U3193, P1_U3524, P2_U3475, P2_U3280, P1_U3462, P3_U3482, U29, P3_U3227, P3_U3278, P2_U3290, P3_U3508, P3_U3228, P2_U3478, P2_U3490, P1_U3273, P2_U3196, P3_U3168, P2_U3417, P1_U3304, P3_U3271, P1_U3248, P3_U3253, P2_U3491, P2_U3186, P1_U3345, P1_U3346, P3_U3193, P3_U3210, P1_U3510, P3_U3201, P1_U3352, P1_U3221, P2_U3536, P3_U3153, P1_U3085, P3_U3191, SUB_1596_U62, P1_U3249, P2_U3201, P1_U3265, P1_U3486, P3_U3264, P1_U3277, P2_U3463, P3_U3292, P3_U3514, P3_U3296, P2_U3192, SUB_1596_U63, P2_U3299, P2_U3261, P1_U3257, P3_U3236, P2_U3543, P1_U3332, P2_U3309, P2_U3529, P1_U3252, P3_U3215, P1_U3474, P3_U3286, P2_U3227, P1_U3285, P1_U3327, P1_U3504, P3_U3500, P2_U3307, P3_U3280, P1_U3566, P3_U3151, P3_U3487, P1_U3220, P3_U3172, P3_U3167, P1_U3579, P2_U3304, P1_U3294, P2_U3507, P3_U3270, P3_U3432, P1_U3219, P1_U3302, P2_U3549, P3_U3455, P1_U3582, P3_U3467, P3_U3202, P2_U3537, SUB_1596_U53, P2_U3320, P1_U3279, P3_U3294, P1_U3575, P1_U3259, P2_U3240, P1_U3266, P2_U3306, P3_U3501, P1_U3528, P2_U3517, P1_U3534, P1_U3243, P2_U3522, P1_U3226, P1_U3330, P1_U3339, P1_U3547, P1_U3574, P1_U3588, P2_U3293, P1_U3303, P2_U3248, P3_U3414, P3_U3470, P3_U3160, P2_U3489, P3_U3411, P3_U3503, P3_U3449, P1_U3315, P2_U3213, P1_U3555, P1_U3585, P2_U3552, P1_U3549, P2_U3297, P1_U3532, P3_U3453, P3_U3206, P2_U3220, SUB_1596_U4, SUB_1596_U70, P1_U3556, P2_U3508, P3_U3515, P2_U3087, P1_U3349, P1_U3316, P1_U3548, P1_U3271, P3_U3204, P1_U3296, P1_U3237, P2_U3538, P2_U3511, SUB_1596_U60, P1_U3298, P1_U3246, P1_U3218, P1_U3477, P1_U3312, P2_U3301, P2_U3554, P3_U3402, P1_U3459, P1_U3533, P2_U3288, P2_U3222, P1_U3544, P2_U3247, P1_U3583, P2_U3194, P1_U3538, P2_U3258, P2_U3305, P1_U3253, P1_U3284, P2_U3287, P2_U3472, P3_U3516, P1_U3531, P3_U3451, P1_U3564, P3_U3200, SUB_1596_U54, P2_U3226, P2_U3556, P2_U3315, P1_U3224, P1_U3445, P1_U3492, P2_U3545, P2_U3200, P2_U3523, P3_U3510, P2_U3451, P3_U3230, P3_U3176, P3_U3512, P2_U3224, P3_U3207, P3_U3182, P1_U3322, P3_U3474, P2_U3445, P2_U3303, P3_U3157, P3_U3220, P3_U3521, P2_U3547, P3_U3447, P2_U3230, P3_U3257, P3_U3173, P2_U3199, P2_U3273, P3_U3496, P3_U3277, P3_U3507, P1_U3340, P3_U3475, P1_U3307, P2_U3481, P1_U3561, P2_U3436, P3_U3283, P2_U3516, P1_U3334, P1_U3270, P3_U3260, P2_U3232, P1_U3323, P3_U3179, P1_U3231, P3_U3408, P3_U3190, P2_U3558, P1_U3262, P3_U3180, P1_U3213, P1_U3539, P2_U3191, P3_U3499, P2_U3231, P1_U3318, P1_U3354, P1_U3268, P2_U3531, P3_U3171, P3_U3291, P2_U3235, P1_U3569, P1_U3570, P3_U3405, P3_U3465, P1_U3227, P3_U3295, P3_U3199, P1_U3465, P1_U3281, P2_U3439, P1_U3521, P3_U3897, P1_U3299, P2_U3509, P3_U3218, P2_U3198, P3_U3161, P2_U3546, P1_U3255, P2_U3245, P3_U3464, P3_U3484, P2_U3506, P1_U3526, P3_U3249, P1_U3540, P3_U3213, P3_U3489, P3_U3174, P1_U3260, P2_U3208, P1_U3516, P1_U3217, P1_U3551, P3_U3505, P1_U3576, P3_U3235, P1_U3276, SUB_1596_U5, P3_U3225, P1_U3306, P1_U3314, P2_U3237, P3_U3454, P1_U3321, P2_U3533, P3_U3238, P1_U3310, SUB_1596_U56, P2_U3286, P1_U3287, P1_U3264, P2_U3496, P1_U3319, P2_U3262, P3_U3237, P2_U3312, P2_U3528, P3_U3265, P1_U3542, P1_U3242, P2_U3448, P3_U3258, P3_U3498, P1_U3297, P3_U3186, P2_U3318, P3_U3217, P1_U3355, P3_U3485, P1_U3320, P1_U3446, P1_U3489, P2_U3319, P2_U3527, P2_U3553, P3_U3417, P3_U3239, P1_U3557, P2_U3298, P1_U3480, P2_U3223, P1_U3288, P2_U3233, P3_U3216, SUB_1596_U66, SUB_1596_U61, P3_U3472, P2_U3327, P3_U3212, P3_U3511, P1_U3214, P3_U3468, P1_U3239, P3_U3495, P3_U3256, P1_U3529, P1_U3546, P1_U3337, P1_U3522, P2_U3242, P1_U3335, P2_U3532, P2_U3215, P2_U3302, P2_U3277, P2_U3197, P2_U3281, P2_U3560, SUB_1596_U59, P2_U3203, P3_U3423, P2_U3518, P3_U3259, P2_U3088, P2_U3534, P1_U3258, P2_U3484, P1_U3589, P2_U3526, P1_U3328, P2_U3267, SUB_1596_U55, P3_U3241, P1_U3342, P2_U3314, P1_U3309, P1_U3518, P2_U3947, P3_U3245, P1_U3348, SUB_1596_U64, P2_U3317, P2_U3218, P2_U3539, P2_U3542, P2_U3321, P2_U3557, P2_U3210, P2_U3271, P3_U3209, P1_U3552, P2_U3469, P2_U3504, P3_U3262, P3_U3189, P1_U3286, P2_U3322, P3_U3234, P1_U3353, P3_U3159, P1_U3498, P3_U3162, P1_U3350, P3_U3435, P1_U3554, P2_U3492, P2_U3204, P2_U3238, P3_U3490, P3_U3177, P1_U3254, P2_U3311, P3_U3255, P2_U3241, P3_U3444, P1_U3251, P1_U3305, P2_U3501, P2_U3283, P1_U3289, P2_U3430, P2_U3515, P2_U3521, P3_U3203, P1_U3317, P2_U3289, P2_U3260, P2_U3219, P2_U3562, P1_U3563, P3_U3266, P3_U3448, P2_U3514, P1_U3225, P3_U3457, P3_U3282, P1_U3329, SUB_1596_U68, P3_U3195, P2_U3266, P3_U3393, P3_U3275, P2_U3209, P2_U3505, P3_U3244, P3_U3192, P2_U3313, P3_U3376, P3_U3293, P2_U3202, P3_U3479, P3_U3276, P3_U3486, P3_U3290, P2_U3253, P1_U3256, P2_U3308, P3_U3274, P1_U3530, P3_U3254, P1_U3525, P2_U3187, P3_U3480, P2_U3229, P2_U3190, P1_U3267, P3_U3240, P1_U3230, P3_U3285, P3_U3261, P1_U3300, P1_U3325, P2_U3323, P2_U3487, P1_U3274, P2_U3561, P1_U3283, P1_U3236, P3_U3231, P1_U3562, P3_U3287, P2_U3221, P2_U3217, P1_U3311, P3_U3488, P1_U3326, P3_U3194, P1_U3295, P2_U3495, P3_U3219, P1_U3301, P1_U3468, P1_U3580, P1_U3331, P2_U3272, P1_U3501, P3_U3169, P2_U3246, P3_U3426, P3_U3420, P1_U3584, P3_U3223, P2_U3249, P2_U3236, P1_U3559, P1_U3351, P1_U3567, P3_U3481, P2_U3326, P2_U3541, P2_U3559, P3_U3281, P2_U3243, P3_U3150, P3_U3476, P3_U3279, P2_U3540, P1_U3471, P1_U3577, P3_U3459, P2_U3328, P2_U3486, P2_U3497, P3_U3504, P2_U3189, P2_U3460, P1_U3247, P1_U3591;
  wire flip_signal;

  b22_C_AntiSAT_128_1 main (P3_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, SI_28_, SI_27_, SI_26_, SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, SI_19_, SI_18_, SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, SI_10_, SI_9_, SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, SI_0_, P3_RD_REG_SCAN_IN, P3_STATE_REG_SCAN_IN, P3_REG3_REG_7__SCAN_IN, P3_REG3_REG_27__SCAN_IN, P3_REG3_REG_14__SCAN_IN, P3_REG3_REG_23__SCAN_IN, P3_REG3_REG_10__SCAN_IN, P3_REG3_REG_3__SCAN_IN, P3_REG3_REG_19__SCAN_IN, P3_REG3_REG_28__SCAN_IN, P3_REG3_REG_8__SCAN_IN, P3_REG3_REG_1__SCAN_IN, P3_REG3_REG_21__SCAN_IN, P3_REG3_REG_12__SCAN_IN, P3_REG3_REG_25__SCAN_IN, P3_REG3_REG_16__SCAN_IN, P3_REG3_REG_5__SCAN_IN, P3_REG3_REG_17__SCAN_IN, P3_REG3_REG_24__SCAN_IN, P3_REG3_REG_4__SCAN_IN, P3_REG3_REG_9__SCAN_IN, P3_REG3_REG_0__SCAN_IN, P3_REG3_REG_20__SCAN_IN, P3_REG3_REG_13__SCAN_IN, P3_REG3_REG_22__SCAN_IN, P3_REG3_REG_11__SCAN_IN, P3_REG3_REG_2__SCAN_IN, P3_REG3_REG_18__SCAN_IN, P3_REG3_REG_6__SCAN_IN, P3_REG3_REG_26__SCAN_IN, P3_REG3_REG_15__SCAN_IN, P3_B_REG_SCAN_IN, P3_DATAO_REG_31__SCAN_IN, P3_DATAO_REG_30__SCAN_IN, P3_DATAO_REG_29__SCAN_IN, P3_DATAO_REG_28__SCAN_IN, P3_DATAO_REG_27__SCAN_IN, P3_DATAO_REG_26__SCAN_IN, P3_DATAO_REG_25__SCAN_IN, P3_DATAO_REG_24__SCAN_IN, P3_DATAO_REG_23__SCAN_IN, P3_DATAO_REG_22__SCAN_IN, P3_DATAO_REG_21__SCAN_IN, P3_DATAO_REG_20__SCAN_IN, P3_DATAO_REG_19__SCAN_IN, P3_DATAO_REG_18__SCAN_IN, P3_DATAO_REG_17__SCAN_IN, P3_DATAO_REG_16__SCAN_IN, P3_DATAO_REG_15__SCAN_IN, P3_DATAO_REG_14__SCAN_IN, P3_DATAO_REG_13__SCAN_IN, P3_DATAO_REG_12__SCAN_IN, P3_DATAO_REG_11__SCAN_IN, P3_DATAO_REG_10__SCAN_IN, P3_DATAO_REG_9__SCAN_IN, P3_DATAO_REG_8__SCAN_IN, P3_DATAO_REG_7__SCAN_IN, P3_DATAO_REG_6__SCAN_IN, P3_DATAO_REG_5__SCAN_IN, P3_DATAO_REG_4__SCAN_IN, P3_DATAO_REG_3__SCAN_IN, P3_DATAO_REG_2__SCAN_IN, P3_DATAO_REG_1__SCAN_IN, P3_DATAO_REG_0__SCAN_IN, P3_ADDR_REG_0__SCAN_IN, P3_ADDR_REG_1__SCAN_IN, P3_ADDR_REG_2__SCAN_IN, P3_ADDR_REG_3__SCAN_IN, P3_ADDR_REG_4__SCAN_IN, P3_ADDR_REG_5__SCAN_IN, P3_ADDR_REG_6__SCAN_IN, P3_ADDR_REG_7__SCAN_IN, P3_ADDR_REG_8__SCAN_IN, P3_ADDR_REG_9__SCAN_IN, P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN, P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN, P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN, P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN, P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN, P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN, P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN, P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN, P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN, P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN, P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN, P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN, P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN, P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN, P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN, P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN, P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN, P1_REG1_REG_3__SCAN_IN, P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN, P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN, P1_REG1_REG_9__SCAN_IN, P1_REG1_REG_10__SCAN_IN, P1_REG1_REG_11__SCAN_IN, P1_REG1_REG_12__SCAN_IN, P1_REG1_REG_13__SCAN_IN, P1_REG1_REG_14__SCAN_IN, P1_REG1_REG_15__SCAN_IN, P1_REG1_REG_16__SCAN_IN, P1_REG1_REG_17__SCAN_IN, P1_REG1_REG_18__SCAN_IN, P1_REG1_REG_19__SCAN_IN, P1_REG1_REG_20__SCAN_IN, P1_REG1_REG_21__SCAN_IN, P1_REG1_REG_22__SCAN_IN, P1_REG1_REG_23__SCAN_IN, P1_REG1_REG_24__SCAN_IN, P1_REG1_REG_25__SCAN_IN, P1_REG1_REG_26__SCAN_IN, P1_REG1_REG_27__SCAN_IN, P1_REG1_REG_28__SCAN_IN, P1_REG1_REG_29__SCAN_IN, P1_REG1_REG_30__SCAN_IN, P1_REG1_REG_31__SCAN_IN, P1_REG2_REG_0__SCAN_IN, P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN, P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN, P1_REG2_REG_6__SCAN_IN, P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN, P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN, P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN, P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN, P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN, P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN, P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN, P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN, P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN, P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN, P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN, P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN, P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN, P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN, P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN, P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN, P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN, P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN, P1_ADDR_REG_6__SCAN_IN, P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN, P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN, P1_ADDR_REG_0__SCAN_IN, P1_DATAO_REG_0__SCAN_IN, P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, P1_REG3_REG_15__SCAN_IN, P1_REG3_REG_26__SCAN_IN, P1_REG3_REG_6__SCAN_IN, P1_REG3_REG_18__SCAN_IN, P1_REG3_REG_2__SCAN_IN, P1_REG3_REG_11__SCAN_IN, P1_REG3_REG_22__SCAN_IN, P1_REG3_REG_13__SCAN_IN, P1_REG3_REG_20__SCAN_IN, P1_REG3_REG_0__SCAN_IN, P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN, P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN, P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN, P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN, P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN, P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN, P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN, P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN, P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN, P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN, P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN, P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN, P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN, P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN, P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN, P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN, P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN, P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN, P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN, P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN, P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN, P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN, P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN, P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN, P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN, P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN, P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN, P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN, P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN, P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN, P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN, P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN, P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN, P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN, P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN, P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN, P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN, P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN, P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN, P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN, P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN, P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN, P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN, P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN, P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN, P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN, P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN, P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN, P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN, P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN, P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN, P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN, P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN, P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN, P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN, P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN, P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN, P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN, P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN, P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN, P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN, P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN, P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN, P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN, P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN, P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN, P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN, P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN, P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN, P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN, P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN, P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN, P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN, P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN, P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN, P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN, P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN, P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN, P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN, P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN, P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN, P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN, P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN, P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN, P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN, P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN, P2_DATAO_REG_5__SCAN_IN, P2_DATAO_REG_6__SCAN_IN, P2_DATAO_REG_7__SCAN_IN, P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_9__SCAN_IN, P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_11__SCAN_IN, P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_13__SCAN_IN, P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_15__SCAN_IN, P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_17__SCAN_IN, P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_19__SCAN_IN, P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_21__SCAN_IN, P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_23__SCAN_IN, P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_25__SCAN_IN, P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_27__SCAN_IN, P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_29__SCAN_IN, P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_31__SCAN_IN, P2_B_REG_SCAN_IN, P2_REG3_REG_15__SCAN_IN, P2_REG3_REG_26__SCAN_IN, P2_REG3_REG_6__SCAN_IN, P2_REG3_REG_18__SCAN_IN, P2_REG3_REG_2__SCAN_IN, P2_REG3_REG_11__SCAN_IN, P2_REG3_REG_22__SCAN_IN, P2_REG3_REG_13__SCAN_IN, P2_REG3_REG_20__SCAN_IN, P2_REG3_REG_0__SCAN_IN, P2_REG3_REG_9__SCAN_IN, P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_24__SCAN_IN, P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_5__SCAN_IN, P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_25__SCAN_IN, P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_21__SCAN_IN, P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_8__SCAN_IN, P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_19__SCAN_IN, P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_10__SCAN_IN, P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_14__SCAN_IN, P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_7__SCAN_IN, P2_STATE_REG_SCAN_IN, P2_RD_REG_SCAN_IN, P2_WR_REG_SCAN_IN, P3_IR_REG_0__SCAN_IN, P3_IR_REG_1__SCAN_IN, P3_IR_REG_2__SCAN_IN, P3_IR_REG_3__SCAN_IN, P3_IR_REG_4__SCAN_IN, P3_IR_REG_5__SCAN_IN, P3_IR_REG_6__SCAN_IN, P3_IR_REG_7__SCAN_IN, P3_IR_REG_8__SCAN_IN, P3_IR_REG_9__SCAN_IN, P3_IR_REG_10__SCAN_IN, P3_IR_REG_11__SCAN_IN, P3_IR_REG_12__SCAN_IN, P3_IR_REG_13__SCAN_IN, P3_IR_REG_14__SCAN_IN, P3_IR_REG_15__SCAN_IN, P3_IR_REG_16__SCAN_IN, P3_IR_REG_17__SCAN_IN, P3_IR_REG_18__SCAN_IN, P3_IR_REG_19__SCAN_IN, P3_IR_REG_20__SCAN_IN, P3_IR_REG_21__SCAN_IN, P3_IR_REG_22__SCAN_IN, P3_IR_REG_23__SCAN_IN, P3_IR_REG_24__SCAN_IN, P3_IR_REG_25__SCAN_IN, P3_IR_REG_26__SCAN_IN, P3_IR_REG_27__SCAN_IN, P3_IR_REG_28__SCAN_IN, P3_IR_REG_29__SCAN_IN, P3_IR_REG_30__SCAN_IN, P3_IR_REG_31__SCAN_IN, P3_D_REG_0__SCAN_IN, P3_D_REG_1__SCAN_IN, P3_D_REG_2__SCAN_IN, P3_D_REG_3__SCAN_IN, P3_D_REG_4__SCAN_IN, P3_D_REG_5__SCAN_IN, P3_D_REG_6__SCAN_IN, P3_D_REG_7__SCAN_IN, P3_D_REG_8__SCAN_IN, P3_D_REG_9__SCAN_IN, P3_D_REG_10__SCAN_IN, P3_D_REG_11__SCAN_IN, P3_D_REG_12__SCAN_IN, P3_D_REG_13__SCAN_IN, P3_D_REG_14__SCAN_IN, P3_D_REG_15__SCAN_IN, P3_D_REG_16__SCAN_IN, P3_D_REG_17__SCAN_IN, P3_D_REG_18__SCAN_IN, P3_D_REG_19__SCAN_IN, P3_D_REG_20__SCAN_IN, P3_D_REG_21__SCAN_IN, P3_D_REG_22__SCAN_IN, P3_D_REG_23__SCAN_IN, P3_D_REG_24__SCAN_IN, P3_D_REG_25__SCAN_IN, P3_D_REG_26__SCAN_IN, P3_D_REG_27__SCAN_IN, P3_D_REG_28__SCAN_IN, P3_D_REG_29__SCAN_IN, P3_D_REG_30__SCAN_IN, P3_D_REG_31__SCAN_IN, P3_REG0_REG_0__SCAN_IN, P3_REG0_REG_1__SCAN_IN, P3_REG0_REG_2__SCAN_IN, P3_REG0_REG_3__SCAN_IN, P3_REG0_REG_4__SCAN_IN, P3_REG0_REG_5__SCAN_IN, P3_REG0_REG_6__SCAN_IN, P3_REG0_REG_7__SCAN_IN, P3_REG0_REG_8__SCAN_IN, P3_REG0_REG_9__SCAN_IN, P3_REG0_REG_10__SCAN_IN, P3_REG0_REG_11__SCAN_IN, P3_REG0_REG_12__SCAN_IN, P3_REG0_REG_13__SCAN_IN, P3_REG0_REG_14__SCAN_IN, P3_REG0_REG_15__SCAN_IN, P3_REG0_REG_16__SCAN_IN, P3_REG0_REG_17__SCAN_IN, P3_REG0_REG_18__SCAN_IN, P3_REG0_REG_19__SCAN_IN, P3_REG0_REG_20__SCAN_IN, P3_REG0_REG_21__SCAN_IN, P3_REG0_REG_22__SCAN_IN, P3_REG0_REG_23__SCAN_IN, P3_REG0_REG_24__SCAN_IN, P3_REG0_REG_25__SCAN_IN, P3_REG0_REG_26__SCAN_IN, P3_REG0_REG_27__SCAN_IN, P3_REG0_REG_28__SCAN_IN, P3_REG0_REG_29__SCAN_IN, P3_REG0_REG_30__SCAN_IN, P3_REG0_REG_31__SCAN_IN, P3_REG1_REG_0__SCAN_IN, P3_REG1_REG_1__SCAN_IN, P3_REG1_REG_2__SCAN_IN, P3_REG1_REG_3__SCAN_IN, P3_REG1_REG_4__SCAN_IN, P3_REG1_REG_5__SCAN_IN, P3_REG1_REG_6__SCAN_IN, P3_REG1_REG_7__SCAN_IN, P3_REG1_REG_8__SCAN_IN, P3_REG1_REG_9__SCAN_IN, P3_REG1_REG_10__SCAN_IN, P3_REG1_REG_11__SCAN_IN, P3_REG1_REG_12__SCAN_IN, P3_REG1_REG_13__SCAN_IN, P3_REG1_REG_14__SCAN_IN, P3_REG1_REG_15__SCAN_IN, P3_REG1_REG_16__SCAN_IN, P3_REG1_REG_17__SCAN_IN, P3_REG1_REG_18__SCAN_IN, P3_REG1_REG_19__SCAN_IN, P3_REG1_REG_20__SCAN_IN, P3_REG1_REG_21__SCAN_IN, P3_REG1_REG_22__SCAN_IN, P3_REG1_REG_23__SCAN_IN, P3_REG1_REG_24__SCAN_IN, P3_REG1_REG_25__SCAN_IN, P3_REG1_REG_26__SCAN_IN, P3_REG1_REG_27__SCAN_IN, P3_REG1_REG_28__SCAN_IN, P3_REG1_REG_29__SCAN_IN, P3_REG1_REG_30__SCAN_IN, P3_REG1_REG_31__SCAN_IN, P3_REG2_REG_0__SCAN_IN, P3_REG2_REG_1__SCAN_IN, P3_REG2_REG_2__SCAN_IN, P3_REG2_REG_3__SCAN_IN, P3_REG2_REG_4__SCAN_IN, P3_REG2_REG_5__SCAN_IN, P3_REG2_REG_6__SCAN_IN, P3_REG2_REG_7__SCAN_IN, P3_REG2_REG_8__SCAN_IN, P3_REG2_REG_9__SCAN_IN, P3_REG2_REG_10__SCAN_IN, P3_REG2_REG_11__SCAN_IN, P3_REG2_REG_12__SCAN_IN, P3_REG2_REG_13__SCAN_IN, P3_REG2_REG_14__SCAN_IN, P3_REG2_REG_15__SCAN_IN, P3_REG2_REG_16__SCAN_IN, P3_REG2_REG_17__SCAN_IN, P3_REG2_REG_18__SCAN_IN, P3_REG2_REG_19__SCAN_IN, P3_REG2_REG_20__SCAN_IN, P3_REG2_REG_21__SCAN_IN, P3_REG2_REG_22__SCAN_IN, P3_REG2_REG_23__SCAN_IN, P3_REG2_REG_24__SCAN_IN, P3_REG2_REG_25__SCAN_IN, P3_REG2_REG_26__SCAN_IN, P3_REG2_REG_27__SCAN_IN, P3_REG2_REG_28__SCAN_IN, P3_REG2_REG_29__SCAN_IN, P3_REG2_REG_30__SCAN_IN, P3_REG2_REG_31__SCAN_IN, P3_ADDR_REG_19__SCAN_IN, P3_ADDR_REG_18__SCAN_IN, P3_ADDR_REG_17__SCAN_IN, P3_ADDR_REG_16__SCAN_IN, P3_ADDR_REG_15__SCAN_IN, P3_ADDR_REG_14__SCAN_IN, P3_ADDR_REG_13__SCAN_IN, P3_ADDR_REG_12__SCAN_IN, P3_ADDR_REG_11__SCAN_IN, P3_ADDR_REG_10__SCAN_IN, flip_signal, SUB_1596_U4, SUB_1596_U62, SUB_1596_U63, SUB_1596_U64, SUB_1596_U65, SUB_1596_U66, SUB_1596_U67, SUB_1596_U68, SUB_1596_U69, SUB_1596_U70, SUB_1596_U54, SUB_1596_U55, SUB_1596_U56, SUB_1596_U57, SUB_1596_U58, SUB_1596_U59, SUB_1596_U60, SUB_1596_U61, SUB_1596_U5, SUB_1596_U53, U29, U28, P1_U3355, P1_U3354, P1_U3353, P1_U3352, P1_U3351, P1_U3350, P1_U3349, P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, P1_U3343, P1_U3342, P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, P1_U3336, P1_U3335, P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, P1_U3329, P1_U3328, P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3445, P1_U3446, P1_U3323, P1_U3322, P1_U3321, P1_U3320, P1_U3319, P1_U3318, P1_U3317, P1_U3316, P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, P1_U3310, P1_U3309, P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, P1_U3303, P1_U3302, P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, P1_U3296, P1_U3295, P1_U3294, P1_U3459, P1_U3462, P1_U3465, P1_U3468, P1_U3471, P1_U3474, P1_U3477, P1_U3480, P1_U3483, P1_U3486, P1_U3489, P1_U3492, P1_U3495, P1_U3498, P1_U3501, P1_U3504, P1_U3507, P1_U3510, P1_U3513, P1_U3515, P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521, P1_U3522, P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528, P1_U3529, P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535, P1_U3536, P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542, P1_U3543, P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549, P1_U3550, P1_U3551, P1_U3552, P1_U3553, P1_U3554, P1_U3555, P1_U3556, P1_U3557, P1_U3558, P1_U3559, P1_U3293, P1_U3292, P1_U3291, P1_U3290, P1_U3289, P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, P1_U3283, P1_U3282, P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, P1_U3276, P1_U3275, P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, P1_U3269, P1_U3268, P1_U3267, P1_U3266, P1_U3265, P1_U3356, P1_U3264, P1_U3263, P1_U3262, P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, P1_U3256, P1_U3255, P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, P1_U3249, P1_U3248, P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, P1_U3560, P1_U3561, P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567, P1_U3568, P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574, P1_U3575, P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581, P1_U3582, P1_U3583, P1_U3584, P1_U3585, P1_U3586, P1_U3587, P1_U3588, P1_U3589, P1_U3590, P1_U3591, P1_U3242, P1_U3241, P1_U3240, P1_U3239, P1_U3238, P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, P1_U3232, P1_U3231, P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, P1_U3225, P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218, P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3086, P1_U3085, P1_U4016, P2_U3327, P2_U3326, P2_U3325, P2_U3324, P2_U3323, P2_U3322, P2_U3321, P2_U3320, P2_U3319, P2_U3318, P2_U3317, P2_U3316, P2_U3315, P2_U3314, P2_U3313, P2_U3312, P2_U3311, P2_U3310, P2_U3309, P2_U3308, P2_U3307, P2_U3306, P2_U3305, P2_U3304, P2_U3303, P2_U3302, P2_U3301, P2_U3300, P2_U3299, P2_U3298, P2_U3297, P2_U3296, P2_U3416, P2_U3417, P2_U3295, P2_U3294, P2_U3293, P2_U3292, P2_U3291, P2_U3290, P2_U3289, P2_U3288, P2_U3287, P2_U3286, P2_U3285, P2_U3284, P2_U3283, P2_U3282, P2_U3281, P2_U3280, P2_U3279, P2_U3278, P2_U3277, P2_U3276, P2_U3275, P2_U3274, P2_U3273, P2_U3272, P2_U3271, P2_U3270, P2_U3269, P2_U3268, P2_U3267, P2_U3266, P2_U3430, P2_U3433, P2_U3436, P2_U3439, P2_U3442, P2_U3445, P2_U3448, P2_U3451, P2_U3454, P2_U3457, P2_U3460, P2_U3463, P2_U3466, P2_U3469, P2_U3472, P2_U3475, P2_U3478, P2_U3481, P2_U3484, P2_U3486, P2_U3487, P2_U3488, P2_U3489, P2_U3490, P2_U3491, P2_U3492, P2_U3493, P2_U3494, P2_U3495, P2_U3496, P2_U3497, P2_U3498, P2_U3499, P2_U3500, P2_U3501, P2_U3502, P2_U3503, P2_U3504, P2_U3505, P2_U3506, P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511, P2_U3512, P2_U3513, P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518, P2_U3519, P2_U3520, P2_U3521, P2_U3522, P2_U3523, P2_U3524, P2_U3525, P2_U3526, P2_U3527, P2_U3528, P2_U3529, P2_U3530, P2_U3265, P2_U3264, P2_U3263, P2_U3262, P2_U3261, P2_U3260, P2_U3259, P2_U3258, P2_U3257, P2_U3256, P2_U3255, P2_U3254, P2_U3253, P2_U3252, P2_U3251, P2_U3250, P2_U3249, P2_U3248, P2_U3247, P2_U3246, P2_U3245, P2_U3244, P2_U3243, P2_U3242, P2_U3241, P2_U3240, P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234, P2_U3233, P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227, P2_U3226, P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220, P2_U3219, P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3214, P2_U3531, P2_U3532, P2_U3533, P2_U3534, P2_U3535, P2_U3536, P2_U3537, P2_U3538, P2_U3539, P2_U3540, P2_U3541, P2_U3542, P2_U3543, P2_U3544, P2_U3545, P2_U3546, P2_U3547, P2_U3548, P2_U3549, P2_U3550, P2_U3551, P2_U3552, P2_U3553, P2_U3554, P2_U3555, P2_U3556, P2_U3557, P2_U3558, P2_U3559, P2_U3560, P2_U3561, P2_U3562, P2_U3328, P2_U3213, P2_U3212, P2_U3211, P2_U3210, P2_U3209, P2_U3208, P2_U3207, P2_U3206, P2_U3205, P2_U3204, P2_U3203, P2_U3202, P2_U3201, P2_U3200, P2_U3199, P2_U3198, P2_U3197, P2_U3196, P2_U3195, P2_U3194, P2_U3193, P2_U3192, P2_U3191, P2_U3190, P2_U3189, P2_U3188, P2_U3187, P2_U3186, P2_U3185, P2_U3088, P2_U3087, P2_U3947, P3_U3295, P3_U3294, P3_U3293, P3_U3292, P3_U3291, P3_U3290, P3_U3289, P3_U3288, P3_U3287, P3_U3286, P3_U3285, P3_U3284, P3_U3283, P3_U3282, P3_U3281, P3_U3280, P3_U3279, P3_U3278, P3_U3277, P3_U3276, P3_U3275, P3_U3274, P3_U3273, P3_U3272, P3_U3271, P3_U3270, P3_U3269, P3_U3268, P3_U3267, P3_U3266, P3_U3265, P3_U3264, P3_U3376, P3_U3377, P3_U3263, P3_U3262, P3_U3261, P3_U3260, P3_U3259, P3_U3258, P3_U3257, P3_U3256, P3_U3255, P3_U3254, P3_U3253, P3_U3252, P3_U3251, P3_U3250, P3_U3249, P3_U3248, P3_U3247, P3_U3246, P3_U3245, P3_U3244, P3_U3243, P3_U3242, P3_U3241, P3_U3240, P3_U3239, P3_U3238, P3_U3237, P3_U3236, P3_U3235, P3_U3234, P3_U3390, P3_U3393, P3_U3396, P3_U3399, P3_U3402, P3_U3405, P3_U3408, P3_U3411, P3_U3414, P3_U3417, P3_U3420, P3_U3423, P3_U3426, P3_U3429, P3_U3432, P3_U3435, P3_U3438, P3_U3441, P3_U3444, P3_U3446, P3_U3447, P3_U3448, P3_U3449, P3_U3450, P3_U3451, P3_U3452, P3_U3453, P3_U3454, P3_U3455, P3_U3456, P3_U3457, P3_U3458, P3_U3459, P3_U3460, P3_U3461, P3_U3462, P3_U3463, P3_U3464, P3_U3465, P3_U3466, P3_U3467, P3_U3468, P3_U3469, P3_U3470, P3_U3471, P3_U3472, P3_U3473, P3_U3474, P3_U3475, P3_U3476, P3_U3477, P3_U3478, P3_U3479, P3_U3480, P3_U3481, P3_U3482, P3_U3483, P3_U3484, P3_U3485, P3_U3486, P3_U3487, P3_U3488, P3_U3489, P3_U3490, P3_U3233, P3_U3232, P3_U3231, P3_U3230, P3_U3229, P3_U3228, P3_U3227, P3_U3226, P3_U3225, P3_U3224, P3_U3223, P3_U3222, P3_U3221, P3_U3220, P3_U3219, P3_U3218, P3_U3217, P3_U3216, P3_U3215, P3_U3214, P3_U3213, P3_U3212, P3_U3211, P3_U3210, P3_U3209, P3_U3208, P3_U3207, P3_U3206, P3_U3205, P3_U3204, P3_U3203, P3_U3202, P3_U3201, P3_U3200, P3_U3199, P3_U3198, P3_U3197, P3_U3196, P3_U3195, P3_U3194, P3_U3193, P3_U3192, P3_U3191, P3_U3190, P3_U3189, P3_U3188, P3_U3187, P3_U3186, P3_U3185, P3_U3184, P3_U3183, P3_U3182, P3_U3491, P3_U3492, P3_U3493, P3_U3494, P3_U3495, P3_U3496, P3_U3497, P3_U3498, P3_U3499, P3_U3500, P3_U3501, P3_U3502, P3_U3503, P3_U3504, P3_U3505, P3_U3506, P3_U3507, P3_U3508, P3_U3509, P3_U3510, P3_U3511, P3_U3512, P3_U3513, P3_U3514, P3_U3515, P3_U3516, P3_U3517, P3_U3518, P3_U3519, P3_U3520, P3_U3521, P3_U3522, P3_U3296, P3_U3181, P3_U3180, P3_U3179, P3_U3178, P3_U3177, P3_U3176, P3_U3175, P3_U3174, P3_U3173, P3_U3172, P3_U3171, P3_U3170, P3_U3169, P3_U3168, P3_U3167, P3_U3166, P3_U3165, P3_U3164, P3_U3163, P3_U3162, P3_U3161, P3_U3160, P3_U3159, P3_U3158, P3_U3157, P3_U3156, P3_U3155, P3_U3154, P3_U3153, P3_U3151, P3_U3150, P3_U3897);
  SatHard flip1 (P2_REG2_REG_9__SCAN_IN, P1_DATAO_REG_0__SCAN_IN, P2_REG2_REG_17__SCAN_IN, P2_D_REG_0__SCAN_IN, P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_18__SCAN_IN, SI_2_, P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_3__SCAN_IN, P2_DATAO_REG_19__SCAN_IN, P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_12__SCAN_IN, P2_DATAO_REG_5__SCAN_IN, P2_DATAO_REG_13__SCAN_IN, P1_RD_REG_SCAN_IN, P1_DATAO_REG_21__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_REG3_REG_22__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_REG3_REG_8__SCAN_IN, P2_IR_REG_7__SCAN_IN, SI_9_, P2_D_REG_11__SCAN_IN, SI_8_, SI_3_, P2_IR_REG_8__SCAN_IN, P1_DATAO_REG_6__SCAN_IN, P2_REG0_REG_2__SCAN_IN, P2_IR_REG_10__SCAN_IN, P1_DATAO_REG_13__SCAN_IN, P2_REG3_REG_20__SCAN_IN, P2_D_REG_2__SCAN_IN, P2_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_5__SCAN_IN, P2_REG0_REG_16__SCAN_IN, P2_DATAO_REG_14__SCAN_IN, P2_REG0_REG_1__SCAN_IN, SI_12_, P2_REG0_REG_0__SCAN_IN, P2_B_REG_SCAN_IN, P2_IR_REG_2__SCAN_IN, P1_DATAO_REG_17__SCAN_IN, P2_REG2_REG_13__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_REG3_REG_16__SCAN_IN, P2_DATAO_REG_1__SCAN_IN, SI_6_, P1_DATAO_REG_10__SCAN_IN, P2_IR_REG_25__SCAN_IN, P2_REG1_REG_9__SCAN_IN, P1_DATAO_REG_7__SCAN_IN, P2_REG0_REG_11__SCAN_IN, P2_D_REG_24__SCAN_IN, P2_IR_REG_5__SCAN_IN, P2_REG2_REG_21__SCAN_IN, P2_REG3_REG_17__SCAN_IN, P2_REG1_REG_8__SCAN_IN, P2_IR_REG_28__SCAN_IN, P2_REG2_REG_16__SCAN_IN, P2_DATAO_REG_11__SCAN_IN, P2_REG3_REG_14__SCAN_IN, P2_REG1_REG_17__SCAN_IN, P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_15__SCAN_IN, keyinput0, keyinput1, keyinput2, keyinput3, keyinput4, keyinput5, keyinput6, keyinput7, keyinput8, keyinput9, keyinput10, keyinput11, keyinput12, keyinput13, keyinput14, keyinput15, keyinput16, keyinput17, keyinput18, keyinput19, keyinput20, keyinput21, keyinput22, keyinput23, keyinput24, keyinput25, keyinput26, keyinput27, keyinput28, keyinput29, keyinput30, keyinput31, keyinput32, keyinput33, keyinput34, keyinput35, keyinput36, keyinput37, keyinput38, keyinput39, keyinput40, keyinput41, keyinput42, keyinput43, keyinput44, keyinput45, keyinput46, keyinput47, keyinput48, keyinput49, keyinput50, keyinput51, keyinput52, keyinput53, keyinput54, keyinput55, keyinput56, keyinput57, keyinput58, keyinput59, keyinput60, keyinput61, keyinput62, keyinput63, keyinput64, keyinput65, keyinput66, keyinput67, keyinput68, keyinput69, keyinput70, keyinput71, keyinput72, keyinput73, keyinput74, keyinput75, keyinput76, keyinput77, keyinput78, keyinput79, keyinput80, keyinput81, keyinput82, keyinput83, keyinput84, keyinput85, keyinput86, keyinput87, keyinput88, keyinput89, keyinput90, keyinput91, keyinput92, keyinput93, keyinput94, keyinput95, keyinput96, keyinput97, keyinput98, keyinput99, keyinput100, keyinput101, keyinput102, keyinput103, keyinput104, keyinput105, keyinput106, keyinput107, keyinput108, keyinput109, keyinput110, keyinput111, keyinput112, keyinput113, keyinput114, keyinput115, keyinput116, keyinput117, keyinput118, keyinput119, keyinput120, keyinput121, keyinput122, keyinput123, keyinput124, keyinput125, keyinput126, keyinput127, flip_signal);
endmodule
/*************** Top Level ***************/

// Main module
module b22_C_AntiSAT_128_1(P3_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, SI_28_, SI_27_, SI_26_, SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, SI_19_, SI_18_, SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, SI_10_, SI_9_, SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, SI_0_, P3_RD_REG_SCAN_IN, P3_STATE_REG_SCAN_IN, P3_REG3_REG_7__SCAN_IN, P3_REG3_REG_27__SCAN_IN, P3_REG3_REG_14__SCAN_IN, P3_REG3_REG_23__SCAN_IN, P3_REG3_REG_10__SCAN_IN, P3_REG3_REG_3__SCAN_IN, P3_REG3_REG_19__SCAN_IN, P3_REG3_REG_28__SCAN_IN, P3_REG3_REG_8__SCAN_IN, P3_REG3_REG_1__SCAN_IN, P3_REG3_REG_21__SCAN_IN, P3_REG3_REG_12__SCAN_IN, P3_REG3_REG_25__SCAN_IN, P3_REG3_REG_16__SCAN_IN, P3_REG3_REG_5__SCAN_IN, P3_REG3_REG_17__SCAN_IN, P3_REG3_REG_24__SCAN_IN, P3_REG3_REG_4__SCAN_IN, P3_REG3_REG_9__SCAN_IN, P3_REG3_REG_0__SCAN_IN, P3_REG3_REG_20__SCAN_IN, P3_REG3_REG_13__SCAN_IN, P3_REG3_REG_22__SCAN_IN, P3_REG3_REG_11__SCAN_IN, P3_REG3_REG_2__SCAN_IN, P3_REG3_REG_18__SCAN_IN, P3_REG3_REG_6__SCAN_IN, P3_REG3_REG_26__SCAN_IN, P3_REG3_REG_15__SCAN_IN, P3_B_REG_SCAN_IN, P3_DATAO_REG_31__SCAN_IN, P3_DATAO_REG_30__SCAN_IN, P3_DATAO_REG_29__SCAN_IN, P3_DATAO_REG_28__SCAN_IN, P3_DATAO_REG_27__SCAN_IN, P3_DATAO_REG_26__SCAN_IN, P3_DATAO_REG_25__SCAN_IN, P3_DATAO_REG_24__SCAN_IN, P3_DATAO_REG_23__SCAN_IN, P3_DATAO_REG_22__SCAN_IN, P3_DATAO_REG_21__SCAN_IN, P3_DATAO_REG_20__SCAN_IN, P3_DATAO_REG_19__SCAN_IN, P3_DATAO_REG_18__SCAN_IN, P3_DATAO_REG_17__SCAN_IN, P3_DATAO_REG_16__SCAN_IN, P3_DATAO_REG_15__SCAN_IN, P3_DATAO_REG_14__SCAN_IN, P3_DATAO_REG_13__SCAN_IN, P3_DATAO_REG_12__SCAN_IN, P3_DATAO_REG_11__SCAN_IN, P3_DATAO_REG_10__SCAN_IN, P3_DATAO_REG_9__SCAN_IN, P3_DATAO_REG_8__SCAN_IN, P3_DATAO_REG_7__SCAN_IN, P3_DATAO_REG_6__SCAN_IN, P3_DATAO_REG_5__SCAN_IN, P3_DATAO_REG_4__SCAN_IN, P3_DATAO_REG_3__SCAN_IN, P3_DATAO_REG_2__SCAN_IN, P3_DATAO_REG_1__SCAN_IN, P3_DATAO_REG_0__SCAN_IN, P3_ADDR_REG_0__SCAN_IN, P3_ADDR_REG_1__SCAN_IN, P3_ADDR_REG_2__SCAN_IN, P3_ADDR_REG_3__SCAN_IN, P3_ADDR_REG_4__SCAN_IN, P3_ADDR_REG_5__SCAN_IN, P3_ADDR_REG_6__SCAN_IN, P3_ADDR_REG_7__SCAN_IN, P3_ADDR_REG_8__SCAN_IN, P3_ADDR_REG_9__SCAN_IN, P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN, P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN, P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN, P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN, P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN, P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN, P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN, P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN, P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN, P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN, P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN, P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN, P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN, P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN, P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN, P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN, P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN, P1_REG1_REG_3__SCAN_IN, P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN, P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN, P1_REG1_REG_9__SCAN_IN, P1_REG1_REG_10__SCAN_IN, P1_REG1_REG_11__SCAN_IN, P1_REG1_REG_12__SCAN_IN, P1_REG1_REG_13__SCAN_IN, P1_REG1_REG_14__SCAN_IN, P1_REG1_REG_15__SCAN_IN, P1_REG1_REG_16__SCAN_IN, P1_REG1_REG_17__SCAN_IN, P1_REG1_REG_18__SCAN_IN, P1_REG1_REG_19__SCAN_IN, P1_REG1_REG_20__SCAN_IN, P1_REG1_REG_21__SCAN_IN, P1_REG1_REG_22__SCAN_IN, P1_REG1_REG_23__SCAN_IN, P1_REG1_REG_24__SCAN_IN, P1_REG1_REG_25__SCAN_IN, P1_REG1_REG_26__SCAN_IN, P1_REG1_REG_27__SCAN_IN, P1_REG1_REG_28__SCAN_IN, P1_REG1_REG_29__SCAN_IN, P1_REG1_REG_30__SCAN_IN, P1_REG1_REG_31__SCAN_IN, P1_REG2_REG_0__SCAN_IN, P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN, P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN, P1_REG2_REG_6__SCAN_IN, P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN, P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN, P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN, P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN, P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN, P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN, P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN, P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN, P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN, P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN, P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN, P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN, P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN, P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN, P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN, P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN, P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN, P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN, P1_ADDR_REG_6__SCAN_IN, P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN, P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN, P1_ADDR_REG_0__SCAN_IN, P1_DATAO_REG_0__SCAN_IN, P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, P1_REG3_REG_15__SCAN_IN, P1_REG3_REG_26__SCAN_IN, P1_REG3_REG_6__SCAN_IN, P1_REG3_REG_18__SCAN_IN, P1_REG3_REG_2__SCAN_IN, P1_REG3_REG_11__SCAN_IN, P1_REG3_REG_22__SCAN_IN, P1_REG3_REG_13__SCAN_IN, P1_REG3_REG_20__SCAN_IN, P1_REG3_REG_0__SCAN_IN, P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN, P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN, P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN, P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN, P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN, P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN, P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN, P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN, P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN, P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN, P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN, P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN, P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN, P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN, P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN, P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN, P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN, P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN, P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN, P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN, P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN, P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN, P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN, P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN, P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN, P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN, P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN, P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN, P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN, P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN, P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN, P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN, P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN, P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN, P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN, P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN, P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN, P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN, P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN, P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN, P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN, P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN, P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN, P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN, P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN, P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN, P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN, P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN, P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN, P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN, P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN, P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN, P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN, P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN, P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN, P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN, P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN, P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN, P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN, P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN, P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN, P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN, P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN, P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN, P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN, P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN, P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN, P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN, P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN, P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN, P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN, P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN, P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN, P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN, P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN, P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN, P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN, P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN, P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN, P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN, P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN, P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN, P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN, P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN, P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN, P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN, P2_DATAO_REG_5__SCAN_IN, P2_DATAO_REG_6__SCAN_IN, P2_DATAO_REG_7__SCAN_IN, P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_9__SCAN_IN, P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_11__SCAN_IN, P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_13__SCAN_IN, P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_15__SCAN_IN, P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_17__SCAN_IN, P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_19__SCAN_IN, P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_21__SCAN_IN, P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_23__SCAN_IN, P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_25__SCAN_IN, P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_27__SCAN_IN, P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_29__SCAN_IN, P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_31__SCAN_IN, P2_B_REG_SCAN_IN, P2_REG3_REG_15__SCAN_IN, P2_REG3_REG_26__SCAN_IN, P2_REG3_REG_6__SCAN_IN, P2_REG3_REG_18__SCAN_IN, P2_REG3_REG_2__SCAN_IN, P2_REG3_REG_11__SCAN_IN, P2_REG3_REG_22__SCAN_IN, P2_REG3_REG_13__SCAN_IN, P2_REG3_REG_20__SCAN_IN, P2_REG3_REG_0__SCAN_IN, P2_REG3_REG_9__SCAN_IN, P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_24__SCAN_IN, P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_5__SCAN_IN, P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_25__SCAN_IN, P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_21__SCAN_IN, P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_8__SCAN_IN, P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_19__SCAN_IN, P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_10__SCAN_IN, P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_14__SCAN_IN, P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_7__SCAN_IN, P2_STATE_REG_SCAN_IN, P2_RD_REG_SCAN_IN, P2_WR_REG_SCAN_IN, P3_IR_REG_0__SCAN_IN, P3_IR_REG_1__SCAN_IN, P3_IR_REG_2__SCAN_IN, P3_IR_REG_3__SCAN_IN, P3_IR_REG_4__SCAN_IN, P3_IR_REG_5__SCAN_IN, P3_IR_REG_6__SCAN_IN, P3_IR_REG_7__SCAN_IN, P3_IR_REG_8__SCAN_IN, P3_IR_REG_9__SCAN_IN, P3_IR_REG_10__SCAN_IN, P3_IR_REG_11__SCAN_IN, P3_IR_REG_12__SCAN_IN, P3_IR_REG_13__SCAN_IN, P3_IR_REG_14__SCAN_IN, P3_IR_REG_15__SCAN_IN, P3_IR_REG_16__SCAN_IN, P3_IR_REG_17__SCAN_IN, P3_IR_REG_18__SCAN_IN, P3_IR_REG_19__SCAN_IN, P3_IR_REG_20__SCAN_IN, P3_IR_REG_21__SCAN_IN, P3_IR_REG_22__SCAN_IN, P3_IR_REG_23__SCAN_IN, P3_IR_REG_24__SCAN_IN, P3_IR_REG_25__SCAN_IN, P3_IR_REG_26__SCAN_IN, P3_IR_REG_27__SCAN_IN, P3_IR_REG_28__SCAN_IN, P3_IR_REG_29__SCAN_IN, P3_IR_REG_30__SCAN_IN, P3_IR_REG_31__SCAN_IN, P3_D_REG_0__SCAN_IN, P3_D_REG_1__SCAN_IN, P3_D_REG_2__SCAN_IN, P3_D_REG_3__SCAN_IN, P3_D_REG_4__SCAN_IN, P3_D_REG_5__SCAN_IN, P3_D_REG_6__SCAN_IN, P3_D_REG_7__SCAN_IN, P3_D_REG_8__SCAN_IN, P3_D_REG_9__SCAN_IN, P3_D_REG_10__SCAN_IN, P3_D_REG_11__SCAN_IN, P3_D_REG_12__SCAN_IN, P3_D_REG_13__SCAN_IN, P3_D_REG_14__SCAN_IN, P3_D_REG_15__SCAN_IN, P3_D_REG_16__SCAN_IN, P3_D_REG_17__SCAN_IN, P3_D_REG_18__SCAN_IN, P3_D_REG_19__SCAN_IN, P3_D_REG_20__SCAN_IN, P3_D_REG_21__SCAN_IN, P3_D_REG_22__SCAN_IN, P3_D_REG_23__SCAN_IN, P3_D_REG_24__SCAN_IN, P3_D_REG_25__SCAN_IN, P3_D_REG_26__SCAN_IN, P3_D_REG_27__SCAN_IN, P3_D_REG_28__SCAN_IN, P3_D_REG_29__SCAN_IN, P3_D_REG_30__SCAN_IN, P3_D_REG_31__SCAN_IN, P3_REG0_REG_0__SCAN_IN, P3_REG0_REG_1__SCAN_IN, P3_REG0_REG_2__SCAN_IN, P3_REG0_REG_3__SCAN_IN, P3_REG0_REG_4__SCAN_IN, P3_REG0_REG_5__SCAN_IN, P3_REG0_REG_6__SCAN_IN, P3_REG0_REG_7__SCAN_IN, P3_REG0_REG_8__SCAN_IN, P3_REG0_REG_9__SCAN_IN, P3_REG0_REG_10__SCAN_IN, P3_REG0_REG_11__SCAN_IN, P3_REG0_REG_12__SCAN_IN, P3_REG0_REG_13__SCAN_IN, P3_REG0_REG_14__SCAN_IN, P3_REG0_REG_15__SCAN_IN, P3_REG0_REG_16__SCAN_IN, P3_REG0_REG_17__SCAN_IN, P3_REG0_REG_18__SCAN_IN, P3_REG0_REG_19__SCAN_IN, P3_REG0_REG_20__SCAN_IN, P3_REG0_REG_21__SCAN_IN, P3_REG0_REG_22__SCAN_IN, P3_REG0_REG_23__SCAN_IN, P3_REG0_REG_24__SCAN_IN, P3_REG0_REG_25__SCAN_IN, P3_REG0_REG_26__SCAN_IN, P3_REG0_REG_27__SCAN_IN, P3_REG0_REG_28__SCAN_IN, P3_REG0_REG_29__SCAN_IN, P3_REG0_REG_30__SCAN_IN, P3_REG0_REG_31__SCAN_IN, P3_REG1_REG_0__SCAN_IN, P3_REG1_REG_1__SCAN_IN, P3_REG1_REG_2__SCAN_IN, P3_REG1_REG_3__SCAN_IN, P3_REG1_REG_4__SCAN_IN, P3_REG1_REG_5__SCAN_IN, P3_REG1_REG_6__SCAN_IN, P3_REG1_REG_7__SCAN_IN, P3_REG1_REG_8__SCAN_IN, P3_REG1_REG_9__SCAN_IN, P3_REG1_REG_10__SCAN_IN, P3_REG1_REG_11__SCAN_IN, P3_REG1_REG_12__SCAN_IN, P3_REG1_REG_13__SCAN_IN, P3_REG1_REG_14__SCAN_IN, P3_REG1_REG_15__SCAN_IN, P3_REG1_REG_16__SCAN_IN, P3_REG1_REG_17__SCAN_IN, P3_REG1_REG_18__SCAN_IN, P3_REG1_REG_19__SCAN_IN, P3_REG1_REG_20__SCAN_IN, P3_REG1_REG_21__SCAN_IN, P3_REG1_REG_22__SCAN_IN, P3_REG1_REG_23__SCAN_IN, P3_REG1_REG_24__SCAN_IN, P3_REG1_REG_25__SCAN_IN, P3_REG1_REG_26__SCAN_IN, P3_REG1_REG_27__SCAN_IN, P3_REG1_REG_28__SCAN_IN, P3_REG1_REG_29__SCAN_IN, P3_REG1_REG_30__SCAN_IN, P3_REG1_REG_31__SCAN_IN, P3_REG2_REG_0__SCAN_IN, P3_REG2_REG_1__SCAN_IN, P3_REG2_REG_2__SCAN_IN, P3_REG2_REG_3__SCAN_IN, P3_REG2_REG_4__SCAN_IN, P3_REG2_REG_5__SCAN_IN, P3_REG2_REG_6__SCAN_IN, P3_REG2_REG_7__SCAN_IN, P3_REG2_REG_8__SCAN_IN, P3_REG2_REG_9__SCAN_IN, P3_REG2_REG_10__SCAN_IN, P3_REG2_REG_11__SCAN_IN, P3_REG2_REG_12__SCAN_IN, P3_REG2_REG_13__SCAN_IN, P3_REG2_REG_14__SCAN_IN, P3_REG2_REG_15__SCAN_IN, P3_REG2_REG_16__SCAN_IN, P3_REG2_REG_17__SCAN_IN, P3_REG2_REG_18__SCAN_IN, P3_REG2_REG_19__SCAN_IN, P3_REG2_REG_20__SCAN_IN, P3_REG2_REG_21__SCAN_IN, P3_REG2_REG_22__SCAN_IN, P3_REG2_REG_23__SCAN_IN, P3_REG2_REG_24__SCAN_IN, P3_REG2_REG_25__SCAN_IN, P3_REG2_REG_26__SCAN_IN, P3_REG2_REG_27__SCAN_IN, P3_REG2_REG_28__SCAN_IN, P3_REG2_REG_29__SCAN_IN, P3_REG2_REG_30__SCAN_IN, P3_REG2_REG_31__SCAN_IN, P3_ADDR_REG_19__SCAN_IN, P3_ADDR_REG_18__SCAN_IN, P3_ADDR_REG_17__SCAN_IN, P3_ADDR_REG_16__SCAN_IN, P3_ADDR_REG_15__SCAN_IN, P3_ADDR_REG_14__SCAN_IN, P3_ADDR_REG_13__SCAN_IN, P3_ADDR_REG_12__SCAN_IN, P3_ADDR_REG_11__SCAN_IN, P3_ADDR_REG_10__SCAN_IN, flip_signal, SUB_1596_U4, SUB_1596_U62, SUB_1596_U63, SUB_1596_U64, SUB_1596_U65, SUB_1596_U66, SUB_1596_U67, SUB_1596_U68, SUB_1596_U69, SUB_1596_U70, SUB_1596_U54, SUB_1596_U55, SUB_1596_U56, SUB_1596_U57, SUB_1596_U58, SUB_1596_U59, SUB_1596_U60, SUB_1596_U61, SUB_1596_U5, SUB_1596_U53, U29, U28, P1_U3355, P1_U3354, P1_U3353, P1_U3352, P1_U3351, P1_U3350, P1_U3349, P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, P1_U3343, P1_U3342, P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, P1_U3336, P1_U3335, P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, P1_U3329, P1_U3328, P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3445, P1_U3446, P1_U3323, P1_U3322, P1_U3321, P1_U3320, P1_U3319, P1_U3318, P1_U3317, P1_U3316, P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, P1_U3310, P1_U3309, P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, P1_U3303, P1_U3302, P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, P1_U3296, P1_U3295, P1_U3294, P1_U3459, P1_U3462, P1_U3465, P1_U3468, P1_U3471, P1_U3474, P1_U3477, P1_U3480, P1_U3483, P1_U3486, P1_U3489, P1_U3492, P1_U3495, P1_U3498, P1_U3501, P1_U3504, P1_U3507, P1_U3510, P1_U3513, P1_U3515, P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521, P1_U3522, P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528, P1_U3529, P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535, P1_U3536, P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542, P1_U3543, P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549, P1_U3550, P1_U3551, P1_U3552, P1_U3553, P1_U3554, P1_U3555, P1_U3556, P1_U3557, P1_U3558, P1_U3559, P1_U3293, P1_U3292, P1_U3291, P1_U3290, P1_U3289, P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, P1_U3283, P1_U3282, P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, P1_U3276, P1_U3275, P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, P1_U3269, P1_U3268, P1_U3267, P1_U3266, P1_U3265, P1_U3356, P1_U3264, P1_U3263, P1_U3262, P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, P1_U3256, P1_U3255, P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, P1_U3249, P1_U3248, P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, P1_U3560, P1_U3561, P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567, P1_U3568, P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574, P1_U3575, P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581, P1_U3582, P1_U3583, P1_U3584, P1_U3585, P1_U3586, P1_U3587, P1_U3588, P1_U3589, P1_U3590, P1_U3591, P1_U3242, P1_U3241, P1_U3240, P1_U3239, P1_U3238, P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, P1_U3232, P1_U3231, P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, P1_U3225, P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218, P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3086, P1_U3085, P1_U4016, P2_U3327, P2_U3326, P2_U3325, P2_U3324, P2_U3323, P2_U3322, P2_U3321, P2_U3320, P2_U3319, P2_U3318, P2_U3317, P2_U3316, P2_U3315, P2_U3314, P2_U3313, P2_U3312, P2_U3311, P2_U3310, P2_U3309, P2_U3308, P2_U3307, P2_U3306, P2_U3305, P2_U3304, P2_U3303, P2_U3302, P2_U3301, P2_U3300, P2_U3299, P2_U3298, P2_U3297, P2_U3296, P2_U3416, P2_U3417, P2_U3295, P2_U3294, P2_U3293, P2_U3292, P2_U3291, P2_U3290, P2_U3289, P2_U3288, P2_U3287, P2_U3286, P2_U3285, P2_U3284, P2_U3283, P2_U3282, P2_U3281, P2_U3280, P2_U3279, P2_U3278, P2_U3277, P2_U3276, P2_U3275, P2_U3274, P2_U3273, P2_U3272, P2_U3271, P2_U3270, P2_U3269, P2_U3268, P2_U3267, P2_U3266, P2_U3430, P2_U3433, P2_U3436, P2_U3439, P2_U3442, P2_U3445, P2_U3448, P2_U3451, P2_U3454, P2_U3457, P2_U3460, P2_U3463, P2_U3466, P2_U3469, P2_U3472, P2_U3475, P2_U3478, P2_U3481, P2_U3484, P2_U3486, P2_U3487, P2_U3488, P2_U3489, P2_U3490, P2_U3491, P2_U3492, P2_U3493, P2_U3494, P2_U3495, P2_U3496, P2_U3497, P2_U3498, P2_U3499, P2_U3500, P2_U3501, P2_U3502, P2_U3503, P2_U3504, P2_U3505, P2_U3506, P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511, P2_U3512, P2_U3513, P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518, P2_U3519, P2_U3520, P2_U3521, P2_U3522, P2_U3523, P2_U3524, P2_U3525, P2_U3526, P2_U3527, P2_U3528, P2_U3529, P2_U3530, P2_U3265, P2_U3264, P2_U3263, P2_U3262, P2_U3261, P2_U3260, P2_U3259, P2_U3258, P2_U3257, P2_U3256, P2_U3255, P2_U3254, P2_U3253, P2_U3252, P2_U3251, P2_U3250, P2_U3249, P2_U3248, P2_U3247, P2_U3246, P2_U3245, P2_U3244, P2_U3243, P2_U3242, P2_U3241, P2_U3240, P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234, P2_U3233, P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227, P2_U3226, P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220, P2_U3219, P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3214, P2_U3531, P2_U3532, P2_U3533, P2_U3534, P2_U3535, P2_U3536, P2_U3537, P2_U3538, P2_U3539, P2_U3540, P2_U3541, P2_U3542, P2_U3543, P2_U3544, P2_U3545, P2_U3546, P2_U3547, P2_U3548, P2_U3549, P2_U3550, P2_U3551, P2_U3552, P2_U3553, P2_U3554, P2_U3555, P2_U3556, P2_U3557, P2_U3558, P2_U3559, P2_U3560, P2_U3561, P2_U3562, P2_U3328, P2_U3213, P2_U3212, P2_U3211, P2_U3210, P2_U3209, P2_U3208, P2_U3207, P2_U3206, P2_U3205, P2_U3204, P2_U3203, P2_U3202, P2_U3201, P2_U3200, P2_U3199, P2_U3198, P2_U3197, P2_U3196, P2_U3195, P2_U3194, P2_U3193, P2_U3192, P2_U3191, P2_U3190, P2_U3189, P2_U3188, P2_U3187, P2_U3186, P2_U3185, P2_U3088, P2_U3087, P2_U3947, P3_U3295, P3_U3294, P3_U3293, P3_U3292, P3_U3291, P3_U3290, P3_U3289, P3_U3288, P3_U3287, P3_U3286, P3_U3285, P3_U3284, P3_U3283, P3_U3282, P3_U3281, P3_U3280, P3_U3279, P3_U3278, P3_U3277, P3_U3276, P3_U3275, P3_U3274, P3_U3273, P3_U3272, P3_U3271, P3_U3270, P3_U3269, P3_U3268, P3_U3267, P3_U3266, P3_U3265, P3_U3264, P3_U3376, P3_U3377, P3_U3263, P3_U3262, P3_U3261, P3_U3260, P3_U3259, P3_U3258, P3_U3257, P3_U3256, P3_U3255, P3_U3254, P3_U3253, P3_U3252, P3_U3251, P3_U3250, P3_U3249, P3_U3248, P3_U3247, P3_U3246, P3_U3245, P3_U3244, P3_U3243, P3_U3242, P3_U3241, P3_U3240, P3_U3239, P3_U3238, P3_U3237, P3_U3236, P3_U3235, P3_U3234, P3_U3390, P3_U3393, P3_U3396, P3_U3399, P3_U3402, P3_U3405, P3_U3408, P3_U3411, P3_U3414, P3_U3417, P3_U3420, P3_U3423, P3_U3426, P3_U3429, P3_U3432, P3_U3435, P3_U3438, P3_U3441, P3_U3444, P3_U3446, P3_U3447, P3_U3448, P3_U3449, P3_U3450, P3_U3451, P3_U3452, P3_U3453, P3_U3454, P3_U3455, P3_U3456, P3_U3457, P3_U3458, P3_U3459, P3_U3460, P3_U3461, P3_U3462, P3_U3463, P3_U3464, P3_U3465, P3_U3466, P3_U3467, P3_U3468, P3_U3469, P3_U3470, P3_U3471, P3_U3472, P3_U3473, P3_U3474, P3_U3475, P3_U3476, P3_U3477, P3_U3478, P3_U3479, P3_U3480, P3_U3481, P3_U3482, P3_U3483, P3_U3484, P3_U3485, P3_U3486, P3_U3487, P3_U3488, P3_U3489, P3_U3490, P3_U3233, P3_U3232, P3_U3231, P3_U3230, P3_U3229, P3_U3228, P3_U3227, P3_U3226, P3_U3225, P3_U3224, P3_U3223, P3_U3222, P3_U3221, P3_U3220, P3_U3219, P3_U3218, P3_U3217, P3_U3216, P3_U3215, P3_U3214, P3_U3213, P3_U3212, P3_U3211, P3_U3210, P3_U3209, P3_U3208, P3_U3207, P3_U3206, P3_U3205, P3_U3204, P3_U3203, P3_U3202, P3_U3201, P3_U3200, P3_U3199, P3_U3198, P3_U3197, P3_U3196, P3_U3195, P3_U3194, P3_U3193, P3_U3192, P3_U3191, P3_U3190, P3_U3189, P3_U3188, P3_U3187, P3_U3186, P3_U3185, P3_U3184, P3_U3183, P3_U3182, P3_U3491, P3_U3492, P3_U3493, P3_U3494, P3_U3495, P3_U3496, P3_U3497, P3_U3498, P3_U3499, P3_U3500, P3_U3501, P3_U3502, P3_U3503, P3_U3504, P3_U3505, P3_U3506, P3_U3507, P3_U3508, P3_U3509, P3_U3510, P3_U3511, P3_U3512, P3_U3513, P3_U3514, P3_U3515, P3_U3516, P3_U3517, P3_U3518, P3_U3519, P3_U3520, P3_U3521, P3_U3522, P3_U3296, P3_U3181, P3_U3180, P3_U3179, P3_U3178, P3_U3177, P3_U3176, P3_U3175, P3_U3174, P3_U3173, P3_U3172, P3_U3171, P3_U3170, P3_U3169, P3_U3168, P3_U3167, P3_U3166, P3_U3165, P3_U3164, P3_U3163, P3_U3162, P3_U3161, P3_U3160, P3_U3159, P3_U3158, P3_U3157, P3_U3156, P3_U3155, P3_U3154, P3_U3153, P3_U3151, P3_U3150, P3_U3897);

  input P3_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, SI_28_, SI_27_, SI_26_, SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, SI_19_, SI_18_, SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, SI_10_, SI_9_, SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, SI_0_, P3_RD_REG_SCAN_IN, P3_STATE_REG_SCAN_IN, P3_REG3_REG_7__SCAN_IN, P3_REG3_REG_27__SCAN_IN, P3_REG3_REG_14__SCAN_IN, P3_REG3_REG_23__SCAN_IN, P3_REG3_REG_10__SCAN_IN, P3_REG3_REG_3__SCAN_IN, P3_REG3_REG_19__SCAN_IN, P3_REG3_REG_28__SCAN_IN, P3_REG3_REG_8__SCAN_IN, P3_REG3_REG_1__SCAN_IN, P3_REG3_REG_21__SCAN_IN, P3_REG3_REG_12__SCAN_IN, P3_REG3_REG_25__SCAN_IN, P3_REG3_REG_16__SCAN_IN, P3_REG3_REG_5__SCAN_IN, P3_REG3_REG_17__SCAN_IN, P3_REG3_REG_24__SCAN_IN, P3_REG3_REG_4__SCAN_IN, P3_REG3_REG_9__SCAN_IN, P3_REG3_REG_0__SCAN_IN, P3_REG3_REG_20__SCAN_IN, P3_REG3_REG_13__SCAN_IN, P3_REG3_REG_22__SCAN_IN, P3_REG3_REG_11__SCAN_IN, P3_REG3_REG_2__SCAN_IN, P3_REG3_REG_18__SCAN_IN, P3_REG3_REG_6__SCAN_IN, P3_REG3_REG_26__SCAN_IN, P3_REG3_REG_15__SCAN_IN, P3_B_REG_SCAN_IN, P3_DATAO_REG_31__SCAN_IN, P3_DATAO_REG_30__SCAN_IN, P3_DATAO_REG_29__SCAN_IN, P3_DATAO_REG_28__SCAN_IN, P3_DATAO_REG_27__SCAN_IN, P3_DATAO_REG_26__SCAN_IN, P3_DATAO_REG_25__SCAN_IN, P3_DATAO_REG_24__SCAN_IN, P3_DATAO_REG_23__SCAN_IN, P3_DATAO_REG_22__SCAN_IN, P3_DATAO_REG_21__SCAN_IN, P3_DATAO_REG_20__SCAN_IN, P3_DATAO_REG_19__SCAN_IN, P3_DATAO_REG_18__SCAN_IN, P3_DATAO_REG_17__SCAN_IN, P3_DATAO_REG_16__SCAN_IN, P3_DATAO_REG_15__SCAN_IN, P3_DATAO_REG_14__SCAN_IN, P3_DATAO_REG_13__SCAN_IN, P3_DATAO_REG_12__SCAN_IN, P3_DATAO_REG_11__SCAN_IN, P3_DATAO_REG_10__SCAN_IN, P3_DATAO_REG_9__SCAN_IN, P3_DATAO_REG_8__SCAN_IN, P3_DATAO_REG_7__SCAN_IN, P3_DATAO_REG_6__SCAN_IN, P3_DATAO_REG_5__SCAN_IN, P3_DATAO_REG_4__SCAN_IN, P3_DATAO_REG_3__SCAN_IN, P3_DATAO_REG_2__SCAN_IN, P3_DATAO_REG_1__SCAN_IN, P3_DATAO_REG_0__SCAN_IN, P3_ADDR_REG_0__SCAN_IN, P3_ADDR_REG_1__SCAN_IN, P3_ADDR_REG_2__SCAN_IN, P3_ADDR_REG_3__SCAN_IN, P3_ADDR_REG_4__SCAN_IN, P3_ADDR_REG_5__SCAN_IN, P3_ADDR_REG_6__SCAN_IN, P3_ADDR_REG_7__SCAN_IN, P3_ADDR_REG_8__SCAN_IN, P3_ADDR_REG_9__SCAN_IN, P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN, P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN, P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN, P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN, P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN, P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN, P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN, P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN, P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN, P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN, P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN, P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN, P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN, P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN, P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN, P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN, P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN, P1_REG1_REG_3__SCAN_IN, P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN, P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN, P1_REG1_REG_9__SCAN_IN, P1_REG1_REG_10__SCAN_IN, P1_REG1_REG_11__SCAN_IN, P1_REG1_REG_12__SCAN_IN, P1_REG1_REG_13__SCAN_IN, P1_REG1_REG_14__SCAN_IN, P1_REG1_REG_15__SCAN_IN, P1_REG1_REG_16__SCAN_IN, P1_REG1_REG_17__SCAN_IN, P1_REG1_REG_18__SCAN_IN, P1_REG1_REG_19__SCAN_IN, P1_REG1_REG_20__SCAN_IN, P1_REG1_REG_21__SCAN_IN, P1_REG1_REG_22__SCAN_IN, P1_REG1_REG_23__SCAN_IN, P1_REG1_REG_24__SCAN_IN, P1_REG1_REG_25__SCAN_IN, P1_REG1_REG_26__SCAN_IN, P1_REG1_REG_27__SCAN_IN, P1_REG1_REG_28__SCAN_IN, P1_REG1_REG_29__SCAN_IN, P1_REG1_REG_30__SCAN_IN, P1_REG1_REG_31__SCAN_IN, P1_REG2_REG_0__SCAN_IN, P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN, P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN, P1_REG2_REG_6__SCAN_IN, P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN, P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN, P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN, P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN, P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN, P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN, P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN, P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN, P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN, P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN, P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN, P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN, P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN, P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN, P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN, P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN, P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN, P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN, P1_ADDR_REG_6__SCAN_IN, P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN, P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN, P1_ADDR_REG_0__SCAN_IN, P1_DATAO_REG_0__SCAN_IN, P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, P1_REG3_REG_15__SCAN_IN, P1_REG3_REG_26__SCAN_IN, P1_REG3_REG_6__SCAN_IN, P1_REG3_REG_18__SCAN_IN, P1_REG3_REG_2__SCAN_IN, P1_REG3_REG_11__SCAN_IN, P1_REG3_REG_22__SCAN_IN, P1_REG3_REG_13__SCAN_IN, P1_REG3_REG_20__SCAN_IN, P1_REG3_REG_0__SCAN_IN, P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN, P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN, P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN, P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN, P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN, P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN, P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN, P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN, P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN, P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN, P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN, P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN, P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN, P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN, P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN, P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN, P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN, P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN, P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN, P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN, P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN, P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN, P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN, P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN, P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN, P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN, P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN, P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN, P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN, P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN, P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN, P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN, P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN, P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN, P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN, P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN, P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN, P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN, P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN, P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN, P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN, P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN, P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN, P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN, P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN, P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN, P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN, P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN, P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN, P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN, P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN, P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN, P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN, P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN, P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN, P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN, P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN, P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN, P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN, P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN, P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN, P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN, P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN, P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN, P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN, P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN, P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN, P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN, P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN, P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN, P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN, P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN, P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN, P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN, P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN, P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN, P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN, P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN, P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN, P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN, P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN, P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN, P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN, P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN, P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN, P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN, P2_DATAO_REG_5__SCAN_IN, P2_DATAO_REG_6__SCAN_IN, P2_DATAO_REG_7__SCAN_IN, P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_9__SCAN_IN, P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_11__SCAN_IN, P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_13__SCAN_IN, P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_15__SCAN_IN, P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_17__SCAN_IN, P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_19__SCAN_IN, P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_21__SCAN_IN, P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_23__SCAN_IN, P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_25__SCAN_IN, P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_27__SCAN_IN, P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_29__SCAN_IN, P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_31__SCAN_IN, P2_B_REG_SCAN_IN, P2_REG3_REG_15__SCAN_IN, P2_REG3_REG_26__SCAN_IN, P2_REG3_REG_6__SCAN_IN, P2_REG3_REG_18__SCAN_IN, P2_REG3_REG_2__SCAN_IN, P2_REG3_REG_11__SCAN_IN, P2_REG3_REG_22__SCAN_IN, P2_REG3_REG_13__SCAN_IN, P2_REG3_REG_20__SCAN_IN, P2_REG3_REG_0__SCAN_IN, P2_REG3_REG_9__SCAN_IN, P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_24__SCAN_IN, P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_5__SCAN_IN, P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_25__SCAN_IN, P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_21__SCAN_IN, P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_8__SCAN_IN, P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_19__SCAN_IN, P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_10__SCAN_IN, P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_14__SCAN_IN, P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_7__SCAN_IN, P2_STATE_REG_SCAN_IN, P2_RD_REG_SCAN_IN, P2_WR_REG_SCAN_IN, P3_IR_REG_0__SCAN_IN, P3_IR_REG_1__SCAN_IN, P3_IR_REG_2__SCAN_IN, P3_IR_REG_3__SCAN_IN, P3_IR_REG_4__SCAN_IN, P3_IR_REG_5__SCAN_IN, P3_IR_REG_6__SCAN_IN, P3_IR_REG_7__SCAN_IN, P3_IR_REG_8__SCAN_IN, P3_IR_REG_9__SCAN_IN, P3_IR_REG_10__SCAN_IN, P3_IR_REG_11__SCAN_IN, P3_IR_REG_12__SCAN_IN, P3_IR_REG_13__SCAN_IN, P3_IR_REG_14__SCAN_IN, P3_IR_REG_15__SCAN_IN, P3_IR_REG_16__SCAN_IN, P3_IR_REG_17__SCAN_IN, P3_IR_REG_18__SCAN_IN, P3_IR_REG_19__SCAN_IN, P3_IR_REG_20__SCAN_IN, P3_IR_REG_21__SCAN_IN, P3_IR_REG_22__SCAN_IN, P3_IR_REG_23__SCAN_IN, P3_IR_REG_24__SCAN_IN, P3_IR_REG_25__SCAN_IN, P3_IR_REG_26__SCAN_IN, P3_IR_REG_27__SCAN_IN, P3_IR_REG_28__SCAN_IN, P3_IR_REG_29__SCAN_IN, P3_IR_REG_30__SCAN_IN, P3_IR_REG_31__SCAN_IN, P3_D_REG_0__SCAN_IN, P3_D_REG_1__SCAN_IN, P3_D_REG_2__SCAN_IN, P3_D_REG_3__SCAN_IN, P3_D_REG_4__SCAN_IN, P3_D_REG_5__SCAN_IN, P3_D_REG_6__SCAN_IN, P3_D_REG_7__SCAN_IN, P3_D_REG_8__SCAN_IN, P3_D_REG_9__SCAN_IN, P3_D_REG_10__SCAN_IN, P3_D_REG_11__SCAN_IN, P3_D_REG_12__SCAN_IN, P3_D_REG_13__SCAN_IN, P3_D_REG_14__SCAN_IN, P3_D_REG_15__SCAN_IN, P3_D_REG_16__SCAN_IN, P3_D_REG_17__SCAN_IN, P3_D_REG_18__SCAN_IN, P3_D_REG_19__SCAN_IN, P3_D_REG_20__SCAN_IN, P3_D_REG_21__SCAN_IN, P3_D_REG_22__SCAN_IN, P3_D_REG_23__SCAN_IN, P3_D_REG_24__SCAN_IN, P3_D_REG_25__SCAN_IN, P3_D_REG_26__SCAN_IN, P3_D_REG_27__SCAN_IN, P3_D_REG_28__SCAN_IN, P3_D_REG_29__SCAN_IN, P3_D_REG_30__SCAN_IN, P3_D_REG_31__SCAN_IN, P3_REG0_REG_0__SCAN_IN, P3_REG0_REG_1__SCAN_IN, P3_REG0_REG_2__SCAN_IN, P3_REG0_REG_3__SCAN_IN, P3_REG0_REG_4__SCAN_IN, P3_REG0_REG_5__SCAN_IN, P3_REG0_REG_6__SCAN_IN, P3_REG0_REG_7__SCAN_IN, P3_REG0_REG_8__SCAN_IN, P3_REG0_REG_9__SCAN_IN, P3_REG0_REG_10__SCAN_IN, P3_REG0_REG_11__SCAN_IN, P3_REG0_REG_12__SCAN_IN, P3_REG0_REG_13__SCAN_IN, P3_REG0_REG_14__SCAN_IN, P3_REG0_REG_15__SCAN_IN, P3_REG0_REG_16__SCAN_IN, P3_REG0_REG_17__SCAN_IN, P3_REG0_REG_18__SCAN_IN, P3_REG0_REG_19__SCAN_IN, P3_REG0_REG_20__SCAN_IN, P3_REG0_REG_21__SCAN_IN, P3_REG0_REG_22__SCAN_IN, P3_REG0_REG_23__SCAN_IN, P3_REG0_REG_24__SCAN_IN, P3_REG0_REG_25__SCAN_IN, P3_REG0_REG_26__SCAN_IN, P3_REG0_REG_27__SCAN_IN, P3_REG0_REG_28__SCAN_IN, P3_REG0_REG_29__SCAN_IN, P3_REG0_REG_30__SCAN_IN, P3_REG0_REG_31__SCAN_IN, P3_REG1_REG_0__SCAN_IN, P3_REG1_REG_1__SCAN_IN, P3_REG1_REG_2__SCAN_IN, P3_REG1_REG_3__SCAN_IN, P3_REG1_REG_4__SCAN_IN, P3_REG1_REG_5__SCAN_IN, P3_REG1_REG_6__SCAN_IN, P3_REG1_REG_7__SCAN_IN, P3_REG1_REG_8__SCAN_IN, P3_REG1_REG_9__SCAN_IN, P3_REG1_REG_10__SCAN_IN, P3_REG1_REG_11__SCAN_IN, P3_REG1_REG_12__SCAN_IN, P3_REG1_REG_13__SCAN_IN, P3_REG1_REG_14__SCAN_IN, P3_REG1_REG_15__SCAN_IN, P3_REG1_REG_16__SCAN_IN, P3_REG1_REG_17__SCAN_IN, P3_REG1_REG_18__SCAN_IN, P3_REG1_REG_19__SCAN_IN, P3_REG1_REG_20__SCAN_IN, P3_REG1_REG_21__SCAN_IN, P3_REG1_REG_22__SCAN_IN, P3_REG1_REG_23__SCAN_IN, P3_REG1_REG_24__SCAN_IN, P3_REG1_REG_25__SCAN_IN, P3_REG1_REG_26__SCAN_IN, P3_REG1_REG_27__SCAN_IN, P3_REG1_REG_28__SCAN_IN, P3_REG1_REG_29__SCAN_IN, P3_REG1_REG_30__SCAN_IN, P3_REG1_REG_31__SCAN_IN, P3_REG2_REG_0__SCAN_IN, P3_REG2_REG_1__SCAN_IN, P3_REG2_REG_2__SCAN_IN, P3_REG2_REG_3__SCAN_IN, P3_REG2_REG_4__SCAN_IN, P3_REG2_REG_5__SCAN_IN, P3_REG2_REG_6__SCAN_IN, P3_REG2_REG_7__SCAN_IN, P3_REG2_REG_8__SCAN_IN, P3_REG2_REG_9__SCAN_IN, P3_REG2_REG_10__SCAN_IN, P3_REG2_REG_11__SCAN_IN, P3_REG2_REG_12__SCAN_IN, P3_REG2_REG_13__SCAN_IN, P3_REG2_REG_14__SCAN_IN, P3_REG2_REG_15__SCAN_IN, P3_REG2_REG_16__SCAN_IN, P3_REG2_REG_17__SCAN_IN, P3_REG2_REG_18__SCAN_IN, P3_REG2_REG_19__SCAN_IN, P3_REG2_REG_20__SCAN_IN, P3_REG2_REG_21__SCAN_IN, P3_REG2_REG_22__SCAN_IN, P3_REG2_REG_23__SCAN_IN, P3_REG2_REG_24__SCAN_IN, P3_REG2_REG_25__SCAN_IN, P3_REG2_REG_26__SCAN_IN, P3_REG2_REG_27__SCAN_IN, P3_REG2_REG_28__SCAN_IN, P3_REG2_REG_29__SCAN_IN, P3_REG2_REG_30__SCAN_IN, P3_REG2_REG_31__SCAN_IN, P3_ADDR_REG_19__SCAN_IN, P3_ADDR_REG_18__SCAN_IN, P3_ADDR_REG_17__SCAN_IN, P3_ADDR_REG_16__SCAN_IN, P3_ADDR_REG_15__SCAN_IN, P3_ADDR_REG_14__SCAN_IN, P3_ADDR_REG_13__SCAN_IN, P3_ADDR_REG_12__SCAN_IN, P3_ADDR_REG_11__SCAN_IN, P3_ADDR_REG_10__SCAN_IN, flip_signal;
  output SUB_1596_U4, SUB_1596_U62, SUB_1596_U63, SUB_1596_U64, SUB_1596_U65, SUB_1596_U66, SUB_1596_U67, SUB_1596_U68, SUB_1596_U69, SUB_1596_U70, SUB_1596_U54, SUB_1596_U55, SUB_1596_U56, SUB_1596_U57, SUB_1596_U58, SUB_1596_U59, SUB_1596_U60, SUB_1596_U61, SUB_1596_U5, SUB_1596_U53, U29, U28, P1_U3355, P1_U3354, P1_U3353, P1_U3352, P1_U3351, P1_U3350, P1_U3349, P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, P1_U3343, P1_U3342, P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, P1_U3336, P1_U3335, P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, P1_U3329, P1_U3328, P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3445, P1_U3446, P1_U3323, P1_U3322, P1_U3321, P1_U3320, P1_U3319, P1_U3318, P1_U3317, P1_U3316, P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, P1_U3310, P1_U3309, P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, P1_U3303, P1_U3302, P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, P1_U3296, P1_U3295, P1_U3294, P1_U3459, P1_U3462, P1_U3465, P1_U3468, P1_U3471, P1_U3474, P1_U3477, P1_U3480, P1_U3483, P1_U3486, P1_U3489, P1_U3492, P1_U3495, P1_U3498, P1_U3501, P1_U3504, P1_U3507, P1_U3510, P1_U3513, P1_U3515, P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521, P1_U3522, P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528, P1_U3529, P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535, P1_U3536, P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542, P1_U3543, P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549, P1_U3550, P1_U3551, P1_U3552, P1_U3553, P1_U3554, P1_U3555, P1_U3556, P1_U3557, P1_U3558, P1_U3559, P1_U3293, P1_U3292, P1_U3291, P1_U3290, P1_U3289, P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, P1_U3283, P1_U3282, P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, P1_U3276, P1_U3275, P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, P1_U3269, P1_U3268, P1_U3267, P1_U3266, P1_U3265, P1_U3356, P1_U3264, P1_U3263, P1_U3262, P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, P1_U3256, P1_U3255, P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, P1_U3249, P1_U3248, P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, P1_U3560, P1_U3561, P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567, P1_U3568, P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574, P1_U3575, P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581, P1_U3582, P1_U3583, P1_U3584, P1_U3585, P1_U3586, P1_U3587, P1_U3588, P1_U3589, P1_U3590, P1_U3591, P1_U3242, P1_U3241, P1_U3240, P1_U3239, P1_U3238, P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, P1_U3232, P1_U3231, P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, P1_U3225, P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218, P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3086, P1_U3085, P1_U4016, P2_U3327, P2_U3326, P2_U3325, P2_U3324, P2_U3323, P2_U3322, P2_U3321, P2_U3320, P2_U3319, P2_U3318, P2_U3317, P2_U3316, P2_U3315, P2_U3314, P2_U3313, P2_U3312, P2_U3311, P2_U3310, P2_U3309, P2_U3308, P2_U3307, P2_U3306, P2_U3305, P2_U3304, P2_U3303, P2_U3302, P2_U3301, P2_U3300, P2_U3299, P2_U3298, P2_U3297, P2_U3296, P2_U3416, P2_U3417, P2_U3295, P2_U3294, P2_U3293, P2_U3292, P2_U3291, P2_U3290, P2_U3289, P2_U3288, P2_U3287, P2_U3286, P2_U3285, P2_U3284, P2_U3283, P2_U3282, P2_U3281, P2_U3280, P2_U3279, P2_U3278, P2_U3277, P2_U3276, P2_U3275, P2_U3274, P2_U3273, P2_U3272, P2_U3271, P2_U3270, P2_U3269, P2_U3268, P2_U3267, P2_U3266, P2_U3430, P2_U3433, P2_U3436, P2_U3439, P2_U3442, P2_U3445, P2_U3448, P2_U3451, P2_U3454, P2_U3457, P2_U3460, P2_U3463, P2_U3466, P2_U3469, P2_U3472, P2_U3475, P2_U3478, P2_U3481, P2_U3484, P2_U3486, P2_U3487, P2_U3488, P2_U3489, P2_U3490, P2_U3491, P2_U3492, P2_U3493, P2_U3494, P2_U3495, P2_U3496, P2_U3497, P2_U3498, P2_U3499, P2_U3500, P2_U3501, P2_U3502, P2_U3503, P2_U3504, P2_U3505, P2_U3506, P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511, P2_U3512, P2_U3513, P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518, P2_U3519, P2_U3520, P2_U3521, P2_U3522, P2_U3523, P2_U3524, P2_U3525, P2_U3526, P2_U3527, P2_U3528, P2_U3529, P2_U3530, P2_U3265, P2_U3264, P2_U3263, P2_U3262, P2_U3261, P2_U3260, P2_U3259, P2_U3258, P2_U3257, P2_U3256, P2_U3255, P2_U3254, P2_U3253, P2_U3252, P2_U3251, P2_U3250, P2_U3249, P2_U3248, P2_U3247, P2_U3246, P2_U3245, P2_U3244, P2_U3243, P2_U3242, P2_U3241, P2_U3240, P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234, P2_U3233, P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227, P2_U3226, P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220, P2_U3219, P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3214, P2_U3531, P2_U3532, P2_U3533, P2_U3534, P2_U3535, P2_U3536, P2_U3537, P2_U3538, P2_U3539, P2_U3540, P2_U3541, P2_U3542, P2_U3543, P2_U3544, P2_U3545, P2_U3546, P2_U3547, P2_U3548, P2_U3549, P2_U3550, P2_U3551, P2_U3552, P2_U3553, P2_U3554, P2_U3555, P2_U3556, P2_U3557, P2_U3558, P2_U3559, P2_U3560, P2_U3561, P2_U3562, P2_U3328, P2_U3213, P2_U3212, P2_U3211, P2_U3210, P2_U3209, P2_U3208, P2_U3207, P2_U3206, P2_U3205, P2_U3204, P2_U3203, P2_U3202, P2_U3201, P2_U3200, P2_U3199, P2_U3198, P2_U3197, P2_U3196, P2_U3195, P2_U3194, P2_U3193, P2_U3192, P2_U3191, P2_U3190, P2_U3189, P2_U3188, P2_U3187, P2_U3186, P2_U3185, P2_U3088, P2_U3087, P2_U3947, P3_U3295, P3_U3294, P3_U3293, P3_U3292, P3_U3291, P3_U3290, P3_U3289, P3_U3288, P3_U3287, P3_U3286, P3_U3285, P3_U3284, P3_U3283, P3_U3282, P3_U3281, P3_U3280, P3_U3279, P3_U3278, P3_U3277, P3_U3276, P3_U3275, P3_U3274, P3_U3273, P3_U3272, P3_U3271, P3_U3270, P3_U3269, P3_U3268, P3_U3267, P3_U3266, P3_U3265, P3_U3264, P3_U3376, P3_U3377, P3_U3263, P3_U3262, P3_U3261, P3_U3260, P3_U3259, P3_U3258, P3_U3257, P3_U3256, P3_U3255, P3_U3254, P3_U3253, P3_U3252, P3_U3251, P3_U3250, P3_U3249, P3_U3248, P3_U3247, P3_U3246, P3_U3245, P3_U3244, P3_U3243, P3_U3242, P3_U3241, P3_U3240, P3_U3239, P3_U3238, P3_U3237, P3_U3236, P3_U3235, P3_U3234, P3_U3390, P3_U3393, P3_U3396, P3_U3399, P3_U3402, P3_U3405, P3_U3408, P3_U3411, P3_U3414, P3_U3417, P3_U3420, P3_U3423, P3_U3426, P3_U3429, P3_U3432, P3_U3435, P3_U3438, P3_U3441, P3_U3444, P3_U3446, P3_U3447, P3_U3448, P3_U3449, P3_U3450, P3_U3451, P3_U3452, P3_U3453, P3_U3454, P3_U3455, P3_U3456, P3_U3457, P3_U3458, P3_U3459, P3_U3460, P3_U3461, P3_U3462, P3_U3463, P3_U3464, P3_U3465, P3_U3466, P3_U3467, P3_U3468, P3_U3469, P3_U3470, P3_U3471, P3_U3472, P3_U3473, P3_U3474, P3_U3475, P3_U3476, P3_U3477, P3_U3478, P3_U3479, P3_U3480, P3_U3481, P3_U3482, P3_U3483, P3_U3484, P3_U3485, P3_U3486, P3_U3487, P3_U3488, P3_U3489, P3_U3490, P3_U3233, P3_U3232, P3_U3231, P3_U3230, P3_U3229, P3_U3228, P3_U3227, P3_U3226, P3_U3225, P3_U3224, P3_U3223, P3_U3222, P3_U3221, P3_U3220, P3_U3219, P3_U3218, P3_U3217, P3_U3216, P3_U3215, P3_U3214, P3_U3213, P3_U3212, P3_U3211, P3_U3210, P3_U3209, P3_U3208, P3_U3207, P3_U3206, P3_U3205, P3_U3204, P3_U3203, P3_U3202, P3_U3201, P3_U3200, P3_U3199, P3_U3198, P3_U3197, P3_U3196, P3_U3195, P3_U3194, P3_U3193, P3_U3192, P3_U3191, P3_U3190, P3_U3189, P3_U3188, P3_U3187, P3_U3186, P3_U3185, P3_U3184, P3_U3183, P3_U3182, P3_U3491, P3_U3492, P3_U3493, P3_U3494, P3_U3495, P3_U3496, P3_U3497, P3_U3498, P3_U3499, P3_U3500, P3_U3501, P3_U3502, P3_U3503, P3_U3504, P3_U3505, P3_U3506, P3_U3507, P3_U3508, P3_U3509, P3_U3510, P3_U3511, P3_U3512, P3_U3513, P3_U3514, P3_U3515, P3_U3516, P3_U3517, P3_U3518, P3_U3519, P3_U3520, P3_U3521, P3_U3522, P3_U3296, P3_U3181, P3_U3180, P3_U3179, P3_U3178, P3_U3177, P3_U3176, P3_U3175, P3_U3174, P3_U3173, P3_U3172, P3_U3171, P3_U3170, P3_U3169, P3_U3168, P3_U3167, P3_U3166, P3_U3165, P3_U3164, P3_U3163, P3_U3162, P3_U3161, P3_U3160, P3_U3159, P3_U3158, P3_U3157, P3_U3156, P3_U3155, P3_U3154, P3_U3153, P3_U3151, P3_U3150, P3_U3897;
  wire ADD_1596_U10, ADD_1596_U100, ADD_1596_U101, ADD_1596_U102, ADD_1596_U103, ADD_1596_U104, ADD_1596_U105, ADD_1596_U106, ADD_1596_U107, ADD_1596_U108, ADD_1596_U109, ADD_1596_U11, ADD_1596_U110, ADD_1596_U111, ADD_1596_U112, ADD_1596_U113, ADD_1596_U114, ADD_1596_U115, ADD_1596_U116, ADD_1596_U117, ADD_1596_U118, ADD_1596_U119, ADD_1596_U12, ADD_1596_U120, ADD_1596_U121, ADD_1596_U122, ADD_1596_U123, ADD_1596_U124, ADD_1596_U125, ADD_1596_U126, ADD_1596_U127, ADD_1596_U128, ADD_1596_U129, ADD_1596_U13, ADD_1596_U130, ADD_1596_U131, ADD_1596_U132, ADD_1596_U133, ADD_1596_U134, ADD_1596_U135, ADD_1596_U136, ADD_1596_U137, ADD_1596_U138, ADD_1596_U139, ADD_1596_U14, ADD_1596_U140, ADD_1596_U141, ADD_1596_U142, ADD_1596_U143, ADD_1596_U144, ADD_1596_U145, ADD_1596_U146, ADD_1596_U147, ADD_1596_U148, ADD_1596_U149, ADD_1596_U15, ADD_1596_U150, ADD_1596_U151, ADD_1596_U152, ADD_1596_U153, ADD_1596_U154, ADD_1596_U155, ADD_1596_U156, ADD_1596_U157, ADD_1596_U158, ADD_1596_U159, ADD_1596_U16, ADD_1596_U160, ADD_1596_U161, ADD_1596_U162, ADD_1596_U163, ADD_1596_U164, ADD_1596_U165, ADD_1596_U166, ADD_1596_U167, ADD_1596_U168, ADD_1596_U169, ADD_1596_U17, ADD_1596_U170, ADD_1596_U171, ADD_1596_U172, ADD_1596_U173, ADD_1596_U174, ADD_1596_U175, ADD_1596_U176, ADD_1596_U177, ADD_1596_U178, ADD_1596_U179, ADD_1596_U18, ADD_1596_U180, ADD_1596_U181, ADD_1596_U182, ADD_1596_U183, ADD_1596_U184, ADD_1596_U185, ADD_1596_U186, ADD_1596_U187, ADD_1596_U188, ADD_1596_U189, ADD_1596_U19, ADD_1596_U190, ADD_1596_U191, ADD_1596_U192, ADD_1596_U193, ADD_1596_U194, ADD_1596_U195, ADD_1596_U196, ADD_1596_U197, ADD_1596_U198, ADD_1596_U199, ADD_1596_U20, ADD_1596_U200, ADD_1596_U201, ADD_1596_U202, ADD_1596_U203, ADD_1596_U204, ADD_1596_U205, ADD_1596_U206, ADD_1596_U207, ADD_1596_U208, ADD_1596_U209, ADD_1596_U21, ADD_1596_U210, ADD_1596_U211, ADD_1596_U212, ADD_1596_U213, ADD_1596_U214, ADD_1596_U215, ADD_1596_U216, ADD_1596_U217, ADD_1596_U218, ADD_1596_U219, ADD_1596_U22, ADD_1596_U220, ADD_1596_U221, ADD_1596_U222, ADD_1596_U223, ADD_1596_U224, ADD_1596_U225, ADD_1596_U226, ADD_1596_U227, ADD_1596_U228, ADD_1596_U229, ADD_1596_U23, ADD_1596_U230, ADD_1596_U231, ADD_1596_U232, ADD_1596_U233, ADD_1596_U234, ADD_1596_U235, ADD_1596_U236, ADD_1596_U237, ADD_1596_U238, ADD_1596_U239, ADD_1596_U24, ADD_1596_U240, ADD_1596_U241, ADD_1596_U242, ADD_1596_U243, ADD_1596_U244, ADD_1596_U245, ADD_1596_U246, ADD_1596_U247, ADD_1596_U248, ADD_1596_U249, ADD_1596_U25, ADD_1596_U250, ADD_1596_U251, ADD_1596_U252, ADD_1596_U253, ADD_1596_U254, ADD_1596_U255, ADD_1596_U256, ADD_1596_U257, ADD_1596_U258, ADD_1596_U259, ADD_1596_U26, ADD_1596_U260, ADD_1596_U261, ADD_1596_U262, ADD_1596_U263, ADD_1596_U264, ADD_1596_U265, ADD_1596_U266, ADD_1596_U267, ADD_1596_U268, ADD_1596_U269, ADD_1596_U27, ADD_1596_U270, ADD_1596_U271, ADD_1596_U272, ADD_1596_U273, ADD_1596_U274, ADD_1596_U28, ADD_1596_U29, ADD_1596_U30, ADD_1596_U31, ADD_1596_U32, ADD_1596_U33, ADD_1596_U34, ADD_1596_U35, ADD_1596_U36, ADD_1596_U37, ADD_1596_U38, ADD_1596_U39, ADD_1596_U40, ADD_1596_U41, ADD_1596_U42, ADD_1596_U43, ADD_1596_U44, ADD_1596_U45, ADD_1596_U46, ADD_1596_U47, ADD_1596_U48, ADD_1596_U49, ADD_1596_U50, ADD_1596_U51, ADD_1596_U52, ADD_1596_U53, ADD_1596_U54, ADD_1596_U55, ADD_1596_U56, ADD_1596_U57, ADD_1596_U58, ADD_1596_U59, ADD_1596_U6, ADD_1596_U60, ADD_1596_U61, ADD_1596_U62, ADD_1596_U63, ADD_1596_U64, ADD_1596_U65, ADD_1596_U66, ADD_1596_U67, ADD_1596_U68, ADD_1596_U69, ADD_1596_U7, ADD_1596_U70, ADD_1596_U71, ADD_1596_U72, ADD_1596_U73, ADD_1596_U74, ADD_1596_U75, ADD_1596_U76, ADD_1596_U77, ADD_1596_U78, ADD_1596_U79, ADD_1596_U8, ADD_1596_U80, ADD_1596_U81, ADD_1596_U82, ADD_1596_U83, ADD_1596_U84, ADD_1596_U85, ADD_1596_U86, ADD_1596_U87, ADD_1596_U88, ADD_1596_U89, ADD_1596_U9, ADD_1596_U90, ADD_1596_U91, ADD_1596_U92, ADD_1596_U93, ADD_1596_U94, ADD_1596_U95, ADD_1596_U96, ADD_1596_U97, ADD_1596_U98, ADD_1596_U99, LT_1601_21_U6, LT_1601_U6, LT_1602_U6, P1_ADD_99_U10, P1_ADD_99_U100, P1_ADD_99_U101, P1_ADD_99_U102, P1_ADD_99_U103, P1_ADD_99_U104, P1_ADD_99_U105, P1_ADD_99_U106, P1_ADD_99_U107, P1_ADD_99_U108, P1_ADD_99_U109, P1_ADD_99_U11, P1_ADD_99_U110, P1_ADD_99_U111, P1_ADD_99_U112, P1_ADD_99_U113, P1_ADD_99_U114, P1_ADD_99_U115, P1_ADD_99_U116, P1_ADD_99_U117, P1_ADD_99_U118, P1_ADD_99_U119, P1_ADD_99_U12, P1_ADD_99_U120, P1_ADD_99_U121, P1_ADD_99_U122, P1_ADD_99_U123, P1_ADD_99_U124, P1_ADD_99_U125, P1_ADD_99_U126, P1_ADD_99_U127, P1_ADD_99_U128, P1_ADD_99_U129, P1_ADD_99_U13, P1_ADD_99_U130, P1_ADD_99_U131, P1_ADD_99_U132, P1_ADD_99_U133, P1_ADD_99_U134, P1_ADD_99_U135, P1_ADD_99_U136, P1_ADD_99_U137, P1_ADD_99_U138, P1_ADD_99_U139, P1_ADD_99_U14, P1_ADD_99_U140, P1_ADD_99_U141, P1_ADD_99_U142, P1_ADD_99_U143, P1_ADD_99_U144, P1_ADD_99_U145, P1_ADD_99_U146, P1_ADD_99_U147, P1_ADD_99_U148, P1_ADD_99_U149, P1_ADD_99_U15, P1_ADD_99_U150, P1_ADD_99_U151, P1_ADD_99_U152, P1_ADD_99_U153, P1_ADD_99_U16, P1_ADD_99_U17, P1_ADD_99_U18, P1_ADD_99_U19, P1_ADD_99_U20, P1_ADD_99_U21, P1_ADD_99_U22, P1_ADD_99_U23, P1_ADD_99_U24, P1_ADD_99_U25, P1_ADD_99_U26, P1_ADD_99_U27, P1_ADD_99_U28, P1_ADD_99_U29, P1_ADD_99_U30, P1_ADD_99_U31, P1_ADD_99_U32, P1_ADD_99_U33, P1_ADD_99_U34, P1_ADD_99_U35, P1_ADD_99_U36, P1_ADD_99_U37, P1_ADD_99_U38, P1_ADD_99_U39, P1_ADD_99_U4, P1_ADD_99_U40, P1_ADD_99_U41, P1_ADD_99_U42, P1_ADD_99_U43, P1_ADD_99_U44, P1_ADD_99_U45, P1_ADD_99_U46, P1_ADD_99_U47, P1_ADD_99_U48, P1_ADD_99_U49, P1_ADD_99_U5, P1_ADD_99_U50, P1_ADD_99_U51, P1_ADD_99_U52, P1_ADD_99_U53, P1_ADD_99_U54, P1_ADD_99_U55, P1_ADD_99_U56, P1_ADD_99_U57, P1_ADD_99_U58, P1_ADD_99_U59, P1_ADD_99_U6, P1_ADD_99_U60, P1_ADD_99_U61, P1_ADD_99_U62, P1_ADD_99_U63, P1_ADD_99_U64, P1_ADD_99_U65, P1_ADD_99_U66, P1_ADD_99_U67, P1_ADD_99_U68, P1_ADD_99_U69, P1_ADD_99_U7, P1_ADD_99_U70, P1_ADD_99_U71, P1_ADD_99_U72, P1_ADD_99_U73, P1_ADD_99_U74, P1_ADD_99_U75, P1_ADD_99_U76, P1_ADD_99_U77, P1_ADD_99_U78, P1_ADD_99_U79, P1_ADD_99_U8, P1_ADD_99_U80, P1_ADD_99_U81, P1_ADD_99_U82, P1_ADD_99_U83, P1_ADD_99_U84, P1_ADD_99_U85, P1_ADD_99_U86, P1_ADD_99_U87, P1_ADD_99_U88, P1_ADD_99_U89, P1_ADD_99_U9, P1_ADD_99_U90, P1_ADD_99_U91, P1_ADD_99_U92, P1_ADD_99_U93, P1_ADD_99_U94, P1_ADD_99_U95, P1_ADD_99_U96, P1_ADD_99_U97, P1_ADD_99_U98, P1_ADD_99_U99, P1_R1105_U10, P1_R1105_U100, P1_R1105_U101, P1_R1105_U102, P1_R1105_U103, P1_R1105_U104, P1_R1105_U105, P1_R1105_U106, P1_R1105_U107, P1_R1105_U108, P1_R1105_U109, P1_R1105_U11, P1_R1105_U110, P1_R1105_U111, P1_R1105_U112, P1_R1105_U113, P1_R1105_U114, P1_R1105_U115, P1_R1105_U116, P1_R1105_U117, P1_R1105_U118, P1_R1105_U119, P1_R1105_U12, P1_R1105_U120, P1_R1105_U121, P1_R1105_U122, P1_R1105_U123, P1_R1105_U124, P1_R1105_U125, P1_R1105_U126, P1_R1105_U127, P1_R1105_U128, P1_R1105_U129, P1_R1105_U13, P1_R1105_U130, P1_R1105_U131, P1_R1105_U132, P1_R1105_U133, P1_R1105_U134, P1_R1105_U135, P1_R1105_U136, P1_R1105_U137, P1_R1105_U138, P1_R1105_U139, P1_R1105_U14, P1_R1105_U140, P1_R1105_U141, P1_R1105_U142, P1_R1105_U143, P1_R1105_U144, P1_R1105_U145, P1_R1105_U146, P1_R1105_U147, P1_R1105_U148, P1_R1105_U149, P1_R1105_U15, P1_R1105_U150, P1_R1105_U151, P1_R1105_U152, P1_R1105_U153, P1_R1105_U154, P1_R1105_U155, P1_R1105_U156, P1_R1105_U157, P1_R1105_U158, P1_R1105_U159, P1_R1105_U16, P1_R1105_U160, P1_R1105_U161, P1_R1105_U162, P1_R1105_U163, P1_R1105_U164, P1_R1105_U165, P1_R1105_U166, P1_R1105_U167, P1_R1105_U168, P1_R1105_U169, P1_R1105_U17, P1_R1105_U170, P1_R1105_U171, P1_R1105_U172, P1_R1105_U173, P1_R1105_U174, P1_R1105_U175, P1_R1105_U176, P1_R1105_U177, P1_R1105_U178, P1_R1105_U179, P1_R1105_U18, P1_R1105_U180, P1_R1105_U181, P1_R1105_U182, P1_R1105_U183, P1_R1105_U184, P1_R1105_U185, P1_R1105_U186, P1_R1105_U187, P1_R1105_U188, P1_R1105_U189, P1_R1105_U19, P1_R1105_U190, P1_R1105_U191, P1_R1105_U192, P1_R1105_U193, P1_R1105_U194, P1_R1105_U195, P1_R1105_U196, P1_R1105_U197, P1_R1105_U198, P1_R1105_U199, P1_R1105_U20, P1_R1105_U200, P1_R1105_U201, P1_R1105_U202, P1_R1105_U203, P1_R1105_U204, P1_R1105_U205, P1_R1105_U206, P1_R1105_U207, P1_R1105_U208, P1_R1105_U209, P1_R1105_U21, P1_R1105_U210, P1_R1105_U211, P1_R1105_U212, P1_R1105_U213, P1_R1105_U214, P1_R1105_U215, P1_R1105_U216, P1_R1105_U217, P1_R1105_U218, P1_R1105_U219, P1_R1105_U22, P1_R1105_U220, P1_R1105_U221, P1_R1105_U222, P1_R1105_U223, P1_R1105_U224, P1_R1105_U225, P1_R1105_U226, P1_R1105_U227, P1_R1105_U228, P1_R1105_U229, P1_R1105_U23, P1_R1105_U230, P1_R1105_U231, P1_R1105_U232, P1_R1105_U233, P1_R1105_U234, P1_R1105_U235, P1_R1105_U236, P1_R1105_U237, P1_R1105_U238, P1_R1105_U239, P1_R1105_U24, P1_R1105_U240, P1_R1105_U241, P1_R1105_U242, P1_R1105_U243, P1_R1105_U244, P1_R1105_U245, P1_R1105_U246, P1_R1105_U247, P1_R1105_U248, P1_R1105_U249, P1_R1105_U25, P1_R1105_U250, P1_R1105_U251, P1_R1105_U252, P1_R1105_U253, P1_R1105_U254, P1_R1105_U255, P1_R1105_U256, P1_R1105_U257, P1_R1105_U258, P1_R1105_U259, P1_R1105_U26, P1_R1105_U260, P1_R1105_U261, P1_R1105_U262, P1_R1105_U263, P1_R1105_U264, P1_R1105_U265, P1_R1105_U266, P1_R1105_U267, P1_R1105_U268, P1_R1105_U269, P1_R1105_U27, P1_R1105_U270, P1_R1105_U271, P1_R1105_U272, P1_R1105_U273, P1_R1105_U274, P1_R1105_U275, P1_R1105_U276, P1_R1105_U277, P1_R1105_U278, P1_R1105_U279, P1_R1105_U28, P1_R1105_U280, P1_R1105_U281, P1_R1105_U282, P1_R1105_U283, P1_R1105_U284, P1_R1105_U285, P1_R1105_U286, P1_R1105_U287, P1_R1105_U288, P1_R1105_U289, P1_R1105_U29, P1_R1105_U290, P1_R1105_U291, P1_R1105_U292, P1_R1105_U293, P1_R1105_U294, P1_R1105_U295, P1_R1105_U296, P1_R1105_U297, P1_R1105_U298, P1_R1105_U299, P1_R1105_U30, P1_R1105_U300, P1_R1105_U301, P1_R1105_U302, P1_R1105_U303, P1_R1105_U304, P1_R1105_U305, P1_R1105_U306, P1_R1105_U307, P1_R1105_U308, P1_R1105_U31, P1_R1105_U32, P1_R1105_U33, P1_R1105_U34, P1_R1105_U35, P1_R1105_U36, P1_R1105_U37, P1_R1105_U38, P1_R1105_U39, P1_R1105_U4, P1_R1105_U40, P1_R1105_U41, P1_R1105_U42, P1_R1105_U43, P1_R1105_U44, P1_R1105_U45, P1_R1105_U46, P1_R1105_U47, P1_R1105_U48, P1_R1105_U49, P1_R1105_U5, P1_R1105_U50, P1_R1105_U51, P1_R1105_U52, P1_R1105_U53, P1_R1105_U54, P1_R1105_U55, P1_R1105_U56, P1_R1105_U57, P1_R1105_U58, P1_R1105_U59, P1_R1105_U6, P1_R1105_U60, P1_R1105_U61, P1_R1105_U62, P1_R1105_U63, P1_R1105_U64, P1_R1105_U65, P1_R1105_U66, P1_R1105_U67, P1_R1105_U68, P1_R1105_U69, P1_R1105_U7, P1_R1105_U70, P1_R1105_U71, P1_R1105_U72, P1_R1105_U73, P1_R1105_U74, P1_R1105_U75, P1_R1105_U76, P1_R1105_U77, P1_R1105_U78, P1_R1105_U79, P1_R1105_U8, P1_R1105_U80, P1_R1105_U81, P1_R1105_U82, P1_R1105_U83, P1_R1105_U84, P1_R1105_U85, P1_R1105_U86, P1_R1105_U87, P1_R1105_U88, P1_R1105_U89, P1_R1105_U9, P1_R1105_U90, P1_R1105_U91, P1_R1105_U92, P1_R1105_U93, P1_R1105_U94, P1_R1105_U95, P1_R1105_U96, P1_R1105_U97, P1_R1105_U98, P1_R1105_U99, P1_R1117_U10, P1_R1117_U100, P1_R1117_U101, P1_R1117_U102, P1_R1117_U103, P1_R1117_U104, P1_R1117_U105, P1_R1117_U106, P1_R1117_U107, P1_R1117_U108, P1_R1117_U109, P1_R1117_U11, P1_R1117_U110, P1_R1117_U111, P1_R1117_U112, P1_R1117_U113, P1_R1117_U114, P1_R1117_U115, P1_R1117_U116, P1_R1117_U117, P1_R1117_U118, P1_R1117_U119, P1_R1117_U12, P1_R1117_U120, P1_R1117_U121, P1_R1117_U122, P1_R1117_U123, P1_R1117_U124, P1_R1117_U125, P1_R1117_U126, P1_R1117_U127, P1_R1117_U128, P1_R1117_U129, P1_R1117_U13, P1_R1117_U130, P1_R1117_U131, P1_R1117_U132, P1_R1117_U133, P1_R1117_U134, P1_R1117_U135, P1_R1117_U136, P1_R1117_U137, P1_R1117_U138, P1_R1117_U139, P1_R1117_U14, P1_R1117_U140, P1_R1117_U141, P1_R1117_U142, P1_R1117_U143, P1_R1117_U144, P1_R1117_U145, P1_R1117_U146, P1_R1117_U147, P1_R1117_U148, P1_R1117_U149, P1_R1117_U15, P1_R1117_U150, P1_R1117_U151, P1_R1117_U152, P1_R1117_U153, P1_R1117_U154, P1_R1117_U155, P1_R1117_U156, P1_R1117_U157, P1_R1117_U158, P1_R1117_U159, P1_R1117_U16, P1_R1117_U160, P1_R1117_U161, P1_R1117_U162, P1_R1117_U163, P1_R1117_U164, P1_R1117_U165, P1_R1117_U166, P1_R1117_U167, P1_R1117_U168, P1_R1117_U169, P1_R1117_U17, P1_R1117_U170, P1_R1117_U171, P1_R1117_U172, P1_R1117_U173, P1_R1117_U174, P1_R1117_U175, P1_R1117_U176, P1_R1117_U177, P1_R1117_U178, P1_R1117_U179, P1_R1117_U18, P1_R1117_U180, P1_R1117_U181, P1_R1117_U182, P1_R1117_U183, P1_R1117_U184, P1_R1117_U185, P1_R1117_U186, P1_R1117_U187, P1_R1117_U188, P1_R1117_U189, P1_R1117_U19, P1_R1117_U190, P1_R1117_U191, P1_R1117_U192, P1_R1117_U193, P1_R1117_U194, P1_R1117_U195, P1_R1117_U196, P1_R1117_U197, P1_R1117_U198, P1_R1117_U199, P1_R1117_U20, P1_R1117_U200, P1_R1117_U201, P1_R1117_U202, P1_R1117_U203, P1_R1117_U204, P1_R1117_U205, P1_R1117_U206, P1_R1117_U207, P1_R1117_U208, P1_R1117_U209, P1_R1117_U21, P1_R1117_U210, P1_R1117_U211, P1_R1117_U212, P1_R1117_U213, P1_R1117_U214, P1_R1117_U215, P1_R1117_U216, P1_R1117_U217, P1_R1117_U218, P1_R1117_U219, P1_R1117_U22, P1_R1117_U220, P1_R1117_U221, P1_R1117_U222, P1_R1117_U223, P1_R1117_U224, P1_R1117_U225, P1_R1117_U226, P1_R1117_U227, P1_R1117_U228, P1_R1117_U229, P1_R1117_U23, P1_R1117_U230, P1_R1117_U231, P1_R1117_U232, P1_R1117_U233, P1_R1117_U234, P1_R1117_U235, P1_R1117_U236, P1_R1117_U237, P1_R1117_U238, P1_R1117_U239, P1_R1117_U24, P1_R1117_U240, P1_R1117_U241, P1_R1117_U242, P1_R1117_U243, P1_R1117_U244, P1_R1117_U245, P1_R1117_U246, P1_R1117_U247, P1_R1117_U248, P1_R1117_U249, P1_R1117_U25, P1_R1117_U250, P1_R1117_U251, P1_R1117_U252, P1_R1117_U253, P1_R1117_U254, P1_R1117_U255, P1_R1117_U256, P1_R1117_U257, P1_R1117_U258, P1_R1117_U259, P1_R1117_U26, P1_R1117_U260, P1_R1117_U261, P1_R1117_U262, P1_R1117_U263, P1_R1117_U264, P1_R1117_U265, P1_R1117_U266, P1_R1117_U267, P1_R1117_U268, P1_R1117_U269, P1_R1117_U27, P1_R1117_U270, P1_R1117_U271, P1_R1117_U272, P1_R1117_U273, P1_R1117_U274, P1_R1117_U275, P1_R1117_U276, P1_R1117_U277, P1_R1117_U278, P1_R1117_U279, P1_R1117_U28, P1_R1117_U280, P1_R1117_U281, P1_R1117_U282, P1_R1117_U283, P1_R1117_U284, P1_R1117_U285, P1_R1117_U286, P1_R1117_U287, P1_R1117_U288, P1_R1117_U289, P1_R1117_U29, P1_R1117_U290, P1_R1117_U291, P1_R1117_U292, P1_R1117_U293, P1_R1117_U294, P1_R1117_U295, P1_R1117_U296, P1_R1117_U297, P1_R1117_U298, P1_R1117_U299, P1_R1117_U30, P1_R1117_U300, P1_R1117_U301, P1_R1117_U302, P1_R1117_U303, P1_R1117_U304, P1_R1117_U305, P1_R1117_U306, P1_R1117_U307, P1_R1117_U308, P1_R1117_U309, P1_R1117_U31, P1_R1117_U310, P1_R1117_U311, P1_R1117_U312, P1_R1117_U313, P1_R1117_U314, P1_R1117_U315, P1_R1117_U316, P1_R1117_U317, P1_R1117_U318, P1_R1117_U319, P1_R1117_U32, P1_R1117_U320, P1_R1117_U321, P1_R1117_U322, P1_R1117_U323, P1_R1117_U324, P1_R1117_U325, P1_R1117_U326, P1_R1117_U327, P1_R1117_U328, P1_R1117_U329, P1_R1117_U33, P1_R1117_U330, P1_R1117_U331, P1_R1117_U332, P1_R1117_U333, P1_R1117_U334, P1_R1117_U335, P1_R1117_U336, P1_R1117_U337, P1_R1117_U338, P1_R1117_U339, P1_R1117_U34, P1_R1117_U340, P1_R1117_U341, P1_R1117_U342, P1_R1117_U343, P1_R1117_U344, P1_R1117_U345, P1_R1117_U346, P1_R1117_U347, P1_R1117_U348, P1_R1117_U349, P1_R1117_U35, P1_R1117_U350, P1_R1117_U351, P1_R1117_U352, P1_R1117_U353, P1_R1117_U354, P1_R1117_U355, P1_R1117_U356, P1_R1117_U357, P1_R1117_U358, P1_R1117_U359, P1_R1117_U36, P1_R1117_U360, P1_R1117_U361, P1_R1117_U362, P1_R1117_U363, P1_R1117_U364, P1_R1117_U365, P1_R1117_U366, P1_R1117_U367, P1_R1117_U368, P1_R1117_U369, P1_R1117_U37, P1_R1117_U370, P1_R1117_U371, P1_R1117_U372, P1_R1117_U373, P1_R1117_U374, P1_R1117_U375, P1_R1117_U376, P1_R1117_U377, P1_R1117_U378, P1_R1117_U379, P1_R1117_U38, P1_R1117_U380, P1_R1117_U381, P1_R1117_U382, P1_R1117_U383, P1_R1117_U384, P1_R1117_U385, P1_R1117_U386, P1_R1117_U387, P1_R1117_U388, P1_R1117_U389, P1_R1117_U39, P1_R1117_U390, P1_R1117_U391, P1_R1117_U392, P1_R1117_U393, P1_R1117_U394, P1_R1117_U395, P1_R1117_U396, P1_R1117_U397, P1_R1117_U398, P1_R1117_U399, P1_R1117_U40, P1_R1117_U400, P1_R1117_U401, P1_R1117_U402, P1_R1117_U403, P1_R1117_U404, P1_R1117_U405, P1_R1117_U406, P1_R1117_U407, P1_R1117_U408, P1_R1117_U409, P1_R1117_U41, P1_R1117_U410, P1_R1117_U411, P1_R1117_U412, P1_R1117_U413, P1_R1117_U414, P1_R1117_U415, P1_R1117_U416, P1_R1117_U417, P1_R1117_U418, P1_R1117_U419, P1_R1117_U42, P1_R1117_U420, P1_R1117_U421, P1_R1117_U422, P1_R1117_U423, P1_R1117_U424, P1_R1117_U425, P1_R1117_U426, P1_R1117_U427, P1_R1117_U428, P1_R1117_U429, P1_R1117_U43, P1_R1117_U430, P1_R1117_U431, P1_R1117_U432, P1_R1117_U433, P1_R1117_U434, P1_R1117_U435, P1_R1117_U436, P1_R1117_U437, P1_R1117_U438, P1_R1117_U439, P1_R1117_U44, P1_R1117_U440, P1_R1117_U441, P1_R1117_U442, P1_R1117_U443, P1_R1117_U444, P1_R1117_U445, P1_R1117_U446, P1_R1117_U447, P1_R1117_U448, P1_R1117_U449, P1_R1117_U45, P1_R1117_U450, P1_R1117_U451, P1_R1117_U452, P1_R1117_U453, P1_R1117_U454, P1_R1117_U455, P1_R1117_U456, P1_R1117_U457, P1_R1117_U458, P1_R1117_U459, P1_R1117_U46, P1_R1117_U460, P1_R1117_U461, P1_R1117_U462, P1_R1117_U463, P1_R1117_U464, P1_R1117_U465, P1_R1117_U466, P1_R1117_U467, P1_R1117_U468, P1_R1117_U469, P1_R1117_U47, P1_R1117_U470, P1_R1117_U471, P1_R1117_U472, P1_R1117_U473, P1_R1117_U474, P1_R1117_U475, P1_R1117_U476, P1_R1117_U48, P1_R1117_U49, P1_R1117_U50, P1_R1117_U51, P1_R1117_U52, P1_R1117_U53, P1_R1117_U54, P1_R1117_U55, P1_R1117_U56, P1_R1117_U57, P1_R1117_U58, P1_R1117_U59, P1_R1117_U6, P1_R1117_U60, P1_R1117_U61, P1_R1117_U62, P1_R1117_U63, P1_R1117_U64, P1_R1117_U65, P1_R1117_U66, P1_R1117_U67, P1_R1117_U68, P1_R1117_U69, P1_R1117_U7, P1_R1117_U70, P1_R1117_U71, P1_R1117_U72, P1_R1117_U73, P1_R1117_U74, P1_R1117_U75, P1_R1117_U76, P1_R1117_U77, P1_R1117_U78, P1_R1117_U79, P1_R1117_U8, P1_R1117_U80, P1_R1117_U81, P1_R1117_U82, P1_R1117_U83, P1_R1117_U84, P1_R1117_U85, P1_R1117_U86, P1_R1117_U87, P1_R1117_U88, P1_R1117_U89, P1_R1117_U9, P1_R1117_U90, P1_R1117_U91, P1_R1117_U92, P1_R1117_U93, P1_R1117_U94, P1_R1117_U95, P1_R1117_U96, P1_R1117_U97, P1_R1117_U98, P1_R1117_U99, P1_R1138_U10, P1_R1138_U100, P1_R1138_U101, P1_R1138_U102, P1_R1138_U103, P1_R1138_U104, P1_R1138_U105, P1_R1138_U106, P1_R1138_U107, P1_R1138_U108, P1_R1138_U109, P1_R1138_U11, P1_R1138_U110, P1_R1138_U111, P1_R1138_U112, P1_R1138_U113, P1_R1138_U114, P1_R1138_U115, P1_R1138_U116, P1_R1138_U117, P1_R1138_U118, P1_R1138_U119, P1_R1138_U12, P1_R1138_U120, P1_R1138_U121, P1_R1138_U122, P1_R1138_U123, P1_R1138_U124, P1_R1138_U125, P1_R1138_U126, P1_R1138_U127, P1_R1138_U128, P1_R1138_U129, P1_R1138_U13, P1_R1138_U130, P1_R1138_U131, P1_R1138_U132, P1_R1138_U133, P1_R1138_U134, P1_R1138_U135, P1_R1138_U136, P1_R1138_U137, P1_R1138_U138, P1_R1138_U139, P1_R1138_U14, P1_R1138_U140, P1_R1138_U141, P1_R1138_U142, P1_R1138_U143, P1_R1138_U144, P1_R1138_U145, P1_R1138_U146, P1_R1138_U147, P1_R1138_U148, P1_R1138_U149, P1_R1138_U15, P1_R1138_U150, P1_R1138_U151, P1_R1138_U152, P1_R1138_U153, P1_R1138_U154, P1_R1138_U155, P1_R1138_U156, P1_R1138_U157, P1_R1138_U158, P1_R1138_U159, P1_R1138_U16, P1_R1138_U160, P1_R1138_U161, P1_R1138_U162, P1_R1138_U163, P1_R1138_U164, P1_R1138_U165, P1_R1138_U166, P1_R1138_U167, P1_R1138_U168, P1_R1138_U169, P1_R1138_U17, P1_R1138_U170, P1_R1138_U171, P1_R1138_U172, P1_R1138_U173, P1_R1138_U174, P1_R1138_U175, P1_R1138_U176, P1_R1138_U177, P1_R1138_U178, P1_R1138_U179, P1_R1138_U18, P1_R1138_U180, P1_R1138_U181, P1_R1138_U182, P1_R1138_U183, P1_R1138_U184, P1_R1138_U185, P1_R1138_U186, P1_R1138_U187, P1_R1138_U188, P1_R1138_U189, P1_R1138_U19, P1_R1138_U190, P1_R1138_U191, P1_R1138_U192, P1_R1138_U193, P1_R1138_U194, P1_R1138_U195, P1_R1138_U196, P1_R1138_U197, P1_R1138_U198, P1_R1138_U199, P1_R1138_U20, P1_R1138_U200, P1_R1138_U201, P1_R1138_U202, P1_R1138_U203, P1_R1138_U204, P1_R1138_U205, P1_R1138_U206, P1_R1138_U207, P1_R1138_U208, P1_R1138_U209, P1_R1138_U21, P1_R1138_U210, P1_R1138_U211, P1_R1138_U212, P1_R1138_U213, P1_R1138_U214, P1_R1138_U215, P1_R1138_U216, P1_R1138_U217, P1_R1138_U218, P1_R1138_U219, P1_R1138_U22, P1_R1138_U220, P1_R1138_U221, P1_R1138_U222, P1_R1138_U223, P1_R1138_U224, P1_R1138_U225, P1_R1138_U226, P1_R1138_U227, P1_R1138_U228, P1_R1138_U229, P1_R1138_U23, P1_R1138_U230, P1_R1138_U231, P1_R1138_U232, P1_R1138_U233, P1_R1138_U234, P1_R1138_U235, P1_R1138_U236, P1_R1138_U237, P1_R1138_U238, P1_R1138_U239, P1_R1138_U24, P1_R1138_U240, P1_R1138_U241, P1_R1138_U242, P1_R1138_U243, P1_R1138_U244, P1_R1138_U245, P1_R1138_U246, P1_R1138_U247, P1_R1138_U248, P1_R1138_U249, P1_R1138_U25, P1_R1138_U250, P1_R1138_U251, P1_R1138_U252, P1_R1138_U253, P1_R1138_U254, P1_R1138_U255, P1_R1138_U256, P1_R1138_U257, P1_R1138_U258, P1_R1138_U259, P1_R1138_U26, P1_R1138_U260, P1_R1138_U261, P1_R1138_U262, P1_R1138_U263, P1_R1138_U264, P1_R1138_U265, P1_R1138_U266, P1_R1138_U267, P1_R1138_U268, P1_R1138_U269, P1_R1138_U27, P1_R1138_U270, P1_R1138_U271, P1_R1138_U272, P1_R1138_U273, P1_R1138_U274, P1_R1138_U275, P1_R1138_U276, P1_R1138_U277, P1_R1138_U278, P1_R1138_U279, P1_R1138_U28, P1_R1138_U280, P1_R1138_U281, P1_R1138_U282, P1_R1138_U283, P1_R1138_U284, P1_R1138_U285, P1_R1138_U286, P1_R1138_U287, P1_R1138_U288, P1_R1138_U289, P1_R1138_U29, P1_R1138_U290, P1_R1138_U291, P1_R1138_U292, P1_R1138_U293, P1_R1138_U294, P1_R1138_U295, P1_R1138_U296, P1_R1138_U297, P1_R1138_U298, P1_R1138_U299, P1_R1138_U30, P1_R1138_U300, P1_R1138_U301, P1_R1138_U302, P1_R1138_U303, P1_R1138_U304, P1_R1138_U305, P1_R1138_U306, P1_R1138_U307, P1_R1138_U308, P1_R1138_U309, P1_R1138_U31, P1_R1138_U310, P1_R1138_U311, P1_R1138_U312, P1_R1138_U313, P1_R1138_U314, P1_R1138_U315, P1_R1138_U316, P1_R1138_U317, P1_R1138_U318, P1_R1138_U319, P1_R1138_U32, P1_R1138_U320, P1_R1138_U321, P1_R1138_U322, P1_R1138_U323, P1_R1138_U324, P1_R1138_U325, P1_R1138_U326, P1_R1138_U327, P1_R1138_U328, P1_R1138_U329, P1_R1138_U33, P1_R1138_U330, P1_R1138_U331, P1_R1138_U332, P1_R1138_U333, P1_R1138_U334, P1_R1138_U335, P1_R1138_U336, P1_R1138_U337, P1_R1138_U338, P1_R1138_U339, P1_R1138_U34, P1_R1138_U340, P1_R1138_U341, P1_R1138_U342, P1_R1138_U343, P1_R1138_U344, P1_R1138_U345, P1_R1138_U346, P1_R1138_U347, P1_R1138_U348, P1_R1138_U349, P1_R1138_U35, P1_R1138_U350, P1_R1138_U351, P1_R1138_U352, P1_R1138_U353, P1_R1138_U354, P1_R1138_U355, P1_R1138_U356, P1_R1138_U357, P1_R1138_U358, P1_R1138_U359, P1_R1138_U36, P1_R1138_U360, P1_R1138_U361, P1_R1138_U362, P1_R1138_U363, P1_R1138_U364, P1_R1138_U365, P1_R1138_U366, P1_R1138_U367, P1_R1138_U368, P1_R1138_U369, P1_R1138_U37, P1_R1138_U370, P1_R1138_U371, P1_R1138_U372, P1_R1138_U373, P1_R1138_U374, P1_R1138_U375, P1_R1138_U376, P1_R1138_U377, P1_R1138_U378, P1_R1138_U379, P1_R1138_U38, P1_R1138_U380, P1_R1138_U381, P1_R1138_U382, P1_R1138_U383, P1_R1138_U384, P1_R1138_U385, P1_R1138_U386, P1_R1138_U387, P1_R1138_U388, P1_R1138_U389, P1_R1138_U39, P1_R1138_U390, P1_R1138_U391, P1_R1138_U392, P1_R1138_U393, P1_R1138_U394, P1_R1138_U395, P1_R1138_U396, P1_R1138_U397, P1_R1138_U398, P1_R1138_U399, P1_R1138_U4, P1_R1138_U40, P1_R1138_U400, P1_R1138_U401, P1_R1138_U402, P1_R1138_U403, P1_R1138_U404, P1_R1138_U405, P1_R1138_U406, P1_R1138_U407, P1_R1138_U408, P1_R1138_U409, P1_R1138_U41, P1_R1138_U410, P1_R1138_U411, P1_R1138_U412, P1_R1138_U413, P1_R1138_U414, P1_R1138_U415, P1_R1138_U416, P1_R1138_U417, P1_R1138_U418, P1_R1138_U419, P1_R1138_U42, P1_R1138_U420, P1_R1138_U421, P1_R1138_U422, P1_R1138_U423, P1_R1138_U424, P1_R1138_U425, P1_R1138_U426, P1_R1138_U427, P1_R1138_U428, P1_R1138_U429, P1_R1138_U43, P1_R1138_U430, P1_R1138_U431, P1_R1138_U432, P1_R1138_U433, P1_R1138_U434, P1_R1138_U435, P1_R1138_U436, P1_R1138_U437, P1_R1138_U438, P1_R1138_U439, P1_R1138_U44, P1_R1138_U440, P1_R1138_U441, P1_R1138_U442, P1_R1138_U443, P1_R1138_U444, P1_R1138_U445, P1_R1138_U446, P1_R1138_U447, P1_R1138_U448, P1_R1138_U449, P1_R1138_U45, P1_R1138_U450, P1_R1138_U451, P1_R1138_U452, P1_R1138_U453, P1_R1138_U454, P1_R1138_U455, P1_R1138_U456, P1_R1138_U457, P1_R1138_U458, P1_R1138_U459, P1_R1138_U46, P1_R1138_U460, P1_R1138_U461, P1_R1138_U462, P1_R1138_U463, P1_R1138_U464, P1_R1138_U465, P1_R1138_U466, P1_R1138_U467, P1_R1138_U468, P1_R1138_U469, P1_R1138_U47, P1_R1138_U470, P1_R1138_U471, P1_R1138_U472, P1_R1138_U473, P1_R1138_U474, P1_R1138_U475, P1_R1138_U476, P1_R1138_U477, P1_R1138_U478, P1_R1138_U479, P1_R1138_U48, P1_R1138_U480, P1_R1138_U481, P1_R1138_U482, P1_R1138_U483, P1_R1138_U484, P1_R1138_U485, P1_R1138_U486, P1_R1138_U487, P1_R1138_U488, P1_R1138_U489, P1_R1138_U49, P1_R1138_U490, P1_R1138_U491, P1_R1138_U492, P1_R1138_U493, P1_R1138_U494, P1_R1138_U495, P1_R1138_U496, P1_R1138_U497, P1_R1138_U498, P1_R1138_U499, P1_R1138_U5, P1_R1138_U50, P1_R1138_U500, P1_R1138_U501, P1_R1138_U51, P1_R1138_U52, P1_R1138_U53, P1_R1138_U54, P1_R1138_U55, P1_R1138_U56, P1_R1138_U57, P1_R1138_U58, P1_R1138_U59, P1_R1138_U6, P1_R1138_U60, P1_R1138_U61, P1_R1138_U62, P1_R1138_U63, P1_R1138_U64, P1_R1138_U65, P1_R1138_U66, P1_R1138_U67, P1_R1138_U68, P1_R1138_U69, P1_R1138_U7, P1_R1138_U70, P1_R1138_U71, P1_R1138_U72, P1_R1138_U73, P1_R1138_U74, P1_R1138_U75, P1_R1138_U76, P1_R1138_U77, P1_R1138_U78, P1_R1138_U79, P1_R1138_U8, P1_R1138_U80, P1_R1138_U81, P1_R1138_U82, P1_R1138_U83, P1_R1138_U84, P1_R1138_U85, P1_R1138_U86, P1_R1138_U87, P1_R1138_U88, P1_R1138_U89, P1_R1138_U9, P1_R1138_U90, P1_R1138_U91, P1_R1138_U92, P1_R1138_U93, P1_R1138_U94, P1_R1138_U95, P1_R1138_U96, P1_R1138_U97, P1_R1138_U98, P1_R1138_U99, P1_R1150_U10, P1_R1150_U100, P1_R1150_U101, P1_R1150_U102, P1_R1150_U103, P1_R1150_U104, P1_R1150_U105, P1_R1150_U106, P1_R1150_U107, P1_R1150_U108, P1_R1150_U109, P1_R1150_U11, P1_R1150_U110, P1_R1150_U111, P1_R1150_U112, P1_R1150_U113, P1_R1150_U114, P1_R1150_U115, P1_R1150_U116, P1_R1150_U117, P1_R1150_U118, P1_R1150_U119, P1_R1150_U12, P1_R1150_U120, P1_R1150_U121, P1_R1150_U122, P1_R1150_U123, P1_R1150_U124, P1_R1150_U125, P1_R1150_U126, P1_R1150_U127, P1_R1150_U128, P1_R1150_U129, P1_R1150_U13, P1_R1150_U130, P1_R1150_U131, P1_R1150_U132, P1_R1150_U133, P1_R1150_U134, P1_R1150_U135, P1_R1150_U136, P1_R1150_U137, P1_R1150_U138, P1_R1150_U139, P1_R1150_U14, P1_R1150_U140, P1_R1150_U141, P1_R1150_U142, P1_R1150_U143, P1_R1150_U144, P1_R1150_U145, P1_R1150_U146, P1_R1150_U147, P1_R1150_U148, P1_R1150_U149, P1_R1150_U15, P1_R1150_U150, P1_R1150_U151, P1_R1150_U152, P1_R1150_U153, P1_R1150_U154, P1_R1150_U155, P1_R1150_U156, P1_R1150_U157, P1_R1150_U158, P1_R1150_U159, P1_R1150_U16, P1_R1150_U160, P1_R1150_U161, P1_R1150_U162, P1_R1150_U163, P1_R1150_U164, P1_R1150_U165, P1_R1150_U166, P1_R1150_U167, P1_R1150_U168, P1_R1150_U169, P1_R1150_U17, P1_R1150_U170, P1_R1150_U171, P1_R1150_U172, P1_R1150_U173, P1_R1150_U174, P1_R1150_U175, P1_R1150_U176, P1_R1150_U177, P1_R1150_U178, P1_R1150_U179, P1_R1150_U18, P1_R1150_U180, P1_R1150_U181, P1_R1150_U182, P1_R1150_U183, P1_R1150_U184, P1_R1150_U185, P1_R1150_U186, P1_R1150_U187, P1_R1150_U188, P1_R1150_U189, P1_R1150_U19, P1_R1150_U190, P1_R1150_U191, P1_R1150_U192, P1_R1150_U193, P1_R1150_U194, P1_R1150_U195, P1_R1150_U196, P1_R1150_U197, P1_R1150_U198, P1_R1150_U199, P1_R1150_U20, P1_R1150_U200, P1_R1150_U201, P1_R1150_U202, P1_R1150_U203, P1_R1150_U204, P1_R1150_U205, P1_R1150_U206, P1_R1150_U207, P1_R1150_U208, P1_R1150_U209, P1_R1150_U21, P1_R1150_U210, P1_R1150_U211, P1_R1150_U212, P1_R1150_U213, P1_R1150_U214, P1_R1150_U215, P1_R1150_U216, P1_R1150_U217, P1_R1150_U218, P1_R1150_U219, P1_R1150_U22, P1_R1150_U220, P1_R1150_U221, P1_R1150_U222, P1_R1150_U223, P1_R1150_U224, P1_R1150_U225, P1_R1150_U226, P1_R1150_U227, P1_R1150_U228, P1_R1150_U229, P1_R1150_U23, P1_R1150_U230, P1_R1150_U231, P1_R1150_U232, P1_R1150_U233, P1_R1150_U234, P1_R1150_U235, P1_R1150_U236, P1_R1150_U237, P1_R1150_U238, P1_R1150_U239, P1_R1150_U24, P1_R1150_U240, P1_R1150_U241, P1_R1150_U242, P1_R1150_U243, P1_R1150_U244, P1_R1150_U245, P1_R1150_U246, P1_R1150_U247, P1_R1150_U248, P1_R1150_U249, P1_R1150_U25, P1_R1150_U250, P1_R1150_U251, P1_R1150_U252, P1_R1150_U253, P1_R1150_U254, P1_R1150_U255, P1_R1150_U256, P1_R1150_U257, P1_R1150_U258, P1_R1150_U259, P1_R1150_U26, P1_R1150_U260, P1_R1150_U261, P1_R1150_U262, P1_R1150_U263, P1_R1150_U264, P1_R1150_U265, P1_R1150_U266, P1_R1150_U267, P1_R1150_U268, P1_R1150_U269, P1_R1150_U27, P1_R1150_U270, P1_R1150_U271, P1_R1150_U272, P1_R1150_U273, P1_R1150_U274, P1_R1150_U275, P1_R1150_U276, P1_R1150_U277, P1_R1150_U278, P1_R1150_U279, P1_R1150_U28, P1_R1150_U280, P1_R1150_U281, P1_R1150_U282, P1_R1150_U283, P1_R1150_U284, P1_R1150_U285, P1_R1150_U286, P1_R1150_U287, P1_R1150_U288, P1_R1150_U289, P1_R1150_U29, P1_R1150_U290, P1_R1150_U291, P1_R1150_U292, P1_R1150_U293, P1_R1150_U294, P1_R1150_U295, P1_R1150_U296, P1_R1150_U297, P1_R1150_U298, P1_R1150_U299, P1_R1150_U30, P1_R1150_U300, P1_R1150_U301, P1_R1150_U302, P1_R1150_U303, P1_R1150_U304, P1_R1150_U305, P1_R1150_U306, P1_R1150_U307, P1_R1150_U308, P1_R1150_U309, P1_R1150_U31, P1_R1150_U310, P1_R1150_U311, P1_R1150_U312, P1_R1150_U313, P1_R1150_U314, P1_R1150_U315, P1_R1150_U316, P1_R1150_U317, P1_R1150_U318, P1_R1150_U319, P1_R1150_U32, P1_R1150_U320, P1_R1150_U321, P1_R1150_U322, P1_R1150_U323, P1_R1150_U324, P1_R1150_U325, P1_R1150_U326, P1_R1150_U327, P1_R1150_U328, P1_R1150_U329, P1_R1150_U33, P1_R1150_U330, P1_R1150_U331, P1_R1150_U332, P1_R1150_U333, P1_R1150_U334, P1_R1150_U335, P1_R1150_U336, P1_R1150_U337, P1_R1150_U338, P1_R1150_U339, P1_R1150_U34, P1_R1150_U340, P1_R1150_U341, P1_R1150_U342, P1_R1150_U343, P1_R1150_U344, P1_R1150_U345, P1_R1150_U346, P1_R1150_U347, P1_R1150_U348, P1_R1150_U349, P1_R1150_U35, P1_R1150_U350, P1_R1150_U351, P1_R1150_U352, P1_R1150_U353, P1_R1150_U354, P1_R1150_U355, P1_R1150_U356, P1_R1150_U357, P1_R1150_U358, P1_R1150_U359, P1_R1150_U36, P1_R1150_U360, P1_R1150_U361, P1_R1150_U362, P1_R1150_U363, P1_R1150_U364, P1_R1150_U365, P1_R1150_U366, P1_R1150_U367, P1_R1150_U368, P1_R1150_U369, P1_R1150_U37, P1_R1150_U370, P1_R1150_U371, P1_R1150_U372, P1_R1150_U373, P1_R1150_U374, P1_R1150_U375, P1_R1150_U376, P1_R1150_U377, P1_R1150_U378, P1_R1150_U379, P1_R1150_U38, P1_R1150_U380, P1_R1150_U381, P1_R1150_U382, P1_R1150_U383, P1_R1150_U384, P1_R1150_U385, P1_R1150_U386, P1_R1150_U387, P1_R1150_U388, P1_R1150_U389, P1_R1150_U39, P1_R1150_U390, P1_R1150_U391, P1_R1150_U392, P1_R1150_U393, P1_R1150_U394, P1_R1150_U395, P1_R1150_U396, P1_R1150_U397, P1_R1150_U398, P1_R1150_U399, P1_R1150_U40, P1_R1150_U400, P1_R1150_U401, P1_R1150_U402, P1_R1150_U403, P1_R1150_U404, P1_R1150_U405, P1_R1150_U406, P1_R1150_U407, P1_R1150_U408, P1_R1150_U409, P1_R1150_U41, P1_R1150_U410, P1_R1150_U411, P1_R1150_U412, P1_R1150_U413, P1_R1150_U414, P1_R1150_U415, P1_R1150_U416, P1_R1150_U417, P1_R1150_U418, P1_R1150_U419, P1_R1150_U42, P1_R1150_U420, P1_R1150_U421, P1_R1150_U422, P1_R1150_U423, P1_R1150_U424, P1_R1150_U425, P1_R1150_U426, P1_R1150_U427, P1_R1150_U428, P1_R1150_U429, P1_R1150_U43, P1_R1150_U430, P1_R1150_U431, P1_R1150_U432, P1_R1150_U433, P1_R1150_U434, P1_R1150_U435, P1_R1150_U436, P1_R1150_U437, P1_R1150_U438, P1_R1150_U439, P1_R1150_U44, P1_R1150_U440, P1_R1150_U441, P1_R1150_U442, P1_R1150_U443, P1_R1150_U444, P1_R1150_U445, P1_R1150_U446, P1_R1150_U447, P1_R1150_U448, P1_R1150_U449, P1_R1150_U45, P1_R1150_U450, P1_R1150_U451, P1_R1150_U452, P1_R1150_U453, P1_R1150_U454, P1_R1150_U455, P1_R1150_U456, P1_R1150_U457, P1_R1150_U458, P1_R1150_U459, P1_R1150_U46, P1_R1150_U460, P1_R1150_U461, P1_R1150_U462, P1_R1150_U463, P1_R1150_U464, P1_R1150_U465, P1_R1150_U466, P1_R1150_U467, P1_R1150_U468, P1_R1150_U469, P1_R1150_U47, P1_R1150_U470, P1_R1150_U471, P1_R1150_U472, P1_R1150_U473, P1_R1150_U474, P1_R1150_U475, P1_R1150_U476, P1_R1150_U48, P1_R1150_U49, P1_R1150_U50, P1_R1150_U51, P1_R1150_U52, P1_R1150_U53, P1_R1150_U54, P1_R1150_U55, P1_R1150_U56, P1_R1150_U57, P1_R1150_U58, P1_R1150_U59, P1_R1150_U6, P1_R1150_U60, P1_R1150_U61, P1_R1150_U62, P1_R1150_U63, P1_R1150_U64, P1_R1150_U65, P1_R1150_U66, P1_R1150_U67, P1_R1150_U68, P1_R1150_U69, P1_R1150_U7, P1_R1150_U70, P1_R1150_U71, P1_R1150_U72, P1_R1150_U73, P1_R1150_U74, P1_R1150_U75, P1_R1150_U76, P1_R1150_U77, P1_R1150_U78, P1_R1150_U79, P1_R1150_U8, P1_R1150_U80, P1_R1150_U81, P1_R1150_U82, P1_R1150_U83, P1_R1150_U84, P1_R1150_U85, P1_R1150_U86, P1_R1150_U87, P1_R1150_U88, P1_R1150_U89, P1_R1150_U9, P1_R1150_U90, P1_R1150_U91, P1_R1150_U92, P1_R1150_U93, P1_R1150_U94, P1_R1150_U95, P1_R1150_U96, P1_R1150_U97, P1_R1150_U98, P1_R1150_U99, P1_R1162_U10, P1_R1162_U100, P1_R1162_U101, P1_R1162_U102, P1_R1162_U103, P1_R1162_U104, P1_R1162_U105, P1_R1162_U106, P1_R1162_U107, P1_R1162_U108, P1_R1162_U109, P1_R1162_U11, P1_R1162_U110, P1_R1162_U111, P1_R1162_U112, P1_R1162_U113, P1_R1162_U114, P1_R1162_U115, P1_R1162_U116, P1_R1162_U117, P1_R1162_U118, P1_R1162_U119, P1_R1162_U12, P1_R1162_U120, P1_R1162_U121, P1_R1162_U122, P1_R1162_U123, P1_R1162_U124, P1_R1162_U125, P1_R1162_U126, P1_R1162_U127, P1_R1162_U128, P1_R1162_U129, P1_R1162_U13, P1_R1162_U130, P1_R1162_U131, P1_R1162_U132, P1_R1162_U133, P1_R1162_U134, P1_R1162_U135, P1_R1162_U136, P1_R1162_U137, P1_R1162_U138, P1_R1162_U139, P1_R1162_U14, P1_R1162_U140, P1_R1162_U141, P1_R1162_U142, P1_R1162_U143, P1_R1162_U144, P1_R1162_U145, P1_R1162_U146, P1_R1162_U147, P1_R1162_U148, P1_R1162_U149, P1_R1162_U15, P1_R1162_U150, P1_R1162_U151, P1_R1162_U152, P1_R1162_U153, P1_R1162_U154, P1_R1162_U155, P1_R1162_U156, P1_R1162_U157, P1_R1162_U158, P1_R1162_U159, P1_R1162_U16, P1_R1162_U160, P1_R1162_U161, P1_R1162_U162, P1_R1162_U163, P1_R1162_U164, P1_R1162_U165, P1_R1162_U166, P1_R1162_U167, P1_R1162_U168, P1_R1162_U169, P1_R1162_U17, P1_R1162_U170, P1_R1162_U171, P1_R1162_U172, P1_R1162_U173, P1_R1162_U174, P1_R1162_U175, P1_R1162_U176, P1_R1162_U177, P1_R1162_U178, P1_R1162_U179, P1_R1162_U18, P1_R1162_U180, P1_R1162_U181, P1_R1162_U182, P1_R1162_U183, P1_R1162_U184, P1_R1162_U185, P1_R1162_U186, P1_R1162_U187, P1_R1162_U188, P1_R1162_U189, P1_R1162_U19, P1_R1162_U190, P1_R1162_U191, P1_R1162_U192, P1_R1162_U193, P1_R1162_U194, P1_R1162_U195, P1_R1162_U196, P1_R1162_U197, P1_R1162_U198, P1_R1162_U199, P1_R1162_U20, P1_R1162_U200, P1_R1162_U201, P1_R1162_U202, P1_R1162_U203, P1_R1162_U204, P1_R1162_U205, P1_R1162_U206, P1_R1162_U207, P1_R1162_U208, P1_R1162_U209, P1_R1162_U21, P1_R1162_U210, P1_R1162_U211, P1_R1162_U212, P1_R1162_U213, P1_R1162_U214, P1_R1162_U215, P1_R1162_U216, P1_R1162_U217, P1_R1162_U218, P1_R1162_U219, P1_R1162_U22, P1_R1162_U220, P1_R1162_U221, P1_R1162_U222, P1_R1162_U223, P1_R1162_U224, P1_R1162_U225, P1_R1162_U226, P1_R1162_U227, P1_R1162_U228, P1_R1162_U229, P1_R1162_U23, P1_R1162_U230, P1_R1162_U231, P1_R1162_U232, P1_R1162_U233, P1_R1162_U234, P1_R1162_U235, P1_R1162_U236, P1_R1162_U237, P1_R1162_U238, P1_R1162_U239, P1_R1162_U24, P1_R1162_U240, P1_R1162_U241, P1_R1162_U242, P1_R1162_U243, P1_R1162_U244, P1_R1162_U245, P1_R1162_U246, P1_R1162_U247, P1_R1162_U248, P1_R1162_U249, P1_R1162_U25, P1_R1162_U250, P1_R1162_U251, P1_R1162_U252, P1_R1162_U253, P1_R1162_U254, P1_R1162_U255, P1_R1162_U256, P1_R1162_U257, P1_R1162_U258, P1_R1162_U259, P1_R1162_U26, P1_R1162_U260, P1_R1162_U261, P1_R1162_U262, P1_R1162_U263, P1_R1162_U264, P1_R1162_U265, P1_R1162_U266, P1_R1162_U267, P1_R1162_U268, P1_R1162_U269, P1_R1162_U27, P1_R1162_U270, P1_R1162_U271, P1_R1162_U272, P1_R1162_U273, P1_R1162_U274, P1_R1162_U275, P1_R1162_U276, P1_R1162_U277, P1_R1162_U278, P1_R1162_U279, P1_R1162_U28, P1_R1162_U280, P1_R1162_U281, P1_R1162_U282, P1_R1162_U283, P1_R1162_U284, P1_R1162_U285, P1_R1162_U286, P1_R1162_U287, P1_R1162_U288, P1_R1162_U289, P1_R1162_U29, P1_R1162_U290, P1_R1162_U291, P1_R1162_U292, P1_R1162_U293, P1_R1162_U294, P1_R1162_U295, P1_R1162_U296, P1_R1162_U297, P1_R1162_U298, P1_R1162_U299, P1_R1162_U30, P1_R1162_U300, P1_R1162_U301, P1_R1162_U302, P1_R1162_U303, P1_R1162_U304, P1_R1162_U305, P1_R1162_U306, P1_R1162_U307, P1_R1162_U308, P1_R1162_U31, P1_R1162_U32, P1_R1162_U33, P1_R1162_U34, P1_R1162_U35, P1_R1162_U36, P1_R1162_U37, P1_R1162_U38, P1_R1162_U39, P1_R1162_U4, P1_R1162_U40, P1_R1162_U41, P1_R1162_U42, P1_R1162_U43, P1_R1162_U44, P1_R1162_U45, P1_R1162_U46, P1_R1162_U47, P1_R1162_U48, P1_R1162_U49, P1_R1162_U5, P1_R1162_U50, P1_R1162_U51, P1_R1162_U52, P1_R1162_U53, P1_R1162_U54, P1_R1162_U55, P1_R1162_U56, P1_R1162_U57, P1_R1162_U58, P1_R1162_U59, P1_R1162_U6, P1_R1162_U60, P1_R1162_U61, P1_R1162_U62, P1_R1162_U63, P1_R1162_U64, P1_R1162_U65, P1_R1162_U66, P1_R1162_U67, P1_R1162_U68, P1_R1162_U69, P1_R1162_U7, P1_R1162_U70, P1_R1162_U71, P1_R1162_U72, P1_R1162_U73, P1_R1162_U74, P1_R1162_U75, P1_R1162_U76, P1_R1162_U77, P1_R1162_U78, P1_R1162_U79, P1_R1162_U8, P1_R1162_U80, P1_R1162_U81, P1_R1162_U82, P1_R1162_U83, P1_R1162_U84, P1_R1162_U85, P1_R1162_U86, P1_R1162_U87, P1_R1162_U88, P1_R1162_U89, P1_R1162_U9, P1_R1162_U90, P1_R1162_U91, P1_R1162_U92, P1_R1162_U93, P1_R1162_U94, P1_R1162_U95, P1_R1162_U96, P1_R1162_U97, P1_R1162_U98, P1_R1162_U99, P1_R1165_U10, P1_R1165_U100, P1_R1165_U101, P1_R1165_U102, P1_R1165_U103, P1_R1165_U104, P1_R1165_U105, P1_R1165_U106, P1_R1165_U107, P1_R1165_U108, P1_R1165_U109, P1_R1165_U11, P1_R1165_U110, P1_R1165_U111, P1_R1165_U112, P1_R1165_U113, P1_R1165_U114, P1_R1165_U115, P1_R1165_U116, P1_R1165_U117, P1_R1165_U118, P1_R1165_U119, P1_R1165_U12, P1_R1165_U120, P1_R1165_U121, P1_R1165_U122, P1_R1165_U123, P1_R1165_U124, P1_R1165_U125, P1_R1165_U126, P1_R1165_U127, P1_R1165_U128, P1_R1165_U129, P1_R1165_U13, P1_R1165_U130, P1_R1165_U131, P1_R1165_U132, P1_R1165_U133, P1_R1165_U134, P1_R1165_U135, P1_R1165_U136, P1_R1165_U137, P1_R1165_U138, P1_R1165_U139, P1_R1165_U14, P1_R1165_U140, P1_R1165_U141, P1_R1165_U142, P1_R1165_U143, P1_R1165_U144, P1_R1165_U145, P1_R1165_U146, P1_R1165_U147, P1_R1165_U148, P1_R1165_U149, P1_R1165_U15, P1_R1165_U150, P1_R1165_U151, P1_R1165_U152, P1_R1165_U153, P1_R1165_U154, P1_R1165_U155, P1_R1165_U156, P1_R1165_U157, P1_R1165_U158, P1_R1165_U159, P1_R1165_U16, P1_R1165_U160, P1_R1165_U161, P1_R1165_U162, P1_R1165_U163, P1_R1165_U164, P1_R1165_U165, P1_R1165_U166, P1_R1165_U167, P1_R1165_U168, P1_R1165_U169, P1_R1165_U17, P1_R1165_U170, P1_R1165_U171, P1_R1165_U172, P1_R1165_U173, P1_R1165_U174, P1_R1165_U175, P1_R1165_U176, P1_R1165_U177, P1_R1165_U178, P1_R1165_U179, P1_R1165_U18, P1_R1165_U180, P1_R1165_U181, P1_R1165_U182, P1_R1165_U183, P1_R1165_U184, P1_R1165_U185, P1_R1165_U186, P1_R1165_U187, P1_R1165_U188, P1_R1165_U189, P1_R1165_U19, P1_R1165_U190, P1_R1165_U191, P1_R1165_U192, P1_R1165_U193, P1_R1165_U194, P1_R1165_U195, P1_R1165_U196, P1_R1165_U197, P1_R1165_U198, P1_R1165_U199, P1_R1165_U20, P1_R1165_U200, P1_R1165_U201, P1_R1165_U202, P1_R1165_U203, P1_R1165_U204, P1_R1165_U205, P1_R1165_U206, P1_R1165_U207, P1_R1165_U208, P1_R1165_U209, P1_R1165_U21, P1_R1165_U210, P1_R1165_U211, P1_R1165_U212, P1_R1165_U213, P1_R1165_U214, P1_R1165_U215, P1_R1165_U216, P1_R1165_U217, P1_R1165_U218, P1_R1165_U219, P1_R1165_U22, P1_R1165_U220, P1_R1165_U221, P1_R1165_U222, P1_R1165_U223, P1_R1165_U224, P1_R1165_U225, P1_R1165_U226, P1_R1165_U227, P1_R1165_U228, P1_R1165_U229, P1_R1165_U23, P1_R1165_U230, P1_R1165_U231, P1_R1165_U232, P1_R1165_U233, P1_R1165_U234, P1_R1165_U235, P1_R1165_U236, P1_R1165_U237, P1_R1165_U238, P1_R1165_U239, P1_R1165_U24, P1_R1165_U240, P1_R1165_U241, P1_R1165_U242, P1_R1165_U243, P1_R1165_U244, P1_R1165_U245, P1_R1165_U246, P1_R1165_U247, P1_R1165_U248, P1_R1165_U249, P1_R1165_U25, P1_R1165_U250, P1_R1165_U251, P1_R1165_U252, P1_R1165_U253, P1_R1165_U254, P1_R1165_U255, P1_R1165_U256, P1_R1165_U257, P1_R1165_U258, P1_R1165_U259, P1_R1165_U26, P1_R1165_U260, P1_R1165_U261, P1_R1165_U262, P1_R1165_U263, P1_R1165_U264, P1_R1165_U265, P1_R1165_U266, P1_R1165_U267, P1_R1165_U268, P1_R1165_U269, P1_R1165_U27, P1_R1165_U270, P1_R1165_U271, P1_R1165_U272, P1_R1165_U273, P1_R1165_U274, P1_R1165_U275, P1_R1165_U276, P1_R1165_U277, P1_R1165_U278, P1_R1165_U279, P1_R1165_U28, P1_R1165_U280, P1_R1165_U281, P1_R1165_U282, P1_R1165_U283, P1_R1165_U284, P1_R1165_U285, P1_R1165_U286, P1_R1165_U287, P1_R1165_U288, P1_R1165_U289, P1_R1165_U29, P1_R1165_U290, P1_R1165_U291, P1_R1165_U292, P1_R1165_U293, P1_R1165_U294, P1_R1165_U295, P1_R1165_U296, P1_R1165_U297, P1_R1165_U298, P1_R1165_U299, P1_R1165_U30, P1_R1165_U300, P1_R1165_U301, P1_R1165_U302, P1_R1165_U303, P1_R1165_U304, P1_R1165_U305, P1_R1165_U306, P1_R1165_U307, P1_R1165_U308, P1_R1165_U309, P1_R1165_U31, P1_R1165_U310, P1_R1165_U311, P1_R1165_U312, P1_R1165_U313, P1_R1165_U314, P1_R1165_U315, P1_R1165_U316, P1_R1165_U317, P1_R1165_U318, P1_R1165_U319, P1_R1165_U32, P1_R1165_U320, P1_R1165_U321, P1_R1165_U322, P1_R1165_U323, P1_R1165_U324, P1_R1165_U325, P1_R1165_U326, P1_R1165_U327, P1_R1165_U328, P1_R1165_U329, P1_R1165_U33, P1_R1165_U330, P1_R1165_U331, P1_R1165_U332, P1_R1165_U333, P1_R1165_U334, P1_R1165_U335, P1_R1165_U336, P1_R1165_U337, P1_R1165_U338, P1_R1165_U339, P1_R1165_U34, P1_R1165_U340, P1_R1165_U341, P1_R1165_U342, P1_R1165_U343, P1_R1165_U344, P1_R1165_U345, P1_R1165_U346, P1_R1165_U347, P1_R1165_U348, P1_R1165_U349, P1_R1165_U35, P1_R1165_U350, P1_R1165_U351, P1_R1165_U352, P1_R1165_U353, P1_R1165_U354, P1_R1165_U355, P1_R1165_U356, P1_R1165_U357, P1_R1165_U358, P1_R1165_U359, P1_R1165_U36, P1_R1165_U360, P1_R1165_U361, P1_R1165_U362, P1_R1165_U363, P1_R1165_U364, P1_R1165_U365, P1_R1165_U366, P1_R1165_U367, P1_R1165_U368, P1_R1165_U369, P1_R1165_U37, P1_R1165_U370, P1_R1165_U371, P1_R1165_U372, P1_R1165_U373, P1_R1165_U374, P1_R1165_U375, P1_R1165_U376, P1_R1165_U377, P1_R1165_U378, P1_R1165_U379, P1_R1165_U38, P1_R1165_U380, P1_R1165_U381, P1_R1165_U382, P1_R1165_U383, P1_R1165_U384, P1_R1165_U385, P1_R1165_U386, P1_R1165_U387, P1_R1165_U388, P1_R1165_U389, P1_R1165_U39, P1_R1165_U390, P1_R1165_U391, P1_R1165_U392, P1_R1165_U393, P1_R1165_U394, P1_R1165_U395, P1_R1165_U396, P1_R1165_U397, P1_R1165_U398, P1_R1165_U399, P1_R1165_U4, P1_R1165_U40, P1_R1165_U400, P1_R1165_U401, P1_R1165_U402, P1_R1165_U403, P1_R1165_U404, P1_R1165_U405, P1_R1165_U406, P1_R1165_U407, P1_R1165_U408, P1_R1165_U409, P1_R1165_U41, P1_R1165_U410, P1_R1165_U411, P1_R1165_U412, P1_R1165_U413, P1_R1165_U414, P1_R1165_U415, P1_R1165_U416, P1_R1165_U417, P1_R1165_U418, P1_R1165_U419, P1_R1165_U42, P1_R1165_U420, P1_R1165_U421, P1_R1165_U422, P1_R1165_U423, P1_R1165_U424, P1_R1165_U425, P1_R1165_U426, P1_R1165_U427, P1_R1165_U428, P1_R1165_U429, P1_R1165_U43, P1_R1165_U430, P1_R1165_U431, P1_R1165_U432, P1_R1165_U433, P1_R1165_U434, P1_R1165_U435, P1_R1165_U436, P1_R1165_U437, P1_R1165_U438, P1_R1165_U439, P1_R1165_U44, P1_R1165_U440, P1_R1165_U441, P1_R1165_U442, P1_R1165_U443, P1_R1165_U444, P1_R1165_U445, P1_R1165_U446, P1_R1165_U447, P1_R1165_U448, P1_R1165_U449, P1_R1165_U45, P1_R1165_U450, P1_R1165_U451, P1_R1165_U452, P1_R1165_U453, P1_R1165_U454, P1_R1165_U455, P1_R1165_U456, P1_R1165_U457, P1_R1165_U458, P1_R1165_U459, P1_R1165_U46, P1_R1165_U460, P1_R1165_U461, P1_R1165_U462, P1_R1165_U463, P1_R1165_U464, P1_R1165_U465, P1_R1165_U466, P1_R1165_U467, P1_R1165_U468, P1_R1165_U469, P1_R1165_U47, P1_R1165_U470, P1_R1165_U471, P1_R1165_U472, P1_R1165_U473, P1_R1165_U474, P1_R1165_U475, P1_R1165_U476, P1_R1165_U477, P1_R1165_U478, P1_R1165_U479, P1_R1165_U48, P1_R1165_U480, P1_R1165_U481, P1_R1165_U482, P1_R1165_U483, P1_R1165_U484, P1_R1165_U485, P1_R1165_U486, P1_R1165_U487, P1_R1165_U488, P1_R1165_U489, P1_R1165_U49, P1_R1165_U490, P1_R1165_U491, P1_R1165_U492, P1_R1165_U493, P1_R1165_U494, P1_R1165_U495, P1_R1165_U496, P1_R1165_U497, P1_R1165_U498, P1_R1165_U499, P1_R1165_U5, P1_R1165_U50, P1_R1165_U500, P1_R1165_U501, P1_R1165_U502, P1_R1165_U503, P1_R1165_U504, P1_R1165_U505, P1_R1165_U506, P1_R1165_U507, P1_R1165_U508, P1_R1165_U509, P1_R1165_U51, P1_R1165_U510, P1_R1165_U511, P1_R1165_U512, P1_R1165_U513, P1_R1165_U514, P1_R1165_U515, P1_R1165_U516, P1_R1165_U517, P1_R1165_U518, P1_R1165_U519, P1_R1165_U52, P1_R1165_U520, P1_R1165_U521, P1_R1165_U522, P1_R1165_U523, P1_R1165_U524, P1_R1165_U525, P1_R1165_U526, P1_R1165_U527, P1_R1165_U528, P1_R1165_U529, P1_R1165_U53, P1_R1165_U530, P1_R1165_U531, P1_R1165_U532, P1_R1165_U533, P1_R1165_U534, P1_R1165_U535, P1_R1165_U536, P1_R1165_U537, P1_R1165_U538, P1_R1165_U539, P1_R1165_U54, P1_R1165_U540, P1_R1165_U541, P1_R1165_U542, P1_R1165_U543, P1_R1165_U544, P1_R1165_U545, P1_R1165_U546, P1_R1165_U547, P1_R1165_U548, P1_R1165_U549, P1_R1165_U55, P1_R1165_U550, P1_R1165_U551, P1_R1165_U552, P1_R1165_U553, P1_R1165_U554, P1_R1165_U555, P1_R1165_U556, P1_R1165_U557, P1_R1165_U558, P1_R1165_U559, P1_R1165_U56, P1_R1165_U560, P1_R1165_U561, P1_R1165_U562, P1_R1165_U563, P1_R1165_U564, P1_R1165_U565, P1_R1165_U566, P1_R1165_U567, P1_R1165_U568, P1_R1165_U569, P1_R1165_U57, P1_R1165_U570, P1_R1165_U571, P1_R1165_U572, P1_R1165_U573, P1_R1165_U574, P1_R1165_U575, P1_R1165_U576, P1_R1165_U577, P1_R1165_U578, P1_R1165_U579, P1_R1165_U58, P1_R1165_U580, P1_R1165_U581, P1_R1165_U582, P1_R1165_U583, P1_R1165_U584, P1_R1165_U585, P1_R1165_U586, P1_R1165_U587, P1_R1165_U588, P1_R1165_U589, P1_R1165_U59, P1_R1165_U590, P1_R1165_U591, P1_R1165_U592, P1_R1165_U593, P1_R1165_U594, P1_R1165_U595, P1_R1165_U6, P1_R1165_U60, P1_R1165_U61, P1_R1165_U62, P1_R1165_U63, P1_R1165_U64, P1_R1165_U65, P1_R1165_U66, P1_R1165_U67, P1_R1165_U68, P1_R1165_U69, P1_R1165_U7, P1_R1165_U70, P1_R1165_U71, P1_R1165_U72, P1_R1165_U73, P1_R1165_U74, P1_R1165_U75, P1_R1165_U76, P1_R1165_U77, P1_R1165_U78, P1_R1165_U79, P1_R1165_U8, P1_R1165_U80, P1_R1165_U81, P1_R1165_U82, P1_R1165_U83, P1_R1165_U84, P1_R1165_U85, P1_R1165_U86, P1_R1165_U87, P1_R1165_U88, P1_R1165_U89, P1_R1165_U9, P1_R1165_U90, P1_R1165_U91, P1_R1165_U92, P1_R1165_U93, P1_R1165_U94, P1_R1165_U95, P1_R1165_U96, P1_R1165_U97, P1_R1165_U98, P1_R1165_U99, P1_R1171_U10, P1_R1171_U100, P1_R1171_U101, P1_R1171_U102, P1_R1171_U103, P1_R1171_U104, P1_R1171_U105, P1_R1171_U106, P1_R1171_U107, P1_R1171_U108, P1_R1171_U109, P1_R1171_U11, P1_R1171_U110, P1_R1171_U111, P1_R1171_U112, P1_R1171_U113, P1_R1171_U114, P1_R1171_U115, P1_R1171_U116, P1_R1171_U117, P1_R1171_U118, P1_R1171_U119, P1_R1171_U12, P1_R1171_U120, P1_R1171_U121, P1_R1171_U122, P1_R1171_U123, P1_R1171_U124, P1_R1171_U125, P1_R1171_U126, P1_R1171_U127, P1_R1171_U128, P1_R1171_U129, P1_R1171_U13, P1_R1171_U130, P1_R1171_U131, P1_R1171_U132, P1_R1171_U133, P1_R1171_U134, P1_R1171_U135, P1_R1171_U136, P1_R1171_U137, P1_R1171_U138, P1_R1171_U139, P1_R1171_U14, P1_R1171_U140, P1_R1171_U141, P1_R1171_U142, P1_R1171_U143, P1_R1171_U144, P1_R1171_U145, P1_R1171_U146, P1_R1171_U147, P1_R1171_U148, P1_R1171_U149, P1_R1171_U15, P1_R1171_U150, P1_R1171_U151, P1_R1171_U152, P1_R1171_U153, P1_R1171_U154, P1_R1171_U155, P1_R1171_U156, P1_R1171_U157, P1_R1171_U158, P1_R1171_U159, P1_R1171_U16, P1_R1171_U160, P1_R1171_U161, P1_R1171_U162, P1_R1171_U163, P1_R1171_U164, P1_R1171_U165, P1_R1171_U166, P1_R1171_U167, P1_R1171_U168, P1_R1171_U169, P1_R1171_U17, P1_R1171_U170, P1_R1171_U171, P1_R1171_U172, P1_R1171_U173, P1_R1171_U174, P1_R1171_U175, P1_R1171_U176, P1_R1171_U177, P1_R1171_U178, P1_R1171_U179, P1_R1171_U18, P1_R1171_U180, P1_R1171_U181, P1_R1171_U182, P1_R1171_U183, P1_R1171_U184, P1_R1171_U185, P1_R1171_U186, P1_R1171_U187, P1_R1171_U188, P1_R1171_U189, P1_R1171_U19, P1_R1171_U190, P1_R1171_U191, P1_R1171_U192, P1_R1171_U193, P1_R1171_U194, P1_R1171_U195, P1_R1171_U196, P1_R1171_U197, P1_R1171_U198, P1_R1171_U199, P1_R1171_U20, P1_R1171_U200, P1_R1171_U201, P1_R1171_U202, P1_R1171_U203, P1_R1171_U204, P1_R1171_U205, P1_R1171_U206, P1_R1171_U207, P1_R1171_U208, P1_R1171_U209, P1_R1171_U21, P1_R1171_U210, P1_R1171_U211, P1_R1171_U212, P1_R1171_U213, P1_R1171_U214, P1_R1171_U215, P1_R1171_U216, P1_R1171_U217, P1_R1171_U218, P1_R1171_U219, P1_R1171_U22, P1_R1171_U220, P1_R1171_U221, P1_R1171_U222, P1_R1171_U223, P1_R1171_U224, P1_R1171_U225, P1_R1171_U226, P1_R1171_U227, P1_R1171_U228, P1_R1171_U229, P1_R1171_U23, P1_R1171_U230, P1_R1171_U231, P1_R1171_U232, P1_R1171_U233, P1_R1171_U234, P1_R1171_U235, P1_R1171_U236, P1_R1171_U237, P1_R1171_U238, P1_R1171_U239, P1_R1171_U24, P1_R1171_U240, P1_R1171_U241, P1_R1171_U242, P1_R1171_U243, P1_R1171_U244, P1_R1171_U245, P1_R1171_U246, P1_R1171_U247, P1_R1171_U248, P1_R1171_U249, P1_R1171_U25, P1_R1171_U250, P1_R1171_U251, P1_R1171_U252, P1_R1171_U253, P1_R1171_U254, P1_R1171_U255, P1_R1171_U256, P1_R1171_U257, P1_R1171_U258, P1_R1171_U259, P1_R1171_U26, P1_R1171_U260, P1_R1171_U261, P1_R1171_U262, P1_R1171_U263, P1_R1171_U264, P1_R1171_U265, P1_R1171_U266, P1_R1171_U267, P1_R1171_U268, P1_R1171_U269, P1_R1171_U27, P1_R1171_U270, P1_R1171_U271, P1_R1171_U272, P1_R1171_U273, P1_R1171_U274, P1_R1171_U275, P1_R1171_U276, P1_R1171_U277, P1_R1171_U278, P1_R1171_U279, P1_R1171_U28, P1_R1171_U280, P1_R1171_U281, P1_R1171_U282, P1_R1171_U283, P1_R1171_U284, P1_R1171_U285, P1_R1171_U286, P1_R1171_U287, P1_R1171_U288, P1_R1171_U289, P1_R1171_U29, P1_R1171_U290, P1_R1171_U291, P1_R1171_U292, P1_R1171_U293, P1_R1171_U294, P1_R1171_U295, P1_R1171_U296, P1_R1171_U297, P1_R1171_U298, P1_R1171_U299, P1_R1171_U30, P1_R1171_U300, P1_R1171_U301, P1_R1171_U302, P1_R1171_U303, P1_R1171_U304, P1_R1171_U305, P1_R1171_U306, P1_R1171_U307, P1_R1171_U308, P1_R1171_U309, P1_R1171_U31, P1_R1171_U310, P1_R1171_U311, P1_R1171_U312, P1_R1171_U313, P1_R1171_U314, P1_R1171_U315, P1_R1171_U316, P1_R1171_U317, P1_R1171_U318, P1_R1171_U319, P1_R1171_U32, P1_R1171_U320, P1_R1171_U321, P1_R1171_U322, P1_R1171_U323, P1_R1171_U324, P1_R1171_U325, P1_R1171_U326, P1_R1171_U327, P1_R1171_U328, P1_R1171_U329, P1_R1171_U33, P1_R1171_U330, P1_R1171_U331, P1_R1171_U332, P1_R1171_U333, P1_R1171_U334, P1_R1171_U335, P1_R1171_U336, P1_R1171_U337, P1_R1171_U338, P1_R1171_U339, P1_R1171_U34, P1_R1171_U340, P1_R1171_U341, P1_R1171_U342, P1_R1171_U343, P1_R1171_U344, P1_R1171_U345, P1_R1171_U346, P1_R1171_U347, P1_R1171_U348, P1_R1171_U349, P1_R1171_U35, P1_R1171_U350, P1_R1171_U351, P1_R1171_U352, P1_R1171_U353, P1_R1171_U354, P1_R1171_U355, P1_R1171_U356, P1_R1171_U357, P1_R1171_U358, P1_R1171_U359, P1_R1171_U36, P1_R1171_U360, P1_R1171_U361, P1_R1171_U362, P1_R1171_U363, P1_R1171_U364, P1_R1171_U365, P1_R1171_U366, P1_R1171_U367, P1_R1171_U368, P1_R1171_U369, P1_R1171_U37, P1_R1171_U370, P1_R1171_U371, P1_R1171_U372, P1_R1171_U373, P1_R1171_U374, P1_R1171_U375, P1_R1171_U376, P1_R1171_U377, P1_R1171_U378, P1_R1171_U379, P1_R1171_U38, P1_R1171_U380, P1_R1171_U381, P1_R1171_U382, P1_R1171_U383, P1_R1171_U384, P1_R1171_U385, P1_R1171_U386, P1_R1171_U387, P1_R1171_U388, P1_R1171_U389, P1_R1171_U39, P1_R1171_U390, P1_R1171_U391, P1_R1171_U392, P1_R1171_U393, P1_R1171_U394, P1_R1171_U395, P1_R1171_U396, P1_R1171_U397, P1_R1171_U398, P1_R1171_U399, P1_R1171_U4, P1_R1171_U40, P1_R1171_U400, P1_R1171_U401, P1_R1171_U402, P1_R1171_U403, P1_R1171_U404, P1_R1171_U405, P1_R1171_U406, P1_R1171_U407, P1_R1171_U408, P1_R1171_U409, P1_R1171_U41, P1_R1171_U410, P1_R1171_U411, P1_R1171_U412, P1_R1171_U413, P1_R1171_U414, P1_R1171_U415, P1_R1171_U416, P1_R1171_U417, P1_R1171_U418, P1_R1171_U419, P1_R1171_U42, P1_R1171_U420, P1_R1171_U421, P1_R1171_U422, P1_R1171_U423, P1_R1171_U424, P1_R1171_U425, P1_R1171_U426, P1_R1171_U427, P1_R1171_U428, P1_R1171_U429, P1_R1171_U43, P1_R1171_U430, P1_R1171_U431, P1_R1171_U432, P1_R1171_U433, P1_R1171_U434, P1_R1171_U435, P1_R1171_U436, P1_R1171_U437, P1_R1171_U438, P1_R1171_U439, P1_R1171_U44, P1_R1171_U440, P1_R1171_U441, P1_R1171_U442, P1_R1171_U443, P1_R1171_U444, P1_R1171_U445, P1_R1171_U446, P1_R1171_U447, P1_R1171_U448, P1_R1171_U449, P1_R1171_U45, P1_R1171_U450, P1_R1171_U451, P1_R1171_U452, P1_R1171_U453, P1_R1171_U454, P1_R1171_U455, P1_R1171_U456, P1_R1171_U457, P1_R1171_U458, P1_R1171_U459, P1_R1171_U46, P1_R1171_U460, P1_R1171_U461, P1_R1171_U462, P1_R1171_U463, P1_R1171_U464, P1_R1171_U465, P1_R1171_U466, P1_R1171_U467, P1_R1171_U468, P1_R1171_U469, P1_R1171_U47, P1_R1171_U470, P1_R1171_U471, P1_R1171_U472, P1_R1171_U473, P1_R1171_U474, P1_R1171_U475, P1_R1171_U476, P1_R1171_U477, P1_R1171_U478, P1_R1171_U479, P1_R1171_U48, P1_R1171_U480, P1_R1171_U481, P1_R1171_U482, P1_R1171_U483, P1_R1171_U484, P1_R1171_U485, P1_R1171_U486, P1_R1171_U487, P1_R1171_U488, P1_R1171_U489, P1_R1171_U49, P1_R1171_U490, P1_R1171_U491, P1_R1171_U492, P1_R1171_U493, P1_R1171_U494, P1_R1171_U495, P1_R1171_U496, P1_R1171_U497, P1_R1171_U498, P1_R1171_U499, P1_R1171_U5, P1_R1171_U50, P1_R1171_U500, P1_R1171_U501, P1_R1171_U51, P1_R1171_U52, P1_R1171_U53, P1_R1171_U54, P1_R1171_U55, P1_R1171_U56, P1_R1171_U57, P1_R1171_U58, P1_R1171_U59, P1_R1171_U6, P1_R1171_U60, P1_R1171_U61, P1_R1171_U62, P1_R1171_U63, P1_R1171_U64, P1_R1171_U65, P1_R1171_U66, P1_R1171_U67, P1_R1171_U68, P1_R1171_U69, P1_R1171_U7, P1_R1171_U70, P1_R1171_U71, P1_R1171_U72, P1_R1171_U73, P1_R1171_U74, P1_R1171_U75, P1_R1171_U76, P1_R1171_U77, P1_R1171_U78, P1_R1171_U79, P1_R1171_U8, P1_R1171_U80, P1_R1171_U81, P1_R1171_U82, P1_R1171_U83, P1_R1171_U84, P1_R1171_U85, P1_R1171_U86, P1_R1171_U87, P1_R1171_U88, P1_R1171_U89, P1_R1171_U9, P1_R1171_U90, P1_R1171_U91, P1_R1171_U92, P1_R1171_U93, P1_R1171_U94, P1_R1171_U95, P1_R1171_U96, P1_R1171_U97, P1_R1171_U98, P1_R1171_U99, P1_R1192_U10, P1_R1192_U100, P1_R1192_U101, P1_R1192_U102, P1_R1192_U103, P1_R1192_U104, P1_R1192_U105, P1_R1192_U106, P1_R1192_U107, P1_R1192_U108, P1_R1192_U109, P1_R1192_U11, P1_R1192_U110, P1_R1192_U111, P1_R1192_U112, P1_R1192_U113, P1_R1192_U114, P1_R1192_U115, P1_R1192_U116, P1_R1192_U117, P1_R1192_U118, P1_R1192_U119, P1_R1192_U12, P1_R1192_U120, P1_R1192_U121, P1_R1192_U122, P1_R1192_U123, P1_R1192_U124, P1_R1192_U125, P1_R1192_U126, P1_R1192_U127, P1_R1192_U128, P1_R1192_U129, P1_R1192_U13, P1_R1192_U130, P1_R1192_U131, P1_R1192_U132, P1_R1192_U133, P1_R1192_U134, P1_R1192_U135, P1_R1192_U136, P1_R1192_U137, P1_R1192_U138, P1_R1192_U139, P1_R1192_U14, P1_R1192_U140, P1_R1192_U141, P1_R1192_U142, P1_R1192_U143, P1_R1192_U144, P1_R1192_U145, P1_R1192_U146, P1_R1192_U147, P1_R1192_U148, P1_R1192_U149, P1_R1192_U15, P1_R1192_U150, P1_R1192_U151, P1_R1192_U152, P1_R1192_U153, P1_R1192_U154, P1_R1192_U155, P1_R1192_U156, P1_R1192_U157, P1_R1192_U158, P1_R1192_U159, P1_R1192_U16, P1_R1192_U160, P1_R1192_U161, P1_R1192_U162, P1_R1192_U163, P1_R1192_U164, P1_R1192_U165, P1_R1192_U166, P1_R1192_U167, P1_R1192_U168, P1_R1192_U169, P1_R1192_U17, P1_R1192_U170, P1_R1192_U171, P1_R1192_U172, P1_R1192_U173, P1_R1192_U174, P1_R1192_U175, P1_R1192_U176, P1_R1192_U177, P1_R1192_U178, P1_R1192_U179, P1_R1192_U18, P1_R1192_U180, P1_R1192_U181, P1_R1192_U182, P1_R1192_U183, P1_R1192_U184, P1_R1192_U185, P1_R1192_U186, P1_R1192_U187, P1_R1192_U188, P1_R1192_U189, P1_R1192_U19, P1_R1192_U190, P1_R1192_U191, P1_R1192_U192, P1_R1192_U193, P1_R1192_U194, P1_R1192_U195, P1_R1192_U196, P1_R1192_U197, P1_R1192_U198, P1_R1192_U199, P1_R1192_U20, P1_R1192_U200, P1_R1192_U201, P1_R1192_U202, P1_R1192_U203, P1_R1192_U204, P1_R1192_U205, P1_R1192_U206, P1_R1192_U207, P1_R1192_U208, P1_R1192_U209, P1_R1192_U21, P1_R1192_U210, P1_R1192_U211, P1_R1192_U212, P1_R1192_U213, P1_R1192_U214, P1_R1192_U215, P1_R1192_U216, P1_R1192_U217, P1_R1192_U218, P1_R1192_U219, P1_R1192_U22, P1_R1192_U220, P1_R1192_U221, P1_R1192_U222, P1_R1192_U223, P1_R1192_U224, P1_R1192_U225, P1_R1192_U226, P1_R1192_U227, P1_R1192_U228, P1_R1192_U229, P1_R1192_U23, P1_R1192_U230, P1_R1192_U231, P1_R1192_U232, P1_R1192_U233, P1_R1192_U234, P1_R1192_U235, P1_R1192_U236, P1_R1192_U237, P1_R1192_U238, P1_R1192_U239, P1_R1192_U24, P1_R1192_U240, P1_R1192_U241, P1_R1192_U242, P1_R1192_U243, P1_R1192_U244, P1_R1192_U245, P1_R1192_U246, P1_R1192_U247, P1_R1192_U248, P1_R1192_U249, P1_R1192_U25, P1_R1192_U250, P1_R1192_U251, P1_R1192_U252, P1_R1192_U253, P1_R1192_U254, P1_R1192_U255, P1_R1192_U256, P1_R1192_U257, P1_R1192_U258, P1_R1192_U259, P1_R1192_U26, P1_R1192_U260, P1_R1192_U261, P1_R1192_U262, P1_R1192_U263, P1_R1192_U264, P1_R1192_U265, P1_R1192_U266, P1_R1192_U267, P1_R1192_U268, P1_R1192_U269, P1_R1192_U27, P1_R1192_U270, P1_R1192_U271, P1_R1192_U272, P1_R1192_U273, P1_R1192_U274, P1_R1192_U275, P1_R1192_U276, P1_R1192_U277, P1_R1192_U278, P1_R1192_U279, P1_R1192_U28, P1_R1192_U280, P1_R1192_U281, P1_R1192_U282, P1_R1192_U283, P1_R1192_U284, P1_R1192_U285, P1_R1192_U286, P1_R1192_U287, P1_R1192_U288, P1_R1192_U289, P1_R1192_U29, P1_R1192_U290, P1_R1192_U291, P1_R1192_U292, P1_R1192_U293, P1_R1192_U294, P1_R1192_U295, P1_R1192_U296, P1_R1192_U297, P1_R1192_U298, P1_R1192_U299, P1_R1192_U30, P1_R1192_U300, P1_R1192_U301, P1_R1192_U302, P1_R1192_U303, P1_R1192_U304, P1_R1192_U305, P1_R1192_U306, P1_R1192_U307, P1_R1192_U308, P1_R1192_U309, P1_R1192_U31, P1_R1192_U310, P1_R1192_U311, P1_R1192_U312, P1_R1192_U313, P1_R1192_U314, P1_R1192_U315, P1_R1192_U316, P1_R1192_U317, P1_R1192_U318, P1_R1192_U319, P1_R1192_U32, P1_R1192_U320, P1_R1192_U321, P1_R1192_U322, P1_R1192_U323, P1_R1192_U324, P1_R1192_U325, P1_R1192_U326, P1_R1192_U327, P1_R1192_U328, P1_R1192_U329, P1_R1192_U33, P1_R1192_U330, P1_R1192_U331, P1_R1192_U332, P1_R1192_U333, P1_R1192_U334, P1_R1192_U335, P1_R1192_U336, P1_R1192_U337, P1_R1192_U338, P1_R1192_U339, P1_R1192_U34, P1_R1192_U340, P1_R1192_U341, P1_R1192_U342, P1_R1192_U343, P1_R1192_U344, P1_R1192_U345, P1_R1192_U346, P1_R1192_U347, P1_R1192_U348, P1_R1192_U349, P1_R1192_U35, P1_R1192_U350, P1_R1192_U351, P1_R1192_U352, P1_R1192_U353, P1_R1192_U354, P1_R1192_U355, P1_R1192_U356, P1_R1192_U357, P1_R1192_U358, P1_R1192_U359, P1_R1192_U36, P1_R1192_U360, P1_R1192_U361, P1_R1192_U362, P1_R1192_U363, P1_R1192_U364, P1_R1192_U365, P1_R1192_U366, P1_R1192_U367, P1_R1192_U368, P1_R1192_U369, P1_R1192_U37, P1_R1192_U370, P1_R1192_U371, P1_R1192_U372, P1_R1192_U373, P1_R1192_U374, P1_R1192_U375, P1_R1192_U376, P1_R1192_U377, P1_R1192_U378, P1_R1192_U379, P1_R1192_U38, P1_R1192_U380, P1_R1192_U381, P1_R1192_U382, P1_R1192_U383, P1_R1192_U384, P1_R1192_U385, P1_R1192_U386, P1_R1192_U387, P1_R1192_U388, P1_R1192_U389, P1_R1192_U39, P1_R1192_U390, P1_R1192_U391, P1_R1192_U392, P1_R1192_U393, P1_R1192_U394, P1_R1192_U395, P1_R1192_U396, P1_R1192_U397, P1_R1192_U398, P1_R1192_U399, P1_R1192_U40, P1_R1192_U400, P1_R1192_U401, P1_R1192_U402, P1_R1192_U403, P1_R1192_U404, P1_R1192_U405, P1_R1192_U406, P1_R1192_U407, P1_R1192_U408, P1_R1192_U409, P1_R1192_U41, P1_R1192_U410, P1_R1192_U411, P1_R1192_U412, P1_R1192_U413, P1_R1192_U414, P1_R1192_U415, P1_R1192_U416, P1_R1192_U417, P1_R1192_U418, P1_R1192_U419, P1_R1192_U42, P1_R1192_U420, P1_R1192_U421, P1_R1192_U422, P1_R1192_U423, P1_R1192_U424, P1_R1192_U425, P1_R1192_U426, P1_R1192_U427, P1_R1192_U428, P1_R1192_U429, P1_R1192_U43, P1_R1192_U430, P1_R1192_U431, P1_R1192_U432, P1_R1192_U433, P1_R1192_U434, P1_R1192_U435, P1_R1192_U436, P1_R1192_U437, P1_R1192_U438, P1_R1192_U439, P1_R1192_U44, P1_R1192_U440, P1_R1192_U441, P1_R1192_U442, P1_R1192_U443, P1_R1192_U444, P1_R1192_U445, P1_R1192_U446, P1_R1192_U447, P1_R1192_U448, P1_R1192_U449, P1_R1192_U45, P1_R1192_U450, P1_R1192_U451, P1_R1192_U452, P1_R1192_U453, P1_R1192_U454, P1_R1192_U455, P1_R1192_U456, P1_R1192_U457, P1_R1192_U458, P1_R1192_U459, P1_R1192_U46, P1_R1192_U460, P1_R1192_U461, P1_R1192_U462, P1_R1192_U463, P1_R1192_U464, P1_R1192_U465, P1_R1192_U466, P1_R1192_U467, P1_R1192_U468, P1_R1192_U469, P1_R1192_U47, P1_R1192_U470, P1_R1192_U471, P1_R1192_U472, P1_R1192_U473, P1_R1192_U474, P1_R1192_U475, P1_R1192_U476, P1_R1192_U48, P1_R1192_U49, P1_R1192_U50, P1_R1192_U51, P1_R1192_U52, P1_R1192_U53, P1_R1192_U54, P1_R1192_U55, P1_R1192_U56, P1_R1192_U57, P1_R1192_U58, P1_R1192_U59, P1_R1192_U6, P1_R1192_U60, P1_R1192_U61, P1_R1192_U62, P1_R1192_U63, P1_R1192_U64, P1_R1192_U65, P1_R1192_U66, P1_R1192_U67, P1_R1192_U68, P1_R1192_U69, P1_R1192_U7, P1_R1192_U70, P1_R1192_U71, P1_R1192_U72, P1_R1192_U73, P1_R1192_U74, P1_R1192_U75, P1_R1192_U76, P1_R1192_U77, P1_R1192_U78, P1_R1192_U79, P1_R1192_U8, P1_R1192_U80, P1_R1192_U81, P1_R1192_U82, P1_R1192_U83, P1_R1192_U84, P1_R1192_U85, P1_R1192_U86, P1_R1192_U87, P1_R1192_U88, P1_R1192_U89, P1_R1192_U9, P1_R1192_U90, P1_R1192_U91, P1_R1192_U92, P1_R1192_U93, P1_R1192_U94, P1_R1192_U95, P1_R1192_U96, P1_R1192_U97, P1_R1192_U98, P1_R1192_U99, P1_R1207_U10, P1_R1207_U100, P1_R1207_U101, P1_R1207_U102, P1_R1207_U103, P1_R1207_U104, P1_R1207_U105, P1_R1207_U106, P1_R1207_U107, P1_R1207_U108, P1_R1207_U109, P1_R1207_U11, P1_R1207_U110, P1_R1207_U111, P1_R1207_U112, P1_R1207_U113, P1_R1207_U114, P1_R1207_U115, P1_R1207_U116, P1_R1207_U117, P1_R1207_U118, P1_R1207_U119, P1_R1207_U12, P1_R1207_U120, P1_R1207_U121, P1_R1207_U122, P1_R1207_U123, P1_R1207_U124, P1_R1207_U125, P1_R1207_U126, P1_R1207_U127, P1_R1207_U128, P1_R1207_U129, P1_R1207_U13, P1_R1207_U130, P1_R1207_U131, P1_R1207_U132, P1_R1207_U133, P1_R1207_U134, P1_R1207_U135, P1_R1207_U136, P1_R1207_U137, P1_R1207_U138, P1_R1207_U139, P1_R1207_U14, P1_R1207_U140, P1_R1207_U141, P1_R1207_U142, P1_R1207_U143, P1_R1207_U144, P1_R1207_U145, P1_R1207_U146, P1_R1207_U147, P1_R1207_U148, P1_R1207_U149, P1_R1207_U15, P1_R1207_U150, P1_R1207_U151, P1_R1207_U152, P1_R1207_U153, P1_R1207_U154, P1_R1207_U155, P1_R1207_U156, P1_R1207_U157, P1_R1207_U158, P1_R1207_U159, P1_R1207_U16, P1_R1207_U160, P1_R1207_U161, P1_R1207_U162, P1_R1207_U163, P1_R1207_U164, P1_R1207_U165, P1_R1207_U166, P1_R1207_U167, P1_R1207_U168, P1_R1207_U169, P1_R1207_U17, P1_R1207_U170, P1_R1207_U171, P1_R1207_U172, P1_R1207_U173, P1_R1207_U174, P1_R1207_U175, P1_R1207_U176, P1_R1207_U177, P1_R1207_U178, P1_R1207_U179, P1_R1207_U18, P1_R1207_U180, P1_R1207_U181, P1_R1207_U182, P1_R1207_U183, P1_R1207_U184, P1_R1207_U185, P1_R1207_U186, P1_R1207_U187, P1_R1207_U188, P1_R1207_U189, P1_R1207_U19, P1_R1207_U190, P1_R1207_U191, P1_R1207_U192, P1_R1207_U193, P1_R1207_U194, P1_R1207_U195, P1_R1207_U196, P1_R1207_U197, P1_R1207_U198, P1_R1207_U199, P1_R1207_U20, P1_R1207_U200, P1_R1207_U201, P1_R1207_U202, P1_R1207_U203, P1_R1207_U204, P1_R1207_U205, P1_R1207_U206, P1_R1207_U207, P1_R1207_U208, P1_R1207_U209, P1_R1207_U21, P1_R1207_U210, P1_R1207_U211, P1_R1207_U212, P1_R1207_U213, P1_R1207_U214, P1_R1207_U215, P1_R1207_U216, P1_R1207_U217, P1_R1207_U218, P1_R1207_U219, P1_R1207_U22, P1_R1207_U220, P1_R1207_U221, P1_R1207_U222, P1_R1207_U223, P1_R1207_U224, P1_R1207_U225, P1_R1207_U226, P1_R1207_U227, P1_R1207_U228, P1_R1207_U229, P1_R1207_U23, P1_R1207_U230, P1_R1207_U231, P1_R1207_U232, P1_R1207_U233, P1_R1207_U234, P1_R1207_U235, P1_R1207_U236, P1_R1207_U237, P1_R1207_U238, P1_R1207_U239, P1_R1207_U24, P1_R1207_U240, P1_R1207_U241, P1_R1207_U242, P1_R1207_U243, P1_R1207_U244, P1_R1207_U245, P1_R1207_U246, P1_R1207_U247, P1_R1207_U248, P1_R1207_U249, P1_R1207_U25, P1_R1207_U250, P1_R1207_U251, P1_R1207_U252, P1_R1207_U253, P1_R1207_U254, P1_R1207_U255, P1_R1207_U256, P1_R1207_U257, P1_R1207_U258, P1_R1207_U259, P1_R1207_U26, P1_R1207_U260, P1_R1207_U261, P1_R1207_U262, P1_R1207_U263, P1_R1207_U264, P1_R1207_U265, P1_R1207_U266, P1_R1207_U267, P1_R1207_U268, P1_R1207_U269, P1_R1207_U27, P1_R1207_U270, P1_R1207_U271, P1_R1207_U272, P1_R1207_U273, P1_R1207_U274, P1_R1207_U275, P1_R1207_U276, P1_R1207_U277, P1_R1207_U278, P1_R1207_U279, P1_R1207_U28, P1_R1207_U280, P1_R1207_U281, P1_R1207_U282, P1_R1207_U283, P1_R1207_U284, P1_R1207_U285, P1_R1207_U286, P1_R1207_U287, P1_R1207_U288, P1_R1207_U289, P1_R1207_U29, P1_R1207_U290, P1_R1207_U291, P1_R1207_U292, P1_R1207_U293, P1_R1207_U294, P1_R1207_U295, P1_R1207_U296, P1_R1207_U297, P1_R1207_U298, P1_R1207_U299, P1_R1207_U30, P1_R1207_U300, P1_R1207_U301, P1_R1207_U302, P1_R1207_U303, P1_R1207_U304, P1_R1207_U305, P1_R1207_U306, P1_R1207_U307, P1_R1207_U308, P1_R1207_U309, P1_R1207_U31, P1_R1207_U310, P1_R1207_U311, P1_R1207_U312, P1_R1207_U313, P1_R1207_U314, P1_R1207_U315, P1_R1207_U316, P1_R1207_U317, P1_R1207_U318, P1_R1207_U319, P1_R1207_U32, P1_R1207_U320, P1_R1207_U321, P1_R1207_U322, P1_R1207_U323, P1_R1207_U324, P1_R1207_U325, P1_R1207_U326, P1_R1207_U327, P1_R1207_U328, P1_R1207_U329, P1_R1207_U33, P1_R1207_U330, P1_R1207_U331, P1_R1207_U332, P1_R1207_U333, P1_R1207_U334, P1_R1207_U335, P1_R1207_U336, P1_R1207_U337, P1_R1207_U338, P1_R1207_U339, P1_R1207_U34, P1_R1207_U340, P1_R1207_U341, P1_R1207_U342, P1_R1207_U343, P1_R1207_U344, P1_R1207_U345, P1_R1207_U346, P1_R1207_U347, P1_R1207_U348, P1_R1207_U349, P1_R1207_U35, P1_R1207_U350, P1_R1207_U351, P1_R1207_U352, P1_R1207_U353, P1_R1207_U354, P1_R1207_U355, P1_R1207_U356, P1_R1207_U357, P1_R1207_U358, P1_R1207_U359, P1_R1207_U36, P1_R1207_U360, P1_R1207_U361, P1_R1207_U362, P1_R1207_U363, P1_R1207_U364, P1_R1207_U365, P1_R1207_U366, P1_R1207_U367, P1_R1207_U368, P1_R1207_U369, P1_R1207_U37, P1_R1207_U370, P1_R1207_U371, P1_R1207_U372, P1_R1207_U373, P1_R1207_U374, P1_R1207_U375, P1_R1207_U376, P1_R1207_U377, P1_R1207_U378, P1_R1207_U379, P1_R1207_U38, P1_R1207_U380, P1_R1207_U381, P1_R1207_U382, P1_R1207_U383, P1_R1207_U384, P1_R1207_U385, P1_R1207_U386, P1_R1207_U387, P1_R1207_U388, P1_R1207_U389, P1_R1207_U39, P1_R1207_U390, P1_R1207_U391, P1_R1207_U392, P1_R1207_U393, P1_R1207_U394, P1_R1207_U395, P1_R1207_U396, P1_R1207_U397, P1_R1207_U398, P1_R1207_U399, P1_R1207_U40, P1_R1207_U400, P1_R1207_U401, P1_R1207_U402, P1_R1207_U403, P1_R1207_U404, P1_R1207_U405, P1_R1207_U406, P1_R1207_U407, P1_R1207_U408, P1_R1207_U409, P1_R1207_U41, P1_R1207_U410, P1_R1207_U411, P1_R1207_U412, P1_R1207_U413, P1_R1207_U414, P1_R1207_U415, P1_R1207_U416, P1_R1207_U417, P1_R1207_U418, P1_R1207_U419, P1_R1207_U42, P1_R1207_U420, P1_R1207_U421, P1_R1207_U422, P1_R1207_U423, P1_R1207_U424, P1_R1207_U425, P1_R1207_U426, P1_R1207_U427, P1_R1207_U428, P1_R1207_U429, P1_R1207_U43, P1_R1207_U430, P1_R1207_U431, P1_R1207_U432, P1_R1207_U433, P1_R1207_U434, P1_R1207_U435, P1_R1207_U436, P1_R1207_U437, P1_R1207_U438, P1_R1207_U439, P1_R1207_U44, P1_R1207_U440, P1_R1207_U441, P1_R1207_U442, P1_R1207_U443, P1_R1207_U444, P1_R1207_U445, P1_R1207_U446, P1_R1207_U447, P1_R1207_U448, P1_R1207_U449, P1_R1207_U45, P1_R1207_U450, P1_R1207_U451, P1_R1207_U452, P1_R1207_U453, P1_R1207_U454, P1_R1207_U455, P1_R1207_U456, P1_R1207_U457, P1_R1207_U458, P1_R1207_U459, P1_R1207_U46, P1_R1207_U460, P1_R1207_U461, P1_R1207_U462, P1_R1207_U463, P1_R1207_U464, P1_R1207_U465, P1_R1207_U466, P1_R1207_U467, P1_R1207_U468, P1_R1207_U469, P1_R1207_U47, P1_R1207_U470, P1_R1207_U471, P1_R1207_U472, P1_R1207_U473, P1_R1207_U474, P1_R1207_U475, P1_R1207_U476, P1_R1207_U48, P1_R1207_U49, P1_R1207_U50, P1_R1207_U51, P1_R1207_U52, P1_R1207_U53, P1_R1207_U54, P1_R1207_U55, P1_R1207_U56, P1_R1207_U57, P1_R1207_U58, P1_R1207_U59, P1_R1207_U6, P1_R1207_U60, P1_R1207_U61, P1_R1207_U62, P1_R1207_U63, P1_R1207_U64, P1_R1207_U65, P1_R1207_U66, P1_R1207_U67, P1_R1207_U68, P1_R1207_U69, P1_R1207_U7, P1_R1207_U70, P1_R1207_U71, P1_R1207_U72, P1_R1207_U73, P1_R1207_U74, P1_R1207_U75, P1_R1207_U76, P1_R1207_U77, P1_R1207_U78, P1_R1207_U79, P1_R1207_U8, P1_R1207_U80, P1_R1207_U81, P1_R1207_U82, P1_R1207_U83, P1_R1207_U84, P1_R1207_U85, P1_R1207_U86, P1_R1207_U87, P1_R1207_U88, P1_R1207_U89, P1_R1207_U9, P1_R1207_U90, P1_R1207_U91, P1_R1207_U92, P1_R1207_U93, P1_R1207_U94, P1_R1207_U95, P1_R1207_U96, P1_R1207_U97, P1_R1207_U98, P1_R1207_U99, P1_R1222_U10, P1_R1222_U100, P1_R1222_U101, P1_R1222_U102, P1_R1222_U103, P1_R1222_U104, P1_R1222_U105, P1_R1222_U106, P1_R1222_U107, P1_R1222_U108, P1_R1222_U109, P1_R1222_U11, P1_R1222_U110, P1_R1222_U111, P1_R1222_U112, P1_R1222_U113, P1_R1222_U114, P1_R1222_U115, P1_R1222_U116, P1_R1222_U117, P1_R1222_U118, P1_R1222_U119, P1_R1222_U12, P1_R1222_U120, P1_R1222_U121, P1_R1222_U122, P1_R1222_U123, P1_R1222_U124, P1_R1222_U125, P1_R1222_U126, P1_R1222_U127, P1_R1222_U128, P1_R1222_U129, P1_R1222_U13, P1_R1222_U130, P1_R1222_U131, P1_R1222_U132, P1_R1222_U133, P1_R1222_U134, P1_R1222_U135, P1_R1222_U136, P1_R1222_U137, P1_R1222_U138, P1_R1222_U139, P1_R1222_U14, P1_R1222_U140, P1_R1222_U141, P1_R1222_U142, P1_R1222_U143, P1_R1222_U144, P1_R1222_U145, P1_R1222_U146, P1_R1222_U147, P1_R1222_U148, P1_R1222_U149, P1_R1222_U15, P1_R1222_U150, P1_R1222_U151, P1_R1222_U152, P1_R1222_U153, P1_R1222_U154, P1_R1222_U155, P1_R1222_U156, P1_R1222_U157, P1_R1222_U158, P1_R1222_U159, P1_R1222_U16, P1_R1222_U160, P1_R1222_U161, P1_R1222_U162, P1_R1222_U163, P1_R1222_U164, P1_R1222_U165, P1_R1222_U166, P1_R1222_U167, P1_R1222_U168, P1_R1222_U169, P1_R1222_U17, P1_R1222_U170, P1_R1222_U171, P1_R1222_U172, P1_R1222_U173, P1_R1222_U174, P1_R1222_U175, P1_R1222_U176, P1_R1222_U177, P1_R1222_U178, P1_R1222_U179, P1_R1222_U18, P1_R1222_U180, P1_R1222_U181, P1_R1222_U182, P1_R1222_U183, P1_R1222_U184, P1_R1222_U185, P1_R1222_U186, P1_R1222_U187, P1_R1222_U188, P1_R1222_U189, P1_R1222_U19, P1_R1222_U190, P1_R1222_U191, P1_R1222_U192, P1_R1222_U193, P1_R1222_U194, P1_R1222_U195, P1_R1222_U196, P1_R1222_U197, P1_R1222_U198, P1_R1222_U199, P1_R1222_U20, P1_R1222_U200, P1_R1222_U201, P1_R1222_U202, P1_R1222_U203, P1_R1222_U204, P1_R1222_U205, P1_R1222_U206, P1_R1222_U207, P1_R1222_U208, P1_R1222_U209, P1_R1222_U21, P1_R1222_U210, P1_R1222_U211, P1_R1222_U212, P1_R1222_U213, P1_R1222_U214, P1_R1222_U215, P1_R1222_U216, P1_R1222_U217, P1_R1222_U218, P1_R1222_U219, P1_R1222_U22, P1_R1222_U220, P1_R1222_U221, P1_R1222_U222, P1_R1222_U223, P1_R1222_U224, P1_R1222_U225, P1_R1222_U226, P1_R1222_U227, P1_R1222_U228, P1_R1222_U229, P1_R1222_U23, P1_R1222_U230, P1_R1222_U231, P1_R1222_U232, P1_R1222_U233, P1_R1222_U234, P1_R1222_U235, P1_R1222_U236, P1_R1222_U237, P1_R1222_U238, P1_R1222_U239, P1_R1222_U24, P1_R1222_U240, P1_R1222_U241, P1_R1222_U242, P1_R1222_U243, P1_R1222_U244, P1_R1222_U245, P1_R1222_U246, P1_R1222_U247, P1_R1222_U248, P1_R1222_U249, P1_R1222_U25, P1_R1222_U250, P1_R1222_U251, P1_R1222_U252, P1_R1222_U253, P1_R1222_U254, P1_R1222_U255, P1_R1222_U256, P1_R1222_U257, P1_R1222_U258, P1_R1222_U259, P1_R1222_U26, P1_R1222_U260, P1_R1222_U261, P1_R1222_U262, P1_R1222_U263, P1_R1222_U264, P1_R1222_U265, P1_R1222_U266, P1_R1222_U267, P1_R1222_U268, P1_R1222_U269, P1_R1222_U27, P1_R1222_U270, P1_R1222_U271, P1_R1222_U272, P1_R1222_U273, P1_R1222_U274, P1_R1222_U275, P1_R1222_U276, P1_R1222_U277, P1_R1222_U278, P1_R1222_U279, P1_R1222_U28, P1_R1222_U280, P1_R1222_U281, P1_R1222_U282, P1_R1222_U283, P1_R1222_U284, P1_R1222_U285, P1_R1222_U286, P1_R1222_U287, P1_R1222_U288, P1_R1222_U289, P1_R1222_U29, P1_R1222_U290, P1_R1222_U291, P1_R1222_U292, P1_R1222_U293, P1_R1222_U294, P1_R1222_U295, P1_R1222_U296, P1_R1222_U297, P1_R1222_U298, P1_R1222_U299, P1_R1222_U30, P1_R1222_U300, P1_R1222_U301, P1_R1222_U302, P1_R1222_U303, P1_R1222_U304, P1_R1222_U305, P1_R1222_U306, P1_R1222_U307, P1_R1222_U308, P1_R1222_U309, P1_R1222_U31, P1_R1222_U310, P1_R1222_U311, P1_R1222_U312, P1_R1222_U313, P1_R1222_U314, P1_R1222_U315, P1_R1222_U316, P1_R1222_U317, P1_R1222_U318, P1_R1222_U319, P1_R1222_U32, P1_R1222_U320, P1_R1222_U321, P1_R1222_U322, P1_R1222_U323, P1_R1222_U324, P1_R1222_U325, P1_R1222_U326, P1_R1222_U327, P1_R1222_U328, P1_R1222_U329, P1_R1222_U33, P1_R1222_U330, P1_R1222_U331, P1_R1222_U332, P1_R1222_U333, P1_R1222_U334, P1_R1222_U335, P1_R1222_U336, P1_R1222_U337, P1_R1222_U338, P1_R1222_U339, P1_R1222_U34, P1_R1222_U340, P1_R1222_U341, P1_R1222_U342, P1_R1222_U343, P1_R1222_U344, P1_R1222_U345, P1_R1222_U346, P1_R1222_U347, P1_R1222_U348, P1_R1222_U349, P1_R1222_U35, P1_R1222_U350, P1_R1222_U351, P1_R1222_U352, P1_R1222_U353, P1_R1222_U354, P1_R1222_U355, P1_R1222_U356, P1_R1222_U357, P1_R1222_U358, P1_R1222_U359, P1_R1222_U36, P1_R1222_U360, P1_R1222_U361, P1_R1222_U362, P1_R1222_U363, P1_R1222_U364, P1_R1222_U365, P1_R1222_U366, P1_R1222_U367, P1_R1222_U368, P1_R1222_U369, P1_R1222_U37, P1_R1222_U370, P1_R1222_U371, P1_R1222_U372, P1_R1222_U373, P1_R1222_U374, P1_R1222_U375, P1_R1222_U376, P1_R1222_U377, P1_R1222_U378, P1_R1222_U379, P1_R1222_U38, P1_R1222_U380, P1_R1222_U381, P1_R1222_U382, P1_R1222_U383, P1_R1222_U384, P1_R1222_U385, P1_R1222_U386, P1_R1222_U387, P1_R1222_U388, P1_R1222_U389, P1_R1222_U39, P1_R1222_U390, P1_R1222_U391, P1_R1222_U392, P1_R1222_U393, P1_R1222_U394, P1_R1222_U395, P1_R1222_U396, P1_R1222_U397, P1_R1222_U398, P1_R1222_U399, P1_R1222_U4, P1_R1222_U40, P1_R1222_U400, P1_R1222_U401, P1_R1222_U402, P1_R1222_U403, P1_R1222_U404, P1_R1222_U405, P1_R1222_U406, P1_R1222_U407, P1_R1222_U408, P1_R1222_U409, P1_R1222_U41, P1_R1222_U410, P1_R1222_U411, P1_R1222_U412, P1_R1222_U413, P1_R1222_U414, P1_R1222_U415, P1_R1222_U416, P1_R1222_U417, P1_R1222_U418, P1_R1222_U419, P1_R1222_U42, P1_R1222_U420, P1_R1222_U421, P1_R1222_U422, P1_R1222_U423, P1_R1222_U424, P1_R1222_U425, P1_R1222_U426, P1_R1222_U427, P1_R1222_U428, P1_R1222_U429, P1_R1222_U43, P1_R1222_U430, P1_R1222_U431, P1_R1222_U432, P1_R1222_U433, P1_R1222_U434, P1_R1222_U435, P1_R1222_U436, P1_R1222_U437, P1_R1222_U438, P1_R1222_U439, P1_R1222_U44, P1_R1222_U440, P1_R1222_U441, P1_R1222_U442, P1_R1222_U443, P1_R1222_U444, P1_R1222_U445, P1_R1222_U446, P1_R1222_U447, P1_R1222_U448, P1_R1222_U449, P1_R1222_U45, P1_R1222_U450, P1_R1222_U451, P1_R1222_U452, P1_R1222_U453, P1_R1222_U454, P1_R1222_U455, P1_R1222_U456, P1_R1222_U457, P1_R1222_U458, P1_R1222_U459, P1_R1222_U46, P1_R1222_U460, P1_R1222_U461, P1_R1222_U462, P1_R1222_U463, P1_R1222_U464, P1_R1222_U465, P1_R1222_U466, P1_R1222_U467, P1_R1222_U468, P1_R1222_U469, P1_R1222_U47, P1_R1222_U470, P1_R1222_U471, P1_R1222_U472, P1_R1222_U473, P1_R1222_U474, P1_R1222_U475, P1_R1222_U476, P1_R1222_U477, P1_R1222_U478, P1_R1222_U479, P1_R1222_U48, P1_R1222_U480, P1_R1222_U481, P1_R1222_U482, P1_R1222_U483, P1_R1222_U484, P1_R1222_U485, P1_R1222_U486, P1_R1222_U487, P1_R1222_U488, P1_R1222_U489, P1_R1222_U49, P1_R1222_U490, P1_R1222_U491, P1_R1222_U492, P1_R1222_U493, P1_R1222_U494, P1_R1222_U495, P1_R1222_U496, P1_R1222_U497, P1_R1222_U498, P1_R1222_U499, P1_R1222_U5, P1_R1222_U50, P1_R1222_U500, P1_R1222_U501, P1_R1222_U51, P1_R1222_U52, P1_R1222_U53, P1_R1222_U54, P1_R1222_U55, P1_R1222_U56, P1_R1222_U57, P1_R1222_U58, P1_R1222_U59, P1_R1222_U6, P1_R1222_U60, P1_R1222_U61, P1_R1222_U62, P1_R1222_U63, P1_R1222_U64, P1_R1222_U65, P1_R1222_U66, P1_R1222_U67, P1_R1222_U68, P1_R1222_U69, P1_R1222_U7, P1_R1222_U70, P1_R1222_U71, P1_R1222_U72, P1_R1222_U73, P1_R1222_U74, P1_R1222_U75, P1_R1222_U76, P1_R1222_U77, P1_R1222_U78, P1_R1222_U79, P1_R1222_U8, P1_R1222_U80, P1_R1222_U81, P1_R1222_U82, P1_R1222_U83, P1_R1222_U84, P1_R1222_U85, P1_R1222_U86, P1_R1222_U87, P1_R1222_U88, P1_R1222_U89, P1_R1222_U9, P1_R1222_U90, P1_R1222_U91, P1_R1222_U92, P1_R1222_U93, P1_R1222_U94, P1_R1222_U95, P1_R1222_U96, P1_R1222_U97, P1_R1222_U98, P1_R1222_U99, P1_R1240_U10, P1_R1240_U100, P1_R1240_U101, P1_R1240_U102, P1_R1240_U103, P1_R1240_U104, P1_R1240_U105, P1_R1240_U106, P1_R1240_U107, P1_R1240_U108, P1_R1240_U109, P1_R1240_U11, P1_R1240_U110, P1_R1240_U111, P1_R1240_U112, P1_R1240_U113, P1_R1240_U114, P1_R1240_U115, P1_R1240_U116, P1_R1240_U117, P1_R1240_U118, P1_R1240_U119, P1_R1240_U12, P1_R1240_U120, P1_R1240_U121, P1_R1240_U122, P1_R1240_U123, P1_R1240_U124, P1_R1240_U125, P1_R1240_U126, P1_R1240_U127, P1_R1240_U128, P1_R1240_U129, P1_R1240_U13, P1_R1240_U130, P1_R1240_U131, P1_R1240_U132, P1_R1240_U133, P1_R1240_U134, P1_R1240_U135, P1_R1240_U136, P1_R1240_U137, P1_R1240_U138, P1_R1240_U139, P1_R1240_U14, P1_R1240_U140, P1_R1240_U141, P1_R1240_U142, P1_R1240_U143, P1_R1240_U144, P1_R1240_U145, P1_R1240_U146, P1_R1240_U147, P1_R1240_U148, P1_R1240_U149, P1_R1240_U15, P1_R1240_U150, P1_R1240_U151, P1_R1240_U152, P1_R1240_U153, P1_R1240_U154, P1_R1240_U155, P1_R1240_U156, P1_R1240_U157, P1_R1240_U158, P1_R1240_U159, P1_R1240_U16, P1_R1240_U160, P1_R1240_U161, P1_R1240_U162, P1_R1240_U163, P1_R1240_U164, P1_R1240_U165, P1_R1240_U166, P1_R1240_U167, P1_R1240_U168, P1_R1240_U169, P1_R1240_U17, P1_R1240_U170, P1_R1240_U171, P1_R1240_U172, P1_R1240_U173, P1_R1240_U174, P1_R1240_U175, P1_R1240_U176, P1_R1240_U177, P1_R1240_U178, P1_R1240_U179, P1_R1240_U18, P1_R1240_U180, P1_R1240_U181, P1_R1240_U182, P1_R1240_U183, P1_R1240_U184, P1_R1240_U185, P1_R1240_U186, P1_R1240_U187, P1_R1240_U188, P1_R1240_U189, P1_R1240_U19, P1_R1240_U190, P1_R1240_U191, P1_R1240_U192, P1_R1240_U193, P1_R1240_U194, P1_R1240_U195, P1_R1240_U196, P1_R1240_U197, P1_R1240_U198, P1_R1240_U199, P1_R1240_U20, P1_R1240_U200, P1_R1240_U201, P1_R1240_U202, P1_R1240_U203, P1_R1240_U204, P1_R1240_U205, P1_R1240_U206, P1_R1240_U207, P1_R1240_U208, P1_R1240_U209, P1_R1240_U21, P1_R1240_U210, P1_R1240_U211, P1_R1240_U212, P1_R1240_U213, P1_R1240_U214, P1_R1240_U215, P1_R1240_U216, P1_R1240_U217, P1_R1240_U218, P1_R1240_U219, P1_R1240_U22, P1_R1240_U220, P1_R1240_U221, P1_R1240_U222, P1_R1240_U223, P1_R1240_U224, P1_R1240_U225, P1_R1240_U226, P1_R1240_U227, P1_R1240_U228, P1_R1240_U229, P1_R1240_U23, P1_R1240_U230, P1_R1240_U231, P1_R1240_U232, P1_R1240_U233, P1_R1240_U234, P1_R1240_U235, P1_R1240_U236, P1_R1240_U237, P1_R1240_U238, P1_R1240_U239, P1_R1240_U24, P1_R1240_U240, P1_R1240_U241, P1_R1240_U242, P1_R1240_U243, P1_R1240_U244, P1_R1240_U245, P1_R1240_U246, P1_R1240_U247, P1_R1240_U248, P1_R1240_U249, P1_R1240_U25, P1_R1240_U250, P1_R1240_U251, P1_R1240_U252, P1_R1240_U253, P1_R1240_U254, P1_R1240_U255, P1_R1240_U256, P1_R1240_U257, P1_R1240_U258, P1_R1240_U259, P1_R1240_U26, P1_R1240_U260, P1_R1240_U261, P1_R1240_U262, P1_R1240_U263, P1_R1240_U264, P1_R1240_U265, P1_R1240_U266, P1_R1240_U267, P1_R1240_U268, P1_R1240_U269, P1_R1240_U27, P1_R1240_U270, P1_R1240_U271, P1_R1240_U272, P1_R1240_U273, P1_R1240_U274, P1_R1240_U275, P1_R1240_U276, P1_R1240_U277, P1_R1240_U278, P1_R1240_U279, P1_R1240_U28, P1_R1240_U280, P1_R1240_U281, P1_R1240_U282, P1_R1240_U283, P1_R1240_U284, P1_R1240_U285, P1_R1240_U286, P1_R1240_U287, P1_R1240_U288, P1_R1240_U289, P1_R1240_U29, P1_R1240_U290, P1_R1240_U291, P1_R1240_U292, P1_R1240_U293, P1_R1240_U294, P1_R1240_U295, P1_R1240_U296, P1_R1240_U297, P1_R1240_U298, P1_R1240_U299, P1_R1240_U30, P1_R1240_U300, P1_R1240_U301, P1_R1240_U302, P1_R1240_U303, P1_R1240_U304, P1_R1240_U305, P1_R1240_U306, P1_R1240_U307, P1_R1240_U308, P1_R1240_U309, P1_R1240_U31, P1_R1240_U310, P1_R1240_U311, P1_R1240_U312, P1_R1240_U313, P1_R1240_U314, P1_R1240_U315, P1_R1240_U316, P1_R1240_U317, P1_R1240_U318, P1_R1240_U319, P1_R1240_U32, P1_R1240_U320, P1_R1240_U321, P1_R1240_U322, P1_R1240_U323, P1_R1240_U324, P1_R1240_U325, P1_R1240_U326, P1_R1240_U327, P1_R1240_U328, P1_R1240_U329, P1_R1240_U33, P1_R1240_U330, P1_R1240_U331, P1_R1240_U332, P1_R1240_U333, P1_R1240_U334, P1_R1240_U335, P1_R1240_U336, P1_R1240_U337, P1_R1240_U338, P1_R1240_U339, P1_R1240_U34, P1_R1240_U340, P1_R1240_U341, P1_R1240_U342, P1_R1240_U343, P1_R1240_U344, P1_R1240_U345, P1_R1240_U346, P1_R1240_U347, P1_R1240_U348, P1_R1240_U349, P1_R1240_U35, P1_R1240_U350, P1_R1240_U351, P1_R1240_U352, P1_R1240_U353, P1_R1240_U354, P1_R1240_U355, P1_R1240_U356, P1_R1240_U357, P1_R1240_U358, P1_R1240_U359, P1_R1240_U36, P1_R1240_U360, P1_R1240_U361, P1_R1240_U362, P1_R1240_U363, P1_R1240_U364, P1_R1240_U365, P1_R1240_U366, P1_R1240_U367, P1_R1240_U368, P1_R1240_U369, P1_R1240_U37, P1_R1240_U370, P1_R1240_U371, P1_R1240_U372, P1_R1240_U373, P1_R1240_U374, P1_R1240_U375, P1_R1240_U376, P1_R1240_U377, P1_R1240_U378, P1_R1240_U379, P1_R1240_U38, P1_R1240_U380, P1_R1240_U381, P1_R1240_U382, P1_R1240_U383, P1_R1240_U384, P1_R1240_U385, P1_R1240_U386, P1_R1240_U387, P1_R1240_U388, P1_R1240_U389, P1_R1240_U39, P1_R1240_U390, P1_R1240_U391, P1_R1240_U392, P1_R1240_U393, P1_R1240_U394, P1_R1240_U395, P1_R1240_U396, P1_R1240_U397, P1_R1240_U398, P1_R1240_U399, P1_R1240_U4, P1_R1240_U40, P1_R1240_U400, P1_R1240_U401, P1_R1240_U402, P1_R1240_U403, P1_R1240_U404, P1_R1240_U405, P1_R1240_U406, P1_R1240_U407, P1_R1240_U408, P1_R1240_U409, P1_R1240_U41, P1_R1240_U410, P1_R1240_U411, P1_R1240_U412, P1_R1240_U413, P1_R1240_U414, P1_R1240_U415, P1_R1240_U416, P1_R1240_U417, P1_R1240_U418, P1_R1240_U419, P1_R1240_U42, P1_R1240_U420, P1_R1240_U421, P1_R1240_U422, P1_R1240_U423, P1_R1240_U424, P1_R1240_U425, P1_R1240_U426, P1_R1240_U427, P1_R1240_U428, P1_R1240_U429, P1_R1240_U43, P1_R1240_U430, P1_R1240_U431, P1_R1240_U432, P1_R1240_U433, P1_R1240_U434, P1_R1240_U435, P1_R1240_U436, P1_R1240_U437, P1_R1240_U438, P1_R1240_U439, P1_R1240_U44, P1_R1240_U440, P1_R1240_U441, P1_R1240_U442, P1_R1240_U443, P1_R1240_U444, P1_R1240_U445, P1_R1240_U446, P1_R1240_U447, P1_R1240_U448, P1_R1240_U449, P1_R1240_U45, P1_R1240_U450, P1_R1240_U451, P1_R1240_U452, P1_R1240_U453, P1_R1240_U454, P1_R1240_U455, P1_R1240_U456, P1_R1240_U457, P1_R1240_U458, P1_R1240_U459, P1_R1240_U46, P1_R1240_U460, P1_R1240_U461, P1_R1240_U462, P1_R1240_U463, P1_R1240_U464, P1_R1240_U465, P1_R1240_U466, P1_R1240_U467, P1_R1240_U468, P1_R1240_U469, P1_R1240_U47, P1_R1240_U470, P1_R1240_U471, P1_R1240_U472, P1_R1240_U473, P1_R1240_U474, P1_R1240_U475, P1_R1240_U476, P1_R1240_U477, P1_R1240_U478, P1_R1240_U479, P1_R1240_U48, P1_R1240_U480, P1_R1240_U481, P1_R1240_U482, P1_R1240_U483, P1_R1240_U484, P1_R1240_U485, P1_R1240_U486, P1_R1240_U487, P1_R1240_U488, P1_R1240_U489, P1_R1240_U49, P1_R1240_U490, P1_R1240_U491, P1_R1240_U492, P1_R1240_U493, P1_R1240_U494, P1_R1240_U495, P1_R1240_U496, P1_R1240_U497, P1_R1240_U498, P1_R1240_U499, P1_R1240_U5, P1_R1240_U50, P1_R1240_U500, P1_R1240_U501, P1_R1240_U51, P1_R1240_U52, P1_R1240_U53, P1_R1240_U54, P1_R1240_U55, P1_R1240_U56, P1_R1240_U57, P1_R1240_U58, P1_R1240_U59, P1_R1240_U6, P1_R1240_U60, P1_R1240_U61, P1_R1240_U62, P1_R1240_U63, P1_R1240_U64, P1_R1240_U65, P1_R1240_U66, P1_R1240_U67, P1_R1240_U68, P1_R1240_U69, P1_R1240_U7, P1_R1240_U70, P1_R1240_U71, P1_R1240_U72, P1_R1240_U73, P1_R1240_U74, P1_R1240_U75, P1_R1240_U76, P1_R1240_U77, P1_R1240_U78, P1_R1240_U79, P1_R1240_U8, P1_R1240_U80, P1_R1240_U81, P1_R1240_U82, P1_R1240_U83, P1_R1240_U84, P1_R1240_U85, P1_R1240_U86, P1_R1240_U87, P1_R1240_U88, P1_R1240_U89, P1_R1240_U9, P1_R1240_U90, P1_R1240_U91, P1_R1240_U92, P1_R1240_U93, P1_R1240_U94, P1_R1240_U95, P1_R1240_U96, P1_R1240_U97, P1_R1240_U98, P1_R1240_U99, P1_R1282_U10, P1_R1282_U100, P1_R1282_U101, P1_R1282_U102, P1_R1282_U103, P1_R1282_U104, P1_R1282_U105, P1_R1282_U106, P1_R1282_U107, P1_R1282_U108, P1_R1282_U109, P1_R1282_U11, P1_R1282_U110, P1_R1282_U111, P1_R1282_U112, P1_R1282_U113, P1_R1282_U114, P1_R1282_U115, P1_R1282_U116, P1_R1282_U117, P1_R1282_U118, P1_R1282_U119, P1_R1282_U12, P1_R1282_U120, P1_R1282_U121, P1_R1282_U122, P1_R1282_U123, P1_R1282_U124, P1_R1282_U125, P1_R1282_U126, P1_R1282_U127, P1_R1282_U128, P1_R1282_U129, P1_R1282_U13, P1_R1282_U130, P1_R1282_U131, P1_R1282_U132, P1_R1282_U133, P1_R1282_U134, P1_R1282_U135, P1_R1282_U136, P1_R1282_U137, P1_R1282_U138, P1_R1282_U139, P1_R1282_U14, P1_R1282_U140, P1_R1282_U141, P1_R1282_U142, P1_R1282_U143, P1_R1282_U144, P1_R1282_U145, P1_R1282_U146, P1_R1282_U147, P1_R1282_U148, P1_R1282_U149, P1_R1282_U15, P1_R1282_U150, P1_R1282_U151, P1_R1282_U152, P1_R1282_U153, P1_R1282_U154, P1_R1282_U155, P1_R1282_U156, P1_R1282_U157, P1_R1282_U158, P1_R1282_U159, P1_R1282_U16, P1_R1282_U17, P1_R1282_U18, P1_R1282_U19, P1_R1282_U20, P1_R1282_U21, P1_R1282_U22, P1_R1282_U23, P1_R1282_U24, P1_R1282_U25, P1_R1282_U26, P1_R1282_U27, P1_R1282_U28, P1_R1282_U29, P1_R1282_U30, P1_R1282_U31, P1_R1282_U32, P1_R1282_U33, P1_R1282_U34, P1_R1282_U35, P1_R1282_U36, P1_R1282_U37, P1_R1282_U38, P1_R1282_U39, P1_R1282_U40, P1_R1282_U41, P1_R1282_U42, P1_R1282_U43, P1_R1282_U44, P1_R1282_U45, P1_R1282_U46, P1_R1282_U47, P1_R1282_U48, P1_R1282_U49, P1_R1282_U50, P1_R1282_U51, P1_R1282_U52, P1_R1282_U53, P1_R1282_U54, P1_R1282_U55, P1_R1282_U56, P1_R1282_U57, P1_R1282_U58, P1_R1282_U59, P1_R1282_U6, P1_R1282_U60, P1_R1282_U61, P1_R1282_U62, P1_R1282_U63, P1_R1282_U64, P1_R1282_U65, P1_R1282_U66, P1_R1282_U67, P1_R1282_U68, P1_R1282_U69, P1_R1282_U7, P1_R1282_U70, P1_R1282_U71, P1_R1282_U72, P1_R1282_U73, P1_R1282_U74, P1_R1282_U75, P1_R1282_U76, P1_R1282_U77, P1_R1282_U78, P1_R1282_U79, P1_R1282_U8, P1_R1282_U80, P1_R1282_U81, P1_R1282_U82, P1_R1282_U83, P1_R1282_U84, P1_R1282_U85, P1_R1282_U86, P1_R1282_U87, P1_R1282_U88, P1_R1282_U89, P1_R1282_U9, P1_R1282_U90, P1_R1282_U91, P1_R1282_U92, P1_R1282_U93, P1_R1282_U94, P1_R1282_U95, P1_R1282_U96, P1_R1282_U97, P1_R1282_U98, P1_R1282_U99, P1_R1309_U10, P1_R1309_U6, P1_R1309_U7, P1_R1309_U8, P1_R1309_U9, P1_R1352_U6, P1_R1352_U7, P1_R1375_U10, P1_R1375_U100, P1_R1375_U101, P1_R1375_U102, P1_R1375_U103, P1_R1375_U104, P1_R1375_U105, P1_R1375_U106, P1_R1375_U107, P1_R1375_U108, P1_R1375_U109, P1_R1375_U11, P1_R1375_U110, P1_R1375_U111, P1_R1375_U112, P1_R1375_U113, P1_R1375_U114, P1_R1375_U115, P1_R1375_U116, P1_R1375_U117, P1_R1375_U118, P1_R1375_U119, P1_R1375_U12, P1_R1375_U120, P1_R1375_U121, P1_R1375_U122, P1_R1375_U123, P1_R1375_U124, P1_R1375_U125, P1_R1375_U126, P1_R1375_U127, P1_R1375_U128, P1_R1375_U129, P1_R1375_U13, P1_R1375_U130, P1_R1375_U131, P1_R1375_U132, P1_R1375_U133, P1_R1375_U134, P1_R1375_U135, P1_R1375_U136, P1_R1375_U137, P1_R1375_U138, P1_R1375_U139, P1_R1375_U14, P1_R1375_U140, P1_R1375_U141, P1_R1375_U142, P1_R1375_U143, P1_R1375_U144, P1_R1375_U145, P1_R1375_U146, P1_R1375_U147, P1_R1375_U148, P1_R1375_U149, P1_R1375_U15, P1_R1375_U150, P1_R1375_U151, P1_R1375_U152, P1_R1375_U153, P1_R1375_U154, P1_R1375_U155, P1_R1375_U156, P1_R1375_U157, P1_R1375_U158, P1_R1375_U159, P1_R1375_U16, P1_R1375_U160, P1_R1375_U161, P1_R1375_U162, P1_R1375_U163, P1_R1375_U164, P1_R1375_U165, P1_R1375_U166, P1_R1375_U167, P1_R1375_U168, P1_R1375_U169, P1_R1375_U17, P1_R1375_U170, P1_R1375_U171, P1_R1375_U172, P1_R1375_U173, P1_R1375_U174, P1_R1375_U175, P1_R1375_U176, P1_R1375_U177, P1_R1375_U178, P1_R1375_U179, P1_R1375_U18, P1_R1375_U180, P1_R1375_U181, P1_R1375_U182, P1_R1375_U183, P1_R1375_U184, P1_R1375_U185, P1_R1375_U186, P1_R1375_U187, P1_R1375_U188, P1_R1375_U189, P1_R1375_U19, P1_R1375_U190, P1_R1375_U191, P1_R1375_U192, P1_R1375_U193, P1_R1375_U194, P1_R1375_U195, P1_R1375_U196, P1_R1375_U197, P1_R1375_U20, P1_R1375_U21, P1_R1375_U22, P1_R1375_U23, P1_R1375_U24, P1_R1375_U25, P1_R1375_U26, P1_R1375_U27, P1_R1375_U28, P1_R1375_U29, P1_R1375_U30, P1_R1375_U31, P1_R1375_U32, P1_R1375_U33, P1_R1375_U34, P1_R1375_U35, P1_R1375_U36, P1_R1375_U37, P1_R1375_U38, P1_R1375_U39, P1_R1375_U40, P1_R1375_U41, P1_R1375_U42, P1_R1375_U43, P1_R1375_U44, P1_R1375_U45, P1_R1375_U46, P1_R1375_U47, P1_R1375_U48, P1_R1375_U49, P1_R1375_U50, P1_R1375_U51, P1_R1375_U52, P1_R1375_U53, P1_R1375_U54, P1_R1375_U55, P1_R1375_U56, P1_R1375_U57, P1_R1375_U58, P1_R1375_U59, P1_R1375_U6, P1_R1375_U60, P1_R1375_U61, P1_R1375_U62, P1_R1375_U63, P1_R1375_U64, P1_R1375_U65, P1_R1375_U66, P1_R1375_U67, P1_R1375_U68, P1_R1375_U69, P1_R1375_U7, P1_R1375_U70, P1_R1375_U71, P1_R1375_U72, P1_R1375_U73, P1_R1375_U74, P1_R1375_U75, P1_R1375_U76, P1_R1375_U77, P1_R1375_U78, P1_R1375_U79, P1_R1375_U8, P1_R1375_U80, P1_R1375_U81, P1_R1375_U82, P1_R1375_U83, P1_R1375_U84, P1_R1375_U85, P1_R1375_U86, P1_R1375_U87, P1_R1375_U88, P1_R1375_U89, P1_R1375_U9, P1_R1375_U90, P1_R1375_U91, P1_R1375_U92, P1_R1375_U93, P1_R1375_U94, P1_R1375_U95, P1_R1375_U96, P1_R1375_U97, P1_R1375_U98, P1_R1375_U99, P1_SUB_88_U10, P1_SUB_88_U100, P1_SUB_88_U101, P1_SUB_88_U102, P1_SUB_88_U103, P1_SUB_88_U104, P1_SUB_88_U105, P1_SUB_88_U106, P1_SUB_88_U107, P1_SUB_88_U108, P1_SUB_88_U109, P1_SUB_88_U11, P1_SUB_88_U110, P1_SUB_88_U111, P1_SUB_88_U112, P1_SUB_88_U113, P1_SUB_88_U114, P1_SUB_88_U115, P1_SUB_88_U116, P1_SUB_88_U117, P1_SUB_88_U118, P1_SUB_88_U119, P1_SUB_88_U12, P1_SUB_88_U120, P1_SUB_88_U121, P1_SUB_88_U122, P1_SUB_88_U123, P1_SUB_88_U124, P1_SUB_88_U125, P1_SUB_88_U126, P1_SUB_88_U127, P1_SUB_88_U128, P1_SUB_88_U129, P1_SUB_88_U13, P1_SUB_88_U130, P1_SUB_88_U131, P1_SUB_88_U132, P1_SUB_88_U133, P1_SUB_88_U134, P1_SUB_88_U135, P1_SUB_88_U136, P1_SUB_88_U137, P1_SUB_88_U138, P1_SUB_88_U139, P1_SUB_88_U14, P1_SUB_88_U140, P1_SUB_88_U141, P1_SUB_88_U142, P1_SUB_88_U143, P1_SUB_88_U144, P1_SUB_88_U145, P1_SUB_88_U146, P1_SUB_88_U147, P1_SUB_88_U148, P1_SUB_88_U149, P1_SUB_88_U15, P1_SUB_88_U150, P1_SUB_88_U151, P1_SUB_88_U152, P1_SUB_88_U153, P1_SUB_88_U154, P1_SUB_88_U155, P1_SUB_88_U156, P1_SUB_88_U157, P1_SUB_88_U158, P1_SUB_88_U159, P1_SUB_88_U16, P1_SUB_88_U160, P1_SUB_88_U161, P1_SUB_88_U162, P1_SUB_88_U163, P1_SUB_88_U164, P1_SUB_88_U165, P1_SUB_88_U166, P1_SUB_88_U167, P1_SUB_88_U168, P1_SUB_88_U169, P1_SUB_88_U17, P1_SUB_88_U170, P1_SUB_88_U171, P1_SUB_88_U172, P1_SUB_88_U173, P1_SUB_88_U174, P1_SUB_88_U175, P1_SUB_88_U176, P1_SUB_88_U177, P1_SUB_88_U178, P1_SUB_88_U179, P1_SUB_88_U18, P1_SUB_88_U180, P1_SUB_88_U181, P1_SUB_88_U182, P1_SUB_88_U183, P1_SUB_88_U184, P1_SUB_88_U185, P1_SUB_88_U186, P1_SUB_88_U187, P1_SUB_88_U188, P1_SUB_88_U189, P1_SUB_88_U19, P1_SUB_88_U190, P1_SUB_88_U191, P1_SUB_88_U192, P1_SUB_88_U193, P1_SUB_88_U194, P1_SUB_88_U195, P1_SUB_88_U196, P1_SUB_88_U197, P1_SUB_88_U198, P1_SUB_88_U199, P1_SUB_88_U20, P1_SUB_88_U200, P1_SUB_88_U201, P1_SUB_88_U202, P1_SUB_88_U203, P1_SUB_88_U204, P1_SUB_88_U205, P1_SUB_88_U206, P1_SUB_88_U207, P1_SUB_88_U208, P1_SUB_88_U209, P1_SUB_88_U21, P1_SUB_88_U210, P1_SUB_88_U211, P1_SUB_88_U212, P1_SUB_88_U213, P1_SUB_88_U214, P1_SUB_88_U215, P1_SUB_88_U216, P1_SUB_88_U217, P1_SUB_88_U218, P1_SUB_88_U219, P1_SUB_88_U22, P1_SUB_88_U220, P1_SUB_88_U221, P1_SUB_88_U222, P1_SUB_88_U223, P1_SUB_88_U224, P1_SUB_88_U225, P1_SUB_88_U226, P1_SUB_88_U227, P1_SUB_88_U228, P1_SUB_88_U229, P1_SUB_88_U23, P1_SUB_88_U230, P1_SUB_88_U231, P1_SUB_88_U232, P1_SUB_88_U233, P1_SUB_88_U234, P1_SUB_88_U235, P1_SUB_88_U236, P1_SUB_88_U237, P1_SUB_88_U238, P1_SUB_88_U239, P1_SUB_88_U24, P1_SUB_88_U240, P1_SUB_88_U241, P1_SUB_88_U242, P1_SUB_88_U243, P1_SUB_88_U244, P1_SUB_88_U245, P1_SUB_88_U246, P1_SUB_88_U247, P1_SUB_88_U248, P1_SUB_88_U249, P1_SUB_88_U25, P1_SUB_88_U250, P1_SUB_88_U251, P1_SUB_88_U26, P1_SUB_88_U27, P1_SUB_88_U28, P1_SUB_88_U29, P1_SUB_88_U30, P1_SUB_88_U31, P1_SUB_88_U32, P1_SUB_88_U33, P1_SUB_88_U34, P1_SUB_88_U35, P1_SUB_88_U36, P1_SUB_88_U37, P1_SUB_88_U38, P1_SUB_88_U39, P1_SUB_88_U40, P1_SUB_88_U41, P1_SUB_88_U42, P1_SUB_88_U43, P1_SUB_88_U44, P1_SUB_88_U45, P1_SUB_88_U46, P1_SUB_88_U47, P1_SUB_88_U48, P1_SUB_88_U49, P1_SUB_88_U50, P1_SUB_88_U51, P1_SUB_88_U52, P1_SUB_88_U53, P1_SUB_88_U54, P1_SUB_88_U55, P1_SUB_88_U56, P1_SUB_88_U57, P1_SUB_88_U58, P1_SUB_88_U59, P1_SUB_88_U6, P1_SUB_88_U60, P1_SUB_88_U61, P1_SUB_88_U62, P1_SUB_88_U63, P1_SUB_88_U64, P1_SUB_88_U65, P1_SUB_88_U66, P1_SUB_88_U67, P1_SUB_88_U68, P1_SUB_88_U69, P1_SUB_88_U7, P1_SUB_88_U70, P1_SUB_88_U71, P1_SUB_88_U72, P1_SUB_88_U73, P1_SUB_88_U74, P1_SUB_88_U75, P1_SUB_88_U76, P1_SUB_88_U77, P1_SUB_88_U78, P1_SUB_88_U79, P1_SUB_88_U8, P1_SUB_88_U80, P1_SUB_88_U81, P1_SUB_88_U82, P1_SUB_88_U83, P1_SUB_88_U84, P1_SUB_88_U85, P1_SUB_88_U86, P1_SUB_88_U87, P1_SUB_88_U88, P1_SUB_88_U89, P1_SUB_88_U9, P1_SUB_88_U90, P1_SUB_88_U91, P1_SUB_88_U92, P1_SUB_88_U93, P1_SUB_88_U94, P1_SUB_88_U95, P1_SUB_88_U96, P1_SUB_88_U97, P1_SUB_88_U98, P1_SUB_88_U99, P1_U3014, P1_U3015, P1_U3016, P1_U3017, P1_U3018, P1_U3019, P1_U3020, P1_U3021, P1_U3022, P1_U3023, P1_U3024, P1_U3025, P1_U3026, P1_U3027, P1_U3028, P1_U3029, P1_U3030, P1_U3031, P1_U3032, P1_U3033, P1_U3034, P1_U3035, P1_U3036, P1_U3037, P1_U3038, P1_U3039, P1_U3040, P1_U3041, P1_U3042, P1_U3043, P1_U3044, P1_U3045, P1_U3046, P1_U3047, P1_U3048, P1_U3049, P1_U3050, P1_U3051, P1_U3052, P1_U3053, P1_U3054, P1_U3055, P1_U3056, P1_U3057, P1_U3058, P1_U3059, P1_U3060, P1_U3061, P1_U3062, P1_U3063, P1_U3064, P1_U3065, P1_U3066, P1_U3067, P1_U3068, P1_U3069, P1_U3070, P1_U3071, P1_U3072, P1_U3073, P1_U3074, P1_U3075, P1_U3076, P1_U3077, P1_U3078, P1_U3079, P1_U3080, P1_U3081, P1_U3082, P1_U3083, P1_U3084, P1_U3087, P1_U3088, P1_U3089, P1_U3090, P1_U3091, P1_U3092, P1_U3093, P1_U3094, P1_U3095, P1_U3096, P1_U3097, P1_U3098, P1_U3099, P1_U3100, P1_U3101, P1_U3102, P1_U3103, P1_U3104, P1_U3105, P1_U3106, P1_U3107, P1_U3108, P1_U3109, P1_U3110, P1_U3111, P1_U3112, P1_U3113, P1_U3114, P1_U3115, P1_U3116, P1_U3117, P1_U3118, P1_U3119, P1_U3120, P1_U3121, P1_U3122, P1_U3123, P1_U3124, P1_U3125, P1_U3126, P1_U3127, P1_U3128, P1_U3129, P1_U3130, P1_U3131, P1_U3132, P1_U3133, P1_U3134, P1_U3135, P1_U3136, P1_U3137, P1_U3138, P1_U3139, P1_U3140, P1_U3141, P1_U3142, P1_U3143, P1_U3144, P1_U3145, P1_U3146, P1_U3147, P1_U3148, P1_U3149, P1_U3150, P1_U3151, P1_U3152, P1_U3153, P1_U3154, P1_U3155, P1_U3156, P1_U3157, P1_U3158, P1_U3159, P1_U3160, P1_U3161, P1_U3162, P1_U3163, P1_U3164, P1_U3165, P1_U3166, P1_U3167, P1_U3168, P1_U3169, P1_U3170, P1_U3171, P1_U3172, P1_U3173, P1_U3174, P1_U3175, P1_U3176, P1_U3177, P1_U3178, P1_U3179, P1_U3180, P1_U3181, P1_U3182, P1_U3183, P1_U3184, P1_U3185, P1_U3186, P1_U3187, P1_U3188, P1_U3189, P1_U3190, P1_U3191, P1_U3192, P1_U3193, P1_U3194, P1_U3195, P1_U3196, P1_U3197, P1_U3198, P1_U3199, P1_U3200, P1_U3201, P1_U3202, P1_U3203, P1_U3204, P1_U3205, P1_U3206, P1_U3207, P1_U3208, P1_U3209, P1_U3210, P1_U3211, P1_U3212, P1_U3357, P1_U3358, P1_U3359, P1_U3360, P1_U3361, P1_U3362, P1_U3363, P1_U3364, P1_U3365, P1_U3366, P1_U3367, P1_U3368, P1_U3369, P1_U3370, P1_U3371, P1_U3372, P1_U3373, P1_U3374, P1_U3375, P1_U3376, P1_U3377, P1_U3378, P1_U3379, P1_U3380, P1_U3381, P1_U3382, P1_U3383, P1_U3384, P1_U3385, P1_U3386, P1_U3387, P1_U3388, P1_U3389, P1_U3390, P1_U3391, P1_U3392, P1_U3393, P1_U3394, P1_U3395, P1_U3396, P1_U3397, P1_U3398, P1_U3399, P1_U3400, P1_U3401, P1_U3402, P1_U3403, P1_U3404, P1_U3405, P1_U3406, P1_U3407, P1_U3408, P1_U3409, P1_U3410, P1_U3411, P1_U3412, P1_U3413, P1_U3414, P1_U3415, P1_U3416, P1_U3417, P1_U3418, P1_U3419, P1_U3420, P1_U3421, P1_U3422, P1_U3423, P1_U3424, P1_U3425, P1_U3426, P1_U3427, P1_U3428, P1_U3429, P1_U3430, P1_U3431, P1_U3432, P1_U3433, P1_U3434, P1_U3435, P1_U3436, P1_U3437, P1_U3438, P1_U3439, P1_U3440, P1_U3441, P1_U3442, P1_U3443, P1_U3444, P1_U3447, P1_U3448, P1_U3449, P1_U3450, P1_U3451, P1_U3452, P1_U3453, P1_U3454, P1_U3455, P1_U3456, P1_U3457, P1_U3458, P1_U3460, P1_U3461, P1_U3463, P1_U3464, P1_U3466, P1_U3467, P1_U3469, P1_U3470, P1_U3472, P1_U3473, P1_U3475, P1_U3476, P1_U3478, P1_U3479, P1_U3481, P1_U3482, P1_U3484, P1_U3485, P1_U3487, P1_U3488, P1_U3490, P1_U3491, P1_U3493, P1_U3494, P1_U3496, P1_U3497, P1_U3499, P1_U3500, P1_U3502, P1_U3503, P1_U3505, P1_U3506, P1_U3508, P1_U3509, P1_U3511, P1_U3512, P1_U3514, P1_U3592, P1_U3593, P1_U3594, P1_U3595, P1_U3596, P1_U3597, P1_U3598, P1_U3599, P1_U3600, P1_U3601, P1_U3602, P1_U3603, P1_U3604, P1_U3605, P1_U3606, P1_U3607, P1_U3608, P1_U3609, P1_U3610, P1_U3611, P1_U3612, P1_U3613, P1_U3614, P1_U3615, P1_U3616, P1_U3617, P1_U3618, P1_U3619, P1_U3620, P1_U3621, P1_U3622, P1_U3623, P1_U3624, P1_U3625, P1_U3626, P1_U3627, P1_U3628, P1_U3629, P1_U3630, P1_U3631, P1_U3632, P1_U3633, P1_U3634, P1_U3635, P1_U3636, P1_U3637, P1_U3638, P1_U3639, P1_U3640, P1_U3641, P1_U3642, P1_U3643, P1_U3644, P1_U3645, P1_U3646, P1_U3647, P1_U3648, P1_U3649, P1_U3650, P1_U3651, P1_U3652, P1_U3653, P1_U3654, P1_U3655, P1_U3656, P1_U3657, P1_U3658, P1_U3659, P1_U3660, P1_U3661, P1_U3662, P1_U3663, P1_U3664, P1_U3665, P1_U3666, P1_U3667, P1_U3668, P1_U3669, P1_U3670, P1_U3671, P1_U3672, P1_U3673, P1_U3674, P1_U3675, P1_U3676, P1_U3677, P1_U3678, P1_U3679, P1_U3680, P1_U3681, P1_U3682, P1_U3683, P1_U3684, P1_U3685, P1_U3686, P1_U3687, P1_U3688, P1_U3689, P1_U3690, P1_U3691, P1_U3692, P1_U3693, P1_U3694, P1_U3695, P1_U3696, P1_U3697, P1_U3698, P1_U3699, P1_U3700, P1_U3701, P1_U3702, P1_U3703, P1_U3704, P1_U3705, P1_U3706, P1_U3707, P1_U3708, P1_U3709, P1_U3710, P1_U3711, P1_U3712, P1_U3713, P1_U3714, P1_U3715, P1_U3716, P1_U3717, P1_U3718, P1_U3719, P1_U3720, P1_U3721, P1_U3722, P1_U3723, P1_U3724, P1_U3725, P1_U3726, P1_U3727, P1_U3728, P1_U3729, P1_U3730, P1_U3731, P1_U3732, P1_U3733, P1_U3734, P1_U3735, P1_U3736, P1_U3737, P1_U3738, P1_U3739, P1_U3740, P1_U3741, P1_U3742, P1_U3743, P1_U3744, P1_U3745, P1_U3746, P1_U3747, P1_U3748, P1_U3749, P1_U3750, P1_U3751, P1_U3752, P1_U3753, P1_U3754, P1_U3755, P1_U3756, P1_U3757, P1_U3758, P1_U3759, P1_U3760, P1_U3761, P1_U3762, P1_U3763, P1_U3764, P1_U3765, P1_U3766, P1_U3767, P1_U3768, P1_U3769, P1_U3770, P1_U3771, P1_U3772, P1_U3773, P1_U3774, P1_U3775, P1_U3776, P1_U3777, P1_U3778, P1_U3779, P1_U3780, P1_U3781, P1_U3782, P1_U3783, P1_U3784, P1_U3785, P1_U3786, P1_U3787, P1_U3788, P1_U3789, P1_U3790, P1_U3791, P1_U3792, P1_U3793, P1_U3794, P1_U3795, P1_U3796, P1_U3797, P1_U3798, P1_U3799, P1_U3800, P1_U3801, P1_U3802, P1_U3803, P1_U3804, P1_U3805, P1_U3806, P1_U3807, P1_U3808, P1_U3809, P1_U3810, P1_U3811, P1_U3812, P1_U3813, P1_U3814, P1_U3815, P1_U3816, P1_U3817, P1_U3818, P1_U3819, P1_U3820, P1_U3821, P1_U3822, P1_U3823, P1_U3824, P1_U3825, P1_U3826, P1_U3827, P1_U3828, P1_U3829, P1_U3830, P1_U3831, P1_U3832, P1_U3833, P1_U3834, P1_U3835, P1_U3836, P1_U3837, P1_U3838, P1_U3839, P1_U3840, P1_U3841, P1_U3842, P1_U3843, P1_U3844, P1_U3845, P1_U3846, P1_U3847, P1_U3848, P1_U3849, P1_U3850, P1_U3851, P1_U3852, P1_U3853, P1_U3854, P1_U3855, P1_U3856, P1_U3857, P1_U3858, P1_U3859, P1_U3860, P1_U3861, P1_U3862, P1_U3863, P1_U3864, P1_U3865, P1_U3866, P1_U3867, P1_U3868, P1_U3869, P1_U3870, P1_U3871, P1_U3872, P1_U3873, P1_U3874, P1_U3875, P1_U3876, P1_U3877, P1_U3878, P1_U3879, P1_U3880, P1_U3881, P1_U3882, P1_U3883, P1_U3884, P1_U3885, P1_U3886, P1_U3887, P1_U3888, P1_U3889, P1_U3890, P1_U3891, P1_U3892, P1_U3893, P1_U3894, P1_U3895, P1_U3896, P1_U3897, P1_U3898, P1_U3899, P1_U3900, P1_U3901, P1_U3902, P1_U3903, P1_U3904, P1_U3905, P1_U3906, P1_U3907, P1_U3908, P1_U3909, P1_U3910, P1_U3911, P1_U3912, P1_U3913, P1_U3914, P1_U3915, P1_U3916, P1_U3917, P1_U3918, P1_U3919, P1_U3920, P1_U3921, P1_U3922, P1_U3923, P1_U3924, P1_U3925, P1_U3926, P1_U3927, P1_U3928, P1_U3929, P1_U3930, P1_U3931, P1_U3932, P1_U3933, P1_U3934, P1_U3935, P1_U3936, P1_U3937, P1_U3938, P1_U3939, P1_U3940, P1_U3941, P1_U3942, P1_U3943, P1_U3944, P1_U3945, P1_U3946, P1_U3947, P1_U3948, P1_U3949, P1_U3950, P1_U3951, P1_U3952, P1_U3953, P1_U3954, P1_U3955, P1_U3956, P1_U3957, P1_U3958, P1_U3959, P1_U3960, P1_U3961, P1_U3962, P1_U3963, P1_U3964, P1_U3965, P1_U3966, P1_U3967, P1_U3968, P1_U3969, P1_U3970, P1_U3971, P1_U3972, P1_U3973, P1_U3974, P1_U3975, P1_U3976, P1_U3977, P1_U3978, P1_U3979, P1_U3980, P1_U3981, P1_U3982, P1_U3983, P1_U3984, P1_U3985, P1_U3986, P1_U3987, P1_U3988, P1_U3989, P1_U3990, P1_U3991, P1_U3992, P1_U3993, P1_U3994, P1_U3995, P1_U3996, P1_U3997, P1_U3998, P1_U3999, P1_U4000, P1_U4001, P1_U4002, P1_U4003, P1_U4004, P1_U4005, P1_U4006, P1_U4007, P1_U4008, P1_U4009, P1_U4010, P1_U4011, P1_U4012, P1_U4013, P1_U4014, P1_U4015, P1_U4017, P1_U4018, P1_U4019, P1_U4020, P1_U4021, P1_U4022, P1_U4023, P1_U4024, P1_U4025, P1_U4026, P1_U4027, P1_U4028, P1_U4029, P1_U4030, P1_U4031, P1_U4032, P1_U4033, P1_U4034, P1_U4035, P1_U4036, P1_U4037, P1_U4038, P1_U4039, P1_U4040, P1_U4041, P1_U4042, P1_U4043, P1_U4044, P1_U4045, P1_U4046, P1_U4047, P1_U4048, P1_U4049, P1_U4050, P1_U4051, P1_U4052, P1_U4053, P1_U4054, P1_U4055, P1_U4056, P1_U4057, P1_U4058, P1_U4059, P1_U4060, P1_U4061, P1_U4062, P1_U4063, P1_U4064, P1_U4065, P1_U4066, P1_U4067, P1_U4068, P1_U4069, P1_U4070, P1_U4071, P1_U4072, P1_U4073, P1_U4074, P1_U4075, P1_U4076, P1_U4077, P1_U4078, P1_U4079, P1_U4080, P1_U4081, P1_U4082, P1_U4083, P1_U4084, P1_U4085, P1_U4086, P1_U4087, P1_U4088, P1_U4089, P1_U4090, P1_U4091, P1_U4092, P1_U4093, P1_U4094, P1_U4095, P1_U4096, P1_U4097, P1_U4098, P1_U4099, P1_U4100, P1_U4101, P1_U4102, P1_U4103, P1_U4104, P1_U4105, P1_U4106, P1_U4107, P1_U4108, P1_U4109, P1_U4110, P1_U4111, P1_U4112, P1_U4113, P1_U4114, P1_U4115, P1_U4116, P1_U4117, P1_U4118, P1_U4119, P1_U4120, P1_U4121, P1_U4122, P1_U4123, P1_U4124, P1_U4125, P1_U4126, P1_U4127, P1_U4128, P1_U4129, P1_U4130, P1_U4131, P1_U4132, P1_U4133, P1_U4134, P1_U4135, P1_U4136, P1_U4137, P1_U4138, P1_U4139, P1_U4140, P1_U4141, P1_U4142, P1_U4143, P1_U4144, P1_U4145, P1_U4146, P1_U4147, P1_U4148, P1_U4149, P1_U4150, P1_U4151, P1_U4152, P1_U4153, P1_U4154, P1_U4155, P1_U4156, P1_U4157, P1_U4158, P1_U4159, P1_U4160, P1_U4161, P1_U4162, P1_U4163, P1_U4164, P1_U4165, P1_U4166, P1_U4167, P1_U4168, P1_U4169, P1_U4170, P1_U4171, P1_U4172, P1_U4173, P1_U4174, P1_U4175, P1_U4176, P1_U4177, P1_U4178, P1_U4179, P1_U4180, P1_U4181, P1_U4182, P1_U4183, P1_U4184, P1_U4185, P1_U4186, P1_U4187, P1_U4188, P1_U4189, P1_U4190, P1_U4191, P1_U4192, P1_U4193, P1_U4194, P1_U4195, P1_U4196, P1_U4197, P1_U4198, P1_U4199, P1_U4200, P1_U4201, P1_U4202, P1_U4203, P1_U4204, P1_U4205, P1_U4206, P1_U4207, P1_U4208, P1_U4209, P1_U4210, P1_U4211, P1_U4212, P1_U4213, P1_U4214, P1_U4215, P1_U4216, P1_U4217, P1_U4218, P1_U4219, P1_U4220, P1_U4221, P1_U4222, P1_U4223, P1_U4224, P1_U4225, P1_U4226, P1_U4227, P1_U4228, P1_U4229, P1_U4230, P1_U4231, P1_U4232, P1_U4233, P1_U4234, P1_U4235, P1_U4236, P1_U4237, P1_U4238, P1_U4239, P1_U4240, P1_U4241, P1_U4242, P1_U4243, P1_U4244, P1_U4245, P1_U4246, P1_U4247, P1_U4248, P1_U4249, P1_U4250, P1_U4251, P1_U4252, P1_U4253, P1_U4254, P1_U4255, P1_U4256, P1_U4257, P1_U4258, P1_U4259, P1_U4260, P1_U4261, P1_U4262, P1_U4263, P1_U4264, P1_U4265, P1_U4266, P1_U4267, P1_U4268, P1_U4269, P1_U4270, P1_U4271, P1_U4272, P1_U4273, P1_U4274, P1_U4275, P1_U4276, P1_U4277, P1_U4278, P1_U4279, P1_U4280, P1_U4281, P1_U4282, P1_U4283, P1_U4284, P1_U4285, P1_U4286, P1_U4287, P1_U4288, P1_U4289, P1_U4290, P1_U4291, P1_U4292, P1_U4293, P1_U4294, P1_U4295, P1_U4296, P1_U4297, P1_U4298, P1_U4299, P1_U4300, P1_U4301, P1_U4302, P1_U4303, P1_U4304, P1_U4305, P1_U4306, P1_U4307, P1_U4308, P1_U4309, P1_U4310, P1_U4311, P1_U4312, P1_U4313, P1_U4314, P1_U4315, P1_U4316, P1_U4317, P1_U4318, P1_U4319, P1_U4320, P1_U4321, P1_U4322, P1_U4323, P1_U4324, P1_U4325, P1_U4326, P1_U4327, P1_U4328, P1_U4329, P1_U4330, P1_U4331, P1_U4332, P1_U4333, P1_U4334, P1_U4335, P1_U4336, P1_U4337, P1_U4338, P1_U4339, P1_U4340, P1_U4341, P1_U4342, P1_U4343, P1_U4344, P1_U4345, P1_U4346, P1_U4347, P1_U4348, P1_U4349, P1_U4350, P1_U4351, P1_U4352, P1_U4353, P1_U4354, P1_U4355, P1_U4356, P1_U4357, P1_U4358, P1_U4359, P1_U4360, P1_U4361, P1_U4362, P1_U4363, P1_U4364, P1_U4365, P1_U4366, P1_U4367, P1_U4368, P1_U4369, P1_U4370, P1_U4371, P1_U4372, P1_U4373, P1_U4374, P1_U4375, P1_U4376, P1_U4377, P1_U4378, P1_U4379, P1_U4380, P1_U4381, P1_U4382, P1_U4383, P1_U4384, P1_U4385, P1_U4386, P1_U4387, P1_U4388, P1_U4389, P1_U4390, P1_U4391, P1_U4392, P1_U4393, P1_U4394, P1_U4395, P1_U4396, P1_U4397, P1_U4398, P1_U4399, P1_U4400, P1_U4401, P1_U4402, P1_U4403, P1_U4404, P1_U4405, P1_U4406, P1_U4407, P1_U4408, P1_U4409, P1_U4410, P1_U4411, P1_U4412, P1_U4413, P1_U4414, P1_U4415, P1_U4416, P1_U4417, P1_U4418, P1_U4419, P1_U4420, P1_U4421, P1_U4422, P1_U4423, P1_U4424, P1_U4425, P1_U4426, P1_U4427, P1_U4428, P1_U4429, P1_U4430, P1_U4431, P1_U4432, P1_U4433, P1_U4434, P1_U4435, P1_U4436, P1_U4437, P1_U4438, P1_U4439, P1_U4440, P1_U4441, P1_U4442, P1_U4443, P1_U4444, P1_U4445, P1_U4446, P1_U4447, P1_U4448, P1_U4449, P1_U4450, P1_U4451, P1_U4452, P1_U4453, P1_U4454, P1_U4455, P1_U4456, P1_U4457, P1_U4458, P1_U4459, P1_U4460, P1_U4461, P1_U4462, P1_U4463, P1_U4464, P1_U4465, P1_U4466, P1_U4467, P1_U4468, P1_U4469, P1_U4470, P1_U4471, P1_U4472, P1_U4473, P1_U4474, P1_U4475, P1_U4476, P1_U4477, P1_U4478, P1_U4479, P1_U4480, P1_U4481, P1_U4482, P1_U4483, P1_U4484, P1_U4485, P1_U4486, P1_U4487, P1_U4488, P1_U4489, P1_U4490, P1_U4491, P1_U4492, P1_U4493, P1_U4494, P1_U4495, P1_U4496, P1_U4497, P1_U4498, P1_U4499, P1_U4500, P1_U4501, P1_U4502, P1_U4503, P1_U4504, P1_U4505, P1_U4506, P1_U4507, P1_U4508, P1_U4509, P1_U4510, P1_U4511, P1_U4512, P1_U4513, P1_U4514, P1_U4515, P1_U4516, P1_U4517, P1_U4518, P1_U4519, P1_U4520, P1_U4521, P1_U4522, P1_U4523, P1_U4524, P1_U4525, P1_U4526, P1_U4527, P1_U4528, P1_U4529, P1_U4530, P1_U4531, P1_U4532, P1_U4533, P1_U4534, P1_U4535, P1_U4536, P1_U4537, P1_U4538, P1_U4539, P1_U4540, P1_U4541, P1_U4542, P1_U4543, P1_U4544, P1_U4545, P1_U4546, P1_U4547, P1_U4548, P1_U4549, P1_U4550, P1_U4551, P1_U4552, P1_U4553, P1_U4554, P1_U4555, P1_U4556, P1_U4557, P1_U4558, P1_U4559, P1_U4560, P1_U4561, P1_U4562, P1_U4563, P1_U4564, P1_U4565, P1_U4566, P1_U4567, P1_U4568, P1_U4569, P1_U4570, P1_U4571, P1_U4572, P1_U4573, P1_U4574, P1_U4575, P1_U4576, P1_U4577, P1_U4578, P1_U4579, P1_U4580, P1_U4581, P1_U4582, P1_U4583, P1_U4584, P1_U4585, P1_U4586, P1_U4587, P1_U4588, P1_U4589, P1_U4590, P1_U4591, P1_U4592, P1_U4593, P1_U4594, P1_U4595, P1_U4596, P1_U4597, P1_U4598, P1_U4599, P1_U4600, P1_U4601, P1_U4602, P1_U4603, P1_U4604, P1_U4605, P1_U4606, P1_U4607, P1_U4608, P1_U4609, P1_U4610, P1_U4611, P1_U4612, P1_U4613, P1_U4614, P1_U4615, P1_U4616, P1_U4617, P1_U4618, P1_U4619, P1_U4620, P1_U4621, P1_U4622, P1_U4623, P1_U4624, P1_U4625, P1_U4626, P1_U4627, P1_U4628, P1_U4629, P1_U4630, P1_U4631, P1_U4632, P1_U4633, P1_U4634, P1_U4635, P1_U4636, P1_U4637, P1_U4638, P1_U4639, P1_U4640, P1_U4641, P1_U4642, P1_U4643, P1_U4644, P1_U4645, P1_U4646, P1_U4647, P1_U4648, P1_U4649, P1_U4650, P1_U4651, P1_U4652, P1_U4653, P1_U4654, P1_U4655, P1_U4656, P1_U4657, P1_U4658, P1_U4659, P1_U4660, P1_U4661, P1_U4662, P1_U4663, P1_U4664, P1_U4665, P1_U4666, P1_U4667, P1_U4668, P1_U4669, P1_U4670, P1_U4671, P1_U4672, P1_U4673, P1_U4674, P1_U4675, P1_U4676, P1_U4677, P1_U4678, P1_U4679, P1_U4680, P1_U4681, P1_U4682, P1_U4683, P1_U4684, P1_U4685, P1_U4686, P1_U4687, P1_U4688, P1_U4689, P1_U4690, P1_U4691, P1_U4692, P1_U4693, P1_U4694, P1_U4695, P1_U4696, P1_U4697, P1_U4698, P1_U4699, P1_U4700, P1_U4701, P1_U4702, P1_U4703, P1_U4704, P1_U4705, P1_U4706, P1_U4707, P1_U4708, P1_U4709, P1_U4710, P1_U4711, P1_U4712, P1_U4713, P1_U4714, P1_U4715, P1_U4716, P1_U4717, P1_U4718, P1_U4719, P1_U4720, P1_U4721, P1_U4722, P1_U4723, P1_U4724, P1_U4725, P1_U4726, P1_U4727, P1_U4728, P1_U4729, P1_U4730, P1_U4731, P1_U4732, P1_U4733, P1_U4734, P1_U4735, P1_U4736, P1_U4737, P1_U4738, P1_U4739, P1_U4740, P1_U4741, P1_U4742, P1_U4743, P1_U4744, P1_U4745, P1_U4746, P1_U4747, P1_U4748, P1_U4749, P1_U4750, P1_U4751, P1_U4752, P1_U4753, P1_U4754, P1_U4755, P1_U4756, P1_U4757, P1_U4758, P1_U4759, P1_U4760, P1_U4761, P1_U4762, P1_U4763, P1_U4764, P1_U4765, P1_U4766, P1_U4767, P1_U4768, P1_U4769, P1_U4770, P1_U4771, P1_U4772, P1_U4773, P1_U4774, P1_U4775, P1_U4776, P1_U4777, P1_U4778, P1_U4779, P1_U4780, P1_U4781, P1_U4782, P1_U4783, P1_U4784, P1_U4785, P1_U4786, P1_U4787, P1_U4788, P1_U4789, P1_U4790, P1_U4791, P1_U4792, P1_U4793, P1_U4794, P1_U4795, P1_U4796, P1_U4797, P1_U4798, P1_U4799, P1_U4800, P1_U4801, P1_U4802, P1_U4803, P1_U4804, P1_U4805, P1_U4806, P1_U4807, P1_U4808, P1_U4809, P1_U4810, P1_U4811, P1_U4812, P1_U4813, P1_U4814, P1_U4815, P1_U4816, P1_U4817, P1_U4818, P1_U4819, P1_U4820, P1_U4821, P1_U4822, P1_U4823, P1_U4824, P1_U4825, P1_U4826, P1_U4827, P1_U4828, P1_U4829, P1_U4830, P1_U4831, P1_U4832, P1_U4833, P1_U4834, P1_U4835, P1_U4836, P1_U4837, P1_U4838, P1_U4839, P1_U4840, P1_U4841, P1_U4842, P1_U4843, P1_U4844, P1_U4845, P1_U4846, P1_U4847, P1_U4848, P1_U4849, P1_U4850, P1_U4851, P1_U4852, P1_U4853, P1_U4854, P1_U4855, P1_U4856, P1_U4857, P1_U4858, P1_U4859, P1_U4860, P1_U4861, P1_U4862, P1_U4863, P1_U4864, P1_U4865, P1_U4866, P1_U4867, P1_U4868, P1_U4869, P1_U4870, P1_U4871, P1_U4872, P1_U4873, P1_U4874, P1_U4875, P1_U4876, P1_U4877, P1_U4878, P1_U4879, P1_U4880, P1_U4881, P1_U4882, P1_U4883, P1_U4884, P1_U4885, P1_U4886, P1_U4887, P1_U4888, P1_U4889, P1_U4890, P1_U4891, P1_U4892, P1_U4893, P1_U4894, P1_U4895, P1_U4896, P1_U4897, P1_U4898, P1_U4899, P1_U4900, P1_U4901, P1_U4902, P1_U4903, P1_U4904, P1_U4905, P1_U4906, P1_U4907, P1_U4908, P1_U4909, P1_U4910, P1_U4911, P1_U4912, P1_U4913, P1_U4914, P1_U4915, P1_U4916, P1_U4917, P1_U4918, P1_U4919, P1_U4920, P1_U4921, P1_U4922, P1_U4923, P1_U4924, P1_U4925, P1_U4926, P1_U4927, P1_U4928, P1_U4929, P1_U4930, P1_U4931, P1_U4932, P1_U4933, P1_U4934, P1_U4935, P1_U4936, P1_U4937, P1_U4938, P1_U4939, P1_U4940, P1_U4941, P1_U4942, P1_U4943, P1_U4944, P1_U4945, P1_U4946, P1_U4947, P1_U4948, P1_U4949, P1_U4950, P1_U4951, P1_U4952, P1_U4953, P1_U4954, P1_U4955, P1_U4956, P1_U4957, P1_U4958, P1_U4959, P1_U4960, P1_U4961, P1_U4962, P1_U4963, P1_U4964, P1_U4965, P1_U4966, P1_U4967, P1_U4968, P1_U4969, P1_U4970, P1_U4971, P1_U4972, P1_U4973, P1_U4974, P1_U4975, P1_U4976, P1_U4977, P1_U4978, P1_U4979, P1_U4980, P1_U4981, P1_U4982, P1_U4983, P1_U4984, P1_U4985, P1_U4986, P1_U4987, P1_U4988, P1_U4989, P1_U4990, P1_U4991, P1_U4992, P1_U4993, P1_U4994, P1_U4995, P1_U4996, P1_U4997, P1_U4998, P1_U4999, P1_U5000, P1_U5001, P1_U5002, P1_U5003, P1_U5004, P1_U5005, P1_U5006, P1_U5007, P1_U5008, P1_U5009, P1_U5010, P1_U5011, P1_U5012, P1_U5013, P1_U5014, P1_U5015, P1_U5016, P1_U5017, P1_U5018, P1_U5019, P1_U5020, P1_U5021, P1_U5022, P1_U5023, P1_U5024, P1_U5025, P1_U5026, P1_U5027, P1_U5028, P1_U5029, P1_U5030, P1_U5031, P1_U5032, P1_U5033, P1_U5034, P1_U5035, P1_U5036, P1_U5037, P1_U5038, P1_U5039, P1_U5040, P1_U5041, P1_U5042, P1_U5043, P1_U5044, P1_U5045, P1_U5046, P1_U5047, P1_U5048, P1_U5049, P1_U5050, P1_U5051, P1_U5052, P1_U5053, P1_U5054, P1_U5055, P1_U5056, P1_U5057, P1_U5058, P1_U5059, P1_U5060, P1_U5061, P1_U5062, P1_U5063, P1_U5064, P1_U5065, P1_U5066, P1_U5067, P1_U5068, P1_U5069, P1_U5070, P1_U5071, P1_U5072, P1_U5073, P1_U5074, P1_U5075, P1_U5076, P1_U5077, P1_U5078, P1_U5079, P1_U5080, P1_U5081, P1_U5082, P1_U5083, P1_U5084, P1_U5085, P1_U5086, P1_U5087, P1_U5088, P1_U5089, P1_U5090, P1_U5091, P1_U5092, P1_U5093, P1_U5094, P1_U5095, P1_U5096, P1_U5097, P1_U5098, P1_U5099, P1_U5100, P1_U5101, P1_U5102, P1_U5103, P1_U5104, P1_U5105, P1_U5106, P1_U5107, P1_U5108, P1_U5109, P1_U5110, P1_U5111, P1_U5112, P1_U5113, P1_U5114, P1_U5115, P1_U5116, P1_U5117, P1_U5118, P1_U5119, P1_U5120, P1_U5121, P1_U5122, P1_U5123, P1_U5124, P1_U5125, P1_U5126, P1_U5127, P1_U5128, P1_U5129, P1_U5130, P1_U5131, P1_U5132, P1_U5133, P1_U5134, P1_U5135, P1_U5136, P1_U5137, P1_U5138, P1_U5139, P1_U5140, P1_U5141, P1_U5142, P1_U5143, P1_U5144, P1_U5145, P1_U5146, P1_U5147, P1_U5148, P1_U5149, P1_U5150, P1_U5151, P1_U5152, P1_U5153, P1_U5154, P1_U5155, P1_U5156, P1_U5157, P1_U5158, P1_U5159, P1_U5160, P1_U5161, P1_U5162, P1_U5163, P1_U5164, P1_U5165, P1_U5166, P1_U5167, P1_U5168, P1_U5169, P1_U5170, P1_U5171, P1_U5172, P1_U5173, P1_U5174, P1_U5175, P1_U5176, P1_U5177, P1_U5178, P1_U5179, P1_U5180, P1_U5181, P1_U5182, P1_U5183, P1_U5184, P1_U5185, P1_U5186, P1_U5187, P1_U5188, P1_U5189, P1_U5190, P1_U5191, P1_U5192, P1_U5193, P1_U5194, P1_U5195, P1_U5196, P1_U5197, P1_U5198, P1_U5199, P1_U5200, P1_U5201, P1_U5202, P1_U5203, P1_U5204, P1_U5205, P1_U5206, P1_U5207, P1_U5208, P1_U5209, P1_U5210, P1_U5211, P1_U5212, P1_U5213, P1_U5214, P1_U5215, P1_U5216, P1_U5217, P1_U5218, P1_U5219, P1_U5220, P1_U5221, P1_U5222, P1_U5223, P1_U5224, P1_U5225, P1_U5226, P1_U5227, P1_U5228, P1_U5229, P1_U5230, P1_U5231, P1_U5232, P1_U5233, P1_U5234, P1_U5235, P1_U5236, P1_U5237, P1_U5238, P1_U5239, P1_U5240, P1_U5241, P1_U5242, P1_U5243, P1_U5244, P1_U5245, P1_U5246, P1_U5247, P1_U5248, P1_U5249, P1_U5250, P1_U5251, P1_U5252, P1_U5253, P1_U5254, P1_U5255, P1_U5256, P1_U5257, P1_U5258, P1_U5259, P1_U5260, P1_U5261, P1_U5262, P1_U5263, P1_U5264, P1_U5265, P1_U5266, P1_U5267, P1_U5268, P1_U5269, P1_U5270, P1_U5271, P1_U5272, P1_U5273, P1_U5274, P1_U5275, P1_U5276, P1_U5277, P1_U5278, P1_U5279, P1_U5280, P1_U5281, P1_U5282, P1_U5283, P1_U5284, P1_U5285, P1_U5286, P1_U5287, P1_U5288, P1_U5289, P1_U5290, P1_U5291, P1_U5292, P1_U5293, P1_U5294, P1_U5295, P1_U5296, P1_U5297, P1_U5298, P1_U5299, P1_U5300, P1_U5301, P1_U5302, P1_U5303, P1_U5304, P1_U5305, P1_U5306, P1_U5307, P1_U5308, P1_U5309, P1_U5310, P1_U5311, P1_U5312, P1_U5313, P1_U5314, P1_U5315, P1_U5316, P1_U5317, P1_U5318, P1_U5319, P1_U5320, P1_U5321, P1_U5322, P1_U5323, P1_U5324, P1_U5325, P1_U5326, P1_U5327, P1_U5328, P1_U5329, P1_U5330, P1_U5331, P1_U5332, P1_U5333, P1_U5334, P1_U5335, P1_U5336, P1_U5337, P1_U5338, P1_U5339, P1_U5340, P1_U5341, P1_U5342, P1_U5343, P1_U5344, P1_U5345, P1_U5346, P1_U5347, P1_U5348, P1_U5349, P1_U5350, P1_U5351, P1_U5352, P1_U5353, P1_U5354, P1_U5355, P1_U5356, P1_U5357, P1_U5358, P1_U5359, P1_U5360, P1_U5361, P1_U5362, P1_U5363, P1_U5364, P1_U5365, P1_U5366, P1_U5367, P1_U5368, P1_U5369, P1_U5370, P1_U5371, P1_U5372, P1_U5373, P1_U5374, P1_U5375, P1_U5376, P1_U5377, P1_U5378, P1_U5379, P1_U5380, P1_U5381, P1_U5382, P1_U5383, P1_U5384, P1_U5385, P1_U5386, P1_U5387, P1_U5388, P1_U5389, P1_U5390, P1_U5391, P1_U5392, P1_U5393, P1_U5394, P1_U5395, P1_U5396, P1_U5397, P1_U5398, P1_U5399, P1_U5400, P1_U5401, P1_U5402, P1_U5403, P1_U5404, P1_U5405, P1_U5406, P1_U5407, P1_U5408, P1_U5409, P1_U5410, P1_U5411, P1_U5412, P1_U5413, P1_U5414, P1_U5415, P1_U5416, P1_U5417, P1_U5418, P1_U5419, P1_U5420, P1_U5421, P1_U5422, P1_U5423, P1_U5424, P1_U5425, P1_U5426, P1_U5427, P1_U5428, P1_U5429, P1_U5430, P1_U5431, P1_U5432, P1_U5433, P1_U5434, P1_U5435, P1_U5436, P1_U5437, P1_U5438, P1_U5439, P1_U5440, P1_U5441, P1_U5442, P1_U5443, P1_U5444, P1_U5445, P1_U5446, P1_U5447, P1_U5448, P1_U5449, P1_U5450, P1_U5451, P1_U5452, P1_U5453, P1_U5454, P1_U5455, P1_U5456, P1_U5457, P1_U5458, P1_U5459, P1_U5460, P1_U5461, P1_U5462, P1_U5463, P1_U5464, P1_U5465, P1_U5466, P1_U5467, P1_U5468, P1_U5469, P1_U5470, P1_U5471, P1_U5472, P1_U5473, P1_U5474, P1_U5475, P1_U5476, P1_U5477, P1_U5478, P1_U5479, P1_U5480, P1_U5481, P1_U5482, P1_U5483, P1_U5484, P1_U5485, P1_U5486, P1_U5487, P1_U5488, P1_U5489, P1_U5490, P1_U5491, P1_U5492, P1_U5493, P1_U5494, P1_U5495, P1_U5496, P1_U5497, P1_U5498, P1_U5499, P1_U5500, P1_U5501, P1_U5502, P1_U5503, P1_U5504, P1_U5505, P1_U5506, P1_U5507, P1_U5508, P1_U5509, P1_U5510, P1_U5511, P1_U5512, P1_U5513, P1_U5514, P1_U5515, P1_U5516, P1_U5517, P1_U5518, P1_U5519, P1_U5520, P1_U5521, P1_U5522, P1_U5523, P1_U5524, P1_U5525, P1_U5526, P1_U5527, P1_U5528, P1_U5529, P1_U5530, P1_U5531, P1_U5532, P1_U5533, P1_U5534, P1_U5535, P1_U5536, P1_U5537, P1_U5538, P1_U5539, P1_U5540, P1_U5541, P1_U5542, P1_U5543, P1_U5544, P1_U5545, P1_U5546, P1_U5547, P1_U5548, P1_U5549, P1_U5550, P1_U5551, P1_U5552, P1_U5553, P1_U5554, P1_U5555, P1_U5556, P1_U5557, P1_U5558, P1_U5559, P1_U5560, P1_U5561, P1_U5562, P1_U5563, P1_U5564, P1_U5565, P1_U5566, P1_U5567, P1_U5568, P1_U5569, P1_U5570, P1_U5571, P1_U5572, P1_U5573, P1_U5574, P1_U5575, P1_U5576, P1_U5577, P1_U5578, P1_U5579, P1_U5580, P1_U5581, P1_U5582, P1_U5583, P1_U5584, P1_U5585, P1_U5586, P1_U5587, P1_U5588, P1_U5589, P1_U5590, P1_U5591, P1_U5592, P1_U5593, P1_U5594, P1_U5595, P1_U5596, P1_U5597, P1_U5598, P1_U5599, P1_U5600, P1_U5601, P1_U5602, P1_U5603, P1_U5604, P1_U5605, P1_U5606, P1_U5607, P1_U5608, P1_U5609, P1_U5610, P1_U5611, P1_U5612, P1_U5613, P1_U5614, P1_U5615, P1_U5616, P1_U5617, P1_U5618, P1_U5619, P1_U5620, P1_U5621, P1_U5622, P1_U5623, P1_U5624, P1_U5625, P1_U5626, P1_U5627, P1_U5628, P1_U5629, P1_U5630, P1_U5631, P1_U5632, P1_U5633, P1_U5634, P1_U5635, P1_U5636, P1_U5637, P1_U5638, P1_U5639, P1_U5640, P1_U5641, P1_U5642, P1_U5643, P1_U5644, P1_U5645, P1_U5646, P1_U5647, P1_U5648, P1_U5649, P1_U5650, P1_U5651, P1_U5652, P1_U5653, P1_U5654, P1_U5655, P1_U5656, P1_U5657, P1_U5658, P1_U5659, P1_U5660, P1_U5661, P1_U5662, P1_U5663, P1_U5664, P1_U5665, P1_U5666, P1_U5667, P1_U5668, P1_U5669, P1_U5670, P1_U5671, P1_U5672, P1_U5673, P1_U5674, P1_U5675, P1_U5676, P1_U5677, P1_U5678, P1_U5679, P1_U5680, P1_U5681, P1_U5682, P1_U5683, P1_U5684, P1_U5685, P1_U5686, P1_U5687, P1_U5688, P1_U5689, P1_U5690, P1_U5691, P1_U5692, P1_U5693, P1_U5694, P1_U5695, P1_U5696, P1_U5697, P1_U5698, P1_U5699, P1_U5700, P1_U5701, P1_U5702, P1_U5703, P1_U5704, P1_U5705, P1_U5706, P1_U5707, P1_U5708, P1_U5709, P1_U5710, P1_U5711, P1_U5712, P1_U5713, P1_U5714, P1_U5715, P1_U5716, P1_U5717, P1_U5718, P1_U5719, P1_U5720, P1_U5721, P1_U5722, P1_U5723, P1_U5724, P1_U5725, P1_U5726, P1_U5727, P1_U5728, P1_U5729, P1_U5730, P1_U5731, P1_U5732, P1_U5733, P1_U5734, P1_U5735, P1_U5736, P1_U5737, P1_U5738, P1_U5739, P1_U5740, P1_U5741, P1_U5742, P1_U5743, P1_U5744, P1_U5745, P1_U5746, P1_U5747, P1_U5748, P1_U5749, P1_U5750, P1_U5751, P1_U5752, P1_U5753, P1_U5754, P1_U5755, P1_U5756, P1_U5757, P1_U5758, P1_U5759, P1_U5760, P1_U5761, P1_U5762, P1_U5763, P1_U5764, P1_U5765, P1_U5766, P1_U5767, P1_U5768, P1_U5769, P1_U5770, P1_U5771, P1_U5772, P1_U5773, P1_U5774, P1_U5775, P1_U5776, P1_U5777, P1_U5778, P1_U5779, P1_U5780, P1_U5781, P1_U5782, P1_U5783, P1_U5784, P1_U5785, P1_U5786, P1_U5787, P1_U5788, P1_U5789, P1_U5790, P1_U5791, P1_U5792, P1_U5793, P1_U5794, P1_U5795, P1_U5796, P1_U5797, P1_U5798, P1_U5799, P1_U5800, P1_U5801, P1_U5802, P1_U5803, P1_U5804, P1_U5805, P1_U5806, P1_U5807, P1_U5808, P1_U5809, P1_U5810, P1_U5811, P1_U5812, P1_U5813, P1_U5814, P1_U5815, P1_U5816, P1_U5817, P1_U5818, P1_U5819, P1_U5820, P1_U5821, P1_U5822, P1_U5823, P1_U5824, P1_U5825, P1_U5826, P1_U5827, P1_U5828, P1_U5829, P1_U5830, P1_U5831, P1_U5832, P1_U5833, P1_U5834, P1_U5835, P1_U5836, P1_U5837, P1_U5838, P1_U5839, P1_U5840, P1_U5841, P1_U5842, P1_U5843, P1_U5844, P1_U5845, P1_U5846, P1_U5847, P1_U5848, P1_U5849, P1_U5850, P1_U5851, P1_U5852, P1_U5853, P1_U5854, P1_U5855, P1_U5856, P1_U5857, P1_U5858, P1_U5859, P1_U5860, P1_U5861, P1_U5862, P1_U5863, P1_U5864, P1_U5865, P1_U5866, P1_U5867, P1_U5868, P1_U5869, P1_U5870, P1_U5871, P1_U5872, P1_U5873, P1_U5874, P1_U5875, P1_U5876, P1_U5877, P1_U5878, P1_U5879, P1_U5880, P1_U5881, P1_U5882, P1_U5883, P1_U5884, P1_U5885, P1_U5886, P1_U5887, P1_U5888, P1_U5889, P1_U5890, P1_U5891, P1_U5892, P1_U5893, P1_U5894, P1_U5895, P1_U5896, P1_U5897, P1_U5898, P1_U5899, P1_U5900, P1_U5901, P1_U5902, P1_U5903, P1_U5904, P1_U5905, P1_U5906, P1_U5907, P1_U5908, P1_U5909, P1_U5910, P1_U5911, P1_U5912, P1_U5913, P1_U5914, P1_U5915, P1_U5916, P1_U5917, P1_U5918, P1_U5919, P1_U5920, P1_U5921, P1_U5922, P1_U5923, P1_U5924, P1_U5925, P1_U5926, P1_U5927, P1_U5928, P1_U5929, P1_U5930, P1_U5931, P1_U5932, P1_U5933, P1_U5934, P1_U5935, P1_U5936, P1_U5937, P1_U5938, P1_U5939, P1_U5940, P1_U5941, P1_U5942, P1_U5943, P1_U5944, P1_U5945, P1_U5946, P1_U5947, P1_U5948, P1_U5949, P1_U5950, P1_U5951, P1_U5952, P1_U5953, P1_U5954, P1_U5955, P1_U5956, P1_U5957, P1_U5958, P1_U5959, P1_U5960, P1_U5961, P1_U5962, P1_U5963, P1_U5964, P1_U5965, P1_U5966, P1_U5967, P1_U5968, P1_U5969, P1_U5970, P1_U5971, P1_U5972, P1_U5973, P1_U5974, P1_U5975, P1_U5976, P1_U5977, P1_U5978, P1_U5979, P1_U5980, P1_U5981, P1_U5982, P1_U5983, P1_U5984, P1_U5985, P1_U5986, P1_U5987, P1_U5988, P1_U5989, P1_U5990, P1_U5991, P1_U5992, P1_U5993, P1_U5994, P1_U5995, P1_U5996, P1_U5997, P1_U5998, P1_U5999, P1_U6000, P1_U6001, P1_U6002, P1_U6003, P1_U6004, P1_U6005, P1_U6006, P1_U6007, P1_U6008, P1_U6009, P1_U6010, P1_U6011, P1_U6012, P1_U6013, P1_U6014, P1_U6015, P1_U6016, P1_U6017, P1_U6018, P1_U6019, P1_U6020, P1_U6021, P1_U6022, P1_U6023, P1_U6024, P1_U6025, P1_U6026, P1_U6027, P1_U6028, P1_U6029, P1_U6030, P1_U6031, P1_U6032, P1_U6033, P1_U6034, P1_U6035, P1_U6036, P1_U6037, P1_U6038, P1_U6039, P1_U6040, P1_U6041, P1_U6042, P1_U6043, P1_U6044, P1_U6045, P1_U6046, P1_U6047, P1_U6048, P1_U6049, P1_U6050, P1_U6051, P1_U6052, P1_U6053, P1_U6054, P1_U6055, P1_U6056, P1_U6057, P1_U6058, P1_U6059, P1_U6060, P1_U6061, P1_U6062, P1_U6063, P1_U6064, P1_U6065, P1_U6066, P1_U6067, P1_U6068, P1_U6069, P1_U6070, P1_U6071, P1_U6072, P1_U6073, P1_U6074, P1_U6075, P1_U6076, P1_U6077, P1_U6078, P1_U6079, P1_U6080, P1_U6081, P1_U6082, P1_U6083, P1_U6084, P1_U6085, P1_U6086, P1_U6087, P1_U6088, P1_U6089, P1_U6090, P1_U6091, P1_U6092, P1_U6093, P1_U6094, P1_U6095, P1_U6096, P1_U6097, P1_U6098, P1_U6099, P1_U6100, P1_U6101, P1_U6102, P1_U6103, P1_U6104, P1_U6105, P1_U6106, P1_U6107, P1_U6108, P1_U6109, P1_U6110, P1_U6111, P1_U6112, P1_U6113, P1_U6114, P1_U6115, P1_U6116, P1_U6117, P1_U6118, P1_U6119, P1_U6120, P1_U6121, P1_U6122, P1_U6123, P1_U6124, P1_U6125, P1_U6126, P1_U6127, P1_U6128, P1_U6129, P1_U6130, P1_U6131, P1_U6132, P1_U6133, P1_U6134, P1_U6135, P1_U6136, P1_U6137, P1_U6138, P1_U6139, P1_U6140, P1_U6141, P1_U6142, P1_U6143, P1_U6144, P1_U6145, P1_U6146, P1_U6147, P1_U6148, P1_U6149, P1_U6150, P1_U6151, P1_U6152, P1_U6153, P1_U6154, P1_U6155, P1_U6156, P1_U6157, P1_U6158, P1_U6159, P1_U6160, P1_U6161, P1_U6162, P1_U6163, P1_U6164, P1_U6165, P1_U6166, P1_U6167, P1_U6168, P1_U6169, P1_U6170, P1_U6171, P1_U6172, P1_U6173, P1_U6174, P1_U6175, P1_U6176, P1_U6177, P1_U6178, P1_U6179, P1_U6180, P1_U6181, P1_U6182, P1_U6183, P1_U6184, P1_U6185, P1_U6186, P1_U6187, P1_U6188, P1_U6189, P1_U6190, P1_U6191, P1_U6192, P1_U6193, P1_U6194, P1_U6195, P1_U6196, P1_U6197, P1_U6198, P1_U6199, P1_U6200, P1_U6201, P1_U6202, P1_U6203, P1_U6204, P1_U6205, P1_U6206, P1_U6207, P1_U6208, P1_U6209, P1_U6210, P1_U6211, P1_U6212, P1_U6213, P1_U6214, P1_U6215, P1_U6216, P1_U6217, P1_U6218, P1_U6219, P1_U6220, P1_U6221, P1_U6222, P1_U6223, P1_U6224, P1_U6225, P1_U6226, P1_U6227, P1_U6228, P1_U6229, P1_U6230, P1_U6231, P1_U6232, P1_U6233, P1_U6234, P1_U6235, P1_U6236, P1_U6237, P1_U6238, P1_U6239, P1_U6240, P1_U6241, P1_U6242, P1_U6243, P1_U6244, P1_U6245, P1_U6246, P1_U6247, P1_U6248, P1_U6249, P1_U6250, P1_U6251, P1_U6252, P1_U6253, P1_U6254, P1_U6255, P1_U6256, P1_U6257, P1_U6258, P1_U6259, P1_U6260, P1_U6261, P1_U6262, P1_U6263, P1_U6264, P1_U6265, P1_U6266, P1_U6267, P1_U6268, P1_U6269, P1_U6270, P1_U6271, P1_U6272, P1_U6273, P1_U6274, P1_U6275, P1_U6276, P1_U6277, P1_U6278, P1_U6279, P1_U6280, P1_U6281, P1_U6282, P1_U6283, P1_U6284, P1_U6285, P2_ADD_1119_U10, P2_ADD_1119_U100, P2_ADD_1119_U101, P2_ADD_1119_U102, P2_ADD_1119_U103, P2_ADD_1119_U104, P2_ADD_1119_U105, P2_ADD_1119_U106, P2_ADD_1119_U107, P2_ADD_1119_U108, P2_ADD_1119_U109, P2_ADD_1119_U11, P2_ADD_1119_U110, P2_ADD_1119_U111, P2_ADD_1119_U112, P2_ADD_1119_U113, P2_ADD_1119_U114, P2_ADD_1119_U115, P2_ADD_1119_U116, P2_ADD_1119_U117, P2_ADD_1119_U118, P2_ADD_1119_U119, P2_ADD_1119_U12, P2_ADD_1119_U120, P2_ADD_1119_U121, P2_ADD_1119_U122, P2_ADD_1119_U123, P2_ADD_1119_U124, P2_ADD_1119_U125, P2_ADD_1119_U126, P2_ADD_1119_U127, P2_ADD_1119_U128, P2_ADD_1119_U129, P2_ADD_1119_U13, P2_ADD_1119_U130, P2_ADD_1119_U131, P2_ADD_1119_U132, P2_ADD_1119_U133, P2_ADD_1119_U134, P2_ADD_1119_U135, P2_ADD_1119_U136, P2_ADD_1119_U137, P2_ADD_1119_U138, P2_ADD_1119_U139, P2_ADD_1119_U14, P2_ADD_1119_U140, P2_ADD_1119_U141, P2_ADD_1119_U142, P2_ADD_1119_U143, P2_ADD_1119_U144, P2_ADD_1119_U145, P2_ADD_1119_U146, P2_ADD_1119_U147, P2_ADD_1119_U148, P2_ADD_1119_U149, P2_ADD_1119_U15, P2_ADD_1119_U150, P2_ADD_1119_U151, P2_ADD_1119_U152, P2_ADD_1119_U153, P2_ADD_1119_U154, P2_ADD_1119_U155, P2_ADD_1119_U156, P2_ADD_1119_U157, P2_ADD_1119_U16, P2_ADD_1119_U17, P2_ADD_1119_U18, P2_ADD_1119_U19, P2_ADD_1119_U20, P2_ADD_1119_U21, P2_ADD_1119_U22, P2_ADD_1119_U23, P2_ADD_1119_U24, P2_ADD_1119_U25, P2_ADD_1119_U26, P2_ADD_1119_U27, P2_ADD_1119_U28, P2_ADD_1119_U29, P2_ADD_1119_U30, P2_ADD_1119_U31, P2_ADD_1119_U32, P2_ADD_1119_U33, P2_ADD_1119_U34, P2_ADD_1119_U35, P2_ADD_1119_U36, P2_ADD_1119_U37, P2_ADD_1119_U38, P2_ADD_1119_U39, P2_ADD_1119_U4, P2_ADD_1119_U40, P2_ADD_1119_U41, P2_ADD_1119_U42, P2_ADD_1119_U43, P2_ADD_1119_U44, P2_ADD_1119_U45, P2_ADD_1119_U46, P2_ADD_1119_U47, P2_ADD_1119_U48, P2_ADD_1119_U49, P2_ADD_1119_U5, P2_ADD_1119_U50, P2_ADD_1119_U51, P2_ADD_1119_U52, P2_ADD_1119_U53, P2_ADD_1119_U54, P2_ADD_1119_U55, P2_ADD_1119_U56, P2_ADD_1119_U57, P2_ADD_1119_U58, P2_ADD_1119_U59, P2_ADD_1119_U6, P2_ADD_1119_U60, P2_ADD_1119_U61, P2_ADD_1119_U62, P2_ADD_1119_U63, P2_ADD_1119_U64, P2_ADD_1119_U65, P2_ADD_1119_U66, P2_ADD_1119_U67, P2_ADD_1119_U68, P2_ADD_1119_U69, P2_ADD_1119_U7, P2_ADD_1119_U70, P2_ADD_1119_U71, P2_ADD_1119_U72, P2_ADD_1119_U73, P2_ADD_1119_U74, P2_ADD_1119_U75, P2_ADD_1119_U76, P2_ADD_1119_U77, P2_ADD_1119_U78, P2_ADD_1119_U79, P2_ADD_1119_U8, P2_ADD_1119_U80, P2_ADD_1119_U81, P2_ADD_1119_U82, P2_ADD_1119_U83, P2_ADD_1119_U84, P2_ADD_1119_U85, P2_ADD_1119_U86, P2_ADD_1119_U87, P2_ADD_1119_U88, P2_ADD_1119_U89, P2_ADD_1119_U9, P2_ADD_1119_U90, P2_ADD_1119_U91, P2_ADD_1119_U92, P2_ADD_1119_U93, P2_ADD_1119_U94, P2_ADD_1119_U95, P2_ADD_1119_U96, P2_ADD_1119_U97, P2_ADD_1119_U98, P2_ADD_1119_U99, P2_R1113_U10, P2_R1113_U100, P2_R1113_U101, P2_R1113_U102, P2_R1113_U103, P2_R1113_U104, P2_R1113_U105, P2_R1113_U106, P2_R1113_U107, P2_R1113_U108, P2_R1113_U109, P2_R1113_U11, P2_R1113_U110, P2_R1113_U111, P2_R1113_U112, P2_R1113_U113, P2_R1113_U114, P2_R1113_U115, P2_R1113_U116, P2_R1113_U117, P2_R1113_U118, P2_R1113_U119, P2_R1113_U12, P2_R1113_U120, P2_R1113_U121, P2_R1113_U122, P2_R1113_U123, P2_R1113_U124, P2_R1113_U125, P2_R1113_U126, P2_R1113_U127, P2_R1113_U128, P2_R1113_U129, P2_R1113_U13, P2_R1113_U130, P2_R1113_U131, P2_R1113_U132, P2_R1113_U133, P2_R1113_U134, P2_R1113_U135, P2_R1113_U136, P2_R1113_U137, P2_R1113_U138, P2_R1113_U139, P2_R1113_U14, P2_R1113_U140, P2_R1113_U141, P2_R1113_U142, P2_R1113_U143, P2_R1113_U144, P2_R1113_U145, P2_R1113_U146, P2_R1113_U147, P2_R1113_U148, P2_R1113_U149, P2_R1113_U15, P2_R1113_U150, P2_R1113_U151, P2_R1113_U152, P2_R1113_U153, P2_R1113_U154, P2_R1113_U155, P2_R1113_U156, P2_R1113_U157, P2_R1113_U158, P2_R1113_U159, P2_R1113_U16, P2_R1113_U160, P2_R1113_U161, P2_R1113_U162, P2_R1113_U163, P2_R1113_U164, P2_R1113_U165, P2_R1113_U166, P2_R1113_U167, P2_R1113_U168, P2_R1113_U169, P2_R1113_U17, P2_R1113_U170, P2_R1113_U171, P2_R1113_U172, P2_R1113_U173, P2_R1113_U174, P2_R1113_U175, P2_R1113_U176, P2_R1113_U177, P2_R1113_U178, P2_R1113_U179, P2_R1113_U18, P2_R1113_U180, P2_R1113_U181, P2_R1113_U182, P2_R1113_U183, P2_R1113_U184, P2_R1113_U185, P2_R1113_U186, P2_R1113_U187, P2_R1113_U188, P2_R1113_U189, P2_R1113_U19, P2_R1113_U190, P2_R1113_U191, P2_R1113_U192, P2_R1113_U193, P2_R1113_U194, P2_R1113_U195, P2_R1113_U196, P2_R1113_U197, P2_R1113_U198, P2_R1113_U199, P2_R1113_U20, P2_R1113_U200, P2_R1113_U201, P2_R1113_U202, P2_R1113_U203, P2_R1113_U204, P2_R1113_U205, P2_R1113_U206, P2_R1113_U207, P2_R1113_U208, P2_R1113_U209, P2_R1113_U21, P2_R1113_U210, P2_R1113_U211, P2_R1113_U212, P2_R1113_U213, P2_R1113_U214, P2_R1113_U215, P2_R1113_U216, P2_R1113_U217, P2_R1113_U218, P2_R1113_U219, P2_R1113_U22, P2_R1113_U220, P2_R1113_U221, P2_R1113_U222, P2_R1113_U223, P2_R1113_U224, P2_R1113_U225, P2_R1113_U226, P2_R1113_U227, P2_R1113_U228, P2_R1113_U229, P2_R1113_U23, P2_R1113_U230, P2_R1113_U231, P2_R1113_U232, P2_R1113_U233, P2_R1113_U234, P2_R1113_U235, P2_R1113_U236, P2_R1113_U237, P2_R1113_U238, P2_R1113_U239, P2_R1113_U24, P2_R1113_U240, P2_R1113_U241, P2_R1113_U242, P2_R1113_U243, P2_R1113_U244, P2_R1113_U245, P2_R1113_U246, P2_R1113_U247, P2_R1113_U248, P2_R1113_U249, P2_R1113_U25, P2_R1113_U250, P2_R1113_U251, P2_R1113_U252, P2_R1113_U253, P2_R1113_U254, P2_R1113_U255, P2_R1113_U256, P2_R1113_U257, P2_R1113_U258, P2_R1113_U259, P2_R1113_U26, P2_R1113_U260, P2_R1113_U261, P2_R1113_U262, P2_R1113_U263, P2_R1113_U264, P2_R1113_U265, P2_R1113_U266, P2_R1113_U267, P2_R1113_U268, P2_R1113_U269, P2_R1113_U27, P2_R1113_U270, P2_R1113_U271, P2_R1113_U272, P2_R1113_U273, P2_R1113_U274, P2_R1113_U275, P2_R1113_U276, P2_R1113_U277, P2_R1113_U278, P2_R1113_U279, P2_R1113_U28, P2_R1113_U280, P2_R1113_U281, P2_R1113_U282, P2_R1113_U283, P2_R1113_U284, P2_R1113_U285, P2_R1113_U286, P2_R1113_U287, P2_R1113_U288, P2_R1113_U289, P2_R1113_U29, P2_R1113_U290, P2_R1113_U291, P2_R1113_U292, P2_R1113_U293, P2_R1113_U294, P2_R1113_U295, P2_R1113_U296, P2_R1113_U297, P2_R1113_U298, P2_R1113_U299, P2_R1113_U30, P2_R1113_U300, P2_R1113_U301, P2_R1113_U302, P2_R1113_U303, P2_R1113_U304, P2_R1113_U305, P2_R1113_U306, P2_R1113_U307, P2_R1113_U308, P2_R1113_U309, P2_R1113_U31, P2_R1113_U310, P2_R1113_U311, P2_R1113_U312, P2_R1113_U313, P2_R1113_U314, P2_R1113_U315, P2_R1113_U316, P2_R1113_U317, P2_R1113_U318, P2_R1113_U319, P2_R1113_U32, P2_R1113_U320, P2_R1113_U321, P2_R1113_U322, P2_R1113_U323, P2_R1113_U324, P2_R1113_U325, P2_R1113_U326, P2_R1113_U327, P2_R1113_U328, P2_R1113_U329, P2_R1113_U33, P2_R1113_U330, P2_R1113_U331, P2_R1113_U332, P2_R1113_U333, P2_R1113_U334, P2_R1113_U335, P2_R1113_U336, P2_R1113_U337, P2_R1113_U338, P2_R1113_U339, P2_R1113_U34, P2_R1113_U340, P2_R1113_U341, P2_R1113_U342, P2_R1113_U343, P2_R1113_U344, P2_R1113_U345, P2_R1113_U346, P2_R1113_U347, P2_R1113_U348, P2_R1113_U349, P2_R1113_U35, P2_R1113_U350, P2_R1113_U351, P2_R1113_U352, P2_R1113_U353, P2_R1113_U354, P2_R1113_U355, P2_R1113_U356, P2_R1113_U357, P2_R1113_U358, P2_R1113_U359, P2_R1113_U36, P2_R1113_U360, P2_R1113_U361, P2_R1113_U362, P2_R1113_U363, P2_R1113_U364, P2_R1113_U365, P2_R1113_U366, P2_R1113_U367, P2_R1113_U368, P2_R1113_U369, P2_R1113_U37, P2_R1113_U370, P2_R1113_U371, P2_R1113_U372, P2_R1113_U373, P2_R1113_U374, P2_R1113_U375, P2_R1113_U376, P2_R1113_U377, P2_R1113_U378, P2_R1113_U379, P2_R1113_U38, P2_R1113_U380, P2_R1113_U381, P2_R1113_U382, P2_R1113_U383, P2_R1113_U384, P2_R1113_U385, P2_R1113_U386, P2_R1113_U387, P2_R1113_U388, P2_R1113_U389, P2_R1113_U39, P2_R1113_U390, P2_R1113_U391, P2_R1113_U392, P2_R1113_U393, P2_R1113_U394, P2_R1113_U395, P2_R1113_U396, P2_R1113_U397, P2_R1113_U398, P2_R1113_U399, P2_R1113_U40, P2_R1113_U400, P2_R1113_U401, P2_R1113_U402, P2_R1113_U403, P2_R1113_U404, P2_R1113_U405, P2_R1113_U406, P2_R1113_U407, P2_R1113_U408, P2_R1113_U409, P2_R1113_U41, P2_R1113_U410, P2_R1113_U411, P2_R1113_U412, P2_R1113_U413, P2_R1113_U414, P2_R1113_U415, P2_R1113_U416, P2_R1113_U417, P2_R1113_U418, P2_R1113_U419, P2_R1113_U42, P2_R1113_U420, P2_R1113_U421, P2_R1113_U422, P2_R1113_U423, P2_R1113_U424, P2_R1113_U425, P2_R1113_U426, P2_R1113_U427, P2_R1113_U428, P2_R1113_U429, P2_R1113_U43, P2_R1113_U430, P2_R1113_U431, P2_R1113_U432, P2_R1113_U433, P2_R1113_U434, P2_R1113_U435, P2_R1113_U436, P2_R1113_U437, P2_R1113_U438, P2_R1113_U439, P2_R1113_U44, P2_R1113_U440, P2_R1113_U441, P2_R1113_U442, P2_R1113_U443, P2_R1113_U444, P2_R1113_U445, P2_R1113_U446, P2_R1113_U447, P2_R1113_U448, P2_R1113_U449, P2_R1113_U45, P2_R1113_U450, P2_R1113_U451, P2_R1113_U452, P2_R1113_U453, P2_R1113_U454, P2_R1113_U455, P2_R1113_U456, P2_R1113_U457, P2_R1113_U458, P2_R1113_U459, P2_R1113_U46, P2_R1113_U460, P2_R1113_U461, P2_R1113_U462, P2_R1113_U463, P2_R1113_U464, P2_R1113_U465, P2_R1113_U466, P2_R1113_U467, P2_R1113_U468, P2_R1113_U469, P2_R1113_U47, P2_R1113_U470, P2_R1113_U471, P2_R1113_U472, P2_R1113_U473, P2_R1113_U474, P2_R1113_U475, P2_R1113_U476, P2_R1113_U477, P2_R1113_U478, P2_R1113_U48, P2_R1113_U49, P2_R1113_U50, P2_R1113_U51, P2_R1113_U52, P2_R1113_U53, P2_R1113_U54, P2_R1113_U55, P2_R1113_U56, P2_R1113_U57, P2_R1113_U58, P2_R1113_U59, P2_R1113_U6, P2_R1113_U60, P2_R1113_U61, P2_R1113_U62, P2_R1113_U63, P2_R1113_U64, P2_R1113_U65, P2_R1113_U66, P2_R1113_U67, P2_R1113_U68, P2_R1113_U69, P2_R1113_U7, P2_R1113_U70, P2_R1113_U71, P2_R1113_U72, P2_R1113_U73, P2_R1113_U74, P2_R1113_U75, P2_R1113_U76, P2_R1113_U77, P2_R1113_U78, P2_R1113_U79, P2_R1113_U8, P2_R1113_U80, P2_R1113_U81, P2_R1113_U82, P2_R1113_U83, P2_R1113_U84, P2_R1113_U85, P2_R1113_U86, P2_R1113_U87, P2_R1113_U88, P2_R1113_U89, P2_R1113_U9, P2_R1113_U90, P2_R1113_U91, P2_R1113_U92, P2_R1113_U93, P2_R1113_U94, P2_R1113_U95, P2_R1113_U96, P2_R1113_U97, P2_R1113_U98, P2_R1113_U99, P2_R1131_U10, P2_R1131_U100, P2_R1131_U101, P2_R1131_U102, P2_R1131_U103, P2_R1131_U104, P2_R1131_U105, P2_R1131_U106, P2_R1131_U107, P2_R1131_U108, P2_R1131_U109, P2_R1131_U11, P2_R1131_U110, P2_R1131_U111, P2_R1131_U112, P2_R1131_U113, P2_R1131_U114, P2_R1131_U115, P2_R1131_U116, P2_R1131_U117, P2_R1131_U118, P2_R1131_U119, P2_R1131_U12, P2_R1131_U120, P2_R1131_U121, P2_R1131_U122, P2_R1131_U123, P2_R1131_U124, P2_R1131_U125, P2_R1131_U126, P2_R1131_U127, P2_R1131_U128, P2_R1131_U129, P2_R1131_U13, P2_R1131_U130, P2_R1131_U131, P2_R1131_U132, P2_R1131_U133, P2_R1131_U134, P2_R1131_U135, P2_R1131_U136, P2_R1131_U137, P2_R1131_U138, P2_R1131_U139, P2_R1131_U14, P2_R1131_U140, P2_R1131_U141, P2_R1131_U142, P2_R1131_U143, P2_R1131_U144, P2_R1131_U145, P2_R1131_U146, P2_R1131_U147, P2_R1131_U148, P2_R1131_U149, P2_R1131_U15, P2_R1131_U150, P2_R1131_U151, P2_R1131_U152, P2_R1131_U153, P2_R1131_U154, P2_R1131_U155, P2_R1131_U156, P2_R1131_U157, P2_R1131_U158, P2_R1131_U159, P2_R1131_U16, P2_R1131_U160, P2_R1131_U161, P2_R1131_U162, P2_R1131_U163, P2_R1131_U164, P2_R1131_U165, P2_R1131_U166, P2_R1131_U167, P2_R1131_U168, P2_R1131_U169, P2_R1131_U17, P2_R1131_U170, P2_R1131_U171, P2_R1131_U172, P2_R1131_U173, P2_R1131_U174, P2_R1131_U175, P2_R1131_U176, P2_R1131_U177, P2_R1131_U178, P2_R1131_U179, P2_R1131_U18, P2_R1131_U180, P2_R1131_U181, P2_R1131_U182, P2_R1131_U183, P2_R1131_U184, P2_R1131_U185, P2_R1131_U186, P2_R1131_U187, P2_R1131_U188, P2_R1131_U189, P2_R1131_U19, P2_R1131_U190, P2_R1131_U191, P2_R1131_U192, P2_R1131_U193, P2_R1131_U194, P2_R1131_U195, P2_R1131_U196, P2_R1131_U197, P2_R1131_U198, P2_R1131_U199, P2_R1131_U20, P2_R1131_U200, P2_R1131_U201, P2_R1131_U202, P2_R1131_U203, P2_R1131_U204, P2_R1131_U205, P2_R1131_U206, P2_R1131_U207, P2_R1131_U208, P2_R1131_U209, P2_R1131_U21, P2_R1131_U210, P2_R1131_U211, P2_R1131_U212, P2_R1131_U213, P2_R1131_U214, P2_R1131_U215, P2_R1131_U216, P2_R1131_U217, P2_R1131_U218, P2_R1131_U219, P2_R1131_U22, P2_R1131_U220, P2_R1131_U221, P2_R1131_U222, P2_R1131_U223, P2_R1131_U224, P2_R1131_U225, P2_R1131_U226, P2_R1131_U227, P2_R1131_U228, P2_R1131_U229, P2_R1131_U23, P2_R1131_U230, P2_R1131_U231, P2_R1131_U232, P2_R1131_U233, P2_R1131_U234, P2_R1131_U235, P2_R1131_U236, P2_R1131_U237, P2_R1131_U238, P2_R1131_U239, P2_R1131_U24, P2_R1131_U240, P2_R1131_U241, P2_R1131_U242, P2_R1131_U243, P2_R1131_U244, P2_R1131_U245, P2_R1131_U246, P2_R1131_U247, P2_R1131_U248, P2_R1131_U249, P2_R1131_U25, P2_R1131_U250, P2_R1131_U251, P2_R1131_U252, P2_R1131_U253, P2_R1131_U254, P2_R1131_U255, P2_R1131_U256, P2_R1131_U257, P2_R1131_U258, P2_R1131_U259, P2_R1131_U26, P2_R1131_U260, P2_R1131_U261, P2_R1131_U262, P2_R1131_U263, P2_R1131_U264, P2_R1131_U265, P2_R1131_U266, P2_R1131_U267, P2_R1131_U268, P2_R1131_U269, P2_R1131_U27, P2_R1131_U270, P2_R1131_U271, P2_R1131_U272, P2_R1131_U273, P2_R1131_U274, P2_R1131_U275, P2_R1131_U276, P2_R1131_U277, P2_R1131_U278, P2_R1131_U279, P2_R1131_U28, P2_R1131_U280, P2_R1131_U281, P2_R1131_U282, P2_R1131_U283, P2_R1131_U284, P2_R1131_U285, P2_R1131_U286, P2_R1131_U287, P2_R1131_U288, P2_R1131_U289, P2_R1131_U29, P2_R1131_U290, P2_R1131_U291, P2_R1131_U292, P2_R1131_U293, P2_R1131_U294, P2_R1131_U295, P2_R1131_U296, P2_R1131_U297, P2_R1131_U298, P2_R1131_U299, P2_R1131_U30, P2_R1131_U300, P2_R1131_U301, P2_R1131_U302, P2_R1131_U303, P2_R1131_U304, P2_R1131_U305, P2_R1131_U306, P2_R1131_U307, P2_R1131_U308, P2_R1131_U309, P2_R1131_U31, P2_R1131_U310, P2_R1131_U311, P2_R1131_U312, P2_R1131_U313, P2_R1131_U314, P2_R1131_U315, P2_R1131_U316, P2_R1131_U317, P2_R1131_U318, P2_R1131_U319, P2_R1131_U32, P2_R1131_U320, P2_R1131_U321, P2_R1131_U322, P2_R1131_U323, P2_R1131_U324, P2_R1131_U325, P2_R1131_U326, P2_R1131_U327, P2_R1131_U328, P2_R1131_U329, P2_R1131_U33, P2_R1131_U330, P2_R1131_U331, P2_R1131_U332, P2_R1131_U333, P2_R1131_U334, P2_R1131_U335, P2_R1131_U336, P2_R1131_U337, P2_R1131_U338, P2_R1131_U339, P2_R1131_U34, P2_R1131_U340, P2_R1131_U341, P2_R1131_U342, P2_R1131_U343, P2_R1131_U344, P2_R1131_U345, P2_R1131_U346, P2_R1131_U347, P2_R1131_U348, P2_R1131_U349, P2_R1131_U35, P2_R1131_U350, P2_R1131_U351, P2_R1131_U352, P2_R1131_U353, P2_R1131_U354, P2_R1131_U355, P2_R1131_U356, P2_R1131_U357, P2_R1131_U358, P2_R1131_U359, P2_R1131_U36, P2_R1131_U360, P2_R1131_U361, P2_R1131_U362, P2_R1131_U363, P2_R1131_U364, P2_R1131_U365, P2_R1131_U366, P2_R1131_U367, P2_R1131_U368, P2_R1131_U369, P2_R1131_U37, P2_R1131_U370, P2_R1131_U371, P2_R1131_U372, P2_R1131_U373, P2_R1131_U374, P2_R1131_U375, P2_R1131_U376, P2_R1131_U377, P2_R1131_U378, P2_R1131_U379, P2_R1131_U38, P2_R1131_U380, P2_R1131_U381, P2_R1131_U382, P2_R1131_U383, P2_R1131_U384, P2_R1131_U385, P2_R1131_U386, P2_R1131_U387, P2_R1131_U388, P2_R1131_U389, P2_R1131_U39, P2_R1131_U390, P2_R1131_U391, P2_R1131_U392, P2_R1131_U393, P2_R1131_U394, P2_R1131_U395, P2_R1131_U396, P2_R1131_U397, P2_R1131_U398, P2_R1131_U399, P2_R1131_U4, P2_R1131_U40, P2_R1131_U400, P2_R1131_U401, P2_R1131_U402, P2_R1131_U403, P2_R1131_U404, P2_R1131_U405, P2_R1131_U406, P2_R1131_U407, P2_R1131_U408, P2_R1131_U409, P2_R1131_U41, P2_R1131_U410, P2_R1131_U411, P2_R1131_U412, P2_R1131_U413, P2_R1131_U414, P2_R1131_U415, P2_R1131_U416, P2_R1131_U417, P2_R1131_U418, P2_R1131_U419, P2_R1131_U42, P2_R1131_U420, P2_R1131_U421, P2_R1131_U422, P2_R1131_U423, P2_R1131_U424, P2_R1131_U425, P2_R1131_U426, P2_R1131_U427, P2_R1131_U428, P2_R1131_U429, P2_R1131_U43, P2_R1131_U430, P2_R1131_U431, P2_R1131_U432, P2_R1131_U433, P2_R1131_U434, P2_R1131_U435, P2_R1131_U436, P2_R1131_U437, P2_R1131_U438, P2_R1131_U439, P2_R1131_U44, P2_R1131_U440, P2_R1131_U441, P2_R1131_U442, P2_R1131_U443, P2_R1131_U444, P2_R1131_U445, P2_R1131_U446, P2_R1131_U447, P2_R1131_U448, P2_R1131_U449, P2_R1131_U45, P2_R1131_U450, P2_R1131_U451, P2_R1131_U452, P2_R1131_U453, P2_R1131_U454, P2_R1131_U455, P2_R1131_U456, P2_R1131_U457, P2_R1131_U458, P2_R1131_U459, P2_R1131_U46, P2_R1131_U460, P2_R1131_U461, P2_R1131_U462, P2_R1131_U463, P2_R1131_U464, P2_R1131_U465, P2_R1131_U466, P2_R1131_U467, P2_R1131_U468, P2_R1131_U469, P2_R1131_U47, P2_R1131_U470, P2_R1131_U471, P2_R1131_U472, P2_R1131_U473, P2_R1131_U474, P2_R1131_U475, P2_R1131_U476, P2_R1131_U477, P2_R1131_U478, P2_R1131_U479, P2_R1131_U48, P2_R1131_U480, P2_R1131_U481, P2_R1131_U482, P2_R1131_U483, P2_R1131_U484, P2_R1131_U485, P2_R1131_U486, P2_R1131_U487, P2_R1131_U488, P2_R1131_U489, P2_R1131_U49, P2_R1131_U490, P2_R1131_U491, P2_R1131_U492, P2_R1131_U493, P2_R1131_U494, P2_R1131_U495, P2_R1131_U496, P2_R1131_U497, P2_R1131_U498, P2_R1131_U499, P2_R1131_U5, P2_R1131_U50, P2_R1131_U500, P2_R1131_U501, P2_R1131_U502, P2_R1131_U503, P2_R1131_U504, P2_R1131_U51, P2_R1131_U52, P2_R1131_U53, P2_R1131_U54, P2_R1131_U55, P2_R1131_U56, P2_R1131_U57, P2_R1131_U58, P2_R1131_U59, P2_R1131_U6, P2_R1131_U60, P2_R1131_U61, P2_R1131_U62, P2_R1131_U63, P2_R1131_U64, P2_R1131_U65, P2_R1131_U66, P2_R1131_U67, P2_R1131_U68, P2_R1131_U69, P2_R1131_U7, P2_R1131_U70, P2_R1131_U71, P2_R1131_U72, P2_R1131_U73, P2_R1131_U74, P2_R1131_U75, P2_R1131_U76, P2_R1131_U77, P2_R1131_U78, P2_R1131_U79, P2_R1131_U8, P2_R1131_U80, P2_R1131_U81, P2_R1131_U82, P2_R1131_U83, P2_R1131_U84, P2_R1131_U85, P2_R1131_U86, P2_R1131_U87, P2_R1131_U88, P2_R1131_U89, P2_R1131_U9, P2_R1131_U90, P2_R1131_U91, P2_R1131_U92, P2_R1131_U93, P2_R1131_U94, P2_R1131_U95, P2_R1131_U96, P2_R1131_U97, P2_R1131_U98, P2_R1131_U99, P2_R1146_U10, P2_R1146_U100, P2_R1146_U101, P2_R1146_U102, P2_R1146_U103, P2_R1146_U104, P2_R1146_U105, P2_R1146_U106, P2_R1146_U107, P2_R1146_U108, P2_R1146_U109, P2_R1146_U11, P2_R1146_U110, P2_R1146_U111, P2_R1146_U112, P2_R1146_U113, P2_R1146_U114, P2_R1146_U115, P2_R1146_U116, P2_R1146_U117, P2_R1146_U118, P2_R1146_U119, P2_R1146_U12, P2_R1146_U120, P2_R1146_U121, P2_R1146_U122, P2_R1146_U123, P2_R1146_U124, P2_R1146_U125, P2_R1146_U126, P2_R1146_U127, P2_R1146_U128, P2_R1146_U129, P2_R1146_U13, P2_R1146_U130, P2_R1146_U131, P2_R1146_U132, P2_R1146_U133, P2_R1146_U134, P2_R1146_U135, P2_R1146_U136, P2_R1146_U137, P2_R1146_U138, P2_R1146_U139, P2_R1146_U14, P2_R1146_U140, P2_R1146_U141, P2_R1146_U142, P2_R1146_U143, P2_R1146_U144, P2_R1146_U145, P2_R1146_U146, P2_R1146_U147, P2_R1146_U148, P2_R1146_U149, P2_R1146_U15, P2_R1146_U150, P2_R1146_U151, P2_R1146_U152, P2_R1146_U153, P2_R1146_U154, P2_R1146_U155, P2_R1146_U156, P2_R1146_U157, P2_R1146_U158, P2_R1146_U159, P2_R1146_U16, P2_R1146_U160, P2_R1146_U161, P2_R1146_U162, P2_R1146_U163, P2_R1146_U164, P2_R1146_U165, P2_R1146_U166, P2_R1146_U167, P2_R1146_U168, P2_R1146_U169, P2_R1146_U17, P2_R1146_U170, P2_R1146_U171, P2_R1146_U172, P2_R1146_U173, P2_R1146_U174, P2_R1146_U175, P2_R1146_U176, P2_R1146_U177, P2_R1146_U178, P2_R1146_U179, P2_R1146_U18, P2_R1146_U180, P2_R1146_U181, P2_R1146_U182, P2_R1146_U183, P2_R1146_U184, P2_R1146_U185, P2_R1146_U186, P2_R1146_U187, P2_R1146_U188, P2_R1146_U189, P2_R1146_U19, P2_R1146_U190, P2_R1146_U191, P2_R1146_U192, P2_R1146_U193, P2_R1146_U194, P2_R1146_U195, P2_R1146_U196, P2_R1146_U197, P2_R1146_U198, P2_R1146_U199, P2_R1146_U20, P2_R1146_U200, P2_R1146_U201, P2_R1146_U202, P2_R1146_U203, P2_R1146_U204, P2_R1146_U205, P2_R1146_U206, P2_R1146_U207, P2_R1146_U208, P2_R1146_U209, P2_R1146_U21, P2_R1146_U210, P2_R1146_U211, P2_R1146_U212, P2_R1146_U213, P2_R1146_U214, P2_R1146_U215, P2_R1146_U216, P2_R1146_U217, P2_R1146_U218, P2_R1146_U219, P2_R1146_U22, P2_R1146_U220, P2_R1146_U221, P2_R1146_U222, P2_R1146_U223, P2_R1146_U224, P2_R1146_U225, P2_R1146_U226, P2_R1146_U227, P2_R1146_U228, P2_R1146_U229, P2_R1146_U23, P2_R1146_U230, P2_R1146_U231, P2_R1146_U232, P2_R1146_U233, P2_R1146_U234, P2_R1146_U235, P2_R1146_U236, P2_R1146_U237, P2_R1146_U238, P2_R1146_U239, P2_R1146_U24, P2_R1146_U240, P2_R1146_U241, P2_R1146_U242, P2_R1146_U243, P2_R1146_U244, P2_R1146_U245, P2_R1146_U246, P2_R1146_U247, P2_R1146_U248, P2_R1146_U249, P2_R1146_U25, P2_R1146_U250, P2_R1146_U251, P2_R1146_U252, P2_R1146_U253, P2_R1146_U254, P2_R1146_U255, P2_R1146_U256, P2_R1146_U257, P2_R1146_U258, P2_R1146_U259, P2_R1146_U26, P2_R1146_U260, P2_R1146_U261, P2_R1146_U262, P2_R1146_U263, P2_R1146_U264, P2_R1146_U265, P2_R1146_U266, P2_R1146_U267, P2_R1146_U268, P2_R1146_U269, P2_R1146_U27, P2_R1146_U270, P2_R1146_U271, P2_R1146_U272, P2_R1146_U273, P2_R1146_U274, P2_R1146_U275, P2_R1146_U276, P2_R1146_U277, P2_R1146_U278, P2_R1146_U279, P2_R1146_U28, P2_R1146_U280, P2_R1146_U281, P2_R1146_U282, P2_R1146_U283, P2_R1146_U284, P2_R1146_U285, P2_R1146_U286, P2_R1146_U287, P2_R1146_U288, P2_R1146_U289, P2_R1146_U29, P2_R1146_U290, P2_R1146_U291, P2_R1146_U292, P2_R1146_U293, P2_R1146_U294, P2_R1146_U295, P2_R1146_U296, P2_R1146_U297, P2_R1146_U298, P2_R1146_U299, P2_R1146_U30, P2_R1146_U300, P2_R1146_U301, P2_R1146_U302, P2_R1146_U303, P2_R1146_U304, P2_R1146_U305, P2_R1146_U306, P2_R1146_U307, P2_R1146_U308, P2_R1146_U309, P2_R1146_U31, P2_R1146_U310, P2_R1146_U311, P2_R1146_U312, P2_R1146_U313, P2_R1146_U314, P2_R1146_U315, P2_R1146_U316, P2_R1146_U317, P2_R1146_U318, P2_R1146_U319, P2_R1146_U32, P2_R1146_U320, P2_R1146_U321, P2_R1146_U322, P2_R1146_U323, P2_R1146_U324, P2_R1146_U325, P2_R1146_U326, P2_R1146_U327, P2_R1146_U328, P2_R1146_U329, P2_R1146_U33, P2_R1146_U330, P2_R1146_U331, P2_R1146_U332, P2_R1146_U333, P2_R1146_U334, P2_R1146_U335, P2_R1146_U336, P2_R1146_U337, P2_R1146_U338, P2_R1146_U339, P2_R1146_U34, P2_R1146_U340, P2_R1146_U341, P2_R1146_U342, P2_R1146_U343, P2_R1146_U344, P2_R1146_U345, P2_R1146_U346, P2_R1146_U347, P2_R1146_U348, P2_R1146_U349, P2_R1146_U35, P2_R1146_U350, P2_R1146_U351, P2_R1146_U352, P2_R1146_U353, P2_R1146_U354, P2_R1146_U355, P2_R1146_U356, P2_R1146_U357, P2_R1146_U358, P2_R1146_U359, P2_R1146_U36, P2_R1146_U360, P2_R1146_U361, P2_R1146_U362, P2_R1146_U363, P2_R1146_U364, P2_R1146_U365, P2_R1146_U366, P2_R1146_U367, P2_R1146_U368, P2_R1146_U369, P2_R1146_U37, P2_R1146_U370, P2_R1146_U371, P2_R1146_U372, P2_R1146_U373, P2_R1146_U374, P2_R1146_U375, P2_R1146_U376, P2_R1146_U377, P2_R1146_U378, P2_R1146_U379, P2_R1146_U38, P2_R1146_U380, P2_R1146_U381, P2_R1146_U382, P2_R1146_U383, P2_R1146_U384, P2_R1146_U385, P2_R1146_U386, P2_R1146_U387, P2_R1146_U388, P2_R1146_U389, P2_R1146_U39, P2_R1146_U390, P2_R1146_U391, P2_R1146_U392, P2_R1146_U393, P2_R1146_U394, P2_R1146_U395, P2_R1146_U396, P2_R1146_U397, P2_R1146_U398, P2_R1146_U399, P2_R1146_U40, P2_R1146_U400, P2_R1146_U401, P2_R1146_U402, P2_R1146_U403, P2_R1146_U404, P2_R1146_U405, P2_R1146_U406, P2_R1146_U407, P2_R1146_U408, P2_R1146_U409, P2_R1146_U41, P2_R1146_U410, P2_R1146_U411, P2_R1146_U412, P2_R1146_U413, P2_R1146_U414, P2_R1146_U415, P2_R1146_U416, P2_R1146_U417, P2_R1146_U418, P2_R1146_U419, P2_R1146_U42, P2_R1146_U420, P2_R1146_U421, P2_R1146_U422, P2_R1146_U423, P2_R1146_U424, P2_R1146_U425, P2_R1146_U426, P2_R1146_U427, P2_R1146_U428, P2_R1146_U429, P2_R1146_U43, P2_R1146_U430, P2_R1146_U431, P2_R1146_U432, P2_R1146_U433, P2_R1146_U434, P2_R1146_U435, P2_R1146_U436, P2_R1146_U437, P2_R1146_U438, P2_R1146_U439, P2_R1146_U44, P2_R1146_U440, P2_R1146_U441, P2_R1146_U442, P2_R1146_U443, P2_R1146_U444, P2_R1146_U445, P2_R1146_U446, P2_R1146_U447, P2_R1146_U448, P2_R1146_U449, P2_R1146_U45, P2_R1146_U450, P2_R1146_U451, P2_R1146_U452, P2_R1146_U453, P2_R1146_U454, P2_R1146_U455, P2_R1146_U456, P2_R1146_U457, P2_R1146_U458, P2_R1146_U459, P2_R1146_U46, P2_R1146_U460, P2_R1146_U461, P2_R1146_U462, P2_R1146_U463, P2_R1146_U464, P2_R1146_U465, P2_R1146_U466, P2_R1146_U467, P2_R1146_U468, P2_R1146_U469, P2_R1146_U47, P2_R1146_U470, P2_R1146_U471, P2_R1146_U472, P2_R1146_U473, P2_R1146_U474, P2_R1146_U475, P2_R1146_U476, P2_R1146_U477, P2_R1146_U478, P2_R1146_U48, P2_R1146_U49, P2_R1146_U50, P2_R1146_U51, P2_R1146_U52, P2_R1146_U53, P2_R1146_U54, P2_R1146_U55, P2_R1146_U56, P2_R1146_U57, P2_R1146_U58, P2_R1146_U59, P2_R1146_U6, P2_R1146_U60, P2_R1146_U61, P2_R1146_U62, P2_R1146_U63, P2_R1146_U64, P2_R1146_U65, P2_R1146_U66, P2_R1146_U67, P2_R1146_U68, P2_R1146_U69, P2_R1146_U7, P2_R1146_U70, P2_R1146_U71, P2_R1146_U72, P2_R1146_U73, P2_R1146_U74, P2_R1146_U75, P2_R1146_U76, P2_R1146_U77, P2_R1146_U78, P2_R1146_U79, P2_R1146_U8, P2_R1146_U80, P2_R1146_U81, P2_R1146_U82, P2_R1146_U83, P2_R1146_U84, P2_R1146_U85, P2_R1146_U86, P2_R1146_U87, P2_R1146_U88, P2_R1146_U89, P2_R1146_U9, P2_R1146_U90, P2_R1146_U91, P2_R1146_U92, P2_R1146_U93, P2_R1146_U94, P2_R1146_U95, P2_R1146_U96, P2_R1146_U97, P2_R1146_U98, P2_R1146_U99, P2_R1164_U10, P2_R1164_U100, P2_R1164_U101, P2_R1164_U102, P2_R1164_U103, P2_R1164_U104, P2_R1164_U105, P2_R1164_U106, P2_R1164_U107, P2_R1164_U108, P2_R1164_U109, P2_R1164_U11, P2_R1164_U110, P2_R1164_U111, P2_R1164_U112, P2_R1164_U113, P2_R1164_U114, P2_R1164_U115, P2_R1164_U116, P2_R1164_U117, P2_R1164_U118, P2_R1164_U119, P2_R1164_U12, P2_R1164_U120, P2_R1164_U121, P2_R1164_U122, P2_R1164_U123, P2_R1164_U124, P2_R1164_U125, P2_R1164_U126, P2_R1164_U127, P2_R1164_U128, P2_R1164_U129, P2_R1164_U13, P2_R1164_U130, P2_R1164_U131, P2_R1164_U132, P2_R1164_U133, P2_R1164_U134, P2_R1164_U135, P2_R1164_U136, P2_R1164_U137, P2_R1164_U138, P2_R1164_U139, P2_R1164_U14, P2_R1164_U140, P2_R1164_U141, P2_R1164_U142, P2_R1164_U143, P2_R1164_U144, P2_R1164_U145, P2_R1164_U146, P2_R1164_U147, P2_R1164_U148, P2_R1164_U149, P2_R1164_U15, P2_R1164_U150, P2_R1164_U151, P2_R1164_U152, P2_R1164_U153, P2_R1164_U154, P2_R1164_U155, P2_R1164_U156, P2_R1164_U157, P2_R1164_U158, P2_R1164_U159, P2_R1164_U16, P2_R1164_U160, P2_R1164_U161, P2_R1164_U162, P2_R1164_U163, P2_R1164_U164, P2_R1164_U165, P2_R1164_U166, P2_R1164_U167, P2_R1164_U168, P2_R1164_U169, P2_R1164_U17, P2_R1164_U170, P2_R1164_U171, P2_R1164_U172, P2_R1164_U173, P2_R1164_U174, P2_R1164_U175, P2_R1164_U176, P2_R1164_U177, P2_R1164_U178, P2_R1164_U179, P2_R1164_U18, P2_R1164_U180, P2_R1164_U181, P2_R1164_U182, P2_R1164_U183, P2_R1164_U184, P2_R1164_U185, P2_R1164_U186, P2_R1164_U187, P2_R1164_U188, P2_R1164_U189, P2_R1164_U19, P2_R1164_U190, P2_R1164_U191, P2_R1164_U192, P2_R1164_U193, P2_R1164_U194, P2_R1164_U195, P2_R1164_U196, P2_R1164_U197, P2_R1164_U198, P2_R1164_U199, P2_R1164_U20, P2_R1164_U200, P2_R1164_U201, P2_R1164_U202, P2_R1164_U203, P2_R1164_U204, P2_R1164_U205, P2_R1164_U206, P2_R1164_U207, P2_R1164_U208, P2_R1164_U209, P2_R1164_U21, P2_R1164_U210, P2_R1164_U211, P2_R1164_U212, P2_R1164_U213, P2_R1164_U214, P2_R1164_U215, P2_R1164_U216, P2_R1164_U217, P2_R1164_U218, P2_R1164_U219, P2_R1164_U22, P2_R1164_U220, P2_R1164_U221, P2_R1164_U222, P2_R1164_U223, P2_R1164_U224, P2_R1164_U225, P2_R1164_U226, P2_R1164_U227, P2_R1164_U228, P2_R1164_U229, P2_R1164_U23, P2_R1164_U230, P2_R1164_U231, P2_R1164_U232, P2_R1164_U233, P2_R1164_U234, P2_R1164_U235, P2_R1164_U236, P2_R1164_U237, P2_R1164_U238, P2_R1164_U239, P2_R1164_U24, P2_R1164_U240, P2_R1164_U241, P2_R1164_U242, P2_R1164_U243, P2_R1164_U244, P2_R1164_U245, P2_R1164_U246, P2_R1164_U247, P2_R1164_U248, P2_R1164_U249, P2_R1164_U25, P2_R1164_U250, P2_R1164_U251, P2_R1164_U252, P2_R1164_U253, P2_R1164_U254, P2_R1164_U255, P2_R1164_U256, P2_R1164_U257, P2_R1164_U258, P2_R1164_U259, P2_R1164_U26, P2_R1164_U260, P2_R1164_U261, P2_R1164_U262, P2_R1164_U263, P2_R1164_U264, P2_R1164_U265, P2_R1164_U266, P2_R1164_U267, P2_R1164_U268, P2_R1164_U269, P2_R1164_U27, P2_R1164_U270, P2_R1164_U271, P2_R1164_U272, P2_R1164_U273, P2_R1164_U274, P2_R1164_U275, P2_R1164_U276, P2_R1164_U277, P2_R1164_U278, P2_R1164_U279, P2_R1164_U28, P2_R1164_U280, P2_R1164_U281, P2_R1164_U282, P2_R1164_U283, P2_R1164_U284, P2_R1164_U285, P2_R1164_U286, P2_R1164_U287, P2_R1164_U288, P2_R1164_U289, P2_R1164_U29, P2_R1164_U290, P2_R1164_U291, P2_R1164_U292, P2_R1164_U293, P2_R1164_U294, P2_R1164_U295, P2_R1164_U296, P2_R1164_U297, P2_R1164_U298, P2_R1164_U299, P2_R1164_U30, P2_R1164_U300, P2_R1164_U301, P2_R1164_U302, P2_R1164_U303, P2_R1164_U304, P2_R1164_U305, P2_R1164_U306, P2_R1164_U307, P2_R1164_U308, P2_R1164_U309, P2_R1164_U31, P2_R1164_U310, P2_R1164_U311, P2_R1164_U312, P2_R1164_U313, P2_R1164_U314, P2_R1164_U315, P2_R1164_U316, P2_R1164_U317, P2_R1164_U318, P2_R1164_U319, P2_R1164_U32, P2_R1164_U320, P2_R1164_U321, P2_R1164_U322, P2_R1164_U323, P2_R1164_U324, P2_R1164_U325, P2_R1164_U326, P2_R1164_U327, P2_R1164_U328, P2_R1164_U329, P2_R1164_U33, P2_R1164_U330, P2_R1164_U331, P2_R1164_U332, P2_R1164_U333, P2_R1164_U334, P2_R1164_U335, P2_R1164_U336, P2_R1164_U337, P2_R1164_U338, P2_R1164_U339, P2_R1164_U34, P2_R1164_U340, P2_R1164_U341, P2_R1164_U342, P2_R1164_U343, P2_R1164_U344, P2_R1164_U345, P2_R1164_U346, P2_R1164_U347, P2_R1164_U348, P2_R1164_U349, P2_R1164_U35, P2_R1164_U350, P2_R1164_U351, P2_R1164_U352, P2_R1164_U353, P2_R1164_U354, P2_R1164_U355, P2_R1164_U356, P2_R1164_U357, P2_R1164_U358, P2_R1164_U359, P2_R1164_U36, P2_R1164_U360, P2_R1164_U361, P2_R1164_U362, P2_R1164_U363, P2_R1164_U364, P2_R1164_U365, P2_R1164_U366, P2_R1164_U367, P2_R1164_U368, P2_R1164_U369, P2_R1164_U37, P2_R1164_U370, P2_R1164_U371, P2_R1164_U372, P2_R1164_U373, P2_R1164_U374, P2_R1164_U375, P2_R1164_U376, P2_R1164_U377, P2_R1164_U378, P2_R1164_U379, P2_R1164_U38, P2_R1164_U380, P2_R1164_U381, P2_R1164_U382, P2_R1164_U383, P2_R1164_U384, P2_R1164_U385, P2_R1164_U386, P2_R1164_U387, P2_R1164_U388, P2_R1164_U389, P2_R1164_U39, P2_R1164_U390, P2_R1164_U391, P2_R1164_U392, P2_R1164_U393, P2_R1164_U394, P2_R1164_U395, P2_R1164_U396, P2_R1164_U397, P2_R1164_U398, P2_R1164_U399, P2_R1164_U4, P2_R1164_U40, P2_R1164_U400, P2_R1164_U401, P2_R1164_U402, P2_R1164_U403, P2_R1164_U404, P2_R1164_U405, P2_R1164_U406, P2_R1164_U407, P2_R1164_U408, P2_R1164_U409, P2_R1164_U41, P2_R1164_U410, P2_R1164_U411, P2_R1164_U412, P2_R1164_U413, P2_R1164_U414, P2_R1164_U415, P2_R1164_U416, P2_R1164_U417, P2_R1164_U418, P2_R1164_U419, P2_R1164_U42, P2_R1164_U420, P2_R1164_U421, P2_R1164_U422, P2_R1164_U423, P2_R1164_U424, P2_R1164_U425, P2_R1164_U426, P2_R1164_U427, P2_R1164_U428, P2_R1164_U429, P2_R1164_U43, P2_R1164_U430, P2_R1164_U431, P2_R1164_U432, P2_R1164_U433, P2_R1164_U434, P2_R1164_U435, P2_R1164_U436, P2_R1164_U437, P2_R1164_U438, P2_R1164_U439, P2_R1164_U44, P2_R1164_U440, P2_R1164_U441, P2_R1164_U442, P2_R1164_U443, P2_R1164_U444, P2_R1164_U445, P2_R1164_U446, P2_R1164_U447, P2_R1164_U448, P2_R1164_U449, P2_R1164_U45, P2_R1164_U450, P2_R1164_U451, P2_R1164_U452, P2_R1164_U453, P2_R1164_U454, P2_R1164_U455, P2_R1164_U456, P2_R1164_U457, P2_R1164_U458, P2_R1164_U459, P2_R1164_U46, P2_R1164_U460, P2_R1164_U461, P2_R1164_U462, P2_R1164_U463, P2_R1164_U464, P2_R1164_U465, P2_R1164_U466, P2_R1164_U467, P2_R1164_U468, P2_R1164_U469, P2_R1164_U47, P2_R1164_U470, P2_R1164_U471, P2_R1164_U472, P2_R1164_U473, P2_R1164_U474, P2_R1164_U475, P2_R1164_U476, P2_R1164_U477, P2_R1164_U478, P2_R1164_U479, P2_R1164_U48, P2_R1164_U480, P2_R1164_U481, P2_R1164_U482, P2_R1164_U483, P2_R1164_U484, P2_R1164_U485, P2_R1164_U486, P2_R1164_U487, P2_R1164_U488, P2_R1164_U489, P2_R1164_U49, P2_R1164_U490, P2_R1164_U491, P2_R1164_U492, P2_R1164_U493, P2_R1164_U494, P2_R1164_U495, P2_R1164_U496, P2_R1164_U497, P2_R1164_U498, P2_R1164_U499, P2_R1164_U5, P2_R1164_U50, P2_R1164_U500, P2_R1164_U501, P2_R1164_U502, P2_R1164_U503, P2_R1164_U504, P2_R1164_U51, P2_R1164_U52, P2_R1164_U53, P2_R1164_U54, P2_R1164_U55, P2_R1164_U56, P2_R1164_U57, P2_R1164_U58, P2_R1164_U59, P2_R1164_U6, P2_R1164_U60, P2_R1164_U61, P2_R1164_U62, P2_R1164_U63, P2_R1164_U64, P2_R1164_U65, P2_R1164_U66, P2_R1164_U67, P2_R1164_U68, P2_R1164_U69, P2_R1164_U7, P2_R1164_U70, P2_R1164_U71, P2_R1164_U72, P2_R1164_U73, P2_R1164_U74, P2_R1164_U75, P2_R1164_U76, P2_R1164_U77, P2_R1164_U78, P2_R1164_U79, P2_R1164_U8, P2_R1164_U80, P2_R1164_U81, P2_R1164_U82, P2_R1164_U83, P2_R1164_U84, P2_R1164_U85, P2_R1164_U86, P2_R1164_U87, P2_R1164_U88, P2_R1164_U89, P2_R1164_U9, P2_R1164_U90, P2_R1164_U91, P2_R1164_U92, P2_R1164_U93, P2_R1164_U94, P2_R1164_U95, P2_R1164_U96, P2_R1164_U97, P2_R1164_U98, P2_R1164_U99, P2_R1170_U10, P2_R1170_U100, P2_R1170_U101, P2_R1170_U102, P2_R1170_U103, P2_R1170_U104, P2_R1170_U105, P2_R1170_U106, P2_R1170_U107, P2_R1170_U108, P2_R1170_U109, P2_R1170_U11, P2_R1170_U110, P2_R1170_U111, P2_R1170_U112, P2_R1170_U113, P2_R1170_U114, P2_R1170_U115, P2_R1170_U116, P2_R1170_U117, P2_R1170_U118, P2_R1170_U119, P2_R1170_U12, P2_R1170_U120, P2_R1170_U121, P2_R1170_U122, P2_R1170_U123, P2_R1170_U124, P2_R1170_U125, P2_R1170_U126, P2_R1170_U127, P2_R1170_U128, P2_R1170_U129, P2_R1170_U13, P2_R1170_U130, P2_R1170_U131, P2_R1170_U132, P2_R1170_U133, P2_R1170_U134, P2_R1170_U135, P2_R1170_U136, P2_R1170_U137, P2_R1170_U138, P2_R1170_U139, P2_R1170_U14, P2_R1170_U140, P2_R1170_U141, P2_R1170_U142, P2_R1170_U143, P2_R1170_U144, P2_R1170_U145, P2_R1170_U146, P2_R1170_U147, P2_R1170_U148, P2_R1170_U149, P2_R1170_U15, P2_R1170_U150, P2_R1170_U151, P2_R1170_U152, P2_R1170_U153, P2_R1170_U154, P2_R1170_U155, P2_R1170_U156, P2_R1170_U157, P2_R1170_U158, P2_R1170_U159, P2_R1170_U16, P2_R1170_U160, P2_R1170_U161, P2_R1170_U162, P2_R1170_U163, P2_R1170_U164, P2_R1170_U165, P2_R1170_U166, P2_R1170_U167, P2_R1170_U168, P2_R1170_U169, P2_R1170_U17, P2_R1170_U170, P2_R1170_U171, P2_R1170_U172, P2_R1170_U173, P2_R1170_U174, P2_R1170_U175, P2_R1170_U176, P2_R1170_U177, P2_R1170_U178, P2_R1170_U179, P2_R1170_U18, P2_R1170_U180, P2_R1170_U181, P2_R1170_U182, P2_R1170_U183, P2_R1170_U184, P2_R1170_U185, P2_R1170_U186, P2_R1170_U187, P2_R1170_U188, P2_R1170_U189, P2_R1170_U19, P2_R1170_U190, P2_R1170_U191, P2_R1170_U192, P2_R1170_U193, P2_R1170_U194, P2_R1170_U195, P2_R1170_U196, P2_R1170_U197, P2_R1170_U198, P2_R1170_U199, P2_R1170_U20, P2_R1170_U200, P2_R1170_U201, P2_R1170_U202, P2_R1170_U203, P2_R1170_U204, P2_R1170_U205, P2_R1170_U206, P2_R1170_U207, P2_R1170_U208, P2_R1170_U209, P2_R1170_U21, P2_R1170_U210, P2_R1170_U211, P2_R1170_U212, P2_R1170_U213, P2_R1170_U214, P2_R1170_U215, P2_R1170_U216, P2_R1170_U217, P2_R1170_U218, P2_R1170_U219, P2_R1170_U22, P2_R1170_U220, P2_R1170_U221, P2_R1170_U222, P2_R1170_U223, P2_R1170_U224, P2_R1170_U225, P2_R1170_U226, P2_R1170_U227, P2_R1170_U228, P2_R1170_U229, P2_R1170_U23, P2_R1170_U230, P2_R1170_U231, P2_R1170_U232, P2_R1170_U233, P2_R1170_U234, P2_R1170_U235, P2_R1170_U236, P2_R1170_U237, P2_R1170_U238, P2_R1170_U239, P2_R1170_U24, P2_R1170_U240, P2_R1170_U241, P2_R1170_U242, P2_R1170_U243, P2_R1170_U244, P2_R1170_U245, P2_R1170_U246, P2_R1170_U247, P2_R1170_U248, P2_R1170_U249, P2_R1170_U25, P2_R1170_U250, P2_R1170_U251, P2_R1170_U252, P2_R1170_U253, P2_R1170_U254, P2_R1170_U255, P2_R1170_U256, P2_R1170_U257, P2_R1170_U258, P2_R1170_U259, P2_R1170_U26, P2_R1170_U260, P2_R1170_U261, P2_R1170_U262, P2_R1170_U263, P2_R1170_U264, P2_R1170_U265, P2_R1170_U266, P2_R1170_U267, P2_R1170_U268, P2_R1170_U269, P2_R1170_U27, P2_R1170_U270, P2_R1170_U271, P2_R1170_U272, P2_R1170_U273, P2_R1170_U274, P2_R1170_U275, P2_R1170_U276, P2_R1170_U277, P2_R1170_U278, P2_R1170_U279, P2_R1170_U28, P2_R1170_U280, P2_R1170_U281, P2_R1170_U282, P2_R1170_U283, P2_R1170_U284, P2_R1170_U285, P2_R1170_U286, P2_R1170_U287, P2_R1170_U288, P2_R1170_U289, P2_R1170_U29, P2_R1170_U290, P2_R1170_U291, P2_R1170_U292, P2_R1170_U293, P2_R1170_U294, P2_R1170_U295, P2_R1170_U296, P2_R1170_U297, P2_R1170_U298, P2_R1170_U299, P2_R1170_U30, P2_R1170_U300, P2_R1170_U301, P2_R1170_U302, P2_R1170_U303, P2_R1170_U304, P2_R1170_U305, P2_R1170_U306, P2_R1170_U307, P2_R1170_U308, P2_R1170_U31, P2_R1170_U32, P2_R1170_U33, P2_R1170_U34, P2_R1170_U35, P2_R1170_U36, P2_R1170_U37, P2_R1170_U38, P2_R1170_U39, P2_R1170_U4, P2_R1170_U40, P2_R1170_U41, P2_R1170_U42, P2_R1170_U43, P2_R1170_U44, P2_R1170_U45, P2_R1170_U46, P2_R1170_U47, P2_R1170_U48, P2_R1170_U49, P2_R1170_U5, P2_R1170_U50, P2_R1170_U51, P2_R1170_U52, P2_R1170_U53, P2_R1170_U54, P2_R1170_U55, P2_R1170_U56, P2_R1170_U57, P2_R1170_U58, P2_R1170_U59, P2_R1170_U6, P2_R1170_U60, P2_R1170_U61, P2_R1170_U62, P2_R1170_U63, P2_R1170_U64, P2_R1170_U65, P2_R1170_U66, P2_R1170_U67, P2_R1170_U68, P2_R1170_U69, P2_R1170_U7, P2_R1170_U70, P2_R1170_U71, P2_R1170_U72, P2_R1170_U73, P2_R1170_U74, P2_R1170_U75, P2_R1170_U76, P2_R1170_U77, P2_R1170_U78, P2_R1170_U79, P2_R1170_U8, P2_R1170_U80, P2_R1170_U81, P2_R1170_U82, P2_R1170_U83, P2_R1170_U84, P2_R1170_U85, P2_R1170_U86, P2_R1170_U87, P2_R1170_U88, P2_R1170_U89, P2_R1170_U9, P2_R1170_U90, P2_R1170_U91, P2_R1170_U92, P2_R1170_U93, P2_R1170_U94, P2_R1170_U95, P2_R1170_U96, P2_R1170_U97, P2_R1170_U98, P2_R1170_U99, P2_R1176_U10, P2_R1176_U100, P2_R1176_U101, P2_R1176_U102, P2_R1176_U103, P2_R1176_U104, P2_R1176_U105, P2_R1176_U106, P2_R1176_U107, P2_R1176_U108, P2_R1176_U109, P2_R1176_U11, P2_R1176_U110, P2_R1176_U111, P2_R1176_U112, P2_R1176_U113, P2_R1176_U114, P2_R1176_U115, P2_R1176_U116, P2_R1176_U117, P2_R1176_U118, P2_R1176_U119, P2_R1176_U12, P2_R1176_U120, P2_R1176_U121, P2_R1176_U122, P2_R1176_U123, P2_R1176_U124, P2_R1176_U125, P2_R1176_U126, P2_R1176_U127, P2_R1176_U128, P2_R1176_U129, P2_R1176_U13, P2_R1176_U130, P2_R1176_U131, P2_R1176_U132, P2_R1176_U133, P2_R1176_U134, P2_R1176_U135, P2_R1176_U136, P2_R1176_U137, P2_R1176_U138, P2_R1176_U139, P2_R1176_U14, P2_R1176_U140, P2_R1176_U141, P2_R1176_U142, P2_R1176_U143, P2_R1176_U144, P2_R1176_U145, P2_R1176_U146, P2_R1176_U147, P2_R1176_U148, P2_R1176_U149, P2_R1176_U15, P2_R1176_U150, P2_R1176_U151, P2_R1176_U152, P2_R1176_U153, P2_R1176_U154, P2_R1176_U155, P2_R1176_U156, P2_R1176_U157, P2_R1176_U158, P2_R1176_U159, P2_R1176_U16, P2_R1176_U160, P2_R1176_U161, P2_R1176_U162, P2_R1176_U163, P2_R1176_U164, P2_R1176_U165, P2_R1176_U166, P2_R1176_U167, P2_R1176_U168, P2_R1176_U169, P2_R1176_U17, P2_R1176_U170, P2_R1176_U171, P2_R1176_U172, P2_R1176_U173, P2_R1176_U174, P2_R1176_U175, P2_R1176_U176, P2_R1176_U177, P2_R1176_U178, P2_R1176_U179, P2_R1176_U18, P2_R1176_U180, P2_R1176_U181, P2_R1176_U182, P2_R1176_U183, P2_R1176_U184, P2_R1176_U185, P2_R1176_U186, P2_R1176_U187, P2_R1176_U188, P2_R1176_U189, P2_R1176_U19, P2_R1176_U190, P2_R1176_U191, P2_R1176_U192, P2_R1176_U193, P2_R1176_U194, P2_R1176_U195, P2_R1176_U196, P2_R1176_U197, P2_R1176_U198, P2_R1176_U199, P2_R1176_U20, P2_R1176_U200, P2_R1176_U201, P2_R1176_U202, P2_R1176_U203, P2_R1176_U204, P2_R1176_U205, P2_R1176_U206, P2_R1176_U207, P2_R1176_U208, P2_R1176_U209, P2_R1176_U21, P2_R1176_U210, P2_R1176_U211, P2_R1176_U212, P2_R1176_U213, P2_R1176_U214, P2_R1176_U215, P2_R1176_U216, P2_R1176_U217, P2_R1176_U218, P2_R1176_U219, P2_R1176_U22, P2_R1176_U220, P2_R1176_U221, P2_R1176_U222, P2_R1176_U223, P2_R1176_U224, P2_R1176_U225, P2_R1176_U226, P2_R1176_U227, P2_R1176_U228, P2_R1176_U229, P2_R1176_U23, P2_R1176_U230, P2_R1176_U231, P2_R1176_U232, P2_R1176_U233, P2_R1176_U234, P2_R1176_U235, P2_R1176_U236, P2_R1176_U237, P2_R1176_U238, P2_R1176_U239, P2_R1176_U24, P2_R1176_U240, P2_R1176_U241, P2_R1176_U242, P2_R1176_U243, P2_R1176_U244, P2_R1176_U245, P2_R1176_U246, P2_R1176_U247, P2_R1176_U248, P2_R1176_U249, P2_R1176_U25, P2_R1176_U250, P2_R1176_U251, P2_R1176_U252, P2_R1176_U253, P2_R1176_U254, P2_R1176_U255, P2_R1176_U256, P2_R1176_U257, P2_R1176_U258, P2_R1176_U259, P2_R1176_U26, P2_R1176_U260, P2_R1176_U261, P2_R1176_U262, P2_R1176_U263, P2_R1176_U264, P2_R1176_U265, P2_R1176_U266, P2_R1176_U267, P2_R1176_U268, P2_R1176_U269, P2_R1176_U27, P2_R1176_U270, P2_R1176_U271, P2_R1176_U272, P2_R1176_U273, P2_R1176_U274, P2_R1176_U275, P2_R1176_U276, P2_R1176_U277, P2_R1176_U278, P2_R1176_U279, P2_R1176_U28, P2_R1176_U280, P2_R1176_U281, P2_R1176_U282, P2_R1176_U283, P2_R1176_U284, P2_R1176_U285, P2_R1176_U286, P2_R1176_U287, P2_R1176_U288, P2_R1176_U289, P2_R1176_U29, P2_R1176_U290, P2_R1176_U291, P2_R1176_U292, P2_R1176_U293, P2_R1176_U294, P2_R1176_U295, P2_R1176_U296, P2_R1176_U297, P2_R1176_U298, P2_R1176_U299, P2_R1176_U30, P2_R1176_U300, P2_R1176_U301, P2_R1176_U302, P2_R1176_U303, P2_R1176_U304, P2_R1176_U305, P2_R1176_U306, P2_R1176_U307, P2_R1176_U308, P2_R1176_U309, P2_R1176_U31, P2_R1176_U310, P2_R1176_U311, P2_R1176_U312, P2_R1176_U313, P2_R1176_U314, P2_R1176_U315, P2_R1176_U316, P2_R1176_U317, P2_R1176_U318, P2_R1176_U319, P2_R1176_U32, P2_R1176_U320, P2_R1176_U321, P2_R1176_U322, P2_R1176_U323, P2_R1176_U324, P2_R1176_U325, P2_R1176_U326, P2_R1176_U327, P2_R1176_U328, P2_R1176_U329, P2_R1176_U33, P2_R1176_U330, P2_R1176_U331, P2_R1176_U332, P2_R1176_U333, P2_R1176_U334, P2_R1176_U335, P2_R1176_U336, P2_R1176_U337, P2_R1176_U338, P2_R1176_U339, P2_R1176_U34, P2_R1176_U340, P2_R1176_U341, P2_R1176_U342, P2_R1176_U343, P2_R1176_U344, P2_R1176_U345, P2_R1176_U346, P2_R1176_U347, P2_R1176_U348, P2_R1176_U349, P2_R1176_U35, P2_R1176_U350, P2_R1176_U351, P2_R1176_U352, P2_R1176_U353, P2_R1176_U354, P2_R1176_U355, P2_R1176_U356, P2_R1176_U357, P2_R1176_U358, P2_R1176_U359, P2_R1176_U36, P2_R1176_U360, P2_R1176_U361, P2_R1176_U362, P2_R1176_U363, P2_R1176_U364, P2_R1176_U365, P2_R1176_U366, P2_R1176_U367, P2_R1176_U368, P2_R1176_U369, P2_R1176_U37, P2_R1176_U370, P2_R1176_U371, P2_R1176_U372, P2_R1176_U373, P2_R1176_U374, P2_R1176_U375, P2_R1176_U376, P2_R1176_U377, P2_R1176_U378, P2_R1176_U379, P2_R1176_U38, P2_R1176_U380, P2_R1176_U381, P2_R1176_U382, P2_R1176_U383, P2_R1176_U384, P2_R1176_U385, P2_R1176_U386, P2_R1176_U387, P2_R1176_U388, P2_R1176_U389, P2_R1176_U39, P2_R1176_U390, P2_R1176_U391, P2_R1176_U392, P2_R1176_U393, P2_R1176_U394, P2_R1176_U395, P2_R1176_U396, P2_R1176_U397, P2_R1176_U398, P2_R1176_U399, P2_R1176_U4, P2_R1176_U40, P2_R1176_U400, P2_R1176_U401, P2_R1176_U402, P2_R1176_U403, P2_R1176_U404, P2_R1176_U405, P2_R1176_U406, P2_R1176_U407, P2_R1176_U408, P2_R1176_U409, P2_R1176_U41, P2_R1176_U410, P2_R1176_U411, P2_R1176_U412, P2_R1176_U413, P2_R1176_U414, P2_R1176_U415, P2_R1176_U416, P2_R1176_U417, P2_R1176_U418, P2_R1176_U419, P2_R1176_U42, P2_R1176_U420, P2_R1176_U421, P2_R1176_U422, P2_R1176_U423, P2_R1176_U424, P2_R1176_U425, P2_R1176_U426, P2_R1176_U427, P2_R1176_U428, P2_R1176_U429, P2_R1176_U43, P2_R1176_U430, P2_R1176_U431, P2_R1176_U432, P2_R1176_U433, P2_R1176_U434, P2_R1176_U435, P2_R1176_U436, P2_R1176_U437, P2_R1176_U438, P2_R1176_U439, P2_R1176_U44, P2_R1176_U440, P2_R1176_U441, P2_R1176_U442, P2_R1176_U443, P2_R1176_U444, P2_R1176_U445, P2_R1176_U446, P2_R1176_U447, P2_R1176_U448, P2_R1176_U449, P2_R1176_U45, P2_R1176_U450, P2_R1176_U451, P2_R1176_U452, P2_R1176_U453, P2_R1176_U454, P2_R1176_U455, P2_R1176_U456, P2_R1176_U457, P2_R1176_U458, P2_R1176_U459, P2_R1176_U46, P2_R1176_U460, P2_R1176_U461, P2_R1176_U462, P2_R1176_U463, P2_R1176_U464, P2_R1176_U465, P2_R1176_U466, P2_R1176_U467, P2_R1176_U468, P2_R1176_U469, P2_R1176_U47, P2_R1176_U470, P2_R1176_U471, P2_R1176_U472, P2_R1176_U473, P2_R1176_U474, P2_R1176_U475, P2_R1176_U476, P2_R1176_U477, P2_R1176_U478, P2_R1176_U479, P2_R1176_U48, P2_R1176_U480, P2_R1176_U481, P2_R1176_U482, P2_R1176_U483, P2_R1176_U484, P2_R1176_U485, P2_R1176_U486, P2_R1176_U487, P2_R1176_U488, P2_R1176_U489, P2_R1176_U49, P2_R1176_U490, P2_R1176_U491, P2_R1176_U492, P2_R1176_U493, P2_R1176_U494, P2_R1176_U495, P2_R1176_U496, P2_R1176_U497, P2_R1176_U498, P2_R1176_U499, P2_R1176_U5, P2_R1176_U50, P2_R1176_U500, P2_R1176_U501, P2_R1176_U502, P2_R1176_U503, P2_R1176_U504, P2_R1176_U505, P2_R1176_U506, P2_R1176_U507, P2_R1176_U508, P2_R1176_U509, P2_R1176_U51, P2_R1176_U510, P2_R1176_U511, P2_R1176_U512, P2_R1176_U513, P2_R1176_U514, P2_R1176_U515, P2_R1176_U516, P2_R1176_U517, P2_R1176_U518, P2_R1176_U519, P2_R1176_U52, P2_R1176_U520, P2_R1176_U521, P2_R1176_U522, P2_R1176_U523, P2_R1176_U524, P2_R1176_U525, P2_R1176_U526, P2_R1176_U527, P2_R1176_U528, P2_R1176_U529, P2_R1176_U53, P2_R1176_U530, P2_R1176_U531, P2_R1176_U532, P2_R1176_U533, P2_R1176_U534, P2_R1176_U535, P2_R1176_U536, P2_R1176_U537, P2_R1176_U538, P2_R1176_U539, P2_R1176_U54, P2_R1176_U540, P2_R1176_U541, P2_R1176_U542, P2_R1176_U543, P2_R1176_U544, P2_R1176_U545, P2_R1176_U546, P2_R1176_U547, P2_R1176_U548, P2_R1176_U549, P2_R1176_U55, P2_R1176_U550, P2_R1176_U551, P2_R1176_U552, P2_R1176_U553, P2_R1176_U554, P2_R1176_U555, P2_R1176_U556, P2_R1176_U557, P2_R1176_U558, P2_R1176_U559, P2_R1176_U56, P2_R1176_U560, P2_R1176_U561, P2_R1176_U562, P2_R1176_U563, P2_R1176_U564, P2_R1176_U565, P2_R1176_U566, P2_R1176_U567, P2_R1176_U568, P2_R1176_U569, P2_R1176_U57, P2_R1176_U570, P2_R1176_U571, P2_R1176_U572, P2_R1176_U573, P2_R1176_U574, P2_R1176_U575, P2_R1176_U576, P2_R1176_U577, P2_R1176_U578, P2_R1176_U579, P2_R1176_U58, P2_R1176_U580, P2_R1176_U581, P2_R1176_U582, P2_R1176_U583, P2_R1176_U584, P2_R1176_U585, P2_R1176_U586, P2_R1176_U587, P2_R1176_U588, P2_R1176_U589, P2_R1176_U59, P2_R1176_U590, P2_R1176_U591, P2_R1176_U592, P2_R1176_U593, P2_R1176_U594, P2_R1176_U595, P2_R1176_U596, P2_R1176_U597, P2_R1176_U598, P2_R1176_U599, P2_R1176_U6, P2_R1176_U60, P2_R1176_U600, P2_R1176_U601, P2_R1176_U602, P2_R1176_U603, P2_R1176_U604, P2_R1176_U605, P2_R1176_U606, P2_R1176_U607, P2_R1176_U608, P2_R1176_U609, P2_R1176_U61, P2_R1176_U610, P2_R1176_U611, P2_R1176_U612, P2_R1176_U613, P2_R1176_U614, P2_R1176_U615, P2_R1176_U616, P2_R1176_U617, P2_R1176_U618, P2_R1176_U619, P2_R1176_U62, P2_R1176_U620, P2_R1176_U621, P2_R1176_U622, P2_R1176_U623, P2_R1176_U63, P2_R1176_U64, P2_R1176_U65, P2_R1176_U66, P2_R1176_U67, P2_R1176_U68, P2_R1176_U69, P2_R1176_U7, P2_R1176_U70, P2_R1176_U71, P2_R1176_U72, P2_R1176_U73, P2_R1176_U74, P2_R1176_U75, P2_R1176_U76, P2_R1176_U77, P2_R1176_U78, P2_R1176_U79, P2_R1176_U8, P2_R1176_U80, P2_R1176_U81, P2_R1176_U82, P2_R1176_U83, P2_R1176_U84, P2_R1176_U85, P2_R1176_U86, P2_R1176_U87, P2_R1176_U88, P2_R1176_U89, P2_R1176_U9, P2_R1176_U90, P2_R1176_U91, P2_R1176_U92, P2_R1176_U93, P2_R1176_U94, P2_R1176_U95, P2_R1176_U96, P2_R1176_U97, P2_R1176_U98, P2_R1176_U99, P2_R1179_U10, P2_R1179_U100, P2_R1179_U101, P2_R1179_U102, P2_R1179_U103, P2_R1179_U104, P2_R1179_U105, P2_R1179_U106, P2_R1179_U107, P2_R1179_U108, P2_R1179_U109, P2_R1179_U11, P2_R1179_U110, P2_R1179_U111, P2_R1179_U112, P2_R1179_U113, P2_R1179_U114, P2_R1179_U115, P2_R1179_U116, P2_R1179_U117, P2_R1179_U118, P2_R1179_U119, P2_R1179_U12, P2_R1179_U120, P2_R1179_U121, P2_R1179_U122, P2_R1179_U123, P2_R1179_U124, P2_R1179_U125, P2_R1179_U126, P2_R1179_U127, P2_R1179_U128, P2_R1179_U129, P2_R1179_U13, P2_R1179_U130, P2_R1179_U131, P2_R1179_U132, P2_R1179_U133, P2_R1179_U134, P2_R1179_U135, P2_R1179_U136, P2_R1179_U137, P2_R1179_U138, P2_R1179_U139, P2_R1179_U14, P2_R1179_U140, P2_R1179_U141, P2_R1179_U142, P2_R1179_U143, P2_R1179_U144, P2_R1179_U145, P2_R1179_U146, P2_R1179_U147, P2_R1179_U148, P2_R1179_U149, P2_R1179_U15, P2_R1179_U150, P2_R1179_U151, P2_R1179_U152, P2_R1179_U153, P2_R1179_U154, P2_R1179_U155, P2_R1179_U156, P2_R1179_U157, P2_R1179_U158, P2_R1179_U159, P2_R1179_U16, P2_R1179_U160, P2_R1179_U161, P2_R1179_U162, P2_R1179_U163, P2_R1179_U164, P2_R1179_U165, P2_R1179_U166, P2_R1179_U167, P2_R1179_U168, P2_R1179_U169, P2_R1179_U17, P2_R1179_U170, P2_R1179_U171, P2_R1179_U172, P2_R1179_U173, P2_R1179_U174, P2_R1179_U175, P2_R1179_U176, P2_R1179_U177, P2_R1179_U178, P2_R1179_U179, P2_R1179_U18, P2_R1179_U180, P2_R1179_U181, P2_R1179_U182, P2_R1179_U183, P2_R1179_U184, P2_R1179_U185, P2_R1179_U186, P2_R1179_U187, P2_R1179_U188, P2_R1179_U189, P2_R1179_U19, P2_R1179_U190, P2_R1179_U191, P2_R1179_U192, P2_R1179_U193, P2_R1179_U194, P2_R1179_U195, P2_R1179_U196, P2_R1179_U197, P2_R1179_U198, P2_R1179_U199, P2_R1179_U20, P2_R1179_U200, P2_R1179_U201, P2_R1179_U202, P2_R1179_U203, P2_R1179_U204, P2_R1179_U205, P2_R1179_U206, P2_R1179_U207, P2_R1179_U208, P2_R1179_U209, P2_R1179_U21, P2_R1179_U210, P2_R1179_U211, P2_R1179_U212, P2_R1179_U213, P2_R1179_U214, P2_R1179_U215, P2_R1179_U216, P2_R1179_U217, P2_R1179_U218, P2_R1179_U219, P2_R1179_U22, P2_R1179_U220, P2_R1179_U221, P2_R1179_U222, P2_R1179_U223, P2_R1179_U224, P2_R1179_U225, P2_R1179_U226, P2_R1179_U227, P2_R1179_U228, P2_R1179_U229, P2_R1179_U23, P2_R1179_U230, P2_R1179_U231, P2_R1179_U232, P2_R1179_U233, P2_R1179_U234, P2_R1179_U235, P2_R1179_U236, P2_R1179_U237, P2_R1179_U238, P2_R1179_U239, P2_R1179_U24, P2_R1179_U240, P2_R1179_U241, P2_R1179_U242, P2_R1179_U243, P2_R1179_U244, P2_R1179_U245, P2_R1179_U246, P2_R1179_U247, P2_R1179_U248, P2_R1179_U249, P2_R1179_U25, P2_R1179_U250, P2_R1179_U251, P2_R1179_U252, P2_R1179_U253, P2_R1179_U254, P2_R1179_U255, P2_R1179_U256, P2_R1179_U257, P2_R1179_U258, P2_R1179_U259, P2_R1179_U26, P2_R1179_U260, P2_R1179_U261, P2_R1179_U262, P2_R1179_U263, P2_R1179_U264, P2_R1179_U265, P2_R1179_U266, P2_R1179_U267, P2_R1179_U268, P2_R1179_U269, P2_R1179_U27, P2_R1179_U270, P2_R1179_U271, P2_R1179_U272, P2_R1179_U273, P2_R1179_U274, P2_R1179_U275, P2_R1179_U276, P2_R1179_U277, P2_R1179_U278, P2_R1179_U279, P2_R1179_U28, P2_R1179_U280, P2_R1179_U281, P2_R1179_U282, P2_R1179_U283, P2_R1179_U284, P2_R1179_U285, P2_R1179_U286, P2_R1179_U287, P2_R1179_U288, P2_R1179_U289, P2_R1179_U29, P2_R1179_U290, P2_R1179_U291, P2_R1179_U292, P2_R1179_U293, P2_R1179_U294, P2_R1179_U295, P2_R1179_U296, P2_R1179_U297, P2_R1179_U298, P2_R1179_U299, P2_R1179_U30, P2_R1179_U300, P2_R1179_U301, P2_R1179_U302, P2_R1179_U303, P2_R1179_U304, P2_R1179_U305, P2_R1179_U306, P2_R1179_U307, P2_R1179_U308, P2_R1179_U309, P2_R1179_U31, P2_R1179_U310, P2_R1179_U311, P2_R1179_U312, P2_R1179_U313, P2_R1179_U314, P2_R1179_U315, P2_R1179_U316, P2_R1179_U317, P2_R1179_U318, P2_R1179_U319, P2_R1179_U32, P2_R1179_U320, P2_R1179_U321, P2_R1179_U322, P2_R1179_U323, P2_R1179_U324, P2_R1179_U325, P2_R1179_U326, P2_R1179_U327, P2_R1179_U328, P2_R1179_U329, P2_R1179_U33, P2_R1179_U330, P2_R1179_U331, P2_R1179_U332, P2_R1179_U333, P2_R1179_U334, P2_R1179_U335, P2_R1179_U336, P2_R1179_U337, P2_R1179_U338, P2_R1179_U339, P2_R1179_U34, P2_R1179_U340, P2_R1179_U341, P2_R1179_U342, P2_R1179_U343, P2_R1179_U344, P2_R1179_U345, P2_R1179_U346, P2_R1179_U347, P2_R1179_U348, P2_R1179_U349, P2_R1179_U35, P2_R1179_U350, P2_R1179_U351, P2_R1179_U352, P2_R1179_U353, P2_R1179_U354, P2_R1179_U355, P2_R1179_U356, P2_R1179_U357, P2_R1179_U358, P2_R1179_U359, P2_R1179_U36, P2_R1179_U360, P2_R1179_U361, P2_R1179_U362, P2_R1179_U363, P2_R1179_U364, P2_R1179_U365, P2_R1179_U366, P2_R1179_U367, P2_R1179_U368, P2_R1179_U369, P2_R1179_U37, P2_R1179_U370, P2_R1179_U371, P2_R1179_U372, P2_R1179_U373, P2_R1179_U374, P2_R1179_U375, P2_R1179_U376, P2_R1179_U377, P2_R1179_U378, P2_R1179_U379, P2_R1179_U38, P2_R1179_U380, P2_R1179_U381, P2_R1179_U382, P2_R1179_U383, P2_R1179_U384, P2_R1179_U385, P2_R1179_U386, P2_R1179_U387, P2_R1179_U388, P2_R1179_U389, P2_R1179_U39, P2_R1179_U390, P2_R1179_U391, P2_R1179_U392, P2_R1179_U393, P2_R1179_U394, P2_R1179_U395, P2_R1179_U396, P2_R1179_U397, P2_R1179_U398, P2_R1179_U399, P2_R1179_U40, P2_R1179_U400, P2_R1179_U401, P2_R1179_U402, P2_R1179_U403, P2_R1179_U404, P2_R1179_U405, P2_R1179_U406, P2_R1179_U407, P2_R1179_U408, P2_R1179_U409, P2_R1179_U41, P2_R1179_U410, P2_R1179_U411, P2_R1179_U412, P2_R1179_U413, P2_R1179_U414, P2_R1179_U415, P2_R1179_U416, P2_R1179_U417, P2_R1179_U418, P2_R1179_U419, P2_R1179_U42, P2_R1179_U420, P2_R1179_U421, P2_R1179_U422, P2_R1179_U423, P2_R1179_U424, P2_R1179_U425, P2_R1179_U426, P2_R1179_U427, P2_R1179_U428, P2_R1179_U429, P2_R1179_U43, P2_R1179_U430, P2_R1179_U431, P2_R1179_U432, P2_R1179_U433, P2_R1179_U434, P2_R1179_U435, P2_R1179_U436, P2_R1179_U437, P2_R1179_U438, P2_R1179_U439, P2_R1179_U44, P2_R1179_U440, P2_R1179_U441, P2_R1179_U442, P2_R1179_U443, P2_R1179_U444, P2_R1179_U445, P2_R1179_U446, P2_R1179_U447, P2_R1179_U448, P2_R1179_U449, P2_R1179_U45, P2_R1179_U450, P2_R1179_U451, P2_R1179_U452, P2_R1179_U453, P2_R1179_U454, P2_R1179_U455, P2_R1179_U456, P2_R1179_U457, P2_R1179_U458, P2_R1179_U459, P2_R1179_U46, P2_R1179_U460, P2_R1179_U461, P2_R1179_U462, P2_R1179_U463, P2_R1179_U464, P2_R1179_U465, P2_R1179_U466, P2_R1179_U467, P2_R1179_U468, P2_R1179_U469, P2_R1179_U47, P2_R1179_U470, P2_R1179_U471, P2_R1179_U472, P2_R1179_U473, P2_R1179_U474, P2_R1179_U475, P2_R1179_U476, P2_R1179_U477, P2_R1179_U478, P2_R1179_U48, P2_R1179_U49, P2_R1179_U50, P2_R1179_U51, P2_R1179_U52, P2_R1179_U53, P2_R1179_U54, P2_R1179_U55, P2_R1179_U56, P2_R1179_U57, P2_R1179_U58, P2_R1179_U59, P2_R1179_U6, P2_R1179_U60, P2_R1179_U61, P2_R1179_U62, P2_R1179_U63, P2_R1179_U64, P2_R1179_U65, P2_R1179_U66, P2_R1179_U67, P2_R1179_U68, P2_R1179_U69, P2_R1179_U7, P2_R1179_U70, P2_R1179_U71, P2_R1179_U72, P2_R1179_U73, P2_R1179_U74, P2_R1179_U75, P2_R1179_U76, P2_R1179_U77, P2_R1179_U78, P2_R1179_U79, P2_R1179_U8, P2_R1179_U80, P2_R1179_U81, P2_R1179_U82, P2_R1179_U83, P2_R1179_U84, P2_R1179_U85, P2_R1179_U86, P2_R1179_U87, P2_R1179_U88, P2_R1179_U89, P2_R1179_U9, P2_R1179_U90, P2_R1179_U91, P2_R1179_U92, P2_R1179_U93, P2_R1179_U94, P2_R1179_U95, P2_R1179_U96, P2_R1179_U97, P2_R1179_U98, P2_R1179_U99, P2_R1203_U10, P2_R1203_U100, P2_R1203_U101, P2_R1203_U102, P2_R1203_U103, P2_R1203_U104, P2_R1203_U105, P2_R1203_U106, P2_R1203_U107, P2_R1203_U108, P2_R1203_U109, P2_R1203_U11, P2_R1203_U110, P2_R1203_U111, P2_R1203_U112, P2_R1203_U113, P2_R1203_U114, P2_R1203_U115, P2_R1203_U116, P2_R1203_U117, P2_R1203_U118, P2_R1203_U119, P2_R1203_U12, P2_R1203_U120, P2_R1203_U121, P2_R1203_U122, P2_R1203_U123, P2_R1203_U124, P2_R1203_U125, P2_R1203_U126, P2_R1203_U127, P2_R1203_U128, P2_R1203_U129, P2_R1203_U13, P2_R1203_U130, P2_R1203_U131, P2_R1203_U132, P2_R1203_U133, P2_R1203_U134, P2_R1203_U135, P2_R1203_U136, P2_R1203_U137, P2_R1203_U138, P2_R1203_U139, P2_R1203_U14, P2_R1203_U140, P2_R1203_U141, P2_R1203_U142, P2_R1203_U143, P2_R1203_U144, P2_R1203_U145, P2_R1203_U146, P2_R1203_U147, P2_R1203_U148, P2_R1203_U149, P2_R1203_U15, P2_R1203_U150, P2_R1203_U151, P2_R1203_U152, P2_R1203_U153, P2_R1203_U154, P2_R1203_U155, P2_R1203_U156, P2_R1203_U157, P2_R1203_U158, P2_R1203_U159, P2_R1203_U16, P2_R1203_U160, P2_R1203_U161, P2_R1203_U162, P2_R1203_U163, P2_R1203_U164, P2_R1203_U165, P2_R1203_U166, P2_R1203_U167, P2_R1203_U168, P2_R1203_U169, P2_R1203_U17, P2_R1203_U170, P2_R1203_U171, P2_R1203_U172, P2_R1203_U173, P2_R1203_U174, P2_R1203_U175, P2_R1203_U176, P2_R1203_U177, P2_R1203_U178, P2_R1203_U179, P2_R1203_U18, P2_R1203_U180, P2_R1203_U181, P2_R1203_U182, P2_R1203_U183, P2_R1203_U184, P2_R1203_U185, P2_R1203_U186, P2_R1203_U187, P2_R1203_U188, P2_R1203_U189, P2_R1203_U19, P2_R1203_U190, P2_R1203_U191, P2_R1203_U192, P2_R1203_U193, P2_R1203_U194, P2_R1203_U195, P2_R1203_U196, P2_R1203_U197, P2_R1203_U198, P2_R1203_U199, P2_R1203_U20, P2_R1203_U200, P2_R1203_U201, P2_R1203_U202, P2_R1203_U203, P2_R1203_U204, P2_R1203_U205, P2_R1203_U206, P2_R1203_U207, P2_R1203_U208, P2_R1203_U209, P2_R1203_U21, P2_R1203_U210, P2_R1203_U211, P2_R1203_U212, P2_R1203_U213, P2_R1203_U214, P2_R1203_U215, P2_R1203_U216, P2_R1203_U217, P2_R1203_U218, P2_R1203_U219, P2_R1203_U22, P2_R1203_U220, P2_R1203_U221, P2_R1203_U222, P2_R1203_U223, P2_R1203_U224, P2_R1203_U225, P2_R1203_U226, P2_R1203_U227, P2_R1203_U228, P2_R1203_U229, P2_R1203_U23, P2_R1203_U230, P2_R1203_U231, P2_R1203_U232, P2_R1203_U233, P2_R1203_U234, P2_R1203_U235, P2_R1203_U236, P2_R1203_U237, P2_R1203_U238, P2_R1203_U239, P2_R1203_U24, P2_R1203_U240, P2_R1203_U241, P2_R1203_U242, P2_R1203_U243, P2_R1203_U244, P2_R1203_U245, P2_R1203_U246, P2_R1203_U247, P2_R1203_U248, P2_R1203_U249, P2_R1203_U25, P2_R1203_U250, P2_R1203_U251, P2_R1203_U252, P2_R1203_U253, P2_R1203_U254, P2_R1203_U255, P2_R1203_U256, P2_R1203_U257, P2_R1203_U258, P2_R1203_U259, P2_R1203_U26, P2_R1203_U260, P2_R1203_U261, P2_R1203_U262, P2_R1203_U263, P2_R1203_U264, P2_R1203_U265, P2_R1203_U266, P2_R1203_U267, P2_R1203_U268, P2_R1203_U269, P2_R1203_U27, P2_R1203_U270, P2_R1203_U271, P2_R1203_U272, P2_R1203_U273, P2_R1203_U274, P2_R1203_U275, P2_R1203_U276, P2_R1203_U277, P2_R1203_U278, P2_R1203_U279, P2_R1203_U28, P2_R1203_U280, P2_R1203_U281, P2_R1203_U282, P2_R1203_U283, P2_R1203_U284, P2_R1203_U285, P2_R1203_U286, P2_R1203_U287, P2_R1203_U288, P2_R1203_U289, P2_R1203_U29, P2_R1203_U290, P2_R1203_U291, P2_R1203_U292, P2_R1203_U293, P2_R1203_U294, P2_R1203_U295, P2_R1203_U296, P2_R1203_U297, P2_R1203_U298, P2_R1203_U299, P2_R1203_U30, P2_R1203_U300, P2_R1203_U301, P2_R1203_U302, P2_R1203_U303, P2_R1203_U304, P2_R1203_U305, P2_R1203_U306, P2_R1203_U307, P2_R1203_U308, P2_R1203_U309, P2_R1203_U31, P2_R1203_U310, P2_R1203_U311, P2_R1203_U312, P2_R1203_U313, P2_R1203_U314, P2_R1203_U315, P2_R1203_U316, P2_R1203_U317, P2_R1203_U318, P2_R1203_U319, P2_R1203_U32, P2_R1203_U320, P2_R1203_U321, P2_R1203_U322, P2_R1203_U323, P2_R1203_U324, P2_R1203_U325, P2_R1203_U326, P2_R1203_U327, P2_R1203_U328, P2_R1203_U329, P2_R1203_U33, P2_R1203_U330, P2_R1203_U331, P2_R1203_U332, P2_R1203_U333, P2_R1203_U334, P2_R1203_U335, P2_R1203_U336, P2_R1203_U337, P2_R1203_U338, P2_R1203_U339, P2_R1203_U34, P2_R1203_U340, P2_R1203_U341, P2_R1203_U342, P2_R1203_U343, P2_R1203_U344, P2_R1203_U345, P2_R1203_U346, P2_R1203_U347, P2_R1203_U348, P2_R1203_U349, P2_R1203_U35, P2_R1203_U350, P2_R1203_U351, P2_R1203_U352, P2_R1203_U353, P2_R1203_U354, P2_R1203_U355, P2_R1203_U356, P2_R1203_U357, P2_R1203_U358, P2_R1203_U359, P2_R1203_U36, P2_R1203_U360, P2_R1203_U361, P2_R1203_U362, P2_R1203_U363, P2_R1203_U364, P2_R1203_U365, P2_R1203_U366, P2_R1203_U367, P2_R1203_U368, P2_R1203_U369, P2_R1203_U37, P2_R1203_U370, P2_R1203_U371, P2_R1203_U372, P2_R1203_U373, P2_R1203_U374, P2_R1203_U375, P2_R1203_U376, P2_R1203_U377, P2_R1203_U378, P2_R1203_U379, P2_R1203_U38, P2_R1203_U380, P2_R1203_U381, P2_R1203_U382, P2_R1203_U383, P2_R1203_U384, P2_R1203_U385, P2_R1203_U386, P2_R1203_U387, P2_R1203_U388, P2_R1203_U389, P2_R1203_U39, P2_R1203_U390, P2_R1203_U391, P2_R1203_U392, P2_R1203_U393, P2_R1203_U394, P2_R1203_U395, P2_R1203_U396, P2_R1203_U397, P2_R1203_U398, P2_R1203_U399, P2_R1203_U40, P2_R1203_U400, P2_R1203_U401, P2_R1203_U402, P2_R1203_U403, P2_R1203_U404, P2_R1203_U405, P2_R1203_U406, P2_R1203_U407, P2_R1203_U408, P2_R1203_U409, P2_R1203_U41, P2_R1203_U410, P2_R1203_U411, P2_R1203_U412, P2_R1203_U413, P2_R1203_U414, P2_R1203_U415, P2_R1203_U416, P2_R1203_U417, P2_R1203_U418, P2_R1203_U419, P2_R1203_U42, P2_R1203_U420, P2_R1203_U421, P2_R1203_U422, P2_R1203_U423, P2_R1203_U424, P2_R1203_U425, P2_R1203_U426, P2_R1203_U427, P2_R1203_U428, P2_R1203_U429, P2_R1203_U43, P2_R1203_U430, P2_R1203_U431, P2_R1203_U432, P2_R1203_U433, P2_R1203_U434, P2_R1203_U435, P2_R1203_U436, P2_R1203_U437, P2_R1203_U438, P2_R1203_U439, P2_R1203_U44, P2_R1203_U440, P2_R1203_U441, P2_R1203_U442, P2_R1203_U443, P2_R1203_U444, P2_R1203_U445, P2_R1203_U446, P2_R1203_U447, P2_R1203_U448, P2_R1203_U449, P2_R1203_U45, P2_R1203_U450, P2_R1203_U451, P2_R1203_U452, P2_R1203_U453, P2_R1203_U454, P2_R1203_U455, P2_R1203_U456, P2_R1203_U457, P2_R1203_U458, P2_R1203_U459, P2_R1203_U46, P2_R1203_U460, P2_R1203_U461, P2_R1203_U462, P2_R1203_U463, P2_R1203_U464, P2_R1203_U465, P2_R1203_U466, P2_R1203_U467, P2_R1203_U468, P2_R1203_U469, P2_R1203_U47, P2_R1203_U470, P2_R1203_U471, P2_R1203_U472, P2_R1203_U473, P2_R1203_U474, P2_R1203_U475, P2_R1203_U476, P2_R1203_U477, P2_R1203_U478, P2_R1203_U48, P2_R1203_U49, P2_R1203_U50, P2_R1203_U51, P2_R1203_U52, P2_R1203_U53, P2_R1203_U54, P2_R1203_U55, P2_R1203_U56, P2_R1203_U57, P2_R1203_U58, P2_R1203_U59, P2_R1203_U6, P2_R1203_U60, P2_R1203_U61, P2_R1203_U62, P2_R1203_U63, P2_R1203_U64, P2_R1203_U65, P2_R1203_U66, P2_R1203_U67, P2_R1203_U68, P2_R1203_U69, P2_R1203_U7, P2_R1203_U70, P2_R1203_U71, P2_R1203_U72, P2_R1203_U73, P2_R1203_U74, P2_R1203_U75, P2_R1203_U76, P2_R1203_U77, P2_R1203_U78, P2_R1203_U79, P2_R1203_U8, P2_R1203_U80, P2_R1203_U81, P2_R1203_U82, P2_R1203_U83, P2_R1203_U84, P2_R1203_U85, P2_R1203_U86, P2_R1203_U87, P2_R1203_U88, P2_R1203_U89, P2_R1203_U9, P2_R1203_U90, P2_R1203_U91, P2_R1203_U92, P2_R1203_U93, P2_R1203_U94, P2_R1203_U95, P2_R1203_U96, P2_R1203_U97, P2_R1203_U98, P2_R1203_U99, P2_R1209_U10, P2_R1209_U100, P2_R1209_U101, P2_R1209_U102, P2_R1209_U103, P2_R1209_U104, P2_R1209_U105, P2_R1209_U106, P2_R1209_U107, P2_R1209_U108, P2_R1209_U109, P2_R1209_U11, P2_R1209_U110, P2_R1209_U111, P2_R1209_U112, P2_R1209_U113, P2_R1209_U114, P2_R1209_U115, P2_R1209_U116, P2_R1209_U117, P2_R1209_U118, P2_R1209_U119, P2_R1209_U12, P2_R1209_U120, P2_R1209_U121, P2_R1209_U122, P2_R1209_U123, P2_R1209_U124, P2_R1209_U125, P2_R1209_U126, P2_R1209_U127, P2_R1209_U128, P2_R1209_U129, P2_R1209_U13, P2_R1209_U130, P2_R1209_U131, P2_R1209_U132, P2_R1209_U133, P2_R1209_U134, P2_R1209_U135, P2_R1209_U136, P2_R1209_U137, P2_R1209_U138, P2_R1209_U139, P2_R1209_U14, P2_R1209_U140, P2_R1209_U141, P2_R1209_U142, P2_R1209_U143, P2_R1209_U144, P2_R1209_U145, P2_R1209_U146, P2_R1209_U147, P2_R1209_U148, P2_R1209_U149, P2_R1209_U15, P2_R1209_U150, P2_R1209_U151, P2_R1209_U152, P2_R1209_U153, P2_R1209_U154, P2_R1209_U155, P2_R1209_U156, P2_R1209_U157, P2_R1209_U158, P2_R1209_U159, P2_R1209_U16, P2_R1209_U160, P2_R1209_U161, P2_R1209_U162, P2_R1209_U163, P2_R1209_U164, P2_R1209_U165, P2_R1209_U166, P2_R1209_U167, P2_R1209_U168, P2_R1209_U169, P2_R1209_U17, P2_R1209_U170, P2_R1209_U171, P2_R1209_U172, P2_R1209_U173, P2_R1209_U174, P2_R1209_U175, P2_R1209_U176, P2_R1209_U177, P2_R1209_U178, P2_R1209_U179, P2_R1209_U18, P2_R1209_U180, P2_R1209_U181, P2_R1209_U182, P2_R1209_U183, P2_R1209_U184, P2_R1209_U185, P2_R1209_U186, P2_R1209_U187, P2_R1209_U188, P2_R1209_U189, P2_R1209_U19, P2_R1209_U190, P2_R1209_U191, P2_R1209_U192, P2_R1209_U193, P2_R1209_U194, P2_R1209_U195, P2_R1209_U196, P2_R1209_U197, P2_R1209_U198, P2_R1209_U199, P2_R1209_U20, P2_R1209_U200, P2_R1209_U201, P2_R1209_U202, P2_R1209_U203, P2_R1209_U204, P2_R1209_U205, P2_R1209_U206, P2_R1209_U207, P2_R1209_U208, P2_R1209_U209, P2_R1209_U21, P2_R1209_U210, P2_R1209_U211, P2_R1209_U212, P2_R1209_U213, P2_R1209_U214, P2_R1209_U215, P2_R1209_U216, P2_R1209_U217, P2_R1209_U218, P2_R1209_U219, P2_R1209_U22, P2_R1209_U220, P2_R1209_U221, P2_R1209_U222, P2_R1209_U223, P2_R1209_U224, P2_R1209_U225, P2_R1209_U226, P2_R1209_U227, P2_R1209_U228, P2_R1209_U229, P2_R1209_U23, P2_R1209_U230, P2_R1209_U231, P2_R1209_U232, P2_R1209_U233, P2_R1209_U234, P2_R1209_U235, P2_R1209_U236, P2_R1209_U237, P2_R1209_U238, P2_R1209_U239, P2_R1209_U24, P2_R1209_U240, P2_R1209_U241, P2_R1209_U242, P2_R1209_U243, P2_R1209_U244, P2_R1209_U245, P2_R1209_U246, P2_R1209_U247, P2_R1209_U248, P2_R1209_U249, P2_R1209_U25, P2_R1209_U250, P2_R1209_U251, P2_R1209_U252, P2_R1209_U253, P2_R1209_U254, P2_R1209_U255, P2_R1209_U256, P2_R1209_U257, P2_R1209_U258, P2_R1209_U259, P2_R1209_U26, P2_R1209_U260, P2_R1209_U261, P2_R1209_U262, P2_R1209_U263, P2_R1209_U264, P2_R1209_U265, P2_R1209_U266, P2_R1209_U267, P2_R1209_U268, P2_R1209_U269, P2_R1209_U27, P2_R1209_U270, P2_R1209_U271, P2_R1209_U272, P2_R1209_U273, P2_R1209_U274, P2_R1209_U275, P2_R1209_U276, P2_R1209_U277, P2_R1209_U278, P2_R1209_U279, P2_R1209_U28, P2_R1209_U280, P2_R1209_U281, P2_R1209_U282, P2_R1209_U283, P2_R1209_U284, P2_R1209_U285, P2_R1209_U286, P2_R1209_U287, P2_R1209_U288, P2_R1209_U289, P2_R1209_U29, P2_R1209_U290, P2_R1209_U291, P2_R1209_U292, P2_R1209_U293, P2_R1209_U294, P2_R1209_U295, P2_R1209_U296, P2_R1209_U297, P2_R1209_U298, P2_R1209_U299, P2_R1209_U30, P2_R1209_U300, P2_R1209_U301, P2_R1209_U302, P2_R1209_U303, P2_R1209_U304, P2_R1209_U305, P2_R1209_U306, P2_R1209_U307, P2_R1209_U308, P2_R1209_U31, P2_R1209_U32, P2_R1209_U33, P2_R1209_U34, P2_R1209_U35, P2_R1209_U36, P2_R1209_U37, P2_R1209_U38, P2_R1209_U39, P2_R1209_U4, P2_R1209_U40, P2_R1209_U41, P2_R1209_U42, P2_R1209_U43, P2_R1209_U44, P2_R1209_U45, P2_R1209_U46, P2_R1209_U47, P2_R1209_U48, P2_R1209_U49, P2_R1209_U5, P2_R1209_U50, P2_R1209_U51, P2_R1209_U52, P2_R1209_U53, P2_R1209_U54, P2_R1209_U55, P2_R1209_U56, P2_R1209_U57, P2_R1209_U58, P2_R1209_U59, P2_R1209_U6, P2_R1209_U60, P2_R1209_U61, P2_R1209_U62, P2_R1209_U63, P2_R1209_U64, P2_R1209_U65, P2_R1209_U66, P2_R1209_U67, P2_R1209_U68, P2_R1209_U69, P2_R1209_U7, P2_R1209_U70, P2_R1209_U71, P2_R1209_U72, P2_R1209_U73, P2_R1209_U74, P2_R1209_U75, P2_R1209_U76, P2_R1209_U77, P2_R1209_U78, P2_R1209_U79, P2_R1209_U8, P2_R1209_U80, P2_R1209_U81, P2_R1209_U82, P2_R1209_U83, P2_R1209_U84, P2_R1209_U85, P2_R1209_U86, P2_R1209_U87, P2_R1209_U88, P2_R1209_U89, P2_R1209_U9, P2_R1209_U90, P2_R1209_U91, P2_R1209_U92, P2_R1209_U93, P2_R1209_U94, P2_R1209_U95, P2_R1209_U96, P2_R1209_U97, P2_R1209_U98, P2_R1209_U99, P2_R1215_U10, P2_R1215_U100, P2_R1215_U101, P2_R1215_U102, P2_R1215_U103, P2_R1215_U104, P2_R1215_U105, P2_R1215_U106, P2_R1215_U107, P2_R1215_U108, P2_R1215_U109, P2_R1215_U11, P2_R1215_U110, P2_R1215_U111, P2_R1215_U112, P2_R1215_U113, P2_R1215_U114, P2_R1215_U115, P2_R1215_U116, P2_R1215_U117, P2_R1215_U118, P2_R1215_U119, P2_R1215_U12, P2_R1215_U120, P2_R1215_U121, P2_R1215_U122, P2_R1215_U123, P2_R1215_U124, P2_R1215_U125, P2_R1215_U126, P2_R1215_U127, P2_R1215_U128, P2_R1215_U129, P2_R1215_U13, P2_R1215_U130, P2_R1215_U131, P2_R1215_U132, P2_R1215_U133, P2_R1215_U134, P2_R1215_U135, P2_R1215_U136, P2_R1215_U137, P2_R1215_U138, P2_R1215_U139, P2_R1215_U14, P2_R1215_U140, P2_R1215_U141, P2_R1215_U142, P2_R1215_U143, P2_R1215_U144, P2_R1215_U145, P2_R1215_U146, P2_R1215_U147, P2_R1215_U148, P2_R1215_U149, P2_R1215_U15, P2_R1215_U150, P2_R1215_U151, P2_R1215_U152, P2_R1215_U153, P2_R1215_U154, P2_R1215_U155, P2_R1215_U156, P2_R1215_U157, P2_R1215_U158, P2_R1215_U159, P2_R1215_U16, P2_R1215_U160, P2_R1215_U161, P2_R1215_U162, P2_R1215_U163, P2_R1215_U164, P2_R1215_U165, P2_R1215_U166, P2_R1215_U167, P2_R1215_U168, P2_R1215_U169, P2_R1215_U17, P2_R1215_U170, P2_R1215_U171, P2_R1215_U172, P2_R1215_U173, P2_R1215_U174, P2_R1215_U175, P2_R1215_U176, P2_R1215_U177, P2_R1215_U178, P2_R1215_U179, P2_R1215_U18, P2_R1215_U180, P2_R1215_U181, P2_R1215_U182, P2_R1215_U183, P2_R1215_U184, P2_R1215_U185, P2_R1215_U186, P2_R1215_U187, P2_R1215_U188, P2_R1215_U189, P2_R1215_U19, P2_R1215_U190, P2_R1215_U191, P2_R1215_U192, P2_R1215_U193, P2_R1215_U194, P2_R1215_U195, P2_R1215_U196, P2_R1215_U197, P2_R1215_U198, P2_R1215_U199, P2_R1215_U20, P2_R1215_U200, P2_R1215_U201, P2_R1215_U202, P2_R1215_U203, P2_R1215_U204, P2_R1215_U205, P2_R1215_U206, P2_R1215_U207, P2_R1215_U208, P2_R1215_U209, P2_R1215_U21, P2_R1215_U210, P2_R1215_U211, P2_R1215_U212, P2_R1215_U213, P2_R1215_U214, P2_R1215_U215, P2_R1215_U216, P2_R1215_U217, P2_R1215_U218, P2_R1215_U219, P2_R1215_U22, P2_R1215_U220, P2_R1215_U221, P2_R1215_U222, P2_R1215_U223, P2_R1215_U224, P2_R1215_U225, P2_R1215_U226, P2_R1215_U227, P2_R1215_U228, P2_R1215_U229, P2_R1215_U23, P2_R1215_U230, P2_R1215_U231, P2_R1215_U232, P2_R1215_U233, P2_R1215_U234, P2_R1215_U235, P2_R1215_U236, P2_R1215_U237, P2_R1215_U238, P2_R1215_U239, P2_R1215_U24, P2_R1215_U240, P2_R1215_U241, P2_R1215_U242, P2_R1215_U243, P2_R1215_U244, P2_R1215_U245, P2_R1215_U246, P2_R1215_U247, P2_R1215_U248, P2_R1215_U249, P2_R1215_U25, P2_R1215_U250, P2_R1215_U251, P2_R1215_U252, P2_R1215_U253, P2_R1215_U254, P2_R1215_U255, P2_R1215_U256, P2_R1215_U257, P2_R1215_U258, P2_R1215_U259, P2_R1215_U26, P2_R1215_U260, P2_R1215_U261, P2_R1215_U262, P2_R1215_U263, P2_R1215_U264, P2_R1215_U265, P2_R1215_U266, P2_R1215_U267, P2_R1215_U268, P2_R1215_U269, P2_R1215_U27, P2_R1215_U270, P2_R1215_U271, P2_R1215_U272, P2_R1215_U273, P2_R1215_U274, P2_R1215_U275, P2_R1215_U276, P2_R1215_U277, P2_R1215_U278, P2_R1215_U279, P2_R1215_U28, P2_R1215_U280, P2_R1215_U281, P2_R1215_U282, P2_R1215_U283, P2_R1215_U284, P2_R1215_U285, P2_R1215_U286, P2_R1215_U287, P2_R1215_U288, P2_R1215_U289, P2_R1215_U29, P2_R1215_U290, P2_R1215_U291, P2_R1215_U292, P2_R1215_U293, P2_R1215_U294, P2_R1215_U295, P2_R1215_U296, P2_R1215_U297, P2_R1215_U298, P2_R1215_U299, P2_R1215_U30, P2_R1215_U300, P2_R1215_U301, P2_R1215_U302, P2_R1215_U303, P2_R1215_U304, P2_R1215_U305, P2_R1215_U306, P2_R1215_U307, P2_R1215_U308, P2_R1215_U309, P2_R1215_U31, P2_R1215_U310, P2_R1215_U311, P2_R1215_U312, P2_R1215_U313, P2_R1215_U314, P2_R1215_U315, P2_R1215_U316, P2_R1215_U317, P2_R1215_U318, P2_R1215_U319, P2_R1215_U32, P2_R1215_U320, P2_R1215_U321, P2_R1215_U322, P2_R1215_U323, P2_R1215_U324, P2_R1215_U325, P2_R1215_U326, P2_R1215_U327, P2_R1215_U328, P2_R1215_U329, P2_R1215_U33, P2_R1215_U330, P2_R1215_U331, P2_R1215_U332, P2_R1215_U333, P2_R1215_U334, P2_R1215_U335, P2_R1215_U336, P2_R1215_U337, P2_R1215_U338, P2_R1215_U339, P2_R1215_U34, P2_R1215_U340, P2_R1215_U341, P2_R1215_U342, P2_R1215_U343, P2_R1215_U344, P2_R1215_U345, P2_R1215_U346, P2_R1215_U347, P2_R1215_U348, P2_R1215_U349, P2_R1215_U35, P2_R1215_U350, P2_R1215_U351, P2_R1215_U352, P2_R1215_U353, P2_R1215_U354, P2_R1215_U355, P2_R1215_U356, P2_R1215_U357, P2_R1215_U358, P2_R1215_U359, P2_R1215_U36, P2_R1215_U360, P2_R1215_U361, P2_R1215_U362, P2_R1215_U363, P2_R1215_U364, P2_R1215_U365, P2_R1215_U366, P2_R1215_U367, P2_R1215_U368, P2_R1215_U369, P2_R1215_U37, P2_R1215_U370, P2_R1215_U371, P2_R1215_U372, P2_R1215_U373, P2_R1215_U374, P2_R1215_U375, P2_R1215_U376, P2_R1215_U377, P2_R1215_U378, P2_R1215_U379, P2_R1215_U38, P2_R1215_U380, P2_R1215_U381, P2_R1215_U382, P2_R1215_U383, P2_R1215_U384, P2_R1215_U385, P2_R1215_U386, P2_R1215_U387, P2_R1215_U388, P2_R1215_U389, P2_R1215_U39, P2_R1215_U390, P2_R1215_U391, P2_R1215_U392, P2_R1215_U393, P2_R1215_U394, P2_R1215_U395, P2_R1215_U396, P2_R1215_U397, P2_R1215_U398, P2_R1215_U399, P2_R1215_U4, P2_R1215_U40, P2_R1215_U400, P2_R1215_U401, P2_R1215_U402, P2_R1215_U403, P2_R1215_U404, P2_R1215_U405, P2_R1215_U406, P2_R1215_U407, P2_R1215_U408, P2_R1215_U409, P2_R1215_U41, P2_R1215_U410, P2_R1215_U411, P2_R1215_U412, P2_R1215_U413, P2_R1215_U414, P2_R1215_U415, P2_R1215_U416, P2_R1215_U417, P2_R1215_U418, P2_R1215_U419, P2_R1215_U42, P2_R1215_U420, P2_R1215_U421, P2_R1215_U422, P2_R1215_U423, P2_R1215_U424, P2_R1215_U425, P2_R1215_U426, P2_R1215_U427, P2_R1215_U428, P2_R1215_U429, P2_R1215_U43, P2_R1215_U430, P2_R1215_U431, P2_R1215_U432, P2_R1215_U433, P2_R1215_U434, P2_R1215_U435, P2_R1215_U436, P2_R1215_U437, P2_R1215_U438, P2_R1215_U439, P2_R1215_U44, P2_R1215_U440, P2_R1215_U441, P2_R1215_U442, P2_R1215_U443, P2_R1215_U444, P2_R1215_U445, P2_R1215_U446, P2_R1215_U447, P2_R1215_U448, P2_R1215_U449, P2_R1215_U45, P2_R1215_U450, P2_R1215_U451, P2_R1215_U452, P2_R1215_U453, P2_R1215_U454, P2_R1215_U455, P2_R1215_U456, P2_R1215_U457, P2_R1215_U458, P2_R1215_U459, P2_R1215_U46, P2_R1215_U460, P2_R1215_U461, P2_R1215_U462, P2_R1215_U463, P2_R1215_U464, P2_R1215_U465, P2_R1215_U466, P2_R1215_U467, P2_R1215_U468, P2_R1215_U469, P2_R1215_U47, P2_R1215_U470, P2_R1215_U471, P2_R1215_U472, P2_R1215_U473, P2_R1215_U474, P2_R1215_U475, P2_R1215_U476, P2_R1215_U477, P2_R1215_U478, P2_R1215_U479, P2_R1215_U48, P2_R1215_U480, P2_R1215_U481, P2_R1215_U482, P2_R1215_U483, P2_R1215_U484, P2_R1215_U485, P2_R1215_U486, P2_R1215_U487, P2_R1215_U488, P2_R1215_U489, P2_R1215_U49, P2_R1215_U490, P2_R1215_U491, P2_R1215_U492, P2_R1215_U493, P2_R1215_U494, P2_R1215_U495, P2_R1215_U496, P2_R1215_U497, P2_R1215_U498, P2_R1215_U499, P2_R1215_U5, P2_R1215_U50, P2_R1215_U500, P2_R1215_U501, P2_R1215_U502, P2_R1215_U503, P2_R1215_U504, P2_R1215_U51, P2_R1215_U52, P2_R1215_U53, P2_R1215_U54, P2_R1215_U55, P2_R1215_U56, P2_R1215_U57, P2_R1215_U58, P2_R1215_U59, P2_R1215_U6, P2_R1215_U60, P2_R1215_U61, P2_R1215_U62, P2_R1215_U63, P2_R1215_U64, P2_R1215_U65, P2_R1215_U66, P2_R1215_U67, P2_R1215_U68, P2_R1215_U69, P2_R1215_U7, P2_R1215_U70, P2_R1215_U71, P2_R1215_U72, P2_R1215_U73, P2_R1215_U74, P2_R1215_U75, P2_R1215_U76, P2_R1215_U77, P2_R1215_U78, P2_R1215_U79, P2_R1215_U8, P2_R1215_U80, P2_R1215_U81, P2_R1215_U82, P2_R1215_U83, P2_R1215_U84, P2_R1215_U85, P2_R1215_U86, P2_R1215_U87, P2_R1215_U88, P2_R1215_U89, P2_R1215_U9, P2_R1215_U90, P2_R1215_U91, P2_R1215_U92, P2_R1215_U93, P2_R1215_U94, P2_R1215_U95, P2_R1215_U96, P2_R1215_U97, P2_R1215_U98, P2_R1215_U99, P2_R1233_U10, P2_R1233_U100, P2_R1233_U101, P2_R1233_U102, P2_R1233_U103, P2_R1233_U104, P2_R1233_U105, P2_R1233_U106, P2_R1233_U107, P2_R1233_U108, P2_R1233_U109, P2_R1233_U11, P2_R1233_U110, P2_R1233_U111, P2_R1233_U112, P2_R1233_U113, P2_R1233_U114, P2_R1233_U115, P2_R1233_U116, P2_R1233_U117, P2_R1233_U118, P2_R1233_U119, P2_R1233_U12, P2_R1233_U120, P2_R1233_U121, P2_R1233_U122, P2_R1233_U123, P2_R1233_U124, P2_R1233_U125, P2_R1233_U126, P2_R1233_U127, P2_R1233_U128, P2_R1233_U129, P2_R1233_U13, P2_R1233_U130, P2_R1233_U131, P2_R1233_U132, P2_R1233_U133, P2_R1233_U134, P2_R1233_U135, P2_R1233_U136, P2_R1233_U137, P2_R1233_U138, P2_R1233_U139, P2_R1233_U14, P2_R1233_U140, P2_R1233_U141, P2_R1233_U142, P2_R1233_U143, P2_R1233_U144, P2_R1233_U145, P2_R1233_U146, P2_R1233_U147, P2_R1233_U148, P2_R1233_U149, P2_R1233_U15, P2_R1233_U150, P2_R1233_U151, P2_R1233_U152, P2_R1233_U153, P2_R1233_U154, P2_R1233_U155, P2_R1233_U156, P2_R1233_U157, P2_R1233_U158, P2_R1233_U159, P2_R1233_U16, P2_R1233_U160, P2_R1233_U161, P2_R1233_U162, P2_R1233_U163, P2_R1233_U164, P2_R1233_U165, P2_R1233_U166, P2_R1233_U167, P2_R1233_U168, P2_R1233_U169, P2_R1233_U17, P2_R1233_U170, P2_R1233_U171, P2_R1233_U172, P2_R1233_U173, P2_R1233_U174, P2_R1233_U175, P2_R1233_U176, P2_R1233_U177, P2_R1233_U178, P2_R1233_U179, P2_R1233_U18, P2_R1233_U180, P2_R1233_U181, P2_R1233_U182, P2_R1233_U183, P2_R1233_U184, P2_R1233_U185, P2_R1233_U186, P2_R1233_U187, P2_R1233_U188, P2_R1233_U189, P2_R1233_U19, P2_R1233_U190, P2_R1233_U191, P2_R1233_U192, P2_R1233_U193, P2_R1233_U194, P2_R1233_U195, P2_R1233_U196, P2_R1233_U197, P2_R1233_U198, P2_R1233_U199, P2_R1233_U20, P2_R1233_U200, P2_R1233_U201, P2_R1233_U202, P2_R1233_U203, P2_R1233_U204, P2_R1233_U205, P2_R1233_U206, P2_R1233_U207, P2_R1233_U208, P2_R1233_U209, P2_R1233_U21, P2_R1233_U210, P2_R1233_U211, P2_R1233_U212, P2_R1233_U213, P2_R1233_U214, P2_R1233_U215, P2_R1233_U216, P2_R1233_U217, P2_R1233_U218, P2_R1233_U219, P2_R1233_U22, P2_R1233_U220, P2_R1233_U221, P2_R1233_U222, P2_R1233_U223, P2_R1233_U224, P2_R1233_U225, P2_R1233_U226, P2_R1233_U227, P2_R1233_U228, P2_R1233_U229, P2_R1233_U23, P2_R1233_U230, P2_R1233_U231, P2_R1233_U232, P2_R1233_U233, P2_R1233_U234, P2_R1233_U235, P2_R1233_U236, P2_R1233_U237, P2_R1233_U238, P2_R1233_U239, P2_R1233_U24, P2_R1233_U240, P2_R1233_U241, P2_R1233_U242, P2_R1233_U243, P2_R1233_U244, P2_R1233_U245, P2_R1233_U246, P2_R1233_U247, P2_R1233_U248, P2_R1233_U249, P2_R1233_U25, P2_R1233_U250, P2_R1233_U251, P2_R1233_U252, P2_R1233_U253, P2_R1233_U254, P2_R1233_U255, P2_R1233_U256, P2_R1233_U257, P2_R1233_U258, P2_R1233_U259, P2_R1233_U26, P2_R1233_U260, P2_R1233_U261, P2_R1233_U262, P2_R1233_U263, P2_R1233_U264, P2_R1233_U265, P2_R1233_U266, P2_R1233_U267, P2_R1233_U268, P2_R1233_U269, P2_R1233_U27, P2_R1233_U270, P2_R1233_U271, P2_R1233_U272, P2_R1233_U273, P2_R1233_U274, P2_R1233_U275, P2_R1233_U276, P2_R1233_U277, P2_R1233_U278, P2_R1233_U279, P2_R1233_U28, P2_R1233_U280, P2_R1233_U281, P2_R1233_U282, P2_R1233_U283, P2_R1233_U284, P2_R1233_U285, P2_R1233_U286, P2_R1233_U287, P2_R1233_U288, P2_R1233_U289, P2_R1233_U29, P2_R1233_U290, P2_R1233_U291, P2_R1233_U292, P2_R1233_U293, P2_R1233_U294, P2_R1233_U295, P2_R1233_U296, P2_R1233_U297, P2_R1233_U298, P2_R1233_U299, P2_R1233_U30, P2_R1233_U300, P2_R1233_U301, P2_R1233_U302, P2_R1233_U303, P2_R1233_U304, P2_R1233_U305, P2_R1233_U306, P2_R1233_U307, P2_R1233_U308, P2_R1233_U309, P2_R1233_U31, P2_R1233_U310, P2_R1233_U311, P2_R1233_U312, P2_R1233_U313, P2_R1233_U314, P2_R1233_U315, P2_R1233_U316, P2_R1233_U317, P2_R1233_U318, P2_R1233_U319, P2_R1233_U32, P2_R1233_U320, P2_R1233_U321, P2_R1233_U322, P2_R1233_U323, P2_R1233_U324, P2_R1233_U325, P2_R1233_U326, P2_R1233_U327, P2_R1233_U328, P2_R1233_U329, P2_R1233_U33, P2_R1233_U330, P2_R1233_U331, P2_R1233_U332, P2_R1233_U333, P2_R1233_U334, P2_R1233_U335, P2_R1233_U336, P2_R1233_U337, P2_R1233_U338, P2_R1233_U339, P2_R1233_U34, P2_R1233_U340, P2_R1233_U341, P2_R1233_U342, P2_R1233_U343, P2_R1233_U344, P2_R1233_U345, P2_R1233_U346, P2_R1233_U347, P2_R1233_U348, P2_R1233_U349, P2_R1233_U35, P2_R1233_U350, P2_R1233_U351, P2_R1233_U352, P2_R1233_U353, P2_R1233_U354, P2_R1233_U355, P2_R1233_U356, P2_R1233_U357, P2_R1233_U358, P2_R1233_U359, P2_R1233_U36, P2_R1233_U360, P2_R1233_U361, P2_R1233_U362, P2_R1233_U363, P2_R1233_U364, P2_R1233_U365, P2_R1233_U366, P2_R1233_U367, P2_R1233_U368, P2_R1233_U369, P2_R1233_U37, P2_R1233_U370, P2_R1233_U371, P2_R1233_U372, P2_R1233_U373, P2_R1233_U374, P2_R1233_U375, P2_R1233_U376, P2_R1233_U377, P2_R1233_U378, P2_R1233_U379, P2_R1233_U38, P2_R1233_U380, P2_R1233_U381, P2_R1233_U382, P2_R1233_U383, P2_R1233_U384, P2_R1233_U385, P2_R1233_U386, P2_R1233_U387, P2_R1233_U388, P2_R1233_U389, P2_R1233_U39, P2_R1233_U390, P2_R1233_U391, P2_R1233_U392, P2_R1233_U393, P2_R1233_U394, P2_R1233_U395, P2_R1233_U396, P2_R1233_U397, P2_R1233_U398, P2_R1233_U399, P2_R1233_U4, P2_R1233_U40, P2_R1233_U400, P2_R1233_U401, P2_R1233_U402, P2_R1233_U403, P2_R1233_U404, P2_R1233_U405, P2_R1233_U406, P2_R1233_U407, P2_R1233_U408, P2_R1233_U409, P2_R1233_U41, P2_R1233_U410, P2_R1233_U411, P2_R1233_U412, P2_R1233_U413, P2_R1233_U414, P2_R1233_U415, P2_R1233_U416, P2_R1233_U417, P2_R1233_U418, P2_R1233_U419, P2_R1233_U42, P2_R1233_U420, P2_R1233_U421, P2_R1233_U422, P2_R1233_U423, P2_R1233_U424, P2_R1233_U425, P2_R1233_U426, P2_R1233_U427, P2_R1233_U428, P2_R1233_U429, P2_R1233_U43, P2_R1233_U430, P2_R1233_U431, P2_R1233_U432, P2_R1233_U433, P2_R1233_U434, P2_R1233_U435, P2_R1233_U436, P2_R1233_U437, P2_R1233_U438, P2_R1233_U439, P2_R1233_U44, P2_R1233_U440, P2_R1233_U441, P2_R1233_U442, P2_R1233_U443, P2_R1233_U444, P2_R1233_U445, P2_R1233_U446, P2_R1233_U447, P2_R1233_U448, P2_R1233_U449, P2_R1233_U45, P2_R1233_U450, P2_R1233_U451, P2_R1233_U452, P2_R1233_U453, P2_R1233_U454, P2_R1233_U455, P2_R1233_U456, P2_R1233_U457, P2_R1233_U458, P2_R1233_U459, P2_R1233_U46, P2_R1233_U460, P2_R1233_U461, P2_R1233_U462, P2_R1233_U463, P2_R1233_U464, P2_R1233_U465, P2_R1233_U466, P2_R1233_U467, P2_R1233_U468, P2_R1233_U469, P2_R1233_U47, P2_R1233_U470, P2_R1233_U471, P2_R1233_U472, P2_R1233_U473, P2_R1233_U474, P2_R1233_U475, P2_R1233_U476, P2_R1233_U477, P2_R1233_U478, P2_R1233_U479, P2_R1233_U48, P2_R1233_U480, P2_R1233_U481, P2_R1233_U482, P2_R1233_U483, P2_R1233_U484, P2_R1233_U485, P2_R1233_U486, P2_R1233_U487, P2_R1233_U488, P2_R1233_U489, P2_R1233_U49, P2_R1233_U490, P2_R1233_U491, P2_R1233_U492, P2_R1233_U493, P2_R1233_U494, P2_R1233_U495, P2_R1233_U496, P2_R1233_U497, P2_R1233_U498, P2_R1233_U499, P2_R1233_U5, P2_R1233_U50, P2_R1233_U500, P2_R1233_U501, P2_R1233_U502, P2_R1233_U503, P2_R1233_U504, P2_R1233_U51, P2_R1233_U52, P2_R1233_U53, P2_R1233_U54, P2_R1233_U55, P2_R1233_U56, P2_R1233_U57, P2_R1233_U58, P2_R1233_U59, P2_R1233_U6, P2_R1233_U60, P2_R1233_U61, P2_R1233_U62, P2_R1233_U63, P2_R1233_U64, P2_R1233_U65, P2_R1233_U66, P2_R1233_U67, P2_R1233_U68, P2_R1233_U69, P2_R1233_U7, P2_R1233_U70, P2_R1233_U71, P2_R1233_U72, P2_R1233_U73, P2_R1233_U74, P2_R1233_U75, P2_R1233_U76, P2_R1233_U77, P2_R1233_U78, P2_R1233_U79, P2_R1233_U8, P2_R1233_U80, P2_R1233_U81, P2_R1233_U82, P2_R1233_U83, P2_R1233_U84, P2_R1233_U85, P2_R1233_U86, P2_R1233_U87, P2_R1233_U88, P2_R1233_U89, P2_R1233_U9, P2_R1233_U90, P2_R1233_U91, P2_R1233_U92, P2_R1233_U93, P2_R1233_U94, P2_R1233_U95, P2_R1233_U96, P2_R1233_U97, P2_R1233_U98, P2_R1233_U99, P2_R1275_U10, P2_R1275_U100, P2_R1275_U101, P2_R1275_U102, P2_R1275_U103, P2_R1275_U104, P2_R1275_U105, P2_R1275_U106, P2_R1275_U107, P2_R1275_U108, P2_R1275_U109, P2_R1275_U11, P2_R1275_U110, P2_R1275_U111, P2_R1275_U112, P2_R1275_U113, P2_R1275_U114, P2_R1275_U115, P2_R1275_U116, P2_R1275_U117, P2_R1275_U118, P2_R1275_U119, P2_R1275_U12, P2_R1275_U120, P2_R1275_U121, P2_R1275_U122, P2_R1275_U123, P2_R1275_U124, P2_R1275_U125, P2_R1275_U126, P2_R1275_U127, P2_R1275_U128, P2_R1275_U129, P2_R1275_U13, P2_R1275_U130, P2_R1275_U131, P2_R1275_U132, P2_R1275_U133, P2_R1275_U134, P2_R1275_U135, P2_R1275_U136, P2_R1275_U137, P2_R1275_U138, P2_R1275_U139, P2_R1275_U14, P2_R1275_U140, P2_R1275_U141, P2_R1275_U142, P2_R1275_U143, P2_R1275_U144, P2_R1275_U145, P2_R1275_U146, P2_R1275_U147, P2_R1275_U148, P2_R1275_U149, P2_R1275_U15, P2_R1275_U150, P2_R1275_U151, P2_R1275_U152, P2_R1275_U153, P2_R1275_U154, P2_R1275_U155, P2_R1275_U156, P2_R1275_U157, P2_R1275_U158, P2_R1275_U159, P2_R1275_U16, P2_R1275_U17, P2_R1275_U18, P2_R1275_U19, P2_R1275_U20, P2_R1275_U21, P2_R1275_U22, P2_R1275_U23, P2_R1275_U24, P2_R1275_U25, P2_R1275_U26, P2_R1275_U27, P2_R1275_U28, P2_R1275_U29, P2_R1275_U30, P2_R1275_U31, P2_R1275_U32, P2_R1275_U33, P2_R1275_U34, P2_R1275_U35, P2_R1275_U36, P2_R1275_U37, P2_R1275_U38, P2_R1275_U39, P2_R1275_U40, P2_R1275_U41, P2_R1275_U42, P2_R1275_U43, P2_R1275_U44, P2_R1275_U45, P2_R1275_U46, P2_R1275_U47, P2_R1275_U48, P2_R1275_U49, P2_R1275_U50, P2_R1275_U51, P2_R1275_U52, P2_R1275_U53, P2_R1275_U54, P2_R1275_U55, P2_R1275_U56, P2_R1275_U57, P2_R1275_U58, P2_R1275_U59, P2_R1275_U6, P2_R1275_U60, P2_R1275_U61, P2_R1275_U62, P2_R1275_U63, P2_R1275_U64, P2_R1275_U65, P2_R1275_U66, P2_R1275_U67, P2_R1275_U68, P2_R1275_U69, P2_R1275_U7, P2_R1275_U70, P2_R1275_U71, P2_R1275_U72, P2_R1275_U73, P2_R1275_U74, P2_R1275_U75, P2_R1275_U76, P2_R1275_U77, P2_R1275_U78, P2_R1275_U79, P2_R1275_U8, P2_R1275_U80, P2_R1275_U81, P2_R1275_U82, P2_R1275_U83, P2_R1275_U84, P2_R1275_U85, P2_R1275_U86, P2_R1275_U87, P2_R1275_U88, P2_R1275_U89, P2_R1275_U9, P2_R1275_U90, P2_R1275_U91, P2_R1275_U92, P2_R1275_U93, P2_R1275_U94, P2_R1275_U95, P2_R1275_U96, P2_R1275_U97, P2_R1275_U98, P2_R1275_U99, P2_R1299_U6, P2_R1299_U7, P2_R1312_U10, P2_R1312_U100, P2_R1312_U101, P2_R1312_U102, P2_R1312_U103, P2_R1312_U104, P2_R1312_U105, P2_R1312_U106, P2_R1312_U107, P2_R1312_U108, P2_R1312_U109, P2_R1312_U11, P2_R1312_U110, P2_R1312_U111, P2_R1312_U112, P2_R1312_U113, P2_R1312_U114, P2_R1312_U115, P2_R1312_U116, P2_R1312_U117, P2_R1312_U118, P2_R1312_U119, P2_R1312_U12, P2_R1312_U120, P2_R1312_U121, P2_R1312_U122, P2_R1312_U123, P2_R1312_U124, P2_R1312_U125, P2_R1312_U126, P2_R1312_U127, P2_R1312_U128, P2_R1312_U129, P2_R1312_U13, P2_R1312_U130, P2_R1312_U131, P2_R1312_U132, P2_R1312_U133, P2_R1312_U134, P2_R1312_U135, P2_R1312_U136, P2_R1312_U137, P2_R1312_U138, P2_R1312_U139, P2_R1312_U14, P2_R1312_U140, P2_R1312_U141, P2_R1312_U142, P2_R1312_U143, P2_R1312_U144, P2_R1312_U145, P2_R1312_U146, P2_R1312_U147, P2_R1312_U148, P2_R1312_U149, P2_R1312_U15, P2_R1312_U150, P2_R1312_U151, P2_R1312_U152, P2_R1312_U153, P2_R1312_U154, P2_R1312_U155, P2_R1312_U156, P2_R1312_U157, P2_R1312_U158, P2_R1312_U159, P2_R1312_U16, P2_R1312_U160, P2_R1312_U161, P2_R1312_U162, P2_R1312_U163, P2_R1312_U164, P2_R1312_U165, P2_R1312_U166, P2_R1312_U167, P2_R1312_U168, P2_R1312_U169, P2_R1312_U17, P2_R1312_U170, P2_R1312_U171, P2_R1312_U172, P2_R1312_U173, P2_R1312_U174, P2_R1312_U175, P2_R1312_U176, P2_R1312_U177, P2_R1312_U178, P2_R1312_U179, P2_R1312_U18, P2_R1312_U180, P2_R1312_U181, P2_R1312_U182, P2_R1312_U183, P2_R1312_U184, P2_R1312_U185, P2_R1312_U186, P2_R1312_U187, P2_R1312_U188, P2_R1312_U189, P2_R1312_U19, P2_R1312_U190, P2_R1312_U191, P2_R1312_U192, P2_R1312_U193, P2_R1312_U194, P2_R1312_U195, P2_R1312_U196, P2_R1312_U197, P2_R1312_U198, P2_R1312_U199, P2_R1312_U20, P2_R1312_U200, P2_R1312_U201, P2_R1312_U202, P2_R1312_U203, P2_R1312_U204, P2_R1312_U205, P2_R1312_U206, P2_R1312_U207, P2_R1312_U208, P2_R1312_U209, P2_R1312_U21, P2_R1312_U210, P2_R1312_U211, P2_R1312_U212, P2_R1312_U213, P2_R1312_U214, P2_R1312_U215, P2_R1312_U216, P2_R1312_U217, P2_R1312_U218, P2_R1312_U219, P2_R1312_U22, P2_R1312_U220, P2_R1312_U221, P2_R1312_U222, P2_R1312_U223, P2_R1312_U224, P2_R1312_U225, P2_R1312_U226, P2_R1312_U227, P2_R1312_U23, P2_R1312_U24, P2_R1312_U25, P2_R1312_U26, P2_R1312_U27, P2_R1312_U28, P2_R1312_U29, P2_R1312_U30, P2_R1312_U31, P2_R1312_U32, P2_R1312_U33, P2_R1312_U34, P2_R1312_U35, P2_R1312_U36, P2_R1312_U37, P2_R1312_U38, P2_R1312_U39, P2_R1312_U40, P2_R1312_U41, P2_R1312_U42, P2_R1312_U43, P2_R1312_U44, P2_R1312_U45, P2_R1312_U46, P2_R1312_U47, P2_R1312_U48, P2_R1312_U49, P2_R1312_U50, P2_R1312_U51, P2_R1312_U52, P2_R1312_U53, P2_R1312_U54, P2_R1312_U55, P2_R1312_U56, P2_R1312_U57, P2_R1312_U58, P2_R1312_U59, P2_R1312_U6, P2_R1312_U60, P2_R1312_U61, P2_R1312_U62, P2_R1312_U63, P2_R1312_U64, P2_R1312_U65, P2_R1312_U66, P2_R1312_U67, P2_R1312_U68, P2_R1312_U69, P2_R1312_U7, P2_R1312_U70, P2_R1312_U71, P2_R1312_U72, P2_R1312_U73, P2_R1312_U74, P2_R1312_U75, P2_R1312_U76, P2_R1312_U77, P2_R1312_U78, P2_R1312_U79, P2_R1312_U8, P2_R1312_U80, P2_R1312_U81, P2_R1312_U82, P2_R1312_U83, P2_R1312_U84, P2_R1312_U85, P2_R1312_U86, P2_R1312_U87, P2_R1312_U88, P2_R1312_U89, P2_R1312_U9, P2_R1312_U90, P2_R1312_U91, P2_R1312_U92, P2_R1312_U93, P2_R1312_U94, P2_R1312_U95, P2_R1312_U96, P2_R1312_U97, P2_R1312_U98, P2_R1312_U99, P2_R1335_U10, P2_R1335_U6, P2_R1335_U7, P2_R1335_U8, P2_R1335_U9, P2_SUB_1108_U10, P2_SUB_1108_U100, P2_SUB_1108_U101, P2_SUB_1108_U102, P2_SUB_1108_U103, P2_SUB_1108_U104, P2_SUB_1108_U105, P2_SUB_1108_U106, P2_SUB_1108_U107, P2_SUB_1108_U108, P2_SUB_1108_U109, P2_SUB_1108_U11, P2_SUB_1108_U110, P2_SUB_1108_U111, P2_SUB_1108_U112, P2_SUB_1108_U113, P2_SUB_1108_U114, P2_SUB_1108_U115, P2_SUB_1108_U116, P2_SUB_1108_U117, P2_SUB_1108_U118, P2_SUB_1108_U119, P2_SUB_1108_U12, P2_SUB_1108_U120, P2_SUB_1108_U121, P2_SUB_1108_U122, P2_SUB_1108_U123, P2_SUB_1108_U124, P2_SUB_1108_U125, P2_SUB_1108_U126, P2_SUB_1108_U127, P2_SUB_1108_U128, P2_SUB_1108_U129, P2_SUB_1108_U13, P2_SUB_1108_U130, P2_SUB_1108_U131, P2_SUB_1108_U132, P2_SUB_1108_U133, P2_SUB_1108_U134, P2_SUB_1108_U135, P2_SUB_1108_U136, P2_SUB_1108_U137, P2_SUB_1108_U138, P2_SUB_1108_U139, P2_SUB_1108_U14, P2_SUB_1108_U140, P2_SUB_1108_U141, P2_SUB_1108_U142, P2_SUB_1108_U143, P2_SUB_1108_U144, P2_SUB_1108_U145, P2_SUB_1108_U146, P2_SUB_1108_U147, P2_SUB_1108_U148, P2_SUB_1108_U149, P2_SUB_1108_U15, P2_SUB_1108_U150, P2_SUB_1108_U151, P2_SUB_1108_U152, P2_SUB_1108_U153, P2_SUB_1108_U154, P2_SUB_1108_U155, P2_SUB_1108_U156, P2_SUB_1108_U157, P2_SUB_1108_U158, P2_SUB_1108_U159, P2_SUB_1108_U16, P2_SUB_1108_U160, P2_SUB_1108_U161, P2_SUB_1108_U162, P2_SUB_1108_U163, P2_SUB_1108_U164, P2_SUB_1108_U165, P2_SUB_1108_U166, P2_SUB_1108_U167, P2_SUB_1108_U168, P2_SUB_1108_U169, P2_SUB_1108_U17, P2_SUB_1108_U170, P2_SUB_1108_U171, P2_SUB_1108_U172, P2_SUB_1108_U173, P2_SUB_1108_U174, P2_SUB_1108_U175, P2_SUB_1108_U176, P2_SUB_1108_U177, P2_SUB_1108_U178, P2_SUB_1108_U179, P2_SUB_1108_U18, P2_SUB_1108_U180, P2_SUB_1108_U181, P2_SUB_1108_U182, P2_SUB_1108_U183, P2_SUB_1108_U184, P2_SUB_1108_U185, P2_SUB_1108_U186, P2_SUB_1108_U187, P2_SUB_1108_U188, P2_SUB_1108_U189, P2_SUB_1108_U19, P2_SUB_1108_U190, P2_SUB_1108_U191, P2_SUB_1108_U192, P2_SUB_1108_U193, P2_SUB_1108_U194, P2_SUB_1108_U195, P2_SUB_1108_U196, P2_SUB_1108_U197, P2_SUB_1108_U198, P2_SUB_1108_U199, P2_SUB_1108_U20, P2_SUB_1108_U200, P2_SUB_1108_U201, P2_SUB_1108_U202, P2_SUB_1108_U21, P2_SUB_1108_U22, P2_SUB_1108_U23, P2_SUB_1108_U24, P2_SUB_1108_U25, P2_SUB_1108_U26, P2_SUB_1108_U27, P2_SUB_1108_U28, P2_SUB_1108_U29, P2_SUB_1108_U30, P2_SUB_1108_U31, P2_SUB_1108_U32, P2_SUB_1108_U33, P2_SUB_1108_U34, P2_SUB_1108_U35, P2_SUB_1108_U36, P2_SUB_1108_U37, P2_SUB_1108_U38, P2_SUB_1108_U39, P2_SUB_1108_U40, P2_SUB_1108_U41, P2_SUB_1108_U42, P2_SUB_1108_U43, P2_SUB_1108_U44, P2_SUB_1108_U45, P2_SUB_1108_U46, P2_SUB_1108_U47, P2_SUB_1108_U48, P2_SUB_1108_U49, P2_SUB_1108_U50, P2_SUB_1108_U51, P2_SUB_1108_U52, P2_SUB_1108_U53, P2_SUB_1108_U54, P2_SUB_1108_U55, P2_SUB_1108_U56, P2_SUB_1108_U57, P2_SUB_1108_U58, P2_SUB_1108_U59, P2_SUB_1108_U6, P2_SUB_1108_U60, P2_SUB_1108_U61, P2_SUB_1108_U62, P2_SUB_1108_U63, P2_SUB_1108_U64, P2_SUB_1108_U65, P2_SUB_1108_U66, P2_SUB_1108_U67, P2_SUB_1108_U68, P2_SUB_1108_U69, P2_SUB_1108_U7, P2_SUB_1108_U70, P2_SUB_1108_U71, P2_SUB_1108_U72, P2_SUB_1108_U73, P2_SUB_1108_U74, P2_SUB_1108_U75, P2_SUB_1108_U76, P2_SUB_1108_U77, P2_SUB_1108_U78, P2_SUB_1108_U79, P2_SUB_1108_U8, P2_SUB_1108_U80, P2_SUB_1108_U81, P2_SUB_1108_U82, P2_SUB_1108_U83, P2_SUB_1108_U84, P2_SUB_1108_U85, P2_SUB_1108_U86, P2_SUB_1108_U87, P2_SUB_1108_U88, P2_SUB_1108_U89, P2_SUB_1108_U9, P2_SUB_1108_U90, P2_SUB_1108_U91, P2_SUB_1108_U92, P2_SUB_1108_U93, P2_SUB_1108_U94, P2_SUB_1108_U95, P2_SUB_1108_U96, P2_SUB_1108_U97, P2_SUB_1108_U98, P2_SUB_1108_U99, P2_U3014, P2_U3015, P2_U3016, P2_U3017, P2_U3018, P2_U3019, P2_U3020, P2_U3021, P2_U3022, P2_U3023, P2_U3024, P2_U3025, P2_U3026, P2_U3027, P2_U3028, P2_U3029, P2_U3030, P2_U3031, P2_U3032, P2_U3033, P2_U3034, P2_U3035, P2_U3036, P2_U3037, P2_U3038, P2_U3039, P2_U3040, P2_U3041, P2_U3042, P2_U3043, P2_U3044, P2_U3045, P2_U3046, P2_U3047, P2_U3048, P2_U3049, P2_U3050, P2_U3051, P2_U3052, P2_U3053, P2_U3054, P2_U3055, P2_U3056, P2_U3057, P2_U3058, P2_U3059, P2_U3060, P2_U3061, P2_U3062, P2_U3063, P2_U3064, P2_U3065, P2_U3066, P2_U3067, P2_U3068, P2_U3069, P2_U3070, P2_U3071, P2_U3072, P2_U3073, P2_U3074, P2_U3075, P2_U3076, P2_U3077, P2_U3078, P2_U3079, P2_U3080, P2_U3081, P2_U3082, P2_U3083, P2_U3084, P2_U3085, P2_U3086, P2_U3089, P2_U3090, P2_U3091, P2_U3092, P2_U3093, P2_U3094, P2_U3095, P2_U3096, P2_U3097, P2_U3098, P2_U3099, P2_U3100, P2_U3101, P2_U3102, P2_U3103, P2_U3104, P2_U3105, P2_U3106, P2_U3107, P2_U3108, P2_U3109, P2_U3110, P2_U3111, P2_U3112, P2_U3113, P2_U3114, P2_U3115, P2_U3116, P2_U3117, P2_U3118, P2_U3119, P2_U3120, P2_U3121, P2_U3122, P2_U3123, P2_U3124, P2_U3125, P2_U3126, P2_U3127, P2_U3128, P2_U3129, P2_U3130, P2_U3131, P2_U3132, P2_U3133, P2_U3134, P2_U3135, P2_U3136, P2_U3137, P2_U3138, P2_U3139, P2_U3140, P2_U3141, P2_U3142, P2_U3143, P2_U3144, P2_U3145, P2_U3146, P2_U3147, P2_U3148, P2_U3149, P2_U3150, P2_U3151, P2_U3152, P2_U3153, P2_U3154, P2_U3155, P2_U3156, P2_U3157, P2_U3158, P2_U3159, P2_U3160, P2_U3161, P2_U3162, P2_U3163, P2_U3164, P2_U3165, P2_U3166, P2_U3167, P2_U3168, P2_U3169, P2_U3170, P2_U3171, P2_U3172, P2_U3173, P2_U3174, P2_U3175, P2_U3176, P2_U3177, P2_U3178, P2_U3179, P2_U3180, P2_U3181, P2_U3182, P2_U3183, P2_U3184, P2_U3329, P2_U3330, P2_U3331, P2_U3332, P2_U3333, P2_U3334, P2_U3335, P2_U3336, P2_U3337, P2_U3338, P2_U3339, P2_U3340, P2_U3341, P2_U3342, P2_U3343, P2_U3344, P2_U3345, P2_U3346, P2_U3347, P2_U3348, P2_U3349, P2_U3350, P2_U3351, P2_U3352, P2_U3353, P2_U3354, P2_U3355, P2_U3356, P2_U3357, P2_U3358, P2_U3359, P2_U3360, P2_U3361, P2_U3362, P2_U3363, P2_U3364, P2_U3365, P2_U3366, P2_U3367, P2_U3368, P2_U3369, P2_U3370, P2_U3371, P2_U3372, P2_U3373, P2_U3374, P2_U3375, P2_U3376, P2_U3377, P2_U3378, P2_U3379, P2_U3380, P2_U3381, P2_U3382, P2_U3383, P2_U3384, P2_U3385, P2_U3386, P2_U3387, P2_U3388, P2_U3389, P2_U3390, P2_U3391, P2_U3392, P2_U3393, P2_U3394, P2_U3395, P2_U3396, P2_U3397, P2_U3398, P2_U3399, P2_U3400, P2_U3401, P2_U3402, P2_U3403, P2_U3404, P2_U3405, P2_U3406, P2_U3407, P2_U3408, P2_U3409, P2_U3410, P2_U3411, P2_U3412, P2_U3413, P2_U3414, P2_U3415, P2_U3418, P2_U3419, P2_U3420, P2_U3421, P2_U3422, P2_U3423, P2_U3424, P2_U3425, P2_U3426, P2_U3427, P2_U3428, P2_U3429, P2_U3431, P2_U3432, P2_U3434, P2_U3435, P2_U3437, P2_U3438, P2_U3440, P2_U3441, P2_U3443, P2_U3444, P2_U3446, P2_U3447, P2_U3449, P2_U3450, P2_U3452, P2_U3453, P2_U3455, P2_U3456, P2_U3458, P2_U3459, P2_U3461, P2_U3462, P2_U3464, P2_U3465, P2_U3467, P2_U3468, P2_U3470, P2_U3471, P2_U3473, P2_U3474, P2_U3476, P2_U3477, P2_U3479, P2_U3480, P2_U3482, P2_U3483, P2_U3485, P2_U3563, P2_U3564, P2_U3565, P2_U3566, P2_U3567, P2_U3568, P2_U3569, P2_U3570, P2_U3571, P2_U3572, P2_U3573, P2_U3574, P2_U3575, P2_U3576, P2_U3577, P2_U3578, P2_U3579, P2_U3580, P2_U3581, P2_U3582, P2_U3583, P2_U3584, P2_U3585, P2_U3586, P2_U3587, P2_U3588, P2_U3589, P2_U3590, P2_U3591, P2_U3592, P2_U3593, P2_U3594, P2_U3595, P2_U3596, P2_U3597, P2_U3598, P2_U3599, P2_U3600, P2_U3601, P2_U3602, P2_U3603, P2_U3604, P2_U3605, P2_U3606, P2_U3607, P2_U3608, P2_U3609, P2_U3610, P2_U3611, P2_U3612, P2_U3613, P2_U3614, P2_U3615, P2_U3616, P2_U3617, P2_U3618, P2_U3619, P2_U3620, P2_U3621, P2_U3622, P2_U3623, P2_U3624, P2_U3625, P2_U3626, P2_U3627, P2_U3628, P2_U3629, P2_U3630, P2_U3631, P2_U3632, P2_U3633, P2_U3634, P2_U3635, P2_U3636, P2_U3637, P2_U3638, P2_U3639, P2_U3640, P2_U3641, P2_U3642, P2_U3643, P2_U3644, P2_U3645, P2_U3646, P2_U3647, P2_U3648, P2_U3649, P2_U3650, P2_U3651, P2_U3652, P2_U3653, P2_U3654, P2_U3655, P2_U3656, P2_U3657, P2_U3658, P2_U3659, P2_U3660, P2_U3661, P2_U3662, P2_U3663, P2_U3664, P2_U3665, P2_U3666, P2_U3667, P2_U3668, P2_U3669, P2_U3670, P2_U3671, P2_U3672, P2_U3673, P2_U3674, P2_U3675, P2_U3676, P2_U3677, P2_U3678, P2_U3679, P2_U3680, P2_U3681, P2_U3682, P2_U3683, P2_U3684, P2_U3685, P2_U3686, P2_U3687, P2_U3688, P2_U3689, P2_U3690, P2_U3691, P2_U3692, P2_U3693, P2_U3694, P2_U3695, P2_U3696, P2_U3697, P2_U3698, P2_U3699, P2_U3700, P2_U3701, P2_U3702, P2_U3703, P2_U3704, P2_U3705, P2_U3706, P2_U3707, P2_U3708, P2_U3709, P2_U3710, P2_U3711, P2_U3712, P2_U3713, P2_U3714, P2_U3715, P2_U3716, P2_U3717, P2_U3718, P2_U3719, P2_U3720, P2_U3721, P2_U3722, P2_U3723, P2_U3724, P2_U3725, P2_U3726, P2_U3727, P2_U3728, P2_U3729, P2_U3730, P2_U3731, P2_U3732, P2_U3733, P2_U3734, P2_U3735, P2_U3736, P2_U3737, P2_U3738, P2_U3739, P2_U3740, P2_U3741, P2_U3742, P2_U3743, P2_U3744, P2_U3745, P2_U3746, P2_U3747, P2_U3748, P2_U3749, P2_U3750, P2_U3751, P2_U3752, P2_U3753, P2_U3754, P2_U3755, P2_U3756, P2_U3757, P2_U3758, P2_U3759, P2_U3760, P2_U3761, P2_U3762, P2_U3763, P2_U3764, P2_U3765, P2_U3766, P2_U3767, P2_U3768, P2_U3769, P2_U3770, P2_U3771, P2_U3772, P2_U3773, P2_U3774, P2_U3775, P2_U3776, P2_U3777, P2_U3778, P2_U3779, P2_U3780, P2_U3781, P2_U3782, P2_U3783, P2_U3784, P2_U3785, P2_U3786, P2_U3787, P2_U3788, P2_U3789, P2_U3790, P2_U3791, P2_U3792, P2_U3793, P2_U3794, P2_U3795, P2_U3796, P2_U3797, P2_U3798, P2_U3799, P2_U3800, P2_U3801, P2_U3802, P2_U3803, P2_U3804, P2_U3805, P2_U3806, P2_U3807, P2_U3808, P2_U3809, P2_U3810, P2_U3811, P2_U3812, P2_U3813, P2_U3814, P2_U3815, P2_U3816, P2_U3817, P2_U3818, P2_U3819, P2_U3820, P2_U3821, P2_U3822, P2_U3823, P2_U3824, P2_U3825, P2_U3826, P2_U3827, P2_U3828, P2_U3829, P2_U3830, P2_U3831, P2_U3832, P2_U3833, P2_U3834, P2_U3835, P2_U3836, P2_U3837, P2_U3838, P2_U3839, P2_U3840, P2_U3841, P2_U3842, P2_U3843, P2_U3844, P2_U3845, P2_U3846, P2_U3847, P2_U3848, P2_U3849, P2_U3850, P2_U3851, P2_U3852, P2_U3853, P2_U3854, P2_U3855, P2_U3856, P2_U3857, P2_U3858, P2_U3859, P2_U3860, P2_U3861, P2_U3862, P2_U3863, P2_U3864, P2_U3865, P2_U3866, P2_U3867, P2_U3868, P2_U3869, P2_U3870, P2_U3871, P2_U3872, P2_U3873, P2_U3874, P2_U3875, P2_U3876, P2_U3877, P2_U3878, P2_U3879, P2_U3880, P2_U3881, P2_U3882, P2_U3883, P2_U3884, P2_U3885, P2_U3886, P2_U3887, P2_U3888, P2_U3889, P2_U3890, P2_U3891, P2_U3892, P2_U3893, P2_U3894, P2_U3895, P2_U3896, P2_U3897, P2_U3898, P2_U3899, P2_U3900, P2_U3901, P2_U3902, P2_U3903, P2_U3904, P2_U3905, P2_U3906, P2_U3907, P2_U3908, P2_U3909, P2_U3910, P2_U3911, P2_U3912, P2_U3913, P2_U3914, P2_U3915, P2_U3916, P2_U3917, P2_U3918, P2_U3919, P2_U3920, P2_U3921, P2_U3922, P2_U3923, P2_U3924, P2_U3925, P2_U3926, P2_U3927, P2_U3928, P2_U3929, P2_U3930, P2_U3931, P2_U3932, P2_U3933, P2_U3934, P2_U3935, P2_U3936, P2_U3937, P2_U3938, P2_U3939, P2_U3940, P2_U3941, P2_U3942, P2_U3943, P2_U3944, P2_U3945, P2_U3946, P2_U3948, P2_U3949, P2_U3950, P2_U3951, P2_U3952, P2_U3953, P2_U3954, P2_U3955, P2_U3956, P2_U3957, P2_U3958, P2_U3959, P2_U3960, P2_U3961, P2_U3962, P2_U3963, P2_U3964, P2_U3965, P2_U3966, P2_U3967, P2_U3968, P2_U3969, P2_U3970, P2_U3971, P2_U3972, P2_U3973, P2_U3974, P2_U3975, P2_U3976, P2_U3977, P2_U3978, P2_U3979, P2_U3980, P2_U3981, P2_U3982, P2_U3983, P2_U3984, P2_U3985, P2_U3986, P2_U3987, P2_U3988, P2_U3989, P2_U3990, P2_U3991, P2_U3992, P2_U3993, P2_U3994, P2_U3995, P2_U3996, P2_U3997, P2_U3998, P2_U3999, P2_U4000, P2_U4001, P2_U4002, P2_U4003, P2_U4004, P2_U4005, P2_U4006, P2_U4007, P2_U4008, P2_U4009, P2_U4010, P2_U4011, P2_U4012, P2_U4013, P2_U4014, P2_U4015, P2_U4016, P2_U4017, P2_U4018, P2_U4019, P2_U4020, P2_U4021, P2_U4022, P2_U4023, P2_U4024, P2_U4025, P2_U4026, P2_U4027, P2_U4028, P2_U4029, P2_U4030, P2_U4031, P2_U4032, P2_U4033, P2_U4034, P2_U4035, P2_U4036, P2_U4037, P2_U4038, P2_U4039, P2_U4040, P2_U4041, P2_U4042, P2_U4043, P2_U4044, P2_U4045, P2_U4046, P2_U4047, P2_U4048, P2_U4049, P2_U4050, P2_U4051, P2_U4052, P2_U4053, P2_U4054, P2_U4055, P2_U4056, P2_U4057, P2_U4058, P2_U4059, P2_U4060, P2_U4061, P2_U4062, P2_U4063, P2_U4064, P2_U4065, P2_U4066, P2_U4067, P2_U4068, P2_U4069, P2_U4070, P2_U4071, P2_U4072, P2_U4073, P2_U4074, P2_U4075, P2_U4076, P2_U4077, P2_U4078, P2_U4079, P2_U4080, P2_U4081, P2_U4082, P2_U4083, P2_U4084, P2_U4085, P2_U4086, P2_U4087, P2_U4088, P2_U4089, P2_U4090, P2_U4091, P2_U4092, P2_U4093, P2_U4094, P2_U4095, P2_U4096, P2_U4097, P2_U4098, P2_U4099, P2_U4100, P2_U4101, P2_U4102, P2_U4103, P2_U4104, P2_U4105, P2_U4106, P2_U4107, P2_U4108, P2_U4109, P2_U4110, P2_U4111, P2_U4112, P2_U4113, P2_U4114, P2_U4115, P2_U4116, P2_U4117, P2_U4118, P2_U4119, P2_U4120, P2_U4121, P2_U4122, P2_U4123, P2_U4124, P2_U4125, P2_U4126, P2_U4127, P2_U4128, P2_U4129, P2_U4130, P2_U4131, P2_U4132, P2_U4133, P2_U4134, P2_U4135, P2_U4136, P2_U4137, P2_U4138, P2_U4139, P2_U4140, P2_U4141, P2_U4142, P2_U4143, P2_U4144, P2_U4145, P2_U4146, P2_U4147, P2_U4148, P2_U4149, P2_U4150, P2_U4151, P2_U4152, P2_U4153, P2_U4154, P2_U4155, P2_U4156, P2_U4157, P2_U4158, P2_U4159, P2_U4160, P2_U4161, P2_U4162, P2_U4163, P2_U4164, P2_U4165, P2_U4166, P2_U4167, P2_U4168, P2_U4169, P2_U4170, P2_U4171, P2_U4172, P2_U4173, P2_U4174, P2_U4175, P2_U4176, P2_U4177, P2_U4178, P2_U4179, P2_U4180, P2_U4181, P2_U4182, P2_U4183, P2_U4184, P2_U4185, P2_U4186, P2_U4187, P2_U4188, P2_U4189, P2_U4190, P2_U4191, P2_U4192, P2_U4193, P2_U4194, P2_U4195, P2_U4196, P2_U4197, P2_U4198, P2_U4199, P2_U4200, P2_U4201, P2_U4202, P2_U4203, P2_U4204, P2_U4205, P2_U4206, P2_U4207, P2_U4208, P2_U4209, P2_U4210, P2_U4211, P2_U4212, P2_U4213, P2_U4214, P2_U4215, P2_U4216, P2_U4217, P2_U4218, P2_U4219, P2_U4220, P2_U4221, P2_U4222, P2_U4223, P2_U4224, P2_U4225, P2_U4226, P2_U4227, P2_U4228, P2_U4229, P2_U4230, P2_U4231, P2_U4232, P2_U4233, P2_U4234, P2_U4235, P2_U4236, P2_U4237, P2_U4238, P2_U4239, P2_U4240, P2_U4241, P2_U4242, P2_U4243, P2_U4244, P2_U4245, P2_U4246, P2_U4247, P2_U4248, P2_U4249, P2_U4250, P2_U4251, P2_U4252, P2_U4253, P2_U4254, P2_U4255, P2_U4256, P2_U4257, P2_U4258, P2_U4259, P2_U4260, P2_U4261, P2_U4262, P2_U4263, P2_U4264, P2_U4265, P2_U4266, P2_U4267, P2_U4268, P2_U4269, P2_U4270, P2_U4271, P2_U4272, P2_U4273, P2_U4274, P2_U4275, P2_U4276, P2_U4277, P2_U4278, P2_U4279, P2_U4280, P2_U4281, P2_U4282, P2_U4283, P2_U4284, P2_U4285, P2_U4286, P2_U4287, P2_U4288, P2_U4289, P2_U4290, P2_U4291, P2_U4292, P2_U4293, P2_U4294, P2_U4295, P2_U4296, P2_U4297, P2_U4298, P2_U4299, P2_U4300, P2_U4301, P2_U4302, P2_U4303, P2_U4304, P2_U4305, P2_U4306, P2_U4307, P2_U4308, P2_U4309, P2_U4310, P2_U4311, P2_U4312, P2_U4313, P2_U4314, P2_U4315, P2_U4316, P2_U4317, P2_U4318, P2_U4319, P2_U4320, P2_U4321, P2_U4322, P2_U4323, P2_U4324, P2_U4325, P2_U4326, P2_U4327, P2_U4328, P2_U4329, P2_U4330, P2_U4331, P2_U4332, P2_U4333, P2_U4334, P2_U4335, P2_U4336, P2_U4337, P2_U4338, P2_U4339, P2_U4340, P2_U4341, P2_U4342, P2_U4343, P2_U4344, P2_U4345, P2_U4346, P2_U4347, P2_U4348, P2_U4349, P2_U4350, P2_U4351, P2_U4352, P2_U4353, P2_U4354, P2_U4355, P2_U4356, P2_U4357, P2_U4358, P2_U4359, P2_U4360, P2_U4361, P2_U4362, P2_U4363, P2_U4364, P2_U4365, P2_U4366, P2_U4367, P2_U4368, P2_U4369, P2_U4370, P2_U4371, P2_U4372, P2_U4373, P2_U4374, P2_U4375, P2_U4376, P2_U4377, P2_U4378, P2_U4379, P2_U4380, P2_U4381, P2_U4382, P2_U4383, P2_U4384, P2_U4385, P2_U4386, P2_U4387, P2_U4388, P2_U4389, P2_U4390, P2_U4391, P2_U4392, P2_U4393, P2_U4394, P2_U4395, P2_U4396, P2_U4397, P2_U4398, P2_U4399, P2_U4400, P2_U4401, P2_U4402, P2_U4403, P2_U4404, P2_U4405, P2_U4406, P2_U4407, P2_U4408, P2_U4409, P2_U4410, P2_U4411, P2_U4412, P2_U4413, P2_U4414, P2_U4415, P2_U4416, P2_U4417, P2_U4418, P2_U4419, P2_U4420, P2_U4421, P2_U4422, P2_U4423, P2_U4424, P2_U4425, P2_U4426, P2_U4427, P2_U4428, P2_U4429, P2_U4430, P2_U4431, P2_U4432, P2_U4433, P2_U4434, P2_U4435, P2_U4436, P2_U4437, P2_U4438, P2_U4439, P2_U4440, P2_U4441, P2_U4442, P2_U4443, P2_U4444, P2_U4445, P2_U4446, P2_U4447, P2_U4448, P2_U4449, P2_U4450, P2_U4451, P2_U4452, P2_U4453, P2_U4454, P2_U4455, P2_U4456, P2_U4457, P2_U4458, P2_U4459, P2_U4460, P2_U4461, P2_U4462, P2_U4463, P2_U4464, P2_U4465, P2_U4466, P2_U4467, P2_U4468, P2_U4469, P2_U4470, P2_U4471, P2_U4472, P2_U4473, P2_U4474, P2_U4475, P2_U4476, P2_U4477, P2_U4478, P2_U4479, P2_U4480, P2_U4481, P2_U4482, P2_U4483, P2_U4484, P2_U4485, P2_U4486, P2_U4487, P2_U4488, P2_U4489, P2_U4490, P2_U4491, P2_U4492, P2_U4493, P2_U4494, P2_U4495, P2_U4496, P2_U4497, P2_U4498, P2_U4499, P2_U4500, P2_U4501, P2_U4502, P2_U4503, P2_U4504, P2_U4505, P2_U4506, P2_U4507, P2_U4508, P2_U4509, P2_U4510, P2_U4511, P2_U4512, P2_U4513, P2_U4514, P2_U4515, P2_U4516, P2_U4517, P2_U4518, P2_U4519, P2_U4520, P2_U4521, P2_U4522, P2_U4523, P2_U4524, P2_U4525, P2_U4526, P2_U4527, P2_U4528, P2_U4529, P2_U4530, P2_U4531, P2_U4532, P2_U4533, P2_U4534, P2_U4535, P2_U4536, P2_U4537, P2_U4538, P2_U4539, P2_U4540, P2_U4541, P2_U4542, P2_U4543, P2_U4544, P2_U4545, P2_U4546, P2_U4547, P2_U4548, P2_U4549, P2_U4550, P2_U4551, P2_U4552, P2_U4553, P2_U4554, P2_U4555, P2_U4556, P2_U4557, P2_U4558, P2_U4559, P2_U4560, P2_U4561, P2_U4562, P2_U4563, P2_U4564, P2_U4565, P2_U4566, P2_U4567, P2_U4568, P2_U4569, P2_U4570, P2_U4571, P2_U4572, P2_U4573, P2_U4574, P2_U4575, P2_U4576, P2_U4577, P2_U4578, P2_U4579, P2_U4580, P2_U4581, P2_U4582, P2_U4583, P2_U4584, P2_U4585, P2_U4586, P2_U4587, P2_U4588, P2_U4589, P2_U4590, P2_U4591, P2_U4592, P2_U4593, P2_U4594, P2_U4595, P2_U4596, P2_U4597, P2_U4598, P2_U4599, P2_U4600, P2_U4601, P2_U4602, P2_U4603, P2_U4604, P2_U4605, P2_U4606, P2_U4607, P2_U4608, P2_U4609, P2_U4610, P2_U4611, P2_U4612, P2_U4613, P2_U4614, P2_U4615, P2_U4616, P2_U4617, P2_U4618, P2_U4619, P2_U4620, P2_U4621, P2_U4622, P2_U4623, P2_U4624, P2_U4625, P2_U4626, P2_U4627, P2_U4628, P2_U4629, P2_U4630, P2_U4631, P2_U4632, P2_U4633, P2_U4634, P2_U4635, P2_U4636, P2_U4637, P2_U4638, P2_U4639, P2_U4640, P2_U4641, P2_U4642, P2_U4643, P2_U4644, P2_U4645, P2_U4646, P2_U4647, P2_U4648, P2_U4649, P2_U4650, P2_U4651, P2_U4652, P2_U4653, P2_U4654, P2_U4655, P2_U4656, P2_U4657, P2_U4658, P2_U4659, P2_U4660, P2_U4661, P2_U4662, P2_U4663, P2_U4664, P2_U4665, P2_U4666, P2_U4667, P2_U4668, P2_U4669, P2_U4670, P2_U4671, P2_U4672, P2_U4673, P2_U4674, P2_U4675, P2_U4676, P2_U4677, P2_U4678, P2_U4679, P2_U4680, P2_U4681, P2_U4682, P2_U4683, P2_U4684, P2_U4685, P2_U4686, P2_U4687, P2_U4688, P2_U4689, P2_U4690, P2_U4691, P2_U4692, P2_U4693, P2_U4694, P2_U4695, P2_U4696, P2_U4697, P2_U4698, P2_U4699, P2_U4700, P2_U4701, P2_U4702, P2_U4703, P2_U4704, P2_U4705, P2_U4706, P2_U4707, P2_U4708, P2_U4709, P2_U4710, P2_U4711, P2_U4712, P2_U4713, P2_U4714, P2_U4715, P2_U4716, P2_U4717, P2_U4718, P2_U4719, P2_U4720, P2_U4721, P2_U4722, P2_U4723, P2_U4724, P2_U4725, P2_U4726, P2_U4727, P2_U4728, P2_U4729, P2_U4730, P2_U4731, P2_U4732, P2_U4733, P2_U4734, P2_U4735, P2_U4736, P2_U4737, P2_U4738, P2_U4739, P2_U4740, P2_U4741, P2_U4742, P2_U4743, P2_U4744, P2_U4745, P2_U4746, P2_U4747, P2_U4748, P2_U4749, P2_U4750, P2_U4751, P2_U4752, P2_U4753, P2_U4754, P2_U4755, P2_U4756, P2_U4757, P2_U4758, P2_U4759, P2_U4760, P2_U4761, P2_U4762, P2_U4763, P2_U4764, P2_U4765, P2_U4766, P2_U4767, P2_U4768, P2_U4769, P2_U4770, P2_U4771, P2_U4772, P2_U4773, P2_U4774, P2_U4775, P2_U4776, P2_U4777, P2_U4778, P2_U4779, P2_U4780, P2_U4781, P2_U4782, P2_U4783, P2_U4784, P2_U4785, P2_U4786, P2_U4787, P2_U4788, P2_U4789, P2_U4790, P2_U4791, P2_U4792, P2_U4793, P2_U4794, P2_U4795, P2_U4796, P2_U4797, P2_U4798, P2_U4799, P2_U4800, P2_U4801, P2_U4802, P2_U4803, P2_U4804, P2_U4805, P2_U4806, P2_U4807, P2_U4808, P2_U4809, P2_U4810, P2_U4811, P2_U4812, P2_U4813, P2_U4814, P2_U4815, P2_U4816, P2_U4817, P2_U4818, P2_U4819, P2_U4820, P2_U4821, P2_U4822, P2_U4823, P2_U4824, P2_U4825, P2_U4826, P2_U4827, P2_U4828, P2_U4829, P2_U4830, P2_U4831, P2_U4832, P2_U4833, P2_U4834, P2_U4835, P2_U4836, P2_U4837, P2_U4838, P2_U4839, P2_U4840, P2_U4841, P2_U4842, P2_U4843, P2_U4844, P2_U4845, P2_U4846, P2_U4847, P2_U4848, P2_U4849, P2_U4850, P2_U4851, P2_U4852, P2_U4853, P2_U4854, P2_U4855, P2_U4856, P2_U4857, P2_U4858, P2_U4859, P2_U4860, P2_U4861, P2_U4862, P2_U4863, P2_U4864, P2_U4865, P2_U4866, P2_U4867, P2_U4868, P2_U4869, P2_U4870, P2_U4871, P2_U4872, P2_U4873, P2_U4874, P2_U4875, P2_U4876, P2_U4877, P2_U4878, P2_U4879, P2_U4880, P2_U4881, P2_U4882, P2_U4883, P2_U4884, P2_U4885, P2_U4886, P2_U4887, P2_U4888, P2_U4889, P2_U4890, P2_U4891, P2_U4892, P2_U4893, P2_U4894, P2_U4895, P2_U4896, P2_U4897, P2_U4898, P2_U4899, P2_U4900, P2_U4901, P2_U4902, P2_U4903, P2_U4904, P2_U4905, P2_U4906, P2_U4907, P2_U4908, P2_U4909, P2_U4910, P2_U4911, P2_U4912, P2_U4913, P2_U4914, P2_U4915, P2_U4916, P2_U4917, P2_U4918, P2_U4919, P2_U4920, P2_U4921, P2_U4922, P2_U4923, P2_U4924, P2_U4925, P2_U4926, P2_U4927, P2_U4928, P2_U4929, P2_U4930, P2_U4931, P2_U4932, P2_U4933, P2_U4934, P2_U4935, P2_U4936, P2_U4937, P2_U4938, P2_U4939, P2_U4940, P2_U4941, P2_U4942, P2_U4943, P2_U4944, P2_U4945, P2_U4946, P2_U4947, P2_U4948, P2_U4949, P2_U4950, P2_U4951, P2_U4952, P2_U4953, P2_U4954, P2_U4955, P2_U4956, P2_U4957, P2_U4958, P2_U4959, P2_U4960, P2_U4961, P2_U4962, P2_U4963, P2_U4964, P2_U4965, P2_U4966, P2_U4967, P2_U4968, P2_U4969, P2_U4970, P2_U4971, P2_U4972, P2_U4973, P2_U4974, P2_U4975, P2_U4976, P2_U4977, P2_U4978, P2_U4979, P2_U4980, P2_U4981, P2_U4982, P2_U4983, P2_U4984, P2_U4985, P2_U4986, P2_U4987, P2_U4988, P2_U4989, P2_U4990, P2_U4991, P2_U4992, P2_U4993, P2_U4994, P2_U4995, P2_U4996, P2_U4997, P2_U4998, P2_U4999, P2_U5000, P2_U5001, P2_U5002, P2_U5003, P2_U5004, P2_U5005, P2_U5006, P2_U5007, P2_U5008, P2_U5009, P2_U5010, P2_U5011, P2_U5012, P2_U5013, P2_U5014, P2_U5015, P2_U5016, P2_U5017, P2_U5018, P2_U5019, P2_U5020, P2_U5021, P2_U5022, P2_U5023, P2_U5024, P2_U5025, P2_U5026, P2_U5027, P2_U5028, P2_U5029, P2_U5030, P2_U5031, P2_U5032, P2_U5033, P2_U5034, P2_U5035, P2_U5036, P2_U5037, P2_U5038, P2_U5039, P2_U5040, P2_U5041, P2_U5042, P2_U5043, P2_U5044, P2_U5045, P2_U5046, P2_U5047, P2_U5048, P2_U5049, P2_U5050, P2_U5051, P2_U5052, P2_U5053, P2_U5054, P2_U5055, P2_U5056, P2_U5057, P2_U5058, P2_U5059, P2_U5060, P2_U5061, P2_U5062, P2_U5063, P2_U5064, P2_U5065, P2_U5066, P2_U5067, P2_U5068, P2_U5069, P2_U5070, P2_U5071, P2_U5072, P2_U5073, P2_U5074, P2_U5075, P2_U5076, P2_U5077, P2_U5078, P2_U5079, P2_U5080, P2_U5081, P2_U5082, P2_U5083, P2_U5084, P2_U5085, P2_U5086, P2_U5087, P2_U5088, P2_U5089, P2_U5090, P2_U5091, P2_U5092, P2_U5093, P2_U5094, P2_U5095, P2_U5096, P2_U5097, P2_U5098, P2_U5099, P2_U5100, P2_U5101, P2_U5102, P2_U5103, P2_U5104, P2_U5105, P2_U5106, P2_U5107, P2_U5108, P2_U5109, P2_U5110, P2_U5111, P2_U5112, P2_U5113, P2_U5114, P2_U5115, P2_U5116, P2_U5117, P2_U5118, P2_U5119, P2_U5120, P2_U5121, P2_U5122, P2_U5123, P2_U5124, P2_U5125, P2_U5126, P2_U5127, P2_U5128, P2_U5129, P2_U5130, P2_U5131, P2_U5132, P2_U5133, P2_U5134, P2_U5135, P2_U5136, P2_U5137, P2_U5138, P2_U5139, P2_U5140, P2_U5141, P2_U5142, P2_U5143, P2_U5144, P2_U5145, P2_U5146, P2_U5147, P2_U5148, P2_U5149, P2_U5150, P2_U5151, P2_U5152, P2_U5153, P2_U5154, P2_U5155, P2_U5156, P2_U5157, P2_U5158, P2_U5159, P2_U5160, P2_U5161, P2_U5162, P2_U5163, P2_U5164, P2_U5165, P2_U5166, P2_U5167, P2_U5168, P2_U5169, P2_U5170, P2_U5171, P2_U5172, P2_U5173, P2_U5174, P2_U5175, P2_U5176, P2_U5177, P2_U5178, P2_U5179, P2_U5180, P2_U5181, P2_U5182, P2_U5183, P2_U5184, P2_U5185, P2_U5186, P2_U5187, P2_U5188, P2_U5189, P2_U5190, P2_U5191, P2_U5192, P2_U5193, P2_U5194, P2_U5195, P2_U5196, P2_U5197, P2_U5198, P2_U5199, P2_U5200, P2_U5201, P2_U5202, P2_U5203, P2_U5204, P2_U5205, P2_U5206, P2_U5207, P2_U5208, P2_U5209, P2_U5210, P2_U5211, P2_U5212, P2_U5213, P2_U5214, P2_U5215, P2_U5216, P2_U5217, P2_U5218, P2_U5219, P2_U5220, P2_U5221, P2_U5222, P2_U5223, P2_U5224, P2_U5225, P2_U5226, P2_U5227, P2_U5228, P2_U5229, P2_U5230, P2_U5231, P2_U5232, P2_U5233, P2_U5234, P2_U5235, P2_U5236, P2_U5237, P2_U5238, P2_U5239, P2_U5240, P2_U5241, P2_U5242, P2_U5243, P2_U5244, P2_U5245, P2_U5246, P2_U5247, P2_U5248, P2_U5249, P2_U5250, P2_U5251, P2_U5252, P2_U5253, P2_U5254, P2_U5255, P2_U5256, P2_U5257, P2_U5258, P2_U5259, P2_U5260, P2_U5261, P2_U5262, P2_U5263, P2_U5264, P2_U5265, P2_U5266, P2_U5267, P2_U5268, P2_U5269, P2_U5270, P2_U5271, P2_U5272, P2_U5273, P2_U5274, P2_U5275, P2_U5276, P2_U5277, P2_U5278, P2_U5279, P2_U5280, P2_U5281, P2_U5282, P2_U5283, P2_U5284, P2_U5285, P2_U5286, P2_U5287, P2_U5288, P2_U5289, P2_U5290, P2_U5291, P2_U5292, P2_U5293, P2_U5294, P2_U5295, P2_U5296, P2_U5297, P2_U5298, P2_U5299, P2_U5300, P2_U5301, P2_U5302, P2_U5303, P2_U5304, P2_U5305, P2_U5306, P2_U5307, P2_U5308, P2_U5309, P2_U5310, P2_U5311, P2_U5312, P2_U5313, P2_U5314, P2_U5315, P2_U5316, P2_U5317, P2_U5318, P2_U5319, P2_U5320, P2_U5321, P2_U5322, P2_U5323, P2_U5324, P2_U5325, P2_U5326, P2_U5327, P2_U5328, P2_U5329, P2_U5330, P2_U5331, P2_U5332, P2_U5333, P2_U5334, P2_U5335, P2_U5336, P2_U5337, P2_U5338, P2_U5339, P2_U5340, P2_U5341, P2_U5342, P2_U5343, P2_U5344, P2_U5345, P2_U5346, P2_U5347, P2_U5348, P2_U5349, P2_U5350, P2_U5351, P2_U5352, P2_U5353, P2_U5354, P2_U5355, P2_U5356, P2_U5357, P2_U5358, P2_U5359, P2_U5360, P2_U5361, P2_U5362, P2_U5363, P2_U5364, P2_U5365, P2_U5366, P2_U5367, P2_U5368, P2_U5369, P2_U5370, P2_U5371, P2_U5372, P2_U5373, P2_U5374, P2_U5375, P2_U5376, P2_U5377, P2_U5378, P2_U5379, P2_U5380, P2_U5381, P2_U5382, P2_U5383, P2_U5384, P2_U5385, P2_U5386, P2_U5387, P2_U5388, P2_U5389, P2_U5390, P2_U5391, P2_U5392, P2_U5393, P2_U5394, P2_U5395, P2_U5396, P2_U5397, P2_U5398, P2_U5399, P2_U5400, P2_U5401, P2_U5402, P2_U5403, P2_U5404, P2_U5405, P2_U5406, P2_U5407, P2_U5408, P2_U5409, P2_U5410, P2_U5411, P2_U5412, P2_U5413, P2_U5414, P2_U5415, P2_U5416, P2_U5417, P2_U5418, P2_U5419, P2_U5420, P2_U5421, P2_U5422, P2_U5423, P2_U5424, P2_U5425, P2_U5426, P2_U5427, P2_U5428, P2_U5429, P2_U5430, P2_U5431, P2_U5432, P2_U5433, P2_U5434, P2_U5435, P2_U5436, P2_U5437, P2_U5438, P2_U5439, P2_U5440, P2_U5441, P2_U5442, P2_U5443, P2_U5444, P2_U5445, P2_U5446, P2_U5447, P2_U5448, P2_U5449, P2_U5450, P2_U5451, P2_U5452, P2_U5453, P2_U5454, P2_U5455, P2_U5456, P2_U5457, P2_U5458, P2_U5459, P2_U5460, P2_U5461, P2_U5462, P2_U5463, P2_U5464, P2_U5465, P2_U5466, P2_U5467, P2_U5468, P2_U5469, P2_U5470, P2_U5471, P2_U5472, P2_U5473, P2_U5474, P2_U5475, P2_U5476, P2_U5477, P2_U5478, P2_U5479, P2_U5480, P2_U5481, P2_U5482, P2_U5483, P2_U5484, P2_U5485, P2_U5486, P2_U5487, P2_U5488, P2_U5489, P2_U5490, P2_U5491, P2_U5492, P2_U5493, P2_U5494, P2_U5495, P2_U5496, P2_U5497, P2_U5498, P2_U5499, P2_U5500, P2_U5501, P2_U5502, P2_U5503, P2_U5504, P2_U5505, P2_U5506, P2_U5507, P2_U5508, P2_U5509, P2_U5510, P2_U5511, P2_U5512, P2_U5513, P2_U5514, P2_U5515, P2_U5516, P2_U5517, P2_U5518, P2_U5519, P2_U5520, P2_U5521, P2_U5522, P2_U5523, P2_U5524, P2_U5525, P2_U5526, P2_U5527, P2_U5528, P2_U5529, P2_U5530, P2_U5531, P2_U5532, P2_U5533, P2_U5534, P2_U5535, P2_U5536, P2_U5537, P2_U5538, P2_U5539, P2_U5540, P2_U5541, P2_U5542, P2_U5543, P2_U5544, P2_U5545, P2_U5546, P2_U5547, P2_U5548, P2_U5549, P2_U5550, P2_U5551, P2_U5552, P2_U5553, P2_U5554, P2_U5555, P2_U5556, P2_U5557, P2_U5558, P2_U5559, P2_U5560, P2_U5561, P2_U5562, P2_U5563, P2_U5564, P2_U5565, P2_U5566, P2_U5567, P2_U5568, P2_U5569, P2_U5570, P2_U5571, P2_U5572, P2_U5573, P2_U5574, P2_U5575, P2_U5576, P2_U5577, P2_U5578, P2_U5579, P2_U5580, P2_U5581, P2_U5582, P2_U5583, P2_U5584, P2_U5585, P2_U5586, P2_U5587, P2_U5588, P2_U5589, P2_U5590, P2_U5591, P2_U5592, P2_U5593, P2_U5594, P2_U5595, P2_U5596, P2_U5597, P2_U5598, P2_U5599, P2_U5600, P2_U5601, P2_U5602, P2_U5603, P2_U5604, P2_U5605, P2_U5606, P2_U5607, P2_U5608, P2_U5609, P2_U5610, P2_U5611, P2_U5612, P2_U5613, P2_U5614, P2_U5615, P2_U5616, P2_U5617, P2_U5618, P2_U5619, P2_U5620, P2_U5621, P2_U5622, P2_U5623, P2_U5624, P2_U5625, P2_U5626, P2_U5627, P2_U5628, P2_U5629, P2_U5630, P2_U5631, P2_U5632, P2_U5633, P2_U5634, P2_U5635, P2_U5636, P2_U5637, P2_U5638, P2_U5639, P2_U5640, P2_U5641, P2_U5642, P2_U5643, P2_U5644, P2_U5645, P2_U5646, P2_U5647, P2_U5648, P2_U5649, P2_U5650, P2_U5651, P2_U5652, P2_U5653, P2_U5654, P2_U5655, P2_U5656, P2_U5657, P2_U5658, P2_U5659, P2_U5660, P2_U5661, P2_U5662, P2_U5663, P2_U5664, P2_U5665, P2_U5666, P2_U5667, P2_U5668, P2_U5669, P2_U5670, P2_U5671, P2_U5672, P2_U5673, P2_U5674, P2_U5675, P2_U5676, P2_U5677, P2_U5678, P2_U5679, P2_U5680, P2_U5681, P2_U5682, P2_U5683, P2_U5684, P2_U5685, P2_U5686, P2_U5687, P2_U5688, P2_U5689, P2_U5690, P2_U5691, P2_U5692, P2_U5693, P2_U5694, P2_U5695, P2_U5696, P2_U5697, P2_U5698, P2_U5699, P2_U5700, P2_U5701, P2_U5702, P2_U5703, P2_U5704, P2_U5705, P2_U5706, P2_U5707, P2_U5708, P2_U5709, P2_U5710, P2_U5711, P2_U5712, P2_U5713, P2_U5714, P2_U5715, P2_U5716, P2_U5717, P2_U5718, P2_U5719, P2_U5720, P2_U5721, P2_U5722, P2_U5723, P2_U5724, P2_U5725, P2_U5726, P2_U5727, P2_U5728, P2_U5729, P2_U5730, P2_U5731, P2_U5732, P2_U5733, P2_U5734, P2_U5735, P2_U5736, P2_U5737, P2_U5738, P2_U5739, P2_U5740, P2_U5741, P2_U5742, P2_U5743, P2_U5744, P2_U5745, P2_U5746, P2_U5747, P2_U5748, P2_U5749, P2_U5750, P2_U5751, P2_U5752, P2_U5753, P2_U5754, P2_U5755, P2_U5756, P2_U5757, P2_U5758, P2_U5759, P2_U5760, P2_U5761, P2_U5762, P2_U5763, P2_U5764, P2_U5765, P2_U5766, P2_U5767, P2_U5768, P2_U5769, P2_U5770, P2_U5771, P2_U5772, P2_U5773, P2_U5774, P2_U5775, P2_U5776, P2_U5777, P2_U5778, P2_U5779, P2_U5780, P2_U5781, P2_U5782, P2_U5783, P2_U5784, P2_U5785, P2_U5786, P2_U5787, P2_U5788, P2_U5789, P2_U5790, P2_U5791, P2_U5792, P2_U5793, P2_U5794, P2_U5795, P2_U5796, P2_U5797, P2_U5798, P2_U5799, P2_U5800, P2_U5801, P2_U5802, P2_U5803, P2_U5804, P2_U5805, P2_U5806, P2_U5807, P2_U5808, P2_U5809, P2_U5810, P2_U5811, P2_U5812, P2_U5813, P2_U5814, P2_U5815, P2_U5816, P2_U5817, P2_U5818, P2_U5819, P2_U5820, P2_U5821, P2_U5822, P2_U5823, P2_U5824, P2_U5825, P2_U5826, P2_U5827, P2_U5828, P2_U5829, P2_U5830, P2_U5831, P2_U5832, P2_U5833, P2_U5834, P2_U5835, P2_U5836, P2_U5837, P2_U5838, P2_U5839, P2_U5840, P2_U5841, P2_U5842, P2_U5843, P2_U5844, P2_U5845, P2_U5846, P2_U5847, P2_U5848, P2_U5849, P2_U5850, P2_U5851, P2_U5852, P2_U5853, P2_U5854, P2_U5855, P2_U5856, P2_U5857, P2_U5858, P2_U5859, P2_U5860, P2_U5861, P2_U5862, P2_U5863, P2_U5864, P2_U5865, P2_U5866, P2_U5867, P2_U5868, P2_U5869, P2_U5870, P2_U5871, P2_U5872, P2_U5873, P2_U5874, P2_U5875, P2_U5876, P2_U5877, P2_U5878, P2_U5879, P2_U5880, P2_U5881, P2_U5882, P2_U5883, P2_U5884, P2_U5885, P2_U5886, P2_U5887, P2_U5888, P2_U5889, P2_U5890, P2_U5891, P2_U5892, P2_U5893, P2_U5894, P2_U5895, P2_U5896, P2_U5897, P2_U5898, P2_U5899, P2_U5900, P2_U5901, P2_U5902, P2_U5903, P2_U5904, P2_U5905, P2_U5906, P2_U5907, P2_U5908, P2_U5909, P2_U5910, P2_U5911, P2_U5912, P2_U5913, P2_U5914, P2_U5915, P2_U5916, P2_U5917, P2_U5918, P2_U5919, P2_U5920, P2_U5921, P2_U5922, P2_U5923, P2_U5924, P2_U5925, P2_U5926, P2_U5927, P2_U5928, P2_U5929, P2_U5930, P2_U5931, P2_U5932, P2_U5933, P2_U5934, P2_U5935, P2_U5936, P2_U5937, P2_U5938, P2_U5939, P2_U5940, P2_U5941, P2_U5942, P2_U5943, P2_U5944, P2_U5945, P2_U5946, P2_U5947, P2_U5948, P2_U5949, P2_U5950, P2_U5951, P2_U5952, P2_U5953, P2_U5954, P2_U5955, P2_U5956, P2_U5957, P2_U5958, P2_U5959, P2_U5960, P2_U5961, P2_U5962, P2_U5963, P2_U5964, P2_U5965, P2_U5966, P2_U5967, P2_U5968, P2_U5969, P2_U5970, P2_U5971, P2_U5972, P2_U5973, P2_U5974, P2_U5975, P2_U5976, P2_U5977, P2_U5978, P2_U5979, P2_U5980, P2_U5981, P2_U5982, P2_U5983, P2_U5984, P2_U5985, P2_U5986, P2_U5987, P2_U5988, P2_U5989, P2_U5990, P2_U5991, P2_U5992, P2_U5993, P2_U5994, P2_U5995, P2_U5996, P2_U5997, P2_U5998, P2_U5999, P2_U6000, P2_U6001, P2_U6002, P2_U6003, P2_U6004, P2_U6005, P2_U6006, P2_U6007, P2_U6008, P2_U6009, P2_U6010, P2_U6011, P2_U6012, P2_U6013, P2_U6014, P2_U6015, P2_U6016, P2_U6017, P2_U6018, P2_U6019, P2_U6020, P2_U6021, P2_U6022, P2_U6023, P2_U6024, P2_U6025, P2_U6026, P2_U6027, P2_U6028, P2_U6029, P2_U6030, P2_U6031, P2_U6032, P2_U6033, P2_U6034, P2_U6035, P2_U6036, P2_U6037, P2_U6038, P2_U6039, P2_U6040, P2_U6041, P2_U6042, P2_U6043, P2_U6044, P2_U6045, P2_U6046, P2_U6047, P2_U6048, P2_U6049, P2_U6050, P2_U6051, P2_U6052, P2_U6053, P2_U6054, P2_U6055, P2_U6056, P2_U6057, P2_U6058, P2_U6059, P2_U6060, P2_U6061, P2_U6062, P2_U6063, P2_U6064, P2_U6065, P2_U6066, P2_U6067, P2_U6068, P2_U6069, P2_U6070, P2_U6071, P2_U6072, P2_U6073, P2_U6074, P2_U6075, P2_U6076, P2_U6077, P2_U6078, P2_U6079, P2_U6080, P2_U6081, P2_U6082, P2_U6083, P2_U6084, P2_U6085, P2_U6086, P2_U6087, P2_U6088, P2_U6089, P2_U6090, P2_U6091, P2_U6092, P2_U6093, P2_U6094, P2_U6095, P2_U6096, P2_U6097, P2_U6098, P2_U6099, P2_U6100, P2_U6101, P2_U6102, P2_U6103, P2_U6104, P2_U6105, P2_U6106, P2_U6107, P2_U6108, P2_U6109, P2_U6110, P2_U6111, P2_U6112, P2_U6113, P2_U6114, P2_U6115, P2_U6116, P2_U6117, P2_U6118, P2_U6119, P2_U6120, P2_U6121, P2_U6122, P2_U6123, P2_U6124, P2_U6125, P2_U6126, P2_U6127, P2_U6128, P2_U6129, P2_U6130, P2_U6131, P2_U6132, P2_U6133, P2_U6134, P2_U6135, P2_U6136, P2_U6137, P2_U6138, P2_U6139, P2_U6140, P2_U6141, P2_U6142, P2_U6143, P2_U6144, P2_U6145, P2_U6146, P2_U6147, P2_U6148, P2_U6149, P2_U6150, P3_R1054_U10, P3_R1054_U100, P3_R1054_U101, P3_R1054_U102, P3_R1054_U103, P3_R1054_U104, P3_R1054_U105, P3_R1054_U106, P3_R1054_U107, P3_R1054_U108, P3_R1054_U109, P3_R1054_U11, P3_R1054_U110, P3_R1054_U111, P3_R1054_U112, P3_R1054_U113, P3_R1054_U114, P3_R1054_U115, P3_R1054_U116, P3_R1054_U117, P3_R1054_U118, P3_R1054_U119, P3_R1054_U12, P3_R1054_U120, P3_R1054_U121, P3_R1054_U122, P3_R1054_U123, P3_R1054_U124, P3_R1054_U125, P3_R1054_U126, P3_R1054_U127, P3_R1054_U128, P3_R1054_U129, P3_R1054_U13, P3_R1054_U130, P3_R1054_U131, P3_R1054_U132, P3_R1054_U133, P3_R1054_U134, P3_R1054_U135, P3_R1054_U136, P3_R1054_U137, P3_R1054_U138, P3_R1054_U139, P3_R1054_U14, P3_R1054_U140, P3_R1054_U141, P3_R1054_U142, P3_R1054_U143, P3_R1054_U144, P3_R1054_U145, P3_R1054_U146, P3_R1054_U147, P3_R1054_U148, P3_R1054_U149, P3_R1054_U15, P3_R1054_U150, P3_R1054_U151, P3_R1054_U152, P3_R1054_U153, P3_R1054_U154, P3_R1054_U155, P3_R1054_U156, P3_R1054_U157, P3_R1054_U158, P3_R1054_U159, P3_R1054_U16, P3_R1054_U160, P3_R1054_U161, P3_R1054_U162, P3_R1054_U163, P3_R1054_U164, P3_R1054_U165, P3_R1054_U166, P3_R1054_U167, P3_R1054_U168, P3_R1054_U169, P3_R1054_U17, P3_R1054_U170, P3_R1054_U171, P3_R1054_U172, P3_R1054_U173, P3_R1054_U174, P3_R1054_U175, P3_R1054_U176, P3_R1054_U177, P3_R1054_U178, P3_R1054_U179, P3_R1054_U18, P3_R1054_U180, P3_R1054_U181, P3_R1054_U182, P3_R1054_U183, P3_R1054_U184, P3_R1054_U185, P3_R1054_U186, P3_R1054_U187, P3_R1054_U188, P3_R1054_U189, P3_R1054_U19, P3_R1054_U190, P3_R1054_U191, P3_R1054_U192, P3_R1054_U193, P3_R1054_U194, P3_R1054_U195, P3_R1054_U196, P3_R1054_U197, P3_R1054_U198, P3_R1054_U199, P3_R1054_U20, P3_R1054_U200, P3_R1054_U201, P3_R1054_U202, P3_R1054_U203, P3_R1054_U204, P3_R1054_U205, P3_R1054_U206, P3_R1054_U207, P3_R1054_U208, P3_R1054_U209, P3_R1054_U21, P3_R1054_U210, P3_R1054_U211, P3_R1054_U212, P3_R1054_U213, P3_R1054_U214, P3_R1054_U215, P3_R1054_U216, P3_R1054_U217, P3_R1054_U218, P3_R1054_U219, P3_R1054_U22, P3_R1054_U220, P3_R1054_U221, P3_R1054_U222, P3_R1054_U223, P3_R1054_U224, P3_R1054_U225, P3_R1054_U226, P3_R1054_U227, P3_R1054_U228, P3_R1054_U229, P3_R1054_U23, P3_R1054_U230, P3_R1054_U231, P3_R1054_U232, P3_R1054_U233, P3_R1054_U234, P3_R1054_U235, P3_R1054_U236, P3_R1054_U237, P3_R1054_U238, P3_R1054_U239, P3_R1054_U24, P3_R1054_U240, P3_R1054_U241, P3_R1054_U242, P3_R1054_U243, P3_R1054_U244, P3_R1054_U245, P3_R1054_U246, P3_R1054_U247, P3_R1054_U248, P3_R1054_U249, P3_R1054_U25, P3_R1054_U250, P3_R1054_U251, P3_R1054_U252, P3_R1054_U253, P3_R1054_U254, P3_R1054_U255, P3_R1054_U256, P3_R1054_U257, P3_R1054_U258, P3_R1054_U259, P3_R1054_U26, P3_R1054_U260, P3_R1054_U261, P3_R1054_U262, P3_R1054_U263, P3_R1054_U264, P3_R1054_U265, P3_R1054_U266, P3_R1054_U267, P3_R1054_U268, P3_R1054_U269, P3_R1054_U27, P3_R1054_U270, P3_R1054_U271, P3_R1054_U272, P3_R1054_U273, P3_R1054_U274, P3_R1054_U275, P3_R1054_U276, P3_R1054_U277, P3_R1054_U278, P3_R1054_U279, P3_R1054_U28, P3_R1054_U280, P3_R1054_U281, P3_R1054_U282, P3_R1054_U283, P3_R1054_U284, P3_R1054_U285, P3_R1054_U286, P3_R1054_U287, P3_R1054_U288, P3_R1054_U289, P3_R1054_U29, P3_R1054_U290, P3_R1054_U291, P3_R1054_U292, P3_R1054_U293, P3_R1054_U294, P3_R1054_U30, P3_R1054_U31, P3_R1054_U32, P3_R1054_U33, P3_R1054_U34, P3_R1054_U35, P3_R1054_U36, P3_R1054_U37, P3_R1054_U38, P3_R1054_U39, P3_R1054_U40, P3_R1054_U41, P3_R1054_U42, P3_R1054_U43, P3_R1054_U44, P3_R1054_U45, P3_R1054_U46, P3_R1054_U47, P3_R1054_U48, P3_R1054_U49, P3_R1054_U50, P3_R1054_U51, P3_R1054_U52, P3_R1054_U53, P3_R1054_U54, P3_R1054_U55, P3_R1054_U56, P3_R1054_U57, P3_R1054_U58, P3_R1054_U59, P3_R1054_U6, P3_R1054_U60, P3_R1054_U61, P3_R1054_U62, P3_R1054_U63, P3_R1054_U64, P3_R1054_U65, P3_R1054_U66, P3_R1054_U67, P3_R1054_U68, P3_R1054_U69, P3_R1054_U7, P3_R1054_U70, P3_R1054_U71, P3_R1054_U72, P3_R1054_U73, P3_R1054_U74, P3_R1054_U75, P3_R1054_U76, P3_R1054_U77, P3_R1054_U78, P3_R1054_U79, P3_R1054_U8, P3_R1054_U80, P3_R1054_U81, P3_R1054_U82, P3_R1054_U83, P3_R1054_U84, P3_R1054_U85, P3_R1054_U86, P3_R1054_U87, P3_R1054_U88, P3_R1054_U89, P3_R1054_U9, P3_R1054_U90, P3_R1054_U91, P3_R1054_U92, P3_R1054_U93, P3_R1054_U94, P3_R1054_U95, P3_R1054_U96, P3_R1054_U97, P3_R1054_U98, P3_R1054_U99, P3_R1077_U10, P3_R1077_U100, P3_R1077_U101, P3_R1077_U102, P3_R1077_U103, P3_R1077_U104, P3_R1077_U105, P3_R1077_U106, P3_R1077_U107, P3_R1077_U108, P3_R1077_U109, P3_R1077_U11, P3_R1077_U110, P3_R1077_U111, P3_R1077_U112, P3_R1077_U113, P3_R1077_U114, P3_R1077_U115, P3_R1077_U116, P3_R1077_U117, P3_R1077_U118, P3_R1077_U119, P3_R1077_U12, P3_R1077_U120, P3_R1077_U121, P3_R1077_U122, P3_R1077_U123, P3_R1077_U124, P3_R1077_U125, P3_R1077_U126, P3_R1077_U127, P3_R1077_U128, P3_R1077_U129, P3_R1077_U13, P3_R1077_U130, P3_R1077_U131, P3_R1077_U132, P3_R1077_U133, P3_R1077_U134, P3_R1077_U135, P3_R1077_U136, P3_R1077_U137, P3_R1077_U138, P3_R1077_U139, P3_R1077_U14, P3_R1077_U140, P3_R1077_U141, P3_R1077_U142, P3_R1077_U143, P3_R1077_U144, P3_R1077_U145, P3_R1077_U146, P3_R1077_U147, P3_R1077_U148, P3_R1077_U149, P3_R1077_U15, P3_R1077_U150, P3_R1077_U151, P3_R1077_U152, P3_R1077_U153, P3_R1077_U154, P3_R1077_U155, P3_R1077_U156, P3_R1077_U157, P3_R1077_U158, P3_R1077_U159, P3_R1077_U16, P3_R1077_U160, P3_R1077_U161, P3_R1077_U162, P3_R1077_U163, P3_R1077_U164, P3_R1077_U165, P3_R1077_U166, P3_R1077_U167, P3_R1077_U168, P3_R1077_U169, P3_R1077_U17, P3_R1077_U170, P3_R1077_U171, P3_R1077_U172, P3_R1077_U173, P3_R1077_U174, P3_R1077_U175, P3_R1077_U176, P3_R1077_U177, P3_R1077_U178, P3_R1077_U179, P3_R1077_U18, P3_R1077_U180, P3_R1077_U181, P3_R1077_U182, P3_R1077_U183, P3_R1077_U184, P3_R1077_U185, P3_R1077_U186, P3_R1077_U187, P3_R1077_U188, P3_R1077_U189, P3_R1077_U19, P3_R1077_U190, P3_R1077_U191, P3_R1077_U192, P3_R1077_U193, P3_R1077_U194, P3_R1077_U195, P3_R1077_U196, P3_R1077_U197, P3_R1077_U198, P3_R1077_U199, P3_R1077_U20, P3_R1077_U200, P3_R1077_U201, P3_R1077_U202, P3_R1077_U203, P3_R1077_U204, P3_R1077_U205, P3_R1077_U206, P3_R1077_U207, P3_R1077_U208, P3_R1077_U209, P3_R1077_U21, P3_R1077_U210, P3_R1077_U211, P3_R1077_U212, P3_R1077_U213, P3_R1077_U214, P3_R1077_U215, P3_R1077_U216, P3_R1077_U217, P3_R1077_U218, P3_R1077_U219, P3_R1077_U22, P3_R1077_U220, P3_R1077_U221, P3_R1077_U222, P3_R1077_U223, P3_R1077_U224, P3_R1077_U225, P3_R1077_U226, P3_R1077_U227, P3_R1077_U228, P3_R1077_U229, P3_R1077_U23, P3_R1077_U230, P3_R1077_U231, P3_R1077_U232, P3_R1077_U233, P3_R1077_U234, P3_R1077_U235, P3_R1077_U236, P3_R1077_U237, P3_R1077_U238, P3_R1077_U239, P3_R1077_U24, P3_R1077_U240, P3_R1077_U241, P3_R1077_U242, P3_R1077_U243, P3_R1077_U244, P3_R1077_U245, P3_R1077_U246, P3_R1077_U247, P3_R1077_U248, P3_R1077_U249, P3_R1077_U25, P3_R1077_U250, P3_R1077_U251, P3_R1077_U252, P3_R1077_U253, P3_R1077_U254, P3_R1077_U255, P3_R1077_U256, P3_R1077_U257, P3_R1077_U258, P3_R1077_U259, P3_R1077_U26, P3_R1077_U260, P3_R1077_U261, P3_R1077_U262, P3_R1077_U263, P3_R1077_U264, P3_R1077_U265, P3_R1077_U266, P3_R1077_U267, P3_R1077_U268, P3_R1077_U269, P3_R1077_U27, P3_R1077_U270, P3_R1077_U271, P3_R1077_U272, P3_R1077_U273, P3_R1077_U274, P3_R1077_U275, P3_R1077_U276, P3_R1077_U277, P3_R1077_U278, P3_R1077_U279, P3_R1077_U28, P3_R1077_U280, P3_R1077_U281, P3_R1077_U282, P3_R1077_U283, P3_R1077_U284, P3_R1077_U285, P3_R1077_U286, P3_R1077_U287, P3_R1077_U288, P3_R1077_U289, P3_R1077_U29, P3_R1077_U290, P3_R1077_U291, P3_R1077_U292, P3_R1077_U293, P3_R1077_U294, P3_R1077_U295, P3_R1077_U296, P3_R1077_U297, P3_R1077_U298, P3_R1077_U299, P3_R1077_U30, P3_R1077_U300, P3_R1077_U301, P3_R1077_U302, P3_R1077_U303, P3_R1077_U304, P3_R1077_U305, P3_R1077_U306, P3_R1077_U307, P3_R1077_U308, P3_R1077_U309, P3_R1077_U31, P3_R1077_U310, P3_R1077_U311, P3_R1077_U312, P3_R1077_U313, P3_R1077_U314, P3_R1077_U315, P3_R1077_U316, P3_R1077_U317, P3_R1077_U318, P3_R1077_U319, P3_R1077_U32, P3_R1077_U320, P3_R1077_U321, P3_R1077_U322, P3_R1077_U323, P3_R1077_U324, P3_R1077_U325, P3_R1077_U326, P3_R1077_U327, P3_R1077_U328, P3_R1077_U329, P3_R1077_U33, P3_R1077_U330, P3_R1077_U331, P3_R1077_U332, P3_R1077_U333, P3_R1077_U334, P3_R1077_U335, P3_R1077_U336, P3_R1077_U337, P3_R1077_U338, P3_R1077_U339, P3_R1077_U34, P3_R1077_U340, P3_R1077_U341, P3_R1077_U342, P3_R1077_U343, P3_R1077_U344, P3_R1077_U345, P3_R1077_U346, P3_R1077_U347, P3_R1077_U348, P3_R1077_U349, P3_R1077_U35, P3_R1077_U350, P3_R1077_U351, P3_R1077_U352, P3_R1077_U353, P3_R1077_U354, P3_R1077_U355, P3_R1077_U356, P3_R1077_U357, P3_R1077_U358, P3_R1077_U359, P3_R1077_U36, P3_R1077_U360, P3_R1077_U361, P3_R1077_U362, P3_R1077_U363, P3_R1077_U364, P3_R1077_U365, P3_R1077_U366, P3_R1077_U367, P3_R1077_U368, P3_R1077_U369, P3_R1077_U37, P3_R1077_U370, P3_R1077_U371, P3_R1077_U372, P3_R1077_U373, P3_R1077_U374, P3_R1077_U375, P3_R1077_U376, P3_R1077_U377, P3_R1077_U378, P3_R1077_U379, P3_R1077_U38, P3_R1077_U380, P3_R1077_U381, P3_R1077_U382, P3_R1077_U383, P3_R1077_U384, P3_R1077_U385, P3_R1077_U386, P3_R1077_U387, P3_R1077_U388, P3_R1077_U389, P3_R1077_U39, P3_R1077_U390, P3_R1077_U391, P3_R1077_U392, P3_R1077_U393, P3_R1077_U394, P3_R1077_U395, P3_R1077_U396, P3_R1077_U397, P3_R1077_U398, P3_R1077_U399, P3_R1077_U4, P3_R1077_U40, P3_R1077_U400, P3_R1077_U401, P3_R1077_U402, P3_R1077_U403, P3_R1077_U404, P3_R1077_U405, P3_R1077_U406, P3_R1077_U407, P3_R1077_U408, P3_R1077_U409, P3_R1077_U41, P3_R1077_U410, P3_R1077_U411, P3_R1077_U412, P3_R1077_U413, P3_R1077_U414, P3_R1077_U415, P3_R1077_U416, P3_R1077_U417, P3_R1077_U418, P3_R1077_U419, P3_R1077_U42, P3_R1077_U420, P3_R1077_U421, P3_R1077_U422, P3_R1077_U423, P3_R1077_U424, P3_R1077_U425, P3_R1077_U426, P3_R1077_U427, P3_R1077_U428, P3_R1077_U429, P3_R1077_U43, P3_R1077_U430, P3_R1077_U431, P3_R1077_U432, P3_R1077_U433, P3_R1077_U434, P3_R1077_U435, P3_R1077_U436, P3_R1077_U437, P3_R1077_U438, P3_R1077_U439, P3_R1077_U44, P3_R1077_U440, P3_R1077_U441, P3_R1077_U442, P3_R1077_U443, P3_R1077_U444, P3_R1077_U445, P3_R1077_U446, P3_R1077_U447, P3_R1077_U448, P3_R1077_U449, P3_R1077_U45, P3_R1077_U450, P3_R1077_U451, P3_R1077_U452, P3_R1077_U453, P3_R1077_U454, P3_R1077_U455, P3_R1077_U456, P3_R1077_U457, P3_R1077_U458, P3_R1077_U459, P3_R1077_U46, P3_R1077_U460, P3_R1077_U461, P3_R1077_U462, P3_R1077_U463, P3_R1077_U464, P3_R1077_U465, P3_R1077_U466, P3_R1077_U467, P3_R1077_U468, P3_R1077_U469, P3_R1077_U47, P3_R1077_U470, P3_R1077_U471, P3_R1077_U472, P3_R1077_U473, P3_R1077_U474, P3_R1077_U475, P3_R1077_U476, P3_R1077_U477, P3_R1077_U478, P3_R1077_U479, P3_R1077_U48, P3_R1077_U480, P3_R1077_U481, P3_R1077_U482, P3_R1077_U483, P3_R1077_U484, P3_R1077_U485, P3_R1077_U486, P3_R1077_U487, P3_R1077_U488, P3_R1077_U489, P3_R1077_U49, P3_R1077_U490, P3_R1077_U491, P3_R1077_U492, P3_R1077_U493, P3_R1077_U494, P3_R1077_U495, P3_R1077_U496, P3_R1077_U497, P3_R1077_U498, P3_R1077_U499, P3_R1077_U5, P3_R1077_U50, P3_R1077_U500, P3_R1077_U501, P3_R1077_U502, P3_R1077_U503, P3_R1077_U504, P3_R1077_U51, P3_R1077_U52, P3_R1077_U53, P3_R1077_U54, P3_R1077_U55, P3_R1077_U56, P3_R1077_U57, P3_R1077_U58, P3_R1077_U59, P3_R1077_U6, P3_R1077_U60, P3_R1077_U61, P3_R1077_U62, P3_R1077_U63, P3_R1077_U64, P3_R1077_U65, P3_R1077_U66, P3_R1077_U67, P3_R1077_U68, P3_R1077_U69, P3_R1077_U7, P3_R1077_U70, P3_R1077_U71, P3_R1077_U72, P3_R1077_U73, P3_R1077_U74, P3_R1077_U75, P3_R1077_U76, P3_R1077_U77, P3_R1077_U78, P3_R1077_U79, P3_R1077_U8, P3_R1077_U80, P3_R1077_U81, P3_R1077_U82, P3_R1077_U83, P3_R1077_U84, P3_R1077_U85, P3_R1077_U86, P3_R1077_U87, P3_R1077_U88, P3_R1077_U89, P3_R1077_U9, P3_R1077_U90, P3_R1077_U91, P3_R1077_U92, P3_R1077_U93, P3_R1077_U94, P3_R1077_U95, P3_R1077_U96, P3_R1077_U97, P3_R1077_U98, P3_R1077_U99, P3_R1095_U10, P3_R1095_U100, P3_R1095_U101, P3_R1095_U102, P3_R1095_U103, P3_R1095_U104, P3_R1095_U105, P3_R1095_U106, P3_R1095_U107, P3_R1095_U108, P3_R1095_U109, P3_R1095_U11, P3_R1095_U110, P3_R1095_U111, P3_R1095_U112, P3_R1095_U113, P3_R1095_U114, P3_R1095_U115, P3_R1095_U116, P3_R1095_U117, P3_R1095_U118, P3_R1095_U119, P3_R1095_U12, P3_R1095_U120, P3_R1095_U121, P3_R1095_U122, P3_R1095_U123, P3_R1095_U124, P3_R1095_U125, P3_R1095_U126, P3_R1095_U127, P3_R1095_U128, P3_R1095_U129, P3_R1095_U13, P3_R1095_U130, P3_R1095_U131, P3_R1095_U132, P3_R1095_U133, P3_R1095_U134, P3_R1095_U135, P3_R1095_U136, P3_R1095_U137, P3_R1095_U138, P3_R1095_U139, P3_R1095_U14, P3_R1095_U140, P3_R1095_U141, P3_R1095_U142, P3_R1095_U143, P3_R1095_U144, P3_R1095_U145, P3_R1095_U146, P3_R1095_U147, P3_R1095_U148, P3_R1095_U149, P3_R1095_U15, P3_R1095_U150, P3_R1095_U151, P3_R1095_U152, P3_R1095_U153, P3_R1095_U154, P3_R1095_U155, P3_R1095_U156, P3_R1095_U157, P3_R1095_U158, P3_R1095_U159, P3_R1095_U16, P3_R1095_U160, P3_R1095_U161, P3_R1095_U162, P3_R1095_U163, P3_R1095_U164, P3_R1095_U165, P3_R1095_U166, P3_R1095_U167, P3_R1095_U168, P3_R1095_U169, P3_R1095_U17, P3_R1095_U170, P3_R1095_U171, P3_R1095_U172, P3_R1095_U173, P3_R1095_U174, P3_R1095_U175, P3_R1095_U176, P3_R1095_U177, P3_R1095_U178, P3_R1095_U179, P3_R1095_U18, P3_R1095_U180, P3_R1095_U181, P3_R1095_U182, P3_R1095_U183, P3_R1095_U184, P3_R1095_U185, P3_R1095_U186, P3_R1095_U187, P3_R1095_U188, P3_R1095_U189, P3_R1095_U19, P3_R1095_U190, P3_R1095_U191, P3_R1095_U192, P3_R1095_U193, P3_R1095_U194, P3_R1095_U195, P3_R1095_U196, P3_R1095_U197, P3_R1095_U198, P3_R1095_U199, P3_R1095_U20, P3_R1095_U200, P3_R1095_U201, P3_R1095_U202, P3_R1095_U203, P3_R1095_U204, P3_R1095_U205, P3_R1095_U206, P3_R1095_U207, P3_R1095_U208, P3_R1095_U209, P3_R1095_U21, P3_R1095_U210, P3_R1095_U211, P3_R1095_U212, P3_R1095_U213, P3_R1095_U214, P3_R1095_U215, P3_R1095_U216, P3_R1095_U217, P3_R1095_U218, P3_R1095_U219, P3_R1095_U22, P3_R1095_U220, P3_R1095_U221, P3_R1095_U222, P3_R1095_U223, P3_R1095_U224, P3_R1095_U225, P3_R1095_U226, P3_R1095_U227, P3_R1095_U228, P3_R1095_U229, P3_R1095_U23, P3_R1095_U230, P3_R1095_U231, P3_R1095_U232, P3_R1095_U233, P3_R1095_U234, P3_R1095_U235, P3_R1095_U236, P3_R1095_U237, P3_R1095_U238, P3_R1095_U239, P3_R1095_U24, P3_R1095_U240, P3_R1095_U241, P3_R1095_U242, P3_R1095_U243, P3_R1095_U244, P3_R1095_U245, P3_R1095_U246, P3_R1095_U247, P3_R1095_U248, P3_R1095_U249, P3_R1095_U25, P3_R1095_U250, P3_R1095_U251, P3_R1095_U252, P3_R1095_U253, P3_R1095_U254, P3_R1095_U255, P3_R1095_U256, P3_R1095_U257, P3_R1095_U258, P3_R1095_U259, P3_R1095_U26, P3_R1095_U260, P3_R1095_U261, P3_R1095_U262, P3_R1095_U263, P3_R1095_U264, P3_R1095_U265, P3_R1095_U266, P3_R1095_U267, P3_R1095_U268, P3_R1095_U269, P3_R1095_U27, P3_R1095_U270, P3_R1095_U271, P3_R1095_U272, P3_R1095_U273, P3_R1095_U274, P3_R1095_U275, P3_R1095_U276, P3_R1095_U277, P3_R1095_U278, P3_R1095_U279, P3_R1095_U28, P3_R1095_U280, P3_R1095_U281, P3_R1095_U282, P3_R1095_U283, P3_R1095_U284, P3_R1095_U285, P3_R1095_U286, P3_R1095_U287, P3_R1095_U288, P3_R1095_U289, P3_R1095_U29, P3_R1095_U290, P3_R1095_U291, P3_R1095_U292, P3_R1095_U293, P3_R1095_U294, P3_R1095_U295, P3_R1095_U296, P3_R1095_U297, P3_R1095_U298, P3_R1095_U299, P3_R1095_U30, P3_R1095_U300, P3_R1095_U301, P3_R1095_U302, P3_R1095_U303, P3_R1095_U304, P3_R1095_U305, P3_R1095_U306, P3_R1095_U307, P3_R1095_U308, P3_R1095_U309, P3_R1095_U31, P3_R1095_U310, P3_R1095_U311, P3_R1095_U312, P3_R1095_U313, P3_R1095_U314, P3_R1095_U315, P3_R1095_U316, P3_R1095_U317, P3_R1095_U318, P3_R1095_U319, P3_R1095_U32, P3_R1095_U320, P3_R1095_U321, P3_R1095_U322, P3_R1095_U323, P3_R1095_U324, P3_R1095_U325, P3_R1095_U326, P3_R1095_U327, P3_R1095_U328, P3_R1095_U329, P3_R1095_U33, P3_R1095_U330, P3_R1095_U331, P3_R1095_U332, P3_R1095_U333, P3_R1095_U334, P3_R1095_U335, P3_R1095_U336, P3_R1095_U337, P3_R1095_U338, P3_R1095_U339, P3_R1095_U34, P3_R1095_U340, P3_R1095_U341, P3_R1095_U342, P3_R1095_U343, P3_R1095_U344, P3_R1095_U345, P3_R1095_U346, P3_R1095_U347, P3_R1095_U348, P3_R1095_U349, P3_R1095_U35, P3_R1095_U350, P3_R1095_U351, P3_R1095_U352, P3_R1095_U353, P3_R1095_U354, P3_R1095_U355, P3_R1095_U356, P3_R1095_U357, P3_R1095_U358, P3_R1095_U359, P3_R1095_U36, P3_R1095_U360, P3_R1095_U361, P3_R1095_U362, P3_R1095_U363, P3_R1095_U364, P3_R1095_U365, P3_R1095_U366, P3_R1095_U367, P3_R1095_U368, P3_R1095_U369, P3_R1095_U37, P3_R1095_U370, P3_R1095_U371, P3_R1095_U372, P3_R1095_U373, P3_R1095_U374, P3_R1095_U375, P3_R1095_U376, P3_R1095_U377, P3_R1095_U378, P3_R1095_U379, P3_R1095_U38, P3_R1095_U380, P3_R1095_U381, P3_R1095_U382, P3_R1095_U383, P3_R1095_U384, P3_R1095_U385, P3_R1095_U386, P3_R1095_U387, P3_R1095_U388, P3_R1095_U389, P3_R1095_U39, P3_R1095_U390, P3_R1095_U391, P3_R1095_U392, P3_R1095_U393, P3_R1095_U394, P3_R1095_U395, P3_R1095_U396, P3_R1095_U397, P3_R1095_U398, P3_R1095_U399, P3_R1095_U40, P3_R1095_U400, P3_R1095_U401, P3_R1095_U402, P3_R1095_U403, P3_R1095_U404, P3_R1095_U405, P3_R1095_U406, P3_R1095_U407, P3_R1095_U408, P3_R1095_U409, P3_R1095_U41, P3_R1095_U410, P3_R1095_U411, P3_R1095_U412, P3_R1095_U413, P3_R1095_U414, P3_R1095_U415, P3_R1095_U416, P3_R1095_U417, P3_R1095_U418, P3_R1095_U419, P3_R1095_U42, P3_R1095_U420, P3_R1095_U421, P3_R1095_U422, P3_R1095_U423, P3_R1095_U424, P3_R1095_U425, P3_R1095_U426, P3_R1095_U427, P3_R1095_U428, P3_R1095_U429, P3_R1095_U43, P3_R1095_U430, P3_R1095_U431, P3_R1095_U432, P3_R1095_U433, P3_R1095_U434, P3_R1095_U435, P3_R1095_U436, P3_R1095_U437, P3_R1095_U438, P3_R1095_U439, P3_R1095_U44, P3_R1095_U440, P3_R1095_U441, P3_R1095_U442, P3_R1095_U443, P3_R1095_U444, P3_R1095_U445, P3_R1095_U446, P3_R1095_U447, P3_R1095_U448, P3_R1095_U449, P3_R1095_U45, P3_R1095_U450, P3_R1095_U451, P3_R1095_U452, P3_R1095_U453, P3_R1095_U454, P3_R1095_U455, P3_R1095_U456, P3_R1095_U457, P3_R1095_U458, P3_R1095_U459, P3_R1095_U46, P3_R1095_U460, P3_R1095_U461, P3_R1095_U462, P3_R1095_U463, P3_R1095_U464, P3_R1095_U465, P3_R1095_U466, P3_R1095_U467, P3_R1095_U468, P3_R1095_U469, P3_R1095_U47, P3_R1095_U470, P3_R1095_U471, P3_R1095_U472, P3_R1095_U473, P3_R1095_U474, P3_R1095_U475, P3_R1095_U476, P3_R1095_U477, P3_R1095_U478, P3_R1095_U479, P3_R1095_U48, P3_R1095_U480, P3_R1095_U481, P3_R1095_U482, P3_R1095_U483, P3_R1095_U484, P3_R1095_U485, P3_R1095_U49, P3_R1095_U50, P3_R1095_U51, P3_R1095_U52, P3_R1095_U53, P3_R1095_U54, P3_R1095_U55, P3_R1095_U56, P3_R1095_U57, P3_R1095_U58, P3_R1095_U59, P3_R1095_U6, P3_R1095_U60, P3_R1095_U61, P3_R1095_U62, P3_R1095_U63, P3_R1095_U64, P3_R1095_U65, P3_R1095_U66, P3_R1095_U67, P3_R1095_U68, P3_R1095_U69, P3_R1095_U7, P3_R1095_U70, P3_R1095_U71, P3_R1095_U72, P3_R1095_U73, P3_R1095_U74, P3_R1095_U75, P3_R1095_U76, P3_R1095_U77, P3_R1095_U78, P3_R1095_U79, P3_R1095_U8, P3_R1095_U80, P3_R1095_U81, P3_R1095_U82, P3_R1095_U83, P3_R1095_U84, P3_R1095_U85, P3_R1095_U86, P3_R1095_U87, P3_R1095_U88, P3_R1095_U89, P3_R1095_U9, P3_R1095_U90, P3_R1095_U91, P3_R1095_U92, P3_R1095_U93, P3_R1095_U94, P3_R1095_U95, P3_R1095_U96, P3_R1095_U97, P3_R1095_U98, P3_R1095_U99, P3_R1110_U10, P3_R1110_U100, P3_R1110_U101, P3_R1110_U102, P3_R1110_U103, P3_R1110_U104, P3_R1110_U105, P3_R1110_U106, P3_R1110_U107, P3_R1110_U108, P3_R1110_U109, P3_R1110_U11, P3_R1110_U110, P3_R1110_U111, P3_R1110_U112, P3_R1110_U113, P3_R1110_U114, P3_R1110_U115, P3_R1110_U116, P3_R1110_U117, P3_R1110_U118, P3_R1110_U119, P3_R1110_U12, P3_R1110_U120, P3_R1110_U121, P3_R1110_U122, P3_R1110_U123, P3_R1110_U124, P3_R1110_U125, P3_R1110_U126, P3_R1110_U127, P3_R1110_U128, P3_R1110_U129, P3_R1110_U13, P3_R1110_U130, P3_R1110_U131, P3_R1110_U132, P3_R1110_U133, P3_R1110_U134, P3_R1110_U135, P3_R1110_U136, P3_R1110_U137, P3_R1110_U138, P3_R1110_U139, P3_R1110_U14, P3_R1110_U140, P3_R1110_U141, P3_R1110_U142, P3_R1110_U143, P3_R1110_U144, P3_R1110_U145, P3_R1110_U146, P3_R1110_U147, P3_R1110_U148, P3_R1110_U149, P3_R1110_U15, P3_R1110_U150, P3_R1110_U151, P3_R1110_U152, P3_R1110_U153, P3_R1110_U154, P3_R1110_U155, P3_R1110_U156, P3_R1110_U157, P3_R1110_U158, P3_R1110_U159, P3_R1110_U16, P3_R1110_U160, P3_R1110_U161, P3_R1110_U162, P3_R1110_U163, P3_R1110_U164, P3_R1110_U165, P3_R1110_U166, P3_R1110_U167, P3_R1110_U168, P3_R1110_U169, P3_R1110_U17, P3_R1110_U170, P3_R1110_U171, P3_R1110_U172, P3_R1110_U173, P3_R1110_U174, P3_R1110_U175, P3_R1110_U176, P3_R1110_U177, P3_R1110_U178, P3_R1110_U179, P3_R1110_U18, P3_R1110_U180, P3_R1110_U181, P3_R1110_U182, P3_R1110_U183, P3_R1110_U184, P3_R1110_U185, P3_R1110_U186, P3_R1110_U187, P3_R1110_U188, P3_R1110_U189, P3_R1110_U19, P3_R1110_U190, P3_R1110_U191, P3_R1110_U192, P3_R1110_U193, P3_R1110_U194, P3_R1110_U195, P3_R1110_U196, P3_R1110_U197, P3_R1110_U198, P3_R1110_U199, P3_R1110_U20, P3_R1110_U200, P3_R1110_U201, P3_R1110_U202, P3_R1110_U203, P3_R1110_U204, P3_R1110_U205, P3_R1110_U206, P3_R1110_U207, P3_R1110_U208, P3_R1110_U209, P3_R1110_U21, P3_R1110_U210, P3_R1110_U211, P3_R1110_U212, P3_R1110_U213, P3_R1110_U214, P3_R1110_U215, P3_R1110_U216, P3_R1110_U217, P3_R1110_U218, P3_R1110_U219, P3_R1110_U22, P3_R1110_U220, P3_R1110_U221, P3_R1110_U222, P3_R1110_U223, P3_R1110_U224, P3_R1110_U225, P3_R1110_U226, P3_R1110_U227, P3_R1110_U228, P3_R1110_U229, P3_R1110_U23, P3_R1110_U230, P3_R1110_U231, P3_R1110_U232, P3_R1110_U233, P3_R1110_U234, P3_R1110_U235, P3_R1110_U236, P3_R1110_U237, P3_R1110_U238, P3_R1110_U239, P3_R1110_U24, P3_R1110_U240, P3_R1110_U241, P3_R1110_U242, P3_R1110_U243, P3_R1110_U244, P3_R1110_U245, P3_R1110_U246, P3_R1110_U247, P3_R1110_U248, P3_R1110_U249, P3_R1110_U25, P3_R1110_U250, P3_R1110_U251, P3_R1110_U252, P3_R1110_U253, P3_R1110_U254, P3_R1110_U255, P3_R1110_U256, P3_R1110_U257, P3_R1110_U258, P3_R1110_U259, P3_R1110_U26, P3_R1110_U260, P3_R1110_U261, P3_R1110_U262, P3_R1110_U263, P3_R1110_U264, P3_R1110_U265, P3_R1110_U266, P3_R1110_U267, P3_R1110_U268, P3_R1110_U269, P3_R1110_U27, P3_R1110_U270, P3_R1110_U271, P3_R1110_U272, P3_R1110_U273, P3_R1110_U274, P3_R1110_U275, P3_R1110_U276, P3_R1110_U277, P3_R1110_U278, P3_R1110_U279, P3_R1110_U28, P3_R1110_U280, P3_R1110_U281, P3_R1110_U282, P3_R1110_U283, P3_R1110_U284, P3_R1110_U285, P3_R1110_U286, P3_R1110_U287, P3_R1110_U288, P3_R1110_U289, P3_R1110_U29, P3_R1110_U290, P3_R1110_U291, P3_R1110_U292, P3_R1110_U293, P3_R1110_U294, P3_R1110_U295, P3_R1110_U296, P3_R1110_U297, P3_R1110_U298, P3_R1110_U299, P3_R1110_U30, P3_R1110_U300, P3_R1110_U301, P3_R1110_U302, P3_R1110_U303, P3_R1110_U304, P3_R1110_U305, P3_R1110_U306, P3_R1110_U307, P3_R1110_U308, P3_R1110_U309, P3_R1110_U31, P3_R1110_U310, P3_R1110_U311, P3_R1110_U312, P3_R1110_U313, P3_R1110_U314, P3_R1110_U315, P3_R1110_U316, P3_R1110_U317, P3_R1110_U318, P3_R1110_U319, P3_R1110_U32, P3_R1110_U320, P3_R1110_U321, P3_R1110_U322, P3_R1110_U323, P3_R1110_U324, P3_R1110_U325, P3_R1110_U326, P3_R1110_U327, P3_R1110_U328, P3_R1110_U329, P3_R1110_U33, P3_R1110_U330, P3_R1110_U331, P3_R1110_U332, P3_R1110_U333, P3_R1110_U334, P3_R1110_U335, P3_R1110_U336, P3_R1110_U337, P3_R1110_U338, P3_R1110_U339, P3_R1110_U34, P3_R1110_U340, P3_R1110_U341, P3_R1110_U342, P3_R1110_U343, P3_R1110_U344, P3_R1110_U345, P3_R1110_U346, P3_R1110_U347, P3_R1110_U348, P3_R1110_U349, P3_R1110_U35, P3_R1110_U350, P3_R1110_U351, P3_R1110_U352, P3_R1110_U353, P3_R1110_U354, P3_R1110_U355, P3_R1110_U356, P3_R1110_U357, P3_R1110_U358, P3_R1110_U359, P3_R1110_U36, P3_R1110_U360, P3_R1110_U361, P3_R1110_U362, P3_R1110_U363, P3_R1110_U364, P3_R1110_U365, P3_R1110_U366, P3_R1110_U367, P3_R1110_U368, P3_R1110_U369, P3_R1110_U37, P3_R1110_U370, P3_R1110_U371, P3_R1110_U372, P3_R1110_U373, P3_R1110_U374, P3_R1110_U375, P3_R1110_U376, P3_R1110_U377, P3_R1110_U378, P3_R1110_U379, P3_R1110_U38, P3_R1110_U380, P3_R1110_U381, P3_R1110_U382, P3_R1110_U383, P3_R1110_U384, P3_R1110_U385, P3_R1110_U386, P3_R1110_U387, P3_R1110_U388, P3_R1110_U389, P3_R1110_U39, P3_R1110_U390, P3_R1110_U391, P3_R1110_U392, P3_R1110_U393, P3_R1110_U394, P3_R1110_U395, P3_R1110_U396, P3_R1110_U397, P3_R1110_U398, P3_R1110_U399, P3_R1110_U4, P3_R1110_U40, P3_R1110_U400, P3_R1110_U401, P3_R1110_U402, P3_R1110_U403, P3_R1110_U404, P3_R1110_U405, P3_R1110_U406, P3_R1110_U407, P3_R1110_U408, P3_R1110_U409, P3_R1110_U41, P3_R1110_U410, P3_R1110_U411, P3_R1110_U412, P3_R1110_U413, P3_R1110_U414, P3_R1110_U415, P3_R1110_U416, P3_R1110_U417, P3_R1110_U418, P3_R1110_U419, P3_R1110_U42, P3_R1110_U420, P3_R1110_U421, P3_R1110_U422, P3_R1110_U423, P3_R1110_U424, P3_R1110_U425, P3_R1110_U426, P3_R1110_U427, P3_R1110_U428, P3_R1110_U429, P3_R1110_U43, P3_R1110_U430, P3_R1110_U431, P3_R1110_U432, P3_R1110_U433, P3_R1110_U434, P3_R1110_U435, P3_R1110_U436, P3_R1110_U437, P3_R1110_U438, P3_R1110_U439, P3_R1110_U44, P3_R1110_U440, P3_R1110_U441, P3_R1110_U442, P3_R1110_U443, P3_R1110_U444, P3_R1110_U445, P3_R1110_U446, P3_R1110_U447, P3_R1110_U448, P3_R1110_U449, P3_R1110_U45, P3_R1110_U450, P3_R1110_U451, P3_R1110_U452, P3_R1110_U453, P3_R1110_U454, P3_R1110_U455, P3_R1110_U456, P3_R1110_U457, P3_R1110_U458, P3_R1110_U459, P3_R1110_U46, P3_R1110_U460, P3_R1110_U461, P3_R1110_U462, P3_R1110_U463, P3_R1110_U464, P3_R1110_U465, P3_R1110_U466, P3_R1110_U467, P3_R1110_U468, P3_R1110_U469, P3_R1110_U47, P3_R1110_U470, P3_R1110_U471, P3_R1110_U472, P3_R1110_U473, P3_R1110_U474, P3_R1110_U475, P3_R1110_U476, P3_R1110_U477, P3_R1110_U478, P3_R1110_U479, P3_R1110_U48, P3_R1110_U480, P3_R1110_U481, P3_R1110_U482, P3_R1110_U483, P3_R1110_U484, P3_R1110_U485, P3_R1110_U486, P3_R1110_U487, P3_R1110_U488, P3_R1110_U489, P3_R1110_U49, P3_R1110_U490, P3_R1110_U491, P3_R1110_U492, P3_R1110_U493, P3_R1110_U494, P3_R1110_U495, P3_R1110_U496, P3_R1110_U497, P3_R1110_U498, P3_R1110_U499, P3_R1110_U5, P3_R1110_U50, P3_R1110_U500, P3_R1110_U501, P3_R1110_U502, P3_R1110_U503, P3_R1110_U504, P3_R1110_U51, P3_R1110_U52, P3_R1110_U53, P3_R1110_U54, P3_R1110_U55, P3_R1110_U56, P3_R1110_U57, P3_R1110_U58, P3_R1110_U59, P3_R1110_U6, P3_R1110_U60, P3_R1110_U61, P3_R1110_U62, P3_R1110_U63, P3_R1110_U64, P3_R1110_U65, P3_R1110_U66, P3_R1110_U67, P3_R1110_U68, P3_R1110_U69, P3_R1110_U7, P3_R1110_U70, P3_R1110_U71, P3_R1110_U72, P3_R1110_U73, P3_R1110_U74, P3_R1110_U75, P3_R1110_U76, P3_R1110_U77, P3_R1110_U78, P3_R1110_U79, P3_R1110_U8, P3_R1110_U80, P3_R1110_U81, P3_R1110_U82, P3_R1110_U83, P3_R1110_U84, P3_R1110_U85, P3_R1110_U86, P3_R1110_U87, P3_R1110_U88, P3_R1110_U89, P3_R1110_U9, P3_R1110_U90, P3_R1110_U91, P3_R1110_U92, P3_R1110_U93, P3_R1110_U94, P3_R1110_U95, P3_R1110_U96, P3_R1110_U97, P3_R1110_U98, P3_R1110_U99, P3_R1131_U10, P3_R1131_U100, P3_R1131_U101, P3_R1131_U102, P3_R1131_U103, P3_R1131_U104, P3_R1131_U105, P3_R1131_U106, P3_R1131_U107, P3_R1131_U108, P3_R1131_U109, P3_R1131_U11, P3_R1131_U110, P3_R1131_U111, P3_R1131_U112, P3_R1131_U113, P3_R1131_U114, P3_R1131_U115, P3_R1131_U116, P3_R1131_U117, P3_R1131_U118, P3_R1131_U119, P3_R1131_U12, P3_R1131_U120, P3_R1131_U121, P3_R1131_U122, P3_R1131_U123, P3_R1131_U124, P3_R1131_U125, P3_R1131_U126, P3_R1131_U127, P3_R1131_U128, P3_R1131_U129, P3_R1131_U13, P3_R1131_U130, P3_R1131_U131, P3_R1131_U132, P3_R1131_U133, P3_R1131_U134, P3_R1131_U135, P3_R1131_U136, P3_R1131_U137, P3_R1131_U138, P3_R1131_U139, P3_R1131_U14, P3_R1131_U140, P3_R1131_U141, P3_R1131_U142, P3_R1131_U143, P3_R1131_U144, P3_R1131_U145, P3_R1131_U146, P3_R1131_U147, P3_R1131_U148, P3_R1131_U149, P3_R1131_U15, P3_R1131_U150, P3_R1131_U151, P3_R1131_U152, P3_R1131_U153, P3_R1131_U154, P3_R1131_U155, P3_R1131_U156, P3_R1131_U157, P3_R1131_U158, P3_R1131_U159, P3_R1131_U16, P3_R1131_U160, P3_R1131_U161, P3_R1131_U162, P3_R1131_U163, P3_R1131_U164, P3_R1131_U165, P3_R1131_U166, P3_R1131_U167, P3_R1131_U168, P3_R1131_U169, P3_R1131_U17, P3_R1131_U170, P3_R1131_U171, P3_R1131_U172, P3_R1131_U173, P3_R1131_U174, P3_R1131_U175, P3_R1131_U176, P3_R1131_U177, P3_R1131_U178, P3_R1131_U179, P3_R1131_U18, P3_R1131_U180, P3_R1131_U181, P3_R1131_U182, P3_R1131_U183, P3_R1131_U184, P3_R1131_U185, P3_R1131_U186, P3_R1131_U187, P3_R1131_U188, P3_R1131_U189, P3_R1131_U19, P3_R1131_U190, P3_R1131_U191, P3_R1131_U192, P3_R1131_U193, P3_R1131_U194, P3_R1131_U195, P3_R1131_U196, P3_R1131_U197, P3_R1131_U198, P3_R1131_U199, P3_R1131_U20, P3_R1131_U200, P3_R1131_U201, P3_R1131_U202, P3_R1131_U203, P3_R1131_U204, P3_R1131_U205, P3_R1131_U206, P3_R1131_U207, P3_R1131_U208, P3_R1131_U209, P3_R1131_U21, P3_R1131_U210, P3_R1131_U211, P3_R1131_U212, P3_R1131_U213, P3_R1131_U214, P3_R1131_U215, P3_R1131_U216, P3_R1131_U217, P3_R1131_U218, P3_R1131_U219, P3_R1131_U22, P3_R1131_U220, P3_R1131_U221, P3_R1131_U222, P3_R1131_U223, P3_R1131_U224, P3_R1131_U225, P3_R1131_U226, P3_R1131_U227, P3_R1131_U228, P3_R1131_U229, P3_R1131_U23, P3_R1131_U230, P3_R1131_U231, P3_R1131_U232, P3_R1131_U233, P3_R1131_U234, P3_R1131_U235, P3_R1131_U236, P3_R1131_U237, P3_R1131_U238, P3_R1131_U239, P3_R1131_U24, P3_R1131_U240, P3_R1131_U241, P3_R1131_U242, P3_R1131_U243, P3_R1131_U244, P3_R1131_U245, P3_R1131_U246, P3_R1131_U247, P3_R1131_U248, P3_R1131_U249, P3_R1131_U25, P3_R1131_U250, P3_R1131_U251, P3_R1131_U252, P3_R1131_U253, P3_R1131_U254, P3_R1131_U255, P3_R1131_U256, P3_R1131_U257, P3_R1131_U258, P3_R1131_U259, P3_R1131_U26, P3_R1131_U260, P3_R1131_U261, P3_R1131_U262, P3_R1131_U263, P3_R1131_U264, P3_R1131_U265, P3_R1131_U266, P3_R1131_U267, P3_R1131_U268, P3_R1131_U269, P3_R1131_U27, P3_R1131_U270, P3_R1131_U271, P3_R1131_U272, P3_R1131_U273, P3_R1131_U274, P3_R1131_U275, P3_R1131_U276, P3_R1131_U277, P3_R1131_U278, P3_R1131_U279, P3_R1131_U28, P3_R1131_U280, P3_R1131_U281, P3_R1131_U282, P3_R1131_U283, P3_R1131_U284, P3_R1131_U285, P3_R1131_U286, P3_R1131_U287, P3_R1131_U288, P3_R1131_U289, P3_R1131_U29, P3_R1131_U290, P3_R1131_U291, P3_R1131_U292, P3_R1131_U293, P3_R1131_U294, P3_R1131_U295, P3_R1131_U296, P3_R1131_U297, P3_R1131_U298, P3_R1131_U299, P3_R1131_U30, P3_R1131_U300, P3_R1131_U301, P3_R1131_U302, P3_R1131_U303, P3_R1131_U304, P3_R1131_U305, P3_R1131_U306, P3_R1131_U307, P3_R1131_U308, P3_R1131_U309, P3_R1131_U31, P3_R1131_U310, P3_R1131_U311, P3_R1131_U312, P3_R1131_U313, P3_R1131_U314, P3_R1131_U315, P3_R1131_U316, P3_R1131_U317, P3_R1131_U318, P3_R1131_U319, P3_R1131_U32, P3_R1131_U320, P3_R1131_U321, P3_R1131_U322, P3_R1131_U323, P3_R1131_U324, P3_R1131_U325, P3_R1131_U326, P3_R1131_U327, P3_R1131_U328, P3_R1131_U329, P3_R1131_U33, P3_R1131_U330, P3_R1131_U331, P3_R1131_U332, P3_R1131_U333, P3_R1131_U334, P3_R1131_U335, P3_R1131_U336, P3_R1131_U337, P3_R1131_U338, P3_R1131_U339, P3_R1131_U34, P3_R1131_U340, P3_R1131_U341, P3_R1131_U342, P3_R1131_U343, P3_R1131_U344, P3_R1131_U345, P3_R1131_U346, P3_R1131_U347, P3_R1131_U348, P3_R1131_U349, P3_R1131_U35, P3_R1131_U350, P3_R1131_U351, P3_R1131_U352, P3_R1131_U353, P3_R1131_U354, P3_R1131_U355, P3_R1131_U356, P3_R1131_U357, P3_R1131_U358, P3_R1131_U359, P3_R1131_U36, P3_R1131_U360, P3_R1131_U361, P3_R1131_U362, P3_R1131_U363, P3_R1131_U364, P3_R1131_U365, P3_R1131_U366, P3_R1131_U367, P3_R1131_U368, P3_R1131_U369, P3_R1131_U37, P3_R1131_U370, P3_R1131_U371, P3_R1131_U372, P3_R1131_U373, P3_R1131_U374, P3_R1131_U375, P3_R1131_U376, P3_R1131_U377, P3_R1131_U378, P3_R1131_U379, P3_R1131_U38, P3_R1131_U380, P3_R1131_U381, P3_R1131_U382, P3_R1131_U383, P3_R1131_U384, P3_R1131_U385, P3_R1131_U386, P3_R1131_U387, P3_R1131_U388, P3_R1131_U389, P3_R1131_U39, P3_R1131_U390, P3_R1131_U391, P3_R1131_U392, P3_R1131_U393, P3_R1131_U394, P3_R1131_U395, P3_R1131_U396, P3_R1131_U397, P3_R1131_U398, P3_R1131_U399, P3_R1131_U40, P3_R1131_U400, P3_R1131_U401, P3_R1131_U402, P3_R1131_U403, P3_R1131_U404, P3_R1131_U405, P3_R1131_U406, P3_R1131_U407, P3_R1131_U408, P3_R1131_U409, P3_R1131_U41, P3_R1131_U410, P3_R1131_U411, P3_R1131_U412, P3_R1131_U413, P3_R1131_U414, P3_R1131_U415, P3_R1131_U416, P3_R1131_U417, P3_R1131_U418, P3_R1131_U419, P3_R1131_U42, P3_R1131_U420, P3_R1131_U421, P3_R1131_U422, P3_R1131_U423, P3_R1131_U424, P3_R1131_U425, P3_R1131_U426, P3_R1131_U427, P3_R1131_U428, P3_R1131_U429, P3_R1131_U43, P3_R1131_U430, P3_R1131_U431, P3_R1131_U432, P3_R1131_U433, P3_R1131_U434, P3_R1131_U435, P3_R1131_U436, P3_R1131_U437, P3_R1131_U438, P3_R1131_U439, P3_R1131_U44, P3_R1131_U440, P3_R1131_U441, P3_R1131_U442, P3_R1131_U443, P3_R1131_U444, P3_R1131_U445, P3_R1131_U446, P3_R1131_U447, P3_R1131_U448, P3_R1131_U449, P3_R1131_U45, P3_R1131_U450, P3_R1131_U451, P3_R1131_U452, P3_R1131_U453, P3_R1131_U454, P3_R1131_U455, P3_R1131_U456, P3_R1131_U457, P3_R1131_U458, P3_R1131_U459, P3_R1131_U46, P3_R1131_U460, P3_R1131_U461, P3_R1131_U462, P3_R1131_U463, P3_R1131_U464, P3_R1131_U465, P3_R1131_U466, P3_R1131_U467, P3_R1131_U468, P3_R1131_U469, P3_R1131_U47, P3_R1131_U470, P3_R1131_U471, P3_R1131_U472, P3_R1131_U473, P3_R1131_U474, P3_R1131_U475, P3_R1131_U476, P3_R1131_U477, P3_R1131_U478, P3_R1131_U479, P3_R1131_U48, P3_R1131_U480, P3_R1131_U481, P3_R1131_U482, P3_R1131_U483, P3_R1131_U484, P3_R1131_U485, P3_R1131_U49, P3_R1131_U50, P3_R1131_U51, P3_R1131_U52, P3_R1131_U53, P3_R1131_U54, P3_R1131_U55, P3_R1131_U56, P3_R1131_U57, P3_R1131_U58, P3_R1131_U59, P3_R1131_U6, P3_R1131_U60, P3_R1131_U61, P3_R1131_U62, P3_R1131_U63, P3_R1131_U64, P3_R1131_U65, P3_R1131_U66, P3_R1131_U67, P3_R1131_U68, P3_R1131_U69, P3_R1131_U7, P3_R1131_U70, P3_R1131_U71, P3_R1131_U72, P3_R1131_U73, P3_R1131_U74, P3_R1131_U75, P3_R1131_U76, P3_R1131_U77, P3_R1131_U78, P3_R1131_U79, P3_R1131_U8, P3_R1131_U80, P3_R1131_U81, P3_R1131_U82, P3_R1131_U83, P3_R1131_U84, P3_R1131_U85, P3_R1131_U86, P3_R1131_U87, P3_R1131_U88, P3_R1131_U89, P3_R1131_U9, P3_R1131_U90, P3_R1131_U91, P3_R1131_U92, P3_R1131_U93, P3_R1131_U94, P3_R1131_U95, P3_R1131_U96, P3_R1131_U97, P3_R1131_U98, P3_R1131_U99, P3_R1143_U10, P3_R1143_U100, P3_R1143_U101, P3_R1143_U102, P3_R1143_U103, P3_R1143_U104, P3_R1143_U105, P3_R1143_U106, P3_R1143_U107, P3_R1143_U108, P3_R1143_U109, P3_R1143_U11, P3_R1143_U110, P3_R1143_U111, P3_R1143_U112, P3_R1143_U113, P3_R1143_U114, P3_R1143_U115, P3_R1143_U116, P3_R1143_U117, P3_R1143_U118, P3_R1143_U119, P3_R1143_U12, P3_R1143_U120, P3_R1143_U121, P3_R1143_U122, P3_R1143_U123, P3_R1143_U124, P3_R1143_U125, P3_R1143_U126, P3_R1143_U127, P3_R1143_U128, P3_R1143_U129, P3_R1143_U13, P3_R1143_U130, P3_R1143_U131, P3_R1143_U132, P3_R1143_U133, P3_R1143_U134, P3_R1143_U135, P3_R1143_U136, P3_R1143_U137, P3_R1143_U138, P3_R1143_U139, P3_R1143_U14, P3_R1143_U140, P3_R1143_U141, P3_R1143_U142, P3_R1143_U143, P3_R1143_U144, P3_R1143_U145, P3_R1143_U146, P3_R1143_U147, P3_R1143_U148, P3_R1143_U149, P3_R1143_U15, P3_R1143_U150, P3_R1143_U151, P3_R1143_U152, P3_R1143_U153, P3_R1143_U154, P3_R1143_U155, P3_R1143_U156, P3_R1143_U157, P3_R1143_U158, P3_R1143_U159, P3_R1143_U16, P3_R1143_U160, P3_R1143_U161, P3_R1143_U162, P3_R1143_U163, P3_R1143_U164, P3_R1143_U165, P3_R1143_U166, P3_R1143_U167, P3_R1143_U168, P3_R1143_U169, P3_R1143_U17, P3_R1143_U170, P3_R1143_U171, P3_R1143_U172, P3_R1143_U173, P3_R1143_U174, P3_R1143_U175, P3_R1143_U176, P3_R1143_U177, P3_R1143_U178, P3_R1143_U179, P3_R1143_U18, P3_R1143_U180, P3_R1143_U181, P3_R1143_U182, P3_R1143_U183, P3_R1143_U184, P3_R1143_U185, P3_R1143_U186, P3_R1143_U187, P3_R1143_U188, P3_R1143_U189, P3_R1143_U19, P3_R1143_U190, P3_R1143_U191, P3_R1143_U192, P3_R1143_U193, P3_R1143_U194, P3_R1143_U195, P3_R1143_U196, P3_R1143_U197, P3_R1143_U198, P3_R1143_U199, P3_R1143_U20, P3_R1143_U200, P3_R1143_U201, P3_R1143_U202, P3_R1143_U203, P3_R1143_U204, P3_R1143_U205, P3_R1143_U206, P3_R1143_U207, P3_R1143_U208, P3_R1143_U209, P3_R1143_U21, P3_R1143_U210, P3_R1143_U211, P3_R1143_U212, P3_R1143_U213, P3_R1143_U214, P3_R1143_U215, P3_R1143_U216, P3_R1143_U217, P3_R1143_U218, P3_R1143_U219, P3_R1143_U22, P3_R1143_U220, P3_R1143_U221, P3_R1143_U222, P3_R1143_U223, P3_R1143_U224, P3_R1143_U225, P3_R1143_U226, P3_R1143_U227, P3_R1143_U228, P3_R1143_U229, P3_R1143_U23, P3_R1143_U230, P3_R1143_U231, P3_R1143_U232, P3_R1143_U233, P3_R1143_U234, P3_R1143_U235, P3_R1143_U236, P3_R1143_U237, P3_R1143_U238, P3_R1143_U239, P3_R1143_U24, P3_R1143_U240, P3_R1143_U241, P3_R1143_U242, P3_R1143_U243, P3_R1143_U244, P3_R1143_U245, P3_R1143_U246, P3_R1143_U247, P3_R1143_U248, P3_R1143_U249, P3_R1143_U25, P3_R1143_U250, P3_R1143_U251, P3_R1143_U252, P3_R1143_U253, P3_R1143_U254, P3_R1143_U255, P3_R1143_U256, P3_R1143_U257, P3_R1143_U258, P3_R1143_U259, P3_R1143_U26, P3_R1143_U260, P3_R1143_U261, P3_R1143_U262, P3_R1143_U263, P3_R1143_U264, P3_R1143_U265, P3_R1143_U266, P3_R1143_U267, P3_R1143_U268, P3_R1143_U269, P3_R1143_U27, P3_R1143_U270, P3_R1143_U271, P3_R1143_U272, P3_R1143_U273, P3_R1143_U274, P3_R1143_U275, P3_R1143_U276, P3_R1143_U277, P3_R1143_U278, P3_R1143_U279, P3_R1143_U28, P3_R1143_U280, P3_R1143_U281, P3_R1143_U282, P3_R1143_U283, P3_R1143_U284, P3_R1143_U285, P3_R1143_U286, P3_R1143_U287, P3_R1143_U288, P3_R1143_U289, P3_R1143_U29, P3_R1143_U290, P3_R1143_U291, P3_R1143_U292, P3_R1143_U293, P3_R1143_U294, P3_R1143_U295, P3_R1143_U296, P3_R1143_U297, P3_R1143_U298, P3_R1143_U299, P3_R1143_U30, P3_R1143_U300, P3_R1143_U301, P3_R1143_U302, P3_R1143_U303, P3_R1143_U304, P3_R1143_U305, P3_R1143_U306, P3_R1143_U307, P3_R1143_U308, P3_R1143_U309, P3_R1143_U31, P3_R1143_U310, P3_R1143_U311, P3_R1143_U312, P3_R1143_U313, P3_R1143_U314, P3_R1143_U315, P3_R1143_U316, P3_R1143_U317, P3_R1143_U318, P3_R1143_U319, P3_R1143_U32, P3_R1143_U320, P3_R1143_U321, P3_R1143_U322, P3_R1143_U323, P3_R1143_U324, P3_R1143_U325, P3_R1143_U326, P3_R1143_U327, P3_R1143_U328, P3_R1143_U329, P3_R1143_U33, P3_R1143_U330, P3_R1143_U331, P3_R1143_U332, P3_R1143_U333, P3_R1143_U334, P3_R1143_U335, P3_R1143_U336, P3_R1143_U337, P3_R1143_U338, P3_R1143_U339, P3_R1143_U34, P3_R1143_U340, P3_R1143_U341, P3_R1143_U342, P3_R1143_U343, P3_R1143_U344, P3_R1143_U345, P3_R1143_U346, P3_R1143_U347, P3_R1143_U348, P3_R1143_U349, P3_R1143_U35, P3_R1143_U350, P3_R1143_U351, P3_R1143_U352, P3_R1143_U353, P3_R1143_U354, P3_R1143_U355, P3_R1143_U356, P3_R1143_U357, P3_R1143_U358, P3_R1143_U359, P3_R1143_U36, P3_R1143_U360, P3_R1143_U361, P3_R1143_U362, P3_R1143_U363, P3_R1143_U364, P3_R1143_U365, P3_R1143_U366, P3_R1143_U367, P3_R1143_U368, P3_R1143_U369, P3_R1143_U37, P3_R1143_U370, P3_R1143_U371, P3_R1143_U372, P3_R1143_U373, P3_R1143_U374, P3_R1143_U375, P3_R1143_U376, P3_R1143_U377, P3_R1143_U378, P3_R1143_U379, P3_R1143_U38, P3_R1143_U380, P3_R1143_U381, P3_R1143_U382, P3_R1143_U383, P3_R1143_U384, P3_R1143_U385, P3_R1143_U386, P3_R1143_U387, P3_R1143_U388, P3_R1143_U389, P3_R1143_U39, P3_R1143_U390, P3_R1143_U391, P3_R1143_U392, P3_R1143_U393, P3_R1143_U394, P3_R1143_U395, P3_R1143_U396, P3_R1143_U397, P3_R1143_U398, P3_R1143_U399, P3_R1143_U4, P3_R1143_U40, P3_R1143_U400, P3_R1143_U401, P3_R1143_U402, P3_R1143_U403, P3_R1143_U404, P3_R1143_U405, P3_R1143_U406, P3_R1143_U407, P3_R1143_U408, P3_R1143_U409, P3_R1143_U41, P3_R1143_U410, P3_R1143_U411, P3_R1143_U412, P3_R1143_U413, P3_R1143_U414, P3_R1143_U415, P3_R1143_U416, P3_R1143_U417, P3_R1143_U418, P3_R1143_U419, P3_R1143_U42, P3_R1143_U420, P3_R1143_U421, P3_R1143_U422, P3_R1143_U423, P3_R1143_U424, P3_R1143_U425, P3_R1143_U426, P3_R1143_U427, P3_R1143_U428, P3_R1143_U429, P3_R1143_U43, P3_R1143_U430, P3_R1143_U431, P3_R1143_U432, P3_R1143_U433, P3_R1143_U434, P3_R1143_U435, P3_R1143_U436, P3_R1143_U437, P3_R1143_U438, P3_R1143_U439, P3_R1143_U44, P3_R1143_U440, P3_R1143_U441, P3_R1143_U442, P3_R1143_U443, P3_R1143_U444, P3_R1143_U445, P3_R1143_U446, P3_R1143_U447, P3_R1143_U448, P3_R1143_U449, P3_R1143_U45, P3_R1143_U450, P3_R1143_U451, P3_R1143_U452, P3_R1143_U453, P3_R1143_U454, P3_R1143_U455, P3_R1143_U456, P3_R1143_U457, P3_R1143_U458, P3_R1143_U459, P3_R1143_U46, P3_R1143_U460, P3_R1143_U461, P3_R1143_U462, P3_R1143_U463, P3_R1143_U464, P3_R1143_U465, P3_R1143_U466, P3_R1143_U467, P3_R1143_U468, P3_R1143_U469, P3_R1143_U47, P3_R1143_U470, P3_R1143_U471, P3_R1143_U472, P3_R1143_U473, P3_R1143_U474, P3_R1143_U475, P3_R1143_U476, P3_R1143_U477, P3_R1143_U478, P3_R1143_U479, P3_R1143_U48, P3_R1143_U480, P3_R1143_U481, P3_R1143_U482, P3_R1143_U483, P3_R1143_U484, P3_R1143_U485, P3_R1143_U486, P3_R1143_U487, P3_R1143_U488, P3_R1143_U489, P3_R1143_U49, P3_R1143_U490, P3_R1143_U491, P3_R1143_U492, P3_R1143_U493, P3_R1143_U494, P3_R1143_U495, P3_R1143_U496, P3_R1143_U497, P3_R1143_U498, P3_R1143_U499, P3_R1143_U5, P3_R1143_U50, P3_R1143_U500, P3_R1143_U501, P3_R1143_U502, P3_R1143_U503, P3_R1143_U504, P3_R1143_U51, P3_R1143_U52, P3_R1143_U53, P3_R1143_U54, P3_R1143_U55, P3_R1143_U56, P3_R1143_U57, P3_R1143_U58, P3_R1143_U59, P3_R1143_U6, P3_R1143_U60, P3_R1143_U61, P3_R1143_U62, P3_R1143_U63, P3_R1143_U64, P3_R1143_U65, P3_R1143_U66, P3_R1143_U67, P3_R1143_U68, P3_R1143_U69, P3_R1143_U7, P3_R1143_U70, P3_R1143_U71, P3_R1143_U72, P3_R1143_U73, P3_R1143_U74, P3_R1143_U75, P3_R1143_U76, P3_R1143_U77, P3_R1143_U78, P3_R1143_U79, P3_R1143_U8, P3_R1143_U80, P3_R1143_U81, P3_R1143_U82, P3_R1143_U83, P3_R1143_U84, P3_R1143_U85, P3_R1143_U86, P3_R1143_U87, P3_R1143_U88, P3_R1143_U89, P3_R1143_U9, P3_R1143_U90, P3_R1143_U91, P3_R1143_U92, P3_R1143_U93, P3_R1143_U94, P3_R1143_U95, P3_R1143_U96, P3_R1143_U97, P3_R1143_U98, P3_R1143_U99, P3_R1158_U10, P3_R1158_U100, P3_R1158_U101, P3_R1158_U102, P3_R1158_U103, P3_R1158_U104, P3_R1158_U105, P3_R1158_U106, P3_R1158_U107, P3_R1158_U108, P3_R1158_U109, P3_R1158_U11, P3_R1158_U110, P3_R1158_U111, P3_R1158_U112, P3_R1158_U113, P3_R1158_U114, P3_R1158_U115, P3_R1158_U116, P3_R1158_U117, P3_R1158_U118, P3_R1158_U119, P3_R1158_U12, P3_R1158_U120, P3_R1158_U121, P3_R1158_U122, P3_R1158_U123, P3_R1158_U124, P3_R1158_U125, P3_R1158_U126, P3_R1158_U127, P3_R1158_U128, P3_R1158_U129, P3_R1158_U13, P3_R1158_U130, P3_R1158_U131, P3_R1158_U132, P3_R1158_U133, P3_R1158_U134, P3_R1158_U135, P3_R1158_U136, P3_R1158_U137, P3_R1158_U138, P3_R1158_U139, P3_R1158_U14, P3_R1158_U140, P3_R1158_U141, P3_R1158_U142, P3_R1158_U143, P3_R1158_U144, P3_R1158_U145, P3_R1158_U146, P3_R1158_U147, P3_R1158_U148, P3_R1158_U149, P3_R1158_U15, P3_R1158_U150, P3_R1158_U151, P3_R1158_U152, P3_R1158_U153, P3_R1158_U154, P3_R1158_U155, P3_R1158_U156, P3_R1158_U157, P3_R1158_U158, P3_R1158_U159, P3_R1158_U16, P3_R1158_U160, P3_R1158_U161, P3_R1158_U162, P3_R1158_U163, P3_R1158_U164, P3_R1158_U165, P3_R1158_U166, P3_R1158_U167, P3_R1158_U168, P3_R1158_U169, P3_R1158_U17, P3_R1158_U170, P3_R1158_U171, P3_R1158_U172, P3_R1158_U173, P3_R1158_U174, P3_R1158_U175, P3_R1158_U176, P3_R1158_U177, P3_R1158_U178, P3_R1158_U179, P3_R1158_U18, P3_R1158_U180, P3_R1158_U181, P3_R1158_U182, P3_R1158_U183, P3_R1158_U184, P3_R1158_U185, P3_R1158_U186, P3_R1158_U187, P3_R1158_U188, P3_R1158_U189, P3_R1158_U19, P3_R1158_U190, P3_R1158_U191, P3_R1158_U192, P3_R1158_U193, P3_R1158_U194, P3_R1158_U195, P3_R1158_U196, P3_R1158_U197, P3_R1158_U198, P3_R1158_U199, P3_R1158_U20, P3_R1158_U200, P3_R1158_U201, P3_R1158_U202, P3_R1158_U203, P3_R1158_U204, P3_R1158_U205, P3_R1158_U206, P3_R1158_U207, P3_R1158_U208, P3_R1158_U209, P3_R1158_U21, P3_R1158_U210, P3_R1158_U211, P3_R1158_U212, P3_R1158_U213, P3_R1158_U214, P3_R1158_U215, P3_R1158_U216, P3_R1158_U217, P3_R1158_U218, P3_R1158_U219, P3_R1158_U22, P3_R1158_U220, P3_R1158_U221, P3_R1158_U222, P3_R1158_U223, P3_R1158_U224, P3_R1158_U225, P3_R1158_U226, P3_R1158_U227, P3_R1158_U228, P3_R1158_U229, P3_R1158_U23, P3_R1158_U230, P3_R1158_U231, P3_R1158_U232, P3_R1158_U233, P3_R1158_U234, P3_R1158_U235, P3_R1158_U236, P3_R1158_U237, P3_R1158_U238, P3_R1158_U239, P3_R1158_U24, P3_R1158_U240, P3_R1158_U241, P3_R1158_U242, P3_R1158_U243, P3_R1158_U244, P3_R1158_U245, P3_R1158_U246, P3_R1158_U247, P3_R1158_U248, P3_R1158_U249, P3_R1158_U25, P3_R1158_U250, P3_R1158_U251, P3_R1158_U252, P3_R1158_U253, P3_R1158_U254, P3_R1158_U255, P3_R1158_U256, P3_R1158_U257, P3_R1158_U258, P3_R1158_U259, P3_R1158_U26, P3_R1158_U260, P3_R1158_U261, P3_R1158_U262, P3_R1158_U263, P3_R1158_U264, P3_R1158_U265, P3_R1158_U266, P3_R1158_U267, P3_R1158_U268, P3_R1158_U269, P3_R1158_U27, P3_R1158_U270, P3_R1158_U271, P3_R1158_U272, P3_R1158_U273, P3_R1158_U274, P3_R1158_U275, P3_R1158_U276, P3_R1158_U277, P3_R1158_U278, P3_R1158_U279, P3_R1158_U28, P3_R1158_U280, P3_R1158_U281, P3_R1158_U282, P3_R1158_U283, P3_R1158_U284, P3_R1158_U285, P3_R1158_U286, P3_R1158_U287, P3_R1158_U288, P3_R1158_U289, P3_R1158_U29, P3_R1158_U290, P3_R1158_U291, P3_R1158_U292, P3_R1158_U293, P3_R1158_U294, P3_R1158_U295, P3_R1158_U296, P3_R1158_U297, P3_R1158_U298, P3_R1158_U299, P3_R1158_U30, P3_R1158_U300, P3_R1158_U301, P3_R1158_U302, P3_R1158_U303, P3_R1158_U304, P3_R1158_U305, P3_R1158_U306, P3_R1158_U307, P3_R1158_U308, P3_R1158_U309, P3_R1158_U31, P3_R1158_U310, P3_R1158_U311, P3_R1158_U312, P3_R1158_U313, P3_R1158_U314, P3_R1158_U315, P3_R1158_U316, P3_R1158_U317, P3_R1158_U318, P3_R1158_U319, P3_R1158_U32, P3_R1158_U320, P3_R1158_U321, P3_R1158_U322, P3_R1158_U323, P3_R1158_U324, P3_R1158_U325, P3_R1158_U326, P3_R1158_U327, P3_R1158_U328, P3_R1158_U329, P3_R1158_U33, P3_R1158_U330, P3_R1158_U331, P3_R1158_U332, P3_R1158_U333, P3_R1158_U334, P3_R1158_U335, P3_R1158_U336, P3_R1158_U337, P3_R1158_U338, P3_R1158_U339, P3_R1158_U34, P3_R1158_U340, P3_R1158_U341, P3_R1158_U342, P3_R1158_U343, P3_R1158_U344, P3_R1158_U345, P3_R1158_U346, P3_R1158_U347, P3_R1158_U348, P3_R1158_U349, P3_R1158_U35, P3_R1158_U350, P3_R1158_U351, P3_R1158_U352, P3_R1158_U353, P3_R1158_U354, P3_R1158_U355, P3_R1158_U356, P3_R1158_U357, P3_R1158_U358, P3_R1158_U359, P3_R1158_U36, P3_R1158_U360, P3_R1158_U361, P3_R1158_U362, P3_R1158_U363, P3_R1158_U364, P3_R1158_U365, P3_R1158_U366, P3_R1158_U367, P3_R1158_U368, P3_R1158_U369, P3_R1158_U37, P3_R1158_U370, P3_R1158_U371, P3_R1158_U372, P3_R1158_U373, P3_R1158_U374, P3_R1158_U375, P3_R1158_U376, P3_R1158_U377, P3_R1158_U378, P3_R1158_U379, P3_R1158_U38, P3_R1158_U380, P3_R1158_U381, P3_R1158_U382, P3_R1158_U383, P3_R1158_U384, P3_R1158_U385, P3_R1158_U386, P3_R1158_U387, P3_R1158_U388, P3_R1158_U389, P3_R1158_U39, P3_R1158_U390, P3_R1158_U391, P3_R1158_U392, P3_R1158_U393, P3_R1158_U394, P3_R1158_U395, P3_R1158_U396, P3_R1158_U397, P3_R1158_U398, P3_R1158_U399, P3_R1158_U4, P3_R1158_U40, P3_R1158_U400, P3_R1158_U401, P3_R1158_U402, P3_R1158_U403, P3_R1158_U404, P3_R1158_U405, P3_R1158_U406, P3_R1158_U407, P3_R1158_U408, P3_R1158_U409, P3_R1158_U41, P3_R1158_U410, P3_R1158_U411, P3_R1158_U412, P3_R1158_U413, P3_R1158_U414, P3_R1158_U415, P3_R1158_U416, P3_R1158_U417, P3_R1158_U418, P3_R1158_U419, P3_R1158_U42, P3_R1158_U420, P3_R1158_U421, P3_R1158_U422, P3_R1158_U423, P3_R1158_U424, P3_R1158_U425, P3_R1158_U426, P3_R1158_U427, P3_R1158_U428, P3_R1158_U429, P3_R1158_U43, P3_R1158_U430, P3_R1158_U431, P3_R1158_U432, P3_R1158_U433, P3_R1158_U434, P3_R1158_U435, P3_R1158_U436, P3_R1158_U437, P3_R1158_U438, P3_R1158_U439, P3_R1158_U44, P3_R1158_U440, P3_R1158_U441, P3_R1158_U442, P3_R1158_U443, P3_R1158_U444, P3_R1158_U445, P3_R1158_U446, P3_R1158_U447, P3_R1158_U448, P3_R1158_U449, P3_R1158_U45, P3_R1158_U450, P3_R1158_U451, P3_R1158_U452, P3_R1158_U453, P3_R1158_U454, P3_R1158_U455, P3_R1158_U456, P3_R1158_U457, P3_R1158_U458, P3_R1158_U459, P3_R1158_U46, P3_R1158_U460, P3_R1158_U461, P3_R1158_U462, P3_R1158_U463, P3_R1158_U464, P3_R1158_U465, P3_R1158_U466, P3_R1158_U467, P3_R1158_U468, P3_R1158_U469, P3_R1158_U47, P3_R1158_U470, P3_R1158_U471, P3_R1158_U472, P3_R1158_U473, P3_R1158_U474, P3_R1158_U475, P3_R1158_U476, P3_R1158_U477, P3_R1158_U478, P3_R1158_U479, P3_R1158_U48, P3_R1158_U480, P3_R1158_U481, P3_R1158_U482, P3_R1158_U483, P3_R1158_U484, P3_R1158_U485, P3_R1158_U486, P3_R1158_U487, P3_R1158_U488, P3_R1158_U489, P3_R1158_U49, P3_R1158_U490, P3_R1158_U491, P3_R1158_U492, P3_R1158_U493, P3_R1158_U494, P3_R1158_U495, P3_R1158_U496, P3_R1158_U497, P3_R1158_U498, P3_R1158_U499, P3_R1158_U5, P3_R1158_U50, P3_R1158_U500, P3_R1158_U501, P3_R1158_U502, P3_R1158_U503, P3_R1158_U504, P3_R1158_U505, P3_R1158_U506, P3_R1158_U507, P3_R1158_U508, P3_R1158_U509, P3_R1158_U51, P3_R1158_U510, P3_R1158_U511, P3_R1158_U512, P3_R1158_U513, P3_R1158_U514, P3_R1158_U515, P3_R1158_U516, P3_R1158_U517, P3_R1158_U518, P3_R1158_U519, P3_R1158_U52, P3_R1158_U520, P3_R1158_U521, P3_R1158_U522, P3_R1158_U523, P3_R1158_U524, P3_R1158_U525, P3_R1158_U526, P3_R1158_U527, P3_R1158_U528, P3_R1158_U529, P3_R1158_U53, P3_R1158_U530, P3_R1158_U531, P3_R1158_U532, P3_R1158_U533, P3_R1158_U534, P3_R1158_U535, P3_R1158_U536, P3_R1158_U537, P3_R1158_U538, P3_R1158_U539, P3_R1158_U54, P3_R1158_U540, P3_R1158_U541, P3_R1158_U542, P3_R1158_U543, P3_R1158_U544, P3_R1158_U545, P3_R1158_U546, P3_R1158_U547, P3_R1158_U548, P3_R1158_U549, P3_R1158_U55, P3_R1158_U550, P3_R1158_U551, P3_R1158_U552, P3_R1158_U553, P3_R1158_U554, P3_R1158_U555, P3_R1158_U556, P3_R1158_U557, P3_R1158_U558, P3_R1158_U559, P3_R1158_U56, P3_R1158_U560, P3_R1158_U561, P3_R1158_U562, P3_R1158_U563, P3_R1158_U564, P3_R1158_U565, P3_R1158_U566, P3_R1158_U567, P3_R1158_U568, P3_R1158_U569, P3_R1158_U57, P3_R1158_U570, P3_R1158_U571, P3_R1158_U572, P3_R1158_U573, P3_R1158_U574, P3_R1158_U575, P3_R1158_U576, P3_R1158_U577, P3_R1158_U578, P3_R1158_U579, P3_R1158_U58, P3_R1158_U580, P3_R1158_U581, P3_R1158_U582, P3_R1158_U583, P3_R1158_U584, P3_R1158_U585, P3_R1158_U586, P3_R1158_U587, P3_R1158_U588, P3_R1158_U589, P3_R1158_U59, P3_R1158_U590, P3_R1158_U591, P3_R1158_U592, P3_R1158_U593, P3_R1158_U594, P3_R1158_U595, P3_R1158_U596, P3_R1158_U597, P3_R1158_U598, P3_R1158_U599, P3_R1158_U6, P3_R1158_U60, P3_R1158_U600, P3_R1158_U601, P3_R1158_U602, P3_R1158_U603, P3_R1158_U604, P3_R1158_U605, P3_R1158_U606, P3_R1158_U607, P3_R1158_U608, P3_R1158_U609, P3_R1158_U61, P3_R1158_U610, P3_R1158_U611, P3_R1158_U612, P3_R1158_U613, P3_R1158_U614, P3_R1158_U615, P3_R1158_U616, P3_R1158_U617, P3_R1158_U618, P3_R1158_U619, P3_R1158_U62, P3_R1158_U620, P3_R1158_U621, P3_R1158_U622, P3_R1158_U623, P3_R1158_U624, P3_R1158_U625, P3_R1158_U626, P3_R1158_U627, P3_R1158_U628, P3_R1158_U629, P3_R1158_U63, P3_R1158_U630, P3_R1158_U631, P3_R1158_U632, P3_R1158_U64, P3_R1158_U65, P3_R1158_U66, P3_R1158_U67, P3_R1158_U68, P3_R1158_U69, P3_R1158_U7, P3_R1158_U70, P3_R1158_U71, P3_R1158_U72, P3_R1158_U73, P3_R1158_U74, P3_R1158_U75, P3_R1158_U76, P3_R1158_U77, P3_R1158_U78, P3_R1158_U79, P3_R1158_U8, P3_R1158_U80, P3_R1158_U81, P3_R1158_U82, P3_R1158_U83, P3_R1158_U84, P3_R1158_U85, P3_R1158_U86, P3_R1158_U87, P3_R1158_U88, P3_R1158_U89, P3_R1158_U9, P3_R1158_U90, P3_R1158_U91, P3_R1158_U92, P3_R1158_U93, P3_R1158_U94, P3_R1158_U95, P3_R1158_U96, P3_R1158_U97, P3_R1158_U98, P3_R1158_U99, P3_R1161_U10, P3_R1161_U100, P3_R1161_U101, P3_R1161_U102, P3_R1161_U103, P3_R1161_U104, P3_R1161_U105, P3_R1161_U106, P3_R1161_U107, P3_R1161_U108, P3_R1161_U109, P3_R1161_U11, P3_R1161_U110, P3_R1161_U111, P3_R1161_U112, P3_R1161_U113, P3_R1161_U114, P3_R1161_U115, P3_R1161_U116, P3_R1161_U117, P3_R1161_U118, P3_R1161_U119, P3_R1161_U12, P3_R1161_U120, P3_R1161_U121, P3_R1161_U122, P3_R1161_U123, P3_R1161_U124, P3_R1161_U125, P3_R1161_U126, P3_R1161_U127, P3_R1161_U128, P3_R1161_U129, P3_R1161_U13, P3_R1161_U130, P3_R1161_U131, P3_R1161_U132, P3_R1161_U133, P3_R1161_U134, P3_R1161_U135, P3_R1161_U136, P3_R1161_U137, P3_R1161_U138, P3_R1161_U139, P3_R1161_U14, P3_R1161_U140, P3_R1161_U141, P3_R1161_U142, P3_R1161_U143, P3_R1161_U144, P3_R1161_U145, P3_R1161_U146, P3_R1161_U147, P3_R1161_U148, P3_R1161_U149, P3_R1161_U15, P3_R1161_U150, P3_R1161_U151, P3_R1161_U152, P3_R1161_U153, P3_R1161_U154, P3_R1161_U155, P3_R1161_U156, P3_R1161_U157, P3_R1161_U158, P3_R1161_U159, P3_R1161_U16, P3_R1161_U160, P3_R1161_U161, P3_R1161_U162, P3_R1161_U163, P3_R1161_U164, P3_R1161_U165, P3_R1161_U166, P3_R1161_U167, P3_R1161_U168, P3_R1161_U169, P3_R1161_U17, P3_R1161_U170, P3_R1161_U171, P3_R1161_U172, P3_R1161_U173, P3_R1161_U174, P3_R1161_U175, P3_R1161_U176, P3_R1161_U177, P3_R1161_U178, P3_R1161_U179, P3_R1161_U18, P3_R1161_U180, P3_R1161_U181, P3_R1161_U182, P3_R1161_U183, P3_R1161_U184, P3_R1161_U185, P3_R1161_U186, P3_R1161_U187, P3_R1161_U188, P3_R1161_U189, P3_R1161_U19, P3_R1161_U190, P3_R1161_U191, P3_R1161_U192, P3_R1161_U193, P3_R1161_U194, P3_R1161_U195, P3_R1161_U196, P3_R1161_U197, P3_R1161_U198, P3_R1161_U199, P3_R1161_U20, P3_R1161_U200, P3_R1161_U201, P3_R1161_U202, P3_R1161_U203, P3_R1161_U204, P3_R1161_U205, P3_R1161_U206, P3_R1161_U207, P3_R1161_U208, P3_R1161_U209, P3_R1161_U21, P3_R1161_U210, P3_R1161_U211, P3_R1161_U212, P3_R1161_U213, P3_R1161_U214, P3_R1161_U215, P3_R1161_U216, P3_R1161_U217, P3_R1161_U218, P3_R1161_U219, P3_R1161_U22, P3_R1161_U220, P3_R1161_U221, P3_R1161_U222, P3_R1161_U223, P3_R1161_U224, P3_R1161_U225, P3_R1161_U226, P3_R1161_U227, P3_R1161_U228, P3_R1161_U229, P3_R1161_U23, P3_R1161_U230, P3_R1161_U231, P3_R1161_U232, P3_R1161_U233, P3_R1161_U234, P3_R1161_U235, P3_R1161_U236, P3_R1161_U237, P3_R1161_U238, P3_R1161_U239, P3_R1161_U24, P3_R1161_U240, P3_R1161_U241, P3_R1161_U242, P3_R1161_U243, P3_R1161_U244, P3_R1161_U245, P3_R1161_U246, P3_R1161_U247, P3_R1161_U248, P3_R1161_U249, P3_R1161_U25, P3_R1161_U250, P3_R1161_U251, P3_R1161_U252, P3_R1161_U253, P3_R1161_U254, P3_R1161_U255, P3_R1161_U256, P3_R1161_U257, P3_R1161_U258, P3_R1161_U259, P3_R1161_U26, P3_R1161_U260, P3_R1161_U261, P3_R1161_U262, P3_R1161_U263, P3_R1161_U264, P3_R1161_U265, P3_R1161_U266, P3_R1161_U267, P3_R1161_U268, P3_R1161_U269, P3_R1161_U27, P3_R1161_U270, P3_R1161_U271, P3_R1161_U272, P3_R1161_U273, P3_R1161_U274, P3_R1161_U275, P3_R1161_U276, P3_R1161_U277, P3_R1161_U278, P3_R1161_U279, P3_R1161_U28, P3_R1161_U280, P3_R1161_U281, P3_R1161_U282, P3_R1161_U283, P3_R1161_U284, P3_R1161_U285, P3_R1161_U286, P3_R1161_U287, P3_R1161_U288, P3_R1161_U289, P3_R1161_U29, P3_R1161_U290, P3_R1161_U291, P3_R1161_U292, P3_R1161_U293, P3_R1161_U294, P3_R1161_U295, P3_R1161_U296, P3_R1161_U297, P3_R1161_U298, P3_R1161_U299, P3_R1161_U30, P3_R1161_U300, P3_R1161_U301, P3_R1161_U302, P3_R1161_U303, P3_R1161_U304, P3_R1161_U305, P3_R1161_U306, P3_R1161_U307, P3_R1161_U308, P3_R1161_U309, P3_R1161_U31, P3_R1161_U310, P3_R1161_U311, P3_R1161_U312, P3_R1161_U313, P3_R1161_U314, P3_R1161_U315, P3_R1161_U316, P3_R1161_U317, P3_R1161_U318, P3_R1161_U319, P3_R1161_U32, P3_R1161_U320, P3_R1161_U321, P3_R1161_U322, P3_R1161_U323, P3_R1161_U324, P3_R1161_U325, P3_R1161_U326, P3_R1161_U327, P3_R1161_U328, P3_R1161_U329, P3_R1161_U33, P3_R1161_U330, P3_R1161_U331, P3_R1161_U332, P3_R1161_U333, P3_R1161_U334, P3_R1161_U335, P3_R1161_U336, P3_R1161_U337, P3_R1161_U338, P3_R1161_U339, P3_R1161_U34, P3_R1161_U340, P3_R1161_U341, P3_R1161_U342, P3_R1161_U343, P3_R1161_U344, P3_R1161_U345, P3_R1161_U346, P3_R1161_U347, P3_R1161_U348, P3_R1161_U349, P3_R1161_U35, P3_R1161_U350, P3_R1161_U351, P3_R1161_U352, P3_R1161_U353, P3_R1161_U354, P3_R1161_U355, P3_R1161_U356, P3_R1161_U357, P3_R1161_U358, P3_R1161_U359, P3_R1161_U36, P3_R1161_U360, P3_R1161_U361, P3_R1161_U362, P3_R1161_U363, P3_R1161_U364, P3_R1161_U365, P3_R1161_U366, P3_R1161_U367, P3_R1161_U368, P3_R1161_U369, P3_R1161_U37, P3_R1161_U370, P3_R1161_U371, P3_R1161_U372, P3_R1161_U373, P3_R1161_U374, P3_R1161_U375, P3_R1161_U376, P3_R1161_U377, P3_R1161_U378, P3_R1161_U379, P3_R1161_U38, P3_R1161_U380, P3_R1161_U381, P3_R1161_U382, P3_R1161_U383, P3_R1161_U384, P3_R1161_U385, P3_R1161_U386, P3_R1161_U387, P3_R1161_U388, P3_R1161_U389, P3_R1161_U39, P3_R1161_U390, P3_R1161_U391, P3_R1161_U392, P3_R1161_U393, P3_R1161_U394, P3_R1161_U395, P3_R1161_U396, P3_R1161_U397, P3_R1161_U398, P3_R1161_U399, P3_R1161_U4, P3_R1161_U40, P3_R1161_U400, P3_R1161_U401, P3_R1161_U402, P3_R1161_U403, P3_R1161_U404, P3_R1161_U405, P3_R1161_U406, P3_R1161_U407, P3_R1161_U408, P3_R1161_U409, P3_R1161_U41, P3_R1161_U410, P3_R1161_U411, P3_R1161_U412, P3_R1161_U413, P3_R1161_U414, P3_R1161_U415, P3_R1161_U416, P3_R1161_U417, P3_R1161_U418, P3_R1161_U419, P3_R1161_U42, P3_R1161_U420, P3_R1161_U421, P3_R1161_U422, P3_R1161_U423, P3_R1161_U424, P3_R1161_U425, P3_R1161_U426, P3_R1161_U427, P3_R1161_U428, P3_R1161_U429, P3_R1161_U43, P3_R1161_U430, P3_R1161_U431, P3_R1161_U432, P3_R1161_U433, P3_R1161_U434, P3_R1161_U435, P3_R1161_U436, P3_R1161_U437, P3_R1161_U438, P3_R1161_U439, P3_R1161_U44, P3_R1161_U440, P3_R1161_U441, P3_R1161_U442, P3_R1161_U443, P3_R1161_U444, P3_R1161_U445, P3_R1161_U446, P3_R1161_U447, P3_R1161_U448, P3_R1161_U449, P3_R1161_U45, P3_R1161_U450, P3_R1161_U451, P3_R1161_U452, P3_R1161_U453, P3_R1161_U454, P3_R1161_U455, P3_R1161_U456, P3_R1161_U457, P3_R1161_U458, P3_R1161_U459, P3_R1161_U46, P3_R1161_U460, P3_R1161_U461, P3_R1161_U462, P3_R1161_U463, P3_R1161_U464, P3_R1161_U465, P3_R1161_U466, P3_R1161_U467, P3_R1161_U468, P3_R1161_U469, P3_R1161_U47, P3_R1161_U470, P3_R1161_U471, P3_R1161_U472, P3_R1161_U473, P3_R1161_U474, P3_R1161_U475, P3_R1161_U476, P3_R1161_U477, P3_R1161_U478, P3_R1161_U479, P3_R1161_U48, P3_R1161_U480, P3_R1161_U481, P3_R1161_U482, P3_R1161_U483, P3_R1161_U484, P3_R1161_U485, P3_R1161_U486, P3_R1161_U487, P3_R1161_U488, P3_R1161_U489, P3_R1161_U49, P3_R1161_U490, P3_R1161_U491, P3_R1161_U492, P3_R1161_U493, P3_R1161_U494, P3_R1161_U495, P3_R1161_U496, P3_R1161_U497, P3_R1161_U498, P3_R1161_U499, P3_R1161_U5, P3_R1161_U50, P3_R1161_U500, P3_R1161_U501, P3_R1161_U502, P3_R1161_U503, P3_R1161_U504, P3_R1161_U51, P3_R1161_U52, P3_R1161_U53, P3_R1161_U54, P3_R1161_U55, P3_R1161_U56, P3_R1161_U57, P3_R1161_U58, P3_R1161_U59, P3_R1161_U6, P3_R1161_U60, P3_R1161_U61, P3_R1161_U62, P3_R1161_U63, P3_R1161_U64, P3_R1161_U65, P3_R1161_U66, P3_R1161_U67, P3_R1161_U68, P3_R1161_U69, P3_R1161_U7, P3_R1161_U70, P3_R1161_U71, P3_R1161_U72, P3_R1161_U73, P3_R1161_U74, P3_R1161_U75, P3_R1161_U76, P3_R1161_U77, P3_R1161_U78, P3_R1161_U79, P3_R1161_U8, P3_R1161_U80, P3_R1161_U81, P3_R1161_U82, P3_R1161_U83, P3_R1161_U84, P3_R1161_U85, P3_R1161_U86, P3_R1161_U87, P3_R1161_U88, P3_R1161_U89, P3_R1161_U9, P3_R1161_U90, P3_R1161_U91, P3_R1161_U92, P3_R1161_U93, P3_R1161_U94, P3_R1161_U95, P3_R1161_U96, P3_R1161_U97, P3_R1161_U98, P3_R1161_U99, P3_R1179_U10, P3_R1179_U100, P3_R1179_U101, P3_R1179_U102, P3_R1179_U103, P3_R1179_U104, P3_R1179_U105, P3_R1179_U106, P3_R1179_U107, P3_R1179_U108, P3_R1179_U109, P3_R1179_U11, P3_R1179_U110, P3_R1179_U111, P3_R1179_U112, P3_R1179_U113, P3_R1179_U114, P3_R1179_U115, P3_R1179_U116, P3_R1179_U117, P3_R1179_U118, P3_R1179_U119, P3_R1179_U12, P3_R1179_U120, P3_R1179_U121, P3_R1179_U122, P3_R1179_U123, P3_R1179_U124, P3_R1179_U125, P3_R1179_U126, P3_R1179_U127, P3_R1179_U128, P3_R1179_U129, P3_R1179_U13, P3_R1179_U130, P3_R1179_U131, P3_R1179_U132, P3_R1179_U133, P3_R1179_U134, P3_R1179_U135, P3_R1179_U136, P3_R1179_U137, P3_R1179_U138, P3_R1179_U139, P3_R1179_U14, P3_R1179_U140, P3_R1179_U141, P3_R1179_U142, P3_R1179_U143, P3_R1179_U144, P3_R1179_U145, P3_R1179_U146, P3_R1179_U147, P3_R1179_U148, P3_R1179_U149, P3_R1179_U15, P3_R1179_U150, P3_R1179_U151, P3_R1179_U152, P3_R1179_U153, P3_R1179_U154, P3_R1179_U155, P3_R1179_U156, P3_R1179_U157, P3_R1179_U158, P3_R1179_U159, P3_R1179_U16, P3_R1179_U160, P3_R1179_U161, P3_R1179_U162, P3_R1179_U163, P3_R1179_U164, P3_R1179_U165, P3_R1179_U166, P3_R1179_U167, P3_R1179_U168, P3_R1179_U169, P3_R1179_U17, P3_R1179_U170, P3_R1179_U171, P3_R1179_U172, P3_R1179_U173, P3_R1179_U174, P3_R1179_U175, P3_R1179_U176, P3_R1179_U177, P3_R1179_U178, P3_R1179_U179, P3_R1179_U18, P3_R1179_U180, P3_R1179_U181, P3_R1179_U182, P3_R1179_U183, P3_R1179_U184, P3_R1179_U185, P3_R1179_U186, P3_R1179_U187, P3_R1179_U188, P3_R1179_U189, P3_R1179_U19, P3_R1179_U190, P3_R1179_U191, P3_R1179_U192, P3_R1179_U193, P3_R1179_U194, P3_R1179_U195, P3_R1179_U196, P3_R1179_U197, P3_R1179_U198, P3_R1179_U199, P3_R1179_U20, P3_R1179_U200, P3_R1179_U201, P3_R1179_U202, P3_R1179_U203, P3_R1179_U204, P3_R1179_U205, P3_R1179_U206, P3_R1179_U207, P3_R1179_U208, P3_R1179_U209, P3_R1179_U21, P3_R1179_U210, P3_R1179_U211, P3_R1179_U212, P3_R1179_U213, P3_R1179_U214, P3_R1179_U215, P3_R1179_U216, P3_R1179_U217, P3_R1179_U218, P3_R1179_U219, P3_R1179_U22, P3_R1179_U220, P3_R1179_U221, P3_R1179_U222, P3_R1179_U223, P3_R1179_U224, P3_R1179_U225, P3_R1179_U226, P3_R1179_U227, P3_R1179_U228, P3_R1179_U229, P3_R1179_U23, P3_R1179_U230, P3_R1179_U231, P3_R1179_U232, P3_R1179_U233, P3_R1179_U234, P3_R1179_U235, P3_R1179_U236, P3_R1179_U237, P3_R1179_U238, P3_R1179_U239, P3_R1179_U24, P3_R1179_U240, P3_R1179_U241, P3_R1179_U242, P3_R1179_U243, P3_R1179_U244, P3_R1179_U245, P3_R1179_U246, P3_R1179_U247, P3_R1179_U248, P3_R1179_U249, P3_R1179_U25, P3_R1179_U250, P3_R1179_U251, P3_R1179_U252, P3_R1179_U253, P3_R1179_U254, P3_R1179_U255, P3_R1179_U256, P3_R1179_U257, P3_R1179_U258, P3_R1179_U259, P3_R1179_U26, P3_R1179_U260, P3_R1179_U261, P3_R1179_U262, P3_R1179_U263, P3_R1179_U264, P3_R1179_U265, P3_R1179_U266, P3_R1179_U267, P3_R1179_U268, P3_R1179_U269, P3_R1179_U27, P3_R1179_U270, P3_R1179_U271, P3_R1179_U272, P3_R1179_U273, P3_R1179_U274, P3_R1179_U275, P3_R1179_U276, P3_R1179_U277, P3_R1179_U278, P3_R1179_U279, P3_R1179_U28, P3_R1179_U280, P3_R1179_U281, P3_R1179_U282, P3_R1179_U283, P3_R1179_U284, P3_R1179_U285, P3_R1179_U286, P3_R1179_U287, P3_R1179_U288, P3_R1179_U289, P3_R1179_U29, P3_R1179_U290, P3_R1179_U291, P3_R1179_U292, P3_R1179_U293, P3_R1179_U294, P3_R1179_U295, P3_R1179_U296, P3_R1179_U297, P3_R1179_U298, P3_R1179_U299, P3_R1179_U30, P3_R1179_U300, P3_R1179_U301, P3_R1179_U302, P3_R1179_U303, P3_R1179_U304, P3_R1179_U305, P3_R1179_U306, P3_R1179_U307, P3_R1179_U308, P3_R1179_U309, P3_R1179_U31, P3_R1179_U310, P3_R1179_U311, P3_R1179_U312, P3_R1179_U313, P3_R1179_U314, P3_R1179_U315, P3_R1179_U316, P3_R1179_U317, P3_R1179_U318, P3_R1179_U319, P3_R1179_U32, P3_R1179_U320, P3_R1179_U321, P3_R1179_U322, P3_R1179_U323, P3_R1179_U324, P3_R1179_U325, P3_R1179_U326, P3_R1179_U327, P3_R1179_U328, P3_R1179_U329, P3_R1179_U33, P3_R1179_U330, P3_R1179_U331, P3_R1179_U332, P3_R1179_U333, P3_R1179_U334, P3_R1179_U335, P3_R1179_U336, P3_R1179_U337, P3_R1179_U338, P3_R1179_U339, P3_R1179_U34, P3_R1179_U340, P3_R1179_U341, P3_R1179_U342, P3_R1179_U343, P3_R1179_U344, P3_R1179_U345, P3_R1179_U346, P3_R1179_U347, P3_R1179_U348, P3_R1179_U349, P3_R1179_U35, P3_R1179_U350, P3_R1179_U351, P3_R1179_U352, P3_R1179_U353, P3_R1179_U354, P3_R1179_U355, P3_R1179_U356, P3_R1179_U357, P3_R1179_U358, P3_R1179_U359, P3_R1179_U36, P3_R1179_U360, P3_R1179_U361, P3_R1179_U362, P3_R1179_U363, P3_R1179_U364, P3_R1179_U365, P3_R1179_U366, P3_R1179_U367, P3_R1179_U368, P3_R1179_U369, P3_R1179_U37, P3_R1179_U370, P3_R1179_U371, P3_R1179_U372, P3_R1179_U373, P3_R1179_U374, P3_R1179_U375, P3_R1179_U376, P3_R1179_U377, P3_R1179_U378, P3_R1179_U379, P3_R1179_U38, P3_R1179_U380, P3_R1179_U381, P3_R1179_U382, P3_R1179_U383, P3_R1179_U384, P3_R1179_U385, P3_R1179_U386, P3_R1179_U387, P3_R1179_U388, P3_R1179_U389, P3_R1179_U39, P3_R1179_U390, P3_R1179_U391, P3_R1179_U392, P3_R1179_U393, P3_R1179_U394, P3_R1179_U395, P3_R1179_U396, P3_R1179_U397, P3_R1179_U398, P3_R1179_U399, P3_R1179_U40, P3_R1179_U400, P3_R1179_U401, P3_R1179_U402, P3_R1179_U403, P3_R1179_U404, P3_R1179_U405, P3_R1179_U406, P3_R1179_U407, P3_R1179_U408, P3_R1179_U409, P3_R1179_U41, P3_R1179_U410, P3_R1179_U411, P3_R1179_U412, P3_R1179_U413, P3_R1179_U414, P3_R1179_U415, P3_R1179_U416, P3_R1179_U417, P3_R1179_U418, P3_R1179_U419, P3_R1179_U42, P3_R1179_U420, P3_R1179_U421, P3_R1179_U422, P3_R1179_U423, P3_R1179_U424, P3_R1179_U425, P3_R1179_U426, P3_R1179_U427, P3_R1179_U428, P3_R1179_U429, P3_R1179_U43, P3_R1179_U430, P3_R1179_U431, P3_R1179_U432, P3_R1179_U433, P3_R1179_U434, P3_R1179_U435, P3_R1179_U436, P3_R1179_U437, P3_R1179_U438, P3_R1179_U439, P3_R1179_U44, P3_R1179_U440, P3_R1179_U441, P3_R1179_U442, P3_R1179_U443, P3_R1179_U444, P3_R1179_U445, P3_R1179_U446, P3_R1179_U447, P3_R1179_U448, P3_R1179_U449, P3_R1179_U45, P3_R1179_U450, P3_R1179_U451, P3_R1179_U452, P3_R1179_U453, P3_R1179_U454, P3_R1179_U455, P3_R1179_U456, P3_R1179_U457, P3_R1179_U458, P3_R1179_U459, P3_R1179_U46, P3_R1179_U460, P3_R1179_U461, P3_R1179_U462, P3_R1179_U463, P3_R1179_U464, P3_R1179_U465, P3_R1179_U466, P3_R1179_U467, P3_R1179_U468, P3_R1179_U469, P3_R1179_U47, P3_R1179_U470, P3_R1179_U471, P3_R1179_U472, P3_R1179_U473, P3_R1179_U474, P3_R1179_U475, P3_R1179_U476, P3_R1179_U477, P3_R1179_U478, P3_R1179_U479, P3_R1179_U48, P3_R1179_U480, P3_R1179_U481, P3_R1179_U482, P3_R1179_U483, P3_R1179_U484, P3_R1179_U485, P3_R1179_U49, P3_R1179_U50, P3_R1179_U51, P3_R1179_U52, P3_R1179_U53, P3_R1179_U54, P3_R1179_U55, P3_R1179_U56, P3_R1179_U57, P3_R1179_U58, P3_R1179_U59, P3_R1179_U6, P3_R1179_U60, P3_R1179_U61, P3_R1179_U62, P3_R1179_U63, P3_R1179_U64, P3_R1179_U65, P3_R1179_U66, P3_R1179_U67, P3_R1179_U68, P3_R1179_U69, P3_R1179_U7, P3_R1179_U70, P3_R1179_U71, P3_R1179_U72, P3_R1179_U73, P3_R1179_U74, P3_R1179_U75, P3_R1179_U76, P3_R1179_U77, P3_R1179_U78, P3_R1179_U79, P3_R1179_U8, P3_R1179_U80, P3_R1179_U81, P3_R1179_U82, P3_R1179_U83, P3_R1179_U84, P3_R1179_U85, P3_R1179_U86, P3_R1179_U87, P3_R1179_U88, P3_R1179_U89, P3_R1179_U9, P3_R1179_U90, P3_R1179_U91, P3_R1179_U92, P3_R1179_U93, P3_R1179_U94, P3_R1179_U95, P3_R1179_U96, P3_R1179_U97, P3_R1179_U98, P3_R1179_U99, P3_R1200_U10, P3_R1200_U100, P3_R1200_U101, P3_R1200_U102, P3_R1200_U103, P3_R1200_U104, P3_R1200_U105, P3_R1200_U106, P3_R1200_U107, P3_R1200_U108, P3_R1200_U109, P3_R1200_U11, P3_R1200_U110, P3_R1200_U111, P3_R1200_U112, P3_R1200_U113, P3_R1200_U114, P3_R1200_U115, P3_R1200_U116, P3_R1200_U117, P3_R1200_U118, P3_R1200_U119, P3_R1200_U12, P3_R1200_U120, P3_R1200_U121, P3_R1200_U122, P3_R1200_U123, P3_R1200_U124, P3_R1200_U125, P3_R1200_U126, P3_R1200_U127, P3_R1200_U128, P3_R1200_U129, P3_R1200_U13, P3_R1200_U130, P3_R1200_U131, P3_R1200_U132, P3_R1200_U133, P3_R1200_U134, P3_R1200_U135, P3_R1200_U136, P3_R1200_U137, P3_R1200_U138, P3_R1200_U139, P3_R1200_U14, P3_R1200_U140, P3_R1200_U141, P3_R1200_U142, P3_R1200_U143, P3_R1200_U144, P3_R1200_U145, P3_R1200_U146, P3_R1200_U147, P3_R1200_U148, P3_R1200_U149, P3_R1200_U15, P3_R1200_U150, P3_R1200_U151, P3_R1200_U152, P3_R1200_U153, P3_R1200_U154, P3_R1200_U155, P3_R1200_U156, P3_R1200_U157, P3_R1200_U158, P3_R1200_U159, P3_R1200_U16, P3_R1200_U160, P3_R1200_U161, P3_R1200_U162, P3_R1200_U163, P3_R1200_U164, P3_R1200_U165, P3_R1200_U166, P3_R1200_U167, P3_R1200_U168, P3_R1200_U169, P3_R1200_U17, P3_R1200_U170, P3_R1200_U171, P3_R1200_U172, P3_R1200_U173, P3_R1200_U174, P3_R1200_U175, P3_R1200_U176, P3_R1200_U177, P3_R1200_U178, P3_R1200_U179, P3_R1200_U18, P3_R1200_U180, P3_R1200_U181, P3_R1200_U182, P3_R1200_U183, P3_R1200_U184, P3_R1200_U185, P3_R1200_U186, P3_R1200_U187, P3_R1200_U188, P3_R1200_U189, P3_R1200_U19, P3_R1200_U190, P3_R1200_U191, P3_R1200_U192, P3_R1200_U193, P3_R1200_U194, P3_R1200_U195, P3_R1200_U196, P3_R1200_U197, P3_R1200_U198, P3_R1200_U199, P3_R1200_U20, P3_R1200_U200, P3_R1200_U201, P3_R1200_U202, P3_R1200_U203, P3_R1200_U204, P3_R1200_U205, P3_R1200_U206, P3_R1200_U207, P3_R1200_U208, P3_R1200_U209, P3_R1200_U21, P3_R1200_U210, P3_R1200_U211, P3_R1200_U212, P3_R1200_U213, P3_R1200_U214, P3_R1200_U215, P3_R1200_U216, P3_R1200_U217, P3_R1200_U218, P3_R1200_U219, P3_R1200_U22, P3_R1200_U220, P3_R1200_U221, P3_R1200_U222, P3_R1200_U223, P3_R1200_U224, P3_R1200_U225, P3_R1200_U226, P3_R1200_U227, P3_R1200_U228, P3_R1200_U229, P3_R1200_U23, P3_R1200_U230, P3_R1200_U231, P3_R1200_U232, P3_R1200_U233, P3_R1200_U234, P3_R1200_U235, P3_R1200_U236, P3_R1200_U237, P3_R1200_U238, P3_R1200_U239, P3_R1200_U24, P3_R1200_U240, P3_R1200_U241, P3_R1200_U242, P3_R1200_U243, P3_R1200_U244, P3_R1200_U245, P3_R1200_U246, P3_R1200_U247, P3_R1200_U248, P3_R1200_U249, P3_R1200_U25, P3_R1200_U250, P3_R1200_U251, P3_R1200_U252, P3_R1200_U253, P3_R1200_U254, P3_R1200_U255, P3_R1200_U256, P3_R1200_U257, P3_R1200_U258, P3_R1200_U259, P3_R1200_U26, P3_R1200_U260, P3_R1200_U261, P3_R1200_U262, P3_R1200_U263, P3_R1200_U264, P3_R1200_U265, P3_R1200_U266, P3_R1200_U267, P3_R1200_U268, P3_R1200_U269, P3_R1200_U27, P3_R1200_U270, P3_R1200_U271, P3_R1200_U272, P3_R1200_U273, P3_R1200_U274, P3_R1200_U275, P3_R1200_U276, P3_R1200_U277, P3_R1200_U278, P3_R1200_U279, P3_R1200_U28, P3_R1200_U280, P3_R1200_U281, P3_R1200_U282, P3_R1200_U283, P3_R1200_U284, P3_R1200_U285, P3_R1200_U286, P3_R1200_U287, P3_R1200_U288, P3_R1200_U289, P3_R1200_U29, P3_R1200_U290, P3_R1200_U291, P3_R1200_U292, P3_R1200_U293, P3_R1200_U294, P3_R1200_U295, P3_R1200_U296, P3_R1200_U297, P3_R1200_U298, P3_R1200_U299, P3_R1200_U30, P3_R1200_U300, P3_R1200_U301, P3_R1200_U302, P3_R1200_U303, P3_R1200_U304, P3_R1200_U305, P3_R1200_U306, P3_R1200_U307, P3_R1200_U308, P3_R1200_U309, P3_R1200_U31, P3_R1200_U310, P3_R1200_U311, P3_R1200_U312, P3_R1200_U313, P3_R1200_U314, P3_R1200_U315, P3_R1200_U316, P3_R1200_U317, P3_R1200_U318, P3_R1200_U319, P3_R1200_U32, P3_R1200_U320, P3_R1200_U321, P3_R1200_U322, P3_R1200_U323, P3_R1200_U324, P3_R1200_U325, P3_R1200_U326, P3_R1200_U327, P3_R1200_U328, P3_R1200_U329, P3_R1200_U33, P3_R1200_U330, P3_R1200_U331, P3_R1200_U332, P3_R1200_U333, P3_R1200_U334, P3_R1200_U335, P3_R1200_U336, P3_R1200_U337, P3_R1200_U338, P3_R1200_U339, P3_R1200_U34, P3_R1200_U340, P3_R1200_U341, P3_R1200_U342, P3_R1200_U343, P3_R1200_U344, P3_R1200_U345, P3_R1200_U346, P3_R1200_U347, P3_R1200_U348, P3_R1200_U349, P3_R1200_U35, P3_R1200_U350, P3_R1200_U351, P3_R1200_U352, P3_R1200_U353, P3_R1200_U354, P3_R1200_U355, P3_R1200_U356, P3_R1200_U357, P3_R1200_U358, P3_R1200_U359, P3_R1200_U36, P3_R1200_U360, P3_R1200_U361, P3_R1200_U362, P3_R1200_U363, P3_R1200_U364, P3_R1200_U365, P3_R1200_U366, P3_R1200_U367, P3_R1200_U368, P3_R1200_U369, P3_R1200_U37, P3_R1200_U370, P3_R1200_U371, P3_R1200_U372, P3_R1200_U373, P3_R1200_U374, P3_R1200_U375, P3_R1200_U376, P3_R1200_U377, P3_R1200_U378, P3_R1200_U379, P3_R1200_U38, P3_R1200_U380, P3_R1200_U381, P3_R1200_U382, P3_R1200_U383, P3_R1200_U384, P3_R1200_U385, P3_R1200_U386, P3_R1200_U387, P3_R1200_U388, P3_R1200_U389, P3_R1200_U39, P3_R1200_U390, P3_R1200_U391, P3_R1200_U392, P3_R1200_U393, P3_R1200_U394, P3_R1200_U395, P3_R1200_U396, P3_R1200_U397, P3_R1200_U398, P3_R1200_U399, P3_R1200_U40, P3_R1200_U400, P3_R1200_U401, P3_R1200_U402, P3_R1200_U403, P3_R1200_U404, P3_R1200_U405, P3_R1200_U406, P3_R1200_U407, P3_R1200_U408, P3_R1200_U409, P3_R1200_U41, P3_R1200_U410, P3_R1200_U411, P3_R1200_U412, P3_R1200_U413, P3_R1200_U414, P3_R1200_U415, P3_R1200_U416, P3_R1200_U417, P3_R1200_U418, P3_R1200_U419, P3_R1200_U42, P3_R1200_U420, P3_R1200_U421, P3_R1200_U422, P3_R1200_U423, P3_R1200_U424, P3_R1200_U425, P3_R1200_U426, P3_R1200_U427, P3_R1200_U428, P3_R1200_U429, P3_R1200_U43, P3_R1200_U430, P3_R1200_U431, P3_R1200_U432, P3_R1200_U433, P3_R1200_U434, P3_R1200_U435, P3_R1200_U436, P3_R1200_U437, P3_R1200_U438, P3_R1200_U439, P3_R1200_U44, P3_R1200_U440, P3_R1200_U441, P3_R1200_U442, P3_R1200_U443, P3_R1200_U444, P3_R1200_U445, P3_R1200_U446, P3_R1200_U447, P3_R1200_U448, P3_R1200_U449, P3_R1200_U45, P3_R1200_U450, P3_R1200_U451, P3_R1200_U452, P3_R1200_U453, P3_R1200_U454, P3_R1200_U455, P3_R1200_U456, P3_R1200_U457, P3_R1200_U458, P3_R1200_U459, P3_R1200_U46, P3_R1200_U460, P3_R1200_U461, P3_R1200_U462, P3_R1200_U463, P3_R1200_U464, P3_R1200_U465, P3_R1200_U466, P3_R1200_U467, P3_R1200_U468, P3_R1200_U469, P3_R1200_U47, P3_R1200_U470, P3_R1200_U471, P3_R1200_U472, P3_R1200_U473, P3_R1200_U474, P3_R1200_U475, P3_R1200_U476, P3_R1200_U477, P3_R1200_U478, P3_R1200_U479, P3_R1200_U48, P3_R1200_U480, P3_R1200_U481, P3_R1200_U482, P3_R1200_U483, P3_R1200_U484, P3_R1200_U485, P3_R1200_U49, P3_R1200_U50, P3_R1200_U51, P3_R1200_U52, P3_R1200_U53, P3_R1200_U54, P3_R1200_U55, P3_R1200_U56, P3_R1200_U57, P3_R1200_U58, P3_R1200_U59, P3_R1200_U6, P3_R1200_U60, P3_R1200_U61, P3_R1200_U62, P3_R1200_U63, P3_R1200_U64, P3_R1200_U65, P3_R1200_U66, P3_R1200_U67, P3_R1200_U68, P3_R1200_U69, P3_R1200_U7, P3_R1200_U70, P3_R1200_U71, P3_R1200_U72, P3_R1200_U73, P3_R1200_U74, P3_R1200_U75, P3_R1200_U76, P3_R1200_U77, P3_R1200_U78, P3_R1200_U79, P3_R1200_U8, P3_R1200_U80, P3_R1200_U81, P3_R1200_U82, P3_R1200_U83, P3_R1200_U84, P3_R1200_U85, P3_R1200_U86, P3_R1200_U87, P3_R1200_U88, P3_R1200_U89, P3_R1200_U9, P3_R1200_U90, P3_R1200_U91, P3_R1200_U92, P3_R1200_U93, P3_R1200_U94, P3_R1200_U95, P3_R1200_U96, P3_R1200_U97, P3_R1200_U98, P3_R1200_U99, P3_R1209_U10, P3_R1209_U100, P3_R1209_U101, P3_R1209_U102, P3_R1209_U103, P3_R1209_U104, P3_R1209_U105, P3_R1209_U106, P3_R1209_U107, P3_R1209_U108, P3_R1209_U109, P3_R1209_U11, P3_R1209_U110, P3_R1209_U111, P3_R1209_U112, P3_R1209_U113, P3_R1209_U114, P3_R1209_U115, P3_R1209_U116, P3_R1209_U117, P3_R1209_U118, P3_R1209_U119, P3_R1209_U12, P3_R1209_U120, P3_R1209_U121, P3_R1209_U122, P3_R1209_U123, P3_R1209_U124, P3_R1209_U125, P3_R1209_U126, P3_R1209_U127, P3_R1209_U128, P3_R1209_U129, P3_R1209_U13, P3_R1209_U130, P3_R1209_U131, P3_R1209_U132, P3_R1209_U133, P3_R1209_U134, P3_R1209_U135, P3_R1209_U136, P3_R1209_U137, P3_R1209_U138, P3_R1209_U139, P3_R1209_U14, P3_R1209_U140, P3_R1209_U141, P3_R1209_U142, P3_R1209_U143, P3_R1209_U144, P3_R1209_U145, P3_R1209_U146, P3_R1209_U147, P3_R1209_U148, P3_R1209_U149, P3_R1209_U15, P3_R1209_U150, P3_R1209_U151, P3_R1209_U152, P3_R1209_U153, P3_R1209_U154, P3_R1209_U155, P3_R1209_U156, P3_R1209_U157, P3_R1209_U158, P3_R1209_U159, P3_R1209_U16, P3_R1209_U160, P3_R1209_U161, P3_R1209_U162, P3_R1209_U163, P3_R1209_U164, P3_R1209_U165, P3_R1209_U166, P3_R1209_U167, P3_R1209_U168, P3_R1209_U169, P3_R1209_U17, P3_R1209_U170, P3_R1209_U171, P3_R1209_U172, P3_R1209_U173, P3_R1209_U174, P3_R1209_U175, P3_R1209_U176, P3_R1209_U177, P3_R1209_U178, P3_R1209_U179, P3_R1209_U18, P3_R1209_U180, P3_R1209_U181, P3_R1209_U182, P3_R1209_U183, P3_R1209_U184, P3_R1209_U185, P3_R1209_U186, P3_R1209_U187, P3_R1209_U188, P3_R1209_U189, P3_R1209_U19, P3_R1209_U190, P3_R1209_U191, P3_R1209_U192, P3_R1209_U193, P3_R1209_U194, P3_R1209_U195, P3_R1209_U196, P3_R1209_U197, P3_R1209_U198, P3_R1209_U199, P3_R1209_U20, P3_R1209_U200, P3_R1209_U201, P3_R1209_U202, P3_R1209_U203, P3_R1209_U204, P3_R1209_U205, P3_R1209_U206, P3_R1209_U207, P3_R1209_U208, P3_R1209_U209, P3_R1209_U21, P3_R1209_U210, P3_R1209_U211, P3_R1209_U212, P3_R1209_U213, P3_R1209_U214, P3_R1209_U215, P3_R1209_U216, P3_R1209_U217, P3_R1209_U218, P3_R1209_U219, P3_R1209_U22, P3_R1209_U220, P3_R1209_U221, P3_R1209_U222, P3_R1209_U223, P3_R1209_U224, P3_R1209_U225, P3_R1209_U226, P3_R1209_U227, P3_R1209_U228, P3_R1209_U229, P3_R1209_U23, P3_R1209_U230, P3_R1209_U231, P3_R1209_U232, P3_R1209_U233, P3_R1209_U234, P3_R1209_U235, P3_R1209_U236, P3_R1209_U237, P3_R1209_U238, P3_R1209_U239, P3_R1209_U24, P3_R1209_U240, P3_R1209_U241, P3_R1209_U242, P3_R1209_U243, P3_R1209_U244, P3_R1209_U245, P3_R1209_U246, P3_R1209_U247, P3_R1209_U248, P3_R1209_U249, P3_R1209_U25, P3_R1209_U250, P3_R1209_U251, P3_R1209_U252, P3_R1209_U253, P3_R1209_U254, P3_R1209_U255, P3_R1209_U256, P3_R1209_U257, P3_R1209_U258, P3_R1209_U259, P3_R1209_U26, P3_R1209_U260, P3_R1209_U261, P3_R1209_U262, P3_R1209_U263, P3_R1209_U264, P3_R1209_U265, P3_R1209_U266, P3_R1209_U267, P3_R1209_U268, P3_R1209_U269, P3_R1209_U27, P3_R1209_U270, P3_R1209_U271, P3_R1209_U272, P3_R1209_U273, P3_R1209_U274, P3_R1209_U275, P3_R1209_U276, P3_R1209_U28, P3_R1209_U29, P3_R1209_U30, P3_R1209_U31, P3_R1209_U32, P3_R1209_U33, P3_R1209_U34, P3_R1209_U35, P3_R1209_U36, P3_R1209_U37, P3_R1209_U38, P3_R1209_U39, P3_R1209_U40, P3_R1209_U41, P3_R1209_U42, P3_R1209_U43, P3_R1209_U44, P3_R1209_U45, P3_R1209_U46, P3_R1209_U47, P3_R1209_U48, P3_R1209_U49, P3_R1209_U50, P3_R1209_U51, P3_R1209_U52, P3_R1209_U53, P3_R1209_U54, P3_R1209_U55, P3_R1209_U56, P3_R1209_U57, P3_R1209_U58, P3_R1209_U59, P3_R1209_U6, P3_R1209_U60, P3_R1209_U61, P3_R1209_U62, P3_R1209_U63, P3_R1209_U64, P3_R1209_U65, P3_R1209_U66, P3_R1209_U67, P3_R1209_U68, P3_R1209_U69, P3_R1209_U7, P3_R1209_U70, P3_R1209_U71, P3_R1209_U72, P3_R1209_U73, P3_R1209_U74, P3_R1209_U75, P3_R1209_U76, P3_R1209_U77, P3_R1209_U78, P3_R1209_U79, P3_R1209_U8, P3_R1209_U80, P3_R1209_U81, P3_R1209_U82, P3_R1209_U83, P3_R1209_U84, P3_R1209_U85, P3_R1209_U86, P3_R1209_U87, P3_R1209_U88, P3_R1209_U89, P3_R1209_U9, P3_R1209_U90, P3_R1209_U91, P3_R1209_U92, P3_R1209_U93, P3_R1209_U94, P3_R1209_U95, P3_R1209_U96, P3_R1209_U97, P3_R1209_U98, P3_R1209_U99, P3_R1212_U10, P3_R1212_U100, P3_R1212_U101, P3_R1212_U102, P3_R1212_U103, P3_R1212_U104, P3_R1212_U105, P3_R1212_U106, P3_R1212_U107, P3_R1212_U108, P3_R1212_U109, P3_R1212_U11, P3_R1212_U110, P3_R1212_U111, P3_R1212_U112, P3_R1212_U113, P3_R1212_U114, P3_R1212_U115, P3_R1212_U116, P3_R1212_U117, P3_R1212_U118, P3_R1212_U119, P3_R1212_U12, P3_R1212_U120, P3_R1212_U121, P3_R1212_U122, P3_R1212_U123, P3_R1212_U124, P3_R1212_U125, P3_R1212_U126, P3_R1212_U127, P3_R1212_U128, P3_R1212_U129, P3_R1212_U13, P3_R1212_U130, P3_R1212_U131, P3_R1212_U132, P3_R1212_U133, P3_R1212_U134, P3_R1212_U135, P3_R1212_U136, P3_R1212_U137, P3_R1212_U138, P3_R1212_U139, P3_R1212_U14, P3_R1212_U140, P3_R1212_U141, P3_R1212_U142, P3_R1212_U143, P3_R1212_U144, P3_R1212_U145, P3_R1212_U146, P3_R1212_U147, P3_R1212_U148, P3_R1212_U149, P3_R1212_U15, P3_R1212_U150, P3_R1212_U151, P3_R1212_U152, P3_R1212_U153, P3_R1212_U154, P3_R1212_U155, P3_R1212_U156, P3_R1212_U157, P3_R1212_U158, P3_R1212_U159, P3_R1212_U16, P3_R1212_U160, P3_R1212_U161, P3_R1212_U162, P3_R1212_U163, P3_R1212_U164, P3_R1212_U165, P3_R1212_U166, P3_R1212_U167, P3_R1212_U168, P3_R1212_U169, P3_R1212_U17, P3_R1212_U170, P3_R1212_U171, P3_R1212_U172, P3_R1212_U173, P3_R1212_U174, P3_R1212_U175, P3_R1212_U176, P3_R1212_U177, P3_R1212_U178, P3_R1212_U179, P3_R1212_U18, P3_R1212_U180, P3_R1212_U181, P3_R1212_U182, P3_R1212_U183, P3_R1212_U184, P3_R1212_U185, P3_R1212_U186, P3_R1212_U187, P3_R1212_U188, P3_R1212_U189, P3_R1212_U19, P3_R1212_U190, P3_R1212_U191, P3_R1212_U192, P3_R1212_U193, P3_R1212_U194, P3_R1212_U195, P3_R1212_U196, P3_R1212_U197, P3_R1212_U198, P3_R1212_U199, P3_R1212_U20, P3_R1212_U200, P3_R1212_U201, P3_R1212_U202, P3_R1212_U203, P3_R1212_U204, P3_R1212_U205, P3_R1212_U206, P3_R1212_U207, P3_R1212_U208, P3_R1212_U209, P3_R1212_U21, P3_R1212_U210, P3_R1212_U211, P3_R1212_U212, P3_R1212_U213, P3_R1212_U214, P3_R1212_U215, P3_R1212_U216, P3_R1212_U217, P3_R1212_U218, P3_R1212_U219, P3_R1212_U22, P3_R1212_U220, P3_R1212_U221, P3_R1212_U222, P3_R1212_U223, P3_R1212_U224, P3_R1212_U225, P3_R1212_U226, P3_R1212_U227, P3_R1212_U228, P3_R1212_U229, P3_R1212_U23, P3_R1212_U230, P3_R1212_U231, P3_R1212_U232, P3_R1212_U233, P3_R1212_U234, P3_R1212_U235, P3_R1212_U236, P3_R1212_U237, P3_R1212_U238, P3_R1212_U239, P3_R1212_U24, P3_R1212_U240, P3_R1212_U241, P3_R1212_U242, P3_R1212_U243, P3_R1212_U244, P3_R1212_U245, P3_R1212_U246, P3_R1212_U247, P3_R1212_U248, P3_R1212_U249, P3_R1212_U25, P3_R1212_U250, P3_R1212_U251, P3_R1212_U252, P3_R1212_U253, P3_R1212_U254, P3_R1212_U255, P3_R1212_U256, P3_R1212_U257, P3_R1212_U258, P3_R1212_U259, P3_R1212_U26, P3_R1212_U260, P3_R1212_U261, P3_R1212_U262, P3_R1212_U263, P3_R1212_U264, P3_R1212_U265, P3_R1212_U266, P3_R1212_U267, P3_R1212_U268, P3_R1212_U269, P3_R1212_U27, P3_R1212_U270, P3_R1212_U271, P3_R1212_U272, P3_R1212_U273, P3_R1212_U274, P3_R1212_U275, P3_R1212_U276, P3_R1212_U28, P3_R1212_U29, P3_R1212_U30, P3_R1212_U31, P3_R1212_U32, P3_R1212_U33, P3_R1212_U34, P3_R1212_U35, P3_R1212_U36, P3_R1212_U37, P3_R1212_U38, P3_R1212_U39, P3_R1212_U40, P3_R1212_U41, P3_R1212_U42, P3_R1212_U43, P3_R1212_U44, P3_R1212_U45, P3_R1212_U46, P3_R1212_U47, P3_R1212_U48, P3_R1212_U49, P3_R1212_U50, P3_R1212_U51, P3_R1212_U52, P3_R1212_U53, P3_R1212_U54, P3_R1212_U55, P3_R1212_U56, P3_R1212_U57, P3_R1212_U58, P3_R1212_U59, P3_R1212_U6, P3_R1212_U60, P3_R1212_U61, P3_R1212_U62, P3_R1212_U63, P3_R1212_U64, P3_R1212_U65, P3_R1212_U66, P3_R1212_U67, P3_R1212_U68, P3_R1212_U69, P3_R1212_U7, P3_R1212_U70, P3_R1212_U71, P3_R1212_U72, P3_R1212_U73, P3_R1212_U74, P3_R1212_U75, P3_R1212_U76, P3_R1212_U77, P3_R1212_U78, P3_R1212_U79, P3_R1212_U8, P3_R1212_U80, P3_R1212_U81, P3_R1212_U82, P3_R1212_U83, P3_R1212_U84, P3_R1212_U85, P3_R1212_U86, P3_R1212_U87, P3_R1212_U88, P3_R1212_U89, P3_R1212_U9, P3_R1212_U90, P3_R1212_U91, P3_R1212_U92, P3_R1212_U93, P3_R1212_U94, P3_R1212_U95, P3_R1212_U96, P3_R1212_U97, P3_R1212_U98, P3_R1212_U99, P3_R1269_U10, P3_R1269_U100, P3_R1269_U101, P3_R1269_U102, P3_R1269_U103, P3_R1269_U104, P3_R1269_U105, P3_R1269_U106, P3_R1269_U107, P3_R1269_U108, P3_R1269_U109, P3_R1269_U11, P3_R1269_U110, P3_R1269_U111, P3_R1269_U112, P3_R1269_U113, P3_R1269_U114, P3_R1269_U115, P3_R1269_U116, P3_R1269_U117, P3_R1269_U118, P3_R1269_U119, P3_R1269_U12, P3_R1269_U120, P3_R1269_U121, P3_R1269_U122, P3_R1269_U123, P3_R1269_U124, P3_R1269_U125, P3_R1269_U126, P3_R1269_U127, P3_R1269_U128, P3_R1269_U129, P3_R1269_U13, P3_R1269_U130, P3_R1269_U131, P3_R1269_U132, P3_R1269_U133, P3_R1269_U134, P3_R1269_U135, P3_R1269_U136, P3_R1269_U137, P3_R1269_U138, P3_R1269_U139, P3_R1269_U14, P3_R1269_U140, P3_R1269_U141, P3_R1269_U142, P3_R1269_U143, P3_R1269_U144, P3_R1269_U145, P3_R1269_U146, P3_R1269_U147, P3_R1269_U148, P3_R1269_U149, P3_R1269_U15, P3_R1269_U150, P3_R1269_U151, P3_R1269_U152, P3_R1269_U153, P3_R1269_U154, P3_R1269_U155, P3_R1269_U156, P3_R1269_U157, P3_R1269_U158, P3_R1269_U159, P3_R1269_U16, P3_R1269_U160, P3_R1269_U161, P3_R1269_U162, P3_R1269_U163, P3_R1269_U164, P3_R1269_U165, P3_R1269_U166, P3_R1269_U167, P3_R1269_U168, P3_R1269_U169, P3_R1269_U17, P3_R1269_U170, P3_R1269_U171, P3_R1269_U172, P3_R1269_U173, P3_R1269_U174, P3_R1269_U175, P3_R1269_U176, P3_R1269_U177, P3_R1269_U178, P3_R1269_U179, P3_R1269_U18, P3_R1269_U180, P3_R1269_U181, P3_R1269_U182, P3_R1269_U183, P3_R1269_U184, P3_R1269_U185, P3_R1269_U186, P3_R1269_U187, P3_R1269_U188, P3_R1269_U189, P3_R1269_U19, P3_R1269_U190, P3_R1269_U191, P3_R1269_U192, P3_R1269_U193, P3_R1269_U194, P3_R1269_U195, P3_R1269_U196, P3_R1269_U197, P3_R1269_U198, P3_R1269_U199, P3_R1269_U20, P3_R1269_U200, P3_R1269_U201, P3_R1269_U202, P3_R1269_U21, P3_R1269_U22, P3_R1269_U23, P3_R1269_U24, P3_R1269_U25, P3_R1269_U26, P3_R1269_U27, P3_R1269_U28, P3_R1269_U29, P3_R1269_U30, P3_R1269_U31, P3_R1269_U32, P3_R1269_U33, P3_R1269_U34, P3_R1269_U35, P3_R1269_U36, P3_R1269_U37, P3_R1269_U38, P3_R1269_U39, P3_R1269_U40, P3_R1269_U41, P3_R1269_U42, P3_R1269_U43, P3_R1269_U44, P3_R1269_U45, P3_R1269_U46, P3_R1269_U47, P3_R1269_U48, P3_R1269_U49, P3_R1269_U50, P3_R1269_U51, P3_R1269_U52, P3_R1269_U53, P3_R1269_U54, P3_R1269_U55, P3_R1269_U56, P3_R1269_U57, P3_R1269_U58, P3_R1269_U59, P3_R1269_U6, P3_R1269_U60, P3_R1269_U61, P3_R1269_U62, P3_R1269_U63, P3_R1269_U64, P3_R1269_U65, P3_R1269_U66, P3_R1269_U67, P3_R1269_U68, P3_R1269_U69, P3_R1269_U7, P3_R1269_U70, P3_R1269_U71, P3_R1269_U72, P3_R1269_U73, P3_R1269_U74, P3_R1269_U75, P3_R1269_U76, P3_R1269_U77, P3_R1269_U78, P3_R1269_U79, P3_R1269_U8, P3_R1269_U80, P3_R1269_U81, P3_R1269_U82, P3_R1269_U83, P3_R1269_U84, P3_R1269_U85, P3_R1269_U86, P3_R1269_U87, P3_R1269_U88, P3_R1269_U89, P3_R1269_U9, P3_R1269_U90, P3_R1269_U91, P3_R1269_U92, P3_R1269_U93, P3_R1269_U94, P3_R1269_U95, P3_R1269_U96, P3_R1269_U97, P3_R1269_U98, P3_R1269_U99, P3_R1297_U6, P3_R1297_U7, P3_R1300_U10, P3_R1300_U6, P3_R1300_U7, P3_R1300_U8, P3_R1300_U9, P3_R693_U10, P3_R693_U100, P3_R693_U101, P3_R693_U102, P3_R693_U103, P3_R693_U104, P3_R693_U105, P3_R693_U106, P3_R693_U107, P3_R693_U108, P3_R693_U109, P3_R693_U11, P3_R693_U110, P3_R693_U111, P3_R693_U112, P3_R693_U113, P3_R693_U114, P3_R693_U115, P3_R693_U116, P3_R693_U117, P3_R693_U118, P3_R693_U119, P3_R693_U12, P3_R693_U120, P3_R693_U121, P3_R693_U122, P3_R693_U123, P3_R693_U124, P3_R693_U125, P3_R693_U126, P3_R693_U127, P3_R693_U128, P3_R693_U129, P3_R693_U13, P3_R693_U130, P3_R693_U131, P3_R693_U132, P3_R693_U133, P3_R693_U134, P3_R693_U135, P3_R693_U136, P3_R693_U137, P3_R693_U138, P3_R693_U139, P3_R693_U14, P3_R693_U140, P3_R693_U141, P3_R693_U142, P3_R693_U143, P3_R693_U144, P3_R693_U145, P3_R693_U146, P3_R693_U147, P3_R693_U148, P3_R693_U149, P3_R693_U15, P3_R693_U150, P3_R693_U151, P3_R693_U152, P3_R693_U153, P3_R693_U154, P3_R693_U155, P3_R693_U156, P3_R693_U157, P3_R693_U158, P3_R693_U159, P3_R693_U16, P3_R693_U160, P3_R693_U161, P3_R693_U162, P3_R693_U163, P3_R693_U164, P3_R693_U165, P3_R693_U166, P3_R693_U167, P3_R693_U168, P3_R693_U169, P3_R693_U17, P3_R693_U170, P3_R693_U171, P3_R693_U172, P3_R693_U173, P3_R693_U174, P3_R693_U175, P3_R693_U176, P3_R693_U177, P3_R693_U178, P3_R693_U179, P3_R693_U18, P3_R693_U180, P3_R693_U181, P3_R693_U182, P3_R693_U183, P3_R693_U184, P3_R693_U185, P3_R693_U186, P3_R693_U187, P3_R693_U188, P3_R693_U189, P3_R693_U19, P3_R693_U190, P3_R693_U191, P3_R693_U192, P3_R693_U193, P3_R693_U194, P3_R693_U195, P3_R693_U196, P3_R693_U20, P3_R693_U21, P3_R693_U22, P3_R693_U23, P3_R693_U24, P3_R693_U25, P3_R693_U26, P3_R693_U27, P3_R693_U28, P3_R693_U29, P3_R693_U30, P3_R693_U31, P3_R693_U32, P3_R693_U33, P3_R693_U34, P3_R693_U35, P3_R693_U36, P3_R693_U37, P3_R693_U38, P3_R693_U39, P3_R693_U40, P3_R693_U41, P3_R693_U42, P3_R693_U43, P3_R693_U44, P3_R693_U45, P3_R693_U46, P3_R693_U47, P3_R693_U48, P3_R693_U49, P3_R693_U50, P3_R693_U51, P3_R693_U52, P3_R693_U53, P3_R693_U54, P3_R693_U55, P3_R693_U56, P3_R693_U57, P3_R693_U58, P3_R693_U59, P3_R693_U6, P3_R693_U60, P3_R693_U61, P3_R693_U62, P3_R693_U63, P3_R693_U64, P3_R693_U65, P3_R693_U66, P3_R693_U67, P3_R693_U68, P3_R693_U69, P3_R693_U7, P3_R693_U70, P3_R693_U71, P3_R693_U72, P3_R693_U73, P3_R693_U74, P3_R693_U75, P3_R693_U76, P3_R693_U77, P3_R693_U78, P3_R693_U79, P3_R693_U8, P3_R693_U80, P3_R693_U81, P3_R693_U82, P3_R693_U83, P3_R693_U84, P3_R693_U85, P3_R693_U86, P3_R693_U87, P3_R693_U88, P3_R693_U89, P3_R693_U9, P3_R693_U90, P3_R693_U91, P3_R693_U92, P3_R693_U93, P3_R693_U94, P3_R693_U95, P3_R693_U96, P3_R693_U97, P3_R693_U98, P3_R693_U99, P3_SUB_598_U10, P3_SUB_598_U100, P3_SUB_598_U101, P3_SUB_598_U102, P3_SUB_598_U103, P3_SUB_598_U104, P3_SUB_598_U105, P3_SUB_598_U106, P3_SUB_598_U107, P3_SUB_598_U108, P3_SUB_598_U109, P3_SUB_598_U11, P3_SUB_598_U110, P3_SUB_598_U111, P3_SUB_598_U112, P3_SUB_598_U113, P3_SUB_598_U114, P3_SUB_598_U115, P3_SUB_598_U116, P3_SUB_598_U117, P3_SUB_598_U118, P3_SUB_598_U119, P3_SUB_598_U12, P3_SUB_598_U120, P3_SUB_598_U121, P3_SUB_598_U122, P3_SUB_598_U123, P3_SUB_598_U124, P3_SUB_598_U125, P3_SUB_598_U126, P3_SUB_598_U127, P3_SUB_598_U128, P3_SUB_598_U129, P3_SUB_598_U13, P3_SUB_598_U130, P3_SUB_598_U131, P3_SUB_598_U132, P3_SUB_598_U133, P3_SUB_598_U134, P3_SUB_598_U135, P3_SUB_598_U136, P3_SUB_598_U137, P3_SUB_598_U138, P3_SUB_598_U139, P3_SUB_598_U14, P3_SUB_598_U140, P3_SUB_598_U141, P3_SUB_598_U142, P3_SUB_598_U143, P3_SUB_598_U144, P3_SUB_598_U145, P3_SUB_598_U146, P3_SUB_598_U147, P3_SUB_598_U148, P3_SUB_598_U149, P3_SUB_598_U15, P3_SUB_598_U150, P3_SUB_598_U151, P3_SUB_598_U152, P3_SUB_598_U153, P3_SUB_598_U154, P3_SUB_598_U155, P3_SUB_598_U156, P3_SUB_598_U157, P3_SUB_598_U158, P3_SUB_598_U159, P3_SUB_598_U16, P3_SUB_598_U160, P3_SUB_598_U17, P3_SUB_598_U18, P3_SUB_598_U19, P3_SUB_598_U20, P3_SUB_598_U21, P3_SUB_598_U22, P3_SUB_598_U23, P3_SUB_598_U24, P3_SUB_598_U25, P3_SUB_598_U26, P3_SUB_598_U27, P3_SUB_598_U28, P3_SUB_598_U29, P3_SUB_598_U30, P3_SUB_598_U31, P3_SUB_598_U32, P3_SUB_598_U33, P3_SUB_598_U34, P3_SUB_598_U35, P3_SUB_598_U36, P3_SUB_598_U37, P3_SUB_598_U38, P3_SUB_598_U39, P3_SUB_598_U40, P3_SUB_598_U41, P3_SUB_598_U42, P3_SUB_598_U43, P3_SUB_598_U44, P3_SUB_598_U45, P3_SUB_598_U46, P3_SUB_598_U47, P3_SUB_598_U48, P3_SUB_598_U49, P3_SUB_598_U50, P3_SUB_598_U51, P3_SUB_598_U52, P3_SUB_598_U53, P3_SUB_598_U54, P3_SUB_598_U55, P3_SUB_598_U56, P3_SUB_598_U57, P3_SUB_598_U58, P3_SUB_598_U59, P3_SUB_598_U6, P3_SUB_598_U60, P3_SUB_598_U61, P3_SUB_598_U62, P3_SUB_598_U63, P3_SUB_598_U64, P3_SUB_598_U65, P3_SUB_598_U66, P3_SUB_598_U67, P3_SUB_598_U68, P3_SUB_598_U69, P3_SUB_598_U7, P3_SUB_598_U70, P3_SUB_598_U71, P3_SUB_598_U72, P3_SUB_598_U73, P3_SUB_598_U74, P3_SUB_598_U75, P3_SUB_598_U76, P3_SUB_598_U77, P3_SUB_598_U78, P3_SUB_598_U79, P3_SUB_598_U8, P3_SUB_598_U80, P3_SUB_598_U81, P3_SUB_598_U82, P3_SUB_598_U83, P3_SUB_598_U84, P3_SUB_598_U85, P3_SUB_598_U86, P3_SUB_598_U87, P3_SUB_598_U88, P3_SUB_598_U89, P3_SUB_598_U9, P3_SUB_598_U90, P3_SUB_598_U91, P3_SUB_598_U92, P3_SUB_598_U93, P3_SUB_598_U94, P3_SUB_598_U95, P3_SUB_598_U96, P3_SUB_598_U97, P3_SUB_598_U98, P3_SUB_598_U99, P3_SUB_609_U10, P3_SUB_609_U100, P3_SUB_609_U101, P3_SUB_609_U102, P3_SUB_609_U103, P3_SUB_609_U104, P3_SUB_609_U105, P3_SUB_609_U106, P3_SUB_609_U107, P3_SUB_609_U108, P3_SUB_609_U109, P3_SUB_609_U11, P3_SUB_609_U110, P3_SUB_609_U111, P3_SUB_609_U112, P3_SUB_609_U113, P3_SUB_609_U114, P3_SUB_609_U115, P3_SUB_609_U12, P3_SUB_609_U13, P3_SUB_609_U14, P3_SUB_609_U15, P3_SUB_609_U16, P3_SUB_609_U17, P3_SUB_609_U18, P3_SUB_609_U19, P3_SUB_609_U20, P3_SUB_609_U21, P3_SUB_609_U22, P3_SUB_609_U23, P3_SUB_609_U24, P3_SUB_609_U25, P3_SUB_609_U26, P3_SUB_609_U27, P3_SUB_609_U28, P3_SUB_609_U29, P3_SUB_609_U30, P3_SUB_609_U31, P3_SUB_609_U32, P3_SUB_609_U33, P3_SUB_609_U34, P3_SUB_609_U35, P3_SUB_609_U36, P3_SUB_609_U37, P3_SUB_609_U38, P3_SUB_609_U39, P3_SUB_609_U40, P3_SUB_609_U41, P3_SUB_609_U42, P3_SUB_609_U43, P3_SUB_609_U44, P3_SUB_609_U45, P3_SUB_609_U46, P3_SUB_609_U47, P3_SUB_609_U48, P3_SUB_609_U49, P3_SUB_609_U50, P3_SUB_609_U51, P3_SUB_609_U52, P3_SUB_609_U53, P3_SUB_609_U54, P3_SUB_609_U55, P3_SUB_609_U56, P3_SUB_609_U57, P3_SUB_609_U58, P3_SUB_609_U59, P3_SUB_609_U6, P3_SUB_609_U60, P3_SUB_609_U61, P3_SUB_609_U62, P3_SUB_609_U63, P3_SUB_609_U64, P3_SUB_609_U65, P3_SUB_609_U66, P3_SUB_609_U67, P3_SUB_609_U68, P3_SUB_609_U69, P3_SUB_609_U7, P3_SUB_609_U70, P3_SUB_609_U71, P3_SUB_609_U72, P3_SUB_609_U73, P3_SUB_609_U74, P3_SUB_609_U75, P3_SUB_609_U76, P3_SUB_609_U77, P3_SUB_609_U78, P3_SUB_609_U79, P3_SUB_609_U8, P3_SUB_609_U80, P3_SUB_609_U81, P3_SUB_609_U82, P3_SUB_609_U83, P3_SUB_609_U84, P3_SUB_609_U85, P3_SUB_609_U86, P3_SUB_609_U87, P3_SUB_609_U88, P3_SUB_609_U89, P3_SUB_609_U9, P3_SUB_609_U90, P3_SUB_609_U91, P3_SUB_609_U92, P3_SUB_609_U93, P3_SUB_609_U94, P3_SUB_609_U95, P3_SUB_609_U96, P3_SUB_609_U97, P3_SUB_609_U98, P3_SUB_609_U99, P3_U3013, P3_U3014, P3_U3015, P3_U3016, P3_U3017, P3_U3018, P3_U3019, P3_U3020, P3_U3021, P3_U3022, P3_U3023, P3_U3024, P3_U3025, P3_U3026, P3_U3027, P3_U3028, P3_U3029, P3_U3030, P3_U3031, P3_U3032, P3_U3033, P3_U3034, P3_U3035, P3_U3036, P3_U3037, P3_U3038, P3_U3039, P3_U3040, P3_U3041, P3_U3042, P3_U3043, P3_U3044, P3_U3045, P3_U3046, P3_U3047, P3_U3048, P3_U3049, P3_U3050, P3_U3051, P3_U3052, P3_U3053, P3_U3054, P3_U3055, P3_U3056, P3_U3057, P3_U3058, P3_U3059, P3_U3060, P3_U3061, P3_U3062, P3_U3063, P3_U3064, P3_U3065, P3_U3066, P3_U3067, P3_U3068, P3_U3069, P3_U3070, P3_U3071, P3_U3072, P3_U3073, P3_U3074, P3_U3075, P3_U3076, P3_U3077, P3_U3078, P3_U3079, P3_U3080, P3_U3081, P3_U3082, P3_U3083, P3_U3084, P3_U3085, P3_U3086, P3_U3087, P3_U3088, P3_U3089, P3_U3090, P3_U3091, P3_U3092, P3_U3093, P3_U3094, P3_U3095, P3_U3096, P3_U3097, P3_U3098, P3_U3099, P3_U3100, P3_U3101, P3_U3102, P3_U3103, P3_U3104, P3_U3105, P3_U3106, P3_U3107, P3_U3108, P3_U3109, P3_U3110, P3_U3111, P3_U3112, P3_U3113, P3_U3114, P3_U3115, P3_U3116, P3_U3117, P3_U3118, P3_U3119, P3_U3120, P3_U3121, P3_U3122, P3_U3123, P3_U3124, P3_U3125, P3_U3126, P3_U3127, P3_U3128, P3_U3129, P3_U3130, P3_U3131, P3_U3132, P3_U3133, P3_U3134, P3_U3135, P3_U3136, P3_U3137, P3_U3138, P3_U3139, P3_U3140, P3_U3141, P3_U3142, P3_U3143, P3_U3144, P3_U3145, P3_U3146, P3_U3147, P3_U3148, P3_U3149, P3_U3152, P3_U3297, P3_U3298, P3_U3299, P3_U3300, P3_U3301, P3_U3302, P3_U3303, P3_U3304, P3_U3305, P3_U3306, P3_U3307, P3_U3308, P3_U3309, P3_U3310, P3_U3311, P3_U3312, P3_U3313, P3_U3314, P3_U3315, P3_U3316, P3_U3317, P3_U3318, P3_U3319, P3_U3320, P3_U3321, P3_U3322, P3_U3323, P3_U3324, P3_U3325, P3_U3326, P3_U3327, P3_U3328, P3_U3329, P3_U3330, P3_U3331, P3_U3332, P3_U3333, P3_U3334, P3_U3335, P3_U3336, P3_U3337, P3_U3338, P3_U3339, P3_U3340, P3_U3341, P3_U3342, P3_U3343, P3_U3344, P3_U3345, P3_U3346, P3_U3347, P3_U3348, P3_U3349, P3_U3350, P3_U3351, P3_U3352, P3_U3353, P3_U3354, P3_U3355, P3_U3356, P3_U3357, P3_U3358, P3_U3359, P3_U3360, P3_U3361, P3_U3362, P3_U3363, P3_U3364, P3_U3365, P3_U3366, P3_U3367, P3_U3368, P3_U3369, P3_U3370, P3_U3371, P3_U3372, P3_U3373, P3_U3374, P3_U3375, P3_U3378, P3_U3379, P3_U3380, P3_U3381, P3_U3382, P3_U3383, P3_U3384, P3_U3385, P3_U3386, P3_U3387, P3_U3388, P3_U3389, P3_U3391, P3_U3392, P3_U3394, P3_U3395, P3_U3397, P3_U3398, P3_U3400, P3_U3401, P3_U3403, P3_U3404, P3_U3406, P3_U3407, P3_U3409, P3_U3410, P3_U3412, P3_U3413, P3_U3415, P3_U3416, P3_U3418, P3_U3419, P3_U3421, P3_U3422, P3_U3424, P3_U3425, P3_U3427, P3_U3428, P3_U3430, P3_U3431, P3_U3433, P3_U3434, P3_U3436, P3_U3437, P3_U3439, P3_U3440, P3_U3442, P3_U3443, P3_U3445, P3_U3523, P3_U3524, P3_U3525, P3_U3526, P3_U3527, P3_U3528, P3_U3529, P3_U3530, P3_U3531, P3_U3532, P3_U3533, P3_U3534, P3_U3535, P3_U3536, P3_U3537, P3_U3538, P3_U3539, P3_U3540, P3_U3541, P3_U3542, P3_U3543, P3_U3544, P3_U3545, P3_U3546, P3_U3547, P3_U3548, P3_U3549, P3_U3550, P3_U3551, P3_U3552, P3_U3553, P3_U3554, P3_U3555, P3_U3556, P3_U3557, P3_U3558, P3_U3559, P3_U3560, P3_U3561, P3_U3562, P3_U3563, P3_U3564, P3_U3565, P3_U3566, P3_U3567, P3_U3568, P3_U3569, P3_U3570, P3_U3571, P3_U3572, P3_U3573, P3_U3574, P3_U3575, P3_U3576, P3_U3577, P3_U3578, P3_U3579, P3_U3580, P3_U3581, P3_U3582, P3_U3583, P3_U3584, P3_U3585, P3_U3586, P3_U3587, P3_U3588, P3_U3589, P3_U3590, P3_U3591, P3_U3592, P3_U3593, P3_U3594, P3_U3595, P3_U3596, P3_U3597, P3_U3598, P3_U3599, P3_U3600, P3_U3601, P3_U3602, P3_U3603, P3_U3604, P3_U3605, P3_U3606, P3_U3607, P3_U3608, P3_U3609, P3_U3610, P3_U3611, P3_U3612, P3_U3613, P3_U3614, P3_U3615, P3_U3616, P3_U3617, P3_U3618, P3_U3619, P3_U3620, P3_U3621, P3_U3622, P3_U3623, P3_U3624, P3_U3625, P3_U3626, P3_U3627, P3_U3628, P3_U3629, P3_U3630, P3_U3631, P3_U3632, P3_U3633, P3_U3634, P3_U3635, P3_U3636, P3_U3637, P3_U3638, P3_U3639, P3_U3640, P3_U3641, P3_U3642, P3_U3643, P3_U3644, P3_U3645, P3_U3646, P3_U3647, P3_U3648, P3_U3649, P3_U3650, P3_U3651, P3_U3652, P3_U3653, P3_U3654, P3_U3655, P3_U3656, P3_U3657, P3_U3658, P3_U3659, P3_U3660, P3_U3661, P3_U3662, P3_U3663, P3_U3664, P3_U3665, P3_U3666, P3_U3667, P3_U3668, P3_U3669, P3_U3670, P3_U3671, P3_U3672, P3_U3673, P3_U3674, P3_U3675, P3_U3676, P3_U3677, P3_U3678, P3_U3679, P3_U3680, P3_U3681, P3_U3682, P3_U3683, P3_U3684, P3_U3685, P3_U3686, P3_U3687, P3_U3688, P3_U3689, P3_U3690, P3_U3691, P3_U3692, P3_U3693, P3_U3694, P3_U3695, P3_U3696, P3_U3697, P3_U3698, P3_U3699, P3_U3700, P3_U3701, P3_U3702, P3_U3703, P3_U3704, P3_U3705, P3_U3706, P3_U3707, P3_U3708, P3_U3709, P3_U3710, P3_U3711, P3_U3712, P3_U3713, P3_U3714, P3_U3715, P3_U3716, P3_U3717, P3_U3718, P3_U3719, P3_U3720, P3_U3721, P3_U3722, P3_U3723, P3_U3724, P3_U3725, P3_U3726, P3_U3727, P3_U3728, P3_U3729, P3_U3730, P3_U3731, P3_U3732, P3_U3733, P3_U3734, P3_U3735, P3_U3736, P3_U3737, P3_U3738, P3_U3739, P3_U3740, P3_U3741, P3_U3742, P3_U3743, P3_U3744, P3_U3745, P3_U3746, P3_U3747, P3_U3748, P3_U3749, P3_U3750, P3_U3751, P3_U3752, P3_U3753, P3_U3754, P3_U3755, P3_U3756, P3_U3757, P3_U3758, P3_U3759, P3_U3760, P3_U3761, P3_U3762, P3_U3763, P3_U3764, P3_U3765, P3_U3766, P3_U3767, P3_U3768, P3_U3769, P3_U3770, P3_U3771, P3_U3772, P3_U3773, P3_U3774, P3_U3775, P3_U3776, P3_U3777, P3_U3778, P3_U3779, P3_U3780, P3_U3781, P3_U3782, P3_U3783, P3_U3784, P3_U3785, P3_U3786, P3_U3787, P3_U3788, P3_U3789, P3_U3790, P3_U3791, P3_U3792, P3_U3793, P3_U3794, P3_U3795, P3_U3796, P3_U3797, P3_U3798, P3_U3799, P3_U3800, P3_U3801, P3_U3802, P3_U3803, P3_U3804, P3_U3805, P3_U3806, P3_U3807, P3_U3808, P3_U3809, P3_U3810, P3_U3811, P3_U3812, P3_U3813, P3_U3814, P3_U3815, P3_U3816, P3_U3817, P3_U3818, P3_U3819, P3_U3820, P3_U3821, P3_U3822, P3_U3823, P3_U3824, P3_U3825, P3_U3826, P3_U3827, P3_U3828, P3_U3829, P3_U3830, P3_U3831, P3_U3832, P3_U3833, P3_U3834, P3_U3835, P3_U3836, P3_U3837, P3_U3838, P3_U3839, P3_U3840, P3_U3841, P3_U3842, P3_U3843, P3_U3844, P3_U3845, P3_U3846, P3_U3847, P3_U3848, P3_U3849, P3_U3850, P3_U3851, P3_U3852, P3_U3853, P3_U3854, P3_U3855, P3_U3856, P3_U3857, P3_U3858, P3_U3859, P3_U3860, P3_U3861, P3_U3862, P3_U3863, P3_U3864, P3_U3865, P3_U3866, P3_U3867, P3_U3868, P3_U3869, P3_U3870, P3_U3871, P3_U3872, P3_U3873, P3_U3874, P3_U3875, P3_U3876, P3_U3877, P3_U3878, P3_U3879, P3_U3880, P3_U3881, P3_U3882, P3_U3883, P3_U3884, P3_U3885, P3_U3886, P3_U3887, P3_U3888, P3_U3889, P3_U3890, P3_U3891, P3_U3892, P3_U3893, P3_U3894, P3_U3895, P3_U3896, P3_U3898, P3_U3899, P3_U3900, P3_U3901, P3_U3902, P3_U3903, P3_U3904, P3_U3905, P3_U3906, P3_U3907, P3_U3908, P3_U3909, P3_U3910, P3_U3911, P3_U3912, P3_U3913, P3_U3914, P3_U3915, P3_U3916, P3_U3917, P3_U3918, P3_U3919, P3_U3920, P3_U3921, P3_U3922, P3_U3923, P3_U3924, P3_U3925, P3_U3926, P3_U3927, P3_U3928, P3_U3929, P3_U3930, P3_U3931, P3_U3932, P3_U3933, P3_U3934, P3_U3935, P3_U3936, P3_U3937, P3_U3938, P3_U3939, P3_U3940, P3_U3941, P3_U3942, P3_U3943, P3_U3944, P3_U3945, P3_U3946, P3_U3947, P3_U3948, P3_U3949, P3_U3950, P3_U3951, P3_U3952, P3_U3953, P3_U3954, P3_U3955, P3_U3956, P3_U3957, P3_U3958, P3_U3959, P3_U3960, P3_U3961, P3_U3962, P3_U3963, P3_U3964, P3_U3965, P3_U3966, P3_U3967, P3_U3968, P3_U3969, P3_U3970, P3_U3971, P3_U3972, P3_U3973, P3_U3974, P3_U3975, P3_U3976, P3_U3977, P3_U3978, P3_U3979, P3_U3980, P3_U3981, P3_U3982, P3_U3983, P3_U3984, P3_U3985, P3_U3986, P3_U3987, P3_U3988, P3_U3989, P3_U3990, P3_U3991, P3_U3992, P3_U3993, P3_U3994, P3_U3995, P3_U3996, P3_U3997, P3_U3998, P3_U3999, P3_U4000, P3_U4001, P3_U4002, P3_U4003, P3_U4004, P3_U4005, P3_U4006, P3_U4007, P3_U4008, P3_U4009, P3_U4010, P3_U4011, P3_U4012, P3_U4013, P3_U4014, P3_U4015, P3_U4016, P3_U4017, P3_U4018, P3_U4019, P3_U4020, P3_U4021, P3_U4022, P3_U4023, P3_U4024, P3_U4025, P3_U4026, P3_U4027, P3_U4028, P3_U4029, P3_U4030, P3_U4031, P3_U4032, P3_U4033, P3_U4034, P3_U4035, P3_U4036, P3_U4037, P3_U4038, P3_U4039, P3_U4040, P3_U4041, P3_U4042, P3_U4043, P3_U4044, P3_U4045, P3_U4046, P3_U4047, P3_U4048, P3_U4049, P3_U4050, P3_U4051, P3_U4052, P3_U4053, P3_U4054, P3_U4055, P3_U4056, P3_U4057, P3_U4058, P3_U4059, P3_U4060, P3_U4061, P3_U4062, P3_U4063, P3_U4064, P3_U4065, P3_U4066, P3_U4067, P3_U4068, P3_U4069, P3_U4070, P3_U4071, P3_U4072, P3_U4073, P3_U4074, P3_U4075, P3_U4076, P3_U4077, P3_U4078, P3_U4079, P3_U4080, P3_U4081, P3_U4082, P3_U4083, P3_U4084, P3_U4085, P3_U4086, P3_U4087, P3_U4088, P3_U4089, P3_U4090, P3_U4091, P3_U4092, P3_U4093, P3_U4094, P3_U4095, P3_U4096, P3_U4097, P3_U4098, P3_U4099, P3_U4100, P3_U4101, P3_U4102, P3_U4103, P3_U4104, P3_U4105, P3_U4106, P3_U4107, P3_U4108, P3_U4109, P3_U4110, P3_U4111, P3_U4112, P3_U4113, P3_U4114, P3_U4115, P3_U4116, P3_U4117, P3_U4118, P3_U4119, P3_U4120, P3_U4121, P3_U4122, P3_U4123, P3_U4124, P3_U4125, P3_U4126, P3_U4127, P3_U4128, P3_U4129, P3_U4130, P3_U4131, P3_U4132, P3_U4133, P3_U4134, P3_U4135, P3_U4136, P3_U4137, P3_U4138, P3_U4139, P3_U4140, P3_U4141, P3_U4142, P3_U4143, P3_U4144, P3_U4145, P3_U4146, P3_U4147, P3_U4148, P3_U4149, P3_U4150, P3_U4151, P3_U4152, P3_U4153, P3_U4154, P3_U4155, P3_U4156, P3_U4157, P3_U4158, P3_U4159, P3_U4160, P3_U4161, P3_U4162, P3_U4163, P3_U4164, P3_U4165, P3_U4166, P3_U4167, P3_U4168, P3_U4169, P3_U4170, P3_U4171, P3_U4172, P3_U4173, P3_U4174, P3_U4175, P3_U4176, P3_U4177, P3_U4178, P3_U4179, P3_U4180, P3_U4181, P3_U4182, P3_U4183, P3_U4184, P3_U4185, P3_U4186, P3_U4187, P3_U4188, P3_U4189, P3_U4190, P3_U4191, P3_U4192, P3_U4193, P3_U4194, P3_U4195, P3_U4196, P3_U4197, P3_U4198, P3_U4199, P3_U4200, P3_U4201, P3_U4202, P3_U4203, P3_U4204, P3_U4205, P3_U4206, P3_U4207, P3_U4208, P3_U4209, P3_U4210, P3_U4211, P3_U4212, P3_U4213, P3_U4214, P3_U4215, P3_U4216, P3_U4217, P3_U4218, P3_U4219, P3_U4220, P3_U4221, P3_U4222, P3_U4223, P3_U4224, P3_U4225, P3_U4226, P3_U4227, P3_U4228, P3_U4229, P3_U4230, P3_U4231, P3_U4232, P3_U4233, P3_U4234, P3_U4235, P3_U4236, P3_U4237, P3_U4238, P3_U4239, P3_U4240, P3_U4241, P3_U4242, P3_U4243, P3_U4244, P3_U4245, P3_U4246, P3_U4247, P3_U4248, P3_U4249, P3_U4250, P3_U4251, P3_U4252, P3_U4253, P3_U4254, P3_U4255, P3_U4256, P3_U4257, P3_U4258, P3_U4259, P3_U4260, P3_U4261, P3_U4262, P3_U4263, P3_U4264, P3_U4265, P3_U4266, P3_U4267, P3_U4268, P3_U4269, P3_U4270, P3_U4271, P3_U4272, P3_U4273, P3_U4274, P3_U4275, P3_U4276, P3_U4277, P3_U4278, P3_U4279, P3_U4280, P3_U4281, P3_U4282, P3_U4283, P3_U4284, P3_U4285, P3_U4286, P3_U4287, P3_U4288, P3_U4289, P3_U4290, P3_U4291, P3_U4292, P3_U4293, P3_U4294, P3_U4295, P3_U4296, P3_U4297, P3_U4298, P3_U4299, P3_U4300, P3_U4301, P3_U4302, P3_U4303, P3_U4304, P3_U4305, P3_U4306, P3_U4307, P3_U4308, P3_U4309, P3_U4310, P3_U4311, P3_U4312, P3_U4313, P3_U4314, P3_U4315, P3_U4316, P3_U4317, P3_U4318, P3_U4319, P3_U4320, P3_U4321, P3_U4322, P3_U4323, P3_U4324, P3_U4325, P3_U4326, P3_U4327, P3_U4328, P3_U4329, P3_U4330, P3_U4331, P3_U4332, P3_U4333, P3_U4334, P3_U4335, P3_U4336, P3_U4337, P3_U4338, P3_U4339, P3_U4340, P3_U4341, P3_U4342, P3_U4343, P3_U4344, P3_U4345, P3_U4346, P3_U4347, P3_U4348, P3_U4349, P3_U4350, P3_U4351, P3_U4352, P3_U4353, P3_U4354, P3_U4355, P3_U4356, P3_U4357, P3_U4358, P3_U4359, P3_U4360, P3_U4361, P3_U4362, P3_U4363, P3_U4364, P3_U4365, P3_U4366, P3_U4367, P3_U4368, P3_U4369, P3_U4370, P3_U4371, P3_U4372, P3_U4373, P3_U4374, P3_U4375, P3_U4376, P3_U4377, P3_U4378, P3_U4379, P3_U4380, P3_U4381, P3_U4382, P3_U4383, P3_U4384, P3_U4385, P3_U4386, P3_U4387, P3_U4388, P3_U4389, P3_U4390, P3_U4391, P3_U4392, P3_U4393, P3_U4394, P3_U4395, P3_U4396, P3_U4397, P3_U4398, P3_U4399, P3_U4400, P3_U4401, P3_U4402, P3_U4403, P3_U4404, P3_U4405, P3_U4406, P3_U4407, P3_U4408, P3_U4409, P3_U4410, P3_U4411, P3_U4412, P3_U4413, P3_U4414, P3_U4415, P3_U4416, P3_U4417, P3_U4418, P3_U4419, P3_U4420, P3_U4421, P3_U4422, P3_U4423, P3_U4424, P3_U4425, P3_U4426, P3_U4427, P3_U4428, P3_U4429, P3_U4430, P3_U4431, P3_U4432, P3_U4433, P3_U4434, P3_U4435, P3_U4436, P3_U4437, P3_U4438, P3_U4439, P3_U4440, P3_U4441, P3_U4442, P3_U4443, P3_U4444, P3_U4445, P3_U4446, P3_U4447, P3_U4448, P3_U4449, P3_U4450, P3_U4451, P3_U4452, P3_U4453, P3_U4454, P3_U4455, P3_U4456, P3_U4457, P3_U4458, P3_U4459, P3_U4460, P3_U4461, P3_U4462, P3_U4463, P3_U4464, P3_U4465, P3_U4466, P3_U4467, P3_U4468, P3_U4469, P3_U4470, P3_U4471, P3_U4472, P3_U4473, P3_U4474, P3_U4475, P3_U4476, P3_U4477, P3_U4478, P3_U4479, P3_U4480, P3_U4481, P3_U4482, P3_U4483, P3_U4484, P3_U4485, P3_U4486, P3_U4487, P3_U4488, P3_U4489, P3_U4490, P3_U4491, P3_U4492, P3_U4493, P3_U4494, P3_U4495, P3_U4496, P3_U4497, P3_U4498, P3_U4499, P3_U4500, P3_U4501, P3_U4502, P3_U4503, P3_U4504, P3_U4505, P3_U4506, P3_U4507, P3_U4508, P3_U4509, P3_U4510, P3_U4511, P3_U4512, P3_U4513, P3_U4514, P3_U4515, P3_U4516, P3_U4517, P3_U4518, P3_U4519, P3_U4520, P3_U4521, P3_U4522, P3_U4523, P3_U4524, P3_U4525, P3_U4526, P3_U4527, P3_U4528, P3_U4529, P3_U4530, P3_U4531, P3_U4532, P3_U4533, P3_U4534, P3_U4535, P3_U4536, P3_U4537, P3_U4538, P3_U4539, P3_U4540, P3_U4541, P3_U4542, P3_U4543, P3_U4544, P3_U4545, P3_U4546, P3_U4547, P3_U4548, P3_U4549, P3_U4550, P3_U4551, P3_U4552, P3_U4553, P3_U4554, P3_U4555, P3_U4556, P3_U4557, P3_U4558, P3_U4559, P3_U4560, P3_U4561, P3_U4562, P3_U4563, P3_U4564, P3_U4565, P3_U4566, P3_U4567, P3_U4568, P3_U4569, P3_U4570, P3_U4571, P3_U4572, P3_U4573, P3_U4574, P3_U4575, P3_U4576, P3_U4577, P3_U4578, P3_U4579, P3_U4580, P3_U4581, P3_U4582, P3_U4583, P3_U4584, P3_U4585, P3_U4586, P3_U4587, P3_U4588, P3_U4589, P3_U4590, P3_U4591, P3_U4592, P3_U4593, P3_U4594, P3_U4595, P3_U4596, P3_U4597, P3_U4598, P3_U4599, P3_U4600, P3_U4601, P3_U4602, P3_U4603, P3_U4604, P3_U4605, P3_U4606, P3_U4607, P3_U4608, P3_U4609, P3_U4610, P3_U4611, P3_U4612, P3_U4613, P3_U4614, P3_U4615, P3_U4616, P3_U4617, P3_U4618, P3_U4619, P3_U4620, P3_U4621, P3_U4622, P3_U4623, P3_U4624, P3_U4625, P3_U4626, P3_U4627, P3_U4628, P3_U4629, P3_U4630, P3_U4631, P3_U4632, P3_U4633, P3_U4634, P3_U4635, P3_U4636, P3_U4637, P3_U4638, P3_U4639, P3_U4640, P3_U4641, P3_U4642, P3_U4643, P3_U4644, P3_U4645, P3_U4646, P3_U4647, P3_U4648, P3_U4649, P3_U4650, P3_U4651, P3_U4652, P3_U4653, P3_U4654, P3_U4655, P3_U4656, P3_U4657, P3_U4658, P3_U4659, P3_U4660, P3_U4661, P3_U4662, P3_U4663, P3_U4664, P3_U4665, P3_U4666, P3_U4667, P3_U4668, P3_U4669, P3_U4670, P3_U4671, P3_U4672, P3_U4673, P3_U4674, P3_U4675, P3_U4676, P3_U4677, P3_U4678, P3_U4679, P3_U4680, P3_U4681, P3_U4682, P3_U4683, P3_U4684, P3_U4685, P3_U4686, P3_U4687, P3_U4688, P3_U4689, P3_U4690, P3_U4691, P3_U4692, P3_U4693, P3_U4694, P3_U4695, P3_U4696, P3_U4697, P3_U4698, P3_U4699, P3_U4700, P3_U4701, P3_U4702, P3_U4703, P3_U4704, P3_U4705, P3_U4706, P3_U4707, P3_U4708, P3_U4709, P3_U4710, P3_U4711, P3_U4712, P3_U4713, P3_U4714, P3_U4715, P3_U4716, P3_U4717, P3_U4718, P3_U4719, P3_U4720, P3_U4721, P3_U4722, P3_U4723, P3_U4724, P3_U4725, P3_U4726, P3_U4727, P3_U4728, P3_U4729, P3_U4730, P3_U4731, P3_U4732, P3_U4733, P3_U4734, P3_U4735, P3_U4736, P3_U4737, P3_U4738, P3_U4739, P3_U4740, P3_U4741, P3_U4742, P3_U4743, P3_U4744, P3_U4745, P3_U4746, P3_U4747, P3_U4748, P3_U4749, P3_U4750, P3_U4751, P3_U4752, P3_U4753, P3_U4754, P3_U4755, P3_U4756, P3_U4757, P3_U4758, P3_U4759, P3_U4760, P3_U4761, P3_U4762, P3_U4763, P3_U4764, P3_U4765, P3_U4766, P3_U4767, P3_U4768, P3_U4769, P3_U4770, P3_U4771, P3_U4772, P3_U4773, P3_U4774, P3_U4775, P3_U4776, P3_U4777, P3_U4778, P3_U4779, P3_U4780, P3_U4781, P3_U4782, P3_U4783, P3_U4784, P3_U4785, P3_U4786, P3_U4787, P3_U4788, P3_U4789, P3_U4790, P3_U4791, P3_U4792, P3_U4793, P3_U4794, P3_U4795, P3_U4796, P3_U4797, P3_U4798, P3_U4799, P3_U4800, P3_U4801, P3_U4802, P3_U4803, P3_U4804, P3_U4805, P3_U4806, P3_U4807, P3_U4808, P3_U4809, P3_U4810, P3_U4811, P3_U4812, P3_U4813, P3_U4814, P3_U4815, P3_U4816, P3_U4817, P3_U4818, P3_U4819, P3_U4820, P3_U4821, P3_U4822, P3_U4823, P3_U4824, P3_U4825, P3_U4826, P3_U4827, P3_U4828, P3_U4829, P3_U4830, P3_U4831, P3_U4832, P3_U4833, P3_U4834, P3_U4835, P3_U4836, P3_U4837, P3_U4838, P3_U4839, P3_U4840, P3_U4841, P3_U4842, P3_U4843, P3_U4844, P3_U4845, P3_U4846, P3_U4847, P3_U4848, P3_U4849, P3_U4850, P3_U4851, P3_U4852, P3_U4853, P3_U4854, P3_U4855, P3_U4856, P3_U4857, P3_U4858, P3_U4859, P3_U4860, P3_U4861, P3_U4862, P3_U4863, P3_U4864, P3_U4865, P3_U4866, P3_U4867, P3_U4868, P3_U4869, P3_U4870, P3_U4871, P3_U4872, P3_U4873, P3_U4874, P3_U4875, P3_U4876, P3_U4877, P3_U4878, P3_U4879, P3_U4880, P3_U4881, P3_U4882, P3_U4883, P3_U4884, P3_U4885, P3_U4886, P3_U4887, P3_U4888, P3_U4889, P3_U4890, P3_U4891, P3_U4892, P3_U4893, P3_U4894, P3_U4895, P3_U4896, P3_U4897, P3_U4898, P3_U4899, P3_U4900, P3_U4901, P3_U4902, P3_U4903, P3_U4904, P3_U4905, P3_U4906, P3_U4907, P3_U4908, P3_U4909, P3_U4910, P3_U4911, P3_U4912, P3_U4913, P3_U4914, P3_U4915, P3_U4916, P3_U4917, P3_U4918, P3_U4919, P3_U4920, P3_U4921, P3_U4922, P3_U4923, P3_U4924, P3_U4925, P3_U4926, P3_U4927, P3_U4928, P3_U4929, P3_U4930, P3_U4931, P3_U4932, P3_U4933, P3_U4934, P3_U4935, P3_U4936, P3_U4937, P3_U4938, P3_U4939, P3_U4940, P3_U4941, P3_U4942, P3_U4943, P3_U4944, P3_U4945, P3_U4946, P3_U4947, P3_U4948, P3_U4949, P3_U4950, P3_U4951, P3_U4952, P3_U4953, P3_U4954, P3_U4955, P3_U4956, P3_U4957, P3_U4958, P3_U4959, P3_U4960, P3_U4961, P3_U4962, P3_U4963, P3_U4964, P3_U4965, P3_U4966, P3_U4967, P3_U4968, P3_U4969, P3_U4970, P3_U4971, P3_U4972, P3_U4973, P3_U4974, P3_U4975, P3_U4976, P3_U4977, P3_U4978, P3_U4979, P3_U4980, P3_U4981, P3_U4982, P3_U4983, P3_U4984, P3_U4985, P3_U4986, P3_U4987, P3_U4988, P3_U4989, P3_U4990, P3_U4991, P3_U4992, P3_U4993, P3_U4994, P3_U4995, P3_U4996, P3_U4997, P3_U4998, P3_U4999, P3_U5000, P3_U5001, P3_U5002, P3_U5003, P3_U5004, P3_U5005, P3_U5006, P3_U5007, P3_U5008, P3_U5009, P3_U5010, P3_U5011, P3_U5012, P3_U5013, P3_U5014, P3_U5015, P3_U5016, P3_U5017, P3_U5018, P3_U5019, P3_U5020, P3_U5021, P3_U5022, P3_U5023, P3_U5024, P3_U5025, P3_U5026, P3_U5027, P3_U5028, P3_U5029, P3_U5030, P3_U5031, P3_U5032, P3_U5033, P3_U5034, P3_U5035, P3_U5036, P3_U5037, P3_U5038, P3_U5039, P3_U5040, P3_U5041, P3_U5042, P3_U5043, P3_U5044, P3_U5045, P3_U5046, P3_U5047, P3_U5048, P3_U5049, P3_U5050, P3_U5051, P3_U5052, P3_U5053, P3_U5054, P3_U5055, P3_U5056, P3_U5057, P3_U5058, P3_U5059, P3_U5060, P3_U5061, P3_U5062, P3_U5063, P3_U5064, P3_U5065, P3_U5066, P3_U5067, P3_U5068, P3_U5069, P3_U5070, P3_U5071, P3_U5072, P3_U5073, P3_U5074, P3_U5075, P3_U5076, P3_U5077, P3_U5078, P3_U5079, P3_U5080, P3_U5081, P3_U5082, P3_U5083, P3_U5084, P3_U5085, P3_U5086, P3_U5087, P3_U5088, P3_U5089, P3_U5090, P3_U5091, P3_U5092, P3_U5093, P3_U5094, P3_U5095, P3_U5096, P3_U5097, P3_U5098, P3_U5099, P3_U5100, P3_U5101, P3_U5102, P3_U5103, P3_U5104, P3_U5105, P3_U5106, P3_U5107, P3_U5108, P3_U5109, P3_U5110, P3_U5111, P3_U5112, P3_U5113, P3_U5114, P3_U5115, P3_U5116, P3_U5117, P3_U5118, P3_U5119, P3_U5120, P3_U5121, P3_U5122, P3_U5123, P3_U5124, P3_U5125, P3_U5126, P3_U5127, P3_U5128, P3_U5129, P3_U5130, P3_U5131, P3_U5132, P3_U5133, P3_U5134, P3_U5135, P3_U5136, P3_U5137, P3_U5138, P3_U5139, P3_U5140, P3_U5141, P3_U5142, P3_U5143, P3_U5144, P3_U5145, P3_U5146, P3_U5147, P3_U5148, P3_U5149, P3_U5150, P3_U5151, P3_U5152, P3_U5153, P3_U5154, P3_U5155, P3_U5156, P3_U5157, P3_U5158, P3_U5159, P3_U5160, P3_U5161, P3_U5162, P3_U5163, P3_U5164, P3_U5165, P3_U5166, P3_U5167, P3_U5168, P3_U5169, P3_U5170, P3_U5171, P3_U5172, P3_U5173, P3_U5174, P3_U5175, P3_U5176, P3_U5177, P3_U5178, P3_U5179, P3_U5180, P3_U5181, P3_U5182, P3_U5183, P3_U5184, P3_U5185, P3_U5186, P3_U5187, P3_U5188, P3_U5189, P3_U5190, P3_U5191, P3_U5192, P3_U5193, P3_U5194, P3_U5195, P3_U5196, P3_U5197, P3_U5198, P3_U5199, P3_U5200, P3_U5201, P3_U5202, P3_U5203, P3_U5204, P3_U5205, P3_U5206, P3_U5207, P3_U5208, P3_U5209, P3_U5210, P3_U5211, P3_U5212, P3_U5213, P3_U5214, P3_U5215, P3_U5216, P3_U5217, P3_U5218, P3_U5219, P3_U5220, P3_U5221, P3_U5222, P3_U5223, P3_U5224, P3_U5225, P3_U5226, P3_U5227, P3_U5228, P3_U5229, P3_U5230, P3_U5231, P3_U5232, P3_U5233, P3_U5234, P3_U5235, P3_U5236, P3_U5237, P3_U5238, P3_U5239, P3_U5240, P3_U5241, P3_U5242, P3_U5243, P3_U5244, P3_U5245, P3_U5246, P3_U5247, P3_U5248, P3_U5249, P3_U5250, P3_U5251, P3_U5252, P3_U5253, P3_U5254, P3_U5255, P3_U5256, P3_U5257, P3_U5258, P3_U5259, P3_U5260, P3_U5261, P3_U5262, P3_U5263, P3_U5264, P3_U5265, P3_U5266, P3_U5267, P3_U5268, P3_U5269, P3_U5270, P3_U5271, P3_U5272, P3_U5273, P3_U5274, P3_U5275, P3_U5276, P3_U5277, P3_U5278, P3_U5279, P3_U5280, P3_U5281, P3_U5282, P3_U5283, P3_U5284, P3_U5285, P3_U5286, P3_U5287, P3_U5288, P3_U5289, P3_U5290, P3_U5291, P3_U5292, P3_U5293, P3_U5294, P3_U5295, P3_U5296, P3_U5297, P3_U5298, P3_U5299, P3_U5300, P3_U5301, P3_U5302, P3_U5303, P3_U5304, P3_U5305, P3_U5306, P3_U5307, P3_U5308, P3_U5309, P3_U5310, P3_U5311, P3_U5312, P3_U5313, P3_U5314, P3_U5315, P3_U5316, P3_U5317, P3_U5318, P3_U5319, P3_U5320, P3_U5321, P3_U5322, P3_U5323, P3_U5324, P3_U5325, P3_U5326, P3_U5327, P3_U5328, P3_U5329, P3_U5330, P3_U5331, P3_U5332, P3_U5333, P3_U5334, P3_U5335, P3_U5336, P3_U5337, P3_U5338, P3_U5339, P3_U5340, P3_U5341, P3_U5342, P3_U5343, P3_U5344, P3_U5345, P3_U5346, P3_U5347, P3_U5348, P3_U5349, P3_U5350, P3_U5351, P3_U5352, P3_U5353, P3_U5354, P3_U5355, P3_U5356, P3_U5357, P3_U5358, P3_U5359, P3_U5360, P3_U5361, P3_U5362, P3_U5363, P3_U5364, P3_U5365, P3_U5366, P3_U5367, P3_U5368, P3_U5369, P3_U5370, P3_U5371, P3_U5372, P3_U5373, P3_U5374, P3_U5375, P3_U5376, P3_U5377, P3_U5378, P3_U5379, P3_U5380, P3_U5381, P3_U5382, P3_U5383, P3_U5384, P3_U5385, P3_U5386, P3_U5387, P3_U5388, P3_U5389, P3_U5390, P3_U5391, P3_U5392, P3_U5393, P3_U5394, P3_U5395, P3_U5396, P3_U5397, P3_U5398, P3_U5399, P3_U5400, P3_U5401, P3_U5402, P3_U5403, P3_U5404, P3_U5405, P3_U5406, P3_U5407, P3_U5408, P3_U5409, P3_U5410, P3_U5411, P3_U5412, P3_U5413, P3_U5414, P3_U5415, P3_U5416, P3_U5417, P3_U5418, P3_U5419, P3_U5420, P3_U5421, P3_U5422, P3_U5423, P3_U5424, P3_U5425, P3_U5426, P3_U5427, P3_U5428, P3_U5429, P3_U5430, P3_U5431, P3_U5432, P3_U5433, P3_U5434, P3_U5435, P3_U5436, P3_U5437, P3_U5438, P3_U5439, P3_U5440, P3_U5441, P3_U5442, P3_U5443, P3_U5444, P3_U5445, P3_U5446, P3_U5447, P3_U5448, P3_U5449, P3_U5450, P3_U5451, P3_U5452, P3_U5453, P3_U5454, P3_U5455, P3_U5456, P3_U5457, P3_U5458, P3_U5459, P3_U5460, P3_U5461, P3_U5462, P3_U5463, P3_U5464, P3_U5465, P3_U5466, P3_U5467, P3_U5468, P3_U5469, P3_U5470, P3_U5471, P3_U5472, P3_U5473, P3_U5474, P3_U5475, P3_U5476, P3_U5477, P3_U5478, P3_U5479, P3_U5480, P3_U5481, P3_U5482, P3_U5483, P3_U5484, P3_U5485, P3_U5486, P3_U5487, P3_U5488, P3_U5489, P3_U5490, P3_U5491, P3_U5492, P3_U5493, P3_U5494, P3_U5495, P3_U5496, P3_U5497, P3_U5498, P3_U5499, P3_U5500, P3_U5501, P3_U5502, P3_U5503, P3_U5504, P3_U5505, P3_U5506, P3_U5507, P3_U5508, P3_U5509, P3_U5510, P3_U5511, P3_U5512, P3_U5513, P3_U5514, P3_U5515, P3_U5516, P3_U5517, P3_U5518, P3_U5519, P3_U5520, P3_U5521, P3_U5522, P3_U5523, P3_U5524, P3_U5525, P3_U5526, P3_U5527, P3_U5528, P3_U5529, P3_U5530, P3_U5531, P3_U5532, P3_U5533, P3_U5534, P3_U5535, P3_U5536, P3_U5537, P3_U5538, P3_U5539, P3_U5540, P3_U5541, P3_U5542, P3_U5543, P3_U5544, P3_U5545, P3_U5546, P3_U5547, P3_U5548, P3_U5549, P3_U5550, P3_U5551, P3_U5552, P3_U5553, P3_U5554, P3_U5555, P3_U5556, P3_U5557, P3_U5558, P3_U5559, P3_U5560, P3_U5561, P3_U5562, P3_U5563, P3_U5564, P3_U5565, P3_U5566, P3_U5567, P3_U5568, P3_U5569, P3_U5570, P3_U5571, P3_U5572, P3_U5573, P3_U5574, P3_U5575, P3_U5576, P3_U5577, P3_U5578, P3_U5579, P3_U5580, P3_U5581, P3_U5582, P3_U5583, P3_U5584, P3_U5585, P3_U5586, P3_U5587, P3_U5588, P3_U5589, P3_U5590, P3_U5591, P3_U5592, P3_U5593, P3_U5594, P3_U5595, P3_U5596, P3_U5597, P3_U5598, P3_U5599, P3_U5600, P3_U5601, P3_U5602, P3_U5603, P3_U5604, P3_U5605, P3_U5606, P3_U5607, P3_U5608, P3_U5609, P3_U5610, P3_U5611, P3_U5612, P3_U5613, P3_U5614, P3_U5615, P3_U5616, P3_U5617, P3_U5618, P3_U5619, P3_U5620, P3_U5621, P3_U5622, P3_U5623, P3_U5624, P3_U5625, P3_U5626, P3_U5627, P3_U5628, P3_U5629, P3_U5630, P3_U5631, P3_U5632, P3_U5633, P3_U5634, P3_U5635, P3_U5636, P3_U5637, P3_U5638, P3_U5639, P3_U5640, P3_U5641, P3_U5642, P3_U5643, P3_U5644, P3_U5645, P3_U5646, P3_U5647, P3_U5648, P3_U5649, P3_U5650, P3_U5651, P3_U5652, P3_U5653, P3_U5654, P3_U5655, P3_U5656, P3_U5657, P3_U5658, P3_U5659, P3_U5660, P3_U5661, P3_U5662, P3_U5663, P3_U5664, P3_U5665, P3_U5666, P3_U5667, P3_U5668, P3_U5669, P3_U5670, P3_U5671, P3_U5672, P3_U5673, P3_U5674, P3_U5675, P3_U5676, P3_U5677, P3_U5678, P3_U5679, P3_U5680, P3_U5681, P3_U5682, P3_U5683, P3_U5684, P3_U5685, P3_U5686, P3_U5687, P3_U5688, P3_U5689, P3_U5690, P3_U5691, P3_U5692, P3_U5693, P3_U5694, P3_U5695, P3_U5696, P3_U5697, P3_U5698, P3_U5699, P3_U5700, P3_U5701, P3_U5702, P3_U5703, P3_U5704, P3_U5705, P3_U5706, P3_U5707, P3_U5708, P3_U5709, P3_U5710, P3_U5711, P3_U5712, P3_U5713, P3_U5714, P3_U5715, P3_U5716, P3_U5717, P3_U5718, P3_U5719, P3_U5720, P3_U5721, P3_U5722, P3_U5723, P3_U5724, P3_U5725, P3_U5726, P3_U5727, P3_U5728, P3_U5729, P3_U5730, P3_U5731, P3_U5732, P3_U5733, P3_U5734, P3_U5735, P3_U5736, P3_U5737, P3_U5738, P3_U5739, P3_U5740, P3_U5741, P3_U5742, P3_U5743, P3_U5744, P3_U5745, P3_U5746, P3_U5747, P3_U5748, P3_U5749, P3_U5750, P3_U5751, P3_U5752, P3_U5753, P3_U5754, P3_U5755, P3_U5756, P3_U5757, P3_U5758, P3_U5759, P3_U5760, P3_U5761, P3_U5762, P3_U5763, P3_U5764, P3_U5765, P3_U5766, P3_U5767, P3_U5768, P3_U5769, P3_U5770, P3_U5771, P3_U5772, P3_U5773, P3_U5774, P3_U5775, P3_U5776, P3_U5777, P3_U5778, P3_U5779, P3_U5780, P3_U5781, P3_U5782, P3_U5783, P3_U5784, P3_U5785, P3_U5786, P3_U5787, P3_U5788, P3_U5789, P3_U5790, P3_U5791, P3_U5792, P3_U5793, P3_U5794, P3_U5795, P3_U5796, P3_U5797, P3_U5798, P3_U5799, P3_U5800, P3_U5801, P3_U5802, P3_U5803, P3_U5804, P3_U5805, P3_U5806, P3_U5807, P3_U5808, P3_U5809, P3_U5810, P3_U5811, P3_U5812, P3_U5813, P3_U5814, P3_U5815, P3_U5816, P3_U5817, P3_U5818, P3_U5819, P3_U5820, P3_U5821, P3_U5822, P3_U5823, P3_U5824, P3_U5825, P3_U5826, P3_U5827, P3_U5828, P3_U5829, P3_U5830, P3_U5831, P3_U5832, P3_U5833, P3_U5834, P3_U5835, P3_U5836, P3_U5837, P3_U5838, P3_U5839, P3_U5840, P3_U5841, P3_U5842, P3_U5843, P3_U5844, P3_U5845, P3_U5846, P3_U5847, P3_U5848, P3_U5849, P3_U5850, P3_U5851, P3_U5852, P3_U5853, P3_U5854, P3_U5855, P3_U5856, P3_U5857, P3_U5858, P3_U5859, P3_U5860, P3_U5861, P3_U5862, P3_U5863, P3_U5864, P3_U5865, P3_U5866, P3_U5867, P3_U5868, P3_U5869, P3_U5870, P3_U5871, P3_U5872, P3_U5873, P3_U5874, P3_U5875, P3_U5876, P3_U5877, P3_U5878, P3_U5879, P3_U5880, P3_U5881, P3_U5882, P3_U5883, P3_U5884, P3_U5885, P3_U5886, P3_U5887, P3_U5888, P3_U5889, P3_U5890, P3_U5891, P3_U5892, P3_U5893, P3_U5894, P3_U5895, P3_U5896, P3_U5897, P3_U5898, P3_U5899, P3_U5900, P3_U5901, P3_U5902, P3_U5903, P3_U5904, P3_U5905, P3_U5906, P3_U5907, P3_U5908, P3_U5909, P3_U5910, P3_U5911, P3_U5912, P3_U5913, P3_U5914, P3_U5915, P3_U5916, P3_U5917, P3_U5918, P3_U5919, P3_U5920, P3_U5921, P3_U5922, P3_U5923, P3_U5924, P3_U5925, P3_U5926, P3_U5927, P3_U5928, P3_U5929, P3_U5930, P3_U5931, P3_U5932, P3_U5933, P3_U5934, P3_U5935, P3_U5936, P3_U5937, P3_U5938, P3_U5939, P3_U5940, P3_U5941, P3_U5942, P3_U5943, P3_U5944, P3_U5945, P3_U5946, P3_U5947, P3_U5948, P3_U5949, P3_U5950, P3_U5951, P3_U5952, P3_U5953, P3_U5954, P3_U5955, P3_U5956, P3_U5957, P3_U5958, P3_U5959, P3_U5960, P3_U5961, P3_U5962, P3_U5963, P3_U5964, P3_U5965, P3_U5966, P3_U5967, P3_U5968, P3_U5969, P3_U5970, P3_U5971, P3_U5972, P3_U5973, P3_U5974, P3_U5975, P3_U5976, P3_U5977, P3_U5978, P3_U5979, P3_U5980, P3_U5981, P3_U5982, P3_U5983, P3_U5984, P3_U5985, P3_U5986, P3_U5987, P3_U5988, P3_U5989, P3_U5990, P3_U5991, P3_U5992, P3_U5993, P3_U5994, P3_U5995, P3_U5996, P3_U5997, P3_U5998, P3_U5999, P3_U6000, P3_U6001, P3_U6002, P3_U6003, P3_U6004, P3_U6005, P3_U6006, P3_U6007, P3_U6008, P3_U6009, P3_U6010, P3_U6011, P3_U6012, P3_U6013, P3_U6014, P3_U6015, P3_U6016, P3_U6017, P3_U6018, P3_U6019, P3_U6020, P3_U6021, P3_U6022, P3_U6023, P3_U6024, P3_U6025, P3_U6026, P3_U6027, P3_U6028, P3_U6029, P3_U6030, P3_U6031, P3_U6032, P3_U6033, P3_U6034, P3_U6035, P3_U6036, P3_U6037, P3_U6038, P3_U6039, P3_U6040, P3_U6041, P3_U6042, P3_U6043, P3_U6044, P3_U6045, P3_U6046, P3_U6047, P3_U6048, R152_U10, R152_U100, R152_U101, R152_U102, R152_U103, R152_U104, R152_U105, R152_U106, R152_U107, R152_U108, R152_U109, R152_U11, R152_U110, R152_U111, R152_U112, R152_U113, R152_U114, R152_U115, R152_U116, R152_U117, R152_U118, R152_U119, R152_U12, R152_U120, R152_U121, R152_U122, R152_U123, R152_U124, R152_U125, R152_U126, R152_U127, R152_U128, R152_U129, R152_U13, R152_U130, R152_U131, R152_U132, R152_U133, R152_U134, R152_U135, R152_U136, R152_U137, R152_U138, R152_U139, R152_U14, R152_U140, R152_U141, R152_U142, R152_U143, R152_U144, R152_U145, R152_U146, R152_U147, R152_U148, R152_U149, R152_U15, R152_U150, R152_U151, R152_U152, R152_U153, R152_U154, R152_U155, R152_U156, R152_U157, R152_U158, R152_U159, R152_U16, R152_U160, R152_U161, R152_U162, R152_U163, R152_U164, R152_U165, R152_U166, R152_U167, R152_U168, R152_U169, R152_U17, R152_U170, R152_U171, R152_U172, R152_U173, R152_U174, R152_U175, R152_U176, R152_U177, R152_U178, R152_U179, R152_U18, R152_U180, R152_U181, R152_U182, R152_U183, R152_U184, R152_U185, R152_U186, R152_U187, R152_U188, R152_U189, R152_U19, R152_U190, R152_U191, R152_U192, R152_U193, R152_U194, R152_U195, R152_U196, R152_U197, R152_U198, R152_U199, R152_U20, R152_U200, R152_U201, R152_U202, R152_U203, R152_U204, R152_U205, R152_U206, R152_U207, R152_U208, R152_U209, R152_U21, R152_U210, R152_U211, R152_U212, R152_U213, R152_U214, R152_U215, R152_U216, R152_U217, R152_U218, R152_U219, R152_U22, R152_U220, R152_U221, R152_U222, R152_U223, R152_U224, R152_U225, R152_U226, R152_U227, R152_U228, R152_U229, R152_U23, R152_U230, R152_U231, R152_U232, R152_U233, R152_U234, R152_U235, R152_U236, R152_U237, R152_U238, R152_U239, R152_U24, R152_U240, R152_U241, R152_U242, R152_U243, R152_U244, R152_U245, R152_U246, R152_U247, R152_U248, R152_U249, R152_U25, R152_U250, R152_U251, R152_U252, R152_U253, R152_U254, R152_U255, R152_U256, R152_U257, R152_U258, R152_U259, R152_U26, R152_U260, R152_U261, R152_U262, R152_U263, R152_U264, R152_U265, R152_U266, R152_U267, R152_U268, R152_U269, R152_U27, R152_U270, R152_U271, R152_U272, R152_U273, R152_U274, R152_U275, R152_U276, R152_U277, R152_U278, R152_U279, R152_U28, R152_U280, R152_U281, R152_U282, R152_U283, R152_U284, R152_U285, R152_U286, R152_U287, R152_U288, R152_U289, R152_U29, R152_U290, R152_U291, R152_U292, R152_U293, R152_U294, R152_U295, R152_U296, R152_U297, R152_U298, R152_U299, R152_U30, R152_U300, R152_U301, R152_U302, R152_U303, R152_U304, R152_U305, R152_U306, R152_U307, R152_U308, R152_U309, R152_U31, R152_U310, R152_U311, R152_U312, R152_U313, R152_U314, R152_U315, R152_U316, R152_U317, R152_U318, R152_U319, R152_U32, R152_U320, R152_U321, R152_U322, R152_U323, R152_U324, R152_U325, R152_U326, R152_U327, R152_U328, R152_U329, R152_U33, R152_U330, R152_U331, R152_U332, R152_U333, R152_U334, R152_U335, R152_U336, R152_U337, R152_U338, R152_U339, R152_U34, R152_U340, R152_U341, R152_U342, R152_U343, R152_U344, R152_U345, R152_U346, R152_U347, R152_U348, R152_U349, R152_U35, R152_U350, R152_U351, R152_U352, R152_U353, R152_U354, R152_U355, R152_U356, R152_U357, R152_U358, R152_U359, R152_U36, R152_U360, R152_U361, R152_U362, R152_U363, R152_U364, R152_U365, R152_U366, R152_U367, R152_U368, R152_U369, R152_U37, R152_U370, R152_U371, R152_U372, R152_U373, R152_U374, R152_U375, R152_U376, R152_U377, R152_U378, R152_U379, R152_U38, R152_U380, R152_U381, R152_U382, R152_U383, R152_U384, R152_U385, R152_U386, R152_U387, R152_U388, R152_U389, R152_U39, R152_U390, R152_U391, R152_U392, R152_U393, R152_U394, R152_U395, R152_U396, R152_U397, R152_U398, R152_U399, R152_U4, R152_U40, R152_U400, R152_U401, R152_U402, R152_U403, R152_U404, R152_U405, R152_U406, R152_U407, R152_U408, R152_U409, R152_U41, R152_U410, R152_U411, R152_U412, R152_U413, R152_U414, R152_U415, R152_U416, R152_U417, R152_U418, R152_U419, R152_U42, R152_U420, R152_U421, R152_U422, R152_U423, R152_U424, R152_U425, R152_U426, R152_U427, R152_U428, R152_U429, R152_U43, R152_U430, R152_U431, R152_U432, R152_U433, R152_U434, R152_U435, R152_U436, R152_U437, R152_U438, R152_U439, R152_U44, R152_U440, R152_U441, R152_U442, R152_U443, R152_U444, R152_U445, R152_U446, R152_U447, R152_U448, R152_U449, R152_U45, R152_U450, R152_U451, R152_U452, R152_U453, R152_U454, R152_U455, R152_U456, R152_U457, R152_U458, R152_U459, R152_U46, R152_U460, R152_U461, R152_U462, R152_U463, R152_U464, R152_U465, R152_U466, R152_U467, R152_U468, R152_U469, R152_U47, R152_U470, R152_U471, R152_U472, R152_U473, R152_U474, R152_U475, R152_U476, R152_U477, R152_U478, R152_U479, R152_U48, R152_U480, R152_U481, R152_U482, R152_U483, R152_U484, R152_U485, R152_U486, R152_U487, R152_U488, R152_U489, R152_U49, R152_U490, R152_U491, R152_U492, R152_U493, R152_U494, R152_U495, R152_U496, R152_U497, R152_U498, R152_U499, R152_U5, R152_U50, R152_U500, R152_U501, R152_U502, R152_U503, R152_U504, R152_U505, R152_U506, R152_U507, R152_U508, R152_U509, R152_U51, R152_U510, R152_U511, R152_U512, R152_U513, R152_U514, R152_U515, R152_U516, R152_U517, R152_U518, R152_U519, R152_U52, R152_U520, R152_U521, R152_U522, R152_U523, R152_U524, R152_U525, R152_U526, R152_U527, R152_U528, R152_U529, R152_U53, R152_U530, R152_U531, R152_U532, R152_U533, R152_U534, R152_U535, R152_U536, R152_U537, R152_U538, R152_U539, R152_U54, R152_U540, R152_U541, R152_U542, R152_U543, R152_U544, R152_U545, R152_U546, R152_U547, R152_U548, R152_U549, R152_U55, R152_U550, R152_U551, R152_U552, R152_U553, R152_U554, R152_U56, R152_U57, R152_U58, R152_U59, R152_U6, R152_U60, R152_U61, R152_U62, R152_U63, R152_U64, R152_U65, R152_U66, R152_U67, R152_U68, R152_U69, R152_U7, R152_U70, R152_U71, R152_U72, R152_U73, R152_U74, R152_U75, R152_U76, R152_U77, R152_U78, R152_U79, R152_U8, R152_U80, R152_U81, R152_U82, R152_U83, R152_U84, R152_U85, R152_U86, R152_U87, R152_U88, R152_U89, R152_U9, R152_U90, R152_U91, R152_U92, R152_U93, R152_U94, R152_U95, R152_U96, R152_U97, R152_U98, R152_U99, SUB_1596_U10, SUB_1596_U100, SUB_1596_U101, SUB_1596_U102, SUB_1596_U103, SUB_1596_U104, SUB_1596_U105, SUB_1596_U106, SUB_1596_U107, SUB_1596_U108, SUB_1596_U109, SUB_1596_U11, SUB_1596_U110, SUB_1596_U111, SUB_1596_U112, SUB_1596_U113, SUB_1596_U114, SUB_1596_U115, SUB_1596_U116, SUB_1596_U117, SUB_1596_U118, SUB_1596_U119, SUB_1596_U12, SUB_1596_U120, SUB_1596_U121, SUB_1596_U122, SUB_1596_U123, SUB_1596_U124, SUB_1596_U125, SUB_1596_U126, SUB_1596_U127, SUB_1596_U128, SUB_1596_U129, SUB_1596_U13, SUB_1596_U130, SUB_1596_U131, SUB_1596_U132, SUB_1596_U133, SUB_1596_U134, SUB_1596_U135, SUB_1596_U136, SUB_1596_U137, SUB_1596_U138, SUB_1596_U139, SUB_1596_U14, SUB_1596_U140, SUB_1596_U141, SUB_1596_U142, SUB_1596_U143, SUB_1596_U144, SUB_1596_U145, SUB_1596_U146, SUB_1596_U147, SUB_1596_U148, SUB_1596_U149, SUB_1596_U15, SUB_1596_U150, SUB_1596_U151, SUB_1596_U152, SUB_1596_U153, SUB_1596_U154, SUB_1596_U155, SUB_1596_U156, SUB_1596_U157, SUB_1596_U158, SUB_1596_U159, SUB_1596_U16, SUB_1596_U160, SUB_1596_U161, SUB_1596_U162, SUB_1596_U163, SUB_1596_U164, SUB_1596_U165, SUB_1596_U166, SUB_1596_U167, SUB_1596_U168, SUB_1596_U169, SUB_1596_U17, SUB_1596_U170, SUB_1596_U171, SUB_1596_U172, SUB_1596_U173, SUB_1596_U174, SUB_1596_U175, SUB_1596_U176, SUB_1596_U177, SUB_1596_U178, SUB_1596_U179, SUB_1596_U18, SUB_1596_U180, SUB_1596_U181, SUB_1596_U182, SUB_1596_U183, SUB_1596_U184, SUB_1596_U185, SUB_1596_U186, SUB_1596_U187, SUB_1596_U188, SUB_1596_U189, SUB_1596_U19, SUB_1596_U190, SUB_1596_U191, SUB_1596_U192, SUB_1596_U193, SUB_1596_U194, SUB_1596_U195, SUB_1596_U196, SUB_1596_U197, SUB_1596_U198, SUB_1596_U199, SUB_1596_U20, SUB_1596_U200, SUB_1596_U201, SUB_1596_U202, SUB_1596_U203, SUB_1596_U204, SUB_1596_U205, SUB_1596_U206, SUB_1596_U207, SUB_1596_U208, SUB_1596_U209, SUB_1596_U21, SUB_1596_U210, SUB_1596_U211, SUB_1596_U212, SUB_1596_U213, SUB_1596_U214, SUB_1596_U215, SUB_1596_U216, SUB_1596_U217, SUB_1596_U218, SUB_1596_U219, SUB_1596_U22, SUB_1596_U220, SUB_1596_U221, SUB_1596_U222, SUB_1596_U223, SUB_1596_U224, SUB_1596_U225, SUB_1596_U226, SUB_1596_U227, SUB_1596_U228, SUB_1596_U229, SUB_1596_U23, SUB_1596_U230, SUB_1596_U231, SUB_1596_U232, SUB_1596_U233, SUB_1596_U234, SUB_1596_U235, SUB_1596_U236, SUB_1596_U237, SUB_1596_U238, SUB_1596_U239, SUB_1596_U24, SUB_1596_U240, SUB_1596_U241, SUB_1596_U242, SUB_1596_U243, SUB_1596_U244, SUB_1596_U245, SUB_1596_U246, SUB_1596_U247, SUB_1596_U248, SUB_1596_U249, SUB_1596_U25, SUB_1596_U250, SUB_1596_U251, SUB_1596_U252, SUB_1596_U253, SUB_1596_U254, SUB_1596_U255, SUB_1596_U256, SUB_1596_U257, SUB_1596_U258, SUB_1596_U259, SUB_1596_U26, SUB_1596_U260, SUB_1596_U261, SUB_1596_U262, SUB_1596_U263, SUB_1596_U264, SUB_1596_U265, SUB_1596_U266, SUB_1596_U267, SUB_1596_U268, SUB_1596_U269, SUB_1596_U27, SUB_1596_U270, SUB_1596_U271, SUB_1596_U272, SUB_1596_U273, SUB_1596_U274, SUB_1596_U275, SUB_1596_U276, SUB_1596_U277, SUB_1596_U278, SUB_1596_U279, SUB_1596_U28, SUB_1596_U280, SUB_1596_U281, SUB_1596_U282, SUB_1596_U283, SUB_1596_U284, SUB_1596_U285, SUB_1596_U286, SUB_1596_U287, SUB_1596_U288, SUB_1596_U289, SUB_1596_U29, SUB_1596_U290, SUB_1596_U291, SUB_1596_U30, SUB_1596_U31, SUB_1596_U32, SUB_1596_U33, SUB_1596_U34, SUB_1596_U35, SUB_1596_U36, SUB_1596_U37, SUB_1596_U38, SUB_1596_U39, SUB_1596_U40, SUB_1596_U41, SUB_1596_U42, SUB_1596_U43, SUB_1596_U44, SUB_1596_U45, SUB_1596_U46, SUB_1596_U47, SUB_1596_U48, SUB_1596_U49, SUB_1596_U50, SUB_1596_U51, SUB_1596_U52, SUB_1596_U6, SUB_1596_U7, SUB_1596_U71, SUB_1596_U72, SUB_1596_U73, SUB_1596_U74, SUB_1596_U75, SUB_1596_U76, SUB_1596_U77, SUB_1596_U78, SUB_1596_U79, SUB_1596_U8, SUB_1596_U80, SUB_1596_U81, SUB_1596_U82, SUB_1596_U83, SUB_1596_U84, SUB_1596_U85, SUB_1596_U86, SUB_1596_U87, SUB_1596_U88, SUB_1596_U89, SUB_1596_U9, SUB_1596_U90, SUB_1596_U91, SUB_1596_U92, SUB_1596_U93, SUB_1596_U94, SUB_1596_U95, SUB_1596_U96, SUB_1596_U97, SUB_1596_U98, SUB_1596_U99, SUB_1605_U10, SUB_1605_U100, SUB_1605_U101, SUB_1605_U102, SUB_1605_U103, SUB_1605_U104, SUB_1605_U105, SUB_1605_U106, SUB_1605_U107, SUB_1605_U108, SUB_1605_U109, SUB_1605_U11, SUB_1605_U110, SUB_1605_U111, SUB_1605_U112, SUB_1605_U113, SUB_1605_U114, SUB_1605_U115, SUB_1605_U116, SUB_1605_U117, SUB_1605_U118, SUB_1605_U119, SUB_1605_U12, SUB_1605_U120, SUB_1605_U121, SUB_1605_U122, SUB_1605_U123, SUB_1605_U124, SUB_1605_U125, SUB_1605_U126, SUB_1605_U127, SUB_1605_U128, SUB_1605_U129, SUB_1605_U13, SUB_1605_U130, SUB_1605_U131, SUB_1605_U132, SUB_1605_U133, SUB_1605_U134, SUB_1605_U135, SUB_1605_U136, SUB_1605_U137, SUB_1605_U138, SUB_1605_U139, SUB_1605_U14, SUB_1605_U140, SUB_1605_U141, SUB_1605_U142, SUB_1605_U143, SUB_1605_U144, SUB_1605_U145, SUB_1605_U146, SUB_1605_U147, SUB_1605_U148, SUB_1605_U149, SUB_1605_U15, SUB_1605_U150, SUB_1605_U151, SUB_1605_U152, SUB_1605_U153, SUB_1605_U154, SUB_1605_U155, SUB_1605_U156, SUB_1605_U157, SUB_1605_U158, SUB_1605_U159, SUB_1605_U16, SUB_1605_U160, SUB_1605_U161, SUB_1605_U162, SUB_1605_U163, SUB_1605_U164, SUB_1605_U165, SUB_1605_U166, SUB_1605_U167, SUB_1605_U168, SUB_1605_U169, SUB_1605_U17, SUB_1605_U170, SUB_1605_U171, SUB_1605_U172, SUB_1605_U173, SUB_1605_U174, SUB_1605_U175, SUB_1605_U176, SUB_1605_U177, SUB_1605_U178, SUB_1605_U179, SUB_1605_U18, SUB_1605_U180, SUB_1605_U181, SUB_1605_U182, SUB_1605_U183, SUB_1605_U184, SUB_1605_U185, SUB_1605_U186, SUB_1605_U187, SUB_1605_U188, SUB_1605_U189, SUB_1605_U19, SUB_1605_U190, SUB_1605_U191, SUB_1605_U192, SUB_1605_U193, SUB_1605_U194, SUB_1605_U195, SUB_1605_U196, SUB_1605_U197, SUB_1605_U198, SUB_1605_U199, SUB_1605_U20, SUB_1605_U200, SUB_1605_U201, SUB_1605_U202, SUB_1605_U203, SUB_1605_U204, SUB_1605_U205, SUB_1605_U206, SUB_1605_U207, SUB_1605_U208, SUB_1605_U209, SUB_1605_U21, SUB_1605_U210, SUB_1605_U211, SUB_1605_U212, SUB_1605_U213, SUB_1605_U214, SUB_1605_U215, SUB_1605_U216, SUB_1605_U217, SUB_1605_U218, SUB_1605_U219, SUB_1605_U22, SUB_1605_U220, SUB_1605_U221, SUB_1605_U222, SUB_1605_U223, SUB_1605_U224, SUB_1605_U225, SUB_1605_U226, SUB_1605_U227, SUB_1605_U228, SUB_1605_U229, SUB_1605_U23, SUB_1605_U230, SUB_1605_U231, SUB_1605_U232, SUB_1605_U233, SUB_1605_U234, SUB_1605_U235, SUB_1605_U236, SUB_1605_U237, SUB_1605_U238, SUB_1605_U239, SUB_1605_U24, SUB_1605_U240, SUB_1605_U241, SUB_1605_U242, SUB_1605_U243, SUB_1605_U244, SUB_1605_U245, SUB_1605_U246, SUB_1605_U247, SUB_1605_U248, SUB_1605_U249, SUB_1605_U25, SUB_1605_U250, SUB_1605_U251, SUB_1605_U252, SUB_1605_U253, SUB_1605_U254, SUB_1605_U255, SUB_1605_U256, SUB_1605_U257, SUB_1605_U258, SUB_1605_U259, SUB_1605_U26, SUB_1605_U260, SUB_1605_U261, SUB_1605_U262, SUB_1605_U263, SUB_1605_U264, SUB_1605_U265, SUB_1605_U266, SUB_1605_U267, SUB_1605_U268, SUB_1605_U269, SUB_1605_U27, SUB_1605_U270, SUB_1605_U271, SUB_1605_U272, SUB_1605_U273, SUB_1605_U274, SUB_1605_U275, SUB_1605_U276, SUB_1605_U277, SUB_1605_U278, SUB_1605_U279, SUB_1605_U28, SUB_1605_U280, SUB_1605_U281, SUB_1605_U282, SUB_1605_U283, SUB_1605_U284, SUB_1605_U285, SUB_1605_U286, SUB_1605_U287, SUB_1605_U288, SUB_1605_U289, SUB_1605_U29, SUB_1605_U290, SUB_1605_U291, SUB_1605_U292, SUB_1605_U293, SUB_1605_U294, SUB_1605_U295, SUB_1605_U296, SUB_1605_U297, SUB_1605_U298, SUB_1605_U299, SUB_1605_U30, SUB_1605_U300, SUB_1605_U301, SUB_1605_U302, SUB_1605_U303, SUB_1605_U304, SUB_1605_U305, SUB_1605_U306, SUB_1605_U307, SUB_1605_U308, SUB_1605_U309, SUB_1605_U31, SUB_1605_U310, SUB_1605_U311, SUB_1605_U312, SUB_1605_U313, SUB_1605_U314, SUB_1605_U315, SUB_1605_U316, SUB_1605_U317, SUB_1605_U318, SUB_1605_U319, SUB_1605_U32, SUB_1605_U320, SUB_1605_U321, SUB_1605_U322, SUB_1605_U323, SUB_1605_U324, SUB_1605_U325, SUB_1605_U326, SUB_1605_U327, SUB_1605_U328, SUB_1605_U329, SUB_1605_U33, SUB_1605_U330, SUB_1605_U331, SUB_1605_U332, SUB_1605_U333, SUB_1605_U334, SUB_1605_U335, SUB_1605_U336, SUB_1605_U337, SUB_1605_U338, SUB_1605_U339, SUB_1605_U34, SUB_1605_U340, SUB_1605_U341, SUB_1605_U342, SUB_1605_U343, SUB_1605_U344, SUB_1605_U345, SUB_1605_U346, SUB_1605_U347, SUB_1605_U348, SUB_1605_U349, SUB_1605_U35, SUB_1605_U350, SUB_1605_U351, SUB_1605_U352, SUB_1605_U353, SUB_1605_U354, SUB_1605_U355, SUB_1605_U356, SUB_1605_U357, SUB_1605_U358, SUB_1605_U359, SUB_1605_U36, SUB_1605_U360, SUB_1605_U361, SUB_1605_U362, SUB_1605_U363, SUB_1605_U364, SUB_1605_U365, SUB_1605_U366, SUB_1605_U367, SUB_1605_U368, SUB_1605_U369, SUB_1605_U37, SUB_1605_U370, SUB_1605_U371, SUB_1605_U372, SUB_1605_U373, SUB_1605_U374, SUB_1605_U375, SUB_1605_U376, SUB_1605_U377, SUB_1605_U378, SUB_1605_U379, SUB_1605_U38, SUB_1605_U380, SUB_1605_U381, SUB_1605_U382, SUB_1605_U383, SUB_1605_U384, SUB_1605_U385, SUB_1605_U386, SUB_1605_U387, SUB_1605_U388, SUB_1605_U389, SUB_1605_U39, SUB_1605_U390, SUB_1605_U391, SUB_1605_U392, SUB_1605_U393, SUB_1605_U394, SUB_1605_U395, SUB_1605_U396, SUB_1605_U397, SUB_1605_U398, SUB_1605_U399, SUB_1605_U40, SUB_1605_U400, SUB_1605_U401, SUB_1605_U402, SUB_1605_U403, SUB_1605_U404, SUB_1605_U405, SUB_1605_U406, SUB_1605_U407, SUB_1605_U408, SUB_1605_U409, SUB_1605_U41, SUB_1605_U410, SUB_1605_U411, SUB_1605_U412, SUB_1605_U413, SUB_1605_U414, SUB_1605_U415, SUB_1605_U416, SUB_1605_U417, SUB_1605_U418, SUB_1605_U419, SUB_1605_U42, SUB_1605_U420, SUB_1605_U421, SUB_1605_U422, SUB_1605_U423, SUB_1605_U424, SUB_1605_U425, SUB_1605_U426, SUB_1605_U427, SUB_1605_U428, SUB_1605_U429, SUB_1605_U43, SUB_1605_U430, SUB_1605_U431, SUB_1605_U432, SUB_1605_U433, SUB_1605_U434, SUB_1605_U435, SUB_1605_U436, SUB_1605_U437, SUB_1605_U438, SUB_1605_U439, SUB_1605_U44, SUB_1605_U440, SUB_1605_U441, SUB_1605_U442, SUB_1605_U443, SUB_1605_U444, SUB_1605_U445, SUB_1605_U446, SUB_1605_U447, SUB_1605_U448, SUB_1605_U449, SUB_1605_U45, SUB_1605_U450, SUB_1605_U451, SUB_1605_U452, SUB_1605_U453, SUB_1605_U454, SUB_1605_U455, SUB_1605_U456, SUB_1605_U457, SUB_1605_U458, SUB_1605_U459, SUB_1605_U46, SUB_1605_U460, SUB_1605_U461, SUB_1605_U462, SUB_1605_U463, SUB_1605_U464, SUB_1605_U465, SUB_1605_U466, SUB_1605_U467, SUB_1605_U468, SUB_1605_U469, SUB_1605_U47, SUB_1605_U470, SUB_1605_U471, SUB_1605_U472, SUB_1605_U473, SUB_1605_U474, SUB_1605_U475, SUB_1605_U476, SUB_1605_U477, SUB_1605_U478, SUB_1605_U479, SUB_1605_U48, SUB_1605_U480, SUB_1605_U49, SUB_1605_U50, SUB_1605_U51, SUB_1605_U52, SUB_1605_U53, SUB_1605_U54, SUB_1605_U55, SUB_1605_U56, SUB_1605_U57, SUB_1605_U58, SUB_1605_U59, SUB_1605_U6, SUB_1605_U60, SUB_1605_U61, SUB_1605_U62, SUB_1605_U63, SUB_1605_U64, SUB_1605_U65, SUB_1605_U66, SUB_1605_U67, SUB_1605_U68, SUB_1605_U69, SUB_1605_U7, SUB_1605_U70, SUB_1605_U71, SUB_1605_U72, SUB_1605_U73, SUB_1605_U74, SUB_1605_U75, SUB_1605_U76, SUB_1605_U77, SUB_1605_U78, SUB_1605_U79, SUB_1605_U8, SUB_1605_U80, SUB_1605_U81, SUB_1605_U82, SUB_1605_U83, SUB_1605_U84, SUB_1605_U85, SUB_1605_U86, SUB_1605_U87, SUB_1605_U88, SUB_1605_U89, SUB_1605_U9, SUB_1605_U90, SUB_1605_U91, SUB_1605_U92, SUB_1605_U93, SUB_1605_U94, SUB_1605_U95, SUB_1605_U96, SUB_1605_U97, SUB_1605_U98, SUB_1605_U99, U100, U101, U102, U103, U104, U105, U106, U107, U108, U109, U110, U111, U112, U113, U114, U115, U116, U117, U118, U119, U120, U121, U122, U123, U124, U125, U126, U127, U128, U129, U130, U131, U132, U133, U134, U135, U136, U137, U138, U139, U140, U141, U142, U143, U144, U145, U146, U147, U148, U149, U150, U151, U152, U153, U154, U155, U156, U157, U158, U159, U160, U161, U162, U163, U164, U165, U166, U167, U168, U169, U170, U171, U172, U173, U174, U175, U176, U177, U178, U179, U180, U181, U182, U183, U184, U185, U186, U187, U188, U189, U190, U191, U192, U193, U194, U195, U196, U197, U198, U199, U200, U201, U202, U203, U204, U205, U206, U207, U208, U209, U210, U211, U212, U213, U214, U215, U216, U217, U218, U219, U220, U221, U222, U223, U224, U225, U226, U227, U228, U229, U230, U231, U232, U233, U234, U235, U236, U237, U238, U239, U240, U241, U242, U243, U244, U245, U246, U247, U248, U249, U250, U251, U252, U253, U254, U255, U256, U257, U258, U259, U260, U261, U262, U263, U264, U265, U266, U267, U268, U269, U270, U271, U272, U273, U274, U275, U276, U277, U278, U279, U280, U281, U282, U283, U284, U285, U286, U287, U288, U289, U290, U291, U292, U293, U294, U295, U296, U297, U298, U299, U30, U300, U301, U302, U303, U304, U305, U306, U307, U308, U309, U31, U310, U311, U312, U313, U314, U315, U316, U317, U318, U319, U32, U320, U321, U322, U323, U324, U325, U326, U327, U328, U329, U33, U330, U331, U332, U333, U334, U335, U336, U337, U338, U339, U34, U340, U341, U342, U343, U344, U345, U346, U347, U348, U349, U35, U350, U351, U352, U353, U354, U355, U356, U357, U358, U359, U36, U360, U361, U362, U363, U364, U365, U366, U367, U368, U369, U37, U370, U371, U372, U373, U374, U375, U376, U377, U378, U379, U38, U380, U381, U382, U383, U384, U385, U386, U387, U388, U389, U39, U390, U391, U392, U393, U394, U395, U396, U397, U398, U399, U40, U400, U401, U402, U403, U404, U405, U406, U407, U408, U409, U41, U410, U411, U412, U413, U414, U415, U416, U417, U418, U419, U42, U420, U421, U422, U423, U424, U425, U426, U427, U43, U44, U45, U46, U47, U48, U49, U50, U51, U52, U53, U54, U55, U56, U57, U58, U59, U60, U61, U62, U63, U64, U65, U66, U67, U68, U69, U70, U71, U72, U73, U74, U75, U76, U77, U78, U79, U80, U81, U82, U83, U84, U85, U86, U87, U88, U89, U90, U91, U92, U93, U94, U95, U96, U97, U98, U99, P2_U3520_in;

  not ginst1 (ADD_1596_U10, P1_ADDR_REG_1__SCAN_IN);
  nand ginst2 (ADD_1596_U100, ADD_1596_U140, ADD_1596_U141);
  nand ginst3 (ADD_1596_U101, ADD_1596_U136, ADD_1596_U137);
  not ginst4 (ADD_1596_U102, ADD_1596_U9);
  nand ginst5 (ADD_1596_U103, ADD_1596_U10, ADD_1596_U102);
  nand ginst6 (ADD_1596_U104, ADD_1596_U103, ADD_1596_U91);
  nand ginst7 (ADD_1596_U105, P1_ADDR_REG_1__SCAN_IN, ADD_1596_U9);
  not ginst8 (ADD_1596_U106, ADD_1596_U90);
  nand ginst9 (ADD_1596_U107, P3_ADDR_REG_2__SCAN_IN, ADD_1596_U12);
  nand ginst10 (ADD_1596_U108, ADD_1596_U107, ADD_1596_U90);
  nand ginst11 (ADD_1596_U109, P1_ADDR_REG_2__SCAN_IN, ADD_1596_U11);
  not ginst12 (ADD_1596_U11, P3_ADDR_REG_2__SCAN_IN);
  not ginst13 (ADD_1596_U110, ADD_1596_U89);
  nand ginst14 (ADD_1596_U111, P3_ADDR_REG_3__SCAN_IN, ADD_1596_U14);
  nand ginst15 (ADD_1596_U112, ADD_1596_U111, ADD_1596_U89);
  nand ginst16 (ADD_1596_U113, P1_ADDR_REG_3__SCAN_IN, ADD_1596_U13);
  not ginst17 (ADD_1596_U114, ADD_1596_U88);
  nand ginst18 (ADD_1596_U115, P3_ADDR_REG_4__SCAN_IN, ADD_1596_U16);
  nand ginst19 (ADD_1596_U116, ADD_1596_U115, ADD_1596_U88);
  nand ginst20 (ADD_1596_U117, P1_ADDR_REG_4__SCAN_IN, ADD_1596_U15);
  not ginst21 (ADD_1596_U118, ADD_1596_U87);
  nand ginst22 (ADD_1596_U119, P3_ADDR_REG_5__SCAN_IN, ADD_1596_U18);
  not ginst23 (ADD_1596_U12, P1_ADDR_REG_2__SCAN_IN);
  nand ginst24 (ADD_1596_U120, ADD_1596_U119, ADD_1596_U87);
  nand ginst25 (ADD_1596_U121, P1_ADDR_REG_5__SCAN_IN, ADD_1596_U17);
  not ginst26 (ADD_1596_U122, ADD_1596_U86);
  nand ginst27 (ADD_1596_U123, P3_ADDR_REG_6__SCAN_IN, ADD_1596_U20);
  nand ginst28 (ADD_1596_U124, ADD_1596_U123, ADD_1596_U86);
  nand ginst29 (ADD_1596_U125, P1_ADDR_REG_6__SCAN_IN, ADD_1596_U19);
  not ginst30 (ADD_1596_U126, ADD_1596_U85);
  nand ginst31 (ADD_1596_U127, P3_ADDR_REG_7__SCAN_IN, ADD_1596_U22);
  nand ginst32 (ADD_1596_U128, ADD_1596_U127, ADD_1596_U85);
  nand ginst33 (ADD_1596_U129, P1_ADDR_REG_7__SCAN_IN, ADD_1596_U21);
  not ginst34 (ADD_1596_U13, P3_ADDR_REG_3__SCAN_IN);
  not ginst35 (ADD_1596_U130, ADD_1596_U84);
  nand ginst36 (ADD_1596_U131, P3_ADDR_REG_8__SCAN_IN, ADD_1596_U24);
  nand ginst37 (ADD_1596_U132, ADD_1596_U131, ADD_1596_U84);
  nand ginst38 (ADD_1596_U133, P1_ADDR_REG_8__SCAN_IN, ADD_1596_U23);
  not ginst39 (ADD_1596_U134, ADD_1596_U83);
  nand ginst40 (ADD_1596_U135, P3_ADDR_REG_9__SCAN_IN, ADD_1596_U26);
  nand ginst41 (ADD_1596_U136, ADD_1596_U135, ADD_1596_U83);
  nand ginst42 (ADD_1596_U137, P1_ADDR_REG_9__SCAN_IN, ADD_1596_U25);
  not ginst43 (ADD_1596_U138, ADD_1596_U101);
  nand ginst44 (ADD_1596_U139, P3_ADDR_REG_10__SCAN_IN, ADD_1596_U28);
  not ginst45 (ADD_1596_U14, P1_ADDR_REG_3__SCAN_IN);
  nand ginst46 (ADD_1596_U140, ADD_1596_U101, ADD_1596_U139);
  nand ginst47 (ADD_1596_U141, P1_ADDR_REG_10__SCAN_IN, ADD_1596_U27);
  not ginst48 (ADD_1596_U142, ADD_1596_U100);
  nand ginst49 (ADD_1596_U143, P3_ADDR_REG_11__SCAN_IN, ADD_1596_U30);
  nand ginst50 (ADD_1596_U144, ADD_1596_U100, ADD_1596_U143);
  nand ginst51 (ADD_1596_U145, P1_ADDR_REG_11__SCAN_IN, ADD_1596_U29);
  not ginst52 (ADD_1596_U146, ADD_1596_U99);
  nand ginst53 (ADD_1596_U147, P3_ADDR_REG_12__SCAN_IN, ADD_1596_U32);
  nand ginst54 (ADD_1596_U148, ADD_1596_U147, ADD_1596_U99);
  nand ginst55 (ADD_1596_U149, P1_ADDR_REG_12__SCAN_IN, ADD_1596_U31);
  not ginst56 (ADD_1596_U15, P3_ADDR_REG_4__SCAN_IN);
  not ginst57 (ADD_1596_U150, ADD_1596_U98);
  nand ginst58 (ADD_1596_U151, P3_ADDR_REG_13__SCAN_IN, ADD_1596_U34);
  nand ginst59 (ADD_1596_U152, ADD_1596_U151, ADD_1596_U98);
  nand ginst60 (ADD_1596_U153, P1_ADDR_REG_13__SCAN_IN, ADD_1596_U33);
  not ginst61 (ADD_1596_U154, ADD_1596_U97);
  nand ginst62 (ADD_1596_U155, P3_ADDR_REG_14__SCAN_IN, ADD_1596_U36);
  nand ginst63 (ADD_1596_U156, ADD_1596_U155, ADD_1596_U97);
  nand ginst64 (ADD_1596_U157, P1_ADDR_REG_14__SCAN_IN, ADD_1596_U35);
  not ginst65 (ADD_1596_U158, ADD_1596_U96);
  nand ginst66 (ADD_1596_U159, P3_ADDR_REG_15__SCAN_IN, ADD_1596_U38);
  not ginst67 (ADD_1596_U16, P1_ADDR_REG_4__SCAN_IN);
  nand ginst68 (ADD_1596_U160, ADD_1596_U159, ADD_1596_U96);
  nand ginst69 (ADD_1596_U161, P1_ADDR_REG_15__SCAN_IN, ADD_1596_U37);
  not ginst70 (ADD_1596_U162, ADD_1596_U95);
  nand ginst71 (ADD_1596_U163, P3_ADDR_REG_16__SCAN_IN, ADD_1596_U40);
  nand ginst72 (ADD_1596_U164, ADD_1596_U163, ADD_1596_U95);
  nand ginst73 (ADD_1596_U165, P1_ADDR_REG_16__SCAN_IN, ADD_1596_U39);
  not ginst74 (ADD_1596_U166, ADD_1596_U94);
  nand ginst75 (ADD_1596_U167, P3_ADDR_REG_17__SCAN_IN, ADD_1596_U42);
  nand ginst76 (ADD_1596_U168, ADD_1596_U167, ADD_1596_U94);
  nand ginst77 (ADD_1596_U169, P1_ADDR_REG_17__SCAN_IN, ADD_1596_U41);
  not ginst78 (ADD_1596_U17, P3_ADDR_REG_5__SCAN_IN);
  not ginst79 (ADD_1596_U170, ADD_1596_U45);
  nand ginst80 (ADD_1596_U171, P1_ADDR_REG_18__SCAN_IN, ADD_1596_U43);
  nand ginst81 (ADD_1596_U172, ADD_1596_U170, ADD_1596_U171);
  nand ginst82 (ADD_1596_U173, P3_ADDR_REG_18__SCAN_IN, ADD_1596_U44);
  nand ginst83 (ADD_1596_U174, ADD_1596_U172, ADD_1596_U173, ADD_1596_U229);
  nand ginst84 (ADD_1596_U175, P3_ADDR_REG_18__SCAN_IN, ADD_1596_U44);
  nand ginst85 (ADD_1596_U176, ADD_1596_U175, ADD_1596_U45);
  nand ginst86 (ADD_1596_U177, P1_ADDR_REG_18__SCAN_IN, ADD_1596_U43);
  nand ginst87 (ADD_1596_U178, ADD_1596_U176, ADD_1596_U177, ADD_1596_U225, ADD_1596_U226);
  nand ginst88 (ADD_1596_U179, P1_ADDR_REG_0__SCAN_IN, ADD_1596_U8);
  not ginst89 (ADD_1596_U18, P1_ADDR_REG_5__SCAN_IN);
  nand ginst90 (ADD_1596_U180, P3_ADDR_REG_9__SCAN_IN, ADD_1596_U26);
  nand ginst91 (ADD_1596_U181, P1_ADDR_REG_9__SCAN_IN, ADD_1596_U25);
  not ginst92 (ADD_1596_U182, ADD_1596_U65);
  nand ginst93 (ADD_1596_U183, ADD_1596_U134, ADD_1596_U182);
  nand ginst94 (ADD_1596_U184, ADD_1596_U65, ADD_1596_U83);
  nand ginst95 (ADD_1596_U185, P3_ADDR_REG_8__SCAN_IN, ADD_1596_U24);
  nand ginst96 (ADD_1596_U186, P1_ADDR_REG_8__SCAN_IN, ADD_1596_U23);
  not ginst97 (ADD_1596_U187, ADD_1596_U66);
  nand ginst98 (ADD_1596_U188, ADD_1596_U130, ADD_1596_U187);
  nand ginst99 (ADD_1596_U189, ADD_1596_U66, ADD_1596_U84);
  not ginst100 (ADD_1596_U19, P3_ADDR_REG_6__SCAN_IN);
  nand ginst101 (ADD_1596_U190, P3_ADDR_REG_7__SCAN_IN, ADD_1596_U22);
  nand ginst102 (ADD_1596_U191, P1_ADDR_REG_7__SCAN_IN, ADD_1596_U21);
  not ginst103 (ADD_1596_U192, ADD_1596_U67);
  nand ginst104 (ADD_1596_U193, ADD_1596_U126, ADD_1596_U192);
  nand ginst105 (ADD_1596_U194, ADD_1596_U67, ADD_1596_U85);
  nand ginst106 (ADD_1596_U195, P3_ADDR_REG_6__SCAN_IN, ADD_1596_U20);
  nand ginst107 (ADD_1596_U196, P1_ADDR_REG_6__SCAN_IN, ADD_1596_U19);
  not ginst108 (ADD_1596_U197, ADD_1596_U68);
  nand ginst109 (ADD_1596_U198, ADD_1596_U122, ADD_1596_U197);
  nand ginst110 (ADD_1596_U199, ADD_1596_U68, ADD_1596_U86);
  not ginst111 (ADD_1596_U20, P1_ADDR_REG_6__SCAN_IN);
  nand ginst112 (ADD_1596_U200, P3_ADDR_REG_5__SCAN_IN, ADD_1596_U18);
  nand ginst113 (ADD_1596_U201, P1_ADDR_REG_5__SCAN_IN, ADD_1596_U17);
  not ginst114 (ADD_1596_U202, ADD_1596_U69);
  nand ginst115 (ADD_1596_U203, ADD_1596_U118, ADD_1596_U202);
  nand ginst116 (ADD_1596_U204, ADD_1596_U69, ADD_1596_U87);
  nand ginst117 (ADD_1596_U205, P3_ADDR_REG_4__SCAN_IN, ADD_1596_U16);
  nand ginst118 (ADD_1596_U206, P1_ADDR_REG_4__SCAN_IN, ADD_1596_U15);
  not ginst119 (ADD_1596_U207, ADD_1596_U70);
  nand ginst120 (ADD_1596_U208, ADD_1596_U114, ADD_1596_U207);
  nand ginst121 (ADD_1596_U209, ADD_1596_U70, ADD_1596_U88);
  not ginst122 (ADD_1596_U21, P3_ADDR_REG_7__SCAN_IN);
  nand ginst123 (ADD_1596_U210, P3_ADDR_REG_3__SCAN_IN, ADD_1596_U14);
  nand ginst124 (ADD_1596_U211, P1_ADDR_REG_3__SCAN_IN, ADD_1596_U13);
  not ginst125 (ADD_1596_U212, ADD_1596_U71);
  nand ginst126 (ADD_1596_U213, ADD_1596_U110, ADD_1596_U212);
  nand ginst127 (ADD_1596_U214, ADD_1596_U71, ADD_1596_U89);
  nand ginst128 (ADD_1596_U215, P3_ADDR_REG_2__SCAN_IN, ADD_1596_U12);
  nand ginst129 (ADD_1596_U216, P1_ADDR_REG_2__SCAN_IN, ADD_1596_U11);
  not ginst130 (ADD_1596_U217, ADD_1596_U72);
  nand ginst131 (ADD_1596_U218, ADD_1596_U106, ADD_1596_U217);
  nand ginst132 (ADD_1596_U219, ADD_1596_U72, ADD_1596_U90);
  not ginst133 (ADD_1596_U22, P1_ADDR_REG_7__SCAN_IN);
  nand ginst134 (ADD_1596_U220, P3_ADDR_REG_1__SCAN_IN, ADD_1596_U10);
  nand ginst135 (ADD_1596_U221, P1_ADDR_REG_1__SCAN_IN, ADD_1596_U91);
  not ginst136 (ADD_1596_U222, ADD_1596_U73);
  nand ginst137 (ADD_1596_U223, ADD_1596_U102, ADD_1596_U222);
  nand ginst138 (ADD_1596_U224, ADD_1596_U73, ADD_1596_U9);
  nand ginst139 (ADD_1596_U225, P3_ADDR_REG_19__SCAN_IN, ADD_1596_U93);
  nand ginst140 (ADD_1596_U226, P1_ADDR_REG_19__SCAN_IN, ADD_1596_U92);
  nand ginst141 (ADD_1596_U227, P3_ADDR_REG_19__SCAN_IN, ADD_1596_U93);
  nand ginst142 (ADD_1596_U228, P1_ADDR_REG_19__SCAN_IN, ADD_1596_U92);
  nand ginst143 (ADD_1596_U229, ADD_1596_U227, ADD_1596_U228);
  not ginst144 (ADD_1596_U23, P3_ADDR_REG_8__SCAN_IN);
  nand ginst145 (ADD_1596_U230, P3_ADDR_REG_18__SCAN_IN, ADD_1596_U44);
  nand ginst146 (ADD_1596_U231, P1_ADDR_REG_18__SCAN_IN, ADD_1596_U43);
  not ginst147 (ADD_1596_U232, ADD_1596_U74);
  nand ginst148 (ADD_1596_U233, ADD_1596_U170, ADD_1596_U232);
  nand ginst149 (ADD_1596_U234, ADD_1596_U45, ADD_1596_U74);
  nand ginst150 (ADD_1596_U235, P3_ADDR_REG_17__SCAN_IN, ADD_1596_U42);
  nand ginst151 (ADD_1596_U236, P1_ADDR_REG_17__SCAN_IN, ADD_1596_U41);
  not ginst152 (ADD_1596_U237, ADD_1596_U75);
  nand ginst153 (ADD_1596_U238, ADD_1596_U166, ADD_1596_U237);
  nand ginst154 (ADD_1596_U239, ADD_1596_U75, ADD_1596_U94);
  not ginst155 (ADD_1596_U24, P1_ADDR_REG_8__SCAN_IN);
  nand ginst156 (ADD_1596_U240, P3_ADDR_REG_16__SCAN_IN, ADD_1596_U40);
  nand ginst157 (ADD_1596_U241, P1_ADDR_REG_16__SCAN_IN, ADD_1596_U39);
  not ginst158 (ADD_1596_U242, ADD_1596_U76);
  nand ginst159 (ADD_1596_U243, ADD_1596_U162, ADD_1596_U242);
  nand ginst160 (ADD_1596_U244, ADD_1596_U76, ADD_1596_U95);
  nand ginst161 (ADD_1596_U245, P3_ADDR_REG_15__SCAN_IN, ADD_1596_U38);
  nand ginst162 (ADD_1596_U246, P1_ADDR_REG_15__SCAN_IN, ADD_1596_U37);
  not ginst163 (ADD_1596_U247, ADD_1596_U77);
  nand ginst164 (ADD_1596_U248, ADD_1596_U158, ADD_1596_U247);
  nand ginst165 (ADD_1596_U249, ADD_1596_U77, ADD_1596_U96);
  not ginst166 (ADD_1596_U25, P3_ADDR_REG_9__SCAN_IN);
  nand ginst167 (ADD_1596_U250, P3_ADDR_REG_14__SCAN_IN, ADD_1596_U36);
  nand ginst168 (ADD_1596_U251, P1_ADDR_REG_14__SCAN_IN, ADD_1596_U35);
  not ginst169 (ADD_1596_U252, ADD_1596_U78);
  nand ginst170 (ADD_1596_U253, ADD_1596_U154, ADD_1596_U252);
  nand ginst171 (ADD_1596_U254, ADD_1596_U78, ADD_1596_U97);
  nand ginst172 (ADD_1596_U255, P3_ADDR_REG_13__SCAN_IN, ADD_1596_U34);
  nand ginst173 (ADD_1596_U256, P1_ADDR_REG_13__SCAN_IN, ADD_1596_U33);
  not ginst174 (ADD_1596_U257, ADD_1596_U79);
  nand ginst175 (ADD_1596_U258, ADD_1596_U150, ADD_1596_U257);
  nand ginst176 (ADD_1596_U259, ADD_1596_U79, ADD_1596_U98);
  not ginst177 (ADD_1596_U26, P1_ADDR_REG_9__SCAN_IN);
  nand ginst178 (ADD_1596_U260, P3_ADDR_REG_12__SCAN_IN, ADD_1596_U32);
  nand ginst179 (ADD_1596_U261, P1_ADDR_REG_12__SCAN_IN, ADD_1596_U31);
  not ginst180 (ADD_1596_U262, ADD_1596_U80);
  nand ginst181 (ADD_1596_U263, ADD_1596_U146, ADD_1596_U262);
  nand ginst182 (ADD_1596_U264, ADD_1596_U80, ADD_1596_U99);
  nand ginst183 (ADD_1596_U265, P3_ADDR_REG_11__SCAN_IN, ADD_1596_U30);
  nand ginst184 (ADD_1596_U266, P1_ADDR_REG_11__SCAN_IN, ADD_1596_U29);
  not ginst185 (ADD_1596_U267, ADD_1596_U81);
  nand ginst186 (ADD_1596_U268, ADD_1596_U142, ADD_1596_U267);
  nand ginst187 (ADD_1596_U269, ADD_1596_U100, ADD_1596_U81);
  not ginst188 (ADD_1596_U27, P3_ADDR_REG_10__SCAN_IN);
  nand ginst189 (ADD_1596_U270, P3_ADDR_REG_10__SCAN_IN, ADD_1596_U28);
  nand ginst190 (ADD_1596_U271, P1_ADDR_REG_10__SCAN_IN, ADD_1596_U27);
  not ginst191 (ADD_1596_U272, ADD_1596_U82);
  nand ginst192 (ADD_1596_U273, ADD_1596_U138, ADD_1596_U272);
  nand ginst193 (ADD_1596_U274, ADD_1596_U101, ADD_1596_U82);
  not ginst194 (ADD_1596_U28, P1_ADDR_REG_10__SCAN_IN);
  not ginst195 (ADD_1596_U29, P3_ADDR_REG_11__SCAN_IN);
  not ginst196 (ADD_1596_U30, P1_ADDR_REG_11__SCAN_IN);
  not ginst197 (ADD_1596_U31, P3_ADDR_REG_12__SCAN_IN);
  not ginst198 (ADD_1596_U32, P1_ADDR_REG_12__SCAN_IN);
  not ginst199 (ADD_1596_U33, P3_ADDR_REG_13__SCAN_IN);
  not ginst200 (ADD_1596_U34, P1_ADDR_REG_13__SCAN_IN);
  not ginst201 (ADD_1596_U35, P3_ADDR_REG_14__SCAN_IN);
  not ginst202 (ADD_1596_U36, P1_ADDR_REG_14__SCAN_IN);
  not ginst203 (ADD_1596_U37, P3_ADDR_REG_15__SCAN_IN);
  not ginst204 (ADD_1596_U38, P1_ADDR_REG_15__SCAN_IN);
  not ginst205 (ADD_1596_U39, P3_ADDR_REG_16__SCAN_IN);
  not ginst206 (ADD_1596_U40, P1_ADDR_REG_16__SCAN_IN);
  not ginst207 (ADD_1596_U41, P3_ADDR_REG_17__SCAN_IN);
  not ginst208 (ADD_1596_U42, P1_ADDR_REG_17__SCAN_IN);
  not ginst209 (ADD_1596_U43, P3_ADDR_REG_18__SCAN_IN);
  not ginst210 (ADD_1596_U44, P1_ADDR_REG_18__SCAN_IN);
  nand ginst211 (ADD_1596_U45, ADD_1596_U168, ADD_1596_U169);
  not ginst212 (ADD_1596_U46, P1_ADDR_REG_0__SCAN_IN);
  nand ginst213 (ADD_1596_U47, ADD_1596_U183, ADD_1596_U184);
  nand ginst214 (ADD_1596_U48, ADD_1596_U188, ADD_1596_U189);
  nand ginst215 (ADD_1596_U49, ADD_1596_U193, ADD_1596_U194);
  nand ginst216 (ADD_1596_U50, ADD_1596_U198, ADD_1596_U199);
  nand ginst217 (ADD_1596_U51, ADD_1596_U203, ADD_1596_U204);
  nand ginst218 (ADD_1596_U52, ADD_1596_U208, ADD_1596_U209);
  nand ginst219 (ADD_1596_U53, ADD_1596_U213, ADD_1596_U214);
  nand ginst220 (ADD_1596_U54, ADD_1596_U218, ADD_1596_U219);
  nand ginst221 (ADD_1596_U55, ADD_1596_U223, ADD_1596_U224);
  nand ginst222 (ADD_1596_U56, ADD_1596_U233, ADD_1596_U234);
  nand ginst223 (ADD_1596_U57, ADD_1596_U238, ADD_1596_U239);
  nand ginst224 (ADD_1596_U58, ADD_1596_U243, ADD_1596_U244);
  nand ginst225 (ADD_1596_U59, ADD_1596_U248, ADD_1596_U249);
  nand ginst226 (ADD_1596_U6, ADD_1596_U174, ADD_1596_U178);
  nand ginst227 (ADD_1596_U60, ADD_1596_U253, ADD_1596_U254);
  nand ginst228 (ADD_1596_U61, ADD_1596_U258, ADD_1596_U259);
  nand ginst229 (ADD_1596_U62, ADD_1596_U263, ADD_1596_U264);
  nand ginst230 (ADD_1596_U63, ADD_1596_U268, ADD_1596_U269);
  nand ginst231 (ADD_1596_U64, ADD_1596_U273, ADD_1596_U274);
  nand ginst232 (ADD_1596_U65, ADD_1596_U180, ADD_1596_U181);
  nand ginst233 (ADD_1596_U66, ADD_1596_U185, ADD_1596_U186);
  nand ginst234 (ADD_1596_U67, ADD_1596_U190, ADD_1596_U191);
  nand ginst235 (ADD_1596_U68, ADD_1596_U195, ADD_1596_U196);
  nand ginst236 (ADD_1596_U69, ADD_1596_U200, ADD_1596_U201);
  nand ginst237 (ADD_1596_U7, ADD_1596_U179, ADD_1596_U9);
  nand ginst238 (ADD_1596_U70, ADD_1596_U205, ADD_1596_U206);
  nand ginst239 (ADD_1596_U71, ADD_1596_U210, ADD_1596_U211);
  nand ginst240 (ADD_1596_U72, ADD_1596_U215, ADD_1596_U216);
  nand ginst241 (ADD_1596_U73, ADD_1596_U220, ADD_1596_U221);
  nand ginst242 (ADD_1596_U74, ADD_1596_U230, ADD_1596_U231);
  nand ginst243 (ADD_1596_U75, ADD_1596_U235, ADD_1596_U236);
  nand ginst244 (ADD_1596_U76, ADD_1596_U240, ADD_1596_U241);
  nand ginst245 (ADD_1596_U77, ADD_1596_U245, ADD_1596_U246);
  nand ginst246 (ADD_1596_U78, ADD_1596_U250, ADD_1596_U251);
  nand ginst247 (ADD_1596_U79, ADD_1596_U255, ADD_1596_U256);
  not ginst248 (ADD_1596_U8, P3_ADDR_REG_0__SCAN_IN);
  nand ginst249 (ADD_1596_U80, ADD_1596_U260, ADD_1596_U261);
  nand ginst250 (ADD_1596_U81, ADD_1596_U265, ADD_1596_U266);
  nand ginst251 (ADD_1596_U82, ADD_1596_U270, ADD_1596_U271);
  nand ginst252 (ADD_1596_U83, ADD_1596_U132, ADD_1596_U133);
  nand ginst253 (ADD_1596_U84, ADD_1596_U128, ADD_1596_U129);
  nand ginst254 (ADD_1596_U85, ADD_1596_U124, ADD_1596_U125);
  nand ginst255 (ADD_1596_U86, ADD_1596_U120, ADD_1596_U121);
  nand ginst256 (ADD_1596_U87, ADD_1596_U116, ADD_1596_U117);
  nand ginst257 (ADD_1596_U88, ADD_1596_U112, ADD_1596_U113);
  nand ginst258 (ADD_1596_U89, ADD_1596_U108, ADD_1596_U109);
  nand ginst259 (ADD_1596_U9, P3_ADDR_REG_0__SCAN_IN, ADD_1596_U46);
  nand ginst260 (ADD_1596_U90, ADD_1596_U104, ADD_1596_U105);
  not ginst261 (ADD_1596_U91, P3_ADDR_REG_1__SCAN_IN);
  not ginst262 (ADD_1596_U92, P3_ADDR_REG_19__SCAN_IN);
  not ginst263 (ADD_1596_U93, P1_ADDR_REG_19__SCAN_IN);
  nand ginst264 (ADD_1596_U94, ADD_1596_U164, ADD_1596_U165);
  nand ginst265 (ADD_1596_U95, ADD_1596_U160, ADD_1596_U161);
  nand ginst266 (ADD_1596_U96, ADD_1596_U156, ADD_1596_U157);
  nand ginst267 (ADD_1596_U97, ADD_1596_U152, ADD_1596_U153);
  nand ginst268 (ADD_1596_U98, ADD_1596_U148, ADD_1596_U149);
  nand ginst269 (ADD_1596_U99, ADD_1596_U144, ADD_1596_U145);
  not ginst270 (LT_1601_21_U6, P2_ADDR_REG_19__SCAN_IN);
  not ginst271 (LT_1601_U6, P1_ADDR_REG_19__SCAN_IN);
  not ginst272 (LT_1602_U6, P3_ADDR_REG_19__SCAN_IN);
  not ginst273 (P1_ADD_99_U10, P1_REG3_REG_6__SCAN_IN);
  not ginst274 (P1_ADD_99_U100, P1_ADD_99_U47);
  not ginst275 (P1_ADD_99_U101, P1_ADD_99_U49);
  not ginst276 (P1_ADD_99_U102, P1_ADD_99_U51);
  not ginst277 (P1_ADD_99_U103, P1_ADD_99_U79);
  nand ginst278 (P1_ADD_99_U104, P1_REG3_REG_9__SCAN_IN, P1_ADD_99_U16);
  nand ginst279 (P1_ADD_99_U105, P1_ADD_99_U15, P1_ADD_99_U84);
  nand ginst280 (P1_ADD_99_U106, P1_REG3_REG_8__SCAN_IN, P1_ADD_99_U13);
  nand ginst281 (P1_ADD_99_U107, P1_ADD_99_U14, P1_ADD_99_U83);
  nand ginst282 (P1_ADD_99_U108, P1_REG3_REG_7__SCAN_IN, P1_ADD_99_U11);
  nand ginst283 (P1_ADD_99_U109, P1_ADD_99_U12, P1_ADD_99_U82);
  nand ginst284 (P1_ADD_99_U11, P1_REG3_REG_6__SCAN_IN, P1_ADD_99_U81);
  nand ginst285 (P1_ADD_99_U110, P1_REG3_REG_6__SCAN_IN, P1_ADD_99_U9);
  nand ginst286 (P1_ADD_99_U111, P1_ADD_99_U10, P1_ADD_99_U81);
  nand ginst287 (P1_ADD_99_U112, P1_REG3_REG_5__SCAN_IN, P1_ADD_99_U7);
  nand ginst288 (P1_ADD_99_U113, P1_ADD_99_U8, P1_ADD_99_U80);
  nand ginst289 (P1_ADD_99_U114, P1_REG3_REG_4__SCAN_IN, P1_ADD_99_U4);
  nand ginst290 (P1_ADD_99_U115, P1_REG3_REG_3__SCAN_IN, P1_ADD_99_U6);
  nand ginst291 (P1_ADD_99_U116, P1_REG3_REG_28__SCAN_IN, P1_ADD_99_U79);
  nand ginst292 (P1_ADD_99_U117, P1_ADD_99_U103, P1_ADD_99_U52);
  nand ginst293 (P1_ADD_99_U118, P1_REG3_REG_27__SCAN_IN, P1_ADD_99_U51);
  nand ginst294 (P1_ADD_99_U119, P1_ADD_99_U102, P1_ADD_99_U53);
  not ginst295 (P1_ADD_99_U12, P1_REG3_REG_7__SCAN_IN);
  nand ginst296 (P1_ADD_99_U120, P1_REG3_REG_26__SCAN_IN, P1_ADD_99_U49);
  nand ginst297 (P1_ADD_99_U121, P1_ADD_99_U101, P1_ADD_99_U50);
  nand ginst298 (P1_ADD_99_U122, P1_REG3_REG_25__SCAN_IN, P1_ADD_99_U47);
  nand ginst299 (P1_ADD_99_U123, P1_ADD_99_U100, P1_ADD_99_U48);
  nand ginst300 (P1_ADD_99_U124, P1_REG3_REG_24__SCAN_IN, P1_ADD_99_U45);
  nand ginst301 (P1_ADD_99_U125, P1_ADD_99_U46, P1_ADD_99_U99);
  nand ginst302 (P1_ADD_99_U126, P1_REG3_REG_23__SCAN_IN, P1_ADD_99_U43);
  nand ginst303 (P1_ADD_99_U127, P1_ADD_99_U44, P1_ADD_99_U98);
  nand ginst304 (P1_ADD_99_U128, P1_REG3_REG_22__SCAN_IN, P1_ADD_99_U41);
  nand ginst305 (P1_ADD_99_U129, P1_ADD_99_U42, P1_ADD_99_U97);
  nand ginst306 (P1_ADD_99_U13, P1_REG3_REG_7__SCAN_IN, P1_ADD_99_U82);
  nand ginst307 (P1_ADD_99_U130, P1_REG3_REG_21__SCAN_IN, P1_ADD_99_U39);
  nand ginst308 (P1_ADD_99_U131, P1_ADD_99_U40, P1_ADD_99_U96);
  nand ginst309 (P1_ADD_99_U132, P1_REG3_REG_20__SCAN_IN, P1_ADD_99_U37);
  nand ginst310 (P1_ADD_99_U133, P1_ADD_99_U38, P1_ADD_99_U95);
  nand ginst311 (P1_ADD_99_U134, P1_REG3_REG_19__SCAN_IN, P1_ADD_99_U35);
  nand ginst312 (P1_ADD_99_U135, P1_ADD_99_U36, P1_ADD_99_U94);
  nand ginst313 (P1_ADD_99_U136, P1_REG3_REG_18__SCAN_IN, P1_ADD_99_U33);
  nand ginst314 (P1_ADD_99_U137, P1_ADD_99_U34, P1_ADD_99_U93);
  nand ginst315 (P1_ADD_99_U138, P1_REG3_REG_17__SCAN_IN, P1_ADD_99_U31);
  nand ginst316 (P1_ADD_99_U139, P1_ADD_99_U32, P1_ADD_99_U92);
  not ginst317 (P1_ADD_99_U14, P1_REG3_REG_8__SCAN_IN);
  nand ginst318 (P1_ADD_99_U140, P1_REG3_REG_16__SCAN_IN, P1_ADD_99_U29);
  nand ginst319 (P1_ADD_99_U141, P1_ADD_99_U30, P1_ADD_99_U91);
  nand ginst320 (P1_ADD_99_U142, P1_REG3_REG_15__SCAN_IN, P1_ADD_99_U27);
  nand ginst321 (P1_ADD_99_U143, P1_ADD_99_U28, P1_ADD_99_U90);
  nand ginst322 (P1_ADD_99_U144, P1_REG3_REG_14__SCAN_IN, P1_ADD_99_U25);
  nand ginst323 (P1_ADD_99_U145, P1_ADD_99_U26, P1_ADD_99_U89);
  nand ginst324 (P1_ADD_99_U146, P1_REG3_REG_13__SCAN_IN, P1_ADD_99_U23);
  nand ginst325 (P1_ADD_99_U147, P1_ADD_99_U24, P1_ADD_99_U88);
  nand ginst326 (P1_ADD_99_U148, P1_REG3_REG_12__SCAN_IN, P1_ADD_99_U21);
  nand ginst327 (P1_ADD_99_U149, P1_ADD_99_U22, P1_ADD_99_U87);
  not ginst328 (P1_ADD_99_U15, P1_REG3_REG_9__SCAN_IN);
  nand ginst329 (P1_ADD_99_U150, P1_REG3_REG_11__SCAN_IN, P1_ADD_99_U19);
  nand ginst330 (P1_ADD_99_U151, P1_ADD_99_U20, P1_ADD_99_U86);
  nand ginst331 (P1_ADD_99_U152, P1_REG3_REG_10__SCAN_IN, P1_ADD_99_U17);
  nand ginst332 (P1_ADD_99_U153, P1_ADD_99_U18, P1_ADD_99_U85);
  nand ginst333 (P1_ADD_99_U16, P1_REG3_REG_8__SCAN_IN, P1_ADD_99_U83);
  nand ginst334 (P1_ADD_99_U17, P1_REG3_REG_9__SCAN_IN, P1_ADD_99_U84);
  not ginst335 (P1_ADD_99_U18, P1_REG3_REG_10__SCAN_IN);
  nand ginst336 (P1_ADD_99_U19, P1_REG3_REG_10__SCAN_IN, P1_ADD_99_U85);
  not ginst337 (P1_ADD_99_U20, P1_REG3_REG_11__SCAN_IN);
  nand ginst338 (P1_ADD_99_U21, P1_REG3_REG_11__SCAN_IN, P1_ADD_99_U86);
  not ginst339 (P1_ADD_99_U22, P1_REG3_REG_12__SCAN_IN);
  nand ginst340 (P1_ADD_99_U23, P1_REG3_REG_12__SCAN_IN, P1_ADD_99_U87);
  not ginst341 (P1_ADD_99_U24, P1_REG3_REG_13__SCAN_IN);
  nand ginst342 (P1_ADD_99_U25, P1_REG3_REG_13__SCAN_IN, P1_ADD_99_U88);
  not ginst343 (P1_ADD_99_U26, P1_REG3_REG_14__SCAN_IN);
  nand ginst344 (P1_ADD_99_U27, P1_REG3_REG_14__SCAN_IN, P1_ADD_99_U89);
  not ginst345 (P1_ADD_99_U28, P1_REG3_REG_15__SCAN_IN);
  nand ginst346 (P1_ADD_99_U29, P1_REG3_REG_15__SCAN_IN, P1_ADD_99_U90);
  not ginst347 (P1_ADD_99_U30, P1_REG3_REG_16__SCAN_IN);
  nand ginst348 (P1_ADD_99_U31, P1_REG3_REG_16__SCAN_IN, P1_ADD_99_U91);
  not ginst349 (P1_ADD_99_U32, P1_REG3_REG_17__SCAN_IN);
  nand ginst350 (P1_ADD_99_U33, P1_REG3_REG_17__SCAN_IN, P1_ADD_99_U92);
  not ginst351 (P1_ADD_99_U34, P1_REG3_REG_18__SCAN_IN);
  nand ginst352 (P1_ADD_99_U35, P1_REG3_REG_18__SCAN_IN, P1_ADD_99_U93);
  not ginst353 (P1_ADD_99_U36, P1_REG3_REG_19__SCAN_IN);
  nand ginst354 (P1_ADD_99_U37, P1_REG3_REG_19__SCAN_IN, P1_ADD_99_U94);
  not ginst355 (P1_ADD_99_U38, P1_REG3_REG_20__SCAN_IN);
  nand ginst356 (P1_ADD_99_U39, P1_REG3_REG_20__SCAN_IN, P1_ADD_99_U95);
  not ginst357 (P1_ADD_99_U4, P1_REG3_REG_3__SCAN_IN);
  not ginst358 (P1_ADD_99_U40, P1_REG3_REG_21__SCAN_IN);
  nand ginst359 (P1_ADD_99_U41, P1_REG3_REG_21__SCAN_IN, P1_ADD_99_U96);
  not ginst360 (P1_ADD_99_U42, P1_REG3_REG_22__SCAN_IN);
  nand ginst361 (P1_ADD_99_U43, P1_REG3_REG_22__SCAN_IN, P1_ADD_99_U97);
  not ginst362 (P1_ADD_99_U44, P1_REG3_REG_23__SCAN_IN);
  nand ginst363 (P1_ADD_99_U45, P1_REG3_REG_23__SCAN_IN, P1_ADD_99_U98);
  not ginst364 (P1_ADD_99_U46, P1_REG3_REG_24__SCAN_IN);
  nand ginst365 (P1_ADD_99_U47, P1_REG3_REG_24__SCAN_IN, P1_ADD_99_U99);
  not ginst366 (P1_ADD_99_U48, P1_REG3_REG_25__SCAN_IN);
  nand ginst367 (P1_ADD_99_U49, P1_REG3_REG_25__SCAN_IN, P1_ADD_99_U100);
  and ginst368 (P1_ADD_99_U5, P1_REG3_REG_28__SCAN_IN, P1_REG3_REG_27__SCAN_IN, P1_ADD_99_U102);
  not ginst369 (P1_ADD_99_U50, P1_REG3_REG_26__SCAN_IN);
  nand ginst370 (P1_ADD_99_U51, P1_REG3_REG_26__SCAN_IN, P1_ADD_99_U101);
  not ginst371 (P1_ADD_99_U52, P1_REG3_REG_28__SCAN_IN);
  not ginst372 (P1_ADD_99_U53, P1_REG3_REG_27__SCAN_IN);
  nand ginst373 (P1_ADD_99_U54, P1_ADD_99_U104, P1_ADD_99_U105);
  nand ginst374 (P1_ADD_99_U55, P1_ADD_99_U106, P1_ADD_99_U107);
  nand ginst375 (P1_ADD_99_U56, P1_ADD_99_U108, P1_ADD_99_U109);
  nand ginst376 (P1_ADD_99_U57, P1_ADD_99_U110, P1_ADD_99_U111);
  nand ginst377 (P1_ADD_99_U58, P1_ADD_99_U112, P1_ADD_99_U113);
  nand ginst378 (P1_ADD_99_U59, P1_ADD_99_U114, P1_ADD_99_U115);
  not ginst379 (P1_ADD_99_U6, P1_REG3_REG_4__SCAN_IN);
  nand ginst380 (P1_ADD_99_U60, P1_ADD_99_U116, P1_ADD_99_U117);
  nand ginst381 (P1_ADD_99_U61, P1_ADD_99_U118, P1_ADD_99_U119);
  nand ginst382 (P1_ADD_99_U62, P1_ADD_99_U120, P1_ADD_99_U121);
  nand ginst383 (P1_ADD_99_U63, P1_ADD_99_U122, P1_ADD_99_U123);
  nand ginst384 (P1_ADD_99_U64, P1_ADD_99_U124, P1_ADD_99_U125);
  nand ginst385 (P1_ADD_99_U65, P1_ADD_99_U126, P1_ADD_99_U127);
  nand ginst386 (P1_ADD_99_U66, P1_ADD_99_U128, P1_ADD_99_U129);
  nand ginst387 (P1_ADD_99_U67, P1_ADD_99_U130, P1_ADD_99_U131);
  nand ginst388 (P1_ADD_99_U68, P1_ADD_99_U132, P1_ADD_99_U133);
  nand ginst389 (P1_ADD_99_U69, P1_ADD_99_U134, P1_ADD_99_U135);
  nand ginst390 (P1_ADD_99_U7, P1_REG3_REG_4__SCAN_IN, P1_REG3_REG_3__SCAN_IN);
  nand ginst391 (P1_ADD_99_U70, P1_ADD_99_U136, P1_ADD_99_U137);
  nand ginst392 (P1_ADD_99_U71, P1_ADD_99_U138, P1_ADD_99_U139);
  nand ginst393 (P1_ADD_99_U72, P1_ADD_99_U140, P1_ADD_99_U141);
  nand ginst394 (P1_ADD_99_U73, P1_ADD_99_U142, P1_ADD_99_U143);
  nand ginst395 (P1_ADD_99_U74, P1_ADD_99_U144, P1_ADD_99_U145);
  nand ginst396 (P1_ADD_99_U75, P1_ADD_99_U146, P1_ADD_99_U147);
  nand ginst397 (P1_ADD_99_U76, P1_ADD_99_U148, P1_ADD_99_U149);
  nand ginst398 (P1_ADD_99_U77, P1_ADD_99_U150, P1_ADD_99_U151);
  nand ginst399 (P1_ADD_99_U78, P1_ADD_99_U152, P1_ADD_99_U153);
  nand ginst400 (P1_ADD_99_U79, P1_REG3_REG_27__SCAN_IN, P1_ADD_99_U102);
  not ginst401 (P1_ADD_99_U8, P1_REG3_REG_5__SCAN_IN);
  not ginst402 (P1_ADD_99_U80, P1_ADD_99_U7);
  not ginst403 (P1_ADD_99_U81, P1_ADD_99_U9);
  not ginst404 (P1_ADD_99_U82, P1_ADD_99_U11);
  not ginst405 (P1_ADD_99_U83, P1_ADD_99_U13);
  not ginst406 (P1_ADD_99_U84, P1_ADD_99_U16);
  not ginst407 (P1_ADD_99_U85, P1_ADD_99_U17);
  not ginst408 (P1_ADD_99_U86, P1_ADD_99_U19);
  not ginst409 (P1_ADD_99_U87, P1_ADD_99_U21);
  not ginst410 (P1_ADD_99_U88, P1_ADD_99_U23);
  not ginst411 (P1_ADD_99_U89, P1_ADD_99_U25);
  nand ginst412 (P1_ADD_99_U9, P1_REG3_REG_5__SCAN_IN, P1_ADD_99_U80);
  not ginst413 (P1_ADD_99_U90, P1_ADD_99_U27);
  not ginst414 (P1_ADD_99_U91, P1_ADD_99_U29);
  not ginst415 (P1_ADD_99_U92, P1_ADD_99_U31);
  not ginst416 (P1_ADD_99_U93, P1_ADD_99_U33);
  not ginst417 (P1_ADD_99_U94, P1_ADD_99_U35);
  not ginst418 (P1_ADD_99_U95, P1_ADD_99_U37);
  not ginst419 (P1_ADD_99_U96, P1_ADD_99_U39);
  not ginst420 (P1_ADD_99_U97, P1_ADD_99_U41);
  not ginst421 (P1_ADD_99_U98, P1_ADD_99_U43);
  not ginst422 (P1_ADD_99_U99, P1_ADD_99_U45);
  and ginst423 (P1_R1105_U10, P1_R1105_U215, P1_R1105_U218);
  not ginst424 (P1_R1105_U100, P1_R1105_U40);
  not ginst425 (P1_R1105_U101, P1_R1105_U41);
  nand ginst426 (P1_R1105_U102, P1_R1105_U40, P1_R1105_U41);
  nand ginst427 (P1_R1105_U103, P1_REG2_REG_2__SCAN_IN, P1_R1105_U96, P1_U3463);
  nand ginst428 (P1_R1105_U104, P1_R1105_U102, P1_R1105_U5);
  nand ginst429 (P1_R1105_U105, P1_REG2_REG_3__SCAN_IN, P1_U3466);
  nand ginst430 (P1_R1105_U106, P1_R1105_U103, P1_R1105_U104, P1_R1105_U105);
  nand ginst431 (P1_R1105_U107, P1_R1105_U32, P1_R1105_U33);
  nand ginst432 (P1_R1105_U108, P1_R1105_U107, P1_U3472);
  nand ginst433 (P1_R1105_U109, P1_R1105_U106, P1_R1105_U4);
  and ginst434 (P1_R1105_U11, P1_R1105_U208, P1_R1105_U211);
  nand ginst435 (P1_R1105_U110, P1_REG2_REG_5__SCAN_IN, P1_R1105_U89);
  not ginst436 (P1_R1105_U111, P1_R1105_U39);
  or ginst437 (P1_R1105_U112, P1_REG2_REG_7__SCAN_IN, P1_U3478);
  or ginst438 (P1_R1105_U113, P1_REG2_REG_6__SCAN_IN, P1_U3475);
  not ginst439 (P1_R1105_U114, P1_R1105_U20);
  nand ginst440 (P1_R1105_U115, P1_R1105_U20, P1_R1105_U21);
  nand ginst441 (P1_R1105_U116, P1_R1105_U115, P1_U3478);
  nand ginst442 (P1_R1105_U117, P1_REG2_REG_7__SCAN_IN, P1_R1105_U114);
  nand ginst443 (P1_R1105_U118, P1_R1105_U39, P1_R1105_U6);
  not ginst444 (P1_R1105_U119, P1_R1105_U81);
  and ginst445 (P1_R1105_U12, P1_R1105_U199, P1_R1105_U202);
  or ginst446 (P1_R1105_U120, P1_REG2_REG_8__SCAN_IN, P1_U3481);
  nand ginst447 (P1_R1105_U121, P1_R1105_U120, P1_R1105_U81);
  not ginst448 (P1_R1105_U122, P1_R1105_U38);
  or ginst449 (P1_R1105_U123, P1_REG2_REG_9__SCAN_IN, P1_U3484);
  or ginst450 (P1_R1105_U124, P1_REG2_REG_6__SCAN_IN, P1_U3475);
  nand ginst451 (P1_R1105_U125, P1_R1105_U124, P1_R1105_U39);
  nand ginst452 (P1_R1105_U126, P1_R1105_U125, P1_R1105_U20, P1_R1105_U237, P1_R1105_U238);
  nand ginst453 (P1_R1105_U127, P1_R1105_U111, P1_R1105_U20);
  nand ginst454 (P1_R1105_U128, P1_REG2_REG_7__SCAN_IN, P1_U3478);
  nand ginst455 (P1_R1105_U129, P1_R1105_U127, P1_R1105_U128, P1_R1105_U6);
  and ginst456 (P1_R1105_U13, P1_R1105_U192, P1_R1105_U196);
  or ginst457 (P1_R1105_U130, P1_REG2_REG_6__SCAN_IN, P1_U3475);
  nand ginst458 (P1_R1105_U131, P1_R1105_U101, P1_R1105_U97);
  nand ginst459 (P1_R1105_U132, P1_REG2_REG_2__SCAN_IN, P1_U3463);
  not ginst460 (P1_R1105_U133, P1_R1105_U43);
  nand ginst461 (P1_R1105_U134, P1_R1105_U100, P1_R1105_U5);
  nand ginst462 (P1_R1105_U135, P1_R1105_U43, P1_R1105_U96);
  nand ginst463 (P1_R1105_U136, P1_REG2_REG_3__SCAN_IN, P1_U3466);
  not ginst464 (P1_R1105_U137, P1_R1105_U42);
  or ginst465 (P1_R1105_U138, P1_REG2_REG_4__SCAN_IN, P1_U3469);
  nand ginst466 (P1_R1105_U139, P1_R1105_U138, P1_R1105_U42);
  and ginst467 (P1_R1105_U14, P1_R1105_U148, P1_R1105_U151);
  nand ginst468 (P1_R1105_U140, P1_R1105_U139, P1_R1105_U244, P1_R1105_U245, P1_R1105_U32);
  nand ginst469 (P1_R1105_U141, P1_R1105_U137, P1_R1105_U32);
  nand ginst470 (P1_R1105_U142, P1_REG2_REG_5__SCAN_IN, P1_U3472);
  nand ginst471 (P1_R1105_U143, P1_R1105_U141, P1_R1105_U142, P1_R1105_U4);
  or ginst472 (P1_R1105_U144, P1_REG2_REG_4__SCAN_IN, P1_U3469);
  nand ginst473 (P1_R1105_U145, P1_R1105_U100, P1_R1105_U97);
  not ginst474 (P1_R1105_U146, P1_R1105_U82);
  nand ginst475 (P1_R1105_U147, P1_REG2_REG_3__SCAN_IN, P1_U3466);
  nand ginst476 (P1_R1105_U148, P1_R1105_U256, P1_R1105_U257, P1_R1105_U40, P1_R1105_U41);
  nand ginst477 (P1_R1105_U149, P1_R1105_U40, P1_R1105_U41);
  and ginst478 (P1_R1105_U15, P1_R1105_U140, P1_R1105_U143);
  nand ginst479 (P1_R1105_U150, P1_REG2_REG_2__SCAN_IN, P1_U3463);
  nand ginst480 (P1_R1105_U151, P1_R1105_U149, P1_R1105_U150, P1_R1105_U97);
  or ginst481 (P1_R1105_U152, P1_REG2_REG_1__SCAN_IN, P1_U3460);
  not ginst482 (P1_R1105_U153, P1_R1105_U83);
  or ginst483 (P1_R1105_U154, P1_REG2_REG_9__SCAN_IN, P1_U3484);
  or ginst484 (P1_R1105_U155, P1_REG2_REG_10__SCAN_IN, P1_U3487);
  nand ginst485 (P1_R1105_U156, P1_R1105_U7, P1_R1105_U93);
  nand ginst486 (P1_R1105_U157, P1_REG2_REG_10__SCAN_IN, P1_U3487);
  nand ginst487 (P1_R1105_U158, P1_R1105_U156, P1_R1105_U157, P1_R1105_U90);
  or ginst488 (P1_R1105_U159, P1_REG2_REG_10__SCAN_IN, P1_U3487);
  and ginst489 (P1_R1105_U16, P1_R1105_U126, P1_R1105_U129);
  nand ginst490 (P1_R1105_U160, P1_R1105_U120, P1_R1105_U7, P1_R1105_U81);
  nand ginst491 (P1_R1105_U161, P1_R1105_U158, P1_R1105_U159);
  not ginst492 (P1_R1105_U162, P1_R1105_U88);
  or ginst493 (P1_R1105_U163, P1_REG2_REG_13__SCAN_IN, P1_U3496);
  or ginst494 (P1_R1105_U164, P1_REG2_REG_12__SCAN_IN, P1_U3493);
  nand ginst495 (P1_R1105_U165, P1_R1105_U8, P1_R1105_U92);
  nand ginst496 (P1_R1105_U166, P1_REG2_REG_13__SCAN_IN, P1_U3496);
  nand ginst497 (P1_R1105_U167, P1_R1105_U165, P1_R1105_U166, P1_R1105_U91);
  or ginst498 (P1_R1105_U168, P1_REG2_REG_11__SCAN_IN, P1_U3490);
  or ginst499 (P1_R1105_U169, P1_REG2_REG_13__SCAN_IN, P1_U3496);
  not ginst500 (P1_R1105_U17, P1_REG2_REG_6__SCAN_IN);
  nand ginst501 (P1_R1105_U170, P1_R1105_U168, P1_R1105_U8, P1_R1105_U88);
  nand ginst502 (P1_R1105_U171, P1_R1105_U167, P1_R1105_U169);
  not ginst503 (P1_R1105_U172, P1_R1105_U87);
  or ginst504 (P1_R1105_U173, P1_REG2_REG_14__SCAN_IN, P1_U3499);
  nand ginst505 (P1_R1105_U174, P1_R1105_U173, P1_R1105_U87);
  nand ginst506 (P1_R1105_U175, P1_REG2_REG_14__SCAN_IN, P1_U3499);
  not ginst507 (P1_R1105_U176, P1_R1105_U86);
  or ginst508 (P1_R1105_U177, P1_REG2_REG_15__SCAN_IN, P1_U3502);
  nand ginst509 (P1_R1105_U178, P1_R1105_U177, P1_R1105_U86);
  nand ginst510 (P1_R1105_U179, P1_REG2_REG_15__SCAN_IN, P1_U3502);
  not ginst511 (P1_R1105_U18, P1_U3475);
  not ginst512 (P1_R1105_U180, P1_R1105_U66);
  or ginst513 (P1_R1105_U181, P1_REG2_REG_17__SCAN_IN, P1_U3508);
  or ginst514 (P1_R1105_U182, P1_REG2_REG_16__SCAN_IN, P1_U3505);
  not ginst515 (P1_R1105_U183, P1_R1105_U47);
  nand ginst516 (P1_R1105_U184, P1_R1105_U47, P1_R1105_U48);
  nand ginst517 (P1_R1105_U185, P1_R1105_U184, P1_U3508);
  nand ginst518 (P1_R1105_U186, P1_REG2_REG_17__SCAN_IN, P1_R1105_U183);
  nand ginst519 (P1_R1105_U187, P1_R1105_U66, P1_R1105_U9);
  not ginst520 (P1_R1105_U188, P1_R1105_U65);
  or ginst521 (P1_R1105_U189, P1_REG2_REG_18__SCAN_IN, P1_U3511);
  not ginst522 (P1_R1105_U19, P1_U3478);
  nand ginst523 (P1_R1105_U190, P1_R1105_U189, P1_R1105_U65);
  nand ginst524 (P1_R1105_U191, P1_REG2_REG_18__SCAN_IN, P1_U3511);
  nand ginst525 (P1_R1105_U192, P1_R1105_U190, P1_R1105_U191, P1_R1105_U260, P1_R1105_U261);
  nand ginst526 (P1_R1105_U193, P1_REG2_REG_18__SCAN_IN, P1_U3511);
  nand ginst527 (P1_R1105_U194, P1_R1105_U188, P1_R1105_U193);
  or ginst528 (P1_R1105_U195, P1_REG2_REG_18__SCAN_IN, P1_U3511);
  nand ginst529 (P1_R1105_U196, P1_R1105_U194, P1_R1105_U195, P1_R1105_U264);
  or ginst530 (P1_R1105_U197, P1_REG2_REG_16__SCAN_IN, P1_U3505);
  nand ginst531 (P1_R1105_U198, P1_R1105_U197, P1_R1105_U66);
  nand ginst532 (P1_R1105_U199, P1_R1105_U198, P1_R1105_U272, P1_R1105_U273, P1_R1105_U47);
  nand ginst533 (P1_R1105_U20, P1_REG2_REG_6__SCAN_IN, P1_U3475);
  nand ginst534 (P1_R1105_U200, P1_R1105_U180, P1_R1105_U47);
  nand ginst535 (P1_R1105_U201, P1_REG2_REG_17__SCAN_IN, P1_U3508);
  nand ginst536 (P1_R1105_U202, P1_R1105_U200, P1_R1105_U201, P1_R1105_U9);
  or ginst537 (P1_R1105_U203, P1_REG2_REG_16__SCAN_IN, P1_U3505);
  nand ginst538 (P1_R1105_U204, P1_R1105_U168, P1_R1105_U88);
  not ginst539 (P1_R1105_U205, P1_R1105_U67);
  or ginst540 (P1_R1105_U206, P1_REG2_REG_12__SCAN_IN, P1_U3493);
  nand ginst541 (P1_R1105_U207, P1_R1105_U206, P1_R1105_U67);
  nand ginst542 (P1_R1105_U208, P1_R1105_U207, P1_R1105_U293, P1_R1105_U294, P1_R1105_U91);
  nand ginst543 (P1_R1105_U209, P1_R1105_U205, P1_R1105_U91);
  not ginst544 (P1_R1105_U21, P1_REG2_REG_7__SCAN_IN);
  nand ginst545 (P1_R1105_U210, P1_REG2_REG_13__SCAN_IN, P1_U3496);
  nand ginst546 (P1_R1105_U211, P1_R1105_U209, P1_R1105_U210, P1_R1105_U8);
  or ginst547 (P1_R1105_U212, P1_REG2_REG_12__SCAN_IN, P1_U3493);
  or ginst548 (P1_R1105_U213, P1_REG2_REG_9__SCAN_IN, P1_U3484);
  nand ginst549 (P1_R1105_U214, P1_R1105_U213, P1_R1105_U38);
  nand ginst550 (P1_R1105_U215, P1_R1105_U214, P1_R1105_U305, P1_R1105_U306, P1_R1105_U90);
  nand ginst551 (P1_R1105_U216, P1_R1105_U122, P1_R1105_U90);
  nand ginst552 (P1_R1105_U217, P1_REG2_REG_10__SCAN_IN, P1_U3487);
  nand ginst553 (P1_R1105_U218, P1_R1105_U216, P1_R1105_U217, P1_R1105_U7);
  nand ginst554 (P1_R1105_U219, P1_R1105_U123, P1_R1105_U90);
  not ginst555 (P1_R1105_U22, P1_REG2_REG_4__SCAN_IN);
  nand ginst556 (P1_R1105_U220, P1_R1105_U120, P1_R1105_U49);
  nand ginst557 (P1_R1105_U221, P1_R1105_U130, P1_R1105_U20);
  nand ginst558 (P1_R1105_U222, P1_R1105_U144, P1_R1105_U32);
  nand ginst559 (P1_R1105_U223, P1_R1105_U147, P1_R1105_U96);
  nand ginst560 (P1_R1105_U224, P1_R1105_U203, P1_R1105_U47);
  nand ginst561 (P1_R1105_U225, P1_R1105_U212, P1_R1105_U91);
  nand ginst562 (P1_R1105_U226, P1_R1105_U168, P1_R1105_U56);
  nand ginst563 (P1_R1105_U227, P1_R1105_U37, P1_U3484);
  nand ginst564 (P1_R1105_U228, P1_REG2_REG_9__SCAN_IN, P1_R1105_U36);
  nand ginst565 (P1_R1105_U229, P1_R1105_U227, P1_R1105_U228);
  not ginst566 (P1_R1105_U23, P1_U3469);
  nand ginst567 (P1_R1105_U230, P1_R1105_U219, P1_R1105_U38);
  nand ginst568 (P1_R1105_U231, P1_R1105_U122, P1_R1105_U229);
  nand ginst569 (P1_R1105_U232, P1_R1105_U34, P1_U3481);
  nand ginst570 (P1_R1105_U233, P1_REG2_REG_8__SCAN_IN, P1_R1105_U35);
  nand ginst571 (P1_R1105_U234, P1_R1105_U232, P1_R1105_U233);
  nand ginst572 (P1_R1105_U235, P1_R1105_U220, P1_R1105_U81);
  nand ginst573 (P1_R1105_U236, P1_R1105_U119, P1_R1105_U234);
  nand ginst574 (P1_R1105_U237, P1_R1105_U21, P1_U3478);
  nand ginst575 (P1_R1105_U238, P1_REG2_REG_7__SCAN_IN, P1_R1105_U19);
  nand ginst576 (P1_R1105_U239, P1_R1105_U17, P1_U3475);
  not ginst577 (P1_R1105_U24, P1_U3472);
  nand ginst578 (P1_R1105_U240, P1_REG2_REG_6__SCAN_IN, P1_R1105_U18);
  nand ginst579 (P1_R1105_U241, P1_R1105_U239, P1_R1105_U240);
  nand ginst580 (P1_R1105_U242, P1_R1105_U221, P1_R1105_U39);
  nand ginst581 (P1_R1105_U243, P1_R1105_U111, P1_R1105_U241);
  nand ginst582 (P1_R1105_U244, P1_R1105_U33, P1_U3472);
  nand ginst583 (P1_R1105_U245, P1_REG2_REG_5__SCAN_IN, P1_R1105_U24);
  nand ginst584 (P1_R1105_U246, P1_R1105_U22, P1_U3469);
  nand ginst585 (P1_R1105_U247, P1_REG2_REG_4__SCAN_IN, P1_R1105_U23);
  nand ginst586 (P1_R1105_U248, P1_R1105_U246, P1_R1105_U247);
  nand ginst587 (P1_R1105_U249, P1_R1105_U222, P1_R1105_U42);
  not ginst588 (P1_R1105_U25, P1_REG2_REG_2__SCAN_IN);
  nand ginst589 (P1_R1105_U250, P1_R1105_U137, P1_R1105_U248);
  nand ginst590 (P1_R1105_U251, P1_R1105_U30, P1_U3466);
  nand ginst591 (P1_R1105_U252, P1_REG2_REG_3__SCAN_IN, P1_R1105_U31);
  nand ginst592 (P1_R1105_U253, P1_R1105_U251, P1_R1105_U252);
  nand ginst593 (P1_R1105_U254, P1_R1105_U223, P1_R1105_U82);
  nand ginst594 (P1_R1105_U255, P1_R1105_U146, P1_R1105_U253);
  nand ginst595 (P1_R1105_U256, P1_R1105_U25, P1_U3463);
  nand ginst596 (P1_R1105_U257, P1_REG2_REG_2__SCAN_IN, P1_R1105_U26);
  nand ginst597 (P1_R1105_U258, P1_R1105_U83, P1_R1105_U98);
  nand ginst598 (P1_R1105_U259, P1_R1105_U153, P1_R1105_U29);
  not ginst599 (P1_R1105_U26, P1_U3463);
  nand ginst600 (P1_R1105_U260, P1_R1105_U85, P1_U3452);
  nand ginst601 (P1_R1105_U261, P1_REG2_REG_19__SCAN_IN, P1_R1105_U84);
  nand ginst602 (P1_R1105_U262, P1_R1105_U85, P1_U3452);
  nand ginst603 (P1_R1105_U263, P1_REG2_REG_19__SCAN_IN, P1_R1105_U84);
  nand ginst604 (P1_R1105_U264, P1_R1105_U262, P1_R1105_U263);
  nand ginst605 (P1_R1105_U265, P1_R1105_U63, P1_U3511);
  nand ginst606 (P1_R1105_U266, P1_REG2_REG_18__SCAN_IN, P1_R1105_U64);
  nand ginst607 (P1_R1105_U267, P1_R1105_U63, P1_U3511);
  nand ginst608 (P1_R1105_U268, P1_REG2_REG_18__SCAN_IN, P1_R1105_U64);
  nand ginst609 (P1_R1105_U269, P1_R1105_U267, P1_R1105_U268);
  not ginst610 (P1_R1105_U27, P1_REG2_REG_0__SCAN_IN);
  nand ginst611 (P1_R1105_U270, P1_R1105_U265, P1_R1105_U266, P1_R1105_U65);
  nand ginst612 (P1_R1105_U271, P1_R1105_U188, P1_R1105_U269);
  nand ginst613 (P1_R1105_U272, P1_R1105_U48, P1_U3508);
  nand ginst614 (P1_R1105_U273, P1_REG2_REG_17__SCAN_IN, P1_R1105_U46);
  nand ginst615 (P1_R1105_U274, P1_R1105_U44, P1_U3505);
  nand ginst616 (P1_R1105_U275, P1_REG2_REG_16__SCAN_IN, P1_R1105_U45);
  nand ginst617 (P1_R1105_U276, P1_R1105_U274, P1_R1105_U275);
  nand ginst618 (P1_R1105_U277, P1_R1105_U224, P1_R1105_U66);
  nand ginst619 (P1_R1105_U278, P1_R1105_U180, P1_R1105_U276);
  nand ginst620 (P1_R1105_U279, P1_R1105_U61, P1_U3502);
  not ginst621 (P1_R1105_U28, P1_U3454);
  nand ginst622 (P1_R1105_U280, P1_REG2_REG_15__SCAN_IN, P1_R1105_U62);
  nand ginst623 (P1_R1105_U281, P1_R1105_U61, P1_U3502);
  nand ginst624 (P1_R1105_U282, P1_REG2_REG_15__SCAN_IN, P1_R1105_U62);
  nand ginst625 (P1_R1105_U283, P1_R1105_U281, P1_R1105_U282);
  nand ginst626 (P1_R1105_U284, P1_R1105_U279, P1_R1105_U280, P1_R1105_U86);
  nand ginst627 (P1_R1105_U285, P1_R1105_U176, P1_R1105_U283);
  nand ginst628 (P1_R1105_U286, P1_R1105_U59, P1_U3499);
  nand ginst629 (P1_R1105_U287, P1_REG2_REG_14__SCAN_IN, P1_R1105_U60);
  nand ginst630 (P1_R1105_U288, P1_R1105_U59, P1_U3499);
  nand ginst631 (P1_R1105_U289, P1_REG2_REG_14__SCAN_IN, P1_R1105_U60);
  nand ginst632 (P1_R1105_U29, P1_REG2_REG_0__SCAN_IN, P1_U3454);
  nand ginst633 (P1_R1105_U290, P1_R1105_U288, P1_R1105_U289);
  nand ginst634 (P1_R1105_U291, P1_R1105_U286, P1_R1105_U287, P1_R1105_U87);
  nand ginst635 (P1_R1105_U292, P1_R1105_U172, P1_R1105_U290);
  nand ginst636 (P1_R1105_U293, P1_R1105_U57, P1_U3496);
  nand ginst637 (P1_R1105_U294, P1_REG2_REG_13__SCAN_IN, P1_R1105_U58);
  nand ginst638 (P1_R1105_U295, P1_R1105_U52, P1_U3493);
  nand ginst639 (P1_R1105_U296, P1_REG2_REG_12__SCAN_IN, P1_R1105_U53);
  nand ginst640 (P1_R1105_U297, P1_R1105_U295, P1_R1105_U296);
  nand ginst641 (P1_R1105_U298, P1_R1105_U225, P1_R1105_U67);
  nand ginst642 (P1_R1105_U299, P1_R1105_U205, P1_R1105_U297);
  not ginst643 (P1_R1105_U30, P1_REG2_REG_3__SCAN_IN);
  nand ginst644 (P1_R1105_U300, P1_R1105_U54, P1_U3490);
  nand ginst645 (P1_R1105_U301, P1_REG2_REG_11__SCAN_IN, P1_R1105_U55);
  nand ginst646 (P1_R1105_U302, P1_R1105_U300, P1_R1105_U301);
  nand ginst647 (P1_R1105_U303, P1_R1105_U226, P1_R1105_U88);
  nand ginst648 (P1_R1105_U304, P1_R1105_U162, P1_R1105_U302);
  nand ginst649 (P1_R1105_U305, P1_R1105_U50, P1_U3487);
  nand ginst650 (P1_R1105_U306, P1_REG2_REG_10__SCAN_IN, P1_R1105_U51);
  nand ginst651 (P1_R1105_U307, P1_R1105_U27, P1_U3454);
  nand ginst652 (P1_R1105_U308, P1_REG2_REG_0__SCAN_IN, P1_R1105_U28);
  not ginst653 (P1_R1105_U31, P1_U3466);
  nand ginst654 (P1_R1105_U32, P1_REG2_REG_4__SCAN_IN, P1_U3469);
  not ginst655 (P1_R1105_U33, P1_REG2_REG_5__SCAN_IN);
  not ginst656 (P1_R1105_U34, P1_REG2_REG_8__SCAN_IN);
  not ginst657 (P1_R1105_U35, P1_U3481);
  not ginst658 (P1_R1105_U36, P1_U3484);
  not ginst659 (P1_R1105_U37, P1_REG2_REG_9__SCAN_IN);
  nand ginst660 (P1_R1105_U38, P1_R1105_U121, P1_R1105_U49);
  nand ginst661 (P1_R1105_U39, P1_R1105_U108, P1_R1105_U109, P1_R1105_U110);
  and ginst662 (P1_R1105_U4, P1_R1105_U94, P1_R1105_U95);
  nand ginst663 (P1_R1105_U40, P1_R1105_U98, P1_R1105_U99);
  nand ginst664 (P1_R1105_U41, P1_REG2_REG_1__SCAN_IN, P1_U3460);
  nand ginst665 (P1_R1105_U42, P1_R1105_U134, P1_R1105_U135, P1_R1105_U136);
  nand ginst666 (P1_R1105_U43, P1_R1105_U131, P1_R1105_U132);
  not ginst667 (P1_R1105_U44, P1_REG2_REG_16__SCAN_IN);
  not ginst668 (P1_R1105_U45, P1_U3505);
  not ginst669 (P1_R1105_U46, P1_U3508);
  nand ginst670 (P1_R1105_U47, P1_REG2_REG_16__SCAN_IN, P1_U3505);
  not ginst671 (P1_R1105_U48, P1_REG2_REG_17__SCAN_IN);
  nand ginst672 (P1_R1105_U49, P1_REG2_REG_8__SCAN_IN, P1_U3481);
  and ginst673 (P1_R1105_U5, P1_R1105_U96, P1_R1105_U97);
  not ginst674 (P1_R1105_U50, P1_REG2_REG_10__SCAN_IN);
  not ginst675 (P1_R1105_U51, P1_U3487);
  not ginst676 (P1_R1105_U52, P1_REG2_REG_12__SCAN_IN);
  not ginst677 (P1_R1105_U53, P1_U3493);
  not ginst678 (P1_R1105_U54, P1_REG2_REG_11__SCAN_IN);
  not ginst679 (P1_R1105_U55, P1_U3490);
  nand ginst680 (P1_R1105_U56, P1_REG2_REG_11__SCAN_IN, P1_U3490);
  not ginst681 (P1_R1105_U57, P1_REG2_REG_13__SCAN_IN);
  not ginst682 (P1_R1105_U58, P1_U3496);
  not ginst683 (P1_R1105_U59, P1_REG2_REG_14__SCAN_IN);
  and ginst684 (P1_R1105_U6, P1_R1105_U112, P1_R1105_U113);
  not ginst685 (P1_R1105_U60, P1_U3499);
  not ginst686 (P1_R1105_U61, P1_REG2_REG_15__SCAN_IN);
  not ginst687 (P1_R1105_U62, P1_U3502);
  not ginst688 (P1_R1105_U63, P1_REG2_REG_18__SCAN_IN);
  not ginst689 (P1_R1105_U64, P1_U3511);
  nand ginst690 (P1_R1105_U65, P1_R1105_U185, P1_R1105_U186, P1_R1105_U187);
  nand ginst691 (P1_R1105_U66, P1_R1105_U178, P1_R1105_U179);
  nand ginst692 (P1_R1105_U67, P1_R1105_U204, P1_R1105_U56);
  nand ginst693 (P1_R1105_U68, P1_R1105_U258, P1_R1105_U259);
  nand ginst694 (P1_R1105_U69, P1_R1105_U307, P1_R1105_U308);
  and ginst695 (P1_R1105_U7, P1_R1105_U154, P1_R1105_U155);
  nand ginst696 (P1_R1105_U70, P1_R1105_U230, P1_R1105_U231);
  nand ginst697 (P1_R1105_U71, P1_R1105_U235, P1_R1105_U236);
  nand ginst698 (P1_R1105_U72, P1_R1105_U242, P1_R1105_U243);
  nand ginst699 (P1_R1105_U73, P1_R1105_U249, P1_R1105_U250);
  nand ginst700 (P1_R1105_U74, P1_R1105_U254, P1_R1105_U255);
  nand ginst701 (P1_R1105_U75, P1_R1105_U270, P1_R1105_U271);
  nand ginst702 (P1_R1105_U76, P1_R1105_U277, P1_R1105_U278);
  nand ginst703 (P1_R1105_U77, P1_R1105_U284, P1_R1105_U285);
  nand ginst704 (P1_R1105_U78, P1_R1105_U291, P1_R1105_U292);
  nand ginst705 (P1_R1105_U79, P1_R1105_U298, P1_R1105_U299);
  and ginst706 (P1_R1105_U8, P1_R1105_U163, P1_R1105_U164);
  nand ginst707 (P1_R1105_U80, P1_R1105_U303, P1_R1105_U304);
  nand ginst708 (P1_R1105_U81, P1_R1105_U116, P1_R1105_U117, P1_R1105_U118);
  nand ginst709 (P1_R1105_U82, P1_R1105_U133, P1_R1105_U145);
  nand ginst710 (P1_R1105_U83, P1_R1105_U152, P1_R1105_U41);
  not ginst711 (P1_R1105_U84, P1_U3452);
  not ginst712 (P1_R1105_U85, P1_REG2_REG_19__SCAN_IN);
  nand ginst713 (P1_R1105_U86, P1_R1105_U174, P1_R1105_U175);
  nand ginst714 (P1_R1105_U87, P1_R1105_U170, P1_R1105_U171);
  nand ginst715 (P1_R1105_U88, P1_R1105_U160, P1_R1105_U161);
  not ginst716 (P1_R1105_U89, P1_R1105_U32);
  and ginst717 (P1_R1105_U9, P1_R1105_U181, P1_R1105_U182);
  nand ginst718 (P1_R1105_U90, P1_REG2_REG_9__SCAN_IN, P1_U3484);
  nand ginst719 (P1_R1105_U91, P1_REG2_REG_12__SCAN_IN, P1_U3493);
  not ginst720 (P1_R1105_U92, P1_R1105_U56);
  not ginst721 (P1_R1105_U93, P1_R1105_U49);
  or ginst722 (P1_R1105_U94, P1_REG2_REG_5__SCAN_IN, P1_U3472);
  or ginst723 (P1_R1105_U95, P1_REG2_REG_4__SCAN_IN, P1_U3469);
  or ginst724 (P1_R1105_U96, P1_REG2_REG_3__SCAN_IN, P1_U3466);
  or ginst725 (P1_R1105_U97, P1_REG2_REG_2__SCAN_IN, P1_U3463);
  not ginst726 (P1_R1105_U98, P1_R1105_U29);
  or ginst727 (P1_R1105_U99, P1_REG2_REG_1__SCAN_IN, P1_U3460);
  and ginst728 (P1_R1117_U10, P1_R1117_U258, P1_R1117_U259);
  nand ginst729 (P1_R1117_U100, P1_R1117_U442, P1_R1117_U443);
  nand ginst730 (P1_R1117_U101, P1_R1117_U447, P1_R1117_U448);
  nand ginst731 (P1_R1117_U102, P1_R1117_U463, P1_R1117_U464);
  nand ginst732 (P1_R1117_U103, P1_R1117_U468, P1_R1117_U469);
  nand ginst733 (P1_R1117_U104, P1_R1117_U351, P1_R1117_U352);
  nand ginst734 (P1_R1117_U105, P1_R1117_U360, P1_R1117_U361);
  nand ginst735 (P1_R1117_U106, P1_R1117_U367, P1_R1117_U368);
  nand ginst736 (P1_R1117_U107, P1_R1117_U371, P1_R1117_U372);
  nand ginst737 (P1_R1117_U108, P1_R1117_U380, P1_R1117_U381);
  nand ginst738 (P1_R1117_U109, P1_R1117_U401, P1_R1117_U402);
  and ginst739 (P1_R1117_U11, P1_R1117_U284, P1_R1117_U285);
  nand ginst740 (P1_R1117_U110, P1_R1117_U418, P1_R1117_U419);
  nand ginst741 (P1_R1117_U111, P1_R1117_U422, P1_R1117_U423);
  nand ginst742 (P1_R1117_U112, P1_R1117_U454, P1_R1117_U455);
  nand ginst743 (P1_R1117_U113, P1_R1117_U458, P1_R1117_U459);
  nand ginst744 (P1_R1117_U114, P1_R1117_U475, P1_R1117_U476);
  and ginst745 (P1_R1117_U115, P1_R1117_U183, P1_R1117_U195);
  and ginst746 (P1_R1117_U116, P1_R1117_U198, P1_R1117_U199);
  and ginst747 (P1_R1117_U117, P1_R1117_U185, P1_R1117_U211);
  and ginst748 (P1_R1117_U118, P1_R1117_U214, P1_R1117_U215);
  and ginst749 (P1_R1117_U119, P1_R1117_U353, P1_R1117_U354, P1_R1117_U40);
  and ginst750 (P1_R1117_U12, P1_R1117_U382, P1_R1117_U383);
  and ginst751 (P1_R1117_U120, P1_R1117_U185, P1_R1117_U357);
  and ginst752 (P1_R1117_U121, P1_R1117_U230, P1_R1117_U7);
  and ginst753 (P1_R1117_U122, P1_R1117_U184, P1_R1117_U364);
  and ginst754 (P1_R1117_U123, P1_R1117_U29, P1_R1117_U373, P1_R1117_U374);
  and ginst755 (P1_R1117_U124, P1_R1117_U183, P1_R1117_U377);
  and ginst756 (P1_R1117_U125, P1_R1117_U217, P1_R1117_U8);
  and ginst757 (P1_R1117_U126, P1_R1117_U180, P1_R1117_U262);
  and ginst758 (P1_R1117_U127, P1_R1117_U181, P1_R1117_U288);
  and ginst759 (P1_R1117_U128, P1_R1117_U304, P1_R1117_U305);
  and ginst760 (P1_R1117_U129, P1_R1117_U307, P1_R1117_U386);
  nand ginst761 (P1_R1117_U13, P1_R1117_U340, P1_R1117_U343);
  and ginst762 (P1_R1117_U130, P1_R1117_U304, P1_R1117_U305, P1_R1117_U308);
  nand ginst763 (P1_R1117_U131, P1_R1117_U389, P1_R1117_U390);
  and ginst764 (P1_R1117_U132, P1_R1117_U394, P1_R1117_U395, P1_R1117_U85);
  and ginst765 (P1_R1117_U133, P1_R1117_U182, P1_R1117_U398);
  nand ginst766 (P1_R1117_U134, P1_R1117_U403, P1_R1117_U404);
  nand ginst767 (P1_R1117_U135, P1_R1117_U408, P1_R1117_U409);
  and ginst768 (P1_R1117_U136, P1_R1117_U181, P1_R1117_U415);
  nand ginst769 (P1_R1117_U137, P1_R1117_U424, P1_R1117_U425);
  nand ginst770 (P1_R1117_U138, P1_R1117_U429, P1_R1117_U430);
  nand ginst771 (P1_R1117_U139, P1_R1117_U434, P1_R1117_U435);
  nand ginst772 (P1_R1117_U14, P1_R1117_U329, P1_R1117_U332);
  nand ginst773 (P1_R1117_U140, P1_R1117_U439, P1_R1117_U440);
  nand ginst774 (P1_R1117_U141, P1_R1117_U444, P1_R1117_U445);
  and ginst775 (P1_R1117_U142, P1_R1117_U180, P1_R1117_U451);
  nand ginst776 (P1_R1117_U143, P1_R1117_U460, P1_R1117_U461);
  nand ginst777 (P1_R1117_U144, P1_R1117_U465, P1_R1117_U466);
  and ginst778 (P1_R1117_U145, P1_R1117_U342, P1_R1117_U9);
  and ginst779 (P1_R1117_U146, P1_R1117_U179, P1_R1117_U472);
  and ginst780 (P1_R1117_U147, P1_R1117_U349, P1_R1117_U350);
  nand ginst781 (P1_R1117_U148, P1_R1117_U118, P1_R1117_U212);
  and ginst782 (P1_R1117_U149, P1_R1117_U358, P1_R1117_U359);
  nand ginst783 (P1_R1117_U15, P1_R1117_U318, P1_R1117_U321);
  and ginst784 (P1_R1117_U150, P1_R1117_U365, P1_R1117_U366);
  and ginst785 (P1_R1117_U151, P1_R1117_U369, P1_R1117_U370);
  nand ginst786 (P1_R1117_U152, P1_R1117_U116, P1_R1117_U196);
  and ginst787 (P1_R1117_U153, P1_R1117_U378, P1_R1117_U379);
  not ginst788 (P1_R1117_U154, P1_U4028);
  not ginst789 (P1_R1117_U155, P1_U3055);
  and ginst790 (P1_R1117_U156, P1_R1117_U387, P1_R1117_U388);
  nand ginst791 (P1_R1117_U157, P1_R1117_U128, P1_R1117_U302);
  and ginst792 (P1_R1117_U158, P1_R1117_U399, P1_R1117_U400);
  nand ginst793 (P1_R1117_U159, P1_R1117_U294, P1_R1117_U295);
  nand ginst794 (P1_R1117_U16, P1_R1117_U310, P1_R1117_U312);
  nand ginst795 (P1_R1117_U160, P1_R1117_U290, P1_R1117_U291);
  and ginst796 (P1_R1117_U161, P1_R1117_U416, P1_R1117_U417);
  and ginst797 (P1_R1117_U162, P1_R1117_U420, P1_R1117_U421);
  nand ginst798 (P1_R1117_U163, P1_R1117_U280, P1_R1117_U281);
  nand ginst799 (P1_R1117_U164, P1_R1117_U276, P1_R1117_U277);
  not ginst800 (P1_R1117_U165, P1_U3461);
  nand ginst801 (P1_R1117_U166, P1_R1117_U272, P1_R1117_U273);
  not ginst802 (P1_R1117_U167, P1_U3512);
  nand ginst803 (P1_R1117_U168, P1_R1117_U264, P1_R1117_U265);
  and ginst804 (P1_R1117_U169, P1_R1117_U452, P1_R1117_U453);
  nand ginst805 (P1_R1117_U17, P1_R1117_U156, P1_R1117_U175, P1_R1117_U348);
  and ginst806 (P1_R1117_U170, P1_R1117_U456, P1_R1117_U457);
  nand ginst807 (P1_R1117_U171, P1_R1117_U254, P1_R1117_U255);
  nand ginst808 (P1_R1117_U172, P1_R1117_U250, P1_R1117_U251);
  nand ginst809 (P1_R1117_U173, P1_R1117_U246, P1_R1117_U247);
  and ginst810 (P1_R1117_U174, P1_R1117_U473, P1_R1117_U474);
  nand ginst811 (P1_R1117_U175, P1_R1117_U129, P1_R1117_U157);
  not ginst812 (P1_R1117_U176, P1_R1117_U85);
  not ginst813 (P1_R1117_U177, P1_R1117_U29);
  not ginst814 (P1_R1117_U178, P1_R1117_U40);
  nand ginst815 (P1_R1117_U179, P1_R1117_U53, P1_U3488);
  nand ginst816 (P1_R1117_U18, P1_R1117_U236, P1_R1117_U238);
  nand ginst817 (P1_R1117_U180, P1_R1117_U62, P1_U3503);
  nand ginst818 (P1_R1117_U181, P1_R1117_U76, P1_U4023);
  nand ginst819 (P1_R1117_U182, P1_R1117_U84, P1_U4019);
  nand ginst820 (P1_R1117_U183, P1_R1117_U28, P1_U3464);
  nand ginst821 (P1_R1117_U184, P1_R1117_U35, P1_U3473);
  nand ginst822 (P1_R1117_U185, P1_R1117_U39, P1_U3479);
  not ginst823 (P1_R1117_U186, P1_R1117_U64);
  not ginst824 (P1_R1117_U187, P1_R1117_U78);
  not ginst825 (P1_R1117_U188, P1_R1117_U37);
  not ginst826 (P1_R1117_U189, P1_R1117_U54);
  nand ginst827 (P1_R1117_U19, P1_R1117_U228, P1_R1117_U231);
  not ginst828 (P1_R1117_U190, P1_R1117_U25);
  nand ginst829 (P1_R1117_U191, P1_R1117_U190, P1_R1117_U26);
  nand ginst830 (P1_R1117_U192, P1_R1117_U165, P1_R1117_U191);
  nand ginst831 (P1_R1117_U193, P1_R1117_U25, P1_U3078);
  not ginst832 (P1_R1117_U194, P1_R1117_U46);
  nand ginst833 (P1_R1117_U195, P1_R1117_U30, P1_U3467);
  nand ginst834 (P1_R1117_U196, P1_R1117_U115, P1_R1117_U46);
  nand ginst835 (P1_R1117_U197, P1_R1117_U29, P1_R1117_U30);
  nand ginst836 (P1_R1117_U198, P1_R1117_U197, P1_R1117_U27);
  nand ginst837 (P1_R1117_U199, P1_R1117_U177, P1_U3064);
  nand ginst838 (P1_R1117_U20, P1_R1117_U220, P1_R1117_U222);
  not ginst839 (P1_R1117_U200, P1_R1117_U152);
  nand ginst840 (P1_R1117_U201, P1_R1117_U34, P1_U3476);
  nand ginst841 (P1_R1117_U202, P1_R1117_U31, P1_U3071);
  nand ginst842 (P1_R1117_U203, P1_R1117_U32, P1_U3067);
  nand ginst843 (P1_R1117_U204, P1_R1117_U188, P1_R1117_U6);
  nand ginst844 (P1_R1117_U205, P1_R1117_U204, P1_R1117_U7);
  nand ginst845 (P1_R1117_U206, P1_R1117_U36, P1_U3470);
  nand ginst846 (P1_R1117_U207, P1_R1117_U34, P1_U3476);
  nand ginst847 (P1_R1117_U208, P1_R1117_U152, P1_R1117_U206, P1_R1117_U6);
  nand ginst848 (P1_R1117_U209, P1_R1117_U205, P1_R1117_U207);
  nand ginst849 (P1_R1117_U21, P1_R1117_U25, P1_R1117_U346);
  not ginst850 (P1_R1117_U210, P1_R1117_U44);
  nand ginst851 (P1_R1117_U211, P1_R1117_U41, P1_U3482);
  nand ginst852 (P1_R1117_U212, P1_R1117_U117, P1_R1117_U44);
  nand ginst853 (P1_R1117_U213, P1_R1117_U40, P1_R1117_U41);
  nand ginst854 (P1_R1117_U214, P1_R1117_U213, P1_R1117_U38);
  nand ginst855 (P1_R1117_U215, P1_R1117_U178, P1_U3084);
  not ginst856 (P1_R1117_U216, P1_R1117_U148);
  nand ginst857 (P1_R1117_U217, P1_R1117_U43, P1_U3485);
  nand ginst858 (P1_R1117_U218, P1_R1117_U217, P1_R1117_U54);
  nand ginst859 (P1_R1117_U219, P1_R1117_U210, P1_R1117_U40);
  not ginst860 (P1_R1117_U22, P1_U3479);
  nand ginst861 (P1_R1117_U220, P1_R1117_U120, P1_R1117_U219);
  nand ginst862 (P1_R1117_U221, P1_R1117_U185, P1_R1117_U44);
  nand ginst863 (P1_R1117_U222, P1_R1117_U119, P1_R1117_U221);
  nand ginst864 (P1_R1117_U223, P1_R1117_U185, P1_R1117_U40);
  nand ginst865 (P1_R1117_U224, P1_R1117_U152, P1_R1117_U206);
  not ginst866 (P1_R1117_U225, P1_R1117_U45);
  nand ginst867 (P1_R1117_U226, P1_R1117_U32, P1_U3067);
  nand ginst868 (P1_R1117_U227, P1_R1117_U225, P1_R1117_U226);
  nand ginst869 (P1_R1117_U228, P1_R1117_U122, P1_R1117_U227);
  nand ginst870 (P1_R1117_U229, P1_R1117_U184, P1_R1117_U45);
  not ginst871 (P1_R1117_U23, P1_U3464);
  nand ginst872 (P1_R1117_U230, P1_R1117_U34, P1_U3476);
  nand ginst873 (P1_R1117_U231, P1_R1117_U121, P1_R1117_U229);
  nand ginst874 (P1_R1117_U232, P1_R1117_U32, P1_U3067);
  nand ginst875 (P1_R1117_U233, P1_R1117_U184, P1_R1117_U232);
  nand ginst876 (P1_R1117_U234, P1_R1117_U206, P1_R1117_U37);
  nand ginst877 (P1_R1117_U235, P1_R1117_U194, P1_R1117_U29);
  nand ginst878 (P1_R1117_U236, P1_R1117_U124, P1_R1117_U235);
  nand ginst879 (P1_R1117_U237, P1_R1117_U183, P1_R1117_U46);
  nand ginst880 (P1_R1117_U238, P1_R1117_U123, P1_R1117_U237);
  nand ginst881 (P1_R1117_U239, P1_R1117_U183, P1_R1117_U29);
  not ginst882 (P1_R1117_U24, P1_U3456);
  nand ginst883 (P1_R1117_U240, P1_R1117_U52, P1_U3491);
  nand ginst884 (P1_R1117_U241, P1_R1117_U50, P1_U3063);
  nand ginst885 (P1_R1117_U242, P1_R1117_U51, P1_U3062);
  nand ginst886 (P1_R1117_U243, P1_R1117_U189, P1_R1117_U8);
  nand ginst887 (P1_R1117_U244, P1_R1117_U243, P1_R1117_U9);
  nand ginst888 (P1_R1117_U245, P1_R1117_U52, P1_U3491);
  nand ginst889 (P1_R1117_U246, P1_R1117_U125, P1_R1117_U148);
  nand ginst890 (P1_R1117_U247, P1_R1117_U244, P1_R1117_U245);
  not ginst891 (P1_R1117_U248, P1_R1117_U173);
  nand ginst892 (P1_R1117_U249, P1_R1117_U56, P1_U3494);
  nand ginst893 (P1_R1117_U25, P1_R1117_U93, P1_U3456);
  nand ginst894 (P1_R1117_U250, P1_R1117_U173, P1_R1117_U249);
  nand ginst895 (P1_R1117_U251, P1_R1117_U55, P1_U3072);
  not ginst896 (P1_R1117_U252, P1_R1117_U172);
  nand ginst897 (P1_R1117_U253, P1_R1117_U58, P1_U3497);
  nand ginst898 (P1_R1117_U254, P1_R1117_U172, P1_R1117_U253);
  nand ginst899 (P1_R1117_U255, P1_R1117_U57, P1_U3080);
  not ginst900 (P1_R1117_U256, P1_R1117_U171);
  nand ginst901 (P1_R1117_U257, P1_R1117_U61, P1_U3506);
  nand ginst902 (P1_R1117_U258, P1_R1117_U59, P1_U3073);
  nand ginst903 (P1_R1117_U259, P1_R1117_U49, P1_U3074);
  not ginst904 (P1_R1117_U26, P1_U3078);
  nand ginst905 (P1_R1117_U260, P1_R1117_U180, P1_R1117_U186);
  nand ginst906 (P1_R1117_U261, P1_R1117_U10, P1_R1117_U260);
  nand ginst907 (P1_R1117_U262, P1_R1117_U63, P1_U3500);
  nand ginst908 (P1_R1117_U263, P1_R1117_U61, P1_U3506);
  nand ginst909 (P1_R1117_U264, P1_R1117_U126, P1_R1117_U171, P1_R1117_U257);
  nand ginst910 (P1_R1117_U265, P1_R1117_U261, P1_R1117_U263);
  not ginst911 (P1_R1117_U266, P1_R1117_U168);
  nand ginst912 (P1_R1117_U267, P1_R1117_U66, P1_U3509);
  nand ginst913 (P1_R1117_U268, P1_R1117_U168, P1_R1117_U267);
  nand ginst914 (P1_R1117_U269, P1_R1117_U65, P1_U3069);
  not ginst915 (P1_R1117_U27, P1_U3467);
  not ginst916 (P1_R1117_U270, P1_R1117_U67);
  nand ginst917 (P1_R1117_U271, P1_R1117_U270, P1_R1117_U68);
  nand ginst918 (P1_R1117_U272, P1_R1117_U167, P1_R1117_U271);
  nand ginst919 (P1_R1117_U273, P1_R1117_U67, P1_U3082);
  not ginst920 (P1_R1117_U274, P1_R1117_U166);
  nand ginst921 (P1_R1117_U275, P1_R1117_U70, P1_U3514);
  nand ginst922 (P1_R1117_U276, P1_R1117_U166, P1_R1117_U275);
  nand ginst923 (P1_R1117_U277, P1_R1117_U69, P1_U3081);
  not ginst924 (P1_R1117_U278, P1_R1117_U164);
  nand ginst925 (P1_R1117_U279, P1_R1117_U72, P1_U4025);
  not ginst926 (P1_R1117_U28, P1_U3068);
  nand ginst927 (P1_R1117_U280, P1_R1117_U164, P1_R1117_U279);
  nand ginst928 (P1_R1117_U281, P1_R1117_U71, P1_U3076);
  not ginst929 (P1_R1117_U282, P1_R1117_U163);
  nand ginst930 (P1_R1117_U283, P1_R1117_U75, P1_U4022);
  nand ginst931 (P1_R1117_U284, P1_R1117_U73, P1_U3066);
  nand ginst932 (P1_R1117_U285, P1_R1117_U48, P1_U3061);
  nand ginst933 (P1_R1117_U286, P1_R1117_U181, P1_R1117_U187);
  nand ginst934 (P1_R1117_U287, P1_R1117_U11, P1_R1117_U286);
  nand ginst935 (P1_R1117_U288, P1_R1117_U77, P1_U4024);
  nand ginst936 (P1_R1117_U289, P1_R1117_U75, P1_U4022);
  nand ginst937 (P1_R1117_U29, P1_R1117_U23, P1_U3068);
  nand ginst938 (P1_R1117_U290, P1_R1117_U127, P1_R1117_U163, P1_R1117_U283);
  nand ginst939 (P1_R1117_U291, P1_R1117_U287, P1_R1117_U289);
  not ginst940 (P1_R1117_U292, P1_R1117_U160);
  nand ginst941 (P1_R1117_U293, P1_R1117_U80, P1_U4021);
  nand ginst942 (P1_R1117_U294, P1_R1117_U160, P1_R1117_U293);
  nand ginst943 (P1_R1117_U295, P1_R1117_U79, P1_U3065);
  not ginst944 (P1_R1117_U296, P1_R1117_U159);
  nand ginst945 (P1_R1117_U297, P1_R1117_U82, P1_U4020);
  nand ginst946 (P1_R1117_U298, P1_R1117_U159, P1_R1117_U297);
  nand ginst947 (P1_R1117_U299, P1_R1117_U81, P1_U3058);
  not ginst948 (P1_R1117_U30, P1_U3064);
  not ginst949 (P1_R1117_U300, P1_R1117_U89);
  nand ginst950 (P1_R1117_U301, P1_R1117_U86, P1_U4018);
  nand ginst951 (P1_R1117_U302, P1_R1117_U182, P1_R1117_U301, P1_R1117_U89);
  nand ginst952 (P1_R1117_U303, P1_R1117_U85, P1_R1117_U86);
  nand ginst953 (P1_R1117_U304, P1_R1117_U303, P1_R1117_U83);
  nand ginst954 (P1_R1117_U305, P1_R1117_U176, P1_U3053);
  not ginst955 (P1_R1117_U306, P1_R1117_U157);
  nand ginst956 (P1_R1117_U307, P1_R1117_U88, P1_U4017);
  nand ginst957 (P1_R1117_U308, P1_R1117_U87, P1_U3054);
  nand ginst958 (P1_R1117_U309, P1_R1117_U300, P1_R1117_U85);
  not ginst959 (P1_R1117_U31, P1_U3476);
  nand ginst960 (P1_R1117_U310, P1_R1117_U133, P1_R1117_U309);
  nand ginst961 (P1_R1117_U311, P1_R1117_U182, P1_R1117_U89);
  nand ginst962 (P1_R1117_U312, P1_R1117_U132, P1_R1117_U311);
  nand ginst963 (P1_R1117_U313, P1_R1117_U182, P1_R1117_U85);
  nand ginst964 (P1_R1117_U314, P1_R1117_U163, P1_R1117_U288);
  not ginst965 (P1_R1117_U315, P1_R1117_U90);
  nand ginst966 (P1_R1117_U316, P1_R1117_U48, P1_U3061);
  nand ginst967 (P1_R1117_U317, P1_R1117_U315, P1_R1117_U316);
  nand ginst968 (P1_R1117_U318, P1_R1117_U136, P1_R1117_U317);
  nand ginst969 (P1_R1117_U319, P1_R1117_U181, P1_R1117_U90);
  not ginst970 (P1_R1117_U32, P1_U3473);
  nand ginst971 (P1_R1117_U320, P1_R1117_U75, P1_U4022);
  nand ginst972 (P1_R1117_U321, P1_R1117_U11, P1_R1117_U319, P1_R1117_U320);
  nand ginst973 (P1_R1117_U322, P1_R1117_U48, P1_U3061);
  nand ginst974 (P1_R1117_U323, P1_R1117_U181, P1_R1117_U322);
  nand ginst975 (P1_R1117_U324, P1_R1117_U288, P1_R1117_U78);
  nand ginst976 (P1_R1117_U325, P1_R1117_U171, P1_R1117_U262);
  not ginst977 (P1_R1117_U326, P1_R1117_U91);
  nand ginst978 (P1_R1117_U327, P1_R1117_U49, P1_U3074);
  nand ginst979 (P1_R1117_U328, P1_R1117_U326, P1_R1117_U327);
  nand ginst980 (P1_R1117_U329, P1_R1117_U142, P1_R1117_U328);
  not ginst981 (P1_R1117_U33, P1_U3470);
  nand ginst982 (P1_R1117_U330, P1_R1117_U180, P1_R1117_U91);
  nand ginst983 (P1_R1117_U331, P1_R1117_U61, P1_U3506);
  nand ginst984 (P1_R1117_U332, P1_R1117_U10, P1_R1117_U330, P1_R1117_U331);
  nand ginst985 (P1_R1117_U333, P1_R1117_U49, P1_U3074);
  nand ginst986 (P1_R1117_U334, P1_R1117_U180, P1_R1117_U333);
  nand ginst987 (P1_R1117_U335, P1_R1117_U262, P1_R1117_U64);
  nand ginst988 (P1_R1117_U336, P1_R1117_U148, P1_R1117_U217);
  not ginst989 (P1_R1117_U337, P1_R1117_U92);
  nand ginst990 (P1_R1117_U338, P1_R1117_U51, P1_U3062);
  nand ginst991 (P1_R1117_U339, P1_R1117_U337, P1_R1117_U338);
  not ginst992 (P1_R1117_U34, P1_U3071);
  nand ginst993 (P1_R1117_U340, P1_R1117_U146, P1_R1117_U339);
  nand ginst994 (P1_R1117_U341, P1_R1117_U179, P1_R1117_U92);
  nand ginst995 (P1_R1117_U342, P1_R1117_U52, P1_U3491);
  nand ginst996 (P1_R1117_U343, P1_R1117_U145, P1_R1117_U341);
  nand ginst997 (P1_R1117_U344, P1_R1117_U51, P1_U3062);
  nand ginst998 (P1_R1117_U345, P1_R1117_U179, P1_R1117_U344);
  nand ginst999 (P1_R1117_U346, P1_R1117_U24, P1_U3077);
  nand ginst1000 (P1_R1117_U347, P1_R1117_U182, P1_R1117_U301, P1_R1117_U89);
  nand ginst1001 (P1_R1117_U348, P1_R1117_U12, P1_R1117_U130, P1_R1117_U347);
  nand ginst1002 (P1_R1117_U349, P1_R1117_U43, P1_U3485);
  not ginst1003 (P1_R1117_U35, P1_U3067);
  nand ginst1004 (P1_R1117_U350, P1_R1117_U42, P1_U3083);
  nand ginst1005 (P1_R1117_U351, P1_R1117_U148, P1_R1117_U218);
  nand ginst1006 (P1_R1117_U352, P1_R1117_U147, P1_R1117_U216);
  nand ginst1007 (P1_R1117_U353, P1_R1117_U41, P1_U3482);
  nand ginst1008 (P1_R1117_U354, P1_R1117_U38, P1_U3084);
  nand ginst1009 (P1_R1117_U355, P1_R1117_U41, P1_U3482);
  nand ginst1010 (P1_R1117_U356, P1_R1117_U38, P1_U3084);
  nand ginst1011 (P1_R1117_U357, P1_R1117_U355, P1_R1117_U356);
  nand ginst1012 (P1_R1117_U358, P1_R1117_U39, P1_U3479);
  nand ginst1013 (P1_R1117_U359, P1_R1117_U22, P1_U3070);
  not ginst1014 (P1_R1117_U36, P1_U3060);
  nand ginst1015 (P1_R1117_U360, P1_R1117_U223, P1_R1117_U44);
  nand ginst1016 (P1_R1117_U361, P1_R1117_U149, P1_R1117_U210);
  nand ginst1017 (P1_R1117_U362, P1_R1117_U34, P1_U3476);
  nand ginst1018 (P1_R1117_U363, P1_R1117_U31, P1_U3071);
  nand ginst1019 (P1_R1117_U364, P1_R1117_U362, P1_R1117_U363);
  nand ginst1020 (P1_R1117_U365, P1_R1117_U35, P1_U3473);
  nand ginst1021 (P1_R1117_U366, P1_R1117_U32, P1_U3067);
  nand ginst1022 (P1_R1117_U367, P1_R1117_U233, P1_R1117_U45);
  nand ginst1023 (P1_R1117_U368, P1_R1117_U150, P1_R1117_U225);
  nand ginst1024 (P1_R1117_U369, P1_R1117_U36, P1_U3470);
  nand ginst1025 (P1_R1117_U37, P1_R1117_U33, P1_U3060);
  nand ginst1026 (P1_R1117_U370, P1_R1117_U33, P1_U3060);
  nand ginst1027 (P1_R1117_U371, P1_R1117_U152, P1_R1117_U234);
  nand ginst1028 (P1_R1117_U372, P1_R1117_U151, P1_R1117_U200);
  nand ginst1029 (P1_R1117_U373, P1_R1117_U30, P1_U3467);
  nand ginst1030 (P1_R1117_U374, P1_R1117_U27, P1_U3064);
  nand ginst1031 (P1_R1117_U375, P1_R1117_U30, P1_U3467);
  nand ginst1032 (P1_R1117_U376, P1_R1117_U27, P1_U3064);
  nand ginst1033 (P1_R1117_U377, P1_R1117_U375, P1_R1117_U376);
  nand ginst1034 (P1_R1117_U378, P1_R1117_U28, P1_U3464);
  nand ginst1035 (P1_R1117_U379, P1_R1117_U23, P1_U3068);
  not ginst1036 (P1_R1117_U38, P1_U3482);
  nand ginst1037 (P1_R1117_U380, P1_R1117_U239, P1_R1117_U46);
  nand ginst1038 (P1_R1117_U381, P1_R1117_U153, P1_R1117_U194);
  nand ginst1039 (P1_R1117_U382, P1_R1117_U155, P1_U4028);
  nand ginst1040 (P1_R1117_U383, P1_R1117_U154, P1_U3055);
  nand ginst1041 (P1_R1117_U384, P1_R1117_U155, P1_U4028);
  nand ginst1042 (P1_R1117_U385, P1_R1117_U154, P1_U3055);
  nand ginst1043 (P1_R1117_U386, P1_R1117_U384, P1_R1117_U385);
  nand ginst1044 (P1_R1117_U387, P1_R1117_U386, P1_R1117_U87, P1_U3054);
  nand ginst1045 (P1_R1117_U388, P1_R1117_U12, P1_R1117_U88, P1_U4017);
  nand ginst1046 (P1_R1117_U389, P1_R1117_U88, P1_U4017);
  not ginst1047 (P1_R1117_U39, P1_U3070);
  nand ginst1048 (P1_R1117_U390, P1_R1117_U87, P1_U3054);
  not ginst1049 (P1_R1117_U391, P1_R1117_U131);
  nand ginst1050 (P1_R1117_U392, P1_R1117_U306, P1_R1117_U391);
  nand ginst1051 (P1_R1117_U393, P1_R1117_U131, P1_R1117_U157);
  nand ginst1052 (P1_R1117_U394, P1_R1117_U86, P1_U4018);
  nand ginst1053 (P1_R1117_U395, P1_R1117_U83, P1_U3053);
  nand ginst1054 (P1_R1117_U396, P1_R1117_U86, P1_U4018);
  nand ginst1055 (P1_R1117_U397, P1_R1117_U83, P1_U3053);
  nand ginst1056 (P1_R1117_U398, P1_R1117_U396, P1_R1117_U397);
  nand ginst1057 (P1_R1117_U399, P1_R1117_U84, P1_U4019);
  nand ginst1058 (P1_R1117_U40, P1_R1117_U22, P1_U3070);
  nand ginst1059 (P1_R1117_U400, P1_R1117_U47, P1_U3057);
  nand ginst1060 (P1_R1117_U401, P1_R1117_U313, P1_R1117_U89);
  nand ginst1061 (P1_R1117_U402, P1_R1117_U158, P1_R1117_U300);
  nand ginst1062 (P1_R1117_U403, P1_R1117_U82, P1_U4020);
  nand ginst1063 (P1_R1117_U404, P1_R1117_U81, P1_U3058);
  not ginst1064 (P1_R1117_U405, P1_R1117_U134);
  nand ginst1065 (P1_R1117_U406, P1_R1117_U296, P1_R1117_U405);
  nand ginst1066 (P1_R1117_U407, P1_R1117_U134, P1_R1117_U159);
  nand ginst1067 (P1_R1117_U408, P1_R1117_U80, P1_U4021);
  nand ginst1068 (P1_R1117_U409, P1_R1117_U79, P1_U3065);
  not ginst1069 (P1_R1117_U41, P1_U3084);
  not ginst1070 (P1_R1117_U410, P1_R1117_U135);
  nand ginst1071 (P1_R1117_U411, P1_R1117_U292, P1_R1117_U410);
  nand ginst1072 (P1_R1117_U412, P1_R1117_U135, P1_R1117_U160);
  nand ginst1073 (P1_R1117_U413, P1_R1117_U75, P1_U4022);
  nand ginst1074 (P1_R1117_U414, P1_R1117_U73, P1_U3066);
  nand ginst1075 (P1_R1117_U415, P1_R1117_U413, P1_R1117_U414);
  nand ginst1076 (P1_R1117_U416, P1_R1117_U76, P1_U4023);
  nand ginst1077 (P1_R1117_U417, P1_R1117_U48, P1_U3061);
  nand ginst1078 (P1_R1117_U418, P1_R1117_U323, P1_R1117_U90);
  nand ginst1079 (P1_R1117_U419, P1_R1117_U161, P1_R1117_U315);
  not ginst1080 (P1_R1117_U42, P1_U3485);
  nand ginst1081 (P1_R1117_U420, P1_R1117_U77, P1_U4024);
  nand ginst1082 (P1_R1117_U421, P1_R1117_U74, P1_U3075);
  nand ginst1083 (P1_R1117_U422, P1_R1117_U163, P1_R1117_U324);
  nand ginst1084 (P1_R1117_U423, P1_R1117_U162, P1_R1117_U282);
  nand ginst1085 (P1_R1117_U424, P1_R1117_U72, P1_U4025);
  nand ginst1086 (P1_R1117_U425, P1_R1117_U71, P1_U3076);
  not ginst1087 (P1_R1117_U426, P1_R1117_U137);
  nand ginst1088 (P1_R1117_U427, P1_R1117_U278, P1_R1117_U426);
  nand ginst1089 (P1_R1117_U428, P1_R1117_U137, P1_R1117_U164);
  nand ginst1090 (P1_R1117_U429, P1_R1117_U26, P1_U3461);
  not ginst1091 (P1_R1117_U43, P1_U3083);
  nand ginst1092 (P1_R1117_U430, P1_R1117_U165, P1_U3078);
  not ginst1093 (P1_R1117_U431, P1_R1117_U138);
  nand ginst1094 (P1_R1117_U432, P1_R1117_U190, P1_R1117_U431);
  nand ginst1095 (P1_R1117_U433, P1_R1117_U138, P1_R1117_U25);
  nand ginst1096 (P1_R1117_U434, P1_R1117_U70, P1_U3514);
  nand ginst1097 (P1_R1117_U435, P1_R1117_U69, P1_U3081);
  not ginst1098 (P1_R1117_U436, P1_R1117_U139);
  nand ginst1099 (P1_R1117_U437, P1_R1117_U274, P1_R1117_U436);
  nand ginst1100 (P1_R1117_U438, P1_R1117_U139, P1_R1117_U166);
  nand ginst1101 (P1_R1117_U439, P1_R1117_U68, P1_U3512);
  nand ginst1102 (P1_R1117_U44, P1_R1117_U208, P1_R1117_U209);
  nand ginst1103 (P1_R1117_U440, P1_R1117_U167, P1_U3082);
  not ginst1104 (P1_R1117_U441, P1_R1117_U140);
  nand ginst1105 (P1_R1117_U442, P1_R1117_U270, P1_R1117_U441);
  nand ginst1106 (P1_R1117_U443, P1_R1117_U140, P1_R1117_U67);
  nand ginst1107 (P1_R1117_U444, P1_R1117_U66, P1_U3509);
  nand ginst1108 (P1_R1117_U445, P1_R1117_U65, P1_U3069);
  not ginst1109 (P1_R1117_U446, P1_R1117_U141);
  nand ginst1110 (P1_R1117_U447, P1_R1117_U266, P1_R1117_U446);
  nand ginst1111 (P1_R1117_U448, P1_R1117_U141, P1_R1117_U168);
  nand ginst1112 (P1_R1117_U449, P1_R1117_U61, P1_U3506);
  nand ginst1113 (P1_R1117_U45, P1_R1117_U224, P1_R1117_U37);
  nand ginst1114 (P1_R1117_U450, P1_R1117_U59, P1_U3073);
  nand ginst1115 (P1_R1117_U451, P1_R1117_U449, P1_R1117_U450);
  nand ginst1116 (P1_R1117_U452, P1_R1117_U62, P1_U3503);
  nand ginst1117 (P1_R1117_U453, P1_R1117_U49, P1_U3074);
  nand ginst1118 (P1_R1117_U454, P1_R1117_U334, P1_R1117_U91);
  nand ginst1119 (P1_R1117_U455, P1_R1117_U169, P1_R1117_U326);
  nand ginst1120 (P1_R1117_U456, P1_R1117_U63, P1_U3500);
  nand ginst1121 (P1_R1117_U457, P1_R1117_U60, P1_U3079);
  nand ginst1122 (P1_R1117_U458, P1_R1117_U171, P1_R1117_U335);
  nand ginst1123 (P1_R1117_U459, P1_R1117_U170, P1_R1117_U256);
  nand ginst1124 (P1_R1117_U46, P1_R1117_U192, P1_R1117_U193);
  nand ginst1125 (P1_R1117_U460, P1_R1117_U58, P1_U3497);
  nand ginst1126 (P1_R1117_U461, P1_R1117_U57, P1_U3080);
  not ginst1127 (P1_R1117_U462, P1_R1117_U143);
  nand ginst1128 (P1_R1117_U463, P1_R1117_U252, P1_R1117_U462);
  nand ginst1129 (P1_R1117_U464, P1_R1117_U143, P1_R1117_U172);
  nand ginst1130 (P1_R1117_U465, P1_R1117_U56, P1_U3494);
  nand ginst1131 (P1_R1117_U466, P1_R1117_U55, P1_U3072);
  not ginst1132 (P1_R1117_U467, P1_R1117_U144);
  nand ginst1133 (P1_R1117_U468, P1_R1117_U248, P1_R1117_U467);
  nand ginst1134 (P1_R1117_U469, P1_R1117_U144, P1_R1117_U173);
  not ginst1135 (P1_R1117_U47, P1_U4019);
  nand ginst1136 (P1_R1117_U470, P1_R1117_U52, P1_U3491);
  nand ginst1137 (P1_R1117_U471, P1_R1117_U50, P1_U3063);
  nand ginst1138 (P1_R1117_U472, P1_R1117_U470, P1_R1117_U471);
  nand ginst1139 (P1_R1117_U473, P1_R1117_U53, P1_U3488);
  nand ginst1140 (P1_R1117_U474, P1_R1117_U51, P1_U3062);
  nand ginst1141 (P1_R1117_U475, P1_R1117_U345, P1_R1117_U92);
  nand ginst1142 (P1_R1117_U476, P1_R1117_U174, P1_R1117_U337);
  not ginst1143 (P1_R1117_U48, P1_U4023);
  not ginst1144 (P1_R1117_U49, P1_U3503);
  not ginst1145 (P1_R1117_U50, P1_U3491);
  not ginst1146 (P1_R1117_U51, P1_U3488);
  not ginst1147 (P1_R1117_U52, P1_U3063);
  not ginst1148 (P1_R1117_U53, P1_U3062);
  nand ginst1149 (P1_R1117_U54, P1_R1117_U42, P1_U3083);
  not ginst1150 (P1_R1117_U55, P1_U3494);
  not ginst1151 (P1_R1117_U56, P1_U3072);
  not ginst1152 (P1_R1117_U57, P1_U3497);
  not ginst1153 (P1_R1117_U58, P1_U3080);
  not ginst1154 (P1_R1117_U59, P1_U3506);
  and ginst1155 (P1_R1117_U6, P1_R1117_U184, P1_R1117_U201);
  not ginst1156 (P1_R1117_U60, P1_U3500);
  not ginst1157 (P1_R1117_U61, P1_U3073);
  not ginst1158 (P1_R1117_U62, P1_U3074);
  not ginst1159 (P1_R1117_U63, P1_U3079);
  nand ginst1160 (P1_R1117_U64, P1_R1117_U60, P1_U3079);
  not ginst1161 (P1_R1117_U65, P1_U3509);
  not ginst1162 (P1_R1117_U66, P1_U3069);
  nand ginst1163 (P1_R1117_U67, P1_R1117_U268, P1_R1117_U269);
  not ginst1164 (P1_R1117_U68, P1_U3082);
  not ginst1165 (P1_R1117_U69, P1_U3514);
  and ginst1166 (P1_R1117_U7, P1_R1117_U202, P1_R1117_U203);
  not ginst1167 (P1_R1117_U70, P1_U3081);
  not ginst1168 (P1_R1117_U71, P1_U4025);
  not ginst1169 (P1_R1117_U72, P1_U3076);
  not ginst1170 (P1_R1117_U73, P1_U4022);
  not ginst1171 (P1_R1117_U74, P1_U4024);
  not ginst1172 (P1_R1117_U75, P1_U3066);
  not ginst1173 (P1_R1117_U76, P1_U3061);
  not ginst1174 (P1_R1117_U77, P1_U3075);
  nand ginst1175 (P1_R1117_U78, P1_R1117_U74, P1_U3075);
  not ginst1176 (P1_R1117_U79, P1_U4021);
  and ginst1177 (P1_R1117_U8, P1_R1117_U179, P1_R1117_U240);
  not ginst1178 (P1_R1117_U80, P1_U3065);
  not ginst1179 (P1_R1117_U81, P1_U4020);
  not ginst1180 (P1_R1117_U82, P1_U3058);
  not ginst1181 (P1_R1117_U83, P1_U4018);
  not ginst1182 (P1_R1117_U84, P1_U3057);
  nand ginst1183 (P1_R1117_U85, P1_R1117_U47, P1_U3057);
  not ginst1184 (P1_R1117_U86, P1_U3053);
  not ginst1185 (P1_R1117_U87, P1_U4017);
  not ginst1186 (P1_R1117_U88, P1_U3054);
  nand ginst1187 (P1_R1117_U89, P1_R1117_U298, P1_R1117_U299);
  and ginst1188 (P1_R1117_U9, P1_R1117_U241, P1_R1117_U242);
  nand ginst1189 (P1_R1117_U90, P1_R1117_U314, P1_R1117_U78);
  nand ginst1190 (P1_R1117_U91, P1_R1117_U325, P1_R1117_U64);
  nand ginst1191 (P1_R1117_U92, P1_R1117_U336, P1_R1117_U54);
  not ginst1192 (P1_R1117_U93, P1_U3077);
  nand ginst1193 (P1_R1117_U94, P1_R1117_U392, P1_R1117_U393);
  nand ginst1194 (P1_R1117_U95, P1_R1117_U406, P1_R1117_U407);
  nand ginst1195 (P1_R1117_U96, P1_R1117_U411, P1_R1117_U412);
  nand ginst1196 (P1_R1117_U97, P1_R1117_U427, P1_R1117_U428);
  nand ginst1197 (P1_R1117_U98, P1_R1117_U432, P1_R1117_U433);
  nand ginst1198 (P1_R1117_U99, P1_R1117_U437, P1_R1117_U438);
  and ginst1199 (P1_R1138_U10, P1_R1138_U268, P1_R1138_U269);
  nand ginst1200 (P1_R1138_U100, P1_R1138_U390, P1_R1138_U391);
  nand ginst1201 (P1_R1138_U101, P1_R1138_U395, P1_R1138_U396);
  nand ginst1202 (P1_R1138_U102, P1_R1138_U404, P1_R1138_U405);
  nand ginst1203 (P1_R1138_U103, P1_R1138_U411, P1_R1138_U412);
  nand ginst1204 (P1_R1138_U104, P1_R1138_U418, P1_R1138_U419);
  nand ginst1205 (P1_R1138_U105, P1_R1138_U425, P1_R1138_U426);
  nand ginst1206 (P1_R1138_U106, P1_R1138_U430, P1_R1138_U431);
  nand ginst1207 (P1_R1138_U107, P1_R1138_U437, P1_R1138_U438);
  nand ginst1208 (P1_R1138_U108, P1_R1138_U444, P1_R1138_U445);
  nand ginst1209 (P1_R1138_U109, P1_R1138_U458, P1_R1138_U459);
  and ginst1210 (P1_R1138_U11, P1_R1138_U345, P1_R1138_U348);
  nand ginst1211 (P1_R1138_U110, P1_R1138_U463, P1_R1138_U464);
  nand ginst1212 (P1_R1138_U111, P1_R1138_U470, P1_R1138_U471);
  nand ginst1213 (P1_R1138_U112, P1_R1138_U477, P1_R1138_U478);
  nand ginst1214 (P1_R1138_U113, P1_R1138_U484, P1_R1138_U485);
  nand ginst1215 (P1_R1138_U114, P1_R1138_U491, P1_R1138_U492);
  nand ginst1216 (P1_R1138_U115, P1_R1138_U496, P1_R1138_U497);
  and ginst1217 (P1_R1138_U116, P1_U3068, P1_U3464);
  and ginst1218 (P1_R1138_U117, P1_R1138_U184, P1_R1138_U186);
  and ginst1219 (P1_R1138_U118, P1_R1138_U189, P1_R1138_U191);
  and ginst1220 (P1_R1138_U119, P1_R1138_U197, P1_R1138_U198);
  and ginst1221 (P1_R1138_U12, P1_R1138_U338, P1_R1138_U341);
  and ginst1222 (P1_R1138_U120, P1_R1138_U23, P1_R1138_U378, P1_R1138_U379);
  and ginst1223 (P1_R1138_U121, P1_R1138_U209, P1_R1138_U6);
  and ginst1224 (P1_R1138_U122, P1_R1138_U215, P1_R1138_U217);
  and ginst1225 (P1_R1138_U123, P1_R1138_U35, P1_R1138_U385, P1_R1138_U386);
  and ginst1226 (P1_R1138_U124, P1_R1138_U223, P1_R1138_U4);
  and ginst1227 (P1_R1138_U125, P1_R1138_U178, P1_R1138_U231);
  and ginst1228 (P1_R1138_U126, P1_R1138_U201, P1_R1138_U7);
  and ginst1229 (P1_R1138_U127, P1_R1138_U168, P1_R1138_U236);
  and ginst1230 (P1_R1138_U128, P1_R1138_U169, P1_R1138_U245);
  and ginst1231 (P1_R1138_U129, P1_R1138_U264, P1_R1138_U265);
  and ginst1232 (P1_R1138_U13, P1_R1138_U329, P1_R1138_U332);
  and ginst1233 (P1_R1138_U130, P1_R1138_U10, P1_R1138_U279);
  and ginst1234 (P1_R1138_U131, P1_R1138_U277, P1_R1138_U282);
  and ginst1235 (P1_R1138_U132, P1_R1138_U295, P1_R1138_U298);
  and ginst1236 (P1_R1138_U133, P1_R1138_U299, P1_R1138_U365);
  and ginst1237 (P1_R1138_U134, P1_R1138_U156, P1_R1138_U275);
  and ginst1238 (P1_R1138_U135, P1_R1138_U465, P1_R1138_U466, P1_R1138_U60);
  and ginst1239 (P1_R1138_U136, P1_R1138_U169, P1_R1138_U486, P1_R1138_U487);
  and ginst1240 (P1_R1138_U137, P1_R1138_U340, P1_R1138_U8);
  and ginst1241 (P1_R1138_U138, P1_R1138_U168, P1_R1138_U498, P1_R1138_U499);
  and ginst1242 (P1_R1138_U139, P1_R1138_U347, P1_R1138_U7);
  and ginst1243 (P1_R1138_U14, P1_R1138_U320, P1_R1138_U323);
  nand ginst1244 (P1_R1138_U140, P1_R1138_U119, P1_R1138_U199);
  nand ginst1245 (P1_R1138_U141, P1_R1138_U214, P1_R1138_U226);
  not ginst1246 (P1_R1138_U142, P1_U3055);
  not ginst1247 (P1_R1138_U143, P1_U4028);
  and ginst1248 (P1_R1138_U144, P1_R1138_U399, P1_R1138_U400);
  nand ginst1249 (P1_R1138_U145, P1_R1138_U166, P1_R1138_U301, P1_R1138_U361);
  and ginst1250 (P1_R1138_U146, P1_R1138_U406, P1_R1138_U407);
  nand ginst1251 (P1_R1138_U147, P1_R1138_U133, P1_R1138_U366, P1_R1138_U367);
  and ginst1252 (P1_R1138_U148, P1_R1138_U413, P1_R1138_U414);
  nand ginst1253 (P1_R1138_U149, P1_R1138_U296, P1_R1138_U362, P1_R1138_U87);
  and ginst1254 (P1_R1138_U15, P1_R1138_U315, P1_R1138_U317);
  and ginst1255 (P1_R1138_U150, P1_R1138_U420, P1_R1138_U421);
  nand ginst1256 (P1_R1138_U151, P1_R1138_U289, P1_R1138_U290);
  and ginst1257 (P1_R1138_U152, P1_R1138_U432, P1_R1138_U433);
  nand ginst1258 (P1_R1138_U153, P1_R1138_U285, P1_R1138_U286);
  and ginst1259 (P1_R1138_U154, P1_R1138_U439, P1_R1138_U440);
  nand ginst1260 (P1_R1138_U155, P1_R1138_U131, P1_R1138_U281);
  and ginst1261 (P1_R1138_U156, P1_R1138_U446, P1_R1138_U447);
  and ginst1262 (P1_R1138_U157, P1_R1138_U451, P1_R1138_U452);
  nand ginst1263 (P1_R1138_U158, P1_R1138_U324, P1_R1138_U44);
  nand ginst1264 (P1_R1138_U159, P1_R1138_U129, P1_R1138_U266);
  and ginst1265 (P1_R1138_U16, P1_R1138_U307, P1_R1138_U310);
  and ginst1266 (P1_R1138_U160, P1_R1138_U472, P1_R1138_U473);
  nand ginst1267 (P1_R1138_U161, P1_R1138_U253, P1_R1138_U254);
  and ginst1268 (P1_R1138_U162, P1_R1138_U479, P1_R1138_U480);
  nand ginst1269 (P1_R1138_U163, P1_R1138_U249, P1_R1138_U250);
  nand ginst1270 (P1_R1138_U164, P1_R1138_U239, P1_R1138_U240);
  nand ginst1271 (P1_R1138_U165, P1_R1138_U363, P1_R1138_U364);
  nand ginst1272 (P1_R1138_U166, P1_R1138_U147, P1_U3054);
  not ginst1273 (P1_R1138_U167, P1_R1138_U35);
  nand ginst1274 (P1_R1138_U168, P1_U3083, P1_U3485);
  nand ginst1275 (P1_R1138_U169, P1_U3072, P1_U3494);
  and ginst1276 (P1_R1138_U17, P1_R1138_U229, P1_R1138_U232);
  nand ginst1277 (P1_R1138_U170, P1_U3058, P1_U4020);
  not ginst1278 (P1_R1138_U171, P1_R1138_U69);
  not ginst1279 (P1_R1138_U172, P1_R1138_U78);
  nand ginst1280 (P1_R1138_U173, P1_U3065, P1_U4021);
  not ginst1281 (P1_R1138_U174, P1_R1138_U62);
  or ginst1282 (P1_R1138_U175, P1_U3067, P1_U3473);
  or ginst1283 (P1_R1138_U176, P1_U3060, P1_U3470);
  or ginst1284 (P1_R1138_U177, P1_U3064, P1_U3467);
  or ginst1285 (P1_R1138_U178, P1_U3068, P1_U3464);
  not ginst1286 (P1_R1138_U179, P1_R1138_U32);
  and ginst1287 (P1_R1138_U18, P1_R1138_U221, P1_R1138_U224);
  or ginst1288 (P1_R1138_U180, P1_U3078, P1_U3461);
  not ginst1289 (P1_R1138_U181, P1_R1138_U43);
  not ginst1290 (P1_R1138_U182, P1_R1138_U44);
  nand ginst1291 (P1_R1138_U183, P1_R1138_U43, P1_R1138_U44);
  nand ginst1292 (P1_R1138_U184, P1_R1138_U116, P1_R1138_U177);
  nand ginst1293 (P1_R1138_U185, P1_R1138_U183, P1_R1138_U5);
  nand ginst1294 (P1_R1138_U186, P1_U3064, P1_U3467);
  nand ginst1295 (P1_R1138_U187, P1_R1138_U117, P1_R1138_U185);
  nand ginst1296 (P1_R1138_U188, P1_R1138_U35, P1_R1138_U36);
  nand ginst1297 (P1_R1138_U189, P1_R1138_U188, P1_U3067);
  and ginst1298 (P1_R1138_U19, P1_R1138_U207, P1_R1138_U210);
  nand ginst1299 (P1_R1138_U190, P1_R1138_U187, P1_R1138_U4);
  nand ginst1300 (P1_R1138_U191, P1_R1138_U167, P1_U3473);
  not ginst1301 (P1_R1138_U192, P1_R1138_U42);
  or ginst1302 (P1_R1138_U193, P1_U3070, P1_U3479);
  or ginst1303 (P1_R1138_U194, P1_U3071, P1_U3476);
  not ginst1304 (P1_R1138_U195, P1_R1138_U23);
  nand ginst1305 (P1_R1138_U196, P1_R1138_U23, P1_R1138_U24);
  nand ginst1306 (P1_R1138_U197, P1_R1138_U196, P1_U3070);
  nand ginst1307 (P1_R1138_U198, P1_R1138_U195, P1_U3479);
  nand ginst1308 (P1_R1138_U199, P1_R1138_U42, P1_R1138_U6);
  not ginst1309 (P1_R1138_U20, P1_U3476);
  not ginst1310 (P1_R1138_U200, P1_R1138_U140);
  or ginst1311 (P1_R1138_U201, P1_U3084, P1_U3482);
  nand ginst1312 (P1_R1138_U202, P1_R1138_U140, P1_R1138_U201);
  not ginst1313 (P1_R1138_U203, P1_R1138_U41);
  or ginst1314 (P1_R1138_U204, P1_U3083, P1_U3485);
  or ginst1315 (P1_R1138_U205, P1_U3071, P1_U3476);
  nand ginst1316 (P1_R1138_U206, P1_R1138_U205, P1_R1138_U42);
  nand ginst1317 (P1_R1138_U207, P1_R1138_U120, P1_R1138_U206);
  nand ginst1318 (P1_R1138_U208, P1_R1138_U192, P1_R1138_U23);
  nand ginst1319 (P1_R1138_U209, P1_U3070, P1_U3479);
  not ginst1320 (P1_R1138_U21, P1_U3071);
  nand ginst1321 (P1_R1138_U210, P1_R1138_U121, P1_R1138_U208);
  or ginst1322 (P1_R1138_U211, P1_U3071, P1_U3476);
  nand ginst1323 (P1_R1138_U212, P1_R1138_U178, P1_R1138_U182);
  nand ginst1324 (P1_R1138_U213, P1_U3068, P1_U3464);
  not ginst1325 (P1_R1138_U214, P1_R1138_U46);
  nand ginst1326 (P1_R1138_U215, P1_R1138_U181, P1_R1138_U5);
  nand ginst1327 (P1_R1138_U216, P1_R1138_U177, P1_R1138_U46);
  nand ginst1328 (P1_R1138_U217, P1_U3064, P1_U3467);
  not ginst1329 (P1_R1138_U218, P1_R1138_U45);
  or ginst1330 (P1_R1138_U219, P1_U3060, P1_U3470);
  not ginst1331 (P1_R1138_U22, P1_U3070);
  nand ginst1332 (P1_R1138_U220, P1_R1138_U219, P1_R1138_U45);
  nand ginst1333 (P1_R1138_U221, P1_R1138_U123, P1_R1138_U220);
  nand ginst1334 (P1_R1138_U222, P1_R1138_U218, P1_R1138_U35);
  nand ginst1335 (P1_R1138_U223, P1_U3067, P1_U3473);
  nand ginst1336 (P1_R1138_U224, P1_R1138_U124, P1_R1138_U222);
  or ginst1337 (P1_R1138_U225, P1_U3060, P1_U3470);
  nand ginst1338 (P1_R1138_U226, P1_R1138_U178, P1_R1138_U181);
  not ginst1339 (P1_R1138_U227, P1_R1138_U141);
  nand ginst1340 (P1_R1138_U228, P1_U3064, P1_U3467);
  nand ginst1341 (P1_R1138_U229, P1_R1138_U397, P1_R1138_U398, P1_R1138_U43, P1_R1138_U44);
  nand ginst1342 (P1_R1138_U23, P1_U3071, P1_U3476);
  nand ginst1343 (P1_R1138_U230, P1_R1138_U43, P1_R1138_U44);
  nand ginst1344 (P1_R1138_U231, P1_U3068, P1_U3464);
  nand ginst1345 (P1_R1138_U232, P1_R1138_U125, P1_R1138_U230);
  or ginst1346 (P1_R1138_U233, P1_U3083, P1_U3485);
  or ginst1347 (P1_R1138_U234, P1_U3062, P1_U3488);
  nand ginst1348 (P1_R1138_U235, P1_R1138_U174, P1_R1138_U7);
  nand ginst1349 (P1_R1138_U236, P1_U3062, P1_U3488);
  nand ginst1350 (P1_R1138_U237, P1_R1138_U127, P1_R1138_U235);
  or ginst1351 (P1_R1138_U238, P1_U3062, P1_U3488);
  nand ginst1352 (P1_R1138_U239, P1_R1138_U126, P1_R1138_U140);
  not ginst1353 (P1_R1138_U24, P1_U3479);
  nand ginst1354 (P1_R1138_U240, P1_R1138_U237, P1_R1138_U238);
  not ginst1355 (P1_R1138_U241, P1_R1138_U164);
  or ginst1356 (P1_R1138_U242, P1_U3080, P1_U3497);
  or ginst1357 (P1_R1138_U243, P1_U3072, P1_U3494);
  nand ginst1358 (P1_R1138_U244, P1_R1138_U171, P1_R1138_U8);
  nand ginst1359 (P1_R1138_U245, P1_U3080, P1_U3497);
  nand ginst1360 (P1_R1138_U246, P1_R1138_U128, P1_R1138_U244);
  or ginst1361 (P1_R1138_U247, P1_U3063, P1_U3491);
  or ginst1362 (P1_R1138_U248, P1_U3080, P1_U3497);
  nand ginst1363 (P1_R1138_U249, P1_R1138_U164, P1_R1138_U247, P1_R1138_U8);
  not ginst1364 (P1_R1138_U25, P1_U3470);
  nand ginst1365 (P1_R1138_U250, P1_R1138_U246, P1_R1138_U248);
  not ginst1366 (P1_R1138_U251, P1_R1138_U163);
  or ginst1367 (P1_R1138_U252, P1_U3079, P1_U3500);
  nand ginst1368 (P1_R1138_U253, P1_R1138_U163, P1_R1138_U252);
  nand ginst1369 (P1_R1138_U254, P1_U3079, P1_U3500);
  not ginst1370 (P1_R1138_U255, P1_R1138_U161);
  or ginst1371 (P1_R1138_U256, P1_U3074, P1_U3503);
  nand ginst1372 (P1_R1138_U257, P1_R1138_U161, P1_R1138_U256);
  nand ginst1373 (P1_R1138_U258, P1_U3074, P1_U3503);
  not ginst1374 (P1_R1138_U259, P1_R1138_U93);
  not ginst1375 (P1_R1138_U26, P1_U3060);
  or ginst1376 (P1_R1138_U260, P1_U3069, P1_U3509);
  or ginst1377 (P1_R1138_U261, P1_U3073, P1_U3506);
  not ginst1378 (P1_R1138_U262, P1_R1138_U60);
  nand ginst1379 (P1_R1138_U263, P1_R1138_U60, P1_R1138_U61);
  nand ginst1380 (P1_R1138_U264, P1_R1138_U263, P1_U3069);
  nand ginst1381 (P1_R1138_U265, P1_R1138_U262, P1_U3509);
  nand ginst1382 (P1_R1138_U266, P1_R1138_U9, P1_R1138_U93);
  not ginst1383 (P1_R1138_U267, P1_R1138_U159);
  or ginst1384 (P1_R1138_U268, P1_U3076, P1_U4025);
  or ginst1385 (P1_R1138_U269, P1_U3081, P1_U3514);
  not ginst1386 (P1_R1138_U27, P1_U3067);
  or ginst1387 (P1_R1138_U270, P1_U3075, P1_U4024);
  not ginst1388 (P1_R1138_U271, P1_R1138_U81);
  nand ginst1389 (P1_R1138_U272, P1_R1138_U271, P1_U4025);
  nand ginst1390 (P1_R1138_U273, P1_R1138_U272, P1_R1138_U91);
  nand ginst1391 (P1_R1138_U274, P1_R1138_U81, P1_R1138_U82);
  nand ginst1392 (P1_R1138_U275, P1_R1138_U273, P1_R1138_U274);
  nand ginst1393 (P1_R1138_U276, P1_R1138_U10, P1_R1138_U172);
  nand ginst1394 (P1_R1138_U277, P1_U3075, P1_U4024);
  nand ginst1395 (P1_R1138_U278, P1_R1138_U275, P1_R1138_U276);
  or ginst1396 (P1_R1138_U279, P1_U3082, P1_U3512);
  not ginst1397 (P1_R1138_U28, P1_U3464);
  or ginst1398 (P1_R1138_U280, P1_U3075, P1_U4024);
  nand ginst1399 (P1_R1138_U281, P1_R1138_U130, P1_R1138_U159, P1_R1138_U270);
  nand ginst1400 (P1_R1138_U282, P1_R1138_U278, P1_R1138_U280);
  not ginst1401 (P1_R1138_U283, P1_R1138_U155);
  or ginst1402 (P1_R1138_U284, P1_U3061, P1_U4023);
  nand ginst1403 (P1_R1138_U285, P1_R1138_U155, P1_R1138_U284);
  nand ginst1404 (P1_R1138_U286, P1_U3061, P1_U4023);
  not ginst1405 (P1_R1138_U287, P1_R1138_U153);
  or ginst1406 (P1_R1138_U288, P1_U3066, P1_U4022);
  nand ginst1407 (P1_R1138_U289, P1_R1138_U153, P1_R1138_U288);
  not ginst1408 (P1_R1138_U29, P1_U3068);
  nand ginst1409 (P1_R1138_U290, P1_U3066, P1_U4022);
  not ginst1410 (P1_R1138_U291, P1_R1138_U151);
  or ginst1411 (P1_R1138_U292, P1_U3058, P1_U4020);
  nand ginst1412 (P1_R1138_U293, P1_R1138_U170, P1_R1138_U173);
  not ginst1413 (P1_R1138_U294, P1_R1138_U87);
  or ginst1414 (P1_R1138_U295, P1_U3065, P1_U4021);
  nand ginst1415 (P1_R1138_U296, P1_R1138_U151, P1_R1138_U165, P1_R1138_U295);
  not ginst1416 (P1_R1138_U297, P1_R1138_U149);
  or ginst1417 (P1_R1138_U298, P1_U3053, P1_U4018);
  nand ginst1418 (P1_R1138_U299, P1_U3053, P1_U4018);
  not ginst1419 (P1_R1138_U30, P1_U3456);
  not ginst1420 (P1_R1138_U300, P1_R1138_U147);
  nand ginst1421 (P1_R1138_U301, P1_R1138_U147, P1_U4017);
  not ginst1422 (P1_R1138_U302, P1_R1138_U145);
  nand ginst1423 (P1_R1138_U303, P1_R1138_U151, P1_R1138_U295);
  not ginst1424 (P1_R1138_U304, P1_R1138_U90);
  or ginst1425 (P1_R1138_U305, P1_U3058, P1_U4020);
  nand ginst1426 (P1_R1138_U306, P1_R1138_U305, P1_R1138_U90);
  nand ginst1427 (P1_R1138_U307, P1_R1138_U150, P1_R1138_U170, P1_R1138_U306);
  nand ginst1428 (P1_R1138_U308, P1_R1138_U170, P1_R1138_U304);
  nand ginst1429 (P1_R1138_U309, P1_U3057, P1_U4019);
  not ginst1430 (P1_R1138_U31, P1_U3077);
  nand ginst1431 (P1_R1138_U310, P1_R1138_U165, P1_R1138_U308, P1_R1138_U309);
  or ginst1432 (P1_R1138_U311, P1_U3058, P1_U4020);
  nand ginst1433 (P1_R1138_U312, P1_R1138_U159, P1_R1138_U279);
  not ginst1434 (P1_R1138_U313, P1_R1138_U92);
  nand ginst1435 (P1_R1138_U314, P1_R1138_U10, P1_R1138_U92);
  nand ginst1436 (P1_R1138_U315, P1_R1138_U134, P1_R1138_U314);
  nand ginst1437 (P1_R1138_U316, P1_R1138_U275, P1_R1138_U314);
  nand ginst1438 (P1_R1138_U317, P1_R1138_U316, P1_R1138_U450);
  or ginst1439 (P1_R1138_U318, P1_U3081, P1_U3514);
  nand ginst1440 (P1_R1138_U319, P1_R1138_U318, P1_R1138_U92);
  nand ginst1441 (P1_R1138_U32, P1_U3077, P1_U3456);
  nand ginst1442 (P1_R1138_U320, P1_R1138_U157, P1_R1138_U319, P1_R1138_U81);
  nand ginst1443 (P1_R1138_U321, P1_R1138_U313, P1_R1138_U81);
  nand ginst1444 (P1_R1138_U322, P1_U3076, P1_U4025);
  nand ginst1445 (P1_R1138_U323, P1_R1138_U10, P1_R1138_U321, P1_R1138_U322);
  or ginst1446 (P1_R1138_U324, P1_U3078, P1_U3461);
  not ginst1447 (P1_R1138_U325, P1_R1138_U158);
  or ginst1448 (P1_R1138_U326, P1_U3081, P1_U3514);
  or ginst1449 (P1_R1138_U327, P1_U3073, P1_U3506);
  nand ginst1450 (P1_R1138_U328, P1_R1138_U327, P1_R1138_U93);
  nand ginst1451 (P1_R1138_U329, P1_R1138_U135, P1_R1138_U328);
  not ginst1452 (P1_R1138_U33, P1_U3467);
  nand ginst1453 (P1_R1138_U330, P1_R1138_U259, P1_R1138_U60);
  nand ginst1454 (P1_R1138_U331, P1_U3069, P1_U3509);
  nand ginst1455 (P1_R1138_U332, P1_R1138_U330, P1_R1138_U331, P1_R1138_U9);
  or ginst1456 (P1_R1138_U333, P1_U3073, P1_U3506);
  nand ginst1457 (P1_R1138_U334, P1_R1138_U164, P1_R1138_U247);
  not ginst1458 (P1_R1138_U335, P1_R1138_U94);
  or ginst1459 (P1_R1138_U336, P1_U3072, P1_U3494);
  nand ginst1460 (P1_R1138_U337, P1_R1138_U336, P1_R1138_U94);
  nand ginst1461 (P1_R1138_U338, P1_R1138_U136, P1_R1138_U337);
  nand ginst1462 (P1_R1138_U339, P1_R1138_U169, P1_R1138_U335);
  not ginst1463 (P1_R1138_U34, P1_U3064);
  nand ginst1464 (P1_R1138_U340, P1_U3080, P1_U3497);
  nand ginst1465 (P1_R1138_U341, P1_R1138_U137, P1_R1138_U339);
  or ginst1466 (P1_R1138_U342, P1_U3072, P1_U3494);
  or ginst1467 (P1_R1138_U343, P1_U3083, P1_U3485);
  nand ginst1468 (P1_R1138_U344, P1_R1138_U343, P1_R1138_U41);
  nand ginst1469 (P1_R1138_U345, P1_R1138_U138, P1_R1138_U344);
  nand ginst1470 (P1_R1138_U346, P1_R1138_U168, P1_R1138_U203);
  nand ginst1471 (P1_R1138_U347, P1_U3062, P1_U3488);
  nand ginst1472 (P1_R1138_U348, P1_R1138_U139, P1_R1138_U346);
  nand ginst1473 (P1_R1138_U349, P1_R1138_U168, P1_R1138_U204);
  nand ginst1474 (P1_R1138_U35, P1_U3060, P1_U3470);
  nand ginst1475 (P1_R1138_U350, P1_R1138_U201, P1_R1138_U62);
  nand ginst1476 (P1_R1138_U351, P1_R1138_U211, P1_R1138_U23);
  nand ginst1477 (P1_R1138_U352, P1_R1138_U225, P1_R1138_U35);
  nand ginst1478 (P1_R1138_U353, P1_R1138_U177, P1_R1138_U228);
  nand ginst1479 (P1_R1138_U354, P1_R1138_U170, P1_R1138_U311);
  nand ginst1480 (P1_R1138_U355, P1_R1138_U173, P1_R1138_U295);
  nand ginst1481 (P1_R1138_U356, P1_R1138_U326, P1_R1138_U81);
  nand ginst1482 (P1_R1138_U357, P1_R1138_U279, P1_R1138_U78);
  nand ginst1483 (P1_R1138_U358, P1_R1138_U333, P1_R1138_U60);
  nand ginst1484 (P1_R1138_U359, P1_R1138_U169, P1_R1138_U342);
  not ginst1485 (P1_R1138_U36, P1_U3473);
  nand ginst1486 (P1_R1138_U360, P1_R1138_U247, P1_R1138_U69);
  nand ginst1487 (P1_R1138_U361, P1_U3054, P1_U4017);
  nand ginst1488 (P1_R1138_U362, P1_R1138_U165, P1_R1138_U293);
  nand ginst1489 (P1_R1138_U363, P1_R1138_U292, P1_U3057);
  nand ginst1490 (P1_R1138_U364, P1_R1138_U292, P1_U4019);
  nand ginst1491 (P1_R1138_U365, P1_R1138_U165, P1_R1138_U293, P1_R1138_U298);
  nand ginst1492 (P1_R1138_U366, P1_R1138_U132, P1_R1138_U151, P1_R1138_U165);
  nand ginst1493 (P1_R1138_U367, P1_R1138_U294, P1_R1138_U298);
  nand ginst1494 (P1_R1138_U368, P1_R1138_U40, P1_U3083);
  nand ginst1495 (P1_R1138_U369, P1_R1138_U39, P1_U3485);
  not ginst1496 (P1_R1138_U37, P1_U3482);
  nand ginst1497 (P1_R1138_U370, P1_R1138_U368, P1_R1138_U369);
  nand ginst1498 (P1_R1138_U371, P1_R1138_U349, P1_R1138_U41);
  nand ginst1499 (P1_R1138_U372, P1_R1138_U203, P1_R1138_U370);
  nand ginst1500 (P1_R1138_U373, P1_R1138_U37, P1_U3084);
  nand ginst1501 (P1_R1138_U374, P1_R1138_U38, P1_U3482);
  nand ginst1502 (P1_R1138_U375, P1_R1138_U373, P1_R1138_U374);
  nand ginst1503 (P1_R1138_U376, P1_R1138_U140, P1_R1138_U350);
  nand ginst1504 (P1_R1138_U377, P1_R1138_U200, P1_R1138_U375);
  nand ginst1505 (P1_R1138_U378, P1_R1138_U24, P1_U3070);
  nand ginst1506 (P1_R1138_U379, P1_R1138_U22, P1_U3479);
  not ginst1507 (P1_R1138_U38, P1_U3084);
  nand ginst1508 (P1_R1138_U380, P1_R1138_U20, P1_U3071);
  nand ginst1509 (P1_R1138_U381, P1_R1138_U21, P1_U3476);
  nand ginst1510 (P1_R1138_U382, P1_R1138_U380, P1_R1138_U381);
  nand ginst1511 (P1_R1138_U383, P1_R1138_U351, P1_R1138_U42);
  nand ginst1512 (P1_R1138_U384, P1_R1138_U192, P1_R1138_U382);
  nand ginst1513 (P1_R1138_U385, P1_R1138_U36, P1_U3067);
  nand ginst1514 (P1_R1138_U386, P1_R1138_U27, P1_U3473);
  nand ginst1515 (P1_R1138_U387, P1_R1138_U25, P1_U3060);
  nand ginst1516 (P1_R1138_U388, P1_R1138_U26, P1_U3470);
  nand ginst1517 (P1_R1138_U389, P1_R1138_U387, P1_R1138_U388);
  not ginst1518 (P1_R1138_U39, P1_U3083);
  nand ginst1519 (P1_R1138_U390, P1_R1138_U352, P1_R1138_U45);
  nand ginst1520 (P1_R1138_U391, P1_R1138_U218, P1_R1138_U389);
  nand ginst1521 (P1_R1138_U392, P1_R1138_U33, P1_U3064);
  nand ginst1522 (P1_R1138_U393, P1_R1138_U34, P1_U3467);
  nand ginst1523 (P1_R1138_U394, P1_R1138_U392, P1_R1138_U393);
  nand ginst1524 (P1_R1138_U395, P1_R1138_U141, P1_R1138_U353);
  nand ginst1525 (P1_R1138_U396, P1_R1138_U227, P1_R1138_U394);
  nand ginst1526 (P1_R1138_U397, P1_R1138_U28, P1_U3068);
  nand ginst1527 (P1_R1138_U398, P1_R1138_U29, P1_U3464);
  nand ginst1528 (P1_R1138_U399, P1_R1138_U143, P1_U3055);
  and ginst1529 (P1_R1138_U4, P1_R1138_U175, P1_R1138_U176);
  not ginst1530 (P1_R1138_U40, P1_U3485);
  nand ginst1531 (P1_R1138_U400, P1_R1138_U142, P1_U4028);
  nand ginst1532 (P1_R1138_U401, P1_R1138_U143, P1_U3055);
  nand ginst1533 (P1_R1138_U402, P1_R1138_U142, P1_U4028);
  nand ginst1534 (P1_R1138_U403, P1_R1138_U401, P1_R1138_U402);
  nand ginst1535 (P1_R1138_U404, P1_R1138_U144, P1_R1138_U145);
  nand ginst1536 (P1_R1138_U405, P1_R1138_U302, P1_R1138_U403);
  nand ginst1537 (P1_R1138_U406, P1_R1138_U89, P1_U3054);
  nand ginst1538 (P1_R1138_U407, P1_R1138_U88, P1_U4017);
  nand ginst1539 (P1_R1138_U408, P1_R1138_U89, P1_U3054);
  nand ginst1540 (P1_R1138_U409, P1_R1138_U88, P1_U4017);
  nand ginst1541 (P1_R1138_U41, P1_R1138_U202, P1_R1138_U62);
  nand ginst1542 (P1_R1138_U410, P1_R1138_U408, P1_R1138_U409);
  nand ginst1543 (P1_R1138_U411, P1_R1138_U146, P1_R1138_U147);
  nand ginst1544 (P1_R1138_U412, P1_R1138_U300, P1_R1138_U410);
  nand ginst1545 (P1_R1138_U413, P1_R1138_U47, P1_U3053);
  nand ginst1546 (P1_R1138_U414, P1_R1138_U48, P1_U4018);
  nand ginst1547 (P1_R1138_U415, P1_R1138_U47, P1_U3053);
  nand ginst1548 (P1_R1138_U416, P1_R1138_U48, P1_U4018);
  nand ginst1549 (P1_R1138_U417, P1_R1138_U415, P1_R1138_U416);
  nand ginst1550 (P1_R1138_U418, P1_R1138_U148, P1_R1138_U149);
  nand ginst1551 (P1_R1138_U419, P1_R1138_U297, P1_R1138_U417);
  nand ginst1552 (P1_R1138_U42, P1_R1138_U118, P1_R1138_U190);
  nand ginst1553 (P1_R1138_U420, P1_R1138_U50, P1_U3057);
  nand ginst1554 (P1_R1138_U421, P1_R1138_U49, P1_U4019);
  nand ginst1555 (P1_R1138_U422, P1_R1138_U51, P1_U3058);
  nand ginst1556 (P1_R1138_U423, P1_R1138_U52, P1_U4020);
  nand ginst1557 (P1_R1138_U424, P1_R1138_U422, P1_R1138_U423);
  nand ginst1558 (P1_R1138_U425, P1_R1138_U354, P1_R1138_U90);
  nand ginst1559 (P1_R1138_U426, P1_R1138_U304, P1_R1138_U424);
  nand ginst1560 (P1_R1138_U427, P1_R1138_U53, P1_U3065);
  nand ginst1561 (P1_R1138_U428, P1_R1138_U54, P1_U4021);
  nand ginst1562 (P1_R1138_U429, P1_R1138_U427, P1_R1138_U428);
  nand ginst1563 (P1_R1138_U43, P1_R1138_U179, P1_R1138_U180);
  nand ginst1564 (P1_R1138_U430, P1_R1138_U151, P1_R1138_U355);
  nand ginst1565 (P1_R1138_U431, P1_R1138_U291, P1_R1138_U429);
  nand ginst1566 (P1_R1138_U432, P1_R1138_U85, P1_U3066);
  nand ginst1567 (P1_R1138_U433, P1_R1138_U86, P1_U4022);
  nand ginst1568 (P1_R1138_U434, P1_R1138_U85, P1_U3066);
  nand ginst1569 (P1_R1138_U435, P1_R1138_U86, P1_U4022);
  nand ginst1570 (P1_R1138_U436, P1_R1138_U434, P1_R1138_U435);
  nand ginst1571 (P1_R1138_U437, P1_R1138_U152, P1_R1138_U153);
  nand ginst1572 (P1_R1138_U438, P1_R1138_U287, P1_R1138_U436);
  nand ginst1573 (P1_R1138_U439, P1_R1138_U83, P1_U3061);
  nand ginst1574 (P1_R1138_U44, P1_U3078, P1_U3461);
  nand ginst1575 (P1_R1138_U440, P1_R1138_U84, P1_U4023);
  nand ginst1576 (P1_R1138_U441, P1_R1138_U83, P1_U3061);
  nand ginst1577 (P1_R1138_U442, P1_R1138_U84, P1_U4023);
  nand ginst1578 (P1_R1138_U443, P1_R1138_U441, P1_R1138_U442);
  nand ginst1579 (P1_R1138_U444, P1_R1138_U154, P1_R1138_U155);
  nand ginst1580 (P1_R1138_U445, P1_R1138_U283, P1_R1138_U443);
  nand ginst1581 (P1_R1138_U446, P1_R1138_U55, P1_U3075);
  nand ginst1582 (P1_R1138_U447, P1_R1138_U56, P1_U4024);
  nand ginst1583 (P1_R1138_U448, P1_R1138_U55, P1_U3075);
  nand ginst1584 (P1_R1138_U449, P1_R1138_U56, P1_U4024);
  nand ginst1585 (P1_R1138_U45, P1_R1138_U122, P1_R1138_U216);
  nand ginst1586 (P1_R1138_U450, P1_R1138_U448, P1_R1138_U449);
  nand ginst1587 (P1_R1138_U451, P1_R1138_U82, P1_U3076);
  nand ginst1588 (P1_R1138_U452, P1_R1138_U91, P1_U4025);
  nand ginst1589 (P1_R1138_U453, P1_R1138_U158, P1_R1138_U179);
  nand ginst1590 (P1_R1138_U454, P1_R1138_U32, P1_R1138_U325);
  nand ginst1591 (P1_R1138_U455, P1_R1138_U79, P1_U3081);
  nand ginst1592 (P1_R1138_U456, P1_R1138_U80, P1_U3514);
  nand ginst1593 (P1_R1138_U457, P1_R1138_U455, P1_R1138_U456);
  nand ginst1594 (P1_R1138_U458, P1_R1138_U356, P1_R1138_U92);
  nand ginst1595 (P1_R1138_U459, P1_R1138_U313, P1_R1138_U457);
  nand ginst1596 (P1_R1138_U46, P1_R1138_U212, P1_R1138_U213);
  nand ginst1597 (P1_R1138_U460, P1_R1138_U76, P1_U3082);
  nand ginst1598 (P1_R1138_U461, P1_R1138_U77, P1_U3512);
  nand ginst1599 (P1_R1138_U462, P1_R1138_U460, P1_R1138_U461);
  nand ginst1600 (P1_R1138_U463, P1_R1138_U159, P1_R1138_U357);
  nand ginst1601 (P1_R1138_U464, P1_R1138_U267, P1_R1138_U462);
  nand ginst1602 (P1_R1138_U465, P1_R1138_U61, P1_U3069);
  nand ginst1603 (P1_R1138_U466, P1_R1138_U59, P1_U3509);
  nand ginst1604 (P1_R1138_U467, P1_R1138_U57, P1_U3073);
  nand ginst1605 (P1_R1138_U468, P1_R1138_U58, P1_U3506);
  nand ginst1606 (P1_R1138_U469, P1_R1138_U467, P1_R1138_U468);
  not ginst1607 (P1_R1138_U47, P1_U4018);
  nand ginst1608 (P1_R1138_U470, P1_R1138_U358, P1_R1138_U93);
  nand ginst1609 (P1_R1138_U471, P1_R1138_U259, P1_R1138_U469);
  nand ginst1610 (P1_R1138_U472, P1_R1138_U74, P1_U3074);
  nand ginst1611 (P1_R1138_U473, P1_R1138_U75, P1_U3503);
  nand ginst1612 (P1_R1138_U474, P1_R1138_U74, P1_U3074);
  nand ginst1613 (P1_R1138_U475, P1_R1138_U75, P1_U3503);
  nand ginst1614 (P1_R1138_U476, P1_R1138_U474, P1_R1138_U475);
  nand ginst1615 (P1_R1138_U477, P1_R1138_U160, P1_R1138_U161);
  nand ginst1616 (P1_R1138_U478, P1_R1138_U255, P1_R1138_U476);
  nand ginst1617 (P1_R1138_U479, P1_R1138_U72, P1_U3079);
  not ginst1618 (P1_R1138_U48, P1_U3053);
  nand ginst1619 (P1_R1138_U480, P1_R1138_U73, P1_U3500);
  nand ginst1620 (P1_R1138_U481, P1_R1138_U72, P1_U3079);
  nand ginst1621 (P1_R1138_U482, P1_R1138_U73, P1_U3500);
  nand ginst1622 (P1_R1138_U483, P1_R1138_U481, P1_R1138_U482);
  nand ginst1623 (P1_R1138_U484, P1_R1138_U162, P1_R1138_U163);
  nand ginst1624 (P1_R1138_U485, P1_R1138_U251, P1_R1138_U483);
  nand ginst1625 (P1_R1138_U486, P1_R1138_U70, P1_U3080);
  nand ginst1626 (P1_R1138_U487, P1_R1138_U71, P1_U3497);
  nand ginst1627 (P1_R1138_U488, P1_R1138_U65, P1_U3072);
  nand ginst1628 (P1_R1138_U489, P1_R1138_U66, P1_U3494);
  not ginst1629 (P1_R1138_U49, P1_U3057);
  nand ginst1630 (P1_R1138_U490, P1_R1138_U488, P1_R1138_U489);
  nand ginst1631 (P1_R1138_U491, P1_R1138_U359, P1_R1138_U94);
  nand ginst1632 (P1_R1138_U492, P1_R1138_U335, P1_R1138_U490);
  nand ginst1633 (P1_R1138_U493, P1_R1138_U67, P1_U3063);
  nand ginst1634 (P1_R1138_U494, P1_R1138_U68, P1_U3491);
  nand ginst1635 (P1_R1138_U495, P1_R1138_U493, P1_R1138_U494);
  nand ginst1636 (P1_R1138_U496, P1_R1138_U164, P1_R1138_U360);
  nand ginst1637 (P1_R1138_U497, P1_R1138_U241, P1_R1138_U495);
  nand ginst1638 (P1_R1138_U498, P1_R1138_U63, P1_U3062);
  nand ginst1639 (P1_R1138_U499, P1_R1138_U64, P1_U3488);
  and ginst1640 (P1_R1138_U5, P1_R1138_U177, P1_R1138_U178);
  not ginst1641 (P1_R1138_U50, P1_U4019);
  nand ginst1642 (P1_R1138_U500, P1_R1138_U30, P1_U3077);
  nand ginst1643 (P1_R1138_U501, P1_R1138_U31, P1_U3456);
  not ginst1644 (P1_R1138_U51, P1_U4020);
  not ginst1645 (P1_R1138_U52, P1_U3058);
  not ginst1646 (P1_R1138_U53, P1_U4021);
  not ginst1647 (P1_R1138_U54, P1_U3065);
  not ginst1648 (P1_R1138_U55, P1_U4024);
  not ginst1649 (P1_R1138_U56, P1_U3075);
  not ginst1650 (P1_R1138_U57, P1_U3506);
  not ginst1651 (P1_R1138_U58, P1_U3073);
  not ginst1652 (P1_R1138_U59, P1_U3069);
  and ginst1653 (P1_R1138_U6, P1_R1138_U193, P1_R1138_U194);
  nand ginst1654 (P1_R1138_U60, P1_U3073, P1_U3506);
  not ginst1655 (P1_R1138_U61, P1_U3509);
  nand ginst1656 (P1_R1138_U62, P1_U3084, P1_U3482);
  not ginst1657 (P1_R1138_U63, P1_U3488);
  not ginst1658 (P1_R1138_U64, P1_U3062);
  not ginst1659 (P1_R1138_U65, P1_U3494);
  not ginst1660 (P1_R1138_U66, P1_U3072);
  not ginst1661 (P1_R1138_U67, P1_U3491);
  not ginst1662 (P1_R1138_U68, P1_U3063);
  nand ginst1663 (P1_R1138_U69, P1_U3063, P1_U3491);
  and ginst1664 (P1_R1138_U7, P1_R1138_U233, P1_R1138_U234);
  not ginst1665 (P1_R1138_U70, P1_U3497);
  not ginst1666 (P1_R1138_U71, P1_U3080);
  not ginst1667 (P1_R1138_U72, P1_U3500);
  not ginst1668 (P1_R1138_U73, P1_U3079);
  not ginst1669 (P1_R1138_U74, P1_U3503);
  not ginst1670 (P1_R1138_U75, P1_U3074);
  not ginst1671 (P1_R1138_U76, P1_U3512);
  not ginst1672 (P1_R1138_U77, P1_U3082);
  nand ginst1673 (P1_R1138_U78, P1_U3082, P1_U3512);
  not ginst1674 (P1_R1138_U79, P1_U3514);
  and ginst1675 (P1_R1138_U8, P1_R1138_U242, P1_R1138_U243);
  not ginst1676 (P1_R1138_U80, P1_U3081);
  nand ginst1677 (P1_R1138_U81, P1_U3081, P1_U3514);
  not ginst1678 (P1_R1138_U82, P1_U4025);
  not ginst1679 (P1_R1138_U83, P1_U4023);
  not ginst1680 (P1_R1138_U84, P1_U3061);
  not ginst1681 (P1_R1138_U85, P1_U4022);
  not ginst1682 (P1_R1138_U86, P1_U3066);
  nand ginst1683 (P1_R1138_U87, P1_U3057, P1_U4019);
  not ginst1684 (P1_R1138_U88, P1_U3054);
  not ginst1685 (P1_R1138_U89, P1_U4017);
  and ginst1686 (P1_R1138_U9, P1_R1138_U260, P1_R1138_U261);
  nand ginst1687 (P1_R1138_U90, P1_R1138_U173, P1_R1138_U303);
  not ginst1688 (P1_R1138_U91, P1_U3076);
  nand ginst1689 (P1_R1138_U92, P1_R1138_U312, P1_R1138_U78);
  nand ginst1690 (P1_R1138_U93, P1_R1138_U257, P1_R1138_U258);
  nand ginst1691 (P1_R1138_U94, P1_R1138_U334, P1_R1138_U69);
  nand ginst1692 (P1_R1138_U95, P1_R1138_U453, P1_R1138_U454);
  nand ginst1693 (P1_R1138_U96, P1_R1138_U500, P1_R1138_U501);
  nand ginst1694 (P1_R1138_U97, P1_R1138_U371, P1_R1138_U372);
  nand ginst1695 (P1_R1138_U98, P1_R1138_U376, P1_R1138_U377);
  nand ginst1696 (P1_R1138_U99, P1_R1138_U383, P1_R1138_U384);
  and ginst1697 (P1_R1150_U10, P1_R1150_U258, P1_R1150_U259);
  nand ginst1698 (P1_R1150_U100, P1_R1150_U442, P1_R1150_U443);
  nand ginst1699 (P1_R1150_U101, P1_R1150_U447, P1_R1150_U448);
  nand ginst1700 (P1_R1150_U102, P1_R1150_U463, P1_R1150_U464);
  nand ginst1701 (P1_R1150_U103, P1_R1150_U468, P1_R1150_U469);
  nand ginst1702 (P1_R1150_U104, P1_R1150_U351, P1_R1150_U352);
  nand ginst1703 (P1_R1150_U105, P1_R1150_U360, P1_R1150_U361);
  nand ginst1704 (P1_R1150_U106, P1_R1150_U367, P1_R1150_U368);
  nand ginst1705 (P1_R1150_U107, P1_R1150_U371, P1_R1150_U372);
  nand ginst1706 (P1_R1150_U108, P1_R1150_U380, P1_R1150_U381);
  nand ginst1707 (P1_R1150_U109, P1_R1150_U401, P1_R1150_U402);
  and ginst1708 (P1_R1150_U11, P1_R1150_U284, P1_R1150_U285);
  nand ginst1709 (P1_R1150_U110, P1_R1150_U418, P1_R1150_U419);
  nand ginst1710 (P1_R1150_U111, P1_R1150_U422, P1_R1150_U423);
  nand ginst1711 (P1_R1150_U112, P1_R1150_U454, P1_R1150_U455);
  nand ginst1712 (P1_R1150_U113, P1_R1150_U458, P1_R1150_U459);
  nand ginst1713 (P1_R1150_U114, P1_R1150_U475, P1_R1150_U476);
  and ginst1714 (P1_R1150_U115, P1_R1150_U183, P1_R1150_U195);
  and ginst1715 (P1_R1150_U116, P1_R1150_U198, P1_R1150_U199);
  and ginst1716 (P1_R1150_U117, P1_R1150_U185, P1_R1150_U211);
  and ginst1717 (P1_R1150_U118, P1_R1150_U214, P1_R1150_U215);
  and ginst1718 (P1_R1150_U119, P1_R1150_U353, P1_R1150_U354, P1_R1150_U40);
  and ginst1719 (P1_R1150_U12, P1_R1150_U382, P1_R1150_U383);
  and ginst1720 (P1_R1150_U120, P1_R1150_U185, P1_R1150_U357);
  and ginst1721 (P1_R1150_U121, P1_R1150_U230, P1_R1150_U7);
  and ginst1722 (P1_R1150_U122, P1_R1150_U184, P1_R1150_U364);
  and ginst1723 (P1_R1150_U123, P1_R1150_U29, P1_R1150_U373, P1_R1150_U374);
  and ginst1724 (P1_R1150_U124, P1_R1150_U183, P1_R1150_U377);
  and ginst1725 (P1_R1150_U125, P1_R1150_U217, P1_R1150_U8);
  and ginst1726 (P1_R1150_U126, P1_R1150_U180, P1_R1150_U262);
  and ginst1727 (P1_R1150_U127, P1_R1150_U181, P1_R1150_U288);
  and ginst1728 (P1_R1150_U128, P1_R1150_U304, P1_R1150_U305);
  and ginst1729 (P1_R1150_U129, P1_R1150_U307, P1_R1150_U386);
  nand ginst1730 (P1_R1150_U13, P1_R1150_U340, P1_R1150_U343);
  and ginst1731 (P1_R1150_U130, P1_R1150_U304, P1_R1150_U305, P1_R1150_U308);
  nand ginst1732 (P1_R1150_U131, P1_R1150_U389, P1_R1150_U390);
  and ginst1733 (P1_R1150_U132, P1_R1150_U394, P1_R1150_U395, P1_R1150_U85);
  and ginst1734 (P1_R1150_U133, P1_R1150_U182, P1_R1150_U398);
  nand ginst1735 (P1_R1150_U134, P1_R1150_U403, P1_R1150_U404);
  nand ginst1736 (P1_R1150_U135, P1_R1150_U408, P1_R1150_U409);
  and ginst1737 (P1_R1150_U136, P1_R1150_U181, P1_R1150_U415);
  nand ginst1738 (P1_R1150_U137, P1_R1150_U424, P1_R1150_U425);
  nand ginst1739 (P1_R1150_U138, P1_R1150_U429, P1_R1150_U430);
  nand ginst1740 (P1_R1150_U139, P1_R1150_U434, P1_R1150_U435);
  nand ginst1741 (P1_R1150_U14, P1_R1150_U329, P1_R1150_U332);
  nand ginst1742 (P1_R1150_U140, P1_R1150_U439, P1_R1150_U440);
  nand ginst1743 (P1_R1150_U141, P1_R1150_U444, P1_R1150_U445);
  and ginst1744 (P1_R1150_U142, P1_R1150_U180, P1_R1150_U451);
  nand ginst1745 (P1_R1150_U143, P1_R1150_U460, P1_R1150_U461);
  nand ginst1746 (P1_R1150_U144, P1_R1150_U465, P1_R1150_U466);
  and ginst1747 (P1_R1150_U145, P1_R1150_U342, P1_R1150_U9);
  and ginst1748 (P1_R1150_U146, P1_R1150_U179, P1_R1150_U472);
  and ginst1749 (P1_R1150_U147, P1_R1150_U349, P1_R1150_U350);
  nand ginst1750 (P1_R1150_U148, P1_R1150_U118, P1_R1150_U212);
  and ginst1751 (P1_R1150_U149, P1_R1150_U358, P1_R1150_U359);
  nand ginst1752 (P1_R1150_U15, P1_R1150_U318, P1_R1150_U321);
  and ginst1753 (P1_R1150_U150, P1_R1150_U365, P1_R1150_U366);
  and ginst1754 (P1_R1150_U151, P1_R1150_U369, P1_R1150_U370);
  nand ginst1755 (P1_R1150_U152, P1_R1150_U116, P1_R1150_U196);
  and ginst1756 (P1_R1150_U153, P1_R1150_U378, P1_R1150_U379);
  not ginst1757 (P1_R1150_U154, P1_U4028);
  not ginst1758 (P1_R1150_U155, P1_U3055);
  and ginst1759 (P1_R1150_U156, P1_R1150_U387, P1_R1150_U388);
  nand ginst1760 (P1_R1150_U157, P1_R1150_U128, P1_R1150_U302);
  and ginst1761 (P1_R1150_U158, P1_R1150_U399, P1_R1150_U400);
  nand ginst1762 (P1_R1150_U159, P1_R1150_U294, P1_R1150_U295);
  nand ginst1763 (P1_R1150_U16, P1_R1150_U310, P1_R1150_U312);
  nand ginst1764 (P1_R1150_U160, P1_R1150_U290, P1_R1150_U291);
  and ginst1765 (P1_R1150_U161, P1_R1150_U416, P1_R1150_U417);
  and ginst1766 (P1_R1150_U162, P1_R1150_U420, P1_R1150_U421);
  nand ginst1767 (P1_R1150_U163, P1_R1150_U280, P1_R1150_U281);
  nand ginst1768 (P1_R1150_U164, P1_R1150_U276, P1_R1150_U277);
  not ginst1769 (P1_R1150_U165, P1_U3461);
  nand ginst1770 (P1_R1150_U166, P1_R1150_U272, P1_R1150_U273);
  not ginst1771 (P1_R1150_U167, P1_U3512);
  nand ginst1772 (P1_R1150_U168, P1_R1150_U264, P1_R1150_U265);
  and ginst1773 (P1_R1150_U169, P1_R1150_U452, P1_R1150_U453);
  nand ginst1774 (P1_R1150_U17, P1_R1150_U156, P1_R1150_U175, P1_R1150_U348);
  and ginst1775 (P1_R1150_U170, P1_R1150_U456, P1_R1150_U457);
  nand ginst1776 (P1_R1150_U171, P1_R1150_U254, P1_R1150_U255);
  nand ginst1777 (P1_R1150_U172, P1_R1150_U250, P1_R1150_U251);
  nand ginst1778 (P1_R1150_U173, P1_R1150_U246, P1_R1150_U247);
  and ginst1779 (P1_R1150_U174, P1_R1150_U473, P1_R1150_U474);
  nand ginst1780 (P1_R1150_U175, P1_R1150_U129, P1_R1150_U157);
  not ginst1781 (P1_R1150_U176, P1_R1150_U85);
  not ginst1782 (P1_R1150_U177, P1_R1150_U29);
  not ginst1783 (P1_R1150_U178, P1_R1150_U40);
  nand ginst1784 (P1_R1150_U179, P1_R1150_U53, P1_U3488);
  nand ginst1785 (P1_R1150_U18, P1_R1150_U236, P1_R1150_U238);
  nand ginst1786 (P1_R1150_U180, P1_R1150_U62, P1_U3503);
  nand ginst1787 (P1_R1150_U181, P1_R1150_U76, P1_U4023);
  nand ginst1788 (P1_R1150_U182, P1_R1150_U84, P1_U4019);
  nand ginst1789 (P1_R1150_U183, P1_R1150_U28, P1_U3464);
  nand ginst1790 (P1_R1150_U184, P1_R1150_U35, P1_U3473);
  nand ginst1791 (P1_R1150_U185, P1_R1150_U39, P1_U3479);
  not ginst1792 (P1_R1150_U186, P1_R1150_U64);
  not ginst1793 (P1_R1150_U187, P1_R1150_U78);
  not ginst1794 (P1_R1150_U188, P1_R1150_U37);
  not ginst1795 (P1_R1150_U189, P1_R1150_U54);
  nand ginst1796 (P1_R1150_U19, P1_R1150_U228, P1_R1150_U231);
  not ginst1797 (P1_R1150_U190, P1_R1150_U25);
  nand ginst1798 (P1_R1150_U191, P1_R1150_U190, P1_R1150_U26);
  nand ginst1799 (P1_R1150_U192, P1_R1150_U165, P1_R1150_U191);
  nand ginst1800 (P1_R1150_U193, P1_R1150_U25, P1_U3078);
  not ginst1801 (P1_R1150_U194, P1_R1150_U46);
  nand ginst1802 (P1_R1150_U195, P1_R1150_U30, P1_U3467);
  nand ginst1803 (P1_R1150_U196, P1_R1150_U115, P1_R1150_U46);
  nand ginst1804 (P1_R1150_U197, P1_R1150_U29, P1_R1150_U30);
  nand ginst1805 (P1_R1150_U198, P1_R1150_U197, P1_R1150_U27);
  nand ginst1806 (P1_R1150_U199, P1_R1150_U177, P1_U3064);
  nand ginst1807 (P1_R1150_U20, P1_R1150_U220, P1_R1150_U222);
  not ginst1808 (P1_R1150_U200, P1_R1150_U152);
  nand ginst1809 (P1_R1150_U201, P1_R1150_U34, P1_U3476);
  nand ginst1810 (P1_R1150_U202, P1_R1150_U31, P1_U3071);
  nand ginst1811 (P1_R1150_U203, P1_R1150_U32, P1_U3067);
  nand ginst1812 (P1_R1150_U204, P1_R1150_U188, P1_R1150_U6);
  nand ginst1813 (P1_R1150_U205, P1_R1150_U204, P1_R1150_U7);
  nand ginst1814 (P1_R1150_U206, P1_R1150_U36, P1_U3470);
  nand ginst1815 (P1_R1150_U207, P1_R1150_U34, P1_U3476);
  nand ginst1816 (P1_R1150_U208, P1_R1150_U152, P1_R1150_U206, P1_R1150_U6);
  nand ginst1817 (P1_R1150_U209, P1_R1150_U205, P1_R1150_U207);
  nand ginst1818 (P1_R1150_U21, P1_R1150_U25, P1_R1150_U346);
  not ginst1819 (P1_R1150_U210, P1_R1150_U44);
  nand ginst1820 (P1_R1150_U211, P1_R1150_U41, P1_U3482);
  nand ginst1821 (P1_R1150_U212, P1_R1150_U117, P1_R1150_U44);
  nand ginst1822 (P1_R1150_U213, P1_R1150_U40, P1_R1150_U41);
  nand ginst1823 (P1_R1150_U214, P1_R1150_U213, P1_R1150_U38);
  nand ginst1824 (P1_R1150_U215, P1_R1150_U178, P1_U3084);
  not ginst1825 (P1_R1150_U216, P1_R1150_U148);
  nand ginst1826 (P1_R1150_U217, P1_R1150_U43, P1_U3485);
  nand ginst1827 (P1_R1150_U218, P1_R1150_U217, P1_R1150_U54);
  nand ginst1828 (P1_R1150_U219, P1_R1150_U210, P1_R1150_U40);
  not ginst1829 (P1_R1150_U22, P1_U3479);
  nand ginst1830 (P1_R1150_U220, P1_R1150_U120, P1_R1150_U219);
  nand ginst1831 (P1_R1150_U221, P1_R1150_U185, P1_R1150_U44);
  nand ginst1832 (P1_R1150_U222, P1_R1150_U119, P1_R1150_U221);
  nand ginst1833 (P1_R1150_U223, P1_R1150_U185, P1_R1150_U40);
  nand ginst1834 (P1_R1150_U224, P1_R1150_U152, P1_R1150_U206);
  not ginst1835 (P1_R1150_U225, P1_R1150_U45);
  nand ginst1836 (P1_R1150_U226, P1_R1150_U32, P1_U3067);
  nand ginst1837 (P1_R1150_U227, P1_R1150_U225, P1_R1150_U226);
  nand ginst1838 (P1_R1150_U228, P1_R1150_U122, P1_R1150_U227);
  nand ginst1839 (P1_R1150_U229, P1_R1150_U184, P1_R1150_U45);
  not ginst1840 (P1_R1150_U23, P1_U3464);
  nand ginst1841 (P1_R1150_U230, P1_R1150_U34, P1_U3476);
  nand ginst1842 (P1_R1150_U231, P1_R1150_U121, P1_R1150_U229);
  nand ginst1843 (P1_R1150_U232, P1_R1150_U32, P1_U3067);
  nand ginst1844 (P1_R1150_U233, P1_R1150_U184, P1_R1150_U232);
  nand ginst1845 (P1_R1150_U234, P1_R1150_U206, P1_R1150_U37);
  nand ginst1846 (P1_R1150_U235, P1_R1150_U194, P1_R1150_U29);
  nand ginst1847 (P1_R1150_U236, P1_R1150_U124, P1_R1150_U235);
  nand ginst1848 (P1_R1150_U237, P1_R1150_U183, P1_R1150_U46);
  nand ginst1849 (P1_R1150_U238, P1_R1150_U123, P1_R1150_U237);
  nand ginst1850 (P1_R1150_U239, P1_R1150_U183, P1_R1150_U29);
  not ginst1851 (P1_R1150_U24, P1_U3456);
  nand ginst1852 (P1_R1150_U240, P1_R1150_U52, P1_U3491);
  nand ginst1853 (P1_R1150_U241, P1_R1150_U50, P1_U3063);
  nand ginst1854 (P1_R1150_U242, P1_R1150_U51, P1_U3062);
  nand ginst1855 (P1_R1150_U243, P1_R1150_U189, P1_R1150_U8);
  nand ginst1856 (P1_R1150_U244, P1_R1150_U243, P1_R1150_U9);
  nand ginst1857 (P1_R1150_U245, P1_R1150_U52, P1_U3491);
  nand ginst1858 (P1_R1150_U246, P1_R1150_U125, P1_R1150_U148);
  nand ginst1859 (P1_R1150_U247, P1_R1150_U244, P1_R1150_U245);
  not ginst1860 (P1_R1150_U248, P1_R1150_U173);
  nand ginst1861 (P1_R1150_U249, P1_R1150_U56, P1_U3494);
  nand ginst1862 (P1_R1150_U25, P1_R1150_U93, P1_U3456);
  nand ginst1863 (P1_R1150_U250, P1_R1150_U173, P1_R1150_U249);
  nand ginst1864 (P1_R1150_U251, P1_R1150_U55, P1_U3072);
  not ginst1865 (P1_R1150_U252, P1_R1150_U172);
  nand ginst1866 (P1_R1150_U253, P1_R1150_U58, P1_U3497);
  nand ginst1867 (P1_R1150_U254, P1_R1150_U172, P1_R1150_U253);
  nand ginst1868 (P1_R1150_U255, P1_R1150_U57, P1_U3080);
  not ginst1869 (P1_R1150_U256, P1_R1150_U171);
  nand ginst1870 (P1_R1150_U257, P1_R1150_U61, P1_U3506);
  nand ginst1871 (P1_R1150_U258, P1_R1150_U59, P1_U3073);
  nand ginst1872 (P1_R1150_U259, P1_R1150_U49, P1_U3074);
  not ginst1873 (P1_R1150_U26, P1_U3078);
  nand ginst1874 (P1_R1150_U260, P1_R1150_U180, P1_R1150_U186);
  nand ginst1875 (P1_R1150_U261, P1_R1150_U10, P1_R1150_U260);
  nand ginst1876 (P1_R1150_U262, P1_R1150_U63, P1_U3500);
  nand ginst1877 (P1_R1150_U263, P1_R1150_U61, P1_U3506);
  nand ginst1878 (P1_R1150_U264, P1_R1150_U126, P1_R1150_U171, P1_R1150_U257);
  nand ginst1879 (P1_R1150_U265, P1_R1150_U261, P1_R1150_U263);
  not ginst1880 (P1_R1150_U266, P1_R1150_U168);
  nand ginst1881 (P1_R1150_U267, P1_R1150_U66, P1_U3509);
  nand ginst1882 (P1_R1150_U268, P1_R1150_U168, P1_R1150_U267);
  nand ginst1883 (P1_R1150_U269, P1_R1150_U65, P1_U3069);
  not ginst1884 (P1_R1150_U27, P1_U3467);
  not ginst1885 (P1_R1150_U270, P1_R1150_U67);
  nand ginst1886 (P1_R1150_U271, P1_R1150_U270, P1_R1150_U68);
  nand ginst1887 (P1_R1150_U272, P1_R1150_U167, P1_R1150_U271);
  nand ginst1888 (P1_R1150_U273, P1_R1150_U67, P1_U3082);
  not ginst1889 (P1_R1150_U274, P1_R1150_U166);
  nand ginst1890 (P1_R1150_U275, P1_R1150_U70, P1_U3514);
  nand ginst1891 (P1_R1150_U276, P1_R1150_U166, P1_R1150_U275);
  nand ginst1892 (P1_R1150_U277, P1_R1150_U69, P1_U3081);
  not ginst1893 (P1_R1150_U278, P1_R1150_U164);
  nand ginst1894 (P1_R1150_U279, P1_R1150_U72, P1_U4025);
  not ginst1895 (P1_R1150_U28, P1_U3068);
  nand ginst1896 (P1_R1150_U280, P1_R1150_U164, P1_R1150_U279);
  nand ginst1897 (P1_R1150_U281, P1_R1150_U71, P1_U3076);
  not ginst1898 (P1_R1150_U282, P1_R1150_U163);
  nand ginst1899 (P1_R1150_U283, P1_R1150_U75, P1_U4022);
  nand ginst1900 (P1_R1150_U284, P1_R1150_U73, P1_U3066);
  nand ginst1901 (P1_R1150_U285, P1_R1150_U48, P1_U3061);
  nand ginst1902 (P1_R1150_U286, P1_R1150_U181, P1_R1150_U187);
  nand ginst1903 (P1_R1150_U287, P1_R1150_U11, P1_R1150_U286);
  nand ginst1904 (P1_R1150_U288, P1_R1150_U77, P1_U4024);
  nand ginst1905 (P1_R1150_U289, P1_R1150_U75, P1_U4022);
  nand ginst1906 (P1_R1150_U29, P1_R1150_U23, P1_U3068);
  nand ginst1907 (P1_R1150_U290, P1_R1150_U127, P1_R1150_U163, P1_R1150_U283);
  nand ginst1908 (P1_R1150_U291, P1_R1150_U287, P1_R1150_U289);
  not ginst1909 (P1_R1150_U292, P1_R1150_U160);
  nand ginst1910 (P1_R1150_U293, P1_R1150_U80, P1_U4021);
  nand ginst1911 (P1_R1150_U294, P1_R1150_U160, P1_R1150_U293);
  nand ginst1912 (P1_R1150_U295, P1_R1150_U79, P1_U3065);
  not ginst1913 (P1_R1150_U296, P1_R1150_U159);
  nand ginst1914 (P1_R1150_U297, P1_R1150_U82, P1_U4020);
  nand ginst1915 (P1_R1150_U298, P1_R1150_U159, P1_R1150_U297);
  nand ginst1916 (P1_R1150_U299, P1_R1150_U81, P1_U3058);
  not ginst1917 (P1_R1150_U30, P1_U3064);
  not ginst1918 (P1_R1150_U300, P1_R1150_U89);
  nand ginst1919 (P1_R1150_U301, P1_R1150_U86, P1_U4018);
  nand ginst1920 (P1_R1150_U302, P1_R1150_U182, P1_R1150_U301, P1_R1150_U89);
  nand ginst1921 (P1_R1150_U303, P1_R1150_U85, P1_R1150_U86);
  nand ginst1922 (P1_R1150_U304, P1_R1150_U303, P1_R1150_U83);
  nand ginst1923 (P1_R1150_U305, P1_R1150_U176, P1_U3053);
  not ginst1924 (P1_R1150_U306, P1_R1150_U157);
  nand ginst1925 (P1_R1150_U307, P1_R1150_U88, P1_U4017);
  nand ginst1926 (P1_R1150_U308, P1_R1150_U87, P1_U3054);
  nand ginst1927 (P1_R1150_U309, P1_R1150_U300, P1_R1150_U85);
  not ginst1928 (P1_R1150_U31, P1_U3476);
  nand ginst1929 (P1_R1150_U310, P1_R1150_U133, P1_R1150_U309);
  nand ginst1930 (P1_R1150_U311, P1_R1150_U182, P1_R1150_U89);
  nand ginst1931 (P1_R1150_U312, P1_R1150_U132, P1_R1150_U311);
  nand ginst1932 (P1_R1150_U313, P1_R1150_U182, P1_R1150_U85);
  nand ginst1933 (P1_R1150_U314, P1_R1150_U163, P1_R1150_U288);
  not ginst1934 (P1_R1150_U315, P1_R1150_U90);
  nand ginst1935 (P1_R1150_U316, P1_R1150_U48, P1_U3061);
  nand ginst1936 (P1_R1150_U317, P1_R1150_U315, P1_R1150_U316);
  nand ginst1937 (P1_R1150_U318, P1_R1150_U136, P1_R1150_U317);
  nand ginst1938 (P1_R1150_U319, P1_R1150_U181, P1_R1150_U90);
  not ginst1939 (P1_R1150_U32, P1_U3473);
  nand ginst1940 (P1_R1150_U320, P1_R1150_U75, P1_U4022);
  nand ginst1941 (P1_R1150_U321, P1_R1150_U11, P1_R1150_U319, P1_R1150_U320);
  nand ginst1942 (P1_R1150_U322, P1_R1150_U48, P1_U3061);
  nand ginst1943 (P1_R1150_U323, P1_R1150_U181, P1_R1150_U322);
  nand ginst1944 (P1_R1150_U324, P1_R1150_U288, P1_R1150_U78);
  nand ginst1945 (P1_R1150_U325, P1_R1150_U171, P1_R1150_U262);
  not ginst1946 (P1_R1150_U326, P1_R1150_U91);
  nand ginst1947 (P1_R1150_U327, P1_R1150_U49, P1_U3074);
  nand ginst1948 (P1_R1150_U328, P1_R1150_U326, P1_R1150_U327);
  nand ginst1949 (P1_R1150_U329, P1_R1150_U142, P1_R1150_U328);
  not ginst1950 (P1_R1150_U33, P1_U3470);
  nand ginst1951 (P1_R1150_U330, P1_R1150_U180, P1_R1150_U91);
  nand ginst1952 (P1_R1150_U331, P1_R1150_U61, P1_U3506);
  nand ginst1953 (P1_R1150_U332, P1_R1150_U10, P1_R1150_U330, P1_R1150_U331);
  nand ginst1954 (P1_R1150_U333, P1_R1150_U49, P1_U3074);
  nand ginst1955 (P1_R1150_U334, P1_R1150_U180, P1_R1150_U333);
  nand ginst1956 (P1_R1150_U335, P1_R1150_U262, P1_R1150_U64);
  nand ginst1957 (P1_R1150_U336, P1_R1150_U148, P1_R1150_U217);
  not ginst1958 (P1_R1150_U337, P1_R1150_U92);
  nand ginst1959 (P1_R1150_U338, P1_R1150_U51, P1_U3062);
  nand ginst1960 (P1_R1150_U339, P1_R1150_U337, P1_R1150_U338);
  not ginst1961 (P1_R1150_U34, P1_U3071);
  nand ginst1962 (P1_R1150_U340, P1_R1150_U146, P1_R1150_U339);
  nand ginst1963 (P1_R1150_U341, P1_R1150_U179, P1_R1150_U92);
  nand ginst1964 (P1_R1150_U342, P1_R1150_U52, P1_U3491);
  nand ginst1965 (P1_R1150_U343, P1_R1150_U145, P1_R1150_U341);
  nand ginst1966 (P1_R1150_U344, P1_R1150_U51, P1_U3062);
  nand ginst1967 (P1_R1150_U345, P1_R1150_U179, P1_R1150_U344);
  nand ginst1968 (P1_R1150_U346, P1_R1150_U24, P1_U3077);
  nand ginst1969 (P1_R1150_U347, P1_R1150_U182, P1_R1150_U301, P1_R1150_U89);
  nand ginst1970 (P1_R1150_U348, P1_R1150_U12, P1_R1150_U130, P1_R1150_U347);
  nand ginst1971 (P1_R1150_U349, P1_R1150_U43, P1_U3485);
  not ginst1972 (P1_R1150_U35, P1_U3067);
  nand ginst1973 (P1_R1150_U350, P1_R1150_U42, P1_U3083);
  nand ginst1974 (P1_R1150_U351, P1_R1150_U148, P1_R1150_U218);
  nand ginst1975 (P1_R1150_U352, P1_R1150_U147, P1_R1150_U216);
  nand ginst1976 (P1_R1150_U353, P1_R1150_U41, P1_U3482);
  nand ginst1977 (P1_R1150_U354, P1_R1150_U38, P1_U3084);
  nand ginst1978 (P1_R1150_U355, P1_R1150_U41, P1_U3482);
  nand ginst1979 (P1_R1150_U356, P1_R1150_U38, P1_U3084);
  nand ginst1980 (P1_R1150_U357, P1_R1150_U355, P1_R1150_U356);
  nand ginst1981 (P1_R1150_U358, P1_R1150_U39, P1_U3479);
  nand ginst1982 (P1_R1150_U359, P1_R1150_U22, P1_U3070);
  not ginst1983 (P1_R1150_U36, P1_U3060);
  nand ginst1984 (P1_R1150_U360, P1_R1150_U223, P1_R1150_U44);
  nand ginst1985 (P1_R1150_U361, P1_R1150_U149, P1_R1150_U210);
  nand ginst1986 (P1_R1150_U362, P1_R1150_U34, P1_U3476);
  nand ginst1987 (P1_R1150_U363, P1_R1150_U31, P1_U3071);
  nand ginst1988 (P1_R1150_U364, P1_R1150_U362, P1_R1150_U363);
  nand ginst1989 (P1_R1150_U365, P1_R1150_U35, P1_U3473);
  nand ginst1990 (P1_R1150_U366, P1_R1150_U32, P1_U3067);
  nand ginst1991 (P1_R1150_U367, P1_R1150_U233, P1_R1150_U45);
  nand ginst1992 (P1_R1150_U368, P1_R1150_U150, P1_R1150_U225);
  nand ginst1993 (P1_R1150_U369, P1_R1150_U36, P1_U3470);
  nand ginst1994 (P1_R1150_U37, P1_R1150_U33, P1_U3060);
  nand ginst1995 (P1_R1150_U370, P1_R1150_U33, P1_U3060);
  nand ginst1996 (P1_R1150_U371, P1_R1150_U152, P1_R1150_U234);
  nand ginst1997 (P1_R1150_U372, P1_R1150_U151, P1_R1150_U200);
  nand ginst1998 (P1_R1150_U373, P1_R1150_U30, P1_U3467);
  nand ginst1999 (P1_R1150_U374, P1_R1150_U27, P1_U3064);
  nand ginst2000 (P1_R1150_U375, P1_R1150_U30, P1_U3467);
  nand ginst2001 (P1_R1150_U376, P1_R1150_U27, P1_U3064);
  nand ginst2002 (P1_R1150_U377, P1_R1150_U375, P1_R1150_U376);
  nand ginst2003 (P1_R1150_U378, P1_R1150_U28, P1_U3464);
  nand ginst2004 (P1_R1150_U379, P1_R1150_U23, P1_U3068);
  not ginst2005 (P1_R1150_U38, P1_U3482);
  nand ginst2006 (P1_R1150_U380, P1_R1150_U239, P1_R1150_U46);
  nand ginst2007 (P1_R1150_U381, P1_R1150_U153, P1_R1150_U194);
  nand ginst2008 (P1_R1150_U382, P1_R1150_U155, P1_U4028);
  nand ginst2009 (P1_R1150_U383, P1_R1150_U154, P1_U3055);
  nand ginst2010 (P1_R1150_U384, P1_R1150_U155, P1_U4028);
  nand ginst2011 (P1_R1150_U385, P1_R1150_U154, P1_U3055);
  nand ginst2012 (P1_R1150_U386, P1_R1150_U384, P1_R1150_U385);
  nand ginst2013 (P1_R1150_U387, P1_R1150_U386, P1_R1150_U87, P1_U3054);
  nand ginst2014 (P1_R1150_U388, P1_R1150_U12, P1_R1150_U88, P1_U4017);
  nand ginst2015 (P1_R1150_U389, P1_R1150_U88, P1_U4017);
  not ginst2016 (P1_R1150_U39, P1_U3070);
  nand ginst2017 (P1_R1150_U390, P1_R1150_U87, P1_U3054);
  not ginst2018 (P1_R1150_U391, P1_R1150_U131);
  nand ginst2019 (P1_R1150_U392, P1_R1150_U306, P1_R1150_U391);
  nand ginst2020 (P1_R1150_U393, P1_R1150_U131, P1_R1150_U157);
  nand ginst2021 (P1_R1150_U394, P1_R1150_U86, P1_U4018);
  nand ginst2022 (P1_R1150_U395, P1_R1150_U83, P1_U3053);
  nand ginst2023 (P1_R1150_U396, P1_R1150_U86, P1_U4018);
  nand ginst2024 (P1_R1150_U397, P1_R1150_U83, P1_U3053);
  nand ginst2025 (P1_R1150_U398, P1_R1150_U396, P1_R1150_U397);
  nand ginst2026 (P1_R1150_U399, P1_R1150_U84, P1_U4019);
  nand ginst2027 (P1_R1150_U40, P1_R1150_U22, P1_U3070);
  nand ginst2028 (P1_R1150_U400, P1_R1150_U47, P1_U3057);
  nand ginst2029 (P1_R1150_U401, P1_R1150_U313, P1_R1150_U89);
  nand ginst2030 (P1_R1150_U402, P1_R1150_U158, P1_R1150_U300);
  nand ginst2031 (P1_R1150_U403, P1_R1150_U82, P1_U4020);
  nand ginst2032 (P1_R1150_U404, P1_R1150_U81, P1_U3058);
  not ginst2033 (P1_R1150_U405, P1_R1150_U134);
  nand ginst2034 (P1_R1150_U406, P1_R1150_U296, P1_R1150_U405);
  nand ginst2035 (P1_R1150_U407, P1_R1150_U134, P1_R1150_U159);
  nand ginst2036 (P1_R1150_U408, P1_R1150_U80, P1_U4021);
  nand ginst2037 (P1_R1150_U409, P1_R1150_U79, P1_U3065);
  not ginst2038 (P1_R1150_U41, P1_U3084);
  not ginst2039 (P1_R1150_U410, P1_R1150_U135);
  nand ginst2040 (P1_R1150_U411, P1_R1150_U292, P1_R1150_U410);
  nand ginst2041 (P1_R1150_U412, P1_R1150_U135, P1_R1150_U160);
  nand ginst2042 (P1_R1150_U413, P1_R1150_U75, P1_U4022);
  nand ginst2043 (P1_R1150_U414, P1_R1150_U73, P1_U3066);
  nand ginst2044 (P1_R1150_U415, P1_R1150_U413, P1_R1150_U414);
  nand ginst2045 (P1_R1150_U416, P1_R1150_U76, P1_U4023);
  nand ginst2046 (P1_R1150_U417, P1_R1150_U48, P1_U3061);
  nand ginst2047 (P1_R1150_U418, P1_R1150_U323, P1_R1150_U90);
  nand ginst2048 (P1_R1150_U419, P1_R1150_U161, P1_R1150_U315);
  not ginst2049 (P1_R1150_U42, P1_U3485);
  nand ginst2050 (P1_R1150_U420, P1_R1150_U77, P1_U4024);
  nand ginst2051 (P1_R1150_U421, P1_R1150_U74, P1_U3075);
  nand ginst2052 (P1_R1150_U422, P1_R1150_U163, P1_R1150_U324);
  nand ginst2053 (P1_R1150_U423, P1_R1150_U162, P1_R1150_U282);
  nand ginst2054 (P1_R1150_U424, P1_R1150_U72, P1_U4025);
  nand ginst2055 (P1_R1150_U425, P1_R1150_U71, P1_U3076);
  not ginst2056 (P1_R1150_U426, P1_R1150_U137);
  nand ginst2057 (P1_R1150_U427, P1_R1150_U278, P1_R1150_U426);
  nand ginst2058 (P1_R1150_U428, P1_R1150_U137, P1_R1150_U164);
  nand ginst2059 (P1_R1150_U429, P1_R1150_U26, P1_U3461);
  not ginst2060 (P1_R1150_U43, P1_U3083);
  nand ginst2061 (P1_R1150_U430, P1_R1150_U165, P1_U3078);
  not ginst2062 (P1_R1150_U431, P1_R1150_U138);
  nand ginst2063 (P1_R1150_U432, P1_R1150_U190, P1_R1150_U431);
  nand ginst2064 (P1_R1150_U433, P1_R1150_U138, P1_R1150_U25);
  nand ginst2065 (P1_R1150_U434, P1_R1150_U70, P1_U3514);
  nand ginst2066 (P1_R1150_U435, P1_R1150_U69, P1_U3081);
  not ginst2067 (P1_R1150_U436, P1_R1150_U139);
  nand ginst2068 (P1_R1150_U437, P1_R1150_U274, P1_R1150_U436);
  nand ginst2069 (P1_R1150_U438, P1_R1150_U139, P1_R1150_U166);
  nand ginst2070 (P1_R1150_U439, P1_R1150_U68, P1_U3512);
  nand ginst2071 (P1_R1150_U44, P1_R1150_U208, P1_R1150_U209);
  nand ginst2072 (P1_R1150_U440, P1_R1150_U167, P1_U3082);
  not ginst2073 (P1_R1150_U441, P1_R1150_U140);
  nand ginst2074 (P1_R1150_U442, P1_R1150_U270, P1_R1150_U441);
  nand ginst2075 (P1_R1150_U443, P1_R1150_U140, P1_R1150_U67);
  nand ginst2076 (P1_R1150_U444, P1_R1150_U66, P1_U3509);
  nand ginst2077 (P1_R1150_U445, P1_R1150_U65, P1_U3069);
  not ginst2078 (P1_R1150_U446, P1_R1150_U141);
  nand ginst2079 (P1_R1150_U447, P1_R1150_U266, P1_R1150_U446);
  nand ginst2080 (P1_R1150_U448, P1_R1150_U141, P1_R1150_U168);
  nand ginst2081 (P1_R1150_U449, P1_R1150_U61, P1_U3506);
  nand ginst2082 (P1_R1150_U45, P1_R1150_U224, P1_R1150_U37);
  nand ginst2083 (P1_R1150_U450, P1_R1150_U59, P1_U3073);
  nand ginst2084 (P1_R1150_U451, P1_R1150_U449, P1_R1150_U450);
  nand ginst2085 (P1_R1150_U452, P1_R1150_U62, P1_U3503);
  nand ginst2086 (P1_R1150_U453, P1_R1150_U49, P1_U3074);
  nand ginst2087 (P1_R1150_U454, P1_R1150_U334, P1_R1150_U91);
  nand ginst2088 (P1_R1150_U455, P1_R1150_U169, P1_R1150_U326);
  nand ginst2089 (P1_R1150_U456, P1_R1150_U63, P1_U3500);
  nand ginst2090 (P1_R1150_U457, P1_R1150_U60, P1_U3079);
  nand ginst2091 (P1_R1150_U458, P1_R1150_U171, P1_R1150_U335);
  nand ginst2092 (P1_R1150_U459, P1_R1150_U170, P1_R1150_U256);
  nand ginst2093 (P1_R1150_U46, P1_R1150_U192, P1_R1150_U193);
  nand ginst2094 (P1_R1150_U460, P1_R1150_U58, P1_U3497);
  nand ginst2095 (P1_R1150_U461, P1_R1150_U57, P1_U3080);
  not ginst2096 (P1_R1150_U462, P1_R1150_U143);
  nand ginst2097 (P1_R1150_U463, P1_R1150_U252, P1_R1150_U462);
  nand ginst2098 (P1_R1150_U464, P1_R1150_U143, P1_R1150_U172);
  nand ginst2099 (P1_R1150_U465, P1_R1150_U56, P1_U3494);
  nand ginst2100 (P1_R1150_U466, P1_R1150_U55, P1_U3072);
  not ginst2101 (P1_R1150_U467, P1_R1150_U144);
  nand ginst2102 (P1_R1150_U468, P1_R1150_U248, P1_R1150_U467);
  nand ginst2103 (P1_R1150_U469, P1_R1150_U144, P1_R1150_U173);
  not ginst2104 (P1_R1150_U47, P1_U4019);
  nand ginst2105 (P1_R1150_U470, P1_R1150_U52, P1_U3491);
  nand ginst2106 (P1_R1150_U471, P1_R1150_U50, P1_U3063);
  nand ginst2107 (P1_R1150_U472, P1_R1150_U470, P1_R1150_U471);
  nand ginst2108 (P1_R1150_U473, P1_R1150_U53, P1_U3488);
  nand ginst2109 (P1_R1150_U474, P1_R1150_U51, P1_U3062);
  nand ginst2110 (P1_R1150_U475, P1_R1150_U345, P1_R1150_U92);
  nand ginst2111 (P1_R1150_U476, P1_R1150_U174, P1_R1150_U337);
  not ginst2112 (P1_R1150_U48, P1_U4023);
  not ginst2113 (P1_R1150_U49, P1_U3503);
  not ginst2114 (P1_R1150_U50, P1_U3491);
  not ginst2115 (P1_R1150_U51, P1_U3488);
  not ginst2116 (P1_R1150_U52, P1_U3063);
  not ginst2117 (P1_R1150_U53, P1_U3062);
  nand ginst2118 (P1_R1150_U54, P1_R1150_U42, P1_U3083);
  not ginst2119 (P1_R1150_U55, P1_U3494);
  not ginst2120 (P1_R1150_U56, P1_U3072);
  not ginst2121 (P1_R1150_U57, P1_U3497);
  not ginst2122 (P1_R1150_U58, P1_U3080);
  not ginst2123 (P1_R1150_U59, P1_U3506);
  and ginst2124 (P1_R1150_U6, P1_R1150_U184, P1_R1150_U201);
  not ginst2125 (P1_R1150_U60, P1_U3500);
  not ginst2126 (P1_R1150_U61, P1_U3073);
  not ginst2127 (P1_R1150_U62, P1_U3074);
  not ginst2128 (P1_R1150_U63, P1_U3079);
  nand ginst2129 (P1_R1150_U64, P1_R1150_U60, P1_U3079);
  not ginst2130 (P1_R1150_U65, P1_U3509);
  not ginst2131 (P1_R1150_U66, P1_U3069);
  nand ginst2132 (P1_R1150_U67, P1_R1150_U268, P1_R1150_U269);
  not ginst2133 (P1_R1150_U68, P1_U3082);
  not ginst2134 (P1_R1150_U69, P1_U3514);
  and ginst2135 (P1_R1150_U7, P1_R1150_U202, P1_R1150_U203);
  not ginst2136 (P1_R1150_U70, P1_U3081);
  not ginst2137 (P1_R1150_U71, P1_U4025);
  not ginst2138 (P1_R1150_U72, P1_U3076);
  not ginst2139 (P1_R1150_U73, P1_U4022);
  not ginst2140 (P1_R1150_U74, P1_U4024);
  not ginst2141 (P1_R1150_U75, P1_U3066);
  not ginst2142 (P1_R1150_U76, P1_U3061);
  not ginst2143 (P1_R1150_U77, P1_U3075);
  nand ginst2144 (P1_R1150_U78, P1_R1150_U74, P1_U3075);
  not ginst2145 (P1_R1150_U79, P1_U4021);
  and ginst2146 (P1_R1150_U8, P1_R1150_U179, P1_R1150_U240);
  not ginst2147 (P1_R1150_U80, P1_U3065);
  not ginst2148 (P1_R1150_U81, P1_U4020);
  not ginst2149 (P1_R1150_U82, P1_U3058);
  not ginst2150 (P1_R1150_U83, P1_U4018);
  not ginst2151 (P1_R1150_U84, P1_U3057);
  nand ginst2152 (P1_R1150_U85, P1_R1150_U47, P1_U3057);
  not ginst2153 (P1_R1150_U86, P1_U3053);
  not ginst2154 (P1_R1150_U87, P1_U4017);
  not ginst2155 (P1_R1150_U88, P1_U3054);
  nand ginst2156 (P1_R1150_U89, P1_R1150_U298, P1_R1150_U299);
  and ginst2157 (P1_R1150_U9, P1_R1150_U241, P1_R1150_U242);
  nand ginst2158 (P1_R1150_U90, P1_R1150_U314, P1_R1150_U78);
  nand ginst2159 (P1_R1150_U91, P1_R1150_U325, P1_R1150_U64);
  nand ginst2160 (P1_R1150_U92, P1_R1150_U336, P1_R1150_U54);
  not ginst2161 (P1_R1150_U93, P1_U3077);
  nand ginst2162 (P1_R1150_U94, P1_R1150_U392, P1_R1150_U393);
  nand ginst2163 (P1_R1150_U95, P1_R1150_U406, P1_R1150_U407);
  nand ginst2164 (P1_R1150_U96, P1_R1150_U411, P1_R1150_U412);
  nand ginst2165 (P1_R1150_U97, P1_R1150_U427, P1_R1150_U428);
  nand ginst2166 (P1_R1150_U98, P1_R1150_U432, P1_R1150_U433);
  nand ginst2167 (P1_R1150_U99, P1_R1150_U437, P1_R1150_U438);
  and ginst2168 (P1_R1162_U10, P1_R1162_U215, P1_R1162_U218);
  not ginst2169 (P1_R1162_U100, P1_R1162_U40);
  not ginst2170 (P1_R1162_U101, P1_R1162_U41);
  nand ginst2171 (P1_R1162_U102, P1_R1162_U40, P1_R1162_U41);
  nand ginst2172 (P1_R1162_U103, P1_REG1_REG_2__SCAN_IN, P1_R1162_U96, P1_U3463);
  nand ginst2173 (P1_R1162_U104, P1_R1162_U102, P1_R1162_U5);
  nand ginst2174 (P1_R1162_U105, P1_REG1_REG_3__SCAN_IN, P1_U3466);
  nand ginst2175 (P1_R1162_U106, P1_R1162_U103, P1_R1162_U104, P1_R1162_U105);
  nand ginst2176 (P1_R1162_U107, P1_R1162_U32, P1_R1162_U33);
  nand ginst2177 (P1_R1162_U108, P1_R1162_U107, P1_U3472);
  nand ginst2178 (P1_R1162_U109, P1_R1162_U106, P1_R1162_U4);
  and ginst2179 (P1_R1162_U11, P1_R1162_U208, P1_R1162_U211);
  nand ginst2180 (P1_R1162_U110, P1_REG1_REG_5__SCAN_IN, P1_R1162_U89);
  not ginst2181 (P1_R1162_U111, P1_R1162_U39);
  or ginst2182 (P1_R1162_U112, P1_REG1_REG_7__SCAN_IN, P1_U3478);
  or ginst2183 (P1_R1162_U113, P1_REG1_REG_6__SCAN_IN, P1_U3475);
  not ginst2184 (P1_R1162_U114, P1_R1162_U20);
  nand ginst2185 (P1_R1162_U115, P1_R1162_U20, P1_R1162_U21);
  nand ginst2186 (P1_R1162_U116, P1_R1162_U115, P1_U3478);
  nand ginst2187 (P1_R1162_U117, P1_REG1_REG_7__SCAN_IN, P1_R1162_U114);
  nand ginst2188 (P1_R1162_U118, P1_R1162_U39, P1_R1162_U6);
  not ginst2189 (P1_R1162_U119, P1_R1162_U81);
  and ginst2190 (P1_R1162_U12, P1_R1162_U199, P1_R1162_U202);
  or ginst2191 (P1_R1162_U120, P1_REG1_REG_8__SCAN_IN, P1_U3481);
  nand ginst2192 (P1_R1162_U121, P1_R1162_U120, P1_R1162_U81);
  not ginst2193 (P1_R1162_U122, P1_R1162_U38);
  or ginst2194 (P1_R1162_U123, P1_REG1_REG_9__SCAN_IN, P1_U3484);
  or ginst2195 (P1_R1162_U124, P1_REG1_REG_6__SCAN_IN, P1_U3475);
  nand ginst2196 (P1_R1162_U125, P1_R1162_U124, P1_R1162_U39);
  nand ginst2197 (P1_R1162_U126, P1_R1162_U125, P1_R1162_U20, P1_R1162_U237, P1_R1162_U238);
  nand ginst2198 (P1_R1162_U127, P1_R1162_U111, P1_R1162_U20);
  nand ginst2199 (P1_R1162_U128, P1_REG1_REG_7__SCAN_IN, P1_U3478);
  nand ginst2200 (P1_R1162_U129, P1_R1162_U127, P1_R1162_U128, P1_R1162_U6);
  and ginst2201 (P1_R1162_U13, P1_R1162_U192, P1_R1162_U196);
  or ginst2202 (P1_R1162_U130, P1_REG1_REG_6__SCAN_IN, P1_U3475);
  nand ginst2203 (P1_R1162_U131, P1_R1162_U101, P1_R1162_U97);
  nand ginst2204 (P1_R1162_U132, P1_REG1_REG_2__SCAN_IN, P1_U3463);
  not ginst2205 (P1_R1162_U133, P1_R1162_U43);
  nand ginst2206 (P1_R1162_U134, P1_R1162_U100, P1_R1162_U5);
  nand ginst2207 (P1_R1162_U135, P1_R1162_U43, P1_R1162_U96);
  nand ginst2208 (P1_R1162_U136, P1_REG1_REG_3__SCAN_IN, P1_U3466);
  not ginst2209 (P1_R1162_U137, P1_R1162_U42);
  or ginst2210 (P1_R1162_U138, P1_REG1_REG_4__SCAN_IN, P1_U3469);
  nand ginst2211 (P1_R1162_U139, P1_R1162_U138, P1_R1162_U42);
  and ginst2212 (P1_R1162_U14, P1_R1162_U148, P1_R1162_U151);
  nand ginst2213 (P1_R1162_U140, P1_R1162_U139, P1_R1162_U244, P1_R1162_U245, P1_R1162_U32);
  nand ginst2214 (P1_R1162_U141, P1_R1162_U137, P1_R1162_U32);
  nand ginst2215 (P1_R1162_U142, P1_REG1_REG_5__SCAN_IN, P1_U3472);
  nand ginst2216 (P1_R1162_U143, P1_R1162_U141, P1_R1162_U142, P1_R1162_U4);
  or ginst2217 (P1_R1162_U144, P1_REG1_REG_4__SCAN_IN, P1_U3469);
  nand ginst2218 (P1_R1162_U145, P1_R1162_U100, P1_R1162_U97);
  not ginst2219 (P1_R1162_U146, P1_R1162_U82);
  nand ginst2220 (P1_R1162_U147, P1_REG1_REG_3__SCAN_IN, P1_U3466);
  nand ginst2221 (P1_R1162_U148, P1_R1162_U256, P1_R1162_U257, P1_R1162_U40, P1_R1162_U41);
  nand ginst2222 (P1_R1162_U149, P1_R1162_U40, P1_R1162_U41);
  and ginst2223 (P1_R1162_U15, P1_R1162_U140, P1_R1162_U143);
  nand ginst2224 (P1_R1162_U150, P1_REG1_REG_2__SCAN_IN, P1_U3463);
  nand ginst2225 (P1_R1162_U151, P1_R1162_U149, P1_R1162_U150, P1_R1162_U97);
  or ginst2226 (P1_R1162_U152, P1_REG1_REG_1__SCAN_IN, P1_U3460);
  not ginst2227 (P1_R1162_U153, P1_R1162_U83);
  or ginst2228 (P1_R1162_U154, P1_REG1_REG_9__SCAN_IN, P1_U3484);
  or ginst2229 (P1_R1162_U155, P1_REG1_REG_10__SCAN_IN, P1_U3487);
  nand ginst2230 (P1_R1162_U156, P1_R1162_U7, P1_R1162_U93);
  nand ginst2231 (P1_R1162_U157, P1_REG1_REG_10__SCAN_IN, P1_U3487);
  nand ginst2232 (P1_R1162_U158, P1_R1162_U156, P1_R1162_U157, P1_R1162_U90);
  or ginst2233 (P1_R1162_U159, P1_REG1_REG_10__SCAN_IN, P1_U3487);
  and ginst2234 (P1_R1162_U16, P1_R1162_U126, P1_R1162_U129);
  nand ginst2235 (P1_R1162_U160, P1_R1162_U120, P1_R1162_U7, P1_R1162_U81);
  nand ginst2236 (P1_R1162_U161, P1_R1162_U158, P1_R1162_U159);
  not ginst2237 (P1_R1162_U162, P1_R1162_U88);
  or ginst2238 (P1_R1162_U163, P1_REG1_REG_13__SCAN_IN, P1_U3496);
  or ginst2239 (P1_R1162_U164, P1_REG1_REG_12__SCAN_IN, P1_U3493);
  nand ginst2240 (P1_R1162_U165, P1_R1162_U8, P1_R1162_U92);
  nand ginst2241 (P1_R1162_U166, P1_REG1_REG_13__SCAN_IN, P1_U3496);
  nand ginst2242 (P1_R1162_U167, P1_R1162_U165, P1_R1162_U166, P1_R1162_U91);
  or ginst2243 (P1_R1162_U168, P1_REG1_REG_11__SCAN_IN, P1_U3490);
  or ginst2244 (P1_R1162_U169, P1_REG1_REG_13__SCAN_IN, P1_U3496);
  not ginst2245 (P1_R1162_U17, P1_REG1_REG_6__SCAN_IN);
  nand ginst2246 (P1_R1162_U170, P1_R1162_U168, P1_R1162_U8, P1_R1162_U88);
  nand ginst2247 (P1_R1162_U171, P1_R1162_U167, P1_R1162_U169);
  not ginst2248 (P1_R1162_U172, P1_R1162_U87);
  or ginst2249 (P1_R1162_U173, P1_REG1_REG_14__SCAN_IN, P1_U3499);
  nand ginst2250 (P1_R1162_U174, P1_R1162_U173, P1_R1162_U87);
  nand ginst2251 (P1_R1162_U175, P1_REG1_REG_14__SCAN_IN, P1_U3499);
  not ginst2252 (P1_R1162_U176, P1_R1162_U86);
  or ginst2253 (P1_R1162_U177, P1_REG1_REG_15__SCAN_IN, P1_U3502);
  nand ginst2254 (P1_R1162_U178, P1_R1162_U177, P1_R1162_U86);
  nand ginst2255 (P1_R1162_U179, P1_REG1_REG_15__SCAN_IN, P1_U3502);
  not ginst2256 (P1_R1162_U18, P1_U3475);
  not ginst2257 (P1_R1162_U180, P1_R1162_U66);
  or ginst2258 (P1_R1162_U181, P1_REG1_REG_17__SCAN_IN, P1_U3508);
  or ginst2259 (P1_R1162_U182, P1_REG1_REG_16__SCAN_IN, P1_U3505);
  not ginst2260 (P1_R1162_U183, P1_R1162_U47);
  nand ginst2261 (P1_R1162_U184, P1_R1162_U47, P1_R1162_U48);
  nand ginst2262 (P1_R1162_U185, P1_R1162_U184, P1_U3508);
  nand ginst2263 (P1_R1162_U186, P1_REG1_REG_17__SCAN_IN, P1_R1162_U183);
  nand ginst2264 (P1_R1162_U187, P1_R1162_U66, P1_R1162_U9);
  not ginst2265 (P1_R1162_U188, P1_R1162_U65);
  or ginst2266 (P1_R1162_U189, P1_REG1_REG_18__SCAN_IN, P1_U3511);
  not ginst2267 (P1_R1162_U19, P1_U3478);
  nand ginst2268 (P1_R1162_U190, P1_R1162_U189, P1_R1162_U65);
  nand ginst2269 (P1_R1162_U191, P1_REG1_REG_18__SCAN_IN, P1_U3511);
  nand ginst2270 (P1_R1162_U192, P1_R1162_U190, P1_R1162_U191, P1_R1162_U260, P1_R1162_U261);
  nand ginst2271 (P1_R1162_U193, P1_REG1_REG_18__SCAN_IN, P1_U3511);
  nand ginst2272 (P1_R1162_U194, P1_R1162_U188, P1_R1162_U193);
  or ginst2273 (P1_R1162_U195, P1_REG1_REG_18__SCAN_IN, P1_U3511);
  nand ginst2274 (P1_R1162_U196, P1_R1162_U194, P1_R1162_U195, P1_R1162_U264);
  or ginst2275 (P1_R1162_U197, P1_REG1_REG_16__SCAN_IN, P1_U3505);
  nand ginst2276 (P1_R1162_U198, P1_R1162_U197, P1_R1162_U66);
  nand ginst2277 (P1_R1162_U199, P1_R1162_U198, P1_R1162_U272, P1_R1162_U273, P1_R1162_U47);
  nand ginst2278 (P1_R1162_U20, P1_REG1_REG_6__SCAN_IN, P1_U3475);
  nand ginst2279 (P1_R1162_U200, P1_R1162_U180, P1_R1162_U47);
  nand ginst2280 (P1_R1162_U201, P1_REG1_REG_17__SCAN_IN, P1_U3508);
  nand ginst2281 (P1_R1162_U202, P1_R1162_U200, P1_R1162_U201, P1_R1162_U9);
  or ginst2282 (P1_R1162_U203, P1_REG1_REG_16__SCAN_IN, P1_U3505);
  nand ginst2283 (P1_R1162_U204, P1_R1162_U168, P1_R1162_U88);
  not ginst2284 (P1_R1162_U205, P1_R1162_U67);
  or ginst2285 (P1_R1162_U206, P1_REG1_REG_12__SCAN_IN, P1_U3493);
  nand ginst2286 (P1_R1162_U207, P1_R1162_U206, P1_R1162_U67);
  nand ginst2287 (P1_R1162_U208, P1_R1162_U207, P1_R1162_U293, P1_R1162_U294, P1_R1162_U91);
  nand ginst2288 (P1_R1162_U209, P1_R1162_U205, P1_R1162_U91);
  not ginst2289 (P1_R1162_U21, P1_REG1_REG_7__SCAN_IN);
  nand ginst2290 (P1_R1162_U210, P1_REG1_REG_13__SCAN_IN, P1_U3496);
  nand ginst2291 (P1_R1162_U211, P1_R1162_U209, P1_R1162_U210, P1_R1162_U8);
  or ginst2292 (P1_R1162_U212, P1_REG1_REG_12__SCAN_IN, P1_U3493);
  or ginst2293 (P1_R1162_U213, P1_REG1_REG_9__SCAN_IN, P1_U3484);
  nand ginst2294 (P1_R1162_U214, P1_R1162_U213, P1_R1162_U38);
  nand ginst2295 (P1_R1162_U215, P1_R1162_U214, P1_R1162_U305, P1_R1162_U306, P1_R1162_U90);
  nand ginst2296 (P1_R1162_U216, P1_R1162_U122, P1_R1162_U90);
  nand ginst2297 (P1_R1162_U217, P1_REG1_REG_10__SCAN_IN, P1_U3487);
  nand ginst2298 (P1_R1162_U218, P1_R1162_U216, P1_R1162_U217, P1_R1162_U7);
  nand ginst2299 (P1_R1162_U219, P1_R1162_U123, P1_R1162_U90);
  not ginst2300 (P1_R1162_U22, P1_REG1_REG_4__SCAN_IN);
  nand ginst2301 (P1_R1162_U220, P1_R1162_U120, P1_R1162_U49);
  nand ginst2302 (P1_R1162_U221, P1_R1162_U130, P1_R1162_U20);
  nand ginst2303 (P1_R1162_U222, P1_R1162_U144, P1_R1162_U32);
  nand ginst2304 (P1_R1162_U223, P1_R1162_U147, P1_R1162_U96);
  nand ginst2305 (P1_R1162_U224, P1_R1162_U203, P1_R1162_U47);
  nand ginst2306 (P1_R1162_U225, P1_R1162_U212, P1_R1162_U91);
  nand ginst2307 (P1_R1162_U226, P1_R1162_U168, P1_R1162_U56);
  nand ginst2308 (P1_R1162_U227, P1_R1162_U37, P1_U3484);
  nand ginst2309 (P1_R1162_U228, P1_REG1_REG_9__SCAN_IN, P1_R1162_U36);
  nand ginst2310 (P1_R1162_U229, P1_R1162_U227, P1_R1162_U228);
  not ginst2311 (P1_R1162_U23, P1_U3469);
  nand ginst2312 (P1_R1162_U230, P1_R1162_U219, P1_R1162_U38);
  nand ginst2313 (P1_R1162_U231, P1_R1162_U122, P1_R1162_U229);
  nand ginst2314 (P1_R1162_U232, P1_R1162_U34, P1_U3481);
  nand ginst2315 (P1_R1162_U233, P1_REG1_REG_8__SCAN_IN, P1_R1162_U35);
  nand ginst2316 (P1_R1162_U234, P1_R1162_U232, P1_R1162_U233);
  nand ginst2317 (P1_R1162_U235, P1_R1162_U220, P1_R1162_U81);
  nand ginst2318 (P1_R1162_U236, P1_R1162_U119, P1_R1162_U234);
  nand ginst2319 (P1_R1162_U237, P1_R1162_U21, P1_U3478);
  nand ginst2320 (P1_R1162_U238, P1_REG1_REG_7__SCAN_IN, P1_R1162_U19);
  nand ginst2321 (P1_R1162_U239, P1_R1162_U17, P1_U3475);
  not ginst2322 (P1_R1162_U24, P1_U3472);
  nand ginst2323 (P1_R1162_U240, P1_REG1_REG_6__SCAN_IN, P1_R1162_U18);
  nand ginst2324 (P1_R1162_U241, P1_R1162_U239, P1_R1162_U240);
  nand ginst2325 (P1_R1162_U242, P1_R1162_U221, P1_R1162_U39);
  nand ginst2326 (P1_R1162_U243, P1_R1162_U111, P1_R1162_U241);
  nand ginst2327 (P1_R1162_U244, P1_R1162_U33, P1_U3472);
  nand ginst2328 (P1_R1162_U245, P1_REG1_REG_5__SCAN_IN, P1_R1162_U24);
  nand ginst2329 (P1_R1162_U246, P1_R1162_U22, P1_U3469);
  nand ginst2330 (P1_R1162_U247, P1_REG1_REG_4__SCAN_IN, P1_R1162_U23);
  nand ginst2331 (P1_R1162_U248, P1_R1162_U246, P1_R1162_U247);
  nand ginst2332 (P1_R1162_U249, P1_R1162_U222, P1_R1162_U42);
  not ginst2333 (P1_R1162_U25, P1_REG1_REG_2__SCAN_IN);
  nand ginst2334 (P1_R1162_U250, P1_R1162_U137, P1_R1162_U248);
  nand ginst2335 (P1_R1162_U251, P1_R1162_U30, P1_U3466);
  nand ginst2336 (P1_R1162_U252, P1_REG1_REG_3__SCAN_IN, P1_R1162_U31);
  nand ginst2337 (P1_R1162_U253, P1_R1162_U251, P1_R1162_U252);
  nand ginst2338 (P1_R1162_U254, P1_R1162_U223, P1_R1162_U82);
  nand ginst2339 (P1_R1162_U255, P1_R1162_U146, P1_R1162_U253);
  nand ginst2340 (P1_R1162_U256, P1_R1162_U25, P1_U3463);
  nand ginst2341 (P1_R1162_U257, P1_REG1_REG_2__SCAN_IN, P1_R1162_U26);
  nand ginst2342 (P1_R1162_U258, P1_R1162_U83, P1_R1162_U98);
  nand ginst2343 (P1_R1162_U259, P1_R1162_U153, P1_R1162_U29);
  not ginst2344 (P1_R1162_U26, P1_U3463);
  nand ginst2345 (P1_R1162_U260, P1_R1162_U85, P1_U3452);
  nand ginst2346 (P1_R1162_U261, P1_REG1_REG_19__SCAN_IN, P1_R1162_U84);
  nand ginst2347 (P1_R1162_U262, P1_R1162_U85, P1_U3452);
  nand ginst2348 (P1_R1162_U263, P1_REG1_REG_19__SCAN_IN, P1_R1162_U84);
  nand ginst2349 (P1_R1162_U264, P1_R1162_U262, P1_R1162_U263);
  nand ginst2350 (P1_R1162_U265, P1_R1162_U63, P1_U3511);
  nand ginst2351 (P1_R1162_U266, P1_REG1_REG_18__SCAN_IN, P1_R1162_U64);
  nand ginst2352 (P1_R1162_U267, P1_R1162_U63, P1_U3511);
  nand ginst2353 (P1_R1162_U268, P1_REG1_REG_18__SCAN_IN, P1_R1162_U64);
  nand ginst2354 (P1_R1162_U269, P1_R1162_U267, P1_R1162_U268);
  not ginst2355 (P1_R1162_U27, P1_REG1_REG_0__SCAN_IN);
  nand ginst2356 (P1_R1162_U270, P1_R1162_U265, P1_R1162_U266, P1_R1162_U65);
  nand ginst2357 (P1_R1162_U271, P1_R1162_U188, P1_R1162_U269);
  nand ginst2358 (P1_R1162_U272, P1_R1162_U48, P1_U3508);
  nand ginst2359 (P1_R1162_U273, P1_REG1_REG_17__SCAN_IN, P1_R1162_U46);
  nand ginst2360 (P1_R1162_U274, P1_R1162_U44, P1_U3505);
  nand ginst2361 (P1_R1162_U275, P1_REG1_REG_16__SCAN_IN, P1_R1162_U45);
  nand ginst2362 (P1_R1162_U276, P1_R1162_U274, P1_R1162_U275);
  nand ginst2363 (P1_R1162_U277, P1_R1162_U224, P1_R1162_U66);
  nand ginst2364 (P1_R1162_U278, P1_R1162_U180, P1_R1162_U276);
  nand ginst2365 (P1_R1162_U279, P1_R1162_U61, P1_U3502);
  not ginst2366 (P1_R1162_U28, P1_U3454);
  nand ginst2367 (P1_R1162_U280, P1_REG1_REG_15__SCAN_IN, P1_R1162_U62);
  nand ginst2368 (P1_R1162_U281, P1_R1162_U61, P1_U3502);
  nand ginst2369 (P1_R1162_U282, P1_REG1_REG_15__SCAN_IN, P1_R1162_U62);
  nand ginst2370 (P1_R1162_U283, P1_R1162_U281, P1_R1162_U282);
  nand ginst2371 (P1_R1162_U284, P1_R1162_U279, P1_R1162_U280, P1_R1162_U86);
  nand ginst2372 (P1_R1162_U285, P1_R1162_U176, P1_R1162_U283);
  nand ginst2373 (P1_R1162_U286, P1_R1162_U59, P1_U3499);
  nand ginst2374 (P1_R1162_U287, P1_REG1_REG_14__SCAN_IN, P1_R1162_U60);
  nand ginst2375 (P1_R1162_U288, P1_R1162_U59, P1_U3499);
  nand ginst2376 (P1_R1162_U289, P1_REG1_REG_14__SCAN_IN, P1_R1162_U60);
  nand ginst2377 (P1_R1162_U29, P1_REG1_REG_0__SCAN_IN, P1_U3454);
  nand ginst2378 (P1_R1162_U290, P1_R1162_U288, P1_R1162_U289);
  nand ginst2379 (P1_R1162_U291, P1_R1162_U286, P1_R1162_U287, P1_R1162_U87);
  nand ginst2380 (P1_R1162_U292, P1_R1162_U172, P1_R1162_U290);
  nand ginst2381 (P1_R1162_U293, P1_R1162_U57, P1_U3496);
  nand ginst2382 (P1_R1162_U294, P1_REG1_REG_13__SCAN_IN, P1_R1162_U58);
  nand ginst2383 (P1_R1162_U295, P1_R1162_U52, P1_U3493);
  nand ginst2384 (P1_R1162_U296, P1_REG1_REG_12__SCAN_IN, P1_R1162_U53);
  nand ginst2385 (P1_R1162_U297, P1_R1162_U295, P1_R1162_U296);
  nand ginst2386 (P1_R1162_U298, P1_R1162_U225, P1_R1162_U67);
  nand ginst2387 (P1_R1162_U299, P1_R1162_U205, P1_R1162_U297);
  not ginst2388 (P1_R1162_U30, P1_REG1_REG_3__SCAN_IN);
  nand ginst2389 (P1_R1162_U300, P1_R1162_U54, P1_U3490);
  nand ginst2390 (P1_R1162_U301, P1_REG1_REG_11__SCAN_IN, P1_R1162_U55);
  nand ginst2391 (P1_R1162_U302, P1_R1162_U300, P1_R1162_U301);
  nand ginst2392 (P1_R1162_U303, P1_R1162_U226, P1_R1162_U88);
  nand ginst2393 (P1_R1162_U304, P1_R1162_U162, P1_R1162_U302);
  nand ginst2394 (P1_R1162_U305, P1_R1162_U50, P1_U3487);
  nand ginst2395 (P1_R1162_U306, P1_REG1_REG_10__SCAN_IN, P1_R1162_U51);
  nand ginst2396 (P1_R1162_U307, P1_R1162_U27, P1_U3454);
  nand ginst2397 (P1_R1162_U308, P1_REG1_REG_0__SCAN_IN, P1_R1162_U28);
  not ginst2398 (P1_R1162_U31, P1_U3466);
  nand ginst2399 (P1_R1162_U32, P1_REG1_REG_4__SCAN_IN, P1_U3469);
  not ginst2400 (P1_R1162_U33, P1_REG1_REG_5__SCAN_IN);
  not ginst2401 (P1_R1162_U34, P1_REG1_REG_8__SCAN_IN);
  not ginst2402 (P1_R1162_U35, P1_U3481);
  not ginst2403 (P1_R1162_U36, P1_U3484);
  not ginst2404 (P1_R1162_U37, P1_REG1_REG_9__SCAN_IN);
  nand ginst2405 (P1_R1162_U38, P1_R1162_U121, P1_R1162_U49);
  nand ginst2406 (P1_R1162_U39, P1_R1162_U108, P1_R1162_U109, P1_R1162_U110);
  and ginst2407 (P1_R1162_U4, P1_R1162_U94, P1_R1162_U95);
  nand ginst2408 (P1_R1162_U40, P1_R1162_U98, P1_R1162_U99);
  nand ginst2409 (P1_R1162_U41, P1_REG1_REG_1__SCAN_IN, P1_U3460);
  nand ginst2410 (P1_R1162_U42, P1_R1162_U134, P1_R1162_U135, P1_R1162_U136);
  nand ginst2411 (P1_R1162_U43, P1_R1162_U131, P1_R1162_U132);
  not ginst2412 (P1_R1162_U44, P1_REG1_REG_16__SCAN_IN);
  not ginst2413 (P1_R1162_U45, P1_U3505);
  not ginst2414 (P1_R1162_U46, P1_U3508);
  nand ginst2415 (P1_R1162_U47, P1_REG1_REG_16__SCAN_IN, P1_U3505);
  not ginst2416 (P1_R1162_U48, P1_REG1_REG_17__SCAN_IN);
  nand ginst2417 (P1_R1162_U49, P1_REG1_REG_8__SCAN_IN, P1_U3481);
  and ginst2418 (P1_R1162_U5, P1_R1162_U96, P1_R1162_U97);
  not ginst2419 (P1_R1162_U50, P1_REG1_REG_10__SCAN_IN);
  not ginst2420 (P1_R1162_U51, P1_U3487);
  not ginst2421 (P1_R1162_U52, P1_REG1_REG_12__SCAN_IN);
  not ginst2422 (P1_R1162_U53, P1_U3493);
  not ginst2423 (P1_R1162_U54, P1_REG1_REG_11__SCAN_IN);
  not ginst2424 (P1_R1162_U55, P1_U3490);
  nand ginst2425 (P1_R1162_U56, P1_REG1_REG_11__SCAN_IN, P1_U3490);
  not ginst2426 (P1_R1162_U57, P1_REG1_REG_13__SCAN_IN);
  not ginst2427 (P1_R1162_U58, P1_U3496);
  not ginst2428 (P1_R1162_U59, P1_REG1_REG_14__SCAN_IN);
  and ginst2429 (P1_R1162_U6, P1_R1162_U112, P1_R1162_U113);
  not ginst2430 (P1_R1162_U60, P1_U3499);
  not ginst2431 (P1_R1162_U61, P1_REG1_REG_15__SCAN_IN);
  not ginst2432 (P1_R1162_U62, P1_U3502);
  not ginst2433 (P1_R1162_U63, P1_REG1_REG_18__SCAN_IN);
  not ginst2434 (P1_R1162_U64, P1_U3511);
  nand ginst2435 (P1_R1162_U65, P1_R1162_U185, P1_R1162_U186, P1_R1162_U187);
  nand ginst2436 (P1_R1162_U66, P1_R1162_U178, P1_R1162_U179);
  nand ginst2437 (P1_R1162_U67, P1_R1162_U204, P1_R1162_U56);
  nand ginst2438 (P1_R1162_U68, P1_R1162_U258, P1_R1162_U259);
  nand ginst2439 (P1_R1162_U69, P1_R1162_U307, P1_R1162_U308);
  and ginst2440 (P1_R1162_U7, P1_R1162_U154, P1_R1162_U155);
  nand ginst2441 (P1_R1162_U70, P1_R1162_U230, P1_R1162_U231);
  nand ginst2442 (P1_R1162_U71, P1_R1162_U235, P1_R1162_U236);
  nand ginst2443 (P1_R1162_U72, P1_R1162_U242, P1_R1162_U243);
  nand ginst2444 (P1_R1162_U73, P1_R1162_U249, P1_R1162_U250);
  nand ginst2445 (P1_R1162_U74, P1_R1162_U254, P1_R1162_U255);
  nand ginst2446 (P1_R1162_U75, P1_R1162_U270, P1_R1162_U271);
  nand ginst2447 (P1_R1162_U76, P1_R1162_U277, P1_R1162_U278);
  nand ginst2448 (P1_R1162_U77, P1_R1162_U284, P1_R1162_U285);
  nand ginst2449 (P1_R1162_U78, P1_R1162_U291, P1_R1162_U292);
  nand ginst2450 (P1_R1162_U79, P1_R1162_U298, P1_R1162_U299);
  and ginst2451 (P1_R1162_U8, P1_R1162_U163, P1_R1162_U164);
  nand ginst2452 (P1_R1162_U80, P1_R1162_U303, P1_R1162_U304);
  nand ginst2453 (P1_R1162_U81, P1_R1162_U116, P1_R1162_U117, P1_R1162_U118);
  nand ginst2454 (P1_R1162_U82, P1_R1162_U133, P1_R1162_U145);
  nand ginst2455 (P1_R1162_U83, P1_R1162_U152, P1_R1162_U41);
  not ginst2456 (P1_R1162_U84, P1_U3452);
  not ginst2457 (P1_R1162_U85, P1_REG1_REG_19__SCAN_IN);
  nand ginst2458 (P1_R1162_U86, P1_R1162_U174, P1_R1162_U175);
  nand ginst2459 (P1_R1162_U87, P1_R1162_U170, P1_R1162_U171);
  nand ginst2460 (P1_R1162_U88, P1_R1162_U160, P1_R1162_U161);
  not ginst2461 (P1_R1162_U89, P1_R1162_U32);
  and ginst2462 (P1_R1162_U9, P1_R1162_U181, P1_R1162_U182);
  nand ginst2463 (P1_R1162_U90, P1_REG1_REG_9__SCAN_IN, P1_U3484);
  nand ginst2464 (P1_R1162_U91, P1_REG1_REG_12__SCAN_IN, P1_U3493);
  not ginst2465 (P1_R1162_U92, P1_R1162_U56);
  not ginst2466 (P1_R1162_U93, P1_R1162_U49);
  or ginst2467 (P1_R1162_U94, P1_REG1_REG_5__SCAN_IN, P1_U3472);
  or ginst2468 (P1_R1162_U95, P1_REG1_REG_4__SCAN_IN, P1_U3469);
  or ginst2469 (P1_R1162_U96, P1_REG1_REG_3__SCAN_IN, P1_U3466);
  or ginst2470 (P1_R1162_U97, P1_REG1_REG_2__SCAN_IN, P1_U3463);
  not ginst2471 (P1_R1162_U98, P1_R1162_U29);
  or ginst2472 (P1_R1162_U99, P1_REG1_REG_1__SCAN_IN, P1_U3460);
  and ginst2473 (P1_R1165_U10, P1_R1165_U327, P1_R1165_U330);
  nand ginst2474 (P1_R1165_U100, P1_R1165_U530, P1_R1165_U531);
  nand ginst2475 (P1_R1165_U101, P1_R1165_U537, P1_R1165_U538);
  nand ginst2476 (P1_R1165_U102, P1_R1165_U542, P1_R1165_U543);
  nand ginst2477 (P1_R1165_U103, P1_R1165_U549, P1_R1165_U550);
  nand ginst2478 (P1_R1165_U104, P1_R1165_U556, P1_R1165_U557);
  nand ginst2479 (P1_R1165_U105, P1_R1165_U563, P1_R1165_U564);
  nand ginst2480 (P1_R1165_U106, P1_R1165_U570, P1_R1165_U571);
  nand ginst2481 (P1_R1165_U107, P1_R1165_U577, P1_R1165_U578);
  nand ginst2482 (P1_R1165_U108, P1_R1165_U582, P1_R1165_U583);
  nand ginst2483 (P1_R1165_U109, P1_R1165_U589, P1_R1165_U590);
  and ginst2484 (P1_R1165_U11, P1_R1165_U320, P1_R1165_U323);
  and ginst2485 (P1_R1165_U110, P1_R1165_U204, P1_R1165_U205);
  and ginst2486 (P1_R1165_U111, P1_R1165_U220, P1_R1165_U221);
  and ginst2487 (P1_R1165_U112, P1_R1165_U17, P1_R1165_U402, P1_R1165_U403);
  and ginst2488 (P1_R1165_U113, P1_R1165_U232, P1_R1165_U5);
  and ginst2489 (P1_R1165_U114, P1_R1165_U20, P1_R1165_U423, P1_R1165_U424);
  and ginst2490 (P1_R1165_U115, P1_R1165_U239, P1_R1165_U4);
  and ginst2491 (P1_R1165_U116, P1_R1165_U255, P1_R1165_U6);
  and ginst2492 (P1_R1165_U117, P1_R1165_U187, P1_R1165_U253);
  and ginst2493 (P1_R1165_U118, P1_R1165_U272, P1_R1165_U273);
  and ginst2494 (P1_R1165_U119, P1_R1165_U357, P1_R1165_U53);
  and ginst2495 (P1_R1165_U12, P1_R1165_U311, P1_R1165_U314);
  and ginst2496 (P1_R1165_U120, P1_R1165_U301, P1_R1165_U306);
  and ginst2497 (P1_R1165_U121, P1_R1165_U305, P1_R1165_U354);
  nand ginst2498 (P1_R1165_U122, P1_R1165_U484, P1_R1165_U485);
  and ginst2499 (P1_R1165_U123, P1_R1165_U189, P1_R1165_U499, P1_R1165_U500);
  and ginst2500 (P1_R1165_U124, P1_R1165_U188, P1_R1165_U525, P1_R1165_U526);
  and ginst2501 (P1_R1165_U125, P1_R1165_U38, P1_R1165_U551, P1_R1165_U552);
  and ginst2502 (P1_R1165_U126, P1_R1165_U329, P1_R1165_U7);
  and ginst2503 (P1_R1165_U127, P1_R1165_U187, P1_R1165_U572, P1_R1165_U573);
  and ginst2504 (P1_R1165_U128, P1_R1165_U338, P1_R1165_U6);
  nand ginst2505 (P1_R1165_U129, P1_R1165_U591, P1_R1165_U592);
  and ginst2506 (P1_R1165_U13, P1_R1165_U237, P1_R1165_U240);
  not ginst2507 (P1_R1165_U130, P1_U3201);
  and ginst2508 (P1_R1165_U131, P1_R1165_U361, P1_R1165_U362);
  not ginst2509 (P1_R1165_U132, P1_U3210);
  not ginst2510 (P1_R1165_U133, P1_U3209);
  not ginst2511 (P1_R1165_U134, P1_U3207);
  not ginst2512 (P1_R1165_U135, P1_U3208);
  not ginst2513 (P1_R1165_U136, P1_U3206);
  not ginst2514 (P1_R1165_U137, P1_U3205);
  not ginst2515 (P1_R1165_U138, P1_U3203);
  not ginst2516 (P1_R1165_U139, P1_U3204);
  and ginst2517 (P1_R1165_U14, P1_R1165_U230, P1_R1165_U233);
  not ginst2518 (P1_R1165_U140, P1_U3202);
  and ginst2519 (P1_R1165_U141, P1_R1165_U395, P1_R1165_U396);
  nand ginst2520 (P1_R1165_U142, P1_R1165_U111, P1_R1165_U222);
  and ginst2521 (P1_R1165_U143, P1_R1165_U409, P1_R1165_U410);
  nand ginst2522 (P1_R1165_U144, P1_R1165_U209, P1_R1165_U210);
  and ginst2523 (P1_R1165_U145, P1_R1165_U416, P1_R1165_U417);
  not ginst2524 (P1_R1165_U146, P1_U3183);
  not ginst2525 (P1_R1165_U147, P1_U3185);
  not ginst2526 (P1_R1165_U148, P1_U3184);
  not ginst2527 (P1_R1165_U149, P1_U3186);
  not ginst2528 (P1_R1165_U15, P1_U3211);
  not ginst2529 (P1_R1165_U150, P1_U3189);
  not ginst2530 (P1_R1165_U151, P1_U3190);
  not ginst2531 (P1_R1165_U152, P1_U3191);
  not ginst2532 (P1_R1165_U153, P1_U3200);
  not ginst2533 (P1_R1165_U154, P1_U3197);
  not ginst2534 (P1_R1165_U155, P1_U3198);
  not ginst2535 (P1_R1165_U156, P1_U3199);
  not ginst2536 (P1_R1165_U157, P1_U3196);
  not ginst2537 (P1_R1165_U158, P1_U3195);
  not ginst2538 (P1_R1165_U159, P1_U3193);
  not ginst2539 (P1_R1165_U16, P1_U3175);
  not ginst2540 (P1_R1165_U160, P1_U3194);
  not ginst2541 (P1_R1165_U161, P1_U3192);
  not ginst2542 (P1_R1165_U162, P1_U3188);
  not ginst2543 (P1_R1165_U163, P1_U3187);
  not ginst2544 (P1_R1165_U164, P1_U3153);
  not ginst2545 (P1_R1165_U165, P1_U3182);
  and ginst2546 (P1_R1165_U166, P1_R1165_U492, P1_R1165_U493);
  nand ginst2547 (P1_R1165_U167, P1_R1165_U302, P1_R1165_U351, P1_R1165_U53);
  nand ginst2548 (P1_R1165_U168, P1_R1165_U295, P1_R1165_U296);
  and ginst2549 (P1_R1165_U169, P1_R1165_U511, P1_R1165_U512);
  nand ginst2550 (P1_R1165_U17, P1_R1165_U59, P1_U3175);
  nand ginst2551 (P1_R1165_U170, P1_R1165_U291, P1_R1165_U292);
  and ginst2552 (P1_R1165_U171, P1_R1165_U518, P1_R1165_U519);
  nand ginst2553 (P1_R1165_U172, P1_R1165_U283, P1_R1165_U287, P1_R1165_U288);
  and ginst2554 (P1_R1165_U173, P1_R1165_U532, P1_R1165_U533);
  nand ginst2555 (P1_R1165_U174, P1_R1165_U194, P1_R1165_U195);
  nand ginst2556 (P1_R1165_U175, P1_R1165_U277, P1_R1165_U278);
  and ginst2557 (P1_R1165_U176, P1_R1165_U544, P1_R1165_U545);
  nand ginst2558 (P1_R1165_U177, P1_R1165_U118, P1_R1165_U274);
  and ginst2559 (P1_R1165_U178, P1_R1165_U558, P1_R1165_U559);
  nand ginst2560 (P1_R1165_U179, P1_R1165_U261, P1_R1165_U262);
  not ginst2561 (P1_R1165_U18, P1_U3174);
  and ginst2562 (P1_R1165_U180, P1_R1165_U565, P1_R1165_U566);
  nand ginst2563 (P1_R1165_U181, P1_R1165_U257, P1_R1165_U258);
  nand ginst2564 (P1_R1165_U182, P1_R1165_U247, P1_R1165_U248);
  and ginst2565 (P1_R1165_U183, P1_R1165_U584, P1_R1165_U585);
  nand ginst2566 (P1_R1165_U184, P1_R1165_U243, P1_R1165_U244);
  nand ginst2567 (P1_R1165_U185, P1_R1165_U352, P1_R1165_U353);
  not ginst2568 (P1_R1165_U186, P1_R1165_U20);
  nand ginst2569 (P1_R1165_U187, P1_R1165_U78, P1_U3169);
  nand ginst2570 (P1_R1165_U188, P1_R1165_U83, P1_U3161);
  nand ginst2571 (P1_R1165_U189, P1_R1165_U69, P1_U3156);
  not ginst2572 (P1_R1165_U19, P1_U3179);
  not ginst2573 (P1_R1165_U190, P1_R1165_U43);
  not ginst2574 (P1_R1165_U191, P1_R1165_U49);
  nand ginst2575 (P1_R1165_U192, P1_R1165_U71, P1_U3157);
  or ginst2576 (P1_R1165_U193, P1_U3181, P1_U3211);
  nand ginst2577 (P1_R1165_U194, P1_R1165_U193, P1_R1165_U63);
  nand ginst2578 (P1_R1165_U195, P1_U3181, P1_U3211);
  not ginst2579 (P1_R1165_U196, P1_R1165_U174);
  nand ginst2580 (P1_R1165_U197, P1_R1165_U23, P1_R1165_U371);
  nand ginst2581 (P1_R1165_U198, P1_R1165_U174, P1_R1165_U197);
  nand ginst2582 (P1_R1165_U199, P1_R1165_U64, P1_U3180);
  nand ginst2583 (P1_R1165_U20, P1_R1165_U61, P1_U3179);
  not ginst2584 (P1_R1165_U200, P1_R1165_U31);
  nand ginst2585 (P1_R1165_U201, P1_R1165_U21, P1_R1165_U374);
  nand ginst2586 (P1_R1165_U202, P1_R1165_U19, P1_R1165_U377);
  nand ginst2587 (P1_R1165_U203, P1_R1165_U20, P1_R1165_U21);
  nand ginst2588 (P1_R1165_U204, P1_R1165_U203, P1_R1165_U62);
  nand ginst2589 (P1_R1165_U205, P1_R1165_U186, P1_U3178);
  nand ginst2590 (P1_R1165_U206, P1_R1165_U31, P1_R1165_U4);
  not ginst2591 (P1_R1165_U207, P1_R1165_U24);
  nand ginst2592 (P1_R1165_U208, P1_R1165_U207, P1_R1165_U25);
  nand ginst2593 (P1_R1165_U209, P1_R1165_U208, P1_R1165_U65);
  not ginst2594 (P1_R1165_U21, P1_U3178);
  nand ginst2595 (P1_R1165_U210, P1_R1165_U24, P1_U3177);
  not ginst2596 (P1_R1165_U211, P1_R1165_U144);
  nand ginst2597 (P1_R1165_U212, P1_R1165_U26, P1_R1165_U383);
  nand ginst2598 (P1_R1165_U213, P1_R1165_U144, P1_R1165_U212);
  nand ginst2599 (P1_R1165_U214, P1_R1165_U66, P1_U3176);
  not ginst2600 (P1_R1165_U215, P1_R1165_U30);
  nand ginst2601 (P1_R1165_U216, P1_R1165_U18, P1_R1165_U386);
  nand ginst2602 (P1_R1165_U217, P1_R1165_U16, P1_R1165_U389);
  not ginst2603 (P1_R1165_U218, P1_R1165_U17);
  nand ginst2604 (P1_R1165_U219, P1_R1165_U17, P1_R1165_U18);
  not ginst2605 (P1_R1165_U22, P1_U3181);
  nand ginst2606 (P1_R1165_U220, P1_R1165_U219, P1_R1165_U60);
  nand ginst2607 (P1_R1165_U221, P1_R1165_U218, P1_U3174);
  nand ginst2608 (P1_R1165_U222, P1_R1165_U30, P1_R1165_U5);
  not ginst2609 (P1_R1165_U223, P1_R1165_U142);
  nand ginst2610 (P1_R1165_U224, P1_R1165_U27, P1_R1165_U392);
  nand ginst2611 (P1_R1165_U225, P1_R1165_U142, P1_R1165_U224);
  nand ginst2612 (P1_R1165_U226, P1_R1165_U67, P1_U3173);
  not ginst2613 (P1_R1165_U227, P1_R1165_U29);
  nand ginst2614 (P1_R1165_U228, P1_R1165_U16, P1_R1165_U389);
  nand ginst2615 (P1_R1165_U229, P1_R1165_U228, P1_R1165_U30);
  not ginst2616 (P1_R1165_U23, P1_U3180);
  nand ginst2617 (P1_R1165_U230, P1_R1165_U112, P1_R1165_U229);
  nand ginst2618 (P1_R1165_U231, P1_R1165_U17, P1_R1165_U215);
  nand ginst2619 (P1_R1165_U232, P1_R1165_U60, P1_U3174);
  nand ginst2620 (P1_R1165_U233, P1_R1165_U113, P1_R1165_U231);
  nand ginst2621 (P1_R1165_U234, P1_R1165_U16, P1_R1165_U389);
  nand ginst2622 (P1_R1165_U235, P1_R1165_U19, P1_R1165_U377);
  nand ginst2623 (P1_R1165_U236, P1_R1165_U235, P1_R1165_U31);
  nand ginst2624 (P1_R1165_U237, P1_R1165_U114, P1_R1165_U236);
  nand ginst2625 (P1_R1165_U238, P1_R1165_U20, P1_R1165_U200);
  nand ginst2626 (P1_R1165_U239, P1_R1165_U62, P1_U3178);
  nand ginst2627 (P1_R1165_U24, P1_R1165_U110, P1_R1165_U206);
  nand ginst2628 (P1_R1165_U240, P1_R1165_U115, P1_R1165_U238);
  nand ginst2629 (P1_R1165_U241, P1_R1165_U19, P1_R1165_U377);
  nand ginst2630 (P1_R1165_U242, P1_R1165_U227, P1_R1165_U28);
  nand ginst2631 (P1_R1165_U243, P1_R1165_U242, P1_R1165_U58);
  nand ginst2632 (P1_R1165_U244, P1_R1165_U29, P1_U3172);
  not ginst2633 (P1_R1165_U245, P1_R1165_U184);
  nand ginst2634 (P1_R1165_U246, P1_R1165_U40, P1_R1165_U453);
  nand ginst2635 (P1_R1165_U247, P1_R1165_U184, P1_R1165_U246);
  nand ginst2636 (P1_R1165_U248, P1_R1165_U75, P1_U3171);
  not ginst2637 (P1_R1165_U249, P1_R1165_U182);
  not ginst2638 (P1_R1165_U25, P1_U3177);
  nand ginst2639 (P1_R1165_U250, P1_R1165_U44, P1_R1165_U456);
  nand ginst2640 (P1_R1165_U251, P1_R1165_U41, P1_R1165_U459);
  nand ginst2641 (P1_R1165_U252, P1_R1165_U190, P1_R1165_U6);
  nand ginst2642 (P1_R1165_U253, P1_R1165_U77, P1_U3168);
  nand ginst2643 (P1_R1165_U254, P1_R1165_U117, P1_R1165_U252);
  nand ginst2644 (P1_R1165_U255, P1_R1165_U42, P1_R1165_U462);
  nand ginst2645 (P1_R1165_U256, P1_R1165_U44, P1_R1165_U456);
  nand ginst2646 (P1_R1165_U257, P1_R1165_U116, P1_R1165_U182);
  nand ginst2647 (P1_R1165_U258, P1_R1165_U254, P1_R1165_U256);
  not ginst2648 (P1_R1165_U259, P1_R1165_U181);
  not ginst2649 (P1_R1165_U26, P1_U3176);
  nand ginst2650 (P1_R1165_U260, P1_R1165_U45, P1_R1165_U465);
  nand ginst2651 (P1_R1165_U261, P1_R1165_U181, P1_R1165_U260);
  nand ginst2652 (P1_R1165_U262, P1_R1165_U79, P1_U3167);
  not ginst2653 (P1_R1165_U263, P1_R1165_U179);
  nand ginst2654 (P1_R1165_U264, P1_R1165_U46, P1_R1165_U468);
  nand ginst2655 (P1_R1165_U265, P1_R1165_U179, P1_R1165_U264);
  nand ginst2656 (P1_R1165_U266, P1_R1165_U80, P1_U3166);
  not ginst2657 (P1_R1165_U267, P1_R1165_U56);
  nand ginst2658 (P1_R1165_U268, P1_R1165_U39, P1_R1165_U471);
  nand ginst2659 (P1_R1165_U269, P1_R1165_U37, P1_R1165_U474);
  not ginst2660 (P1_R1165_U27, P1_U3173);
  not ginst2661 (P1_R1165_U270, P1_R1165_U38);
  nand ginst2662 (P1_R1165_U271, P1_R1165_U38, P1_R1165_U39);
  nand ginst2663 (P1_R1165_U272, P1_R1165_U271, P1_R1165_U74);
  nand ginst2664 (P1_R1165_U273, P1_R1165_U270, P1_U3164);
  nand ginst2665 (P1_R1165_U274, P1_R1165_U56, P1_R1165_U7);
  not ginst2666 (P1_R1165_U275, P1_R1165_U177);
  nand ginst2667 (P1_R1165_U276, P1_R1165_U47, P1_R1165_U477);
  nand ginst2668 (P1_R1165_U277, P1_R1165_U177, P1_R1165_U276);
  nand ginst2669 (P1_R1165_U278, P1_R1165_U81, P1_U3163);
  not ginst2670 (P1_R1165_U279, P1_R1165_U175);
  not ginst2671 (P1_R1165_U28, P1_U3172);
  nand ginst2672 (P1_R1165_U280, P1_R1165_U36, P1_R1165_U444);
  nand ginst2673 (P1_R1165_U281, P1_R1165_U447, P1_R1165_U50);
  nand ginst2674 (P1_R1165_U282, P1_R1165_U191, P1_R1165_U8);
  nand ginst2675 (P1_R1165_U283, P1_R1165_U72, P1_U3160);
  nand ginst2676 (P1_R1165_U284, P1_R1165_U188, P1_R1165_U282);
  nand ginst2677 (P1_R1165_U285, P1_R1165_U450, P1_R1165_U48);
  nand ginst2678 (P1_R1165_U286, P1_R1165_U36, P1_R1165_U444);
  nand ginst2679 (P1_R1165_U287, P1_R1165_U175, P1_R1165_U285, P1_R1165_U8);
  nand ginst2680 (P1_R1165_U288, P1_R1165_U284, P1_R1165_U286);
  not ginst2681 (P1_R1165_U289, P1_R1165_U172);
  nand ginst2682 (P1_R1165_U29, P1_R1165_U225, P1_R1165_U226);
  nand ginst2683 (P1_R1165_U290, P1_R1165_U480, P1_R1165_U51);
  nand ginst2684 (P1_R1165_U291, P1_R1165_U172, P1_R1165_U290);
  nand ginst2685 (P1_R1165_U292, P1_R1165_U84, P1_U3159);
  not ginst2686 (P1_R1165_U293, P1_R1165_U170);
  nand ginst2687 (P1_R1165_U294, P1_R1165_U483, P1_R1165_U52);
  nand ginst2688 (P1_R1165_U295, P1_R1165_U170, P1_R1165_U294);
  nand ginst2689 (P1_R1165_U296, P1_R1165_U85, P1_U3158);
  not ginst2690 (P1_R1165_U297, P1_R1165_U168);
  nand ginst2691 (P1_R1165_U298, P1_R1165_U34, P1_R1165_U435);
  nand ginst2692 (P1_R1165_U299, P1_R1165_U189, P1_R1165_U192);
  nand ginst2693 (P1_R1165_U30, P1_R1165_U213, P1_R1165_U214);
  not ginst2694 (P1_R1165_U300, P1_R1165_U53);
  nand ginst2695 (P1_R1165_U301, P1_R1165_U35, P1_R1165_U441);
  nand ginst2696 (P1_R1165_U302, P1_R1165_U168, P1_R1165_U185, P1_R1165_U301);
  not ginst2697 (P1_R1165_U303, P1_R1165_U167);
  nand ginst2698 (P1_R1165_U304, P1_R1165_U32, P1_R1165_U432);
  nand ginst2699 (P1_R1165_U305, P1_R1165_U68, P1_U3154);
  nand ginst2700 (P1_R1165_U306, P1_R1165_U32, P1_R1165_U432);
  nand ginst2701 (P1_R1165_U307, P1_R1165_U168, P1_R1165_U301);
  not ginst2702 (P1_R1165_U308, P1_R1165_U54);
  nand ginst2703 (P1_R1165_U309, P1_R1165_U34, P1_R1165_U435);
  nand ginst2704 (P1_R1165_U31, P1_R1165_U198, P1_R1165_U199);
  nand ginst2705 (P1_R1165_U310, P1_R1165_U309, P1_R1165_U54);
  nand ginst2706 (P1_R1165_U311, P1_R1165_U123, P1_R1165_U310);
  nand ginst2707 (P1_R1165_U312, P1_R1165_U189, P1_R1165_U308);
  nand ginst2708 (P1_R1165_U313, P1_R1165_U70, P1_U3155);
  nand ginst2709 (P1_R1165_U314, P1_R1165_U185, P1_R1165_U312, P1_R1165_U313);
  nand ginst2710 (P1_R1165_U315, P1_R1165_U34, P1_R1165_U435);
  nand ginst2711 (P1_R1165_U316, P1_R1165_U175, P1_R1165_U285);
  not ginst2712 (P1_R1165_U317, P1_R1165_U55);
  nand ginst2713 (P1_R1165_U318, P1_R1165_U447, P1_R1165_U50);
  nand ginst2714 (P1_R1165_U319, P1_R1165_U318, P1_R1165_U55);
  not ginst2715 (P1_R1165_U32, P1_U3154);
  nand ginst2716 (P1_R1165_U320, P1_R1165_U124, P1_R1165_U319);
  nand ginst2717 (P1_R1165_U321, P1_R1165_U188, P1_R1165_U317);
  nand ginst2718 (P1_R1165_U322, P1_R1165_U72, P1_U3160);
  nand ginst2719 (P1_R1165_U323, P1_R1165_U321, P1_R1165_U322, P1_R1165_U8);
  nand ginst2720 (P1_R1165_U324, P1_R1165_U447, P1_R1165_U50);
  nand ginst2721 (P1_R1165_U325, P1_R1165_U37, P1_R1165_U474);
  nand ginst2722 (P1_R1165_U326, P1_R1165_U325, P1_R1165_U56);
  nand ginst2723 (P1_R1165_U327, P1_R1165_U125, P1_R1165_U326);
  nand ginst2724 (P1_R1165_U328, P1_R1165_U267, P1_R1165_U38);
  nand ginst2725 (P1_R1165_U329, P1_R1165_U74, P1_U3164);
  not ginst2726 (P1_R1165_U33, P1_U3155);
  nand ginst2727 (P1_R1165_U330, P1_R1165_U126, P1_R1165_U328);
  nand ginst2728 (P1_R1165_U331, P1_R1165_U37, P1_R1165_U474);
  nand ginst2729 (P1_R1165_U332, P1_R1165_U182, P1_R1165_U255);
  not ginst2730 (P1_R1165_U333, P1_R1165_U57);
  nand ginst2731 (P1_R1165_U334, P1_R1165_U41, P1_R1165_U459);
  nand ginst2732 (P1_R1165_U335, P1_R1165_U334, P1_R1165_U57);
  nand ginst2733 (P1_R1165_U336, P1_R1165_U127, P1_R1165_U335);
  nand ginst2734 (P1_R1165_U337, P1_R1165_U187, P1_R1165_U333);
  nand ginst2735 (P1_R1165_U338, P1_R1165_U77, P1_U3168);
  nand ginst2736 (P1_R1165_U339, P1_R1165_U128, P1_R1165_U337);
  not ginst2737 (P1_R1165_U34, P1_U3156);
  nand ginst2738 (P1_R1165_U340, P1_R1165_U41, P1_R1165_U459);
  nand ginst2739 (P1_R1165_U341, P1_R1165_U17, P1_R1165_U234);
  nand ginst2740 (P1_R1165_U342, P1_R1165_U20, P1_R1165_U241);
  nand ginst2741 (P1_R1165_U343, P1_R1165_U189, P1_R1165_U315);
  nand ginst2742 (P1_R1165_U344, P1_R1165_U192, P1_R1165_U301);
  nand ginst2743 (P1_R1165_U345, P1_R1165_U188, P1_R1165_U324);
  nand ginst2744 (P1_R1165_U346, P1_R1165_U285, P1_R1165_U49);
  nand ginst2745 (P1_R1165_U347, P1_R1165_U331, P1_R1165_U38);
  nand ginst2746 (P1_R1165_U348, P1_R1165_U187, P1_R1165_U340);
  nand ginst2747 (P1_R1165_U349, P1_R1165_U255, P1_R1165_U43);
  not ginst2748 (P1_R1165_U35, P1_U3157);
  nand ginst2749 (P1_R1165_U350, P1_R1165_U119, P1_R1165_U302, P1_R1165_U351);
  nand ginst2750 (P1_R1165_U351, P1_R1165_U185, P1_R1165_U299);
  nand ginst2751 (P1_R1165_U352, P1_R1165_U298, P1_R1165_U70);
  nand ginst2752 (P1_R1165_U353, P1_R1165_U298, P1_U3155);
  nand ginst2753 (P1_R1165_U354, P1_R1165_U185, P1_R1165_U299, P1_R1165_U306);
  nand ginst2754 (P1_R1165_U355, P1_R1165_U120, P1_R1165_U168, P1_R1165_U185);
  nand ginst2755 (P1_R1165_U356, P1_R1165_U300, P1_R1165_U306);
  nand ginst2756 (P1_R1165_U357, P1_R1165_U68, P1_U3154);
  nand ginst2757 (P1_R1165_U358, P1_R1165_U130, P1_U3211);
  nand ginst2758 (P1_R1165_U359, P1_R1165_U15, P1_U3201);
  not ginst2759 (P1_R1165_U36, P1_U3160);
  not ginst2760 (P1_R1165_U360, P1_R1165_U58);
  nand ginst2761 (P1_R1165_U361, P1_R1165_U360, P1_U3172);
  nand ginst2762 (P1_R1165_U362, P1_R1165_U28, P1_R1165_U58);
  nand ginst2763 (P1_R1165_U363, P1_R1165_U360, P1_U3172);
  nand ginst2764 (P1_R1165_U364, P1_R1165_U28, P1_R1165_U58);
  nand ginst2765 (P1_R1165_U365, P1_R1165_U363, P1_R1165_U364);
  nand ginst2766 (P1_R1165_U366, P1_R1165_U132, P1_U3211);
  nand ginst2767 (P1_R1165_U367, P1_R1165_U15, P1_U3210);
  not ginst2768 (P1_R1165_U368, P1_R1165_U63);
  nand ginst2769 (P1_R1165_U369, P1_R1165_U133, P1_U3211);
  not ginst2770 (P1_R1165_U37, P1_U3165);
  nand ginst2771 (P1_R1165_U370, P1_R1165_U15, P1_U3209);
  not ginst2772 (P1_R1165_U371, P1_R1165_U64);
  nand ginst2773 (P1_R1165_U372, P1_R1165_U134, P1_U3211);
  nand ginst2774 (P1_R1165_U373, P1_R1165_U15, P1_U3207);
  not ginst2775 (P1_R1165_U374, P1_R1165_U62);
  nand ginst2776 (P1_R1165_U375, P1_R1165_U135, P1_U3211);
  nand ginst2777 (P1_R1165_U376, P1_R1165_U15, P1_U3208);
  not ginst2778 (P1_R1165_U377, P1_R1165_U61);
  nand ginst2779 (P1_R1165_U378, P1_R1165_U136, P1_U3211);
  nand ginst2780 (P1_R1165_U379, P1_R1165_U15, P1_U3206);
  nand ginst2781 (P1_R1165_U38, P1_R1165_U73, P1_U3165);
  not ginst2782 (P1_R1165_U380, P1_R1165_U65);
  nand ginst2783 (P1_R1165_U381, P1_R1165_U137, P1_U3211);
  nand ginst2784 (P1_R1165_U382, P1_R1165_U15, P1_U3205);
  not ginst2785 (P1_R1165_U383, P1_R1165_U66);
  nand ginst2786 (P1_R1165_U384, P1_R1165_U138, P1_U3211);
  nand ginst2787 (P1_R1165_U385, P1_R1165_U15, P1_U3203);
  not ginst2788 (P1_R1165_U386, P1_R1165_U60);
  nand ginst2789 (P1_R1165_U387, P1_R1165_U139, P1_U3211);
  nand ginst2790 (P1_R1165_U388, P1_R1165_U15, P1_U3204);
  not ginst2791 (P1_R1165_U389, P1_R1165_U59);
  not ginst2792 (P1_R1165_U39, P1_U3164);
  nand ginst2793 (P1_R1165_U390, P1_R1165_U140, P1_U3211);
  nand ginst2794 (P1_R1165_U391, P1_R1165_U15, P1_U3202);
  not ginst2795 (P1_R1165_U392, P1_R1165_U67);
  nand ginst2796 (P1_R1165_U393, P1_R1165_U131, P1_R1165_U29);
  nand ginst2797 (P1_R1165_U394, P1_R1165_U227, P1_R1165_U365);
  nand ginst2798 (P1_R1165_U395, P1_R1165_U392, P1_U3173);
  nand ginst2799 (P1_R1165_U396, P1_R1165_U27, P1_R1165_U67);
  nand ginst2800 (P1_R1165_U397, P1_R1165_U392, P1_U3173);
  nand ginst2801 (P1_R1165_U398, P1_R1165_U27, P1_R1165_U67);
  nand ginst2802 (P1_R1165_U399, P1_R1165_U397, P1_R1165_U398);
  and ginst2803 (P1_R1165_U4, P1_R1165_U201, P1_R1165_U202);
  not ginst2804 (P1_R1165_U40, P1_U3171);
  nand ginst2805 (P1_R1165_U400, P1_R1165_U141, P1_R1165_U142);
  nand ginst2806 (P1_R1165_U401, P1_R1165_U223, P1_R1165_U399);
  nand ginst2807 (P1_R1165_U402, P1_R1165_U386, P1_U3174);
  nand ginst2808 (P1_R1165_U403, P1_R1165_U18, P1_R1165_U60);
  nand ginst2809 (P1_R1165_U404, P1_R1165_U389, P1_U3175);
  nand ginst2810 (P1_R1165_U405, P1_R1165_U16, P1_R1165_U59);
  nand ginst2811 (P1_R1165_U406, P1_R1165_U404, P1_R1165_U405);
  nand ginst2812 (P1_R1165_U407, P1_R1165_U30, P1_R1165_U341);
  nand ginst2813 (P1_R1165_U408, P1_R1165_U215, P1_R1165_U406);
  nand ginst2814 (P1_R1165_U409, P1_R1165_U383, P1_U3176);
  not ginst2815 (P1_R1165_U41, P1_U3169);
  nand ginst2816 (P1_R1165_U410, P1_R1165_U26, P1_R1165_U66);
  nand ginst2817 (P1_R1165_U411, P1_R1165_U383, P1_U3176);
  nand ginst2818 (P1_R1165_U412, P1_R1165_U26, P1_R1165_U66);
  nand ginst2819 (P1_R1165_U413, P1_R1165_U411, P1_R1165_U412);
  nand ginst2820 (P1_R1165_U414, P1_R1165_U143, P1_R1165_U144);
  nand ginst2821 (P1_R1165_U415, P1_R1165_U211, P1_R1165_U413);
  nand ginst2822 (P1_R1165_U416, P1_R1165_U380, P1_U3177);
  nand ginst2823 (P1_R1165_U417, P1_R1165_U25, P1_R1165_U65);
  nand ginst2824 (P1_R1165_U418, P1_R1165_U380, P1_U3177);
  nand ginst2825 (P1_R1165_U419, P1_R1165_U25, P1_R1165_U65);
  not ginst2826 (P1_R1165_U42, P1_U3170);
  nand ginst2827 (P1_R1165_U420, P1_R1165_U418, P1_R1165_U419);
  nand ginst2828 (P1_R1165_U421, P1_R1165_U145, P1_R1165_U24);
  nand ginst2829 (P1_R1165_U422, P1_R1165_U207, P1_R1165_U420);
  nand ginst2830 (P1_R1165_U423, P1_R1165_U374, P1_U3178);
  nand ginst2831 (P1_R1165_U424, P1_R1165_U21, P1_R1165_U62);
  nand ginst2832 (P1_R1165_U425, P1_R1165_U377, P1_U3179);
  nand ginst2833 (P1_R1165_U426, P1_R1165_U19, P1_R1165_U61);
  nand ginst2834 (P1_R1165_U427, P1_R1165_U425, P1_R1165_U426);
  nand ginst2835 (P1_R1165_U428, P1_R1165_U31, P1_R1165_U342);
  nand ginst2836 (P1_R1165_U429, P1_R1165_U200, P1_R1165_U427);
  nand ginst2837 (P1_R1165_U43, P1_R1165_U76, P1_U3170);
  nand ginst2838 (P1_R1165_U430, P1_R1165_U146, P1_U3211);
  nand ginst2839 (P1_R1165_U431, P1_R1165_U15, P1_U3183);
  not ginst2840 (P1_R1165_U432, P1_R1165_U68);
  nand ginst2841 (P1_R1165_U433, P1_R1165_U147, P1_U3211);
  nand ginst2842 (P1_R1165_U434, P1_R1165_U15, P1_U3185);
  not ginst2843 (P1_R1165_U435, P1_R1165_U69);
  nand ginst2844 (P1_R1165_U436, P1_R1165_U148, P1_U3211);
  nand ginst2845 (P1_R1165_U437, P1_R1165_U15, P1_U3184);
  not ginst2846 (P1_R1165_U438, P1_R1165_U70);
  nand ginst2847 (P1_R1165_U439, P1_R1165_U149, P1_U3211);
  not ginst2848 (P1_R1165_U44, P1_U3168);
  nand ginst2849 (P1_R1165_U440, P1_R1165_U15, P1_U3186);
  not ginst2850 (P1_R1165_U441, P1_R1165_U71);
  nand ginst2851 (P1_R1165_U442, P1_R1165_U150, P1_U3211);
  nand ginst2852 (P1_R1165_U443, P1_R1165_U15, P1_U3189);
  not ginst2853 (P1_R1165_U444, P1_R1165_U72);
  nand ginst2854 (P1_R1165_U445, P1_R1165_U151, P1_U3211);
  nand ginst2855 (P1_R1165_U446, P1_R1165_U15, P1_U3190);
  not ginst2856 (P1_R1165_U447, P1_R1165_U83);
  nand ginst2857 (P1_R1165_U448, P1_R1165_U152, P1_U3211);
  nand ginst2858 (P1_R1165_U449, P1_R1165_U15, P1_U3191);
  not ginst2859 (P1_R1165_U45, P1_U3167);
  not ginst2860 (P1_R1165_U450, P1_R1165_U82);
  nand ginst2861 (P1_R1165_U451, P1_R1165_U153, P1_U3211);
  nand ginst2862 (P1_R1165_U452, P1_R1165_U15, P1_U3200);
  not ginst2863 (P1_R1165_U453, P1_R1165_U75);
  nand ginst2864 (P1_R1165_U454, P1_R1165_U154, P1_U3211);
  nand ginst2865 (P1_R1165_U455, P1_R1165_U15, P1_U3197);
  not ginst2866 (P1_R1165_U456, P1_R1165_U77);
  nand ginst2867 (P1_R1165_U457, P1_R1165_U155, P1_U3211);
  nand ginst2868 (P1_R1165_U458, P1_R1165_U15, P1_U3198);
  not ginst2869 (P1_R1165_U459, P1_R1165_U78);
  not ginst2870 (P1_R1165_U46, P1_U3166);
  nand ginst2871 (P1_R1165_U460, P1_R1165_U156, P1_U3211);
  nand ginst2872 (P1_R1165_U461, P1_R1165_U15, P1_U3199);
  not ginst2873 (P1_R1165_U462, P1_R1165_U76);
  nand ginst2874 (P1_R1165_U463, P1_R1165_U157, P1_U3211);
  nand ginst2875 (P1_R1165_U464, P1_R1165_U15, P1_U3196);
  not ginst2876 (P1_R1165_U465, P1_R1165_U79);
  nand ginst2877 (P1_R1165_U466, P1_R1165_U158, P1_U3211);
  nand ginst2878 (P1_R1165_U467, P1_R1165_U15, P1_U3195);
  not ginst2879 (P1_R1165_U468, P1_R1165_U80);
  nand ginst2880 (P1_R1165_U469, P1_R1165_U159, P1_U3211);
  not ginst2881 (P1_R1165_U47, P1_U3163);
  nand ginst2882 (P1_R1165_U470, P1_R1165_U15, P1_U3193);
  not ginst2883 (P1_R1165_U471, P1_R1165_U74);
  nand ginst2884 (P1_R1165_U472, P1_R1165_U160, P1_U3211);
  nand ginst2885 (P1_R1165_U473, P1_R1165_U15, P1_U3194);
  not ginst2886 (P1_R1165_U474, P1_R1165_U73);
  nand ginst2887 (P1_R1165_U475, P1_R1165_U161, P1_U3211);
  nand ginst2888 (P1_R1165_U476, P1_R1165_U15, P1_U3192);
  not ginst2889 (P1_R1165_U477, P1_R1165_U81);
  nand ginst2890 (P1_R1165_U478, P1_R1165_U162, P1_U3211);
  nand ginst2891 (P1_R1165_U479, P1_R1165_U15, P1_U3188);
  not ginst2892 (P1_R1165_U48, P1_U3162);
  not ginst2893 (P1_R1165_U480, P1_R1165_U84);
  nand ginst2894 (P1_R1165_U481, P1_R1165_U163, P1_U3211);
  nand ginst2895 (P1_R1165_U482, P1_R1165_U15, P1_U3187);
  not ginst2896 (P1_R1165_U483, P1_R1165_U85);
  nand ginst2897 (P1_R1165_U484, P1_R1165_U164, P1_U3211);
  nand ginst2898 (P1_R1165_U485, P1_R1165_U15, P1_U3153);
  not ginst2899 (P1_R1165_U486, P1_R1165_U122);
  nand ginst2900 (P1_R1165_U487, P1_R1165_U486, P1_U3182);
  nand ginst2901 (P1_R1165_U488, P1_R1165_U122, P1_R1165_U165);
  not ginst2902 (P1_R1165_U489, P1_R1165_U86);
  nand ginst2903 (P1_R1165_U49, P1_R1165_U82, P1_U3162);
  nand ginst2904 (P1_R1165_U490, P1_R1165_U304, P1_R1165_U350, P1_R1165_U489);
  nand ginst2905 (P1_R1165_U491, P1_R1165_U121, P1_R1165_U355, P1_R1165_U356, P1_R1165_U86);
  nand ginst2906 (P1_R1165_U492, P1_R1165_U432, P1_U3154);
  nand ginst2907 (P1_R1165_U493, P1_R1165_U32, P1_R1165_U68);
  nand ginst2908 (P1_R1165_U494, P1_R1165_U432, P1_U3154);
  nand ginst2909 (P1_R1165_U495, P1_R1165_U32, P1_R1165_U68);
  nand ginst2910 (P1_R1165_U496, P1_R1165_U494, P1_R1165_U495);
  nand ginst2911 (P1_R1165_U497, P1_R1165_U166, P1_R1165_U167);
  nand ginst2912 (P1_R1165_U498, P1_R1165_U303, P1_R1165_U496);
  nand ginst2913 (P1_R1165_U499, P1_R1165_U438, P1_U3155);
  and ginst2914 (P1_R1165_U5, P1_R1165_U216, P1_R1165_U217);
  not ginst2915 (P1_R1165_U50, P1_U3161);
  nand ginst2916 (P1_R1165_U500, P1_R1165_U33, P1_R1165_U70);
  nand ginst2917 (P1_R1165_U501, P1_R1165_U435, P1_U3156);
  nand ginst2918 (P1_R1165_U502, P1_R1165_U34, P1_R1165_U69);
  nand ginst2919 (P1_R1165_U503, P1_R1165_U501, P1_R1165_U502);
  nand ginst2920 (P1_R1165_U504, P1_R1165_U343, P1_R1165_U54);
  nand ginst2921 (P1_R1165_U505, P1_R1165_U308, P1_R1165_U503);
  nand ginst2922 (P1_R1165_U506, P1_R1165_U441, P1_U3157);
  nand ginst2923 (P1_R1165_U507, P1_R1165_U35, P1_R1165_U71);
  nand ginst2924 (P1_R1165_U508, P1_R1165_U506, P1_R1165_U507);
  nand ginst2925 (P1_R1165_U509, P1_R1165_U168, P1_R1165_U344);
  not ginst2926 (P1_R1165_U51, P1_U3159);
  nand ginst2927 (P1_R1165_U510, P1_R1165_U297, P1_R1165_U508);
  nand ginst2928 (P1_R1165_U511, P1_R1165_U483, P1_U3158);
  nand ginst2929 (P1_R1165_U512, P1_R1165_U52, P1_R1165_U85);
  nand ginst2930 (P1_R1165_U513, P1_R1165_U483, P1_U3158);
  nand ginst2931 (P1_R1165_U514, P1_R1165_U52, P1_R1165_U85);
  nand ginst2932 (P1_R1165_U515, P1_R1165_U513, P1_R1165_U514);
  nand ginst2933 (P1_R1165_U516, P1_R1165_U169, P1_R1165_U170);
  nand ginst2934 (P1_R1165_U517, P1_R1165_U293, P1_R1165_U515);
  nand ginst2935 (P1_R1165_U518, P1_R1165_U480, P1_U3159);
  nand ginst2936 (P1_R1165_U519, P1_R1165_U51, P1_R1165_U84);
  not ginst2937 (P1_R1165_U52, P1_U3158);
  nand ginst2938 (P1_R1165_U520, P1_R1165_U480, P1_U3159);
  nand ginst2939 (P1_R1165_U521, P1_R1165_U51, P1_R1165_U84);
  nand ginst2940 (P1_R1165_U522, P1_R1165_U520, P1_R1165_U521);
  nand ginst2941 (P1_R1165_U523, P1_R1165_U171, P1_R1165_U172);
  nand ginst2942 (P1_R1165_U524, P1_R1165_U289, P1_R1165_U522);
  nand ginst2943 (P1_R1165_U525, P1_R1165_U444, P1_U3160);
  nand ginst2944 (P1_R1165_U526, P1_R1165_U36, P1_R1165_U72);
  nand ginst2945 (P1_R1165_U527, P1_R1165_U447, P1_U3161);
  nand ginst2946 (P1_R1165_U528, P1_R1165_U50, P1_R1165_U83);
  nand ginst2947 (P1_R1165_U529, P1_R1165_U527, P1_R1165_U528);
  nand ginst2948 (P1_R1165_U53, P1_R1165_U70, P1_U3155);
  nand ginst2949 (P1_R1165_U530, P1_R1165_U345, P1_R1165_U55);
  nand ginst2950 (P1_R1165_U531, P1_R1165_U317, P1_R1165_U529);
  nand ginst2951 (P1_R1165_U532, P1_R1165_U371, P1_U3180);
  nand ginst2952 (P1_R1165_U533, P1_R1165_U23, P1_R1165_U64);
  nand ginst2953 (P1_R1165_U534, P1_R1165_U371, P1_U3180);
  nand ginst2954 (P1_R1165_U535, P1_R1165_U23, P1_R1165_U64);
  nand ginst2955 (P1_R1165_U536, P1_R1165_U534, P1_R1165_U535);
  nand ginst2956 (P1_R1165_U537, P1_R1165_U173, P1_R1165_U174);
  nand ginst2957 (P1_R1165_U538, P1_R1165_U196, P1_R1165_U536);
  nand ginst2958 (P1_R1165_U539, P1_R1165_U450, P1_U3162);
  nand ginst2959 (P1_R1165_U54, P1_R1165_U192, P1_R1165_U307);
  nand ginst2960 (P1_R1165_U540, P1_R1165_U48, P1_R1165_U82);
  nand ginst2961 (P1_R1165_U541, P1_R1165_U539, P1_R1165_U540);
  nand ginst2962 (P1_R1165_U542, P1_R1165_U175, P1_R1165_U346);
  nand ginst2963 (P1_R1165_U543, P1_R1165_U279, P1_R1165_U541);
  nand ginst2964 (P1_R1165_U544, P1_R1165_U477, P1_U3163);
  nand ginst2965 (P1_R1165_U545, P1_R1165_U47, P1_R1165_U81);
  nand ginst2966 (P1_R1165_U546, P1_R1165_U477, P1_U3163);
  nand ginst2967 (P1_R1165_U547, P1_R1165_U47, P1_R1165_U81);
  nand ginst2968 (P1_R1165_U548, P1_R1165_U546, P1_R1165_U547);
  nand ginst2969 (P1_R1165_U549, P1_R1165_U176, P1_R1165_U177);
  nand ginst2970 (P1_R1165_U55, P1_R1165_U316, P1_R1165_U49);
  nand ginst2971 (P1_R1165_U550, P1_R1165_U275, P1_R1165_U548);
  nand ginst2972 (P1_R1165_U551, P1_R1165_U471, P1_U3164);
  nand ginst2973 (P1_R1165_U552, P1_R1165_U39, P1_R1165_U74);
  nand ginst2974 (P1_R1165_U553, P1_R1165_U474, P1_U3165);
  nand ginst2975 (P1_R1165_U554, P1_R1165_U37, P1_R1165_U73);
  nand ginst2976 (P1_R1165_U555, P1_R1165_U553, P1_R1165_U554);
  nand ginst2977 (P1_R1165_U556, P1_R1165_U347, P1_R1165_U56);
  nand ginst2978 (P1_R1165_U557, P1_R1165_U267, P1_R1165_U555);
  nand ginst2979 (P1_R1165_U558, P1_R1165_U468, P1_U3166);
  nand ginst2980 (P1_R1165_U559, P1_R1165_U46, P1_R1165_U80);
  nand ginst2981 (P1_R1165_U56, P1_R1165_U265, P1_R1165_U266);
  nand ginst2982 (P1_R1165_U560, P1_R1165_U468, P1_U3166);
  nand ginst2983 (P1_R1165_U561, P1_R1165_U46, P1_R1165_U80);
  nand ginst2984 (P1_R1165_U562, P1_R1165_U560, P1_R1165_U561);
  nand ginst2985 (P1_R1165_U563, P1_R1165_U178, P1_R1165_U179);
  nand ginst2986 (P1_R1165_U564, P1_R1165_U263, P1_R1165_U562);
  nand ginst2987 (P1_R1165_U565, P1_R1165_U465, P1_U3167);
  nand ginst2988 (P1_R1165_U566, P1_R1165_U45, P1_R1165_U79);
  nand ginst2989 (P1_R1165_U567, P1_R1165_U465, P1_U3167);
  nand ginst2990 (P1_R1165_U568, P1_R1165_U45, P1_R1165_U79);
  nand ginst2991 (P1_R1165_U569, P1_R1165_U567, P1_R1165_U568);
  nand ginst2992 (P1_R1165_U57, P1_R1165_U332, P1_R1165_U43);
  nand ginst2993 (P1_R1165_U570, P1_R1165_U180, P1_R1165_U181);
  nand ginst2994 (P1_R1165_U571, P1_R1165_U259, P1_R1165_U569);
  nand ginst2995 (P1_R1165_U572, P1_R1165_U456, P1_U3168);
  nand ginst2996 (P1_R1165_U573, P1_R1165_U44, P1_R1165_U77);
  nand ginst2997 (P1_R1165_U574, P1_R1165_U459, P1_U3169);
  nand ginst2998 (P1_R1165_U575, P1_R1165_U41, P1_R1165_U78);
  nand ginst2999 (P1_R1165_U576, P1_R1165_U574, P1_R1165_U575);
  nand ginst3000 (P1_R1165_U577, P1_R1165_U348, P1_R1165_U57);
  nand ginst3001 (P1_R1165_U578, P1_R1165_U333, P1_R1165_U576);
  nand ginst3002 (P1_R1165_U579, P1_R1165_U462, P1_U3170);
  nand ginst3003 (P1_R1165_U58, P1_R1165_U358, P1_R1165_U359);
  nand ginst3004 (P1_R1165_U580, P1_R1165_U42, P1_R1165_U76);
  nand ginst3005 (P1_R1165_U581, P1_R1165_U579, P1_R1165_U580);
  nand ginst3006 (P1_R1165_U582, P1_R1165_U182, P1_R1165_U349);
  nand ginst3007 (P1_R1165_U583, P1_R1165_U249, P1_R1165_U581);
  nand ginst3008 (P1_R1165_U584, P1_R1165_U453, P1_U3171);
  nand ginst3009 (P1_R1165_U585, P1_R1165_U40, P1_R1165_U75);
  nand ginst3010 (P1_R1165_U586, P1_R1165_U453, P1_U3171);
  nand ginst3011 (P1_R1165_U587, P1_R1165_U40, P1_R1165_U75);
  nand ginst3012 (P1_R1165_U588, P1_R1165_U586, P1_R1165_U587);
  nand ginst3013 (P1_R1165_U589, P1_R1165_U183, P1_R1165_U184);
  nand ginst3014 (P1_R1165_U59, P1_R1165_U387, P1_R1165_U388);
  nand ginst3015 (P1_R1165_U590, P1_R1165_U245, P1_R1165_U588);
  nand ginst3016 (P1_R1165_U591, P1_R1165_U15, P1_U3181);
  nand ginst3017 (P1_R1165_U592, P1_R1165_U22, P1_U3211);
  not ginst3018 (P1_R1165_U593, P1_R1165_U129);
  nand ginst3019 (P1_R1165_U594, P1_R1165_U593, P1_R1165_U63);
  nand ginst3020 (P1_R1165_U595, P1_R1165_U129, P1_R1165_U368);
  and ginst3021 (P1_R1165_U6, P1_R1165_U250, P1_R1165_U251);
  nand ginst3022 (P1_R1165_U60, P1_R1165_U384, P1_R1165_U385);
  nand ginst3023 (P1_R1165_U61, P1_R1165_U375, P1_R1165_U376);
  nand ginst3024 (P1_R1165_U62, P1_R1165_U372, P1_R1165_U373);
  nand ginst3025 (P1_R1165_U63, P1_R1165_U366, P1_R1165_U367);
  nand ginst3026 (P1_R1165_U64, P1_R1165_U369, P1_R1165_U370);
  nand ginst3027 (P1_R1165_U65, P1_R1165_U378, P1_R1165_U379);
  nand ginst3028 (P1_R1165_U66, P1_R1165_U381, P1_R1165_U382);
  nand ginst3029 (P1_R1165_U67, P1_R1165_U390, P1_R1165_U391);
  nand ginst3030 (P1_R1165_U68, P1_R1165_U430, P1_R1165_U431);
  nand ginst3031 (P1_R1165_U69, P1_R1165_U433, P1_R1165_U434);
  and ginst3032 (P1_R1165_U7, P1_R1165_U268, P1_R1165_U269);
  nand ginst3033 (P1_R1165_U70, P1_R1165_U436, P1_R1165_U437);
  nand ginst3034 (P1_R1165_U71, P1_R1165_U439, P1_R1165_U440);
  nand ginst3035 (P1_R1165_U72, P1_R1165_U442, P1_R1165_U443);
  nand ginst3036 (P1_R1165_U73, P1_R1165_U472, P1_R1165_U473);
  nand ginst3037 (P1_R1165_U74, P1_R1165_U469, P1_R1165_U470);
  nand ginst3038 (P1_R1165_U75, P1_R1165_U451, P1_R1165_U452);
  nand ginst3039 (P1_R1165_U76, P1_R1165_U460, P1_R1165_U461);
  nand ginst3040 (P1_R1165_U77, P1_R1165_U454, P1_R1165_U455);
  nand ginst3041 (P1_R1165_U78, P1_R1165_U457, P1_R1165_U458);
  nand ginst3042 (P1_R1165_U79, P1_R1165_U463, P1_R1165_U464);
  and ginst3043 (P1_R1165_U8, P1_R1165_U280, P1_R1165_U281);
  nand ginst3044 (P1_R1165_U80, P1_R1165_U466, P1_R1165_U467);
  nand ginst3045 (P1_R1165_U81, P1_R1165_U475, P1_R1165_U476);
  nand ginst3046 (P1_R1165_U82, P1_R1165_U448, P1_R1165_U449);
  nand ginst3047 (P1_R1165_U83, P1_R1165_U445, P1_R1165_U446);
  nand ginst3048 (P1_R1165_U84, P1_R1165_U478, P1_R1165_U479);
  nand ginst3049 (P1_R1165_U85, P1_R1165_U481, P1_R1165_U482);
  nand ginst3050 (P1_R1165_U86, P1_R1165_U487, P1_R1165_U488);
  nand ginst3051 (P1_R1165_U87, P1_R1165_U594, P1_R1165_U595);
  nand ginst3052 (P1_R1165_U88, P1_R1165_U393, P1_R1165_U394);
  nand ginst3053 (P1_R1165_U89, P1_R1165_U400, P1_R1165_U401);
  and ginst3054 (P1_R1165_U9, P1_R1165_U336, P1_R1165_U339);
  nand ginst3055 (P1_R1165_U90, P1_R1165_U407, P1_R1165_U408);
  nand ginst3056 (P1_R1165_U91, P1_R1165_U414, P1_R1165_U415);
  nand ginst3057 (P1_R1165_U92, P1_R1165_U421, P1_R1165_U422);
  nand ginst3058 (P1_R1165_U93, P1_R1165_U428, P1_R1165_U429);
  nand ginst3059 (P1_R1165_U94, P1_R1165_U490, P1_R1165_U491);
  nand ginst3060 (P1_R1165_U95, P1_R1165_U497, P1_R1165_U498);
  nand ginst3061 (P1_R1165_U96, P1_R1165_U504, P1_R1165_U505);
  nand ginst3062 (P1_R1165_U97, P1_R1165_U509, P1_R1165_U510);
  nand ginst3063 (P1_R1165_U98, P1_R1165_U516, P1_R1165_U517);
  nand ginst3064 (P1_R1165_U99, P1_R1165_U523, P1_R1165_U524);
  and ginst3065 (P1_R1171_U10, P1_R1171_U268, P1_R1171_U269);
  nand ginst3066 (P1_R1171_U100, P1_R1171_U390, P1_R1171_U391);
  nand ginst3067 (P1_R1171_U101, P1_R1171_U395, P1_R1171_U396);
  nand ginst3068 (P1_R1171_U102, P1_R1171_U404, P1_R1171_U405);
  nand ginst3069 (P1_R1171_U103, P1_R1171_U411, P1_R1171_U412);
  nand ginst3070 (P1_R1171_U104, P1_R1171_U418, P1_R1171_U419);
  nand ginst3071 (P1_R1171_U105, P1_R1171_U425, P1_R1171_U426);
  nand ginst3072 (P1_R1171_U106, P1_R1171_U430, P1_R1171_U431);
  nand ginst3073 (P1_R1171_U107, P1_R1171_U437, P1_R1171_U438);
  nand ginst3074 (P1_R1171_U108, P1_R1171_U444, P1_R1171_U445);
  nand ginst3075 (P1_R1171_U109, P1_R1171_U458, P1_R1171_U459);
  and ginst3076 (P1_R1171_U11, P1_R1171_U345, P1_R1171_U348);
  nand ginst3077 (P1_R1171_U110, P1_R1171_U463, P1_R1171_U464);
  nand ginst3078 (P1_R1171_U111, P1_R1171_U470, P1_R1171_U471);
  nand ginst3079 (P1_R1171_U112, P1_R1171_U477, P1_R1171_U478);
  nand ginst3080 (P1_R1171_U113, P1_R1171_U484, P1_R1171_U485);
  nand ginst3081 (P1_R1171_U114, P1_R1171_U491, P1_R1171_U492);
  nand ginst3082 (P1_R1171_U115, P1_R1171_U496, P1_R1171_U497);
  and ginst3083 (P1_R1171_U116, P1_U3068, P1_U3464);
  and ginst3084 (P1_R1171_U117, P1_R1171_U184, P1_R1171_U186);
  and ginst3085 (P1_R1171_U118, P1_R1171_U189, P1_R1171_U191);
  and ginst3086 (P1_R1171_U119, P1_R1171_U197, P1_R1171_U198);
  and ginst3087 (P1_R1171_U12, P1_R1171_U338, P1_R1171_U341);
  and ginst3088 (P1_R1171_U120, P1_R1171_U23, P1_R1171_U378, P1_R1171_U379);
  and ginst3089 (P1_R1171_U121, P1_R1171_U209, P1_R1171_U6);
  and ginst3090 (P1_R1171_U122, P1_R1171_U215, P1_R1171_U217);
  and ginst3091 (P1_R1171_U123, P1_R1171_U35, P1_R1171_U385, P1_R1171_U386);
  and ginst3092 (P1_R1171_U124, P1_R1171_U223, P1_R1171_U4);
  and ginst3093 (P1_R1171_U125, P1_R1171_U178, P1_R1171_U231);
  and ginst3094 (P1_R1171_U126, P1_R1171_U201, P1_R1171_U7);
  and ginst3095 (P1_R1171_U127, P1_R1171_U168, P1_R1171_U236);
  and ginst3096 (P1_R1171_U128, P1_R1171_U169, P1_R1171_U245);
  and ginst3097 (P1_R1171_U129, P1_R1171_U264, P1_R1171_U265);
  and ginst3098 (P1_R1171_U13, P1_R1171_U329, P1_R1171_U332);
  and ginst3099 (P1_R1171_U130, P1_R1171_U10, P1_R1171_U279);
  and ginst3100 (P1_R1171_U131, P1_R1171_U277, P1_R1171_U282);
  and ginst3101 (P1_R1171_U132, P1_R1171_U295, P1_R1171_U298);
  and ginst3102 (P1_R1171_U133, P1_R1171_U299, P1_R1171_U365);
  and ginst3103 (P1_R1171_U134, P1_R1171_U156, P1_R1171_U275);
  and ginst3104 (P1_R1171_U135, P1_R1171_U465, P1_R1171_U466, P1_R1171_U60);
  and ginst3105 (P1_R1171_U136, P1_R1171_U169, P1_R1171_U486, P1_R1171_U487);
  and ginst3106 (P1_R1171_U137, P1_R1171_U340, P1_R1171_U8);
  and ginst3107 (P1_R1171_U138, P1_R1171_U168, P1_R1171_U498, P1_R1171_U499);
  and ginst3108 (P1_R1171_U139, P1_R1171_U347, P1_R1171_U7);
  and ginst3109 (P1_R1171_U14, P1_R1171_U320, P1_R1171_U323);
  nand ginst3110 (P1_R1171_U140, P1_R1171_U119, P1_R1171_U199);
  nand ginst3111 (P1_R1171_U141, P1_R1171_U214, P1_R1171_U226);
  not ginst3112 (P1_R1171_U142, P1_U3055);
  not ginst3113 (P1_R1171_U143, P1_U4028);
  and ginst3114 (P1_R1171_U144, P1_R1171_U399, P1_R1171_U400);
  nand ginst3115 (P1_R1171_U145, P1_R1171_U166, P1_R1171_U301, P1_R1171_U361);
  and ginst3116 (P1_R1171_U146, P1_R1171_U406, P1_R1171_U407);
  nand ginst3117 (P1_R1171_U147, P1_R1171_U133, P1_R1171_U366, P1_R1171_U367);
  and ginst3118 (P1_R1171_U148, P1_R1171_U413, P1_R1171_U414);
  nand ginst3119 (P1_R1171_U149, P1_R1171_U296, P1_R1171_U362, P1_R1171_U87);
  and ginst3120 (P1_R1171_U15, P1_R1171_U315, P1_R1171_U317);
  and ginst3121 (P1_R1171_U150, P1_R1171_U420, P1_R1171_U421);
  nand ginst3122 (P1_R1171_U151, P1_R1171_U289, P1_R1171_U290);
  and ginst3123 (P1_R1171_U152, P1_R1171_U432, P1_R1171_U433);
  nand ginst3124 (P1_R1171_U153, P1_R1171_U285, P1_R1171_U286);
  and ginst3125 (P1_R1171_U154, P1_R1171_U439, P1_R1171_U440);
  nand ginst3126 (P1_R1171_U155, P1_R1171_U131, P1_R1171_U281);
  and ginst3127 (P1_R1171_U156, P1_R1171_U446, P1_R1171_U447);
  and ginst3128 (P1_R1171_U157, P1_R1171_U451, P1_R1171_U452);
  nand ginst3129 (P1_R1171_U158, P1_R1171_U324, P1_R1171_U44);
  nand ginst3130 (P1_R1171_U159, P1_R1171_U129, P1_R1171_U266);
  and ginst3131 (P1_R1171_U16, P1_R1171_U307, P1_R1171_U310);
  and ginst3132 (P1_R1171_U160, P1_R1171_U472, P1_R1171_U473);
  nand ginst3133 (P1_R1171_U161, P1_R1171_U253, P1_R1171_U254);
  and ginst3134 (P1_R1171_U162, P1_R1171_U479, P1_R1171_U480);
  nand ginst3135 (P1_R1171_U163, P1_R1171_U249, P1_R1171_U250);
  nand ginst3136 (P1_R1171_U164, P1_R1171_U239, P1_R1171_U240);
  nand ginst3137 (P1_R1171_U165, P1_R1171_U363, P1_R1171_U364);
  nand ginst3138 (P1_R1171_U166, P1_R1171_U147, P1_U3054);
  not ginst3139 (P1_R1171_U167, P1_R1171_U35);
  nand ginst3140 (P1_R1171_U168, P1_U3083, P1_U3485);
  nand ginst3141 (P1_R1171_U169, P1_U3072, P1_U3494);
  and ginst3142 (P1_R1171_U17, P1_R1171_U229, P1_R1171_U232);
  nand ginst3143 (P1_R1171_U170, P1_U3058, P1_U4020);
  not ginst3144 (P1_R1171_U171, P1_R1171_U69);
  not ginst3145 (P1_R1171_U172, P1_R1171_U78);
  nand ginst3146 (P1_R1171_U173, P1_U3065, P1_U4021);
  not ginst3147 (P1_R1171_U174, P1_R1171_U62);
  or ginst3148 (P1_R1171_U175, P1_U3067, P1_U3473);
  or ginst3149 (P1_R1171_U176, P1_U3060, P1_U3470);
  or ginst3150 (P1_R1171_U177, P1_U3064, P1_U3467);
  or ginst3151 (P1_R1171_U178, P1_U3068, P1_U3464);
  not ginst3152 (P1_R1171_U179, P1_R1171_U32);
  and ginst3153 (P1_R1171_U18, P1_R1171_U221, P1_R1171_U224);
  or ginst3154 (P1_R1171_U180, P1_U3078, P1_U3461);
  not ginst3155 (P1_R1171_U181, P1_R1171_U43);
  not ginst3156 (P1_R1171_U182, P1_R1171_U44);
  nand ginst3157 (P1_R1171_U183, P1_R1171_U43, P1_R1171_U44);
  nand ginst3158 (P1_R1171_U184, P1_R1171_U116, P1_R1171_U177);
  nand ginst3159 (P1_R1171_U185, P1_R1171_U183, P1_R1171_U5);
  nand ginst3160 (P1_R1171_U186, P1_U3064, P1_U3467);
  nand ginst3161 (P1_R1171_U187, P1_R1171_U117, P1_R1171_U185);
  nand ginst3162 (P1_R1171_U188, P1_R1171_U35, P1_R1171_U36);
  nand ginst3163 (P1_R1171_U189, P1_R1171_U188, P1_U3067);
  and ginst3164 (P1_R1171_U19, P1_R1171_U207, P1_R1171_U210);
  nand ginst3165 (P1_R1171_U190, P1_R1171_U187, P1_R1171_U4);
  nand ginst3166 (P1_R1171_U191, P1_R1171_U167, P1_U3473);
  not ginst3167 (P1_R1171_U192, P1_R1171_U42);
  or ginst3168 (P1_R1171_U193, P1_U3070, P1_U3479);
  or ginst3169 (P1_R1171_U194, P1_U3071, P1_U3476);
  not ginst3170 (P1_R1171_U195, P1_R1171_U23);
  nand ginst3171 (P1_R1171_U196, P1_R1171_U23, P1_R1171_U24);
  nand ginst3172 (P1_R1171_U197, P1_R1171_U196, P1_U3070);
  nand ginst3173 (P1_R1171_U198, P1_R1171_U195, P1_U3479);
  nand ginst3174 (P1_R1171_U199, P1_R1171_U42, P1_R1171_U6);
  not ginst3175 (P1_R1171_U20, P1_U3476);
  not ginst3176 (P1_R1171_U200, P1_R1171_U140);
  or ginst3177 (P1_R1171_U201, P1_U3084, P1_U3482);
  nand ginst3178 (P1_R1171_U202, P1_R1171_U140, P1_R1171_U201);
  not ginst3179 (P1_R1171_U203, P1_R1171_U41);
  or ginst3180 (P1_R1171_U204, P1_U3083, P1_U3485);
  or ginst3181 (P1_R1171_U205, P1_U3071, P1_U3476);
  nand ginst3182 (P1_R1171_U206, P1_R1171_U205, P1_R1171_U42);
  nand ginst3183 (P1_R1171_U207, P1_R1171_U120, P1_R1171_U206);
  nand ginst3184 (P1_R1171_U208, P1_R1171_U192, P1_R1171_U23);
  nand ginst3185 (P1_R1171_U209, P1_U3070, P1_U3479);
  not ginst3186 (P1_R1171_U21, P1_U3071);
  nand ginst3187 (P1_R1171_U210, P1_R1171_U121, P1_R1171_U208);
  or ginst3188 (P1_R1171_U211, P1_U3071, P1_U3476);
  nand ginst3189 (P1_R1171_U212, P1_R1171_U178, P1_R1171_U182);
  nand ginst3190 (P1_R1171_U213, P1_U3068, P1_U3464);
  not ginst3191 (P1_R1171_U214, P1_R1171_U46);
  nand ginst3192 (P1_R1171_U215, P1_R1171_U181, P1_R1171_U5);
  nand ginst3193 (P1_R1171_U216, P1_R1171_U177, P1_R1171_U46);
  nand ginst3194 (P1_R1171_U217, P1_U3064, P1_U3467);
  not ginst3195 (P1_R1171_U218, P1_R1171_U45);
  or ginst3196 (P1_R1171_U219, P1_U3060, P1_U3470);
  not ginst3197 (P1_R1171_U22, P1_U3070);
  nand ginst3198 (P1_R1171_U220, P1_R1171_U219, P1_R1171_U45);
  nand ginst3199 (P1_R1171_U221, P1_R1171_U123, P1_R1171_U220);
  nand ginst3200 (P1_R1171_U222, P1_R1171_U218, P1_R1171_U35);
  nand ginst3201 (P1_R1171_U223, P1_U3067, P1_U3473);
  nand ginst3202 (P1_R1171_U224, P1_R1171_U124, P1_R1171_U222);
  or ginst3203 (P1_R1171_U225, P1_U3060, P1_U3470);
  nand ginst3204 (P1_R1171_U226, P1_R1171_U178, P1_R1171_U181);
  not ginst3205 (P1_R1171_U227, P1_R1171_U141);
  nand ginst3206 (P1_R1171_U228, P1_U3064, P1_U3467);
  nand ginst3207 (P1_R1171_U229, P1_R1171_U397, P1_R1171_U398, P1_R1171_U43, P1_R1171_U44);
  nand ginst3208 (P1_R1171_U23, P1_U3071, P1_U3476);
  nand ginst3209 (P1_R1171_U230, P1_R1171_U43, P1_R1171_U44);
  nand ginst3210 (P1_R1171_U231, P1_U3068, P1_U3464);
  nand ginst3211 (P1_R1171_U232, P1_R1171_U125, P1_R1171_U230);
  or ginst3212 (P1_R1171_U233, P1_U3083, P1_U3485);
  or ginst3213 (P1_R1171_U234, P1_U3062, P1_U3488);
  nand ginst3214 (P1_R1171_U235, P1_R1171_U174, P1_R1171_U7);
  nand ginst3215 (P1_R1171_U236, P1_U3062, P1_U3488);
  nand ginst3216 (P1_R1171_U237, P1_R1171_U127, P1_R1171_U235);
  or ginst3217 (P1_R1171_U238, P1_U3062, P1_U3488);
  nand ginst3218 (P1_R1171_U239, P1_R1171_U126, P1_R1171_U140);
  not ginst3219 (P1_R1171_U24, P1_U3479);
  nand ginst3220 (P1_R1171_U240, P1_R1171_U237, P1_R1171_U238);
  not ginst3221 (P1_R1171_U241, P1_R1171_U164);
  or ginst3222 (P1_R1171_U242, P1_U3080, P1_U3497);
  or ginst3223 (P1_R1171_U243, P1_U3072, P1_U3494);
  nand ginst3224 (P1_R1171_U244, P1_R1171_U171, P1_R1171_U8);
  nand ginst3225 (P1_R1171_U245, P1_U3080, P1_U3497);
  nand ginst3226 (P1_R1171_U246, P1_R1171_U128, P1_R1171_U244);
  or ginst3227 (P1_R1171_U247, P1_U3063, P1_U3491);
  or ginst3228 (P1_R1171_U248, P1_U3080, P1_U3497);
  nand ginst3229 (P1_R1171_U249, P1_R1171_U164, P1_R1171_U247, P1_R1171_U8);
  not ginst3230 (P1_R1171_U25, P1_U3470);
  nand ginst3231 (P1_R1171_U250, P1_R1171_U246, P1_R1171_U248);
  not ginst3232 (P1_R1171_U251, P1_R1171_U163);
  or ginst3233 (P1_R1171_U252, P1_U3079, P1_U3500);
  nand ginst3234 (P1_R1171_U253, P1_R1171_U163, P1_R1171_U252);
  nand ginst3235 (P1_R1171_U254, P1_U3079, P1_U3500);
  not ginst3236 (P1_R1171_U255, P1_R1171_U161);
  or ginst3237 (P1_R1171_U256, P1_U3074, P1_U3503);
  nand ginst3238 (P1_R1171_U257, P1_R1171_U161, P1_R1171_U256);
  nand ginst3239 (P1_R1171_U258, P1_U3074, P1_U3503);
  not ginst3240 (P1_R1171_U259, P1_R1171_U93);
  not ginst3241 (P1_R1171_U26, P1_U3060);
  or ginst3242 (P1_R1171_U260, P1_U3069, P1_U3509);
  or ginst3243 (P1_R1171_U261, P1_U3073, P1_U3506);
  not ginst3244 (P1_R1171_U262, P1_R1171_U60);
  nand ginst3245 (P1_R1171_U263, P1_R1171_U60, P1_R1171_U61);
  nand ginst3246 (P1_R1171_U264, P1_R1171_U263, P1_U3069);
  nand ginst3247 (P1_R1171_U265, P1_R1171_U262, P1_U3509);
  nand ginst3248 (P1_R1171_U266, P1_R1171_U9, P1_R1171_U93);
  not ginst3249 (P1_R1171_U267, P1_R1171_U159);
  or ginst3250 (P1_R1171_U268, P1_U3076, P1_U4025);
  or ginst3251 (P1_R1171_U269, P1_U3081, P1_U3514);
  not ginst3252 (P1_R1171_U27, P1_U3067);
  or ginst3253 (P1_R1171_U270, P1_U3075, P1_U4024);
  not ginst3254 (P1_R1171_U271, P1_R1171_U81);
  nand ginst3255 (P1_R1171_U272, P1_R1171_U271, P1_U4025);
  nand ginst3256 (P1_R1171_U273, P1_R1171_U272, P1_R1171_U91);
  nand ginst3257 (P1_R1171_U274, P1_R1171_U81, P1_R1171_U82);
  nand ginst3258 (P1_R1171_U275, P1_R1171_U273, P1_R1171_U274);
  nand ginst3259 (P1_R1171_U276, P1_R1171_U10, P1_R1171_U172);
  nand ginst3260 (P1_R1171_U277, P1_U3075, P1_U4024);
  nand ginst3261 (P1_R1171_U278, P1_R1171_U275, P1_R1171_U276);
  or ginst3262 (P1_R1171_U279, P1_U3082, P1_U3512);
  not ginst3263 (P1_R1171_U28, P1_U3464);
  or ginst3264 (P1_R1171_U280, P1_U3075, P1_U4024);
  nand ginst3265 (P1_R1171_U281, P1_R1171_U130, P1_R1171_U159, P1_R1171_U270);
  nand ginst3266 (P1_R1171_U282, P1_R1171_U278, P1_R1171_U280);
  not ginst3267 (P1_R1171_U283, P1_R1171_U155);
  or ginst3268 (P1_R1171_U284, P1_U3061, P1_U4023);
  nand ginst3269 (P1_R1171_U285, P1_R1171_U155, P1_R1171_U284);
  nand ginst3270 (P1_R1171_U286, P1_U3061, P1_U4023);
  not ginst3271 (P1_R1171_U287, P1_R1171_U153);
  or ginst3272 (P1_R1171_U288, P1_U3066, P1_U4022);
  nand ginst3273 (P1_R1171_U289, P1_R1171_U153, P1_R1171_U288);
  not ginst3274 (P1_R1171_U29, P1_U3068);
  nand ginst3275 (P1_R1171_U290, P1_U3066, P1_U4022);
  not ginst3276 (P1_R1171_U291, P1_R1171_U151);
  or ginst3277 (P1_R1171_U292, P1_U3058, P1_U4020);
  nand ginst3278 (P1_R1171_U293, P1_R1171_U170, P1_R1171_U173);
  not ginst3279 (P1_R1171_U294, P1_R1171_U87);
  or ginst3280 (P1_R1171_U295, P1_U3065, P1_U4021);
  nand ginst3281 (P1_R1171_U296, P1_R1171_U151, P1_R1171_U165, P1_R1171_U295);
  not ginst3282 (P1_R1171_U297, P1_R1171_U149);
  or ginst3283 (P1_R1171_U298, P1_U3053, P1_U4018);
  nand ginst3284 (P1_R1171_U299, P1_U3053, P1_U4018);
  not ginst3285 (P1_R1171_U30, P1_U3456);
  not ginst3286 (P1_R1171_U300, P1_R1171_U147);
  nand ginst3287 (P1_R1171_U301, P1_R1171_U147, P1_U4017);
  not ginst3288 (P1_R1171_U302, P1_R1171_U145);
  nand ginst3289 (P1_R1171_U303, P1_R1171_U151, P1_R1171_U295);
  not ginst3290 (P1_R1171_U304, P1_R1171_U90);
  or ginst3291 (P1_R1171_U305, P1_U3058, P1_U4020);
  nand ginst3292 (P1_R1171_U306, P1_R1171_U305, P1_R1171_U90);
  nand ginst3293 (P1_R1171_U307, P1_R1171_U150, P1_R1171_U170, P1_R1171_U306);
  nand ginst3294 (P1_R1171_U308, P1_R1171_U170, P1_R1171_U304);
  nand ginst3295 (P1_R1171_U309, P1_U3057, P1_U4019);
  not ginst3296 (P1_R1171_U31, P1_U3077);
  nand ginst3297 (P1_R1171_U310, P1_R1171_U165, P1_R1171_U308, P1_R1171_U309);
  or ginst3298 (P1_R1171_U311, P1_U3058, P1_U4020);
  nand ginst3299 (P1_R1171_U312, P1_R1171_U159, P1_R1171_U279);
  not ginst3300 (P1_R1171_U313, P1_R1171_U92);
  nand ginst3301 (P1_R1171_U314, P1_R1171_U10, P1_R1171_U92);
  nand ginst3302 (P1_R1171_U315, P1_R1171_U134, P1_R1171_U314);
  nand ginst3303 (P1_R1171_U316, P1_R1171_U275, P1_R1171_U314);
  nand ginst3304 (P1_R1171_U317, P1_R1171_U316, P1_R1171_U450);
  or ginst3305 (P1_R1171_U318, P1_U3081, P1_U3514);
  nand ginst3306 (P1_R1171_U319, P1_R1171_U318, P1_R1171_U92);
  nand ginst3307 (P1_R1171_U32, P1_U3077, P1_U3456);
  nand ginst3308 (P1_R1171_U320, P1_R1171_U157, P1_R1171_U319, P1_R1171_U81);
  nand ginst3309 (P1_R1171_U321, P1_R1171_U313, P1_R1171_U81);
  nand ginst3310 (P1_R1171_U322, P1_U3076, P1_U4025);
  nand ginst3311 (P1_R1171_U323, P1_R1171_U10, P1_R1171_U321, P1_R1171_U322);
  or ginst3312 (P1_R1171_U324, P1_U3078, P1_U3461);
  not ginst3313 (P1_R1171_U325, P1_R1171_U158);
  or ginst3314 (P1_R1171_U326, P1_U3081, P1_U3514);
  or ginst3315 (P1_R1171_U327, P1_U3073, P1_U3506);
  nand ginst3316 (P1_R1171_U328, P1_R1171_U327, P1_R1171_U93);
  nand ginst3317 (P1_R1171_U329, P1_R1171_U135, P1_R1171_U328);
  not ginst3318 (P1_R1171_U33, P1_U3467);
  nand ginst3319 (P1_R1171_U330, P1_R1171_U259, P1_R1171_U60);
  nand ginst3320 (P1_R1171_U331, P1_U3069, P1_U3509);
  nand ginst3321 (P1_R1171_U332, P1_R1171_U330, P1_R1171_U331, P1_R1171_U9);
  or ginst3322 (P1_R1171_U333, P1_U3073, P1_U3506);
  nand ginst3323 (P1_R1171_U334, P1_R1171_U164, P1_R1171_U247);
  not ginst3324 (P1_R1171_U335, P1_R1171_U94);
  or ginst3325 (P1_R1171_U336, P1_U3072, P1_U3494);
  nand ginst3326 (P1_R1171_U337, P1_R1171_U336, P1_R1171_U94);
  nand ginst3327 (P1_R1171_U338, P1_R1171_U136, P1_R1171_U337);
  nand ginst3328 (P1_R1171_U339, P1_R1171_U169, P1_R1171_U335);
  not ginst3329 (P1_R1171_U34, P1_U3064);
  nand ginst3330 (P1_R1171_U340, P1_U3080, P1_U3497);
  nand ginst3331 (P1_R1171_U341, P1_R1171_U137, P1_R1171_U339);
  or ginst3332 (P1_R1171_U342, P1_U3072, P1_U3494);
  or ginst3333 (P1_R1171_U343, P1_U3083, P1_U3485);
  nand ginst3334 (P1_R1171_U344, P1_R1171_U343, P1_R1171_U41);
  nand ginst3335 (P1_R1171_U345, P1_R1171_U138, P1_R1171_U344);
  nand ginst3336 (P1_R1171_U346, P1_R1171_U168, P1_R1171_U203);
  nand ginst3337 (P1_R1171_U347, P1_U3062, P1_U3488);
  nand ginst3338 (P1_R1171_U348, P1_R1171_U139, P1_R1171_U346);
  nand ginst3339 (P1_R1171_U349, P1_R1171_U168, P1_R1171_U204);
  nand ginst3340 (P1_R1171_U35, P1_U3060, P1_U3470);
  nand ginst3341 (P1_R1171_U350, P1_R1171_U201, P1_R1171_U62);
  nand ginst3342 (P1_R1171_U351, P1_R1171_U211, P1_R1171_U23);
  nand ginst3343 (P1_R1171_U352, P1_R1171_U225, P1_R1171_U35);
  nand ginst3344 (P1_R1171_U353, P1_R1171_U177, P1_R1171_U228);
  nand ginst3345 (P1_R1171_U354, P1_R1171_U170, P1_R1171_U311);
  nand ginst3346 (P1_R1171_U355, P1_R1171_U173, P1_R1171_U295);
  nand ginst3347 (P1_R1171_U356, P1_R1171_U326, P1_R1171_U81);
  nand ginst3348 (P1_R1171_U357, P1_R1171_U279, P1_R1171_U78);
  nand ginst3349 (P1_R1171_U358, P1_R1171_U333, P1_R1171_U60);
  nand ginst3350 (P1_R1171_U359, P1_R1171_U169, P1_R1171_U342);
  not ginst3351 (P1_R1171_U36, P1_U3473);
  nand ginst3352 (P1_R1171_U360, P1_R1171_U247, P1_R1171_U69);
  nand ginst3353 (P1_R1171_U361, P1_U3054, P1_U4017);
  nand ginst3354 (P1_R1171_U362, P1_R1171_U165, P1_R1171_U293);
  nand ginst3355 (P1_R1171_U363, P1_R1171_U292, P1_U3057);
  nand ginst3356 (P1_R1171_U364, P1_R1171_U292, P1_U4019);
  nand ginst3357 (P1_R1171_U365, P1_R1171_U165, P1_R1171_U293, P1_R1171_U298);
  nand ginst3358 (P1_R1171_U366, P1_R1171_U132, P1_R1171_U151, P1_R1171_U165);
  nand ginst3359 (P1_R1171_U367, P1_R1171_U294, P1_R1171_U298);
  nand ginst3360 (P1_R1171_U368, P1_R1171_U40, P1_U3083);
  nand ginst3361 (P1_R1171_U369, P1_R1171_U39, P1_U3485);
  not ginst3362 (P1_R1171_U37, P1_U3482);
  nand ginst3363 (P1_R1171_U370, P1_R1171_U368, P1_R1171_U369);
  nand ginst3364 (P1_R1171_U371, P1_R1171_U349, P1_R1171_U41);
  nand ginst3365 (P1_R1171_U372, P1_R1171_U203, P1_R1171_U370);
  nand ginst3366 (P1_R1171_U373, P1_R1171_U37, P1_U3084);
  nand ginst3367 (P1_R1171_U374, P1_R1171_U38, P1_U3482);
  nand ginst3368 (P1_R1171_U375, P1_R1171_U373, P1_R1171_U374);
  nand ginst3369 (P1_R1171_U376, P1_R1171_U140, P1_R1171_U350);
  nand ginst3370 (P1_R1171_U377, P1_R1171_U200, P1_R1171_U375);
  nand ginst3371 (P1_R1171_U378, P1_R1171_U24, P1_U3070);
  nand ginst3372 (P1_R1171_U379, P1_R1171_U22, P1_U3479);
  not ginst3373 (P1_R1171_U38, P1_U3084);
  nand ginst3374 (P1_R1171_U380, P1_R1171_U20, P1_U3071);
  nand ginst3375 (P1_R1171_U381, P1_R1171_U21, P1_U3476);
  nand ginst3376 (P1_R1171_U382, P1_R1171_U380, P1_R1171_U381);
  nand ginst3377 (P1_R1171_U383, P1_R1171_U351, P1_R1171_U42);
  nand ginst3378 (P1_R1171_U384, P1_R1171_U192, P1_R1171_U382);
  nand ginst3379 (P1_R1171_U385, P1_R1171_U36, P1_U3067);
  nand ginst3380 (P1_R1171_U386, P1_R1171_U27, P1_U3473);
  nand ginst3381 (P1_R1171_U387, P1_R1171_U25, P1_U3060);
  nand ginst3382 (P1_R1171_U388, P1_R1171_U26, P1_U3470);
  nand ginst3383 (P1_R1171_U389, P1_R1171_U387, P1_R1171_U388);
  not ginst3384 (P1_R1171_U39, P1_U3083);
  nand ginst3385 (P1_R1171_U390, P1_R1171_U352, P1_R1171_U45);
  nand ginst3386 (P1_R1171_U391, P1_R1171_U218, P1_R1171_U389);
  nand ginst3387 (P1_R1171_U392, P1_R1171_U33, P1_U3064);
  nand ginst3388 (P1_R1171_U393, P1_R1171_U34, P1_U3467);
  nand ginst3389 (P1_R1171_U394, P1_R1171_U392, P1_R1171_U393);
  nand ginst3390 (P1_R1171_U395, P1_R1171_U141, P1_R1171_U353);
  nand ginst3391 (P1_R1171_U396, P1_R1171_U227, P1_R1171_U394);
  nand ginst3392 (P1_R1171_U397, P1_R1171_U28, P1_U3068);
  nand ginst3393 (P1_R1171_U398, P1_R1171_U29, P1_U3464);
  nand ginst3394 (P1_R1171_U399, P1_R1171_U143, P1_U3055);
  and ginst3395 (P1_R1171_U4, P1_R1171_U175, P1_R1171_U176);
  not ginst3396 (P1_R1171_U40, P1_U3485);
  nand ginst3397 (P1_R1171_U400, P1_R1171_U142, P1_U4028);
  nand ginst3398 (P1_R1171_U401, P1_R1171_U143, P1_U3055);
  nand ginst3399 (P1_R1171_U402, P1_R1171_U142, P1_U4028);
  nand ginst3400 (P1_R1171_U403, P1_R1171_U401, P1_R1171_U402);
  nand ginst3401 (P1_R1171_U404, P1_R1171_U144, P1_R1171_U145);
  nand ginst3402 (P1_R1171_U405, P1_R1171_U302, P1_R1171_U403);
  nand ginst3403 (P1_R1171_U406, P1_R1171_U89, P1_U3054);
  nand ginst3404 (P1_R1171_U407, P1_R1171_U88, P1_U4017);
  nand ginst3405 (P1_R1171_U408, P1_R1171_U89, P1_U3054);
  nand ginst3406 (P1_R1171_U409, P1_R1171_U88, P1_U4017);
  nand ginst3407 (P1_R1171_U41, P1_R1171_U202, P1_R1171_U62);
  nand ginst3408 (P1_R1171_U410, P1_R1171_U408, P1_R1171_U409);
  nand ginst3409 (P1_R1171_U411, P1_R1171_U146, P1_R1171_U147);
  nand ginst3410 (P1_R1171_U412, P1_R1171_U300, P1_R1171_U410);
  nand ginst3411 (P1_R1171_U413, P1_R1171_U47, P1_U3053);
  nand ginst3412 (P1_R1171_U414, P1_R1171_U48, P1_U4018);
  nand ginst3413 (P1_R1171_U415, P1_R1171_U47, P1_U3053);
  nand ginst3414 (P1_R1171_U416, P1_R1171_U48, P1_U4018);
  nand ginst3415 (P1_R1171_U417, P1_R1171_U415, P1_R1171_U416);
  nand ginst3416 (P1_R1171_U418, P1_R1171_U148, P1_R1171_U149);
  nand ginst3417 (P1_R1171_U419, P1_R1171_U297, P1_R1171_U417);
  nand ginst3418 (P1_R1171_U42, P1_R1171_U118, P1_R1171_U190);
  nand ginst3419 (P1_R1171_U420, P1_R1171_U50, P1_U3057);
  nand ginst3420 (P1_R1171_U421, P1_R1171_U49, P1_U4019);
  nand ginst3421 (P1_R1171_U422, P1_R1171_U51, P1_U3058);
  nand ginst3422 (P1_R1171_U423, P1_R1171_U52, P1_U4020);
  nand ginst3423 (P1_R1171_U424, P1_R1171_U422, P1_R1171_U423);
  nand ginst3424 (P1_R1171_U425, P1_R1171_U354, P1_R1171_U90);
  nand ginst3425 (P1_R1171_U426, P1_R1171_U304, P1_R1171_U424);
  nand ginst3426 (P1_R1171_U427, P1_R1171_U53, P1_U3065);
  nand ginst3427 (P1_R1171_U428, P1_R1171_U54, P1_U4021);
  nand ginst3428 (P1_R1171_U429, P1_R1171_U427, P1_R1171_U428);
  nand ginst3429 (P1_R1171_U43, P1_R1171_U179, P1_R1171_U180);
  nand ginst3430 (P1_R1171_U430, P1_R1171_U151, P1_R1171_U355);
  nand ginst3431 (P1_R1171_U431, P1_R1171_U291, P1_R1171_U429);
  nand ginst3432 (P1_R1171_U432, P1_R1171_U85, P1_U3066);
  nand ginst3433 (P1_R1171_U433, P1_R1171_U86, P1_U4022);
  nand ginst3434 (P1_R1171_U434, P1_R1171_U85, P1_U3066);
  nand ginst3435 (P1_R1171_U435, P1_R1171_U86, P1_U4022);
  nand ginst3436 (P1_R1171_U436, P1_R1171_U434, P1_R1171_U435);
  nand ginst3437 (P1_R1171_U437, P1_R1171_U152, P1_R1171_U153);
  nand ginst3438 (P1_R1171_U438, P1_R1171_U287, P1_R1171_U436);
  nand ginst3439 (P1_R1171_U439, P1_R1171_U83, P1_U3061);
  nand ginst3440 (P1_R1171_U44, P1_U3078, P1_U3461);
  nand ginst3441 (P1_R1171_U440, P1_R1171_U84, P1_U4023);
  nand ginst3442 (P1_R1171_U441, P1_R1171_U83, P1_U3061);
  nand ginst3443 (P1_R1171_U442, P1_R1171_U84, P1_U4023);
  nand ginst3444 (P1_R1171_U443, P1_R1171_U441, P1_R1171_U442);
  nand ginst3445 (P1_R1171_U444, P1_R1171_U154, P1_R1171_U155);
  nand ginst3446 (P1_R1171_U445, P1_R1171_U283, P1_R1171_U443);
  nand ginst3447 (P1_R1171_U446, P1_R1171_U55, P1_U3075);
  nand ginst3448 (P1_R1171_U447, P1_R1171_U56, P1_U4024);
  nand ginst3449 (P1_R1171_U448, P1_R1171_U55, P1_U3075);
  nand ginst3450 (P1_R1171_U449, P1_R1171_U56, P1_U4024);
  nand ginst3451 (P1_R1171_U45, P1_R1171_U122, P1_R1171_U216);
  nand ginst3452 (P1_R1171_U450, P1_R1171_U448, P1_R1171_U449);
  nand ginst3453 (P1_R1171_U451, P1_R1171_U82, P1_U3076);
  nand ginst3454 (P1_R1171_U452, P1_R1171_U91, P1_U4025);
  nand ginst3455 (P1_R1171_U453, P1_R1171_U158, P1_R1171_U179);
  nand ginst3456 (P1_R1171_U454, P1_R1171_U32, P1_R1171_U325);
  nand ginst3457 (P1_R1171_U455, P1_R1171_U79, P1_U3081);
  nand ginst3458 (P1_R1171_U456, P1_R1171_U80, P1_U3514);
  nand ginst3459 (P1_R1171_U457, P1_R1171_U455, P1_R1171_U456);
  nand ginst3460 (P1_R1171_U458, P1_R1171_U356, P1_R1171_U92);
  nand ginst3461 (P1_R1171_U459, P1_R1171_U313, P1_R1171_U457);
  nand ginst3462 (P1_R1171_U46, P1_R1171_U212, P1_R1171_U213);
  nand ginst3463 (P1_R1171_U460, P1_R1171_U76, P1_U3082);
  nand ginst3464 (P1_R1171_U461, P1_R1171_U77, P1_U3512);
  nand ginst3465 (P1_R1171_U462, P1_R1171_U460, P1_R1171_U461);
  nand ginst3466 (P1_R1171_U463, P1_R1171_U159, P1_R1171_U357);
  nand ginst3467 (P1_R1171_U464, P1_R1171_U267, P1_R1171_U462);
  nand ginst3468 (P1_R1171_U465, P1_R1171_U61, P1_U3069);
  nand ginst3469 (P1_R1171_U466, P1_R1171_U59, P1_U3509);
  nand ginst3470 (P1_R1171_U467, P1_R1171_U57, P1_U3073);
  nand ginst3471 (P1_R1171_U468, P1_R1171_U58, P1_U3506);
  nand ginst3472 (P1_R1171_U469, P1_R1171_U467, P1_R1171_U468);
  not ginst3473 (P1_R1171_U47, P1_U4018);
  nand ginst3474 (P1_R1171_U470, P1_R1171_U358, P1_R1171_U93);
  nand ginst3475 (P1_R1171_U471, P1_R1171_U259, P1_R1171_U469);
  nand ginst3476 (P1_R1171_U472, P1_R1171_U74, P1_U3074);
  nand ginst3477 (P1_R1171_U473, P1_R1171_U75, P1_U3503);
  nand ginst3478 (P1_R1171_U474, P1_R1171_U74, P1_U3074);
  nand ginst3479 (P1_R1171_U475, P1_R1171_U75, P1_U3503);
  nand ginst3480 (P1_R1171_U476, P1_R1171_U474, P1_R1171_U475);
  nand ginst3481 (P1_R1171_U477, P1_R1171_U160, P1_R1171_U161);
  nand ginst3482 (P1_R1171_U478, P1_R1171_U255, P1_R1171_U476);
  nand ginst3483 (P1_R1171_U479, P1_R1171_U72, P1_U3079);
  not ginst3484 (P1_R1171_U48, P1_U3053);
  nand ginst3485 (P1_R1171_U480, P1_R1171_U73, P1_U3500);
  nand ginst3486 (P1_R1171_U481, P1_R1171_U72, P1_U3079);
  nand ginst3487 (P1_R1171_U482, P1_R1171_U73, P1_U3500);
  nand ginst3488 (P1_R1171_U483, P1_R1171_U481, P1_R1171_U482);
  nand ginst3489 (P1_R1171_U484, P1_R1171_U162, P1_R1171_U163);
  nand ginst3490 (P1_R1171_U485, P1_R1171_U251, P1_R1171_U483);
  nand ginst3491 (P1_R1171_U486, P1_R1171_U70, P1_U3080);
  nand ginst3492 (P1_R1171_U487, P1_R1171_U71, P1_U3497);
  nand ginst3493 (P1_R1171_U488, P1_R1171_U65, P1_U3072);
  nand ginst3494 (P1_R1171_U489, P1_R1171_U66, P1_U3494);
  not ginst3495 (P1_R1171_U49, P1_U3057);
  nand ginst3496 (P1_R1171_U490, P1_R1171_U488, P1_R1171_U489);
  nand ginst3497 (P1_R1171_U491, P1_R1171_U359, P1_R1171_U94);
  nand ginst3498 (P1_R1171_U492, P1_R1171_U335, P1_R1171_U490);
  nand ginst3499 (P1_R1171_U493, P1_R1171_U67, P1_U3063);
  nand ginst3500 (P1_R1171_U494, P1_R1171_U68, P1_U3491);
  nand ginst3501 (P1_R1171_U495, P1_R1171_U493, P1_R1171_U494);
  nand ginst3502 (P1_R1171_U496, P1_R1171_U164, P1_R1171_U360);
  nand ginst3503 (P1_R1171_U497, P1_R1171_U241, P1_R1171_U495);
  nand ginst3504 (P1_R1171_U498, P1_R1171_U63, P1_U3062);
  nand ginst3505 (P1_R1171_U499, P1_R1171_U64, P1_U3488);
  and ginst3506 (P1_R1171_U5, P1_R1171_U177, P1_R1171_U178);
  not ginst3507 (P1_R1171_U50, P1_U4019);
  nand ginst3508 (P1_R1171_U500, P1_R1171_U30, P1_U3077);
  nand ginst3509 (P1_R1171_U501, P1_R1171_U31, P1_U3456);
  not ginst3510 (P1_R1171_U51, P1_U4020);
  not ginst3511 (P1_R1171_U52, P1_U3058);
  not ginst3512 (P1_R1171_U53, P1_U4021);
  not ginst3513 (P1_R1171_U54, P1_U3065);
  not ginst3514 (P1_R1171_U55, P1_U4024);
  not ginst3515 (P1_R1171_U56, P1_U3075);
  not ginst3516 (P1_R1171_U57, P1_U3506);
  not ginst3517 (P1_R1171_U58, P1_U3073);
  not ginst3518 (P1_R1171_U59, P1_U3069);
  and ginst3519 (P1_R1171_U6, P1_R1171_U193, P1_R1171_U194);
  nand ginst3520 (P1_R1171_U60, P1_U3073, P1_U3506);
  not ginst3521 (P1_R1171_U61, P1_U3509);
  nand ginst3522 (P1_R1171_U62, P1_U3084, P1_U3482);
  not ginst3523 (P1_R1171_U63, P1_U3488);
  not ginst3524 (P1_R1171_U64, P1_U3062);
  not ginst3525 (P1_R1171_U65, P1_U3494);
  not ginst3526 (P1_R1171_U66, P1_U3072);
  not ginst3527 (P1_R1171_U67, P1_U3491);
  not ginst3528 (P1_R1171_U68, P1_U3063);
  nand ginst3529 (P1_R1171_U69, P1_U3063, P1_U3491);
  and ginst3530 (P1_R1171_U7, P1_R1171_U233, P1_R1171_U234);
  not ginst3531 (P1_R1171_U70, P1_U3497);
  not ginst3532 (P1_R1171_U71, P1_U3080);
  not ginst3533 (P1_R1171_U72, P1_U3500);
  not ginst3534 (P1_R1171_U73, P1_U3079);
  not ginst3535 (P1_R1171_U74, P1_U3503);
  not ginst3536 (P1_R1171_U75, P1_U3074);
  not ginst3537 (P1_R1171_U76, P1_U3512);
  not ginst3538 (P1_R1171_U77, P1_U3082);
  nand ginst3539 (P1_R1171_U78, P1_U3082, P1_U3512);
  not ginst3540 (P1_R1171_U79, P1_U3514);
  and ginst3541 (P1_R1171_U8, P1_R1171_U242, P1_R1171_U243);
  not ginst3542 (P1_R1171_U80, P1_U3081);
  nand ginst3543 (P1_R1171_U81, P1_U3081, P1_U3514);
  not ginst3544 (P1_R1171_U82, P1_U4025);
  not ginst3545 (P1_R1171_U83, P1_U4023);
  not ginst3546 (P1_R1171_U84, P1_U3061);
  not ginst3547 (P1_R1171_U85, P1_U4022);
  not ginst3548 (P1_R1171_U86, P1_U3066);
  nand ginst3549 (P1_R1171_U87, P1_U3057, P1_U4019);
  not ginst3550 (P1_R1171_U88, P1_U3054);
  not ginst3551 (P1_R1171_U89, P1_U4017);
  and ginst3552 (P1_R1171_U9, P1_R1171_U260, P1_R1171_U261);
  nand ginst3553 (P1_R1171_U90, P1_R1171_U173, P1_R1171_U303);
  not ginst3554 (P1_R1171_U91, P1_U3076);
  nand ginst3555 (P1_R1171_U92, P1_R1171_U312, P1_R1171_U78);
  nand ginst3556 (P1_R1171_U93, P1_R1171_U257, P1_R1171_U258);
  nand ginst3557 (P1_R1171_U94, P1_R1171_U334, P1_R1171_U69);
  nand ginst3558 (P1_R1171_U95, P1_R1171_U453, P1_R1171_U454);
  nand ginst3559 (P1_R1171_U96, P1_R1171_U500, P1_R1171_U501);
  nand ginst3560 (P1_R1171_U97, P1_R1171_U371, P1_R1171_U372);
  nand ginst3561 (P1_R1171_U98, P1_R1171_U376, P1_R1171_U377);
  nand ginst3562 (P1_R1171_U99, P1_R1171_U383, P1_R1171_U384);
  and ginst3563 (P1_R1192_U10, P1_R1192_U258, P1_R1192_U259);
  nand ginst3564 (P1_R1192_U100, P1_R1192_U442, P1_R1192_U443);
  nand ginst3565 (P1_R1192_U101, P1_R1192_U447, P1_R1192_U448);
  nand ginst3566 (P1_R1192_U102, P1_R1192_U463, P1_R1192_U464);
  nand ginst3567 (P1_R1192_U103, P1_R1192_U468, P1_R1192_U469);
  nand ginst3568 (P1_R1192_U104, P1_R1192_U351, P1_R1192_U352);
  nand ginst3569 (P1_R1192_U105, P1_R1192_U360, P1_R1192_U361);
  nand ginst3570 (P1_R1192_U106, P1_R1192_U367, P1_R1192_U368);
  nand ginst3571 (P1_R1192_U107, P1_R1192_U371, P1_R1192_U372);
  nand ginst3572 (P1_R1192_U108, P1_R1192_U380, P1_R1192_U381);
  nand ginst3573 (P1_R1192_U109, P1_R1192_U401, P1_R1192_U402);
  and ginst3574 (P1_R1192_U11, P1_R1192_U284, P1_R1192_U285);
  nand ginst3575 (P1_R1192_U110, P1_R1192_U418, P1_R1192_U419);
  nand ginst3576 (P1_R1192_U111, P1_R1192_U422, P1_R1192_U423);
  nand ginst3577 (P1_R1192_U112, P1_R1192_U454, P1_R1192_U455);
  nand ginst3578 (P1_R1192_U113, P1_R1192_U458, P1_R1192_U459);
  nand ginst3579 (P1_R1192_U114, P1_R1192_U475, P1_R1192_U476);
  and ginst3580 (P1_R1192_U115, P1_R1192_U183, P1_R1192_U195);
  and ginst3581 (P1_R1192_U116, P1_R1192_U198, P1_R1192_U199);
  and ginst3582 (P1_R1192_U117, P1_R1192_U185, P1_R1192_U211);
  and ginst3583 (P1_R1192_U118, P1_R1192_U214, P1_R1192_U215);
  and ginst3584 (P1_R1192_U119, P1_R1192_U353, P1_R1192_U354, P1_R1192_U40);
  and ginst3585 (P1_R1192_U12, P1_R1192_U382, P1_R1192_U383);
  and ginst3586 (P1_R1192_U120, P1_R1192_U185, P1_R1192_U357);
  and ginst3587 (P1_R1192_U121, P1_R1192_U230, P1_R1192_U7);
  and ginst3588 (P1_R1192_U122, P1_R1192_U184, P1_R1192_U364);
  and ginst3589 (P1_R1192_U123, P1_R1192_U29, P1_R1192_U373, P1_R1192_U374);
  and ginst3590 (P1_R1192_U124, P1_R1192_U183, P1_R1192_U377);
  and ginst3591 (P1_R1192_U125, P1_R1192_U217, P1_R1192_U8);
  and ginst3592 (P1_R1192_U126, P1_R1192_U180, P1_R1192_U262);
  and ginst3593 (P1_R1192_U127, P1_R1192_U181, P1_R1192_U288);
  and ginst3594 (P1_R1192_U128, P1_R1192_U304, P1_R1192_U305);
  and ginst3595 (P1_R1192_U129, P1_R1192_U307, P1_R1192_U386);
  nand ginst3596 (P1_R1192_U13, P1_R1192_U340, P1_R1192_U343);
  and ginst3597 (P1_R1192_U130, P1_R1192_U304, P1_R1192_U305, P1_R1192_U308);
  nand ginst3598 (P1_R1192_U131, P1_R1192_U389, P1_R1192_U390);
  and ginst3599 (P1_R1192_U132, P1_R1192_U394, P1_R1192_U395, P1_R1192_U85);
  and ginst3600 (P1_R1192_U133, P1_R1192_U182, P1_R1192_U398);
  nand ginst3601 (P1_R1192_U134, P1_R1192_U403, P1_R1192_U404);
  nand ginst3602 (P1_R1192_U135, P1_R1192_U408, P1_R1192_U409);
  and ginst3603 (P1_R1192_U136, P1_R1192_U181, P1_R1192_U415);
  nand ginst3604 (P1_R1192_U137, P1_R1192_U424, P1_R1192_U425);
  nand ginst3605 (P1_R1192_U138, P1_R1192_U429, P1_R1192_U430);
  nand ginst3606 (P1_R1192_U139, P1_R1192_U434, P1_R1192_U435);
  nand ginst3607 (P1_R1192_U14, P1_R1192_U329, P1_R1192_U332);
  nand ginst3608 (P1_R1192_U140, P1_R1192_U439, P1_R1192_U440);
  nand ginst3609 (P1_R1192_U141, P1_R1192_U444, P1_R1192_U445);
  and ginst3610 (P1_R1192_U142, P1_R1192_U180, P1_R1192_U451);
  nand ginst3611 (P1_R1192_U143, P1_R1192_U460, P1_R1192_U461);
  nand ginst3612 (P1_R1192_U144, P1_R1192_U465, P1_R1192_U466);
  and ginst3613 (P1_R1192_U145, P1_R1192_U342, P1_R1192_U9);
  and ginst3614 (P1_R1192_U146, P1_R1192_U179, P1_R1192_U472);
  and ginst3615 (P1_R1192_U147, P1_R1192_U349, P1_R1192_U350);
  nand ginst3616 (P1_R1192_U148, P1_R1192_U118, P1_R1192_U212);
  and ginst3617 (P1_R1192_U149, P1_R1192_U358, P1_R1192_U359);
  nand ginst3618 (P1_R1192_U15, P1_R1192_U318, P1_R1192_U321);
  and ginst3619 (P1_R1192_U150, P1_R1192_U365, P1_R1192_U366);
  and ginst3620 (P1_R1192_U151, P1_R1192_U369, P1_R1192_U370);
  nand ginst3621 (P1_R1192_U152, P1_R1192_U116, P1_R1192_U196);
  and ginst3622 (P1_R1192_U153, P1_R1192_U378, P1_R1192_U379);
  not ginst3623 (P1_R1192_U154, P1_U4028);
  not ginst3624 (P1_R1192_U155, P1_U3055);
  and ginst3625 (P1_R1192_U156, P1_R1192_U387, P1_R1192_U388);
  nand ginst3626 (P1_R1192_U157, P1_R1192_U128, P1_R1192_U302);
  and ginst3627 (P1_R1192_U158, P1_R1192_U399, P1_R1192_U400);
  nand ginst3628 (P1_R1192_U159, P1_R1192_U294, P1_R1192_U295);
  nand ginst3629 (P1_R1192_U16, P1_R1192_U310, P1_R1192_U312);
  nand ginst3630 (P1_R1192_U160, P1_R1192_U290, P1_R1192_U291);
  and ginst3631 (P1_R1192_U161, P1_R1192_U416, P1_R1192_U417);
  and ginst3632 (P1_R1192_U162, P1_R1192_U420, P1_R1192_U421);
  nand ginst3633 (P1_R1192_U163, P1_R1192_U280, P1_R1192_U281);
  nand ginst3634 (P1_R1192_U164, P1_R1192_U276, P1_R1192_U277);
  not ginst3635 (P1_R1192_U165, P1_U3461);
  nand ginst3636 (P1_R1192_U166, P1_R1192_U272, P1_R1192_U273);
  not ginst3637 (P1_R1192_U167, P1_U3512);
  nand ginst3638 (P1_R1192_U168, P1_R1192_U264, P1_R1192_U265);
  and ginst3639 (P1_R1192_U169, P1_R1192_U452, P1_R1192_U453);
  nand ginst3640 (P1_R1192_U17, P1_R1192_U156, P1_R1192_U175, P1_R1192_U348);
  and ginst3641 (P1_R1192_U170, P1_R1192_U456, P1_R1192_U457);
  nand ginst3642 (P1_R1192_U171, P1_R1192_U254, P1_R1192_U255);
  nand ginst3643 (P1_R1192_U172, P1_R1192_U250, P1_R1192_U251);
  nand ginst3644 (P1_R1192_U173, P1_R1192_U246, P1_R1192_U247);
  and ginst3645 (P1_R1192_U174, P1_R1192_U473, P1_R1192_U474);
  nand ginst3646 (P1_R1192_U175, P1_R1192_U129, P1_R1192_U157);
  not ginst3647 (P1_R1192_U176, P1_R1192_U85);
  not ginst3648 (P1_R1192_U177, P1_R1192_U29);
  not ginst3649 (P1_R1192_U178, P1_R1192_U40);
  nand ginst3650 (P1_R1192_U179, P1_R1192_U53, P1_U3488);
  nand ginst3651 (P1_R1192_U18, P1_R1192_U236, P1_R1192_U238);
  nand ginst3652 (P1_R1192_U180, P1_R1192_U62, P1_U3503);
  nand ginst3653 (P1_R1192_U181, P1_R1192_U76, P1_U4023);
  nand ginst3654 (P1_R1192_U182, P1_R1192_U84, P1_U4019);
  nand ginst3655 (P1_R1192_U183, P1_R1192_U28, P1_U3464);
  nand ginst3656 (P1_R1192_U184, P1_R1192_U35, P1_U3473);
  nand ginst3657 (P1_R1192_U185, P1_R1192_U39, P1_U3479);
  not ginst3658 (P1_R1192_U186, P1_R1192_U64);
  not ginst3659 (P1_R1192_U187, P1_R1192_U78);
  not ginst3660 (P1_R1192_U188, P1_R1192_U37);
  not ginst3661 (P1_R1192_U189, P1_R1192_U54);
  nand ginst3662 (P1_R1192_U19, P1_R1192_U228, P1_R1192_U231);
  not ginst3663 (P1_R1192_U190, P1_R1192_U25);
  nand ginst3664 (P1_R1192_U191, P1_R1192_U190, P1_R1192_U26);
  nand ginst3665 (P1_R1192_U192, P1_R1192_U165, P1_R1192_U191);
  nand ginst3666 (P1_R1192_U193, P1_R1192_U25, P1_U3078);
  not ginst3667 (P1_R1192_U194, P1_R1192_U46);
  nand ginst3668 (P1_R1192_U195, P1_R1192_U30, P1_U3467);
  nand ginst3669 (P1_R1192_U196, P1_R1192_U115, P1_R1192_U46);
  nand ginst3670 (P1_R1192_U197, P1_R1192_U29, P1_R1192_U30);
  nand ginst3671 (P1_R1192_U198, P1_R1192_U197, P1_R1192_U27);
  nand ginst3672 (P1_R1192_U199, P1_R1192_U177, P1_U3064);
  nand ginst3673 (P1_R1192_U20, P1_R1192_U220, P1_R1192_U222);
  not ginst3674 (P1_R1192_U200, P1_R1192_U152);
  nand ginst3675 (P1_R1192_U201, P1_R1192_U34, P1_U3476);
  nand ginst3676 (P1_R1192_U202, P1_R1192_U31, P1_U3071);
  nand ginst3677 (P1_R1192_U203, P1_R1192_U32, P1_U3067);
  nand ginst3678 (P1_R1192_U204, P1_R1192_U188, P1_R1192_U6);
  nand ginst3679 (P1_R1192_U205, P1_R1192_U204, P1_R1192_U7);
  nand ginst3680 (P1_R1192_U206, P1_R1192_U36, P1_U3470);
  nand ginst3681 (P1_R1192_U207, P1_R1192_U34, P1_U3476);
  nand ginst3682 (P1_R1192_U208, P1_R1192_U152, P1_R1192_U206, P1_R1192_U6);
  nand ginst3683 (P1_R1192_U209, P1_R1192_U205, P1_R1192_U207);
  nand ginst3684 (P1_R1192_U21, P1_R1192_U25, P1_R1192_U346);
  not ginst3685 (P1_R1192_U210, P1_R1192_U44);
  nand ginst3686 (P1_R1192_U211, P1_R1192_U41, P1_U3482);
  nand ginst3687 (P1_R1192_U212, P1_R1192_U117, P1_R1192_U44);
  nand ginst3688 (P1_R1192_U213, P1_R1192_U40, P1_R1192_U41);
  nand ginst3689 (P1_R1192_U214, P1_R1192_U213, P1_R1192_U38);
  nand ginst3690 (P1_R1192_U215, P1_R1192_U178, P1_U3084);
  not ginst3691 (P1_R1192_U216, P1_R1192_U148);
  nand ginst3692 (P1_R1192_U217, P1_R1192_U43, P1_U3485);
  nand ginst3693 (P1_R1192_U218, P1_R1192_U217, P1_R1192_U54);
  nand ginst3694 (P1_R1192_U219, P1_R1192_U210, P1_R1192_U40);
  not ginst3695 (P1_R1192_U22, P1_U3479);
  nand ginst3696 (P1_R1192_U220, P1_R1192_U120, P1_R1192_U219);
  nand ginst3697 (P1_R1192_U221, P1_R1192_U185, P1_R1192_U44);
  nand ginst3698 (P1_R1192_U222, P1_R1192_U119, P1_R1192_U221);
  nand ginst3699 (P1_R1192_U223, P1_R1192_U185, P1_R1192_U40);
  nand ginst3700 (P1_R1192_U224, P1_R1192_U152, P1_R1192_U206);
  not ginst3701 (P1_R1192_U225, P1_R1192_U45);
  nand ginst3702 (P1_R1192_U226, P1_R1192_U32, P1_U3067);
  nand ginst3703 (P1_R1192_U227, P1_R1192_U225, P1_R1192_U226);
  nand ginst3704 (P1_R1192_U228, P1_R1192_U122, P1_R1192_U227);
  nand ginst3705 (P1_R1192_U229, P1_R1192_U184, P1_R1192_U45);
  not ginst3706 (P1_R1192_U23, P1_U3464);
  nand ginst3707 (P1_R1192_U230, P1_R1192_U34, P1_U3476);
  nand ginst3708 (P1_R1192_U231, P1_R1192_U121, P1_R1192_U229);
  nand ginst3709 (P1_R1192_U232, P1_R1192_U32, P1_U3067);
  nand ginst3710 (P1_R1192_U233, P1_R1192_U184, P1_R1192_U232);
  nand ginst3711 (P1_R1192_U234, P1_R1192_U206, P1_R1192_U37);
  nand ginst3712 (P1_R1192_U235, P1_R1192_U194, P1_R1192_U29);
  nand ginst3713 (P1_R1192_U236, P1_R1192_U124, P1_R1192_U235);
  nand ginst3714 (P1_R1192_U237, P1_R1192_U183, P1_R1192_U46);
  nand ginst3715 (P1_R1192_U238, P1_R1192_U123, P1_R1192_U237);
  nand ginst3716 (P1_R1192_U239, P1_R1192_U183, P1_R1192_U29);
  not ginst3717 (P1_R1192_U24, P1_U3456);
  nand ginst3718 (P1_R1192_U240, P1_R1192_U52, P1_U3491);
  nand ginst3719 (P1_R1192_U241, P1_R1192_U50, P1_U3063);
  nand ginst3720 (P1_R1192_U242, P1_R1192_U51, P1_U3062);
  nand ginst3721 (P1_R1192_U243, P1_R1192_U189, P1_R1192_U8);
  nand ginst3722 (P1_R1192_U244, P1_R1192_U243, P1_R1192_U9);
  nand ginst3723 (P1_R1192_U245, P1_R1192_U52, P1_U3491);
  nand ginst3724 (P1_R1192_U246, P1_R1192_U125, P1_R1192_U148);
  nand ginst3725 (P1_R1192_U247, P1_R1192_U244, P1_R1192_U245);
  not ginst3726 (P1_R1192_U248, P1_R1192_U173);
  nand ginst3727 (P1_R1192_U249, P1_R1192_U56, P1_U3494);
  nand ginst3728 (P1_R1192_U25, P1_R1192_U93, P1_U3456);
  nand ginst3729 (P1_R1192_U250, P1_R1192_U173, P1_R1192_U249);
  nand ginst3730 (P1_R1192_U251, P1_R1192_U55, P1_U3072);
  not ginst3731 (P1_R1192_U252, P1_R1192_U172);
  nand ginst3732 (P1_R1192_U253, P1_R1192_U58, P1_U3497);
  nand ginst3733 (P1_R1192_U254, P1_R1192_U172, P1_R1192_U253);
  nand ginst3734 (P1_R1192_U255, P1_R1192_U57, P1_U3080);
  not ginst3735 (P1_R1192_U256, P1_R1192_U171);
  nand ginst3736 (P1_R1192_U257, P1_R1192_U61, P1_U3506);
  nand ginst3737 (P1_R1192_U258, P1_R1192_U59, P1_U3073);
  nand ginst3738 (P1_R1192_U259, P1_R1192_U49, P1_U3074);
  not ginst3739 (P1_R1192_U26, P1_U3078);
  nand ginst3740 (P1_R1192_U260, P1_R1192_U180, P1_R1192_U186);
  nand ginst3741 (P1_R1192_U261, P1_R1192_U10, P1_R1192_U260);
  nand ginst3742 (P1_R1192_U262, P1_R1192_U63, P1_U3500);
  nand ginst3743 (P1_R1192_U263, P1_R1192_U61, P1_U3506);
  nand ginst3744 (P1_R1192_U264, P1_R1192_U126, P1_R1192_U171, P1_R1192_U257);
  nand ginst3745 (P1_R1192_U265, P1_R1192_U261, P1_R1192_U263);
  not ginst3746 (P1_R1192_U266, P1_R1192_U168);
  nand ginst3747 (P1_R1192_U267, P1_R1192_U66, P1_U3509);
  nand ginst3748 (P1_R1192_U268, P1_R1192_U168, P1_R1192_U267);
  nand ginst3749 (P1_R1192_U269, P1_R1192_U65, P1_U3069);
  not ginst3750 (P1_R1192_U27, P1_U3467);
  not ginst3751 (P1_R1192_U270, P1_R1192_U67);
  nand ginst3752 (P1_R1192_U271, P1_R1192_U270, P1_R1192_U68);
  nand ginst3753 (P1_R1192_U272, P1_R1192_U167, P1_R1192_U271);
  nand ginst3754 (P1_R1192_U273, P1_R1192_U67, P1_U3082);
  not ginst3755 (P1_R1192_U274, P1_R1192_U166);
  nand ginst3756 (P1_R1192_U275, P1_R1192_U70, P1_U3514);
  nand ginst3757 (P1_R1192_U276, P1_R1192_U166, P1_R1192_U275);
  nand ginst3758 (P1_R1192_U277, P1_R1192_U69, P1_U3081);
  not ginst3759 (P1_R1192_U278, P1_R1192_U164);
  nand ginst3760 (P1_R1192_U279, P1_R1192_U72, P1_U4025);
  not ginst3761 (P1_R1192_U28, P1_U3068);
  nand ginst3762 (P1_R1192_U280, P1_R1192_U164, P1_R1192_U279);
  nand ginst3763 (P1_R1192_U281, P1_R1192_U71, P1_U3076);
  not ginst3764 (P1_R1192_U282, P1_R1192_U163);
  nand ginst3765 (P1_R1192_U283, P1_R1192_U75, P1_U4022);
  nand ginst3766 (P1_R1192_U284, P1_R1192_U73, P1_U3066);
  nand ginst3767 (P1_R1192_U285, P1_R1192_U48, P1_U3061);
  nand ginst3768 (P1_R1192_U286, P1_R1192_U181, P1_R1192_U187);
  nand ginst3769 (P1_R1192_U287, P1_R1192_U11, P1_R1192_U286);
  nand ginst3770 (P1_R1192_U288, P1_R1192_U77, P1_U4024);
  nand ginst3771 (P1_R1192_U289, P1_R1192_U75, P1_U4022);
  nand ginst3772 (P1_R1192_U29, P1_R1192_U23, P1_U3068);
  nand ginst3773 (P1_R1192_U290, P1_R1192_U127, P1_R1192_U163, P1_R1192_U283);
  nand ginst3774 (P1_R1192_U291, P1_R1192_U287, P1_R1192_U289);
  not ginst3775 (P1_R1192_U292, P1_R1192_U160);
  nand ginst3776 (P1_R1192_U293, P1_R1192_U80, P1_U4021);
  nand ginst3777 (P1_R1192_U294, P1_R1192_U160, P1_R1192_U293);
  nand ginst3778 (P1_R1192_U295, P1_R1192_U79, P1_U3065);
  not ginst3779 (P1_R1192_U296, P1_R1192_U159);
  nand ginst3780 (P1_R1192_U297, P1_R1192_U82, P1_U4020);
  nand ginst3781 (P1_R1192_U298, P1_R1192_U159, P1_R1192_U297);
  nand ginst3782 (P1_R1192_U299, P1_R1192_U81, P1_U3058);
  not ginst3783 (P1_R1192_U30, P1_U3064);
  not ginst3784 (P1_R1192_U300, P1_R1192_U89);
  nand ginst3785 (P1_R1192_U301, P1_R1192_U86, P1_U4018);
  nand ginst3786 (P1_R1192_U302, P1_R1192_U182, P1_R1192_U301, P1_R1192_U89);
  nand ginst3787 (P1_R1192_U303, P1_R1192_U85, P1_R1192_U86);
  nand ginst3788 (P1_R1192_U304, P1_R1192_U303, P1_R1192_U83);
  nand ginst3789 (P1_R1192_U305, P1_R1192_U176, P1_U3053);
  not ginst3790 (P1_R1192_U306, P1_R1192_U157);
  nand ginst3791 (P1_R1192_U307, P1_R1192_U88, P1_U4017);
  nand ginst3792 (P1_R1192_U308, P1_R1192_U87, P1_U3054);
  nand ginst3793 (P1_R1192_U309, P1_R1192_U300, P1_R1192_U85);
  not ginst3794 (P1_R1192_U31, P1_U3476);
  nand ginst3795 (P1_R1192_U310, P1_R1192_U133, P1_R1192_U309);
  nand ginst3796 (P1_R1192_U311, P1_R1192_U182, P1_R1192_U89);
  nand ginst3797 (P1_R1192_U312, P1_R1192_U132, P1_R1192_U311);
  nand ginst3798 (P1_R1192_U313, P1_R1192_U182, P1_R1192_U85);
  nand ginst3799 (P1_R1192_U314, P1_R1192_U163, P1_R1192_U288);
  not ginst3800 (P1_R1192_U315, P1_R1192_U90);
  nand ginst3801 (P1_R1192_U316, P1_R1192_U48, P1_U3061);
  nand ginst3802 (P1_R1192_U317, P1_R1192_U315, P1_R1192_U316);
  nand ginst3803 (P1_R1192_U318, P1_R1192_U136, P1_R1192_U317);
  nand ginst3804 (P1_R1192_U319, P1_R1192_U181, P1_R1192_U90);
  not ginst3805 (P1_R1192_U32, P1_U3473);
  nand ginst3806 (P1_R1192_U320, P1_R1192_U75, P1_U4022);
  nand ginst3807 (P1_R1192_U321, P1_R1192_U11, P1_R1192_U319, P1_R1192_U320);
  nand ginst3808 (P1_R1192_U322, P1_R1192_U48, P1_U3061);
  nand ginst3809 (P1_R1192_U323, P1_R1192_U181, P1_R1192_U322);
  nand ginst3810 (P1_R1192_U324, P1_R1192_U288, P1_R1192_U78);
  nand ginst3811 (P1_R1192_U325, P1_R1192_U171, P1_R1192_U262);
  not ginst3812 (P1_R1192_U326, P1_R1192_U91);
  nand ginst3813 (P1_R1192_U327, P1_R1192_U49, P1_U3074);
  nand ginst3814 (P1_R1192_U328, P1_R1192_U326, P1_R1192_U327);
  nand ginst3815 (P1_R1192_U329, P1_R1192_U142, P1_R1192_U328);
  not ginst3816 (P1_R1192_U33, P1_U3470);
  nand ginst3817 (P1_R1192_U330, P1_R1192_U180, P1_R1192_U91);
  nand ginst3818 (P1_R1192_U331, P1_R1192_U61, P1_U3506);
  nand ginst3819 (P1_R1192_U332, P1_R1192_U10, P1_R1192_U330, P1_R1192_U331);
  nand ginst3820 (P1_R1192_U333, P1_R1192_U49, P1_U3074);
  nand ginst3821 (P1_R1192_U334, P1_R1192_U180, P1_R1192_U333);
  nand ginst3822 (P1_R1192_U335, P1_R1192_U262, P1_R1192_U64);
  nand ginst3823 (P1_R1192_U336, P1_R1192_U148, P1_R1192_U217);
  not ginst3824 (P1_R1192_U337, P1_R1192_U92);
  nand ginst3825 (P1_R1192_U338, P1_R1192_U51, P1_U3062);
  nand ginst3826 (P1_R1192_U339, P1_R1192_U337, P1_R1192_U338);
  not ginst3827 (P1_R1192_U34, P1_U3071);
  nand ginst3828 (P1_R1192_U340, P1_R1192_U146, P1_R1192_U339);
  nand ginst3829 (P1_R1192_U341, P1_R1192_U179, P1_R1192_U92);
  nand ginst3830 (P1_R1192_U342, P1_R1192_U52, P1_U3491);
  nand ginst3831 (P1_R1192_U343, P1_R1192_U145, P1_R1192_U341);
  nand ginst3832 (P1_R1192_U344, P1_R1192_U51, P1_U3062);
  nand ginst3833 (P1_R1192_U345, P1_R1192_U179, P1_R1192_U344);
  nand ginst3834 (P1_R1192_U346, P1_R1192_U24, P1_U3077);
  nand ginst3835 (P1_R1192_U347, P1_R1192_U182, P1_R1192_U301, P1_R1192_U89);
  nand ginst3836 (P1_R1192_U348, P1_R1192_U12, P1_R1192_U130, P1_R1192_U347);
  nand ginst3837 (P1_R1192_U349, P1_R1192_U43, P1_U3485);
  not ginst3838 (P1_R1192_U35, P1_U3067);
  nand ginst3839 (P1_R1192_U350, P1_R1192_U42, P1_U3083);
  nand ginst3840 (P1_R1192_U351, P1_R1192_U148, P1_R1192_U218);
  nand ginst3841 (P1_R1192_U352, P1_R1192_U147, P1_R1192_U216);
  nand ginst3842 (P1_R1192_U353, P1_R1192_U41, P1_U3482);
  nand ginst3843 (P1_R1192_U354, P1_R1192_U38, P1_U3084);
  nand ginst3844 (P1_R1192_U355, P1_R1192_U41, P1_U3482);
  nand ginst3845 (P1_R1192_U356, P1_R1192_U38, P1_U3084);
  nand ginst3846 (P1_R1192_U357, P1_R1192_U355, P1_R1192_U356);
  nand ginst3847 (P1_R1192_U358, P1_R1192_U39, P1_U3479);
  nand ginst3848 (P1_R1192_U359, P1_R1192_U22, P1_U3070);
  not ginst3849 (P1_R1192_U36, P1_U3060);
  nand ginst3850 (P1_R1192_U360, P1_R1192_U223, P1_R1192_U44);
  nand ginst3851 (P1_R1192_U361, P1_R1192_U149, P1_R1192_U210);
  nand ginst3852 (P1_R1192_U362, P1_R1192_U34, P1_U3476);
  nand ginst3853 (P1_R1192_U363, P1_R1192_U31, P1_U3071);
  nand ginst3854 (P1_R1192_U364, P1_R1192_U362, P1_R1192_U363);
  nand ginst3855 (P1_R1192_U365, P1_R1192_U35, P1_U3473);
  nand ginst3856 (P1_R1192_U366, P1_R1192_U32, P1_U3067);
  nand ginst3857 (P1_R1192_U367, P1_R1192_U233, P1_R1192_U45);
  nand ginst3858 (P1_R1192_U368, P1_R1192_U150, P1_R1192_U225);
  nand ginst3859 (P1_R1192_U369, P1_R1192_U36, P1_U3470);
  nand ginst3860 (P1_R1192_U37, P1_R1192_U33, P1_U3060);
  nand ginst3861 (P1_R1192_U370, P1_R1192_U33, P1_U3060);
  nand ginst3862 (P1_R1192_U371, P1_R1192_U152, P1_R1192_U234);
  nand ginst3863 (P1_R1192_U372, P1_R1192_U151, P1_R1192_U200);
  nand ginst3864 (P1_R1192_U373, P1_R1192_U30, P1_U3467);
  nand ginst3865 (P1_R1192_U374, P1_R1192_U27, P1_U3064);
  nand ginst3866 (P1_R1192_U375, P1_R1192_U30, P1_U3467);
  nand ginst3867 (P1_R1192_U376, P1_R1192_U27, P1_U3064);
  nand ginst3868 (P1_R1192_U377, P1_R1192_U375, P1_R1192_U376);
  nand ginst3869 (P1_R1192_U378, P1_R1192_U28, P1_U3464);
  nand ginst3870 (P1_R1192_U379, P1_R1192_U23, P1_U3068);
  not ginst3871 (P1_R1192_U38, P1_U3482);
  nand ginst3872 (P1_R1192_U380, P1_R1192_U239, P1_R1192_U46);
  nand ginst3873 (P1_R1192_U381, P1_R1192_U153, P1_R1192_U194);
  nand ginst3874 (P1_R1192_U382, P1_R1192_U155, P1_U4028);
  nand ginst3875 (P1_R1192_U383, P1_R1192_U154, P1_U3055);
  nand ginst3876 (P1_R1192_U384, P1_R1192_U155, P1_U4028);
  nand ginst3877 (P1_R1192_U385, P1_R1192_U154, P1_U3055);
  nand ginst3878 (P1_R1192_U386, P1_R1192_U384, P1_R1192_U385);
  nand ginst3879 (P1_R1192_U387, P1_R1192_U386, P1_R1192_U87, P1_U3054);
  nand ginst3880 (P1_R1192_U388, P1_R1192_U12, P1_R1192_U88, P1_U4017);
  nand ginst3881 (P1_R1192_U389, P1_R1192_U88, P1_U4017);
  not ginst3882 (P1_R1192_U39, P1_U3070);
  nand ginst3883 (P1_R1192_U390, P1_R1192_U87, P1_U3054);
  not ginst3884 (P1_R1192_U391, P1_R1192_U131);
  nand ginst3885 (P1_R1192_U392, P1_R1192_U306, P1_R1192_U391);
  nand ginst3886 (P1_R1192_U393, P1_R1192_U131, P1_R1192_U157);
  nand ginst3887 (P1_R1192_U394, P1_R1192_U86, P1_U4018);
  nand ginst3888 (P1_R1192_U395, P1_R1192_U83, P1_U3053);
  nand ginst3889 (P1_R1192_U396, P1_R1192_U86, P1_U4018);
  nand ginst3890 (P1_R1192_U397, P1_R1192_U83, P1_U3053);
  nand ginst3891 (P1_R1192_U398, P1_R1192_U396, P1_R1192_U397);
  nand ginst3892 (P1_R1192_U399, P1_R1192_U84, P1_U4019);
  nand ginst3893 (P1_R1192_U40, P1_R1192_U22, P1_U3070);
  nand ginst3894 (P1_R1192_U400, P1_R1192_U47, P1_U3057);
  nand ginst3895 (P1_R1192_U401, P1_R1192_U313, P1_R1192_U89);
  nand ginst3896 (P1_R1192_U402, P1_R1192_U158, P1_R1192_U300);
  nand ginst3897 (P1_R1192_U403, P1_R1192_U82, P1_U4020);
  nand ginst3898 (P1_R1192_U404, P1_R1192_U81, P1_U3058);
  not ginst3899 (P1_R1192_U405, P1_R1192_U134);
  nand ginst3900 (P1_R1192_U406, P1_R1192_U296, P1_R1192_U405);
  nand ginst3901 (P1_R1192_U407, P1_R1192_U134, P1_R1192_U159);
  nand ginst3902 (P1_R1192_U408, P1_R1192_U80, P1_U4021);
  nand ginst3903 (P1_R1192_U409, P1_R1192_U79, P1_U3065);
  not ginst3904 (P1_R1192_U41, P1_U3084);
  not ginst3905 (P1_R1192_U410, P1_R1192_U135);
  nand ginst3906 (P1_R1192_U411, P1_R1192_U292, P1_R1192_U410);
  nand ginst3907 (P1_R1192_U412, P1_R1192_U135, P1_R1192_U160);
  nand ginst3908 (P1_R1192_U413, P1_R1192_U75, P1_U4022);
  nand ginst3909 (P1_R1192_U414, P1_R1192_U73, P1_U3066);
  nand ginst3910 (P1_R1192_U415, P1_R1192_U413, P1_R1192_U414);
  nand ginst3911 (P1_R1192_U416, P1_R1192_U76, P1_U4023);
  nand ginst3912 (P1_R1192_U417, P1_R1192_U48, P1_U3061);
  nand ginst3913 (P1_R1192_U418, P1_R1192_U323, P1_R1192_U90);
  nand ginst3914 (P1_R1192_U419, P1_R1192_U161, P1_R1192_U315);
  not ginst3915 (P1_R1192_U42, P1_U3485);
  nand ginst3916 (P1_R1192_U420, P1_R1192_U77, P1_U4024);
  nand ginst3917 (P1_R1192_U421, P1_R1192_U74, P1_U3075);
  nand ginst3918 (P1_R1192_U422, P1_R1192_U163, P1_R1192_U324);
  nand ginst3919 (P1_R1192_U423, P1_R1192_U162, P1_R1192_U282);
  nand ginst3920 (P1_R1192_U424, P1_R1192_U72, P1_U4025);
  nand ginst3921 (P1_R1192_U425, P1_R1192_U71, P1_U3076);
  not ginst3922 (P1_R1192_U426, P1_R1192_U137);
  nand ginst3923 (P1_R1192_U427, P1_R1192_U278, P1_R1192_U426);
  nand ginst3924 (P1_R1192_U428, P1_R1192_U137, P1_R1192_U164);
  nand ginst3925 (P1_R1192_U429, P1_R1192_U26, P1_U3461);
  not ginst3926 (P1_R1192_U43, P1_U3083);
  nand ginst3927 (P1_R1192_U430, P1_R1192_U165, P1_U3078);
  not ginst3928 (P1_R1192_U431, P1_R1192_U138);
  nand ginst3929 (P1_R1192_U432, P1_R1192_U190, P1_R1192_U431);
  nand ginst3930 (P1_R1192_U433, P1_R1192_U138, P1_R1192_U25);
  nand ginst3931 (P1_R1192_U434, P1_R1192_U70, P1_U3514);
  nand ginst3932 (P1_R1192_U435, P1_R1192_U69, P1_U3081);
  not ginst3933 (P1_R1192_U436, P1_R1192_U139);
  nand ginst3934 (P1_R1192_U437, P1_R1192_U274, P1_R1192_U436);
  nand ginst3935 (P1_R1192_U438, P1_R1192_U139, P1_R1192_U166);
  nand ginst3936 (P1_R1192_U439, P1_R1192_U68, P1_U3512);
  nand ginst3937 (P1_R1192_U44, P1_R1192_U208, P1_R1192_U209);
  nand ginst3938 (P1_R1192_U440, P1_R1192_U167, P1_U3082);
  not ginst3939 (P1_R1192_U441, P1_R1192_U140);
  nand ginst3940 (P1_R1192_U442, P1_R1192_U270, P1_R1192_U441);
  nand ginst3941 (P1_R1192_U443, P1_R1192_U140, P1_R1192_U67);
  nand ginst3942 (P1_R1192_U444, P1_R1192_U66, P1_U3509);
  nand ginst3943 (P1_R1192_U445, P1_R1192_U65, P1_U3069);
  not ginst3944 (P1_R1192_U446, P1_R1192_U141);
  nand ginst3945 (P1_R1192_U447, P1_R1192_U266, P1_R1192_U446);
  nand ginst3946 (P1_R1192_U448, P1_R1192_U141, P1_R1192_U168);
  nand ginst3947 (P1_R1192_U449, P1_R1192_U61, P1_U3506);
  nand ginst3948 (P1_R1192_U45, P1_R1192_U224, P1_R1192_U37);
  nand ginst3949 (P1_R1192_U450, P1_R1192_U59, P1_U3073);
  nand ginst3950 (P1_R1192_U451, P1_R1192_U449, P1_R1192_U450);
  nand ginst3951 (P1_R1192_U452, P1_R1192_U62, P1_U3503);
  nand ginst3952 (P1_R1192_U453, P1_R1192_U49, P1_U3074);
  nand ginst3953 (P1_R1192_U454, P1_R1192_U334, P1_R1192_U91);
  nand ginst3954 (P1_R1192_U455, P1_R1192_U169, P1_R1192_U326);
  nand ginst3955 (P1_R1192_U456, P1_R1192_U63, P1_U3500);
  nand ginst3956 (P1_R1192_U457, P1_R1192_U60, P1_U3079);
  nand ginst3957 (P1_R1192_U458, P1_R1192_U171, P1_R1192_U335);
  nand ginst3958 (P1_R1192_U459, P1_R1192_U170, P1_R1192_U256);
  nand ginst3959 (P1_R1192_U46, P1_R1192_U192, P1_R1192_U193);
  nand ginst3960 (P1_R1192_U460, P1_R1192_U58, P1_U3497);
  nand ginst3961 (P1_R1192_U461, P1_R1192_U57, P1_U3080);
  not ginst3962 (P1_R1192_U462, P1_R1192_U143);
  nand ginst3963 (P1_R1192_U463, P1_R1192_U252, P1_R1192_U462);
  nand ginst3964 (P1_R1192_U464, P1_R1192_U143, P1_R1192_U172);
  nand ginst3965 (P1_R1192_U465, P1_R1192_U56, P1_U3494);
  nand ginst3966 (P1_R1192_U466, P1_R1192_U55, P1_U3072);
  not ginst3967 (P1_R1192_U467, P1_R1192_U144);
  nand ginst3968 (P1_R1192_U468, P1_R1192_U248, P1_R1192_U467);
  nand ginst3969 (P1_R1192_U469, P1_R1192_U144, P1_R1192_U173);
  not ginst3970 (P1_R1192_U47, P1_U4019);
  nand ginst3971 (P1_R1192_U470, P1_R1192_U52, P1_U3491);
  nand ginst3972 (P1_R1192_U471, P1_R1192_U50, P1_U3063);
  nand ginst3973 (P1_R1192_U472, P1_R1192_U470, P1_R1192_U471);
  nand ginst3974 (P1_R1192_U473, P1_R1192_U53, P1_U3488);
  nand ginst3975 (P1_R1192_U474, P1_R1192_U51, P1_U3062);
  nand ginst3976 (P1_R1192_U475, P1_R1192_U345, P1_R1192_U92);
  nand ginst3977 (P1_R1192_U476, P1_R1192_U174, P1_R1192_U337);
  not ginst3978 (P1_R1192_U48, P1_U4023);
  not ginst3979 (P1_R1192_U49, P1_U3503);
  not ginst3980 (P1_R1192_U50, P1_U3491);
  not ginst3981 (P1_R1192_U51, P1_U3488);
  not ginst3982 (P1_R1192_U52, P1_U3063);
  not ginst3983 (P1_R1192_U53, P1_U3062);
  nand ginst3984 (P1_R1192_U54, P1_R1192_U42, P1_U3083);
  not ginst3985 (P1_R1192_U55, P1_U3494);
  not ginst3986 (P1_R1192_U56, P1_U3072);
  not ginst3987 (P1_R1192_U57, P1_U3497);
  not ginst3988 (P1_R1192_U58, P1_U3080);
  not ginst3989 (P1_R1192_U59, P1_U3506);
  and ginst3990 (P1_R1192_U6, P1_R1192_U184, P1_R1192_U201);
  not ginst3991 (P1_R1192_U60, P1_U3500);
  not ginst3992 (P1_R1192_U61, P1_U3073);
  not ginst3993 (P1_R1192_U62, P1_U3074);
  not ginst3994 (P1_R1192_U63, P1_U3079);
  nand ginst3995 (P1_R1192_U64, P1_R1192_U60, P1_U3079);
  not ginst3996 (P1_R1192_U65, P1_U3509);
  not ginst3997 (P1_R1192_U66, P1_U3069);
  nand ginst3998 (P1_R1192_U67, P1_R1192_U268, P1_R1192_U269);
  not ginst3999 (P1_R1192_U68, P1_U3082);
  not ginst4000 (P1_R1192_U69, P1_U3514);
  and ginst4001 (P1_R1192_U7, P1_R1192_U202, P1_R1192_U203);
  not ginst4002 (P1_R1192_U70, P1_U3081);
  not ginst4003 (P1_R1192_U71, P1_U4025);
  not ginst4004 (P1_R1192_U72, P1_U3076);
  not ginst4005 (P1_R1192_U73, P1_U4022);
  not ginst4006 (P1_R1192_U74, P1_U4024);
  not ginst4007 (P1_R1192_U75, P1_U3066);
  not ginst4008 (P1_R1192_U76, P1_U3061);
  not ginst4009 (P1_R1192_U77, P1_U3075);
  nand ginst4010 (P1_R1192_U78, P1_R1192_U74, P1_U3075);
  not ginst4011 (P1_R1192_U79, P1_U4021);
  and ginst4012 (P1_R1192_U8, P1_R1192_U179, P1_R1192_U240);
  not ginst4013 (P1_R1192_U80, P1_U3065);
  not ginst4014 (P1_R1192_U81, P1_U4020);
  not ginst4015 (P1_R1192_U82, P1_U3058);
  not ginst4016 (P1_R1192_U83, P1_U4018);
  not ginst4017 (P1_R1192_U84, P1_U3057);
  nand ginst4018 (P1_R1192_U85, P1_R1192_U47, P1_U3057);
  not ginst4019 (P1_R1192_U86, P1_U3053);
  not ginst4020 (P1_R1192_U87, P1_U4017);
  not ginst4021 (P1_R1192_U88, P1_U3054);
  nand ginst4022 (P1_R1192_U89, P1_R1192_U298, P1_R1192_U299);
  and ginst4023 (P1_R1192_U9, P1_R1192_U241, P1_R1192_U242);
  nand ginst4024 (P1_R1192_U90, P1_R1192_U314, P1_R1192_U78);
  nand ginst4025 (P1_R1192_U91, P1_R1192_U325, P1_R1192_U64);
  nand ginst4026 (P1_R1192_U92, P1_R1192_U336, P1_R1192_U54);
  not ginst4027 (P1_R1192_U93, P1_U3077);
  nand ginst4028 (P1_R1192_U94, P1_R1192_U392, P1_R1192_U393);
  nand ginst4029 (P1_R1192_U95, P1_R1192_U406, P1_R1192_U407);
  nand ginst4030 (P1_R1192_U96, P1_R1192_U411, P1_R1192_U412);
  nand ginst4031 (P1_R1192_U97, P1_R1192_U427, P1_R1192_U428);
  nand ginst4032 (P1_R1192_U98, P1_R1192_U432, P1_R1192_U433);
  nand ginst4033 (P1_R1192_U99, P1_R1192_U437, P1_R1192_U438);
  and ginst4034 (P1_R1207_U10, P1_R1207_U258, P1_R1207_U259);
  nand ginst4035 (P1_R1207_U100, P1_R1207_U442, P1_R1207_U443);
  nand ginst4036 (P1_R1207_U101, P1_R1207_U447, P1_R1207_U448);
  nand ginst4037 (P1_R1207_U102, P1_R1207_U463, P1_R1207_U464);
  nand ginst4038 (P1_R1207_U103, P1_R1207_U468, P1_R1207_U469);
  nand ginst4039 (P1_R1207_U104, P1_R1207_U351, P1_R1207_U352);
  nand ginst4040 (P1_R1207_U105, P1_R1207_U360, P1_R1207_U361);
  nand ginst4041 (P1_R1207_U106, P1_R1207_U367, P1_R1207_U368);
  nand ginst4042 (P1_R1207_U107, P1_R1207_U371, P1_R1207_U372);
  nand ginst4043 (P1_R1207_U108, P1_R1207_U380, P1_R1207_U381);
  nand ginst4044 (P1_R1207_U109, P1_R1207_U401, P1_R1207_U402);
  and ginst4045 (P1_R1207_U11, P1_R1207_U284, P1_R1207_U285);
  nand ginst4046 (P1_R1207_U110, P1_R1207_U418, P1_R1207_U419);
  nand ginst4047 (P1_R1207_U111, P1_R1207_U422, P1_R1207_U423);
  nand ginst4048 (P1_R1207_U112, P1_R1207_U454, P1_R1207_U455);
  nand ginst4049 (P1_R1207_U113, P1_R1207_U458, P1_R1207_U459);
  nand ginst4050 (P1_R1207_U114, P1_R1207_U475, P1_R1207_U476);
  and ginst4051 (P1_R1207_U115, P1_R1207_U183, P1_R1207_U195);
  and ginst4052 (P1_R1207_U116, P1_R1207_U198, P1_R1207_U199);
  and ginst4053 (P1_R1207_U117, P1_R1207_U185, P1_R1207_U211);
  and ginst4054 (P1_R1207_U118, P1_R1207_U214, P1_R1207_U215);
  and ginst4055 (P1_R1207_U119, P1_R1207_U353, P1_R1207_U354, P1_R1207_U40);
  and ginst4056 (P1_R1207_U12, P1_R1207_U382, P1_R1207_U383);
  and ginst4057 (P1_R1207_U120, P1_R1207_U185, P1_R1207_U357);
  and ginst4058 (P1_R1207_U121, P1_R1207_U230, P1_R1207_U7);
  and ginst4059 (P1_R1207_U122, P1_R1207_U184, P1_R1207_U364);
  and ginst4060 (P1_R1207_U123, P1_R1207_U29, P1_R1207_U373, P1_R1207_U374);
  and ginst4061 (P1_R1207_U124, P1_R1207_U183, P1_R1207_U377);
  and ginst4062 (P1_R1207_U125, P1_R1207_U217, P1_R1207_U8);
  and ginst4063 (P1_R1207_U126, P1_R1207_U180, P1_R1207_U262);
  and ginst4064 (P1_R1207_U127, P1_R1207_U181, P1_R1207_U288);
  and ginst4065 (P1_R1207_U128, P1_R1207_U304, P1_R1207_U305);
  and ginst4066 (P1_R1207_U129, P1_R1207_U307, P1_R1207_U386);
  nand ginst4067 (P1_R1207_U13, P1_R1207_U340, P1_R1207_U343);
  and ginst4068 (P1_R1207_U130, P1_R1207_U304, P1_R1207_U305, P1_R1207_U308);
  nand ginst4069 (P1_R1207_U131, P1_R1207_U389, P1_R1207_U390);
  and ginst4070 (P1_R1207_U132, P1_R1207_U394, P1_R1207_U395, P1_R1207_U85);
  and ginst4071 (P1_R1207_U133, P1_R1207_U182, P1_R1207_U398);
  nand ginst4072 (P1_R1207_U134, P1_R1207_U403, P1_R1207_U404);
  nand ginst4073 (P1_R1207_U135, P1_R1207_U408, P1_R1207_U409);
  and ginst4074 (P1_R1207_U136, P1_R1207_U181, P1_R1207_U415);
  nand ginst4075 (P1_R1207_U137, P1_R1207_U424, P1_R1207_U425);
  nand ginst4076 (P1_R1207_U138, P1_R1207_U429, P1_R1207_U430);
  nand ginst4077 (P1_R1207_U139, P1_R1207_U434, P1_R1207_U435);
  nand ginst4078 (P1_R1207_U14, P1_R1207_U329, P1_R1207_U332);
  nand ginst4079 (P1_R1207_U140, P1_R1207_U439, P1_R1207_U440);
  nand ginst4080 (P1_R1207_U141, P1_R1207_U444, P1_R1207_U445);
  and ginst4081 (P1_R1207_U142, P1_R1207_U180, P1_R1207_U451);
  nand ginst4082 (P1_R1207_U143, P1_R1207_U460, P1_R1207_U461);
  nand ginst4083 (P1_R1207_U144, P1_R1207_U465, P1_R1207_U466);
  and ginst4084 (P1_R1207_U145, P1_R1207_U342, P1_R1207_U9);
  and ginst4085 (P1_R1207_U146, P1_R1207_U179, P1_R1207_U472);
  and ginst4086 (P1_R1207_U147, P1_R1207_U349, P1_R1207_U350);
  nand ginst4087 (P1_R1207_U148, P1_R1207_U118, P1_R1207_U212);
  and ginst4088 (P1_R1207_U149, P1_R1207_U358, P1_R1207_U359);
  nand ginst4089 (P1_R1207_U15, P1_R1207_U318, P1_R1207_U321);
  and ginst4090 (P1_R1207_U150, P1_R1207_U365, P1_R1207_U366);
  and ginst4091 (P1_R1207_U151, P1_R1207_U369, P1_R1207_U370);
  nand ginst4092 (P1_R1207_U152, P1_R1207_U116, P1_R1207_U196);
  and ginst4093 (P1_R1207_U153, P1_R1207_U378, P1_R1207_U379);
  not ginst4094 (P1_R1207_U154, P1_U4028);
  not ginst4095 (P1_R1207_U155, P1_U3055);
  and ginst4096 (P1_R1207_U156, P1_R1207_U387, P1_R1207_U388);
  nand ginst4097 (P1_R1207_U157, P1_R1207_U128, P1_R1207_U302);
  and ginst4098 (P1_R1207_U158, P1_R1207_U399, P1_R1207_U400);
  nand ginst4099 (P1_R1207_U159, P1_R1207_U294, P1_R1207_U295);
  nand ginst4100 (P1_R1207_U16, P1_R1207_U310, P1_R1207_U312);
  nand ginst4101 (P1_R1207_U160, P1_R1207_U290, P1_R1207_U291);
  and ginst4102 (P1_R1207_U161, P1_R1207_U416, P1_R1207_U417);
  and ginst4103 (P1_R1207_U162, P1_R1207_U420, P1_R1207_U421);
  nand ginst4104 (P1_R1207_U163, P1_R1207_U280, P1_R1207_U281);
  nand ginst4105 (P1_R1207_U164, P1_R1207_U276, P1_R1207_U277);
  not ginst4106 (P1_R1207_U165, P1_U3461);
  nand ginst4107 (P1_R1207_U166, P1_R1207_U272, P1_R1207_U273);
  not ginst4108 (P1_R1207_U167, P1_U3512);
  nand ginst4109 (P1_R1207_U168, P1_R1207_U264, P1_R1207_U265);
  and ginst4110 (P1_R1207_U169, P1_R1207_U452, P1_R1207_U453);
  nand ginst4111 (P1_R1207_U17, P1_R1207_U156, P1_R1207_U175, P1_R1207_U348);
  and ginst4112 (P1_R1207_U170, P1_R1207_U456, P1_R1207_U457);
  nand ginst4113 (P1_R1207_U171, P1_R1207_U254, P1_R1207_U255);
  nand ginst4114 (P1_R1207_U172, P1_R1207_U250, P1_R1207_U251);
  nand ginst4115 (P1_R1207_U173, P1_R1207_U246, P1_R1207_U247);
  and ginst4116 (P1_R1207_U174, P1_R1207_U473, P1_R1207_U474);
  nand ginst4117 (P1_R1207_U175, P1_R1207_U129, P1_R1207_U157);
  not ginst4118 (P1_R1207_U176, P1_R1207_U85);
  not ginst4119 (P1_R1207_U177, P1_R1207_U29);
  not ginst4120 (P1_R1207_U178, P1_R1207_U40);
  nand ginst4121 (P1_R1207_U179, P1_R1207_U53, P1_U3488);
  nand ginst4122 (P1_R1207_U18, P1_R1207_U236, P1_R1207_U238);
  nand ginst4123 (P1_R1207_U180, P1_R1207_U62, P1_U3503);
  nand ginst4124 (P1_R1207_U181, P1_R1207_U76, P1_U4023);
  nand ginst4125 (P1_R1207_U182, P1_R1207_U84, P1_U4019);
  nand ginst4126 (P1_R1207_U183, P1_R1207_U28, P1_U3464);
  nand ginst4127 (P1_R1207_U184, P1_R1207_U35, P1_U3473);
  nand ginst4128 (P1_R1207_U185, P1_R1207_U39, P1_U3479);
  not ginst4129 (P1_R1207_U186, P1_R1207_U64);
  not ginst4130 (P1_R1207_U187, P1_R1207_U78);
  not ginst4131 (P1_R1207_U188, P1_R1207_U37);
  not ginst4132 (P1_R1207_U189, P1_R1207_U54);
  nand ginst4133 (P1_R1207_U19, P1_R1207_U228, P1_R1207_U231);
  not ginst4134 (P1_R1207_U190, P1_R1207_U25);
  nand ginst4135 (P1_R1207_U191, P1_R1207_U190, P1_R1207_U26);
  nand ginst4136 (P1_R1207_U192, P1_R1207_U165, P1_R1207_U191);
  nand ginst4137 (P1_R1207_U193, P1_R1207_U25, P1_U3078);
  not ginst4138 (P1_R1207_U194, P1_R1207_U46);
  nand ginst4139 (P1_R1207_U195, P1_R1207_U30, P1_U3467);
  nand ginst4140 (P1_R1207_U196, P1_R1207_U115, P1_R1207_U46);
  nand ginst4141 (P1_R1207_U197, P1_R1207_U29, P1_R1207_U30);
  nand ginst4142 (P1_R1207_U198, P1_R1207_U197, P1_R1207_U27);
  nand ginst4143 (P1_R1207_U199, P1_R1207_U177, P1_U3064);
  nand ginst4144 (P1_R1207_U20, P1_R1207_U220, P1_R1207_U222);
  not ginst4145 (P1_R1207_U200, P1_R1207_U152);
  nand ginst4146 (P1_R1207_U201, P1_R1207_U34, P1_U3476);
  nand ginst4147 (P1_R1207_U202, P1_R1207_U31, P1_U3071);
  nand ginst4148 (P1_R1207_U203, P1_R1207_U32, P1_U3067);
  nand ginst4149 (P1_R1207_U204, P1_R1207_U188, P1_R1207_U6);
  nand ginst4150 (P1_R1207_U205, P1_R1207_U204, P1_R1207_U7);
  nand ginst4151 (P1_R1207_U206, P1_R1207_U36, P1_U3470);
  nand ginst4152 (P1_R1207_U207, P1_R1207_U34, P1_U3476);
  nand ginst4153 (P1_R1207_U208, P1_R1207_U152, P1_R1207_U206, P1_R1207_U6);
  nand ginst4154 (P1_R1207_U209, P1_R1207_U205, P1_R1207_U207);
  nand ginst4155 (P1_R1207_U21, P1_R1207_U25, P1_R1207_U346);
  not ginst4156 (P1_R1207_U210, P1_R1207_U44);
  nand ginst4157 (P1_R1207_U211, P1_R1207_U41, P1_U3482);
  nand ginst4158 (P1_R1207_U212, P1_R1207_U117, P1_R1207_U44);
  nand ginst4159 (P1_R1207_U213, P1_R1207_U40, P1_R1207_U41);
  nand ginst4160 (P1_R1207_U214, P1_R1207_U213, P1_R1207_U38);
  nand ginst4161 (P1_R1207_U215, P1_R1207_U178, P1_U3084);
  not ginst4162 (P1_R1207_U216, P1_R1207_U148);
  nand ginst4163 (P1_R1207_U217, P1_R1207_U43, P1_U3485);
  nand ginst4164 (P1_R1207_U218, P1_R1207_U217, P1_R1207_U54);
  nand ginst4165 (P1_R1207_U219, P1_R1207_U210, P1_R1207_U40);
  not ginst4166 (P1_R1207_U22, P1_U3479);
  nand ginst4167 (P1_R1207_U220, P1_R1207_U120, P1_R1207_U219);
  nand ginst4168 (P1_R1207_U221, P1_R1207_U185, P1_R1207_U44);
  nand ginst4169 (P1_R1207_U222, P1_R1207_U119, P1_R1207_U221);
  nand ginst4170 (P1_R1207_U223, P1_R1207_U185, P1_R1207_U40);
  nand ginst4171 (P1_R1207_U224, P1_R1207_U152, P1_R1207_U206);
  not ginst4172 (P1_R1207_U225, P1_R1207_U45);
  nand ginst4173 (P1_R1207_U226, P1_R1207_U32, P1_U3067);
  nand ginst4174 (P1_R1207_U227, P1_R1207_U225, P1_R1207_U226);
  nand ginst4175 (P1_R1207_U228, P1_R1207_U122, P1_R1207_U227);
  nand ginst4176 (P1_R1207_U229, P1_R1207_U184, P1_R1207_U45);
  not ginst4177 (P1_R1207_U23, P1_U3464);
  nand ginst4178 (P1_R1207_U230, P1_R1207_U34, P1_U3476);
  nand ginst4179 (P1_R1207_U231, P1_R1207_U121, P1_R1207_U229);
  nand ginst4180 (P1_R1207_U232, P1_R1207_U32, P1_U3067);
  nand ginst4181 (P1_R1207_U233, P1_R1207_U184, P1_R1207_U232);
  nand ginst4182 (P1_R1207_U234, P1_R1207_U206, P1_R1207_U37);
  nand ginst4183 (P1_R1207_U235, P1_R1207_U194, P1_R1207_U29);
  nand ginst4184 (P1_R1207_U236, P1_R1207_U124, P1_R1207_U235);
  nand ginst4185 (P1_R1207_U237, P1_R1207_U183, P1_R1207_U46);
  nand ginst4186 (P1_R1207_U238, P1_R1207_U123, P1_R1207_U237);
  nand ginst4187 (P1_R1207_U239, P1_R1207_U183, P1_R1207_U29);
  not ginst4188 (P1_R1207_U24, P1_U3456);
  nand ginst4189 (P1_R1207_U240, P1_R1207_U52, P1_U3491);
  nand ginst4190 (P1_R1207_U241, P1_R1207_U50, P1_U3063);
  nand ginst4191 (P1_R1207_U242, P1_R1207_U51, P1_U3062);
  nand ginst4192 (P1_R1207_U243, P1_R1207_U189, P1_R1207_U8);
  nand ginst4193 (P1_R1207_U244, P1_R1207_U243, P1_R1207_U9);
  nand ginst4194 (P1_R1207_U245, P1_R1207_U52, P1_U3491);
  nand ginst4195 (P1_R1207_U246, P1_R1207_U125, P1_R1207_U148);
  nand ginst4196 (P1_R1207_U247, P1_R1207_U244, P1_R1207_U245);
  not ginst4197 (P1_R1207_U248, P1_R1207_U173);
  nand ginst4198 (P1_R1207_U249, P1_R1207_U56, P1_U3494);
  nand ginst4199 (P1_R1207_U25, P1_R1207_U93, P1_U3456);
  nand ginst4200 (P1_R1207_U250, P1_R1207_U173, P1_R1207_U249);
  nand ginst4201 (P1_R1207_U251, P1_R1207_U55, P1_U3072);
  not ginst4202 (P1_R1207_U252, P1_R1207_U172);
  nand ginst4203 (P1_R1207_U253, P1_R1207_U58, P1_U3497);
  nand ginst4204 (P1_R1207_U254, P1_R1207_U172, P1_R1207_U253);
  nand ginst4205 (P1_R1207_U255, P1_R1207_U57, P1_U3080);
  not ginst4206 (P1_R1207_U256, P1_R1207_U171);
  nand ginst4207 (P1_R1207_U257, P1_R1207_U61, P1_U3506);
  nand ginst4208 (P1_R1207_U258, P1_R1207_U59, P1_U3073);
  nand ginst4209 (P1_R1207_U259, P1_R1207_U49, P1_U3074);
  not ginst4210 (P1_R1207_U26, P1_U3078);
  nand ginst4211 (P1_R1207_U260, P1_R1207_U180, P1_R1207_U186);
  nand ginst4212 (P1_R1207_U261, P1_R1207_U10, P1_R1207_U260);
  nand ginst4213 (P1_R1207_U262, P1_R1207_U63, P1_U3500);
  nand ginst4214 (P1_R1207_U263, P1_R1207_U61, P1_U3506);
  nand ginst4215 (P1_R1207_U264, P1_R1207_U126, P1_R1207_U171, P1_R1207_U257);
  nand ginst4216 (P1_R1207_U265, P1_R1207_U261, P1_R1207_U263);
  not ginst4217 (P1_R1207_U266, P1_R1207_U168);
  nand ginst4218 (P1_R1207_U267, P1_R1207_U66, P1_U3509);
  nand ginst4219 (P1_R1207_U268, P1_R1207_U168, P1_R1207_U267);
  nand ginst4220 (P1_R1207_U269, P1_R1207_U65, P1_U3069);
  not ginst4221 (P1_R1207_U27, P1_U3467);
  not ginst4222 (P1_R1207_U270, P1_R1207_U67);
  nand ginst4223 (P1_R1207_U271, P1_R1207_U270, P1_R1207_U68);
  nand ginst4224 (P1_R1207_U272, P1_R1207_U167, P1_R1207_U271);
  nand ginst4225 (P1_R1207_U273, P1_R1207_U67, P1_U3082);
  not ginst4226 (P1_R1207_U274, P1_R1207_U166);
  nand ginst4227 (P1_R1207_U275, P1_R1207_U70, P1_U3514);
  nand ginst4228 (P1_R1207_U276, P1_R1207_U166, P1_R1207_U275);
  nand ginst4229 (P1_R1207_U277, P1_R1207_U69, P1_U3081);
  not ginst4230 (P1_R1207_U278, P1_R1207_U164);
  nand ginst4231 (P1_R1207_U279, P1_R1207_U72, P1_U4025);
  not ginst4232 (P1_R1207_U28, P1_U3068);
  nand ginst4233 (P1_R1207_U280, P1_R1207_U164, P1_R1207_U279);
  nand ginst4234 (P1_R1207_U281, P1_R1207_U71, P1_U3076);
  not ginst4235 (P1_R1207_U282, P1_R1207_U163);
  nand ginst4236 (P1_R1207_U283, P1_R1207_U75, P1_U4022);
  nand ginst4237 (P1_R1207_U284, P1_R1207_U73, P1_U3066);
  nand ginst4238 (P1_R1207_U285, P1_R1207_U48, P1_U3061);
  nand ginst4239 (P1_R1207_U286, P1_R1207_U181, P1_R1207_U187);
  nand ginst4240 (P1_R1207_U287, P1_R1207_U11, P1_R1207_U286);
  nand ginst4241 (P1_R1207_U288, P1_R1207_U77, P1_U4024);
  nand ginst4242 (P1_R1207_U289, P1_R1207_U75, P1_U4022);
  nand ginst4243 (P1_R1207_U29, P1_R1207_U23, P1_U3068);
  nand ginst4244 (P1_R1207_U290, P1_R1207_U127, P1_R1207_U163, P1_R1207_U283);
  nand ginst4245 (P1_R1207_U291, P1_R1207_U287, P1_R1207_U289);
  not ginst4246 (P1_R1207_U292, P1_R1207_U160);
  nand ginst4247 (P1_R1207_U293, P1_R1207_U80, P1_U4021);
  nand ginst4248 (P1_R1207_U294, P1_R1207_U160, P1_R1207_U293);
  nand ginst4249 (P1_R1207_U295, P1_R1207_U79, P1_U3065);
  not ginst4250 (P1_R1207_U296, P1_R1207_U159);
  nand ginst4251 (P1_R1207_U297, P1_R1207_U82, P1_U4020);
  nand ginst4252 (P1_R1207_U298, P1_R1207_U159, P1_R1207_U297);
  nand ginst4253 (P1_R1207_U299, P1_R1207_U81, P1_U3058);
  not ginst4254 (P1_R1207_U30, P1_U3064);
  not ginst4255 (P1_R1207_U300, P1_R1207_U89);
  nand ginst4256 (P1_R1207_U301, P1_R1207_U86, P1_U4018);
  nand ginst4257 (P1_R1207_U302, P1_R1207_U182, P1_R1207_U301, P1_R1207_U89);
  nand ginst4258 (P1_R1207_U303, P1_R1207_U85, P1_R1207_U86);
  nand ginst4259 (P1_R1207_U304, P1_R1207_U303, P1_R1207_U83);
  nand ginst4260 (P1_R1207_U305, P1_R1207_U176, P1_U3053);
  not ginst4261 (P1_R1207_U306, P1_R1207_U157);
  nand ginst4262 (P1_R1207_U307, P1_R1207_U88, P1_U4017);
  nand ginst4263 (P1_R1207_U308, P1_R1207_U87, P1_U3054);
  nand ginst4264 (P1_R1207_U309, P1_R1207_U300, P1_R1207_U85);
  not ginst4265 (P1_R1207_U31, P1_U3476);
  nand ginst4266 (P1_R1207_U310, P1_R1207_U133, P1_R1207_U309);
  nand ginst4267 (P1_R1207_U311, P1_R1207_U182, P1_R1207_U89);
  nand ginst4268 (P1_R1207_U312, P1_R1207_U132, P1_R1207_U311);
  nand ginst4269 (P1_R1207_U313, P1_R1207_U182, P1_R1207_U85);
  nand ginst4270 (P1_R1207_U314, P1_R1207_U163, P1_R1207_U288);
  not ginst4271 (P1_R1207_U315, P1_R1207_U90);
  nand ginst4272 (P1_R1207_U316, P1_R1207_U48, P1_U3061);
  nand ginst4273 (P1_R1207_U317, P1_R1207_U315, P1_R1207_U316);
  nand ginst4274 (P1_R1207_U318, P1_R1207_U136, P1_R1207_U317);
  nand ginst4275 (P1_R1207_U319, P1_R1207_U181, P1_R1207_U90);
  not ginst4276 (P1_R1207_U32, P1_U3473);
  nand ginst4277 (P1_R1207_U320, P1_R1207_U75, P1_U4022);
  nand ginst4278 (P1_R1207_U321, P1_R1207_U11, P1_R1207_U319, P1_R1207_U320);
  nand ginst4279 (P1_R1207_U322, P1_R1207_U48, P1_U3061);
  nand ginst4280 (P1_R1207_U323, P1_R1207_U181, P1_R1207_U322);
  nand ginst4281 (P1_R1207_U324, P1_R1207_U288, P1_R1207_U78);
  nand ginst4282 (P1_R1207_U325, P1_R1207_U171, P1_R1207_U262);
  not ginst4283 (P1_R1207_U326, P1_R1207_U91);
  nand ginst4284 (P1_R1207_U327, P1_R1207_U49, P1_U3074);
  nand ginst4285 (P1_R1207_U328, P1_R1207_U326, P1_R1207_U327);
  nand ginst4286 (P1_R1207_U329, P1_R1207_U142, P1_R1207_U328);
  not ginst4287 (P1_R1207_U33, P1_U3470);
  nand ginst4288 (P1_R1207_U330, P1_R1207_U180, P1_R1207_U91);
  nand ginst4289 (P1_R1207_U331, P1_R1207_U61, P1_U3506);
  nand ginst4290 (P1_R1207_U332, P1_R1207_U10, P1_R1207_U330, P1_R1207_U331);
  nand ginst4291 (P1_R1207_U333, P1_R1207_U49, P1_U3074);
  nand ginst4292 (P1_R1207_U334, P1_R1207_U180, P1_R1207_U333);
  nand ginst4293 (P1_R1207_U335, P1_R1207_U262, P1_R1207_U64);
  nand ginst4294 (P1_R1207_U336, P1_R1207_U148, P1_R1207_U217);
  not ginst4295 (P1_R1207_U337, P1_R1207_U92);
  nand ginst4296 (P1_R1207_U338, P1_R1207_U51, P1_U3062);
  nand ginst4297 (P1_R1207_U339, P1_R1207_U337, P1_R1207_U338);
  not ginst4298 (P1_R1207_U34, P1_U3071);
  nand ginst4299 (P1_R1207_U340, P1_R1207_U146, P1_R1207_U339);
  nand ginst4300 (P1_R1207_U341, P1_R1207_U179, P1_R1207_U92);
  nand ginst4301 (P1_R1207_U342, P1_R1207_U52, P1_U3491);
  nand ginst4302 (P1_R1207_U343, P1_R1207_U145, P1_R1207_U341);
  nand ginst4303 (P1_R1207_U344, P1_R1207_U51, P1_U3062);
  nand ginst4304 (P1_R1207_U345, P1_R1207_U179, P1_R1207_U344);
  nand ginst4305 (P1_R1207_U346, P1_R1207_U24, P1_U3077);
  nand ginst4306 (P1_R1207_U347, P1_R1207_U182, P1_R1207_U301, P1_R1207_U89);
  nand ginst4307 (P1_R1207_U348, P1_R1207_U12, P1_R1207_U130, P1_R1207_U347);
  nand ginst4308 (P1_R1207_U349, P1_R1207_U43, P1_U3485);
  not ginst4309 (P1_R1207_U35, P1_U3067);
  nand ginst4310 (P1_R1207_U350, P1_R1207_U42, P1_U3083);
  nand ginst4311 (P1_R1207_U351, P1_R1207_U148, P1_R1207_U218);
  nand ginst4312 (P1_R1207_U352, P1_R1207_U147, P1_R1207_U216);
  nand ginst4313 (P1_R1207_U353, P1_R1207_U41, P1_U3482);
  nand ginst4314 (P1_R1207_U354, P1_R1207_U38, P1_U3084);
  nand ginst4315 (P1_R1207_U355, P1_R1207_U41, P1_U3482);
  nand ginst4316 (P1_R1207_U356, P1_R1207_U38, P1_U3084);
  nand ginst4317 (P1_R1207_U357, P1_R1207_U355, P1_R1207_U356);
  nand ginst4318 (P1_R1207_U358, P1_R1207_U39, P1_U3479);
  nand ginst4319 (P1_R1207_U359, P1_R1207_U22, P1_U3070);
  not ginst4320 (P1_R1207_U36, P1_U3060);
  nand ginst4321 (P1_R1207_U360, P1_R1207_U223, P1_R1207_U44);
  nand ginst4322 (P1_R1207_U361, P1_R1207_U149, P1_R1207_U210);
  nand ginst4323 (P1_R1207_U362, P1_R1207_U34, P1_U3476);
  nand ginst4324 (P1_R1207_U363, P1_R1207_U31, P1_U3071);
  nand ginst4325 (P1_R1207_U364, P1_R1207_U362, P1_R1207_U363);
  nand ginst4326 (P1_R1207_U365, P1_R1207_U35, P1_U3473);
  nand ginst4327 (P1_R1207_U366, P1_R1207_U32, P1_U3067);
  nand ginst4328 (P1_R1207_U367, P1_R1207_U233, P1_R1207_U45);
  nand ginst4329 (P1_R1207_U368, P1_R1207_U150, P1_R1207_U225);
  nand ginst4330 (P1_R1207_U369, P1_R1207_U36, P1_U3470);
  nand ginst4331 (P1_R1207_U37, P1_R1207_U33, P1_U3060);
  nand ginst4332 (P1_R1207_U370, P1_R1207_U33, P1_U3060);
  nand ginst4333 (P1_R1207_U371, P1_R1207_U152, P1_R1207_U234);
  nand ginst4334 (P1_R1207_U372, P1_R1207_U151, P1_R1207_U200);
  nand ginst4335 (P1_R1207_U373, P1_R1207_U30, P1_U3467);
  nand ginst4336 (P1_R1207_U374, P1_R1207_U27, P1_U3064);
  nand ginst4337 (P1_R1207_U375, P1_R1207_U30, P1_U3467);
  nand ginst4338 (P1_R1207_U376, P1_R1207_U27, P1_U3064);
  nand ginst4339 (P1_R1207_U377, P1_R1207_U375, P1_R1207_U376);
  nand ginst4340 (P1_R1207_U378, P1_R1207_U28, P1_U3464);
  nand ginst4341 (P1_R1207_U379, P1_R1207_U23, P1_U3068);
  not ginst4342 (P1_R1207_U38, P1_U3482);
  nand ginst4343 (P1_R1207_U380, P1_R1207_U239, P1_R1207_U46);
  nand ginst4344 (P1_R1207_U381, P1_R1207_U153, P1_R1207_U194);
  nand ginst4345 (P1_R1207_U382, P1_R1207_U155, P1_U4028);
  nand ginst4346 (P1_R1207_U383, P1_R1207_U154, P1_U3055);
  nand ginst4347 (P1_R1207_U384, P1_R1207_U155, P1_U4028);
  nand ginst4348 (P1_R1207_U385, P1_R1207_U154, P1_U3055);
  nand ginst4349 (P1_R1207_U386, P1_R1207_U384, P1_R1207_U385);
  nand ginst4350 (P1_R1207_U387, P1_R1207_U386, P1_R1207_U87, P1_U3054);
  nand ginst4351 (P1_R1207_U388, P1_R1207_U12, P1_R1207_U88, P1_U4017);
  nand ginst4352 (P1_R1207_U389, P1_R1207_U88, P1_U4017);
  not ginst4353 (P1_R1207_U39, P1_U3070);
  nand ginst4354 (P1_R1207_U390, P1_R1207_U87, P1_U3054);
  not ginst4355 (P1_R1207_U391, P1_R1207_U131);
  nand ginst4356 (P1_R1207_U392, P1_R1207_U306, P1_R1207_U391);
  nand ginst4357 (P1_R1207_U393, P1_R1207_U131, P1_R1207_U157);
  nand ginst4358 (P1_R1207_U394, P1_R1207_U86, P1_U4018);
  nand ginst4359 (P1_R1207_U395, P1_R1207_U83, P1_U3053);
  nand ginst4360 (P1_R1207_U396, P1_R1207_U86, P1_U4018);
  nand ginst4361 (P1_R1207_U397, P1_R1207_U83, P1_U3053);
  nand ginst4362 (P1_R1207_U398, P1_R1207_U396, P1_R1207_U397);
  nand ginst4363 (P1_R1207_U399, P1_R1207_U84, P1_U4019);
  nand ginst4364 (P1_R1207_U40, P1_R1207_U22, P1_U3070);
  nand ginst4365 (P1_R1207_U400, P1_R1207_U47, P1_U3057);
  nand ginst4366 (P1_R1207_U401, P1_R1207_U313, P1_R1207_U89);
  nand ginst4367 (P1_R1207_U402, P1_R1207_U158, P1_R1207_U300);
  nand ginst4368 (P1_R1207_U403, P1_R1207_U82, P1_U4020);
  nand ginst4369 (P1_R1207_U404, P1_R1207_U81, P1_U3058);
  not ginst4370 (P1_R1207_U405, P1_R1207_U134);
  nand ginst4371 (P1_R1207_U406, P1_R1207_U296, P1_R1207_U405);
  nand ginst4372 (P1_R1207_U407, P1_R1207_U134, P1_R1207_U159);
  nand ginst4373 (P1_R1207_U408, P1_R1207_U80, P1_U4021);
  nand ginst4374 (P1_R1207_U409, P1_R1207_U79, P1_U3065);
  not ginst4375 (P1_R1207_U41, P1_U3084);
  not ginst4376 (P1_R1207_U410, P1_R1207_U135);
  nand ginst4377 (P1_R1207_U411, P1_R1207_U292, P1_R1207_U410);
  nand ginst4378 (P1_R1207_U412, P1_R1207_U135, P1_R1207_U160);
  nand ginst4379 (P1_R1207_U413, P1_R1207_U75, P1_U4022);
  nand ginst4380 (P1_R1207_U414, P1_R1207_U73, P1_U3066);
  nand ginst4381 (P1_R1207_U415, P1_R1207_U413, P1_R1207_U414);
  nand ginst4382 (P1_R1207_U416, P1_R1207_U76, P1_U4023);
  nand ginst4383 (P1_R1207_U417, P1_R1207_U48, P1_U3061);
  nand ginst4384 (P1_R1207_U418, P1_R1207_U323, P1_R1207_U90);
  nand ginst4385 (P1_R1207_U419, P1_R1207_U161, P1_R1207_U315);
  not ginst4386 (P1_R1207_U42, P1_U3485);
  nand ginst4387 (P1_R1207_U420, P1_R1207_U77, P1_U4024);
  nand ginst4388 (P1_R1207_U421, P1_R1207_U74, P1_U3075);
  nand ginst4389 (P1_R1207_U422, P1_R1207_U163, P1_R1207_U324);
  nand ginst4390 (P1_R1207_U423, P1_R1207_U162, P1_R1207_U282);
  nand ginst4391 (P1_R1207_U424, P1_R1207_U72, P1_U4025);
  nand ginst4392 (P1_R1207_U425, P1_R1207_U71, P1_U3076);
  not ginst4393 (P1_R1207_U426, P1_R1207_U137);
  nand ginst4394 (P1_R1207_U427, P1_R1207_U278, P1_R1207_U426);
  nand ginst4395 (P1_R1207_U428, P1_R1207_U137, P1_R1207_U164);
  nand ginst4396 (P1_R1207_U429, P1_R1207_U26, P1_U3461);
  not ginst4397 (P1_R1207_U43, P1_U3083);
  nand ginst4398 (P1_R1207_U430, P1_R1207_U165, P1_U3078);
  not ginst4399 (P1_R1207_U431, P1_R1207_U138);
  nand ginst4400 (P1_R1207_U432, P1_R1207_U190, P1_R1207_U431);
  nand ginst4401 (P1_R1207_U433, P1_R1207_U138, P1_R1207_U25);
  nand ginst4402 (P1_R1207_U434, P1_R1207_U70, P1_U3514);
  nand ginst4403 (P1_R1207_U435, P1_R1207_U69, P1_U3081);
  not ginst4404 (P1_R1207_U436, P1_R1207_U139);
  nand ginst4405 (P1_R1207_U437, P1_R1207_U274, P1_R1207_U436);
  nand ginst4406 (P1_R1207_U438, P1_R1207_U139, P1_R1207_U166);
  nand ginst4407 (P1_R1207_U439, P1_R1207_U68, P1_U3512);
  nand ginst4408 (P1_R1207_U44, P1_R1207_U208, P1_R1207_U209);
  nand ginst4409 (P1_R1207_U440, P1_R1207_U167, P1_U3082);
  not ginst4410 (P1_R1207_U441, P1_R1207_U140);
  nand ginst4411 (P1_R1207_U442, P1_R1207_U270, P1_R1207_U441);
  nand ginst4412 (P1_R1207_U443, P1_R1207_U140, P1_R1207_U67);
  nand ginst4413 (P1_R1207_U444, P1_R1207_U66, P1_U3509);
  nand ginst4414 (P1_R1207_U445, P1_R1207_U65, P1_U3069);
  not ginst4415 (P1_R1207_U446, P1_R1207_U141);
  nand ginst4416 (P1_R1207_U447, P1_R1207_U266, P1_R1207_U446);
  nand ginst4417 (P1_R1207_U448, P1_R1207_U141, P1_R1207_U168);
  nand ginst4418 (P1_R1207_U449, P1_R1207_U61, P1_U3506);
  nand ginst4419 (P1_R1207_U45, P1_R1207_U224, P1_R1207_U37);
  nand ginst4420 (P1_R1207_U450, P1_R1207_U59, P1_U3073);
  nand ginst4421 (P1_R1207_U451, P1_R1207_U449, P1_R1207_U450);
  nand ginst4422 (P1_R1207_U452, P1_R1207_U62, P1_U3503);
  nand ginst4423 (P1_R1207_U453, P1_R1207_U49, P1_U3074);
  nand ginst4424 (P1_R1207_U454, P1_R1207_U334, P1_R1207_U91);
  nand ginst4425 (P1_R1207_U455, P1_R1207_U169, P1_R1207_U326);
  nand ginst4426 (P1_R1207_U456, P1_R1207_U63, P1_U3500);
  nand ginst4427 (P1_R1207_U457, P1_R1207_U60, P1_U3079);
  nand ginst4428 (P1_R1207_U458, P1_R1207_U171, P1_R1207_U335);
  nand ginst4429 (P1_R1207_U459, P1_R1207_U170, P1_R1207_U256);
  nand ginst4430 (P1_R1207_U46, P1_R1207_U192, P1_R1207_U193);
  nand ginst4431 (P1_R1207_U460, P1_R1207_U58, P1_U3497);
  nand ginst4432 (P1_R1207_U461, P1_R1207_U57, P1_U3080);
  not ginst4433 (P1_R1207_U462, P1_R1207_U143);
  nand ginst4434 (P1_R1207_U463, P1_R1207_U252, P1_R1207_U462);
  nand ginst4435 (P1_R1207_U464, P1_R1207_U143, P1_R1207_U172);
  nand ginst4436 (P1_R1207_U465, P1_R1207_U56, P1_U3494);
  nand ginst4437 (P1_R1207_U466, P1_R1207_U55, P1_U3072);
  not ginst4438 (P1_R1207_U467, P1_R1207_U144);
  nand ginst4439 (P1_R1207_U468, P1_R1207_U248, P1_R1207_U467);
  nand ginst4440 (P1_R1207_U469, P1_R1207_U144, P1_R1207_U173);
  not ginst4441 (P1_R1207_U47, P1_U4019);
  nand ginst4442 (P1_R1207_U470, P1_R1207_U52, P1_U3491);
  nand ginst4443 (P1_R1207_U471, P1_R1207_U50, P1_U3063);
  nand ginst4444 (P1_R1207_U472, P1_R1207_U470, P1_R1207_U471);
  nand ginst4445 (P1_R1207_U473, P1_R1207_U53, P1_U3488);
  nand ginst4446 (P1_R1207_U474, P1_R1207_U51, P1_U3062);
  nand ginst4447 (P1_R1207_U475, P1_R1207_U345, P1_R1207_U92);
  nand ginst4448 (P1_R1207_U476, P1_R1207_U174, P1_R1207_U337);
  not ginst4449 (P1_R1207_U48, P1_U4023);
  not ginst4450 (P1_R1207_U49, P1_U3503);
  not ginst4451 (P1_R1207_U50, P1_U3491);
  not ginst4452 (P1_R1207_U51, P1_U3488);
  not ginst4453 (P1_R1207_U52, P1_U3063);
  not ginst4454 (P1_R1207_U53, P1_U3062);
  nand ginst4455 (P1_R1207_U54, P1_R1207_U42, P1_U3083);
  not ginst4456 (P1_R1207_U55, P1_U3494);
  not ginst4457 (P1_R1207_U56, P1_U3072);
  not ginst4458 (P1_R1207_U57, P1_U3497);
  not ginst4459 (P1_R1207_U58, P1_U3080);
  not ginst4460 (P1_R1207_U59, P1_U3506);
  and ginst4461 (P1_R1207_U6, P1_R1207_U184, P1_R1207_U201);
  not ginst4462 (P1_R1207_U60, P1_U3500);
  not ginst4463 (P1_R1207_U61, P1_U3073);
  not ginst4464 (P1_R1207_U62, P1_U3074);
  not ginst4465 (P1_R1207_U63, P1_U3079);
  nand ginst4466 (P1_R1207_U64, P1_R1207_U60, P1_U3079);
  not ginst4467 (P1_R1207_U65, P1_U3509);
  not ginst4468 (P1_R1207_U66, P1_U3069);
  nand ginst4469 (P1_R1207_U67, P1_R1207_U268, P1_R1207_U269);
  not ginst4470 (P1_R1207_U68, P1_U3082);
  not ginst4471 (P1_R1207_U69, P1_U3514);
  and ginst4472 (P1_R1207_U7, P1_R1207_U202, P1_R1207_U203);
  not ginst4473 (P1_R1207_U70, P1_U3081);
  not ginst4474 (P1_R1207_U71, P1_U4025);
  not ginst4475 (P1_R1207_U72, P1_U3076);
  not ginst4476 (P1_R1207_U73, P1_U4022);
  not ginst4477 (P1_R1207_U74, P1_U4024);
  not ginst4478 (P1_R1207_U75, P1_U3066);
  not ginst4479 (P1_R1207_U76, P1_U3061);
  not ginst4480 (P1_R1207_U77, P1_U3075);
  nand ginst4481 (P1_R1207_U78, P1_R1207_U74, P1_U3075);
  not ginst4482 (P1_R1207_U79, P1_U4021);
  and ginst4483 (P1_R1207_U8, P1_R1207_U179, P1_R1207_U240);
  not ginst4484 (P1_R1207_U80, P1_U3065);
  not ginst4485 (P1_R1207_U81, P1_U4020);
  not ginst4486 (P1_R1207_U82, P1_U3058);
  not ginst4487 (P1_R1207_U83, P1_U4018);
  not ginst4488 (P1_R1207_U84, P1_U3057);
  nand ginst4489 (P1_R1207_U85, P1_R1207_U47, P1_U3057);
  not ginst4490 (P1_R1207_U86, P1_U3053);
  not ginst4491 (P1_R1207_U87, P1_U4017);
  not ginst4492 (P1_R1207_U88, P1_U3054);
  nand ginst4493 (P1_R1207_U89, P1_R1207_U298, P1_R1207_U299);
  and ginst4494 (P1_R1207_U9, P1_R1207_U241, P1_R1207_U242);
  nand ginst4495 (P1_R1207_U90, P1_R1207_U314, P1_R1207_U78);
  nand ginst4496 (P1_R1207_U91, P1_R1207_U325, P1_R1207_U64);
  nand ginst4497 (P1_R1207_U92, P1_R1207_U336, P1_R1207_U54);
  not ginst4498 (P1_R1207_U93, P1_U3077);
  nand ginst4499 (P1_R1207_U94, P1_R1207_U392, P1_R1207_U393);
  nand ginst4500 (P1_R1207_U95, P1_R1207_U406, P1_R1207_U407);
  nand ginst4501 (P1_R1207_U96, P1_R1207_U411, P1_R1207_U412);
  nand ginst4502 (P1_R1207_U97, P1_R1207_U427, P1_R1207_U428);
  nand ginst4503 (P1_R1207_U98, P1_R1207_U432, P1_R1207_U433);
  nand ginst4504 (P1_R1207_U99, P1_R1207_U437, P1_R1207_U438);
  and ginst4505 (P1_R1222_U10, P1_R1222_U268, P1_R1222_U269);
  nand ginst4506 (P1_R1222_U100, P1_R1222_U390, P1_R1222_U391);
  nand ginst4507 (P1_R1222_U101, P1_R1222_U395, P1_R1222_U396);
  nand ginst4508 (P1_R1222_U102, P1_R1222_U404, P1_R1222_U405);
  nand ginst4509 (P1_R1222_U103, P1_R1222_U411, P1_R1222_U412);
  nand ginst4510 (P1_R1222_U104, P1_R1222_U418, P1_R1222_U419);
  nand ginst4511 (P1_R1222_U105, P1_R1222_U425, P1_R1222_U426);
  nand ginst4512 (P1_R1222_U106, P1_R1222_U430, P1_R1222_U431);
  nand ginst4513 (P1_R1222_U107, P1_R1222_U437, P1_R1222_U438);
  nand ginst4514 (P1_R1222_U108, P1_R1222_U444, P1_R1222_U445);
  nand ginst4515 (P1_R1222_U109, P1_R1222_U458, P1_R1222_U459);
  and ginst4516 (P1_R1222_U11, P1_R1222_U345, P1_R1222_U348);
  nand ginst4517 (P1_R1222_U110, P1_R1222_U463, P1_R1222_U464);
  nand ginst4518 (P1_R1222_U111, P1_R1222_U470, P1_R1222_U471);
  nand ginst4519 (P1_R1222_U112, P1_R1222_U477, P1_R1222_U478);
  nand ginst4520 (P1_R1222_U113, P1_R1222_U484, P1_R1222_U485);
  nand ginst4521 (P1_R1222_U114, P1_R1222_U491, P1_R1222_U492);
  nand ginst4522 (P1_R1222_U115, P1_R1222_U496, P1_R1222_U497);
  and ginst4523 (P1_R1222_U116, P1_U3068, P1_U3464);
  and ginst4524 (P1_R1222_U117, P1_R1222_U184, P1_R1222_U186);
  and ginst4525 (P1_R1222_U118, P1_R1222_U189, P1_R1222_U191);
  and ginst4526 (P1_R1222_U119, P1_R1222_U197, P1_R1222_U198);
  and ginst4527 (P1_R1222_U12, P1_R1222_U338, P1_R1222_U341);
  and ginst4528 (P1_R1222_U120, P1_R1222_U23, P1_R1222_U378, P1_R1222_U379);
  and ginst4529 (P1_R1222_U121, P1_R1222_U209, P1_R1222_U6);
  and ginst4530 (P1_R1222_U122, P1_R1222_U215, P1_R1222_U217);
  and ginst4531 (P1_R1222_U123, P1_R1222_U35, P1_R1222_U385, P1_R1222_U386);
  and ginst4532 (P1_R1222_U124, P1_R1222_U223, P1_R1222_U4);
  and ginst4533 (P1_R1222_U125, P1_R1222_U178, P1_R1222_U231);
  and ginst4534 (P1_R1222_U126, P1_R1222_U201, P1_R1222_U7);
  and ginst4535 (P1_R1222_U127, P1_R1222_U168, P1_R1222_U236);
  and ginst4536 (P1_R1222_U128, P1_R1222_U169, P1_R1222_U245);
  and ginst4537 (P1_R1222_U129, P1_R1222_U264, P1_R1222_U265);
  and ginst4538 (P1_R1222_U13, P1_R1222_U329, P1_R1222_U332);
  and ginst4539 (P1_R1222_U130, P1_R1222_U10, P1_R1222_U279);
  and ginst4540 (P1_R1222_U131, P1_R1222_U277, P1_R1222_U282);
  and ginst4541 (P1_R1222_U132, P1_R1222_U295, P1_R1222_U298);
  and ginst4542 (P1_R1222_U133, P1_R1222_U299, P1_R1222_U365);
  and ginst4543 (P1_R1222_U134, P1_R1222_U156, P1_R1222_U275);
  and ginst4544 (P1_R1222_U135, P1_R1222_U465, P1_R1222_U466, P1_R1222_U60);
  and ginst4545 (P1_R1222_U136, P1_R1222_U169, P1_R1222_U486, P1_R1222_U487);
  and ginst4546 (P1_R1222_U137, P1_R1222_U340, P1_R1222_U8);
  and ginst4547 (P1_R1222_U138, P1_R1222_U168, P1_R1222_U498, P1_R1222_U499);
  and ginst4548 (P1_R1222_U139, P1_R1222_U347, P1_R1222_U7);
  and ginst4549 (P1_R1222_U14, P1_R1222_U320, P1_R1222_U323);
  nand ginst4550 (P1_R1222_U140, P1_R1222_U119, P1_R1222_U199);
  nand ginst4551 (P1_R1222_U141, P1_R1222_U214, P1_R1222_U226);
  not ginst4552 (P1_R1222_U142, P1_U3055);
  not ginst4553 (P1_R1222_U143, P1_U4028);
  and ginst4554 (P1_R1222_U144, P1_R1222_U399, P1_R1222_U400);
  nand ginst4555 (P1_R1222_U145, P1_R1222_U166, P1_R1222_U301, P1_R1222_U361);
  and ginst4556 (P1_R1222_U146, P1_R1222_U406, P1_R1222_U407);
  nand ginst4557 (P1_R1222_U147, P1_R1222_U133, P1_R1222_U366, P1_R1222_U367);
  and ginst4558 (P1_R1222_U148, P1_R1222_U413, P1_R1222_U414);
  nand ginst4559 (P1_R1222_U149, P1_R1222_U296, P1_R1222_U362, P1_R1222_U87);
  and ginst4560 (P1_R1222_U15, P1_R1222_U315, P1_R1222_U317);
  and ginst4561 (P1_R1222_U150, P1_R1222_U420, P1_R1222_U421);
  nand ginst4562 (P1_R1222_U151, P1_R1222_U289, P1_R1222_U290);
  and ginst4563 (P1_R1222_U152, P1_R1222_U432, P1_R1222_U433);
  nand ginst4564 (P1_R1222_U153, P1_R1222_U285, P1_R1222_U286);
  and ginst4565 (P1_R1222_U154, P1_R1222_U439, P1_R1222_U440);
  nand ginst4566 (P1_R1222_U155, P1_R1222_U131, P1_R1222_U281);
  and ginst4567 (P1_R1222_U156, P1_R1222_U446, P1_R1222_U447);
  and ginst4568 (P1_R1222_U157, P1_R1222_U451, P1_R1222_U452);
  nand ginst4569 (P1_R1222_U158, P1_R1222_U324, P1_R1222_U44);
  nand ginst4570 (P1_R1222_U159, P1_R1222_U129, P1_R1222_U266);
  and ginst4571 (P1_R1222_U16, P1_R1222_U307, P1_R1222_U310);
  and ginst4572 (P1_R1222_U160, P1_R1222_U472, P1_R1222_U473);
  nand ginst4573 (P1_R1222_U161, P1_R1222_U253, P1_R1222_U254);
  and ginst4574 (P1_R1222_U162, P1_R1222_U479, P1_R1222_U480);
  nand ginst4575 (P1_R1222_U163, P1_R1222_U249, P1_R1222_U250);
  nand ginst4576 (P1_R1222_U164, P1_R1222_U239, P1_R1222_U240);
  nand ginst4577 (P1_R1222_U165, P1_R1222_U363, P1_R1222_U364);
  nand ginst4578 (P1_R1222_U166, P1_R1222_U147, P1_U3054);
  not ginst4579 (P1_R1222_U167, P1_R1222_U35);
  nand ginst4580 (P1_R1222_U168, P1_U3083, P1_U3485);
  nand ginst4581 (P1_R1222_U169, P1_U3072, P1_U3494);
  and ginst4582 (P1_R1222_U17, P1_R1222_U229, P1_R1222_U232);
  nand ginst4583 (P1_R1222_U170, P1_U3058, P1_U4020);
  not ginst4584 (P1_R1222_U171, P1_R1222_U69);
  not ginst4585 (P1_R1222_U172, P1_R1222_U78);
  nand ginst4586 (P1_R1222_U173, P1_U3065, P1_U4021);
  not ginst4587 (P1_R1222_U174, P1_R1222_U62);
  or ginst4588 (P1_R1222_U175, P1_U3067, P1_U3473);
  or ginst4589 (P1_R1222_U176, P1_U3060, P1_U3470);
  or ginst4590 (P1_R1222_U177, P1_U3064, P1_U3467);
  or ginst4591 (P1_R1222_U178, P1_U3068, P1_U3464);
  not ginst4592 (P1_R1222_U179, P1_R1222_U32);
  and ginst4593 (P1_R1222_U18, P1_R1222_U221, P1_R1222_U224);
  or ginst4594 (P1_R1222_U180, P1_U3078, P1_U3461);
  not ginst4595 (P1_R1222_U181, P1_R1222_U43);
  not ginst4596 (P1_R1222_U182, P1_R1222_U44);
  nand ginst4597 (P1_R1222_U183, P1_R1222_U43, P1_R1222_U44);
  nand ginst4598 (P1_R1222_U184, P1_R1222_U116, P1_R1222_U177);
  nand ginst4599 (P1_R1222_U185, P1_R1222_U183, P1_R1222_U5);
  nand ginst4600 (P1_R1222_U186, P1_U3064, P1_U3467);
  nand ginst4601 (P1_R1222_U187, P1_R1222_U117, P1_R1222_U185);
  nand ginst4602 (P1_R1222_U188, P1_R1222_U35, P1_R1222_U36);
  nand ginst4603 (P1_R1222_U189, P1_R1222_U188, P1_U3067);
  and ginst4604 (P1_R1222_U19, P1_R1222_U207, P1_R1222_U210);
  nand ginst4605 (P1_R1222_U190, P1_R1222_U187, P1_R1222_U4);
  nand ginst4606 (P1_R1222_U191, P1_R1222_U167, P1_U3473);
  not ginst4607 (P1_R1222_U192, P1_R1222_U42);
  or ginst4608 (P1_R1222_U193, P1_U3070, P1_U3479);
  or ginst4609 (P1_R1222_U194, P1_U3071, P1_U3476);
  not ginst4610 (P1_R1222_U195, P1_R1222_U23);
  nand ginst4611 (P1_R1222_U196, P1_R1222_U23, P1_R1222_U24);
  nand ginst4612 (P1_R1222_U197, P1_R1222_U196, P1_U3070);
  nand ginst4613 (P1_R1222_U198, P1_R1222_U195, P1_U3479);
  nand ginst4614 (P1_R1222_U199, P1_R1222_U42, P1_R1222_U6);
  not ginst4615 (P1_R1222_U20, P1_U3476);
  not ginst4616 (P1_R1222_U200, P1_R1222_U140);
  or ginst4617 (P1_R1222_U201, P1_U3084, P1_U3482);
  nand ginst4618 (P1_R1222_U202, P1_R1222_U140, P1_R1222_U201);
  not ginst4619 (P1_R1222_U203, P1_R1222_U41);
  or ginst4620 (P1_R1222_U204, P1_U3083, P1_U3485);
  or ginst4621 (P1_R1222_U205, P1_U3071, P1_U3476);
  nand ginst4622 (P1_R1222_U206, P1_R1222_U205, P1_R1222_U42);
  nand ginst4623 (P1_R1222_U207, P1_R1222_U120, P1_R1222_U206);
  nand ginst4624 (P1_R1222_U208, P1_R1222_U192, P1_R1222_U23);
  nand ginst4625 (P1_R1222_U209, P1_U3070, P1_U3479);
  not ginst4626 (P1_R1222_U21, P1_U3071);
  nand ginst4627 (P1_R1222_U210, P1_R1222_U121, P1_R1222_U208);
  or ginst4628 (P1_R1222_U211, P1_U3071, P1_U3476);
  nand ginst4629 (P1_R1222_U212, P1_R1222_U178, P1_R1222_U182);
  nand ginst4630 (P1_R1222_U213, P1_U3068, P1_U3464);
  not ginst4631 (P1_R1222_U214, P1_R1222_U46);
  nand ginst4632 (P1_R1222_U215, P1_R1222_U181, P1_R1222_U5);
  nand ginst4633 (P1_R1222_U216, P1_R1222_U177, P1_R1222_U46);
  nand ginst4634 (P1_R1222_U217, P1_U3064, P1_U3467);
  not ginst4635 (P1_R1222_U218, P1_R1222_U45);
  or ginst4636 (P1_R1222_U219, P1_U3060, P1_U3470);
  not ginst4637 (P1_R1222_U22, P1_U3070);
  nand ginst4638 (P1_R1222_U220, P1_R1222_U219, P1_R1222_U45);
  nand ginst4639 (P1_R1222_U221, P1_R1222_U123, P1_R1222_U220);
  nand ginst4640 (P1_R1222_U222, P1_R1222_U218, P1_R1222_U35);
  nand ginst4641 (P1_R1222_U223, P1_U3067, P1_U3473);
  nand ginst4642 (P1_R1222_U224, P1_R1222_U124, P1_R1222_U222);
  or ginst4643 (P1_R1222_U225, P1_U3060, P1_U3470);
  nand ginst4644 (P1_R1222_U226, P1_R1222_U178, P1_R1222_U181);
  not ginst4645 (P1_R1222_U227, P1_R1222_U141);
  nand ginst4646 (P1_R1222_U228, P1_U3064, P1_U3467);
  nand ginst4647 (P1_R1222_U229, P1_R1222_U397, P1_R1222_U398, P1_R1222_U43, P1_R1222_U44);
  nand ginst4648 (P1_R1222_U23, P1_U3071, P1_U3476);
  nand ginst4649 (P1_R1222_U230, P1_R1222_U43, P1_R1222_U44);
  nand ginst4650 (P1_R1222_U231, P1_U3068, P1_U3464);
  nand ginst4651 (P1_R1222_U232, P1_R1222_U125, P1_R1222_U230);
  or ginst4652 (P1_R1222_U233, P1_U3083, P1_U3485);
  or ginst4653 (P1_R1222_U234, P1_U3062, P1_U3488);
  nand ginst4654 (P1_R1222_U235, P1_R1222_U174, P1_R1222_U7);
  nand ginst4655 (P1_R1222_U236, P1_U3062, P1_U3488);
  nand ginst4656 (P1_R1222_U237, P1_R1222_U127, P1_R1222_U235);
  or ginst4657 (P1_R1222_U238, P1_U3062, P1_U3488);
  nand ginst4658 (P1_R1222_U239, P1_R1222_U126, P1_R1222_U140);
  not ginst4659 (P1_R1222_U24, P1_U3479);
  nand ginst4660 (P1_R1222_U240, P1_R1222_U237, P1_R1222_U238);
  not ginst4661 (P1_R1222_U241, P1_R1222_U164);
  or ginst4662 (P1_R1222_U242, P1_U3080, P1_U3497);
  or ginst4663 (P1_R1222_U243, P1_U3072, P1_U3494);
  nand ginst4664 (P1_R1222_U244, P1_R1222_U171, P1_R1222_U8);
  nand ginst4665 (P1_R1222_U245, P1_U3080, P1_U3497);
  nand ginst4666 (P1_R1222_U246, P1_R1222_U128, P1_R1222_U244);
  or ginst4667 (P1_R1222_U247, P1_U3063, P1_U3491);
  or ginst4668 (P1_R1222_U248, P1_U3080, P1_U3497);
  nand ginst4669 (P1_R1222_U249, P1_R1222_U164, P1_R1222_U247, P1_R1222_U8);
  not ginst4670 (P1_R1222_U25, P1_U3470);
  nand ginst4671 (P1_R1222_U250, P1_R1222_U246, P1_R1222_U248);
  not ginst4672 (P1_R1222_U251, P1_R1222_U163);
  or ginst4673 (P1_R1222_U252, P1_U3079, P1_U3500);
  nand ginst4674 (P1_R1222_U253, P1_R1222_U163, P1_R1222_U252);
  nand ginst4675 (P1_R1222_U254, P1_U3079, P1_U3500);
  not ginst4676 (P1_R1222_U255, P1_R1222_U161);
  or ginst4677 (P1_R1222_U256, P1_U3074, P1_U3503);
  nand ginst4678 (P1_R1222_U257, P1_R1222_U161, P1_R1222_U256);
  nand ginst4679 (P1_R1222_U258, P1_U3074, P1_U3503);
  not ginst4680 (P1_R1222_U259, P1_R1222_U93);
  not ginst4681 (P1_R1222_U26, P1_U3060);
  or ginst4682 (P1_R1222_U260, P1_U3069, P1_U3509);
  or ginst4683 (P1_R1222_U261, P1_U3073, P1_U3506);
  not ginst4684 (P1_R1222_U262, P1_R1222_U60);
  nand ginst4685 (P1_R1222_U263, P1_R1222_U60, P1_R1222_U61);
  nand ginst4686 (P1_R1222_U264, P1_R1222_U263, P1_U3069);
  nand ginst4687 (P1_R1222_U265, P1_R1222_U262, P1_U3509);
  nand ginst4688 (P1_R1222_U266, P1_R1222_U9, P1_R1222_U93);
  not ginst4689 (P1_R1222_U267, P1_R1222_U159);
  or ginst4690 (P1_R1222_U268, P1_U3076, P1_U4025);
  or ginst4691 (P1_R1222_U269, P1_U3081, P1_U3514);
  not ginst4692 (P1_R1222_U27, P1_U3067);
  or ginst4693 (P1_R1222_U270, P1_U3075, P1_U4024);
  not ginst4694 (P1_R1222_U271, P1_R1222_U81);
  nand ginst4695 (P1_R1222_U272, P1_R1222_U271, P1_U4025);
  nand ginst4696 (P1_R1222_U273, P1_R1222_U272, P1_R1222_U91);
  nand ginst4697 (P1_R1222_U274, P1_R1222_U81, P1_R1222_U82);
  nand ginst4698 (P1_R1222_U275, P1_R1222_U273, P1_R1222_U274);
  nand ginst4699 (P1_R1222_U276, P1_R1222_U10, P1_R1222_U172);
  nand ginst4700 (P1_R1222_U277, P1_U3075, P1_U4024);
  nand ginst4701 (P1_R1222_U278, P1_R1222_U275, P1_R1222_U276);
  or ginst4702 (P1_R1222_U279, P1_U3082, P1_U3512);
  not ginst4703 (P1_R1222_U28, P1_U3464);
  or ginst4704 (P1_R1222_U280, P1_U3075, P1_U4024);
  nand ginst4705 (P1_R1222_U281, P1_R1222_U130, P1_R1222_U159, P1_R1222_U270);
  nand ginst4706 (P1_R1222_U282, P1_R1222_U278, P1_R1222_U280);
  not ginst4707 (P1_R1222_U283, P1_R1222_U155);
  or ginst4708 (P1_R1222_U284, P1_U3061, P1_U4023);
  nand ginst4709 (P1_R1222_U285, P1_R1222_U155, P1_R1222_U284);
  nand ginst4710 (P1_R1222_U286, P1_U3061, P1_U4023);
  not ginst4711 (P1_R1222_U287, P1_R1222_U153);
  or ginst4712 (P1_R1222_U288, P1_U3066, P1_U4022);
  nand ginst4713 (P1_R1222_U289, P1_R1222_U153, P1_R1222_U288);
  not ginst4714 (P1_R1222_U29, P1_U3068);
  nand ginst4715 (P1_R1222_U290, P1_U3066, P1_U4022);
  not ginst4716 (P1_R1222_U291, P1_R1222_U151);
  or ginst4717 (P1_R1222_U292, P1_U3058, P1_U4020);
  nand ginst4718 (P1_R1222_U293, P1_R1222_U170, P1_R1222_U173);
  not ginst4719 (P1_R1222_U294, P1_R1222_U87);
  or ginst4720 (P1_R1222_U295, P1_U3065, P1_U4021);
  nand ginst4721 (P1_R1222_U296, P1_R1222_U151, P1_R1222_U165, P1_R1222_U295);
  not ginst4722 (P1_R1222_U297, P1_R1222_U149);
  or ginst4723 (P1_R1222_U298, P1_U3053, P1_U4018);
  nand ginst4724 (P1_R1222_U299, P1_U3053, P1_U4018);
  not ginst4725 (P1_R1222_U30, P1_U3456);
  not ginst4726 (P1_R1222_U300, P1_R1222_U147);
  nand ginst4727 (P1_R1222_U301, P1_R1222_U147, P1_U4017);
  not ginst4728 (P1_R1222_U302, P1_R1222_U145);
  nand ginst4729 (P1_R1222_U303, P1_R1222_U151, P1_R1222_U295);
  not ginst4730 (P1_R1222_U304, P1_R1222_U90);
  or ginst4731 (P1_R1222_U305, P1_U3058, P1_U4020);
  nand ginst4732 (P1_R1222_U306, P1_R1222_U305, P1_R1222_U90);
  nand ginst4733 (P1_R1222_U307, P1_R1222_U150, P1_R1222_U170, P1_R1222_U306);
  nand ginst4734 (P1_R1222_U308, P1_R1222_U170, P1_R1222_U304);
  nand ginst4735 (P1_R1222_U309, P1_U3057, P1_U4019);
  not ginst4736 (P1_R1222_U31, P1_U3077);
  nand ginst4737 (P1_R1222_U310, P1_R1222_U165, P1_R1222_U308, P1_R1222_U309);
  or ginst4738 (P1_R1222_U311, P1_U3058, P1_U4020);
  nand ginst4739 (P1_R1222_U312, P1_R1222_U159, P1_R1222_U279);
  not ginst4740 (P1_R1222_U313, P1_R1222_U92);
  nand ginst4741 (P1_R1222_U314, P1_R1222_U10, P1_R1222_U92);
  nand ginst4742 (P1_R1222_U315, P1_R1222_U134, P1_R1222_U314);
  nand ginst4743 (P1_R1222_U316, P1_R1222_U275, P1_R1222_U314);
  nand ginst4744 (P1_R1222_U317, P1_R1222_U316, P1_R1222_U450);
  or ginst4745 (P1_R1222_U318, P1_U3081, P1_U3514);
  nand ginst4746 (P1_R1222_U319, P1_R1222_U318, P1_R1222_U92);
  nand ginst4747 (P1_R1222_U32, P1_U3077, P1_U3456);
  nand ginst4748 (P1_R1222_U320, P1_R1222_U157, P1_R1222_U319, P1_R1222_U81);
  nand ginst4749 (P1_R1222_U321, P1_R1222_U313, P1_R1222_U81);
  nand ginst4750 (P1_R1222_U322, P1_U3076, P1_U4025);
  nand ginst4751 (P1_R1222_U323, P1_R1222_U10, P1_R1222_U321, P1_R1222_U322);
  or ginst4752 (P1_R1222_U324, P1_U3078, P1_U3461);
  not ginst4753 (P1_R1222_U325, P1_R1222_U158);
  or ginst4754 (P1_R1222_U326, P1_U3081, P1_U3514);
  or ginst4755 (P1_R1222_U327, P1_U3073, P1_U3506);
  nand ginst4756 (P1_R1222_U328, P1_R1222_U327, P1_R1222_U93);
  nand ginst4757 (P1_R1222_U329, P1_R1222_U135, P1_R1222_U328);
  not ginst4758 (P1_R1222_U33, P1_U3467);
  nand ginst4759 (P1_R1222_U330, P1_R1222_U259, P1_R1222_U60);
  nand ginst4760 (P1_R1222_U331, P1_U3069, P1_U3509);
  nand ginst4761 (P1_R1222_U332, P1_R1222_U330, P1_R1222_U331, P1_R1222_U9);
  or ginst4762 (P1_R1222_U333, P1_U3073, P1_U3506);
  nand ginst4763 (P1_R1222_U334, P1_R1222_U164, P1_R1222_U247);
  not ginst4764 (P1_R1222_U335, P1_R1222_U94);
  or ginst4765 (P1_R1222_U336, P1_U3072, P1_U3494);
  nand ginst4766 (P1_R1222_U337, P1_R1222_U336, P1_R1222_U94);
  nand ginst4767 (P1_R1222_U338, P1_R1222_U136, P1_R1222_U337);
  nand ginst4768 (P1_R1222_U339, P1_R1222_U169, P1_R1222_U335);
  not ginst4769 (P1_R1222_U34, P1_U3064);
  nand ginst4770 (P1_R1222_U340, P1_U3080, P1_U3497);
  nand ginst4771 (P1_R1222_U341, P1_R1222_U137, P1_R1222_U339);
  or ginst4772 (P1_R1222_U342, P1_U3072, P1_U3494);
  or ginst4773 (P1_R1222_U343, P1_U3083, P1_U3485);
  nand ginst4774 (P1_R1222_U344, P1_R1222_U343, P1_R1222_U41);
  nand ginst4775 (P1_R1222_U345, P1_R1222_U138, P1_R1222_U344);
  nand ginst4776 (P1_R1222_U346, P1_R1222_U168, P1_R1222_U203);
  nand ginst4777 (P1_R1222_U347, P1_U3062, P1_U3488);
  nand ginst4778 (P1_R1222_U348, P1_R1222_U139, P1_R1222_U346);
  nand ginst4779 (P1_R1222_U349, P1_R1222_U168, P1_R1222_U204);
  nand ginst4780 (P1_R1222_U35, P1_U3060, P1_U3470);
  nand ginst4781 (P1_R1222_U350, P1_R1222_U201, P1_R1222_U62);
  nand ginst4782 (P1_R1222_U351, P1_R1222_U211, P1_R1222_U23);
  nand ginst4783 (P1_R1222_U352, P1_R1222_U225, P1_R1222_U35);
  nand ginst4784 (P1_R1222_U353, P1_R1222_U177, P1_R1222_U228);
  nand ginst4785 (P1_R1222_U354, P1_R1222_U170, P1_R1222_U311);
  nand ginst4786 (P1_R1222_U355, P1_R1222_U173, P1_R1222_U295);
  nand ginst4787 (P1_R1222_U356, P1_R1222_U326, P1_R1222_U81);
  nand ginst4788 (P1_R1222_U357, P1_R1222_U279, P1_R1222_U78);
  nand ginst4789 (P1_R1222_U358, P1_R1222_U333, P1_R1222_U60);
  nand ginst4790 (P1_R1222_U359, P1_R1222_U169, P1_R1222_U342);
  not ginst4791 (P1_R1222_U36, P1_U3473);
  nand ginst4792 (P1_R1222_U360, P1_R1222_U247, P1_R1222_U69);
  nand ginst4793 (P1_R1222_U361, P1_U3054, P1_U4017);
  nand ginst4794 (P1_R1222_U362, P1_R1222_U165, P1_R1222_U293);
  nand ginst4795 (P1_R1222_U363, P1_R1222_U292, P1_U3057);
  nand ginst4796 (P1_R1222_U364, P1_R1222_U292, P1_U4019);
  nand ginst4797 (P1_R1222_U365, P1_R1222_U165, P1_R1222_U293, P1_R1222_U298);
  nand ginst4798 (P1_R1222_U366, P1_R1222_U132, P1_R1222_U151, P1_R1222_U165);
  nand ginst4799 (P1_R1222_U367, P1_R1222_U294, P1_R1222_U298);
  nand ginst4800 (P1_R1222_U368, P1_R1222_U40, P1_U3083);
  nand ginst4801 (P1_R1222_U369, P1_R1222_U39, P1_U3485);
  not ginst4802 (P1_R1222_U37, P1_U3482);
  nand ginst4803 (P1_R1222_U370, P1_R1222_U368, P1_R1222_U369);
  nand ginst4804 (P1_R1222_U371, P1_R1222_U349, P1_R1222_U41);
  nand ginst4805 (P1_R1222_U372, P1_R1222_U203, P1_R1222_U370);
  nand ginst4806 (P1_R1222_U373, P1_R1222_U37, P1_U3084);
  nand ginst4807 (P1_R1222_U374, P1_R1222_U38, P1_U3482);
  nand ginst4808 (P1_R1222_U375, P1_R1222_U373, P1_R1222_U374);
  nand ginst4809 (P1_R1222_U376, P1_R1222_U140, P1_R1222_U350);
  nand ginst4810 (P1_R1222_U377, P1_R1222_U200, P1_R1222_U375);
  nand ginst4811 (P1_R1222_U378, P1_R1222_U24, P1_U3070);
  nand ginst4812 (P1_R1222_U379, P1_R1222_U22, P1_U3479);
  not ginst4813 (P1_R1222_U38, P1_U3084);
  nand ginst4814 (P1_R1222_U380, P1_R1222_U20, P1_U3071);
  nand ginst4815 (P1_R1222_U381, P1_R1222_U21, P1_U3476);
  nand ginst4816 (P1_R1222_U382, P1_R1222_U380, P1_R1222_U381);
  nand ginst4817 (P1_R1222_U383, P1_R1222_U351, P1_R1222_U42);
  nand ginst4818 (P1_R1222_U384, P1_R1222_U192, P1_R1222_U382);
  nand ginst4819 (P1_R1222_U385, P1_R1222_U36, P1_U3067);
  nand ginst4820 (P1_R1222_U386, P1_R1222_U27, P1_U3473);
  nand ginst4821 (P1_R1222_U387, P1_R1222_U25, P1_U3060);
  nand ginst4822 (P1_R1222_U388, P1_R1222_U26, P1_U3470);
  nand ginst4823 (P1_R1222_U389, P1_R1222_U387, P1_R1222_U388);
  not ginst4824 (P1_R1222_U39, P1_U3083);
  nand ginst4825 (P1_R1222_U390, P1_R1222_U352, P1_R1222_U45);
  nand ginst4826 (P1_R1222_U391, P1_R1222_U218, P1_R1222_U389);
  nand ginst4827 (P1_R1222_U392, P1_R1222_U33, P1_U3064);
  nand ginst4828 (P1_R1222_U393, P1_R1222_U34, P1_U3467);
  nand ginst4829 (P1_R1222_U394, P1_R1222_U392, P1_R1222_U393);
  nand ginst4830 (P1_R1222_U395, P1_R1222_U141, P1_R1222_U353);
  nand ginst4831 (P1_R1222_U396, P1_R1222_U227, P1_R1222_U394);
  nand ginst4832 (P1_R1222_U397, P1_R1222_U28, P1_U3068);
  nand ginst4833 (P1_R1222_U398, P1_R1222_U29, P1_U3464);
  nand ginst4834 (P1_R1222_U399, P1_R1222_U143, P1_U3055);
  and ginst4835 (P1_R1222_U4, P1_R1222_U175, P1_R1222_U176);
  not ginst4836 (P1_R1222_U40, P1_U3485);
  nand ginst4837 (P1_R1222_U400, P1_R1222_U142, P1_U4028);
  nand ginst4838 (P1_R1222_U401, P1_R1222_U143, P1_U3055);
  nand ginst4839 (P1_R1222_U402, P1_R1222_U142, P1_U4028);
  nand ginst4840 (P1_R1222_U403, P1_R1222_U401, P1_R1222_U402);
  nand ginst4841 (P1_R1222_U404, P1_R1222_U144, P1_R1222_U145);
  nand ginst4842 (P1_R1222_U405, P1_R1222_U302, P1_R1222_U403);
  nand ginst4843 (P1_R1222_U406, P1_R1222_U89, P1_U3054);
  nand ginst4844 (P1_R1222_U407, P1_R1222_U88, P1_U4017);
  nand ginst4845 (P1_R1222_U408, P1_R1222_U89, P1_U3054);
  nand ginst4846 (P1_R1222_U409, P1_R1222_U88, P1_U4017);
  nand ginst4847 (P1_R1222_U41, P1_R1222_U202, P1_R1222_U62);
  nand ginst4848 (P1_R1222_U410, P1_R1222_U408, P1_R1222_U409);
  nand ginst4849 (P1_R1222_U411, P1_R1222_U146, P1_R1222_U147);
  nand ginst4850 (P1_R1222_U412, P1_R1222_U300, P1_R1222_U410);
  nand ginst4851 (P1_R1222_U413, P1_R1222_U47, P1_U3053);
  nand ginst4852 (P1_R1222_U414, P1_R1222_U48, P1_U4018);
  nand ginst4853 (P1_R1222_U415, P1_R1222_U47, P1_U3053);
  nand ginst4854 (P1_R1222_U416, P1_R1222_U48, P1_U4018);
  nand ginst4855 (P1_R1222_U417, P1_R1222_U415, P1_R1222_U416);
  nand ginst4856 (P1_R1222_U418, P1_R1222_U148, P1_R1222_U149);
  nand ginst4857 (P1_R1222_U419, P1_R1222_U297, P1_R1222_U417);
  nand ginst4858 (P1_R1222_U42, P1_R1222_U118, P1_R1222_U190);
  nand ginst4859 (P1_R1222_U420, P1_R1222_U50, P1_U3057);
  nand ginst4860 (P1_R1222_U421, P1_R1222_U49, P1_U4019);
  nand ginst4861 (P1_R1222_U422, P1_R1222_U51, P1_U3058);
  nand ginst4862 (P1_R1222_U423, P1_R1222_U52, P1_U4020);
  nand ginst4863 (P1_R1222_U424, P1_R1222_U422, P1_R1222_U423);
  nand ginst4864 (P1_R1222_U425, P1_R1222_U354, P1_R1222_U90);
  nand ginst4865 (P1_R1222_U426, P1_R1222_U304, P1_R1222_U424);
  nand ginst4866 (P1_R1222_U427, P1_R1222_U53, P1_U3065);
  nand ginst4867 (P1_R1222_U428, P1_R1222_U54, P1_U4021);
  nand ginst4868 (P1_R1222_U429, P1_R1222_U427, P1_R1222_U428);
  nand ginst4869 (P1_R1222_U43, P1_R1222_U179, P1_R1222_U180);
  nand ginst4870 (P1_R1222_U430, P1_R1222_U151, P1_R1222_U355);
  nand ginst4871 (P1_R1222_U431, P1_R1222_U291, P1_R1222_U429);
  nand ginst4872 (P1_R1222_U432, P1_R1222_U85, P1_U3066);
  nand ginst4873 (P1_R1222_U433, P1_R1222_U86, P1_U4022);
  nand ginst4874 (P1_R1222_U434, P1_R1222_U85, P1_U3066);
  nand ginst4875 (P1_R1222_U435, P1_R1222_U86, P1_U4022);
  nand ginst4876 (P1_R1222_U436, P1_R1222_U434, P1_R1222_U435);
  nand ginst4877 (P1_R1222_U437, P1_R1222_U152, P1_R1222_U153);
  nand ginst4878 (P1_R1222_U438, P1_R1222_U287, P1_R1222_U436);
  nand ginst4879 (P1_R1222_U439, P1_R1222_U83, P1_U3061);
  nand ginst4880 (P1_R1222_U44, P1_U3078, P1_U3461);
  nand ginst4881 (P1_R1222_U440, P1_R1222_U84, P1_U4023);
  nand ginst4882 (P1_R1222_U441, P1_R1222_U83, P1_U3061);
  nand ginst4883 (P1_R1222_U442, P1_R1222_U84, P1_U4023);
  nand ginst4884 (P1_R1222_U443, P1_R1222_U441, P1_R1222_U442);
  nand ginst4885 (P1_R1222_U444, P1_R1222_U154, P1_R1222_U155);
  nand ginst4886 (P1_R1222_U445, P1_R1222_U283, P1_R1222_U443);
  nand ginst4887 (P1_R1222_U446, P1_R1222_U55, P1_U3075);
  nand ginst4888 (P1_R1222_U447, P1_R1222_U56, P1_U4024);
  nand ginst4889 (P1_R1222_U448, P1_R1222_U55, P1_U3075);
  nand ginst4890 (P1_R1222_U449, P1_R1222_U56, P1_U4024);
  nand ginst4891 (P1_R1222_U45, P1_R1222_U122, P1_R1222_U216);
  nand ginst4892 (P1_R1222_U450, P1_R1222_U448, P1_R1222_U449);
  nand ginst4893 (P1_R1222_U451, P1_R1222_U82, P1_U3076);
  nand ginst4894 (P1_R1222_U452, P1_R1222_U91, P1_U4025);
  nand ginst4895 (P1_R1222_U453, P1_R1222_U158, P1_R1222_U179);
  nand ginst4896 (P1_R1222_U454, P1_R1222_U32, P1_R1222_U325);
  nand ginst4897 (P1_R1222_U455, P1_R1222_U79, P1_U3081);
  nand ginst4898 (P1_R1222_U456, P1_R1222_U80, P1_U3514);
  nand ginst4899 (P1_R1222_U457, P1_R1222_U455, P1_R1222_U456);
  nand ginst4900 (P1_R1222_U458, P1_R1222_U356, P1_R1222_U92);
  nand ginst4901 (P1_R1222_U459, P1_R1222_U313, P1_R1222_U457);
  nand ginst4902 (P1_R1222_U46, P1_R1222_U212, P1_R1222_U213);
  nand ginst4903 (P1_R1222_U460, P1_R1222_U76, P1_U3082);
  nand ginst4904 (P1_R1222_U461, P1_R1222_U77, P1_U3512);
  nand ginst4905 (P1_R1222_U462, P1_R1222_U460, P1_R1222_U461);
  nand ginst4906 (P1_R1222_U463, P1_R1222_U159, P1_R1222_U357);
  nand ginst4907 (P1_R1222_U464, P1_R1222_U267, P1_R1222_U462);
  nand ginst4908 (P1_R1222_U465, P1_R1222_U61, P1_U3069);
  nand ginst4909 (P1_R1222_U466, P1_R1222_U59, P1_U3509);
  nand ginst4910 (P1_R1222_U467, P1_R1222_U57, P1_U3073);
  nand ginst4911 (P1_R1222_U468, P1_R1222_U58, P1_U3506);
  nand ginst4912 (P1_R1222_U469, P1_R1222_U467, P1_R1222_U468);
  not ginst4913 (P1_R1222_U47, P1_U4018);
  nand ginst4914 (P1_R1222_U470, P1_R1222_U358, P1_R1222_U93);
  nand ginst4915 (P1_R1222_U471, P1_R1222_U259, P1_R1222_U469);
  nand ginst4916 (P1_R1222_U472, P1_R1222_U74, P1_U3074);
  nand ginst4917 (P1_R1222_U473, P1_R1222_U75, P1_U3503);
  nand ginst4918 (P1_R1222_U474, P1_R1222_U74, P1_U3074);
  nand ginst4919 (P1_R1222_U475, P1_R1222_U75, P1_U3503);
  nand ginst4920 (P1_R1222_U476, P1_R1222_U474, P1_R1222_U475);
  nand ginst4921 (P1_R1222_U477, P1_R1222_U160, P1_R1222_U161);
  nand ginst4922 (P1_R1222_U478, P1_R1222_U255, P1_R1222_U476);
  nand ginst4923 (P1_R1222_U479, P1_R1222_U72, P1_U3079);
  not ginst4924 (P1_R1222_U48, P1_U3053);
  nand ginst4925 (P1_R1222_U480, P1_R1222_U73, P1_U3500);
  nand ginst4926 (P1_R1222_U481, P1_R1222_U72, P1_U3079);
  nand ginst4927 (P1_R1222_U482, P1_R1222_U73, P1_U3500);
  nand ginst4928 (P1_R1222_U483, P1_R1222_U481, P1_R1222_U482);
  nand ginst4929 (P1_R1222_U484, P1_R1222_U162, P1_R1222_U163);
  nand ginst4930 (P1_R1222_U485, P1_R1222_U251, P1_R1222_U483);
  nand ginst4931 (P1_R1222_U486, P1_R1222_U70, P1_U3080);
  nand ginst4932 (P1_R1222_U487, P1_R1222_U71, P1_U3497);
  nand ginst4933 (P1_R1222_U488, P1_R1222_U65, P1_U3072);
  nand ginst4934 (P1_R1222_U489, P1_R1222_U66, P1_U3494);
  not ginst4935 (P1_R1222_U49, P1_U3057);
  nand ginst4936 (P1_R1222_U490, P1_R1222_U488, P1_R1222_U489);
  nand ginst4937 (P1_R1222_U491, P1_R1222_U359, P1_R1222_U94);
  nand ginst4938 (P1_R1222_U492, P1_R1222_U335, P1_R1222_U490);
  nand ginst4939 (P1_R1222_U493, P1_R1222_U67, P1_U3063);
  nand ginst4940 (P1_R1222_U494, P1_R1222_U68, P1_U3491);
  nand ginst4941 (P1_R1222_U495, P1_R1222_U493, P1_R1222_U494);
  nand ginst4942 (P1_R1222_U496, P1_R1222_U164, P1_R1222_U360);
  nand ginst4943 (P1_R1222_U497, P1_R1222_U241, P1_R1222_U495);
  nand ginst4944 (P1_R1222_U498, P1_R1222_U63, P1_U3062);
  nand ginst4945 (P1_R1222_U499, P1_R1222_U64, P1_U3488);
  and ginst4946 (P1_R1222_U5, P1_R1222_U177, P1_R1222_U178);
  not ginst4947 (P1_R1222_U50, P1_U4019);
  nand ginst4948 (P1_R1222_U500, P1_R1222_U30, P1_U3077);
  nand ginst4949 (P1_R1222_U501, P1_R1222_U31, P1_U3456);
  not ginst4950 (P1_R1222_U51, P1_U4020);
  not ginst4951 (P1_R1222_U52, P1_U3058);
  not ginst4952 (P1_R1222_U53, P1_U4021);
  not ginst4953 (P1_R1222_U54, P1_U3065);
  not ginst4954 (P1_R1222_U55, P1_U4024);
  not ginst4955 (P1_R1222_U56, P1_U3075);
  not ginst4956 (P1_R1222_U57, P1_U3506);
  not ginst4957 (P1_R1222_U58, P1_U3073);
  not ginst4958 (P1_R1222_U59, P1_U3069);
  and ginst4959 (P1_R1222_U6, P1_R1222_U193, P1_R1222_U194);
  nand ginst4960 (P1_R1222_U60, P1_U3073, P1_U3506);
  not ginst4961 (P1_R1222_U61, P1_U3509);
  nand ginst4962 (P1_R1222_U62, P1_U3084, P1_U3482);
  not ginst4963 (P1_R1222_U63, P1_U3488);
  not ginst4964 (P1_R1222_U64, P1_U3062);
  not ginst4965 (P1_R1222_U65, P1_U3494);
  not ginst4966 (P1_R1222_U66, P1_U3072);
  not ginst4967 (P1_R1222_U67, P1_U3491);
  not ginst4968 (P1_R1222_U68, P1_U3063);
  nand ginst4969 (P1_R1222_U69, P1_U3063, P1_U3491);
  and ginst4970 (P1_R1222_U7, P1_R1222_U233, P1_R1222_U234);
  not ginst4971 (P1_R1222_U70, P1_U3497);
  not ginst4972 (P1_R1222_U71, P1_U3080);
  not ginst4973 (P1_R1222_U72, P1_U3500);
  not ginst4974 (P1_R1222_U73, P1_U3079);
  not ginst4975 (P1_R1222_U74, P1_U3503);
  not ginst4976 (P1_R1222_U75, P1_U3074);
  not ginst4977 (P1_R1222_U76, P1_U3512);
  not ginst4978 (P1_R1222_U77, P1_U3082);
  nand ginst4979 (P1_R1222_U78, P1_U3082, P1_U3512);
  not ginst4980 (P1_R1222_U79, P1_U3514);
  and ginst4981 (P1_R1222_U8, P1_R1222_U242, P1_R1222_U243);
  not ginst4982 (P1_R1222_U80, P1_U3081);
  nand ginst4983 (P1_R1222_U81, P1_U3081, P1_U3514);
  not ginst4984 (P1_R1222_U82, P1_U4025);
  not ginst4985 (P1_R1222_U83, P1_U4023);
  not ginst4986 (P1_R1222_U84, P1_U3061);
  not ginst4987 (P1_R1222_U85, P1_U4022);
  not ginst4988 (P1_R1222_U86, P1_U3066);
  nand ginst4989 (P1_R1222_U87, P1_U3057, P1_U4019);
  not ginst4990 (P1_R1222_U88, P1_U3054);
  not ginst4991 (P1_R1222_U89, P1_U4017);
  and ginst4992 (P1_R1222_U9, P1_R1222_U260, P1_R1222_U261);
  nand ginst4993 (P1_R1222_U90, P1_R1222_U173, P1_R1222_U303);
  not ginst4994 (P1_R1222_U91, P1_U3076);
  nand ginst4995 (P1_R1222_U92, P1_R1222_U312, P1_R1222_U78);
  nand ginst4996 (P1_R1222_U93, P1_R1222_U257, P1_R1222_U258);
  nand ginst4997 (P1_R1222_U94, P1_R1222_U334, P1_R1222_U69);
  nand ginst4998 (P1_R1222_U95, P1_R1222_U453, P1_R1222_U454);
  nand ginst4999 (P1_R1222_U96, P1_R1222_U500, P1_R1222_U501);
  nand ginst5000 (P1_R1222_U97, P1_R1222_U371, P1_R1222_U372);
  nand ginst5001 (P1_R1222_U98, P1_R1222_U376, P1_R1222_U377);
  nand ginst5002 (P1_R1222_U99, P1_R1222_U383, P1_R1222_U384);
  and ginst5003 (P1_R1240_U10, P1_R1240_U268, P1_R1240_U269);
  nand ginst5004 (P1_R1240_U100, P1_R1240_U390, P1_R1240_U391);
  nand ginst5005 (P1_R1240_U101, P1_R1240_U395, P1_R1240_U396);
  nand ginst5006 (P1_R1240_U102, P1_R1240_U404, P1_R1240_U405);
  nand ginst5007 (P1_R1240_U103, P1_R1240_U411, P1_R1240_U412);
  nand ginst5008 (P1_R1240_U104, P1_R1240_U418, P1_R1240_U419);
  nand ginst5009 (P1_R1240_U105, P1_R1240_U425, P1_R1240_U426);
  nand ginst5010 (P1_R1240_U106, P1_R1240_U430, P1_R1240_U431);
  nand ginst5011 (P1_R1240_U107, P1_R1240_U437, P1_R1240_U438);
  nand ginst5012 (P1_R1240_U108, P1_R1240_U444, P1_R1240_U445);
  nand ginst5013 (P1_R1240_U109, P1_R1240_U458, P1_R1240_U459);
  and ginst5014 (P1_R1240_U11, P1_R1240_U345, P1_R1240_U348);
  nand ginst5015 (P1_R1240_U110, P1_R1240_U463, P1_R1240_U464);
  nand ginst5016 (P1_R1240_U111, P1_R1240_U470, P1_R1240_U471);
  nand ginst5017 (P1_R1240_U112, P1_R1240_U477, P1_R1240_U478);
  nand ginst5018 (P1_R1240_U113, P1_R1240_U484, P1_R1240_U485);
  nand ginst5019 (P1_R1240_U114, P1_R1240_U491, P1_R1240_U492);
  nand ginst5020 (P1_R1240_U115, P1_R1240_U496, P1_R1240_U497);
  and ginst5021 (P1_R1240_U116, P1_U3068, P1_U3464);
  and ginst5022 (P1_R1240_U117, P1_R1240_U184, P1_R1240_U186);
  and ginst5023 (P1_R1240_U118, P1_R1240_U189, P1_R1240_U191);
  and ginst5024 (P1_R1240_U119, P1_R1240_U197, P1_R1240_U198);
  and ginst5025 (P1_R1240_U12, P1_R1240_U338, P1_R1240_U341);
  and ginst5026 (P1_R1240_U120, P1_R1240_U23, P1_R1240_U378, P1_R1240_U379);
  and ginst5027 (P1_R1240_U121, P1_R1240_U209, P1_R1240_U6);
  and ginst5028 (P1_R1240_U122, P1_R1240_U215, P1_R1240_U217);
  and ginst5029 (P1_R1240_U123, P1_R1240_U35, P1_R1240_U385, P1_R1240_U386);
  and ginst5030 (P1_R1240_U124, P1_R1240_U223, P1_R1240_U4);
  and ginst5031 (P1_R1240_U125, P1_R1240_U178, P1_R1240_U231);
  and ginst5032 (P1_R1240_U126, P1_R1240_U201, P1_R1240_U7);
  and ginst5033 (P1_R1240_U127, P1_R1240_U168, P1_R1240_U236);
  and ginst5034 (P1_R1240_U128, P1_R1240_U169, P1_R1240_U245);
  and ginst5035 (P1_R1240_U129, P1_R1240_U264, P1_R1240_U265);
  and ginst5036 (P1_R1240_U13, P1_R1240_U329, P1_R1240_U332);
  and ginst5037 (P1_R1240_U130, P1_R1240_U10, P1_R1240_U279);
  and ginst5038 (P1_R1240_U131, P1_R1240_U277, P1_R1240_U282);
  and ginst5039 (P1_R1240_U132, P1_R1240_U295, P1_R1240_U298);
  and ginst5040 (P1_R1240_U133, P1_R1240_U299, P1_R1240_U365);
  and ginst5041 (P1_R1240_U134, P1_R1240_U156, P1_R1240_U275);
  and ginst5042 (P1_R1240_U135, P1_R1240_U465, P1_R1240_U466, P1_R1240_U60);
  and ginst5043 (P1_R1240_U136, P1_R1240_U169, P1_R1240_U486, P1_R1240_U487);
  and ginst5044 (P1_R1240_U137, P1_R1240_U340, P1_R1240_U8);
  and ginst5045 (P1_R1240_U138, P1_R1240_U168, P1_R1240_U498, P1_R1240_U499);
  and ginst5046 (P1_R1240_U139, P1_R1240_U347, P1_R1240_U7);
  and ginst5047 (P1_R1240_U14, P1_R1240_U320, P1_R1240_U323);
  nand ginst5048 (P1_R1240_U140, P1_R1240_U119, P1_R1240_U199);
  nand ginst5049 (P1_R1240_U141, P1_R1240_U214, P1_R1240_U226);
  not ginst5050 (P1_R1240_U142, P1_U3055);
  not ginst5051 (P1_R1240_U143, P1_U4028);
  and ginst5052 (P1_R1240_U144, P1_R1240_U399, P1_R1240_U400);
  nand ginst5053 (P1_R1240_U145, P1_R1240_U166, P1_R1240_U301, P1_R1240_U361);
  and ginst5054 (P1_R1240_U146, P1_R1240_U406, P1_R1240_U407);
  nand ginst5055 (P1_R1240_U147, P1_R1240_U133, P1_R1240_U366, P1_R1240_U367);
  and ginst5056 (P1_R1240_U148, P1_R1240_U413, P1_R1240_U414);
  nand ginst5057 (P1_R1240_U149, P1_R1240_U296, P1_R1240_U362, P1_R1240_U87);
  and ginst5058 (P1_R1240_U15, P1_R1240_U315, P1_R1240_U317);
  and ginst5059 (P1_R1240_U150, P1_R1240_U420, P1_R1240_U421);
  nand ginst5060 (P1_R1240_U151, P1_R1240_U289, P1_R1240_U290);
  and ginst5061 (P1_R1240_U152, P1_R1240_U432, P1_R1240_U433);
  nand ginst5062 (P1_R1240_U153, P1_R1240_U285, P1_R1240_U286);
  and ginst5063 (P1_R1240_U154, P1_R1240_U439, P1_R1240_U440);
  nand ginst5064 (P1_R1240_U155, P1_R1240_U131, P1_R1240_U281);
  and ginst5065 (P1_R1240_U156, P1_R1240_U446, P1_R1240_U447);
  and ginst5066 (P1_R1240_U157, P1_R1240_U451, P1_R1240_U452);
  nand ginst5067 (P1_R1240_U158, P1_R1240_U324, P1_R1240_U44);
  nand ginst5068 (P1_R1240_U159, P1_R1240_U129, P1_R1240_U266);
  and ginst5069 (P1_R1240_U16, P1_R1240_U307, P1_R1240_U310);
  and ginst5070 (P1_R1240_U160, P1_R1240_U472, P1_R1240_U473);
  nand ginst5071 (P1_R1240_U161, P1_R1240_U253, P1_R1240_U254);
  and ginst5072 (P1_R1240_U162, P1_R1240_U479, P1_R1240_U480);
  nand ginst5073 (P1_R1240_U163, P1_R1240_U249, P1_R1240_U250);
  nand ginst5074 (P1_R1240_U164, P1_R1240_U239, P1_R1240_U240);
  nand ginst5075 (P1_R1240_U165, P1_R1240_U363, P1_R1240_U364);
  nand ginst5076 (P1_R1240_U166, P1_R1240_U147, P1_U3054);
  not ginst5077 (P1_R1240_U167, P1_R1240_U35);
  nand ginst5078 (P1_R1240_U168, P1_U3083, P1_U3485);
  nand ginst5079 (P1_R1240_U169, P1_U3072, P1_U3494);
  and ginst5080 (P1_R1240_U17, P1_R1240_U229, P1_R1240_U232);
  nand ginst5081 (P1_R1240_U170, P1_U3058, P1_U4020);
  not ginst5082 (P1_R1240_U171, P1_R1240_U69);
  not ginst5083 (P1_R1240_U172, P1_R1240_U78);
  nand ginst5084 (P1_R1240_U173, P1_U3065, P1_U4021);
  not ginst5085 (P1_R1240_U174, P1_R1240_U62);
  or ginst5086 (P1_R1240_U175, P1_U3067, P1_U3473);
  or ginst5087 (P1_R1240_U176, P1_U3060, P1_U3470);
  or ginst5088 (P1_R1240_U177, P1_U3064, P1_U3467);
  or ginst5089 (P1_R1240_U178, P1_U3068, P1_U3464);
  not ginst5090 (P1_R1240_U179, P1_R1240_U32);
  and ginst5091 (P1_R1240_U18, P1_R1240_U221, P1_R1240_U224);
  or ginst5092 (P1_R1240_U180, P1_U3078, P1_U3461);
  not ginst5093 (P1_R1240_U181, P1_R1240_U43);
  not ginst5094 (P1_R1240_U182, P1_R1240_U44);
  nand ginst5095 (P1_R1240_U183, P1_R1240_U43, P1_R1240_U44);
  nand ginst5096 (P1_R1240_U184, P1_R1240_U116, P1_R1240_U177);
  nand ginst5097 (P1_R1240_U185, P1_R1240_U183, P1_R1240_U5);
  nand ginst5098 (P1_R1240_U186, P1_U3064, P1_U3467);
  nand ginst5099 (P1_R1240_U187, P1_R1240_U117, P1_R1240_U185);
  nand ginst5100 (P1_R1240_U188, P1_R1240_U35, P1_R1240_U36);
  nand ginst5101 (P1_R1240_U189, P1_R1240_U188, P1_U3067);
  and ginst5102 (P1_R1240_U19, P1_R1240_U207, P1_R1240_U210);
  nand ginst5103 (P1_R1240_U190, P1_R1240_U187, P1_R1240_U4);
  nand ginst5104 (P1_R1240_U191, P1_R1240_U167, P1_U3473);
  not ginst5105 (P1_R1240_U192, P1_R1240_U42);
  or ginst5106 (P1_R1240_U193, P1_U3070, P1_U3479);
  or ginst5107 (P1_R1240_U194, P1_U3071, P1_U3476);
  not ginst5108 (P1_R1240_U195, P1_R1240_U23);
  nand ginst5109 (P1_R1240_U196, P1_R1240_U23, P1_R1240_U24);
  nand ginst5110 (P1_R1240_U197, P1_R1240_U196, P1_U3070);
  nand ginst5111 (P1_R1240_U198, P1_R1240_U195, P1_U3479);
  nand ginst5112 (P1_R1240_U199, P1_R1240_U42, P1_R1240_U6);
  not ginst5113 (P1_R1240_U20, P1_U3476);
  not ginst5114 (P1_R1240_U200, P1_R1240_U140);
  or ginst5115 (P1_R1240_U201, P1_U3084, P1_U3482);
  nand ginst5116 (P1_R1240_U202, P1_R1240_U140, P1_R1240_U201);
  not ginst5117 (P1_R1240_U203, P1_R1240_U41);
  or ginst5118 (P1_R1240_U204, P1_U3083, P1_U3485);
  or ginst5119 (P1_R1240_U205, P1_U3071, P1_U3476);
  nand ginst5120 (P1_R1240_U206, P1_R1240_U205, P1_R1240_U42);
  nand ginst5121 (P1_R1240_U207, P1_R1240_U120, P1_R1240_U206);
  nand ginst5122 (P1_R1240_U208, P1_R1240_U192, P1_R1240_U23);
  nand ginst5123 (P1_R1240_U209, P1_U3070, P1_U3479);
  not ginst5124 (P1_R1240_U21, P1_U3071);
  nand ginst5125 (P1_R1240_U210, P1_R1240_U121, P1_R1240_U208);
  or ginst5126 (P1_R1240_U211, P1_U3071, P1_U3476);
  nand ginst5127 (P1_R1240_U212, P1_R1240_U178, P1_R1240_U182);
  nand ginst5128 (P1_R1240_U213, P1_U3068, P1_U3464);
  not ginst5129 (P1_R1240_U214, P1_R1240_U46);
  nand ginst5130 (P1_R1240_U215, P1_R1240_U181, P1_R1240_U5);
  nand ginst5131 (P1_R1240_U216, P1_R1240_U177, P1_R1240_U46);
  nand ginst5132 (P1_R1240_U217, P1_U3064, P1_U3467);
  not ginst5133 (P1_R1240_U218, P1_R1240_U45);
  or ginst5134 (P1_R1240_U219, P1_U3060, P1_U3470);
  not ginst5135 (P1_R1240_U22, P1_U3070);
  nand ginst5136 (P1_R1240_U220, P1_R1240_U219, P1_R1240_U45);
  nand ginst5137 (P1_R1240_U221, P1_R1240_U123, P1_R1240_U220);
  nand ginst5138 (P1_R1240_U222, P1_R1240_U218, P1_R1240_U35);
  nand ginst5139 (P1_R1240_U223, P1_U3067, P1_U3473);
  nand ginst5140 (P1_R1240_U224, P1_R1240_U124, P1_R1240_U222);
  or ginst5141 (P1_R1240_U225, P1_U3060, P1_U3470);
  nand ginst5142 (P1_R1240_U226, P1_R1240_U178, P1_R1240_U181);
  not ginst5143 (P1_R1240_U227, P1_R1240_U141);
  nand ginst5144 (P1_R1240_U228, P1_U3064, P1_U3467);
  nand ginst5145 (P1_R1240_U229, P1_R1240_U397, P1_R1240_U398, P1_R1240_U43, P1_R1240_U44);
  nand ginst5146 (P1_R1240_U23, P1_U3071, P1_U3476);
  nand ginst5147 (P1_R1240_U230, P1_R1240_U43, P1_R1240_U44);
  nand ginst5148 (P1_R1240_U231, P1_U3068, P1_U3464);
  nand ginst5149 (P1_R1240_U232, P1_R1240_U125, P1_R1240_U230);
  or ginst5150 (P1_R1240_U233, P1_U3083, P1_U3485);
  or ginst5151 (P1_R1240_U234, P1_U3062, P1_U3488);
  nand ginst5152 (P1_R1240_U235, P1_R1240_U174, P1_R1240_U7);
  nand ginst5153 (P1_R1240_U236, P1_U3062, P1_U3488);
  nand ginst5154 (P1_R1240_U237, P1_R1240_U127, P1_R1240_U235);
  or ginst5155 (P1_R1240_U238, P1_U3062, P1_U3488);
  nand ginst5156 (P1_R1240_U239, P1_R1240_U126, P1_R1240_U140);
  not ginst5157 (P1_R1240_U24, P1_U3479);
  nand ginst5158 (P1_R1240_U240, P1_R1240_U237, P1_R1240_U238);
  not ginst5159 (P1_R1240_U241, P1_R1240_U164);
  or ginst5160 (P1_R1240_U242, P1_U3080, P1_U3497);
  or ginst5161 (P1_R1240_U243, P1_U3072, P1_U3494);
  nand ginst5162 (P1_R1240_U244, P1_R1240_U171, P1_R1240_U8);
  nand ginst5163 (P1_R1240_U245, P1_U3080, P1_U3497);
  nand ginst5164 (P1_R1240_U246, P1_R1240_U128, P1_R1240_U244);
  or ginst5165 (P1_R1240_U247, P1_U3063, P1_U3491);
  or ginst5166 (P1_R1240_U248, P1_U3080, P1_U3497);
  nand ginst5167 (P1_R1240_U249, P1_R1240_U164, P1_R1240_U247, P1_R1240_U8);
  not ginst5168 (P1_R1240_U25, P1_U3470);
  nand ginst5169 (P1_R1240_U250, P1_R1240_U246, P1_R1240_U248);
  not ginst5170 (P1_R1240_U251, P1_R1240_U163);
  or ginst5171 (P1_R1240_U252, P1_U3079, P1_U3500);
  nand ginst5172 (P1_R1240_U253, P1_R1240_U163, P1_R1240_U252);
  nand ginst5173 (P1_R1240_U254, P1_U3079, P1_U3500);
  not ginst5174 (P1_R1240_U255, P1_R1240_U161);
  or ginst5175 (P1_R1240_U256, P1_U3074, P1_U3503);
  nand ginst5176 (P1_R1240_U257, P1_R1240_U161, P1_R1240_U256);
  nand ginst5177 (P1_R1240_U258, P1_U3074, P1_U3503);
  not ginst5178 (P1_R1240_U259, P1_R1240_U93);
  not ginst5179 (P1_R1240_U26, P1_U3060);
  or ginst5180 (P1_R1240_U260, P1_U3069, P1_U3509);
  or ginst5181 (P1_R1240_U261, P1_U3073, P1_U3506);
  not ginst5182 (P1_R1240_U262, P1_R1240_U60);
  nand ginst5183 (P1_R1240_U263, P1_R1240_U60, P1_R1240_U61);
  nand ginst5184 (P1_R1240_U264, P1_R1240_U263, P1_U3069);
  nand ginst5185 (P1_R1240_U265, P1_R1240_U262, P1_U3509);
  nand ginst5186 (P1_R1240_U266, P1_R1240_U9, P1_R1240_U93);
  not ginst5187 (P1_R1240_U267, P1_R1240_U159);
  or ginst5188 (P1_R1240_U268, P1_U3076, P1_U4025);
  or ginst5189 (P1_R1240_U269, P1_U3081, P1_U3514);
  not ginst5190 (P1_R1240_U27, P1_U3067);
  or ginst5191 (P1_R1240_U270, P1_U3075, P1_U4024);
  not ginst5192 (P1_R1240_U271, P1_R1240_U81);
  nand ginst5193 (P1_R1240_U272, P1_R1240_U271, P1_U4025);
  nand ginst5194 (P1_R1240_U273, P1_R1240_U272, P1_R1240_U91);
  nand ginst5195 (P1_R1240_U274, P1_R1240_U81, P1_R1240_U82);
  nand ginst5196 (P1_R1240_U275, P1_R1240_U273, P1_R1240_U274);
  nand ginst5197 (P1_R1240_U276, P1_R1240_U10, P1_R1240_U172);
  nand ginst5198 (P1_R1240_U277, P1_U3075, P1_U4024);
  nand ginst5199 (P1_R1240_U278, P1_R1240_U275, P1_R1240_U276);
  or ginst5200 (P1_R1240_U279, P1_U3082, P1_U3512);
  not ginst5201 (P1_R1240_U28, P1_U3464);
  or ginst5202 (P1_R1240_U280, P1_U3075, P1_U4024);
  nand ginst5203 (P1_R1240_U281, P1_R1240_U130, P1_R1240_U159, P1_R1240_U270);
  nand ginst5204 (P1_R1240_U282, P1_R1240_U278, P1_R1240_U280);
  not ginst5205 (P1_R1240_U283, P1_R1240_U155);
  or ginst5206 (P1_R1240_U284, P1_U3061, P1_U4023);
  nand ginst5207 (P1_R1240_U285, P1_R1240_U155, P1_R1240_U284);
  nand ginst5208 (P1_R1240_U286, P1_U3061, P1_U4023);
  not ginst5209 (P1_R1240_U287, P1_R1240_U153);
  or ginst5210 (P1_R1240_U288, P1_U3066, P1_U4022);
  nand ginst5211 (P1_R1240_U289, P1_R1240_U153, P1_R1240_U288);
  not ginst5212 (P1_R1240_U29, P1_U3068);
  nand ginst5213 (P1_R1240_U290, P1_U3066, P1_U4022);
  not ginst5214 (P1_R1240_U291, P1_R1240_U151);
  or ginst5215 (P1_R1240_U292, P1_U3058, P1_U4020);
  nand ginst5216 (P1_R1240_U293, P1_R1240_U170, P1_R1240_U173);
  not ginst5217 (P1_R1240_U294, P1_R1240_U87);
  or ginst5218 (P1_R1240_U295, P1_U3065, P1_U4021);
  nand ginst5219 (P1_R1240_U296, P1_R1240_U151, P1_R1240_U165, P1_R1240_U295);
  not ginst5220 (P1_R1240_U297, P1_R1240_U149);
  or ginst5221 (P1_R1240_U298, P1_U3053, P1_U4018);
  nand ginst5222 (P1_R1240_U299, P1_U3053, P1_U4018);
  not ginst5223 (P1_R1240_U30, P1_U3456);
  not ginst5224 (P1_R1240_U300, P1_R1240_U147);
  nand ginst5225 (P1_R1240_U301, P1_R1240_U147, P1_U4017);
  not ginst5226 (P1_R1240_U302, P1_R1240_U145);
  nand ginst5227 (P1_R1240_U303, P1_R1240_U151, P1_R1240_U295);
  not ginst5228 (P1_R1240_U304, P1_R1240_U90);
  or ginst5229 (P1_R1240_U305, P1_U3058, P1_U4020);
  nand ginst5230 (P1_R1240_U306, P1_R1240_U305, P1_R1240_U90);
  nand ginst5231 (P1_R1240_U307, P1_R1240_U150, P1_R1240_U170, P1_R1240_U306);
  nand ginst5232 (P1_R1240_U308, P1_R1240_U170, P1_R1240_U304);
  nand ginst5233 (P1_R1240_U309, P1_U3057, P1_U4019);
  not ginst5234 (P1_R1240_U31, P1_U3077);
  nand ginst5235 (P1_R1240_U310, P1_R1240_U165, P1_R1240_U308, P1_R1240_U309);
  or ginst5236 (P1_R1240_U311, P1_U3058, P1_U4020);
  nand ginst5237 (P1_R1240_U312, P1_R1240_U159, P1_R1240_U279);
  not ginst5238 (P1_R1240_U313, P1_R1240_U92);
  nand ginst5239 (P1_R1240_U314, P1_R1240_U10, P1_R1240_U92);
  nand ginst5240 (P1_R1240_U315, P1_R1240_U134, P1_R1240_U314);
  nand ginst5241 (P1_R1240_U316, P1_R1240_U275, P1_R1240_U314);
  nand ginst5242 (P1_R1240_U317, P1_R1240_U316, P1_R1240_U450);
  or ginst5243 (P1_R1240_U318, P1_U3081, P1_U3514);
  nand ginst5244 (P1_R1240_U319, P1_R1240_U318, P1_R1240_U92);
  nand ginst5245 (P1_R1240_U32, P1_U3077, P1_U3456);
  nand ginst5246 (P1_R1240_U320, P1_R1240_U157, P1_R1240_U319, P1_R1240_U81);
  nand ginst5247 (P1_R1240_U321, P1_R1240_U313, P1_R1240_U81);
  nand ginst5248 (P1_R1240_U322, P1_U3076, P1_U4025);
  nand ginst5249 (P1_R1240_U323, P1_R1240_U10, P1_R1240_U321, P1_R1240_U322);
  or ginst5250 (P1_R1240_U324, P1_U3078, P1_U3461);
  not ginst5251 (P1_R1240_U325, P1_R1240_U158);
  or ginst5252 (P1_R1240_U326, P1_U3081, P1_U3514);
  or ginst5253 (P1_R1240_U327, P1_U3073, P1_U3506);
  nand ginst5254 (P1_R1240_U328, P1_R1240_U327, P1_R1240_U93);
  nand ginst5255 (P1_R1240_U329, P1_R1240_U135, P1_R1240_U328);
  not ginst5256 (P1_R1240_U33, P1_U3467);
  nand ginst5257 (P1_R1240_U330, P1_R1240_U259, P1_R1240_U60);
  nand ginst5258 (P1_R1240_U331, P1_U3069, P1_U3509);
  nand ginst5259 (P1_R1240_U332, P1_R1240_U330, P1_R1240_U331, P1_R1240_U9);
  or ginst5260 (P1_R1240_U333, P1_U3073, P1_U3506);
  nand ginst5261 (P1_R1240_U334, P1_R1240_U164, P1_R1240_U247);
  not ginst5262 (P1_R1240_U335, P1_R1240_U94);
  or ginst5263 (P1_R1240_U336, P1_U3072, P1_U3494);
  nand ginst5264 (P1_R1240_U337, P1_R1240_U336, P1_R1240_U94);
  nand ginst5265 (P1_R1240_U338, P1_R1240_U136, P1_R1240_U337);
  nand ginst5266 (P1_R1240_U339, P1_R1240_U169, P1_R1240_U335);
  not ginst5267 (P1_R1240_U34, P1_U3064);
  nand ginst5268 (P1_R1240_U340, P1_U3080, P1_U3497);
  nand ginst5269 (P1_R1240_U341, P1_R1240_U137, P1_R1240_U339);
  or ginst5270 (P1_R1240_U342, P1_U3072, P1_U3494);
  or ginst5271 (P1_R1240_U343, P1_U3083, P1_U3485);
  nand ginst5272 (P1_R1240_U344, P1_R1240_U343, P1_R1240_U41);
  nand ginst5273 (P1_R1240_U345, P1_R1240_U138, P1_R1240_U344);
  nand ginst5274 (P1_R1240_U346, P1_R1240_U168, P1_R1240_U203);
  nand ginst5275 (P1_R1240_U347, P1_U3062, P1_U3488);
  nand ginst5276 (P1_R1240_U348, P1_R1240_U139, P1_R1240_U346);
  nand ginst5277 (P1_R1240_U349, P1_R1240_U168, P1_R1240_U204);
  nand ginst5278 (P1_R1240_U35, P1_U3060, P1_U3470);
  nand ginst5279 (P1_R1240_U350, P1_R1240_U201, P1_R1240_U62);
  nand ginst5280 (P1_R1240_U351, P1_R1240_U211, P1_R1240_U23);
  nand ginst5281 (P1_R1240_U352, P1_R1240_U225, P1_R1240_U35);
  nand ginst5282 (P1_R1240_U353, P1_R1240_U177, P1_R1240_U228);
  nand ginst5283 (P1_R1240_U354, P1_R1240_U170, P1_R1240_U311);
  nand ginst5284 (P1_R1240_U355, P1_R1240_U173, P1_R1240_U295);
  nand ginst5285 (P1_R1240_U356, P1_R1240_U326, P1_R1240_U81);
  nand ginst5286 (P1_R1240_U357, P1_R1240_U279, P1_R1240_U78);
  nand ginst5287 (P1_R1240_U358, P1_R1240_U333, P1_R1240_U60);
  nand ginst5288 (P1_R1240_U359, P1_R1240_U169, P1_R1240_U342);
  not ginst5289 (P1_R1240_U36, P1_U3473);
  nand ginst5290 (P1_R1240_U360, P1_R1240_U247, P1_R1240_U69);
  nand ginst5291 (P1_R1240_U361, P1_U3054, P1_U4017);
  nand ginst5292 (P1_R1240_U362, P1_R1240_U165, P1_R1240_U293);
  nand ginst5293 (P1_R1240_U363, P1_R1240_U292, P1_U3057);
  nand ginst5294 (P1_R1240_U364, P1_R1240_U292, P1_U4019);
  nand ginst5295 (P1_R1240_U365, P1_R1240_U165, P1_R1240_U293, P1_R1240_U298);
  nand ginst5296 (P1_R1240_U366, P1_R1240_U132, P1_R1240_U151, P1_R1240_U165);
  nand ginst5297 (P1_R1240_U367, P1_R1240_U294, P1_R1240_U298);
  nand ginst5298 (P1_R1240_U368, P1_R1240_U40, P1_U3083);
  nand ginst5299 (P1_R1240_U369, P1_R1240_U39, P1_U3485);
  not ginst5300 (P1_R1240_U37, P1_U3482);
  nand ginst5301 (P1_R1240_U370, P1_R1240_U368, P1_R1240_U369);
  nand ginst5302 (P1_R1240_U371, P1_R1240_U349, P1_R1240_U41);
  nand ginst5303 (P1_R1240_U372, P1_R1240_U203, P1_R1240_U370);
  nand ginst5304 (P1_R1240_U373, P1_R1240_U37, P1_U3084);
  nand ginst5305 (P1_R1240_U374, P1_R1240_U38, P1_U3482);
  nand ginst5306 (P1_R1240_U375, P1_R1240_U373, P1_R1240_U374);
  nand ginst5307 (P1_R1240_U376, P1_R1240_U140, P1_R1240_U350);
  nand ginst5308 (P1_R1240_U377, P1_R1240_U200, P1_R1240_U375);
  nand ginst5309 (P1_R1240_U378, P1_R1240_U24, P1_U3070);
  nand ginst5310 (P1_R1240_U379, P1_R1240_U22, P1_U3479);
  not ginst5311 (P1_R1240_U38, P1_U3084);
  nand ginst5312 (P1_R1240_U380, P1_R1240_U20, P1_U3071);
  nand ginst5313 (P1_R1240_U381, P1_R1240_U21, P1_U3476);
  nand ginst5314 (P1_R1240_U382, P1_R1240_U380, P1_R1240_U381);
  nand ginst5315 (P1_R1240_U383, P1_R1240_U351, P1_R1240_U42);
  nand ginst5316 (P1_R1240_U384, P1_R1240_U192, P1_R1240_U382);
  nand ginst5317 (P1_R1240_U385, P1_R1240_U36, P1_U3067);
  nand ginst5318 (P1_R1240_U386, P1_R1240_U27, P1_U3473);
  nand ginst5319 (P1_R1240_U387, P1_R1240_U25, P1_U3060);
  nand ginst5320 (P1_R1240_U388, P1_R1240_U26, P1_U3470);
  nand ginst5321 (P1_R1240_U389, P1_R1240_U387, P1_R1240_U388);
  not ginst5322 (P1_R1240_U39, P1_U3083);
  nand ginst5323 (P1_R1240_U390, P1_R1240_U352, P1_R1240_U45);
  nand ginst5324 (P1_R1240_U391, P1_R1240_U218, P1_R1240_U389);
  nand ginst5325 (P1_R1240_U392, P1_R1240_U33, P1_U3064);
  nand ginst5326 (P1_R1240_U393, P1_R1240_U34, P1_U3467);
  nand ginst5327 (P1_R1240_U394, P1_R1240_U392, P1_R1240_U393);
  nand ginst5328 (P1_R1240_U395, P1_R1240_U141, P1_R1240_U353);
  nand ginst5329 (P1_R1240_U396, P1_R1240_U227, P1_R1240_U394);
  nand ginst5330 (P1_R1240_U397, P1_R1240_U28, P1_U3068);
  nand ginst5331 (P1_R1240_U398, P1_R1240_U29, P1_U3464);
  nand ginst5332 (P1_R1240_U399, P1_R1240_U143, P1_U3055);
  and ginst5333 (P1_R1240_U4, P1_R1240_U175, P1_R1240_U176);
  not ginst5334 (P1_R1240_U40, P1_U3485);
  nand ginst5335 (P1_R1240_U400, P1_R1240_U142, P1_U4028);
  nand ginst5336 (P1_R1240_U401, P1_R1240_U143, P1_U3055);
  nand ginst5337 (P1_R1240_U402, P1_R1240_U142, P1_U4028);
  nand ginst5338 (P1_R1240_U403, P1_R1240_U401, P1_R1240_U402);
  nand ginst5339 (P1_R1240_U404, P1_R1240_U144, P1_R1240_U145);
  nand ginst5340 (P1_R1240_U405, P1_R1240_U302, P1_R1240_U403);
  nand ginst5341 (P1_R1240_U406, P1_R1240_U89, P1_U3054);
  nand ginst5342 (P1_R1240_U407, P1_R1240_U88, P1_U4017);
  nand ginst5343 (P1_R1240_U408, P1_R1240_U89, P1_U3054);
  nand ginst5344 (P1_R1240_U409, P1_R1240_U88, P1_U4017);
  nand ginst5345 (P1_R1240_U41, P1_R1240_U202, P1_R1240_U62);
  nand ginst5346 (P1_R1240_U410, P1_R1240_U408, P1_R1240_U409);
  nand ginst5347 (P1_R1240_U411, P1_R1240_U146, P1_R1240_U147);
  nand ginst5348 (P1_R1240_U412, P1_R1240_U300, P1_R1240_U410);
  nand ginst5349 (P1_R1240_U413, P1_R1240_U47, P1_U3053);
  nand ginst5350 (P1_R1240_U414, P1_R1240_U48, P1_U4018);
  nand ginst5351 (P1_R1240_U415, P1_R1240_U47, P1_U3053);
  nand ginst5352 (P1_R1240_U416, P1_R1240_U48, P1_U4018);
  nand ginst5353 (P1_R1240_U417, P1_R1240_U415, P1_R1240_U416);
  nand ginst5354 (P1_R1240_U418, P1_R1240_U148, P1_R1240_U149);
  nand ginst5355 (P1_R1240_U419, P1_R1240_U297, P1_R1240_U417);
  nand ginst5356 (P1_R1240_U42, P1_R1240_U118, P1_R1240_U190);
  nand ginst5357 (P1_R1240_U420, P1_R1240_U50, P1_U3057);
  nand ginst5358 (P1_R1240_U421, P1_R1240_U49, P1_U4019);
  nand ginst5359 (P1_R1240_U422, P1_R1240_U51, P1_U3058);
  nand ginst5360 (P1_R1240_U423, P1_R1240_U52, P1_U4020);
  nand ginst5361 (P1_R1240_U424, P1_R1240_U422, P1_R1240_U423);
  nand ginst5362 (P1_R1240_U425, P1_R1240_U354, P1_R1240_U90);
  nand ginst5363 (P1_R1240_U426, P1_R1240_U304, P1_R1240_U424);
  nand ginst5364 (P1_R1240_U427, P1_R1240_U53, P1_U3065);
  nand ginst5365 (P1_R1240_U428, P1_R1240_U54, P1_U4021);
  nand ginst5366 (P1_R1240_U429, P1_R1240_U427, P1_R1240_U428);
  nand ginst5367 (P1_R1240_U43, P1_R1240_U179, P1_R1240_U180);
  nand ginst5368 (P1_R1240_U430, P1_R1240_U151, P1_R1240_U355);
  nand ginst5369 (P1_R1240_U431, P1_R1240_U291, P1_R1240_U429);
  nand ginst5370 (P1_R1240_U432, P1_R1240_U85, P1_U3066);
  nand ginst5371 (P1_R1240_U433, P1_R1240_U86, P1_U4022);
  nand ginst5372 (P1_R1240_U434, P1_R1240_U85, P1_U3066);
  nand ginst5373 (P1_R1240_U435, P1_R1240_U86, P1_U4022);
  nand ginst5374 (P1_R1240_U436, P1_R1240_U434, P1_R1240_U435);
  nand ginst5375 (P1_R1240_U437, P1_R1240_U152, P1_R1240_U153);
  nand ginst5376 (P1_R1240_U438, P1_R1240_U287, P1_R1240_U436);
  nand ginst5377 (P1_R1240_U439, P1_R1240_U83, P1_U3061);
  nand ginst5378 (P1_R1240_U44, P1_U3078, P1_U3461);
  nand ginst5379 (P1_R1240_U440, P1_R1240_U84, P1_U4023);
  nand ginst5380 (P1_R1240_U441, P1_R1240_U83, P1_U3061);
  nand ginst5381 (P1_R1240_U442, P1_R1240_U84, P1_U4023);
  nand ginst5382 (P1_R1240_U443, P1_R1240_U441, P1_R1240_U442);
  nand ginst5383 (P1_R1240_U444, P1_R1240_U154, P1_R1240_U155);
  nand ginst5384 (P1_R1240_U445, P1_R1240_U283, P1_R1240_U443);
  nand ginst5385 (P1_R1240_U446, P1_R1240_U55, P1_U3075);
  nand ginst5386 (P1_R1240_U447, P1_R1240_U56, P1_U4024);
  nand ginst5387 (P1_R1240_U448, P1_R1240_U55, P1_U3075);
  nand ginst5388 (P1_R1240_U449, P1_R1240_U56, P1_U4024);
  nand ginst5389 (P1_R1240_U45, P1_R1240_U122, P1_R1240_U216);
  nand ginst5390 (P1_R1240_U450, P1_R1240_U448, P1_R1240_U449);
  nand ginst5391 (P1_R1240_U451, P1_R1240_U82, P1_U3076);
  nand ginst5392 (P1_R1240_U452, P1_R1240_U91, P1_U4025);
  nand ginst5393 (P1_R1240_U453, P1_R1240_U158, P1_R1240_U179);
  nand ginst5394 (P1_R1240_U454, P1_R1240_U32, P1_R1240_U325);
  nand ginst5395 (P1_R1240_U455, P1_R1240_U79, P1_U3081);
  nand ginst5396 (P1_R1240_U456, P1_R1240_U80, P1_U3514);
  nand ginst5397 (P1_R1240_U457, P1_R1240_U455, P1_R1240_U456);
  nand ginst5398 (P1_R1240_U458, P1_R1240_U356, P1_R1240_U92);
  nand ginst5399 (P1_R1240_U459, P1_R1240_U313, P1_R1240_U457);
  nand ginst5400 (P1_R1240_U46, P1_R1240_U212, P1_R1240_U213);
  nand ginst5401 (P1_R1240_U460, P1_R1240_U76, P1_U3082);
  nand ginst5402 (P1_R1240_U461, P1_R1240_U77, P1_U3512);
  nand ginst5403 (P1_R1240_U462, P1_R1240_U460, P1_R1240_U461);
  nand ginst5404 (P1_R1240_U463, P1_R1240_U159, P1_R1240_U357);
  nand ginst5405 (P1_R1240_U464, P1_R1240_U267, P1_R1240_U462);
  nand ginst5406 (P1_R1240_U465, P1_R1240_U61, P1_U3069);
  nand ginst5407 (P1_R1240_U466, P1_R1240_U59, P1_U3509);
  nand ginst5408 (P1_R1240_U467, P1_R1240_U57, P1_U3073);
  nand ginst5409 (P1_R1240_U468, P1_R1240_U58, P1_U3506);
  nand ginst5410 (P1_R1240_U469, P1_R1240_U467, P1_R1240_U468);
  not ginst5411 (P1_R1240_U47, P1_U4018);
  nand ginst5412 (P1_R1240_U470, P1_R1240_U358, P1_R1240_U93);
  nand ginst5413 (P1_R1240_U471, P1_R1240_U259, P1_R1240_U469);
  nand ginst5414 (P1_R1240_U472, P1_R1240_U74, P1_U3074);
  nand ginst5415 (P1_R1240_U473, P1_R1240_U75, P1_U3503);
  nand ginst5416 (P1_R1240_U474, P1_R1240_U74, P1_U3074);
  nand ginst5417 (P1_R1240_U475, P1_R1240_U75, P1_U3503);
  nand ginst5418 (P1_R1240_U476, P1_R1240_U474, P1_R1240_U475);
  nand ginst5419 (P1_R1240_U477, P1_R1240_U160, P1_R1240_U161);
  nand ginst5420 (P1_R1240_U478, P1_R1240_U255, P1_R1240_U476);
  nand ginst5421 (P1_R1240_U479, P1_R1240_U72, P1_U3079);
  not ginst5422 (P1_R1240_U48, P1_U3053);
  nand ginst5423 (P1_R1240_U480, P1_R1240_U73, P1_U3500);
  nand ginst5424 (P1_R1240_U481, P1_R1240_U72, P1_U3079);
  nand ginst5425 (P1_R1240_U482, P1_R1240_U73, P1_U3500);
  nand ginst5426 (P1_R1240_U483, P1_R1240_U481, P1_R1240_U482);
  nand ginst5427 (P1_R1240_U484, P1_R1240_U162, P1_R1240_U163);
  nand ginst5428 (P1_R1240_U485, P1_R1240_U251, P1_R1240_U483);
  nand ginst5429 (P1_R1240_U486, P1_R1240_U70, P1_U3080);
  nand ginst5430 (P1_R1240_U487, P1_R1240_U71, P1_U3497);
  nand ginst5431 (P1_R1240_U488, P1_R1240_U65, P1_U3072);
  nand ginst5432 (P1_R1240_U489, P1_R1240_U66, P1_U3494);
  not ginst5433 (P1_R1240_U49, P1_U3057);
  nand ginst5434 (P1_R1240_U490, P1_R1240_U488, P1_R1240_U489);
  nand ginst5435 (P1_R1240_U491, P1_R1240_U359, P1_R1240_U94);
  nand ginst5436 (P1_R1240_U492, P1_R1240_U335, P1_R1240_U490);
  nand ginst5437 (P1_R1240_U493, P1_R1240_U67, P1_U3063);
  nand ginst5438 (P1_R1240_U494, P1_R1240_U68, P1_U3491);
  nand ginst5439 (P1_R1240_U495, P1_R1240_U493, P1_R1240_U494);
  nand ginst5440 (P1_R1240_U496, P1_R1240_U164, P1_R1240_U360);
  nand ginst5441 (P1_R1240_U497, P1_R1240_U241, P1_R1240_U495);
  nand ginst5442 (P1_R1240_U498, P1_R1240_U63, P1_U3062);
  nand ginst5443 (P1_R1240_U499, P1_R1240_U64, P1_U3488);
  and ginst5444 (P1_R1240_U5, P1_R1240_U177, P1_R1240_U178);
  not ginst5445 (P1_R1240_U50, P1_U4019);
  nand ginst5446 (P1_R1240_U500, P1_R1240_U30, P1_U3077);
  nand ginst5447 (P1_R1240_U501, P1_R1240_U31, P1_U3456);
  not ginst5448 (P1_R1240_U51, P1_U4020);
  not ginst5449 (P1_R1240_U52, P1_U3058);
  not ginst5450 (P1_R1240_U53, P1_U4021);
  not ginst5451 (P1_R1240_U54, P1_U3065);
  not ginst5452 (P1_R1240_U55, P1_U4024);
  not ginst5453 (P1_R1240_U56, P1_U3075);
  not ginst5454 (P1_R1240_U57, P1_U3506);
  not ginst5455 (P1_R1240_U58, P1_U3073);
  not ginst5456 (P1_R1240_U59, P1_U3069);
  and ginst5457 (P1_R1240_U6, P1_R1240_U193, P1_R1240_U194);
  nand ginst5458 (P1_R1240_U60, P1_U3073, P1_U3506);
  not ginst5459 (P1_R1240_U61, P1_U3509);
  nand ginst5460 (P1_R1240_U62, P1_U3084, P1_U3482);
  not ginst5461 (P1_R1240_U63, P1_U3488);
  not ginst5462 (P1_R1240_U64, P1_U3062);
  not ginst5463 (P1_R1240_U65, P1_U3494);
  not ginst5464 (P1_R1240_U66, P1_U3072);
  not ginst5465 (P1_R1240_U67, P1_U3491);
  not ginst5466 (P1_R1240_U68, P1_U3063);
  nand ginst5467 (P1_R1240_U69, P1_U3063, P1_U3491);
  and ginst5468 (P1_R1240_U7, P1_R1240_U233, P1_R1240_U234);
  not ginst5469 (P1_R1240_U70, P1_U3497);
  not ginst5470 (P1_R1240_U71, P1_U3080);
  not ginst5471 (P1_R1240_U72, P1_U3500);
  not ginst5472 (P1_R1240_U73, P1_U3079);
  not ginst5473 (P1_R1240_U74, P1_U3503);
  not ginst5474 (P1_R1240_U75, P1_U3074);
  not ginst5475 (P1_R1240_U76, P1_U3512);
  not ginst5476 (P1_R1240_U77, P1_U3082);
  nand ginst5477 (P1_R1240_U78, P1_U3082, P1_U3512);
  not ginst5478 (P1_R1240_U79, P1_U3514);
  and ginst5479 (P1_R1240_U8, P1_R1240_U242, P1_R1240_U243);
  not ginst5480 (P1_R1240_U80, P1_U3081);
  nand ginst5481 (P1_R1240_U81, P1_U3081, P1_U3514);
  not ginst5482 (P1_R1240_U82, P1_U4025);
  not ginst5483 (P1_R1240_U83, P1_U4023);
  not ginst5484 (P1_R1240_U84, P1_U3061);
  not ginst5485 (P1_R1240_U85, P1_U4022);
  not ginst5486 (P1_R1240_U86, P1_U3066);
  nand ginst5487 (P1_R1240_U87, P1_U3057, P1_U4019);
  not ginst5488 (P1_R1240_U88, P1_U3054);
  not ginst5489 (P1_R1240_U89, P1_U4017);
  and ginst5490 (P1_R1240_U9, P1_R1240_U260, P1_R1240_U261);
  nand ginst5491 (P1_R1240_U90, P1_R1240_U173, P1_R1240_U303);
  not ginst5492 (P1_R1240_U91, P1_U3076);
  nand ginst5493 (P1_R1240_U92, P1_R1240_U312, P1_R1240_U78);
  nand ginst5494 (P1_R1240_U93, P1_R1240_U257, P1_R1240_U258);
  nand ginst5495 (P1_R1240_U94, P1_R1240_U334, P1_R1240_U69);
  nand ginst5496 (P1_R1240_U95, P1_R1240_U453, P1_R1240_U454);
  nand ginst5497 (P1_R1240_U96, P1_R1240_U500, P1_R1240_U501);
  nand ginst5498 (P1_R1240_U97, P1_R1240_U371, P1_R1240_U372);
  nand ginst5499 (P1_R1240_U98, P1_R1240_U376, P1_R1240_U377);
  nand ginst5500 (P1_R1240_U99, P1_R1240_U383, P1_R1240_U384);
  and ginst5501 (P1_R1282_U10, P1_R1282_U129, P1_R1282_U39);
  not ginst5502 (P1_R1282_U100, P1_R1282_U36);
  not ginst5503 (P1_R1282_U101, P1_R1282_U37);
  not ginst5504 (P1_R1282_U102, P1_R1282_U38);
  not ginst5505 (P1_R1282_U103, P1_R1282_U39);
  not ginst5506 (P1_R1282_U104, P1_R1282_U40);
  not ginst5507 (P1_R1282_U105, P1_R1282_U41);
  not ginst5508 (P1_R1282_U106, P1_R1282_U42);
  not ginst5509 (P1_R1282_U107, P1_R1282_U43);
  not ginst5510 (P1_R1282_U108, P1_R1282_U44);
  not ginst5511 (P1_R1282_U109, P1_R1282_U45);
  and ginst5512 (P1_R1282_U11, P1_R1282_U128, P1_R1282_U40);
  not ginst5513 (P1_R1282_U110, P1_R1282_U46);
  not ginst5514 (P1_R1282_U111, P1_R1282_U67);
  nand ginst5515 (P1_R1282_U112, P1_R1282_U110, P1_R1282_U69);
  nand ginst5516 (P1_R1282_U113, P1_R1282_U112, P1_U4027);
  or ginst5517 (P1_R1282_U114, P1_U3456, P1_U3461);
  nand ginst5518 (P1_R1282_U115, P1_R1282_U114, P1_U3464);
  nand ginst5519 (P1_R1282_U116, P1_R1282_U109, P1_R1282_U71);
  nand ginst5520 (P1_R1282_U117, P1_R1282_U116, P1_U4017);
  nand ginst5521 (P1_R1282_U118, P1_R1282_U108, P1_R1282_U73);
  nand ginst5522 (P1_R1282_U119, P1_R1282_U118, P1_U4019);
  and ginst5523 (P1_R1282_U12, P1_R1282_U127, P1_R1282_U41);
  nand ginst5524 (P1_R1282_U120, P1_R1282_U107, P1_R1282_U75);
  nand ginst5525 (P1_R1282_U121, P1_R1282_U120, P1_U4021);
  nand ginst5526 (P1_R1282_U122, P1_R1282_U106, P1_R1282_U77);
  nand ginst5527 (P1_R1282_U123, P1_R1282_U122, P1_U4023);
  nand ginst5528 (P1_R1282_U124, P1_R1282_U105, P1_R1282_U81);
  nand ginst5529 (P1_R1282_U125, P1_R1282_U124, P1_U4025);
  nand ginst5530 (P1_R1282_U126, P1_R1282_U104, P1_R1282_U83);
  nand ginst5531 (P1_R1282_U127, P1_R1282_U126, P1_U3512);
  nand ginst5532 (P1_R1282_U128, P1_R1282_U39, P1_U3506);
  nand ginst5533 (P1_R1282_U129, P1_R1282_U38, P1_U3503);
  and ginst5534 (P1_R1282_U13, P1_R1282_U125, P1_R1282_U42);
  nand ginst5535 (P1_R1282_U130, P1_R1282_U101, P1_R1282_U85);
  nand ginst5536 (P1_R1282_U131, P1_R1282_U130, P1_U3500);
  nand ginst5537 (P1_R1282_U132, P1_R1282_U36, P1_U3494);
  nand ginst5538 (P1_R1282_U133, P1_R1282_U35, P1_U3491);
  nand ginst5539 (P1_R1282_U134, P1_R1282_U62, P1_R1282_U92);
  nand ginst5540 (P1_R1282_U135, P1_R1282_U134, P1_U3488);
  nand ginst5541 (P1_R1282_U136, P1_R1282_U30, P1_U3485);
  nand ginst5542 (P1_R1282_U137, P1_R1282_U62, P1_R1282_U92);
  nand ginst5543 (P1_R1282_U138, P1_R1282_U27, P1_U3473);
  nand ginst5544 (P1_R1282_U139, P1_R1282_U64, P1_R1282_U89);
  and ginst5545 (P1_R1282_U14, P1_R1282_U123, P1_R1282_U43);
  nand ginst5546 (P1_R1282_U140, P1_R1282_U67, P1_U4026);
  nand ginst5547 (P1_R1282_U141, P1_R1282_U111, P1_R1282_U66);
  nand ginst5548 (P1_R1282_U142, P1_R1282_U46, P1_U4028);
  nand ginst5549 (P1_R1282_U143, P1_R1282_U110, P1_R1282_U69);
  nand ginst5550 (P1_R1282_U144, P1_R1282_U45, P1_U4018);
  nand ginst5551 (P1_R1282_U145, P1_R1282_U109, P1_R1282_U71);
  nand ginst5552 (P1_R1282_U146, P1_R1282_U44, P1_U4020);
  nand ginst5553 (P1_R1282_U147, P1_R1282_U108, P1_R1282_U73);
  nand ginst5554 (P1_R1282_U148, P1_R1282_U43, P1_U4022);
  nand ginst5555 (P1_R1282_U149, P1_R1282_U107, P1_R1282_U75);
  and ginst5556 (P1_R1282_U15, P1_R1282_U121, P1_R1282_U44);
  nand ginst5557 (P1_R1282_U150, P1_R1282_U42, P1_U4024);
  nand ginst5558 (P1_R1282_U151, P1_R1282_U106, P1_R1282_U77);
  nand ginst5559 (P1_R1282_U152, P1_R1282_U80, P1_U3461);
  nand ginst5560 (P1_R1282_U153, P1_R1282_U79, P1_U3456);
  nand ginst5561 (P1_R1282_U154, P1_R1282_U41, P1_U3514);
  nand ginst5562 (P1_R1282_U155, P1_R1282_U105, P1_R1282_U81);
  nand ginst5563 (P1_R1282_U156, P1_R1282_U40, P1_U3509);
  nand ginst5564 (P1_R1282_U157, P1_R1282_U104, P1_R1282_U83);
  nand ginst5565 (P1_R1282_U158, P1_R1282_U37, P1_U3497);
  nand ginst5566 (P1_R1282_U159, P1_R1282_U101, P1_R1282_U85);
  and ginst5567 (P1_R1282_U16, P1_R1282_U119, P1_R1282_U45);
  and ginst5568 (P1_R1282_U17, P1_R1282_U117, P1_R1282_U46);
  and ginst5569 (P1_R1282_U18, P1_R1282_U115, P1_R1282_U25);
  and ginst5570 (P1_R1282_U19, P1_R1282_U113, P1_R1282_U67);
  and ginst5571 (P1_R1282_U20, P1_R1282_U26, P1_R1282_U98);
  and ginst5572 (P1_R1282_U21, P1_R1282_U27, P1_R1282_U97);
  and ginst5573 (P1_R1282_U22, P1_R1282_U28, P1_R1282_U96);
  and ginst5574 (P1_R1282_U23, P1_R1282_U29, P1_R1282_U94);
  and ginst5575 (P1_R1282_U24, P1_R1282_U30, P1_R1282_U93);
  or ginst5576 (P1_R1282_U25, P1_U3456, P1_U3461, P1_U3464);
  nand ginst5577 (P1_R1282_U26, P1_R1282_U34, P1_R1282_U87);
  nand ginst5578 (P1_R1282_U27, P1_R1282_U33, P1_R1282_U88);
  nand ginst5579 (P1_R1282_U28, P1_R1282_U57, P1_R1282_U89);
  nand ginst5580 (P1_R1282_U29, P1_R1282_U32, P1_R1282_U90);
  nand ginst5581 (P1_R1282_U30, P1_R1282_U31, P1_R1282_U91);
  not ginst5582 (P1_R1282_U31, P1_U3482);
  not ginst5583 (P1_R1282_U32, P1_U3479);
  not ginst5584 (P1_R1282_U33, P1_U3470);
  not ginst5585 (P1_R1282_U34, P1_U3467);
  nand ginst5586 (P1_R1282_U35, P1_R1282_U58, P1_R1282_U92);
  nand ginst5587 (P1_R1282_U36, P1_R1282_U55, P1_R1282_U99);
  nand ginst5588 (P1_R1282_U37, P1_R1282_U100, P1_R1282_U54);
  nand ginst5589 (P1_R1282_U38, P1_R1282_U101, P1_R1282_U59);
  nand ginst5590 (P1_R1282_U39, P1_R1282_U102, P1_R1282_U53);
  nand ginst5591 (P1_R1282_U40, P1_R1282_U103, P1_R1282_U52);
  nand ginst5592 (P1_R1282_U41, P1_R1282_U104, P1_R1282_U60);
  nand ginst5593 (P1_R1282_U42, P1_R1282_U105, P1_R1282_U61);
  nand ginst5594 (P1_R1282_U43, P1_R1282_U106, P1_R1282_U51, P1_R1282_U77);
  nand ginst5595 (P1_R1282_U44, P1_R1282_U107, P1_R1282_U50, P1_R1282_U75);
  nand ginst5596 (P1_R1282_U45, P1_R1282_U108, P1_R1282_U49, P1_R1282_U73);
  nand ginst5597 (P1_R1282_U46, P1_R1282_U109, P1_R1282_U48, P1_R1282_U71);
  not ginst5598 (P1_R1282_U47, P1_U4027);
  not ginst5599 (P1_R1282_U48, P1_U4017);
  not ginst5600 (P1_R1282_U49, P1_U4019);
  not ginst5601 (P1_R1282_U50, P1_U4021);
  not ginst5602 (P1_R1282_U51, P1_U4023);
  not ginst5603 (P1_R1282_U52, P1_U3506);
  not ginst5604 (P1_R1282_U53, P1_U3503);
  not ginst5605 (P1_R1282_U54, P1_U3494);
  not ginst5606 (P1_R1282_U55, P1_U3491);
  nand ginst5607 (P1_R1282_U56, P1_R1282_U152, P1_R1282_U153);
  nor ginst5608 (P1_R1282_U57, P1_U3473, P1_U3476);
  nor ginst5609 (P1_R1282_U58, P1_U3485, P1_U3488);
  nor ginst5610 (P1_R1282_U59, P1_U3497, P1_U3500);
  and ginst5611 (P1_R1282_U6, P1_R1282_U135, P1_R1282_U35);
  nor ginst5612 (P1_R1282_U60, P1_U3509, P1_U3512);
  nor ginst5613 (P1_R1282_U61, P1_U3514, P1_U4025);
  not ginst5614 (P1_R1282_U62, P1_U3485);
  and ginst5615 (P1_R1282_U63, P1_R1282_U136, P1_R1282_U137);
  not ginst5616 (P1_R1282_U64, P1_U3473);
  and ginst5617 (P1_R1282_U65, P1_R1282_U138, P1_R1282_U139);
  not ginst5618 (P1_R1282_U66, P1_U4026);
  nand ginst5619 (P1_R1282_U67, P1_R1282_U110, P1_R1282_U47, P1_R1282_U69);
  and ginst5620 (P1_R1282_U68, P1_R1282_U140, P1_R1282_U141);
  not ginst5621 (P1_R1282_U69, P1_U4028);
  and ginst5622 (P1_R1282_U7, P1_R1282_U133, P1_R1282_U36);
  and ginst5623 (P1_R1282_U70, P1_R1282_U142, P1_R1282_U143);
  not ginst5624 (P1_R1282_U71, P1_U4018);
  and ginst5625 (P1_R1282_U72, P1_R1282_U144, P1_R1282_U145);
  not ginst5626 (P1_R1282_U73, P1_U4020);
  and ginst5627 (P1_R1282_U74, P1_R1282_U146, P1_R1282_U147);
  not ginst5628 (P1_R1282_U75, P1_U4022);
  and ginst5629 (P1_R1282_U76, P1_R1282_U148, P1_R1282_U149);
  not ginst5630 (P1_R1282_U77, P1_U4024);
  and ginst5631 (P1_R1282_U78, P1_R1282_U150, P1_R1282_U151);
  not ginst5632 (P1_R1282_U79, P1_U3461);
  and ginst5633 (P1_R1282_U8, P1_R1282_U132, P1_R1282_U37);
  not ginst5634 (P1_R1282_U80, P1_U3456);
  not ginst5635 (P1_R1282_U81, P1_U3514);
  and ginst5636 (P1_R1282_U82, P1_R1282_U154, P1_R1282_U155);
  not ginst5637 (P1_R1282_U83, P1_U3509);
  and ginst5638 (P1_R1282_U84, P1_R1282_U156, P1_R1282_U157);
  not ginst5639 (P1_R1282_U85, P1_U3497);
  and ginst5640 (P1_R1282_U86, P1_R1282_U158, P1_R1282_U159);
  not ginst5641 (P1_R1282_U87, P1_R1282_U25);
  not ginst5642 (P1_R1282_U88, P1_R1282_U26);
  not ginst5643 (P1_R1282_U89, P1_R1282_U27);
  and ginst5644 (P1_R1282_U9, P1_R1282_U131, P1_R1282_U38);
  not ginst5645 (P1_R1282_U90, P1_R1282_U28);
  not ginst5646 (P1_R1282_U91, P1_R1282_U29);
  not ginst5647 (P1_R1282_U92, P1_R1282_U30);
  nand ginst5648 (P1_R1282_U93, P1_R1282_U29, P1_U3482);
  nand ginst5649 (P1_R1282_U94, P1_R1282_U28, P1_U3479);
  nand ginst5650 (P1_R1282_U95, P1_R1282_U64, P1_R1282_U89);
  nand ginst5651 (P1_R1282_U96, P1_R1282_U95, P1_U3476);
  nand ginst5652 (P1_R1282_U97, P1_R1282_U26, P1_U3470);
  nand ginst5653 (P1_R1282_U98, P1_R1282_U25, P1_U3467);
  not ginst5654 (P1_R1282_U99, P1_R1282_U35);
  nand ginst5655 (P1_R1309_U10, P1_R1309_U7, P1_U3059);
  not ginst5656 (P1_R1309_U6, P1_U3059);
  not ginst5657 (P1_R1309_U7, P1_U3056);
  and ginst5658 (P1_R1309_U8, P1_R1309_U10, P1_R1309_U9);
  nand ginst5659 (P1_R1309_U9, P1_R1309_U6, P1_U3056);
  and ginst5660 (P1_R1352_U6, P1_R1352_U7, P1_U3059);
  not ginst5661 (P1_R1352_U7, P1_U3056);
  not ginst5662 (P1_R1375_U10, P1_U3088);
  and ginst5663 (P1_R1375_U100, P1_R1375_U196, P1_R1375_U197);
  not ginst5664 (P1_R1375_U101, P1_U3122);
  nand ginst5665 (P1_R1375_U102, P1_U3150, P1_U3151);
  nand ginst5666 (P1_R1375_U103, P1_R1375_U102, P1_U3118);
  or ginst5667 (P1_R1375_U104, P1_U3150, P1_U3151);
  nand ginst5668 (P1_R1375_U105, P1_R1375_U16, P1_U3117);
  nand ginst5669 (P1_R1375_U106, P1_R1375_U103, P1_R1375_U104, P1_R1375_U105);
  nand ginst5670 (P1_R1375_U107, P1_R1375_U15, P1_U3149);
  nand ginst5671 (P1_R1375_U108, P1_R1375_U18, P1_U3148);
  nand ginst5672 (P1_R1375_U109, P1_R1375_U106, P1_R1375_U70);
  not ginst5673 (P1_R1375_U11, P1_U3087);
  nand ginst5674 (P1_R1375_U110, P1_R1375_U17, P1_U3116);
  nand ginst5675 (P1_R1375_U111, P1_R1375_U20, P1_U3115);
  nand ginst5676 (P1_R1375_U112, P1_R1375_U109, P1_R1375_U71);
  nand ginst5677 (P1_R1375_U113, P1_R1375_U19, P1_U3147);
  nand ginst5678 (P1_R1375_U114, P1_R1375_U22, P1_U3146);
  nand ginst5679 (P1_R1375_U115, P1_R1375_U112, P1_R1375_U72);
  nand ginst5680 (P1_R1375_U116, P1_R1375_U21, P1_U3114);
  nand ginst5681 (P1_R1375_U117, P1_R1375_U24, P1_U3113);
  nand ginst5682 (P1_R1375_U118, P1_R1375_U115, P1_R1375_U73);
  nand ginst5683 (P1_R1375_U119, P1_R1375_U23, P1_U3145);
  not ginst5684 (P1_R1375_U12, P1_U3121);
  nand ginst5685 (P1_R1375_U120, P1_R1375_U26, P1_U3144);
  nand ginst5686 (P1_R1375_U121, P1_R1375_U118, P1_R1375_U74);
  nand ginst5687 (P1_R1375_U122, P1_R1375_U25, P1_U3112);
  nand ginst5688 (P1_R1375_U123, P1_R1375_U28, P1_U3111);
  nand ginst5689 (P1_R1375_U124, P1_R1375_U121, P1_R1375_U75);
  nand ginst5690 (P1_R1375_U125, P1_R1375_U27, P1_U3143);
  nand ginst5691 (P1_R1375_U126, P1_R1375_U30, P1_U3142);
  nand ginst5692 (P1_R1375_U127, P1_R1375_U124, P1_R1375_U76);
  nand ginst5693 (P1_R1375_U128, P1_R1375_U29, P1_U3110);
  nand ginst5694 (P1_R1375_U129, P1_R1375_U32, P1_U3109);
  not ginst5695 (P1_R1375_U13, P1_U3120);
  nand ginst5696 (P1_R1375_U130, P1_R1375_U127, P1_R1375_U77);
  nand ginst5697 (P1_R1375_U131, P1_R1375_U31, P1_U3141);
  nand ginst5698 (P1_R1375_U132, P1_R1375_U34, P1_U3140);
  nand ginst5699 (P1_R1375_U133, P1_R1375_U130, P1_R1375_U78);
  nand ginst5700 (P1_R1375_U134, P1_R1375_U33, P1_U3108);
  nand ginst5701 (P1_R1375_U135, P1_R1375_U36, P1_U3107);
  nand ginst5702 (P1_R1375_U136, P1_R1375_U133, P1_R1375_U79);
  nand ginst5703 (P1_R1375_U137, P1_R1375_U35, P1_U3139);
  nand ginst5704 (P1_R1375_U138, P1_R1375_U38, P1_U3138);
  nand ginst5705 (P1_R1375_U139, P1_R1375_U136, P1_R1375_U80);
  not ginst5706 (P1_R1375_U14, P1_U3152);
  nand ginst5707 (P1_R1375_U140, P1_R1375_U37, P1_U3106);
  nand ginst5708 (P1_R1375_U141, P1_R1375_U40, P1_U3105);
  nand ginst5709 (P1_R1375_U142, P1_R1375_U139, P1_R1375_U81);
  nand ginst5710 (P1_R1375_U143, P1_R1375_U39, P1_U3137);
  nand ginst5711 (P1_R1375_U144, P1_R1375_U42, P1_U3136);
  nand ginst5712 (P1_R1375_U145, P1_R1375_U142, P1_R1375_U82);
  nand ginst5713 (P1_R1375_U146, P1_R1375_U41, P1_U3104);
  nand ginst5714 (P1_R1375_U147, P1_R1375_U44, P1_U3103);
  nand ginst5715 (P1_R1375_U148, P1_R1375_U145, P1_R1375_U83);
  nand ginst5716 (P1_R1375_U149, P1_R1375_U43, P1_U3135);
  not ginst5717 (P1_R1375_U15, P1_U3117);
  nand ginst5718 (P1_R1375_U150, P1_R1375_U46, P1_U3134);
  nand ginst5719 (P1_R1375_U151, P1_R1375_U148, P1_R1375_U84);
  nand ginst5720 (P1_R1375_U152, P1_R1375_U45, P1_U3102);
  nand ginst5721 (P1_R1375_U153, P1_R1375_U48, P1_U3101);
  nand ginst5722 (P1_R1375_U154, P1_R1375_U151, P1_R1375_U85);
  nand ginst5723 (P1_R1375_U155, P1_R1375_U47, P1_U3133);
  nand ginst5724 (P1_R1375_U156, P1_R1375_U50, P1_U3132);
  nand ginst5725 (P1_R1375_U157, P1_R1375_U154, P1_R1375_U86);
  nand ginst5726 (P1_R1375_U158, P1_R1375_U49, P1_U3100);
  nand ginst5727 (P1_R1375_U159, P1_R1375_U52, P1_U3099);
  not ginst5728 (P1_R1375_U16, P1_U3149);
  nand ginst5729 (P1_R1375_U160, P1_R1375_U157, P1_R1375_U87);
  nand ginst5730 (P1_R1375_U161, P1_R1375_U51, P1_U3131);
  nand ginst5731 (P1_R1375_U162, P1_R1375_U54, P1_U3130);
  nand ginst5732 (P1_R1375_U163, P1_R1375_U160, P1_R1375_U88);
  nand ginst5733 (P1_R1375_U164, P1_R1375_U53, P1_U3098);
  nand ginst5734 (P1_R1375_U165, P1_R1375_U56, P1_U3097);
  nand ginst5735 (P1_R1375_U166, P1_R1375_U163, P1_R1375_U89);
  nand ginst5736 (P1_R1375_U167, P1_R1375_U55, P1_U3129);
  nand ginst5737 (P1_R1375_U168, P1_R1375_U58, P1_U3128);
  nand ginst5738 (P1_R1375_U169, P1_R1375_U166, P1_R1375_U90);
  not ginst5739 (P1_R1375_U17, P1_U3148);
  nand ginst5740 (P1_R1375_U170, P1_R1375_U57, P1_U3096);
  nand ginst5741 (P1_R1375_U171, P1_R1375_U60, P1_U3095);
  nand ginst5742 (P1_R1375_U172, P1_R1375_U169, P1_R1375_U91);
  nand ginst5743 (P1_R1375_U173, P1_R1375_U59, P1_U3127);
  nand ginst5744 (P1_R1375_U174, P1_R1375_U62, P1_U3126);
  nand ginst5745 (P1_R1375_U175, P1_R1375_U172, P1_R1375_U92);
  nand ginst5746 (P1_R1375_U176, P1_R1375_U61, P1_U3094);
  nand ginst5747 (P1_R1375_U177, P1_R1375_U64, P1_U3093);
  nand ginst5748 (P1_R1375_U178, P1_R1375_U175, P1_R1375_U93);
  nand ginst5749 (P1_R1375_U179, P1_R1375_U63, P1_U3125);
  not ginst5750 (P1_R1375_U18, P1_U3116);
  nand ginst5751 (P1_R1375_U180, P1_R1375_U66, P1_U3124);
  nand ginst5752 (P1_R1375_U181, P1_R1375_U178, P1_R1375_U94);
  nand ginst5753 (P1_R1375_U182, P1_R1375_U65, P1_U3092);
  nand ginst5754 (P1_R1375_U183, P1_R1375_U68, P1_U3091);
  nand ginst5755 (P1_R1375_U184, P1_R1375_U181, P1_R1375_U95);
  nand ginst5756 (P1_R1375_U185, P1_R1375_U184, P1_R1375_U96);
  nand ginst5757 (P1_R1375_U186, P1_R1375_U67, P1_U3123);
  nand ginst5758 (P1_R1375_U187, P1_R1375_U101, P1_U3090);
  nand ginst5759 (P1_R1375_U188, P1_R1375_U12, P1_U3089);
  nand ginst5760 (P1_R1375_U189, P1_R1375_U191, P1_R1375_U69, P1_R1375_U8, P1_U3121);
  not ginst5761 (P1_R1375_U19, P1_U3115);
  nand ginst5762 (P1_R1375_U190, P1_R1375_U10, P1_R1375_U8, P1_U3120);
  nand ginst5763 (P1_R1375_U191, P1_R1375_U13, P1_U3088);
  nand ginst5764 (P1_R1375_U192, P1_R1375_U185, P1_R1375_U193, P1_R1375_U6, P1_R1375_U98);
  nand ginst5765 (P1_R1375_U193, P1_R1375_U184, P1_R1375_U97);
  nand ginst5766 (P1_R1375_U194, P1_R1375_U99, P1_U3087);
  nand ginst5767 (P1_R1375_U195, P1_R1375_U11, P1_U3119);
  nand ginst5768 (P1_R1375_U196, P1_R1375_U99, P1_U3087, P1_U3152);
  nand ginst5769 (P1_R1375_U197, P1_R1375_U11, P1_R1375_U14, P1_U3119);
  not ginst5770 (P1_R1375_U20, P1_U3147);
  not ginst5771 (P1_R1375_U21, P1_U3146);
  not ginst5772 (P1_R1375_U22, P1_U3114);
  not ginst5773 (P1_R1375_U23, P1_U3113);
  not ginst5774 (P1_R1375_U24, P1_U3145);
  not ginst5775 (P1_R1375_U25, P1_U3144);
  not ginst5776 (P1_R1375_U26, P1_U3112);
  not ginst5777 (P1_R1375_U27, P1_U3111);
  not ginst5778 (P1_R1375_U28, P1_U3143);
  not ginst5779 (P1_R1375_U29, P1_U3142);
  not ginst5780 (P1_R1375_U30, P1_U3110);
  not ginst5781 (P1_R1375_U31, P1_U3109);
  not ginst5782 (P1_R1375_U32, P1_U3141);
  not ginst5783 (P1_R1375_U33, P1_U3140);
  not ginst5784 (P1_R1375_U34, P1_U3108);
  not ginst5785 (P1_R1375_U35, P1_U3107);
  not ginst5786 (P1_R1375_U36, P1_U3139);
  not ginst5787 (P1_R1375_U37, P1_U3138);
  not ginst5788 (P1_R1375_U38, P1_U3106);
  not ginst5789 (P1_R1375_U39, P1_U3105);
  not ginst5790 (P1_R1375_U40, P1_U3137);
  not ginst5791 (P1_R1375_U41, P1_U3136);
  not ginst5792 (P1_R1375_U42, P1_U3104);
  not ginst5793 (P1_R1375_U43, P1_U3103);
  not ginst5794 (P1_R1375_U44, P1_U3135);
  not ginst5795 (P1_R1375_U45, P1_U3134);
  not ginst5796 (P1_R1375_U46, P1_U3102);
  not ginst5797 (P1_R1375_U47, P1_U3101);
  not ginst5798 (P1_R1375_U48, P1_U3133);
  not ginst5799 (P1_R1375_U49, P1_U3132);
  not ginst5800 (P1_R1375_U50, P1_U3100);
  not ginst5801 (P1_R1375_U51, P1_U3099);
  not ginst5802 (P1_R1375_U52, P1_U3131);
  not ginst5803 (P1_R1375_U53, P1_U3130);
  not ginst5804 (P1_R1375_U54, P1_U3098);
  not ginst5805 (P1_R1375_U55, P1_U3097);
  not ginst5806 (P1_R1375_U56, P1_U3129);
  not ginst5807 (P1_R1375_U57, P1_U3128);
  not ginst5808 (P1_R1375_U58, P1_U3096);
  not ginst5809 (P1_R1375_U59, P1_U3095);
  and ginst5810 (P1_R1375_U6, P1_R1375_U191, P1_R1375_U8);
  not ginst5811 (P1_R1375_U60, P1_U3127);
  not ginst5812 (P1_R1375_U61, P1_U3126);
  not ginst5813 (P1_R1375_U62, P1_U3094);
  not ginst5814 (P1_R1375_U63, P1_U3093);
  not ginst5815 (P1_R1375_U64, P1_U3125);
  not ginst5816 (P1_R1375_U65, P1_U3124);
  not ginst5817 (P1_R1375_U66, P1_U3092);
  not ginst5818 (P1_R1375_U67, P1_U3091);
  not ginst5819 (P1_R1375_U68, P1_U3123);
  not ginst5820 (P1_R1375_U69, P1_U3089);
  and ginst5821 (P1_R1375_U7, P1_R1375_U100, P1_R1375_U189, P1_R1375_U190);
  and ginst5822 (P1_R1375_U70, P1_R1375_U107, P1_R1375_U108);
  and ginst5823 (P1_R1375_U71, P1_R1375_U110, P1_R1375_U111);
  and ginst5824 (P1_R1375_U72, P1_R1375_U113, P1_R1375_U114);
  and ginst5825 (P1_R1375_U73, P1_R1375_U116, P1_R1375_U117);
  and ginst5826 (P1_R1375_U74, P1_R1375_U119, P1_R1375_U120);
  and ginst5827 (P1_R1375_U75, P1_R1375_U122, P1_R1375_U123);
  and ginst5828 (P1_R1375_U76, P1_R1375_U125, P1_R1375_U126);
  and ginst5829 (P1_R1375_U77, P1_R1375_U128, P1_R1375_U129);
  and ginst5830 (P1_R1375_U78, P1_R1375_U131, P1_R1375_U132);
  and ginst5831 (P1_R1375_U79, P1_R1375_U134, P1_R1375_U135);
  and ginst5832 (P1_R1375_U8, P1_R1375_U194, P1_R1375_U195);
  and ginst5833 (P1_R1375_U80, P1_R1375_U137, P1_R1375_U138);
  and ginst5834 (P1_R1375_U81, P1_R1375_U140, P1_R1375_U141);
  and ginst5835 (P1_R1375_U82, P1_R1375_U143, P1_R1375_U144);
  and ginst5836 (P1_R1375_U83, P1_R1375_U146, P1_R1375_U147);
  and ginst5837 (P1_R1375_U84, P1_R1375_U149, P1_R1375_U150);
  and ginst5838 (P1_R1375_U85, P1_R1375_U152, P1_R1375_U153);
  and ginst5839 (P1_R1375_U86, P1_R1375_U155, P1_R1375_U156);
  and ginst5840 (P1_R1375_U87, P1_R1375_U158, P1_R1375_U159);
  and ginst5841 (P1_R1375_U88, P1_R1375_U161, P1_R1375_U162);
  and ginst5842 (P1_R1375_U89, P1_R1375_U164, P1_R1375_U165);
  nand ginst5843 (P1_R1375_U9, P1_R1375_U192, P1_R1375_U7);
  and ginst5844 (P1_R1375_U90, P1_R1375_U167, P1_R1375_U168);
  and ginst5845 (P1_R1375_U91, P1_R1375_U170, P1_R1375_U171);
  and ginst5846 (P1_R1375_U92, P1_R1375_U173, P1_R1375_U174);
  and ginst5847 (P1_R1375_U93, P1_R1375_U176, P1_R1375_U177);
  and ginst5848 (P1_R1375_U94, P1_R1375_U179, P1_R1375_U180);
  and ginst5849 (P1_R1375_U95, P1_R1375_U182, P1_R1375_U183);
  and ginst5850 (P1_R1375_U96, P1_R1375_U101, P1_R1375_U186);
  and ginst5851 (P1_R1375_U97, P1_R1375_U186, P1_U3090);
  and ginst5852 (P1_R1375_U98, P1_R1375_U187, P1_R1375_U188);
  not ginst5853 (P1_R1375_U99, P1_U3119);
  and ginst5854 (P1_SUB_88_U10, P1_SUB_88_U195, P1_SUB_88_U221);
  nor ginst5855 (P1_SUB_88_U100, P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN, P1_IR_REG_20__SCAN_IN);
  and ginst5856 (P1_SUB_88_U101, P1_SUB_88_U100, P1_SUB_88_U97, P1_SUB_88_U98, P1_SUB_88_U99);
  nor ginst5857 (P1_SUB_88_U102, P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN);
  nor ginst5858 (P1_SUB_88_U103, P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN, P1_IR_REG_25__SCAN_IN);
  nor ginst5859 (P1_SUB_88_U104, P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN);
  nor ginst5860 (P1_SUB_88_U105, P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN);
  and ginst5861 (P1_SUB_88_U106, P1_SUB_88_U102, P1_SUB_88_U103, P1_SUB_88_U104, P1_SUB_88_U105);
  nor ginst5862 (P1_SUB_88_U107, P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN);
  nor ginst5863 (P1_SUB_88_U108, P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN);
  nor ginst5864 (P1_SUB_88_U109, P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN);
  and ginst5865 (P1_SUB_88_U11, P1_SUB_88_U220, P1_SUB_88_U34);
  nor ginst5866 (P1_SUB_88_U110, P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN, P1_IR_REG_20__SCAN_IN);
  and ginst5867 (P1_SUB_88_U111, P1_SUB_88_U107, P1_SUB_88_U108, P1_SUB_88_U109, P1_SUB_88_U110);
  nor ginst5868 (P1_SUB_88_U112, P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN);
  nor ginst5869 (P1_SUB_88_U113, P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN, P1_IR_REG_24__SCAN_IN);
  nor ginst5870 (P1_SUB_88_U114, P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN);
  nor ginst5871 (P1_SUB_88_U115, P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN);
  and ginst5872 (P1_SUB_88_U116, P1_SUB_88_U112, P1_SUB_88_U113, P1_SUB_88_U114, P1_SUB_88_U115);
  nor ginst5873 (P1_SUB_88_U117, P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN);
  nor ginst5874 (P1_SUB_88_U118, P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN);
  nor ginst5875 (P1_SUB_88_U119, P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN);
  and ginst5876 (P1_SUB_88_U12, P1_SUB_88_U197, P1_SUB_88_U219);
  nor ginst5877 (P1_SUB_88_U120, P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN, P1_IR_REG_19__SCAN_IN);
  and ginst5878 (P1_SUB_88_U121, P1_SUB_88_U117, P1_SUB_88_U118, P1_SUB_88_U119, P1_SUB_88_U120);
  nor ginst5879 (P1_SUB_88_U122, P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN);
  nor ginst5880 (P1_SUB_88_U123, P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN, P1_IR_REG_23__SCAN_IN);
  nor ginst5881 (P1_SUB_88_U124, P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN);
  nor ginst5882 (P1_SUB_88_U125, P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN);
  and ginst5883 (P1_SUB_88_U126, P1_SUB_88_U122, P1_SUB_88_U123, P1_SUB_88_U124, P1_SUB_88_U125);
  nor ginst5884 (P1_SUB_88_U127, P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN);
  nor ginst5885 (P1_SUB_88_U128, P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN, P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN);
  nor ginst5886 (P1_SUB_88_U129, P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN);
  and ginst5887 (P1_SUB_88_U13, P1_SUB_88_U198, P1_SUB_88_U217);
  nor ginst5888 (P1_SUB_88_U130, P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN);
  nor ginst5889 (P1_SUB_88_U131, P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN);
  nor ginst5890 (P1_SUB_88_U132, P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN);
  nor ginst5891 (P1_SUB_88_U133, P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN);
  and ginst5892 (P1_SUB_88_U134, P1_SUB_88_U131, P1_SUB_88_U132, P1_SUB_88_U133);
  nor ginst5893 (P1_SUB_88_U135, P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN);
  nor ginst5894 (P1_SUB_88_U136, P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN);
  and ginst5895 (P1_SUB_88_U137, P1_SUB_88_U135, P1_SUB_88_U136);
  nor ginst5896 (P1_SUB_88_U138, P1_IR_REG_1__SCAN_IN, P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN);
  nor ginst5897 (P1_SUB_88_U139, P1_IR_REG_0__SCAN_IN, P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN);
  and ginst5898 (P1_SUB_88_U14, P1_SUB_88_U172, P1_SUB_88_U216);
  nor ginst5899 (P1_SUB_88_U140, P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN);
  and ginst5900 (P1_SUB_88_U141, P1_SUB_88_U139, P1_SUB_88_U140);
  nor ginst5901 (P1_SUB_88_U142, P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN);
  nor ginst5902 (P1_SUB_88_U143, P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN);
  nor ginst5903 (P1_SUB_88_U144, P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN);
  nor ginst5904 (P1_SUB_88_U145, P1_IR_REG_1__SCAN_IN, P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN);
  nor ginst5905 (P1_SUB_88_U146, P1_IR_REG_0__SCAN_IN, P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN, P1_IR_REG_20__SCAN_IN);
  nor ginst5906 (P1_SUB_88_U147, P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN);
  nor ginst5907 (P1_SUB_88_U148, P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN);
  nor ginst5908 (P1_SUB_88_U149, P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN);
  and ginst5909 (P1_SUB_88_U15, P1_SUB_88_U200, P1_SUB_88_U215);
  nor ginst5910 (P1_SUB_88_U150, P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN);
  nor ginst5911 (P1_SUB_88_U151, P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN);
  nor ginst5912 (P1_SUB_88_U152, P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN);
  nor ginst5913 (P1_SUB_88_U153, P1_IR_REG_1__SCAN_IN, P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN);
  nor ginst5914 (P1_SUB_88_U154, P1_IR_REG_0__SCAN_IN, P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN);
  nor ginst5915 (P1_SUB_88_U155, P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN);
  nor ginst5916 (P1_SUB_88_U156, P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN);
  nor ginst5917 (P1_SUB_88_U157, P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN);
  nor ginst5918 (P1_SUB_88_U158, P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN);
  not ginst5919 (P1_SUB_88_U159, P1_IR_REG_9__SCAN_IN);
  and ginst5920 (P1_SUB_88_U16, P1_SUB_88_U201, P1_SUB_88_U213);
  and ginst5921 (P1_SUB_88_U160, P1_SUB_88_U232, P1_SUB_88_U233);
  not ginst5922 (P1_SUB_88_U161, P1_IR_REG_5__SCAN_IN);
  and ginst5923 (P1_SUB_88_U162, P1_SUB_88_U234, P1_SUB_88_U235);
  not ginst5924 (P1_SUB_88_U163, P1_IR_REG_31__SCAN_IN);
  not ginst5925 (P1_SUB_88_U164, P1_IR_REG_30__SCAN_IN);
  and ginst5926 (P1_SUB_88_U165, P1_SUB_88_U238, P1_SUB_88_U239);
  not ginst5927 (P1_SUB_88_U166, P1_IR_REG_27__SCAN_IN);
  nand ginst5928 (P1_SUB_88_U167, P1_SUB_88_U91, P1_SUB_88_U96);
  not ginst5929 (P1_SUB_88_U168, P1_IR_REG_25__SCAN_IN);
  nand ginst5930 (P1_SUB_88_U169, P1_SUB_88_U111, P1_SUB_88_U116);
  and ginst5931 (P1_SUB_88_U17, P1_SUB_88_U169, P1_SUB_88_U212);
  and ginst5932 (P1_SUB_88_U170, P1_SUB_88_U242, P1_SUB_88_U243);
  not ginst5933 (P1_SUB_88_U171, P1_IR_REG_21__SCAN_IN);
  nand ginst5934 (P1_SUB_88_U172, P1_SUB_88_U143, P1_SUB_88_U144, P1_SUB_88_U145, P1_SUB_88_U146, P1_SUB_88_U147);
  and ginst5935 (P1_SUB_88_U173, P1_SUB_88_U244, P1_SUB_88_U245);
  not ginst5936 (P1_SUB_88_U174, P1_IR_REG_1__SCAN_IN);
  not ginst5937 (P1_SUB_88_U175, P1_IR_REG_0__SCAN_IN);
  not ginst5938 (P1_SUB_88_U176, P1_IR_REG_17__SCAN_IN);
  and ginst5939 (P1_SUB_88_U177, P1_SUB_88_U248, P1_SUB_88_U249);
  not ginst5940 (P1_SUB_88_U178, P1_IR_REG_13__SCAN_IN);
  and ginst5941 (P1_SUB_88_U179, P1_SUB_88_U250, P1_SUB_88_U251);
  and ginst5942 (P1_SUB_88_U18, P1_SUB_88_U167, P1_SUB_88_U211);
  nand ginst5943 (P1_SUB_88_U180, P1_SUB_88_U230, P1_SUB_88_U32);
  not ginst5944 (P1_SUB_88_U181, P1_SUB_88_U29);
  not ginst5945 (P1_SUB_88_U182, P1_SUB_88_U30);
  nand ginst5946 (P1_SUB_88_U183, P1_SUB_88_U182, P1_SUB_88_U31);
  not ginst5947 (P1_SUB_88_U184, P1_SUB_88_U28);
  nand ginst5948 (P1_SUB_88_U185, P1_IR_REG_8__SCAN_IN, P1_SUB_88_U183);
  nand ginst5949 (P1_SUB_88_U186, P1_IR_REG_7__SCAN_IN, P1_SUB_88_U30);
  nand ginst5950 (P1_SUB_88_U187, P1_SUB_88_U161, P1_SUB_88_U181);
  nand ginst5951 (P1_SUB_88_U188, P1_IR_REG_6__SCAN_IN, P1_SUB_88_U187);
  nand ginst5952 (P1_SUB_88_U189, P1_IR_REG_4__SCAN_IN, P1_SUB_88_U180);
  and ginst5953 (P1_SUB_88_U19, P1_SUB_88_U204, P1_SUB_88_U209);
  nand ginst5954 (P1_SUB_88_U190, P1_IR_REG_3__SCAN_IN, P1_SUB_88_U27);
  not ginst5955 (P1_SUB_88_U191, P1_SUB_88_U38);
  nand ginst5956 (P1_SUB_88_U192, P1_SUB_88_U191, P1_SUB_88_U39);
  not ginst5957 (P1_SUB_88_U193, P1_SUB_88_U35);
  not ginst5958 (P1_SUB_88_U194, P1_SUB_88_U36);
  nand ginst5959 (P1_SUB_88_U195, P1_SUB_88_U194, P1_SUB_88_U37);
  not ginst5960 (P1_SUB_88_U196, P1_SUB_88_U34);
  nand ginst5961 (P1_SUB_88_U197, P1_SUB_88_U152, P1_SUB_88_U153, P1_SUB_88_U154, P1_SUB_88_U155);
  nand ginst5962 (P1_SUB_88_U198, P1_SUB_88_U148, P1_SUB_88_U149, P1_SUB_88_U150, P1_SUB_88_U151);
  not ginst5963 (P1_SUB_88_U199, P1_SUB_88_U172);
  and ginst5964 (P1_SUB_88_U20, P1_SUB_88_U208, P1_SUB_88_U33);
  nand ginst5965 (P1_SUB_88_U200, P1_SUB_88_U134, P1_SUB_88_U196);
  nand ginst5966 (P1_SUB_88_U201, P1_SUB_88_U121, P1_SUB_88_U126);
  not ginst5967 (P1_SUB_88_U202, P1_SUB_88_U169);
  not ginst5968 (P1_SUB_88_U203, P1_SUB_88_U167);
  nand ginst5969 (P1_SUB_88_U204, P1_SUB_88_U61, P1_SUB_88_U66);
  not ginst5970 (P1_SUB_88_U205, P1_SUB_88_U33);
  or ginst5971 (P1_SUB_88_U206, P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN);
  nand ginst5972 (P1_SUB_88_U207, P1_IR_REG_2__SCAN_IN, P1_SUB_88_U206);
  nand ginst5973 (P1_SUB_88_U208, P1_IR_REG_29__SCAN_IN, P1_SUB_88_U204);
  nand ginst5974 (P1_SUB_88_U209, P1_IR_REG_28__SCAN_IN, P1_SUB_88_U229);
  and ginst5975 (P1_SUB_88_U21, P1_SUB_88_U207, P1_SUB_88_U27);
  nand ginst5976 (P1_SUB_88_U210, P1_SUB_88_U101, P1_SUB_88_U106);
  nand ginst5977 (P1_SUB_88_U211, P1_IR_REG_26__SCAN_IN, P1_SUB_88_U210);
  nand ginst5978 (P1_SUB_88_U212, P1_IR_REG_24__SCAN_IN, P1_SUB_88_U201);
  nand ginst5979 (P1_SUB_88_U213, P1_IR_REG_23__SCAN_IN, P1_SUB_88_U200);
  nand ginst5980 (P1_SUB_88_U214, P1_SUB_88_U137, P1_SUB_88_U138, P1_SUB_88_U141, P1_SUB_88_U142);
  nand ginst5981 (P1_SUB_88_U215, P1_IR_REG_22__SCAN_IN, P1_SUB_88_U214);
  nand ginst5982 (P1_SUB_88_U216, P1_IR_REG_20__SCAN_IN, P1_SUB_88_U198);
  nand ginst5983 (P1_SUB_88_U217, P1_IR_REG_19__SCAN_IN, P1_SUB_88_U197);
  nand ginst5984 (P1_SUB_88_U218, P1_SUB_88_U176, P1_SUB_88_U196);
  nand ginst5985 (P1_SUB_88_U219, P1_IR_REG_18__SCAN_IN, P1_SUB_88_U218);
  and ginst5986 (P1_SUB_88_U22, P1_SUB_88_U180, P1_SUB_88_U190);
  nand ginst5987 (P1_SUB_88_U220, P1_IR_REG_16__SCAN_IN, P1_SUB_88_U195);
  nand ginst5988 (P1_SUB_88_U221, P1_IR_REG_15__SCAN_IN, P1_SUB_88_U36);
  nand ginst5989 (P1_SUB_88_U222, P1_SUB_88_U178, P1_SUB_88_U193);
  nand ginst5990 (P1_SUB_88_U223, P1_IR_REG_14__SCAN_IN, P1_SUB_88_U222);
  nand ginst5991 (P1_SUB_88_U224, P1_IR_REG_12__SCAN_IN, P1_SUB_88_U192);
  nand ginst5992 (P1_SUB_88_U225, P1_IR_REG_11__SCAN_IN, P1_SUB_88_U38);
  nand ginst5993 (P1_SUB_88_U226, P1_SUB_88_U159, P1_SUB_88_U184);
  nand ginst5994 (P1_SUB_88_U227, P1_IR_REG_10__SCAN_IN, P1_SUB_88_U226);
  nand ginst5995 (P1_SUB_88_U228, P1_SUB_88_U164, P1_SUB_88_U205);
  nand ginst5996 (P1_SUB_88_U229, P1_SUB_88_U71, P1_SUB_88_U76);
  and ginst5997 (P1_SUB_88_U23, P1_SUB_88_U189, P1_SUB_88_U29);
  not ginst5998 (P1_SUB_88_U230, P1_SUB_88_U27);
  nand ginst5999 (P1_SUB_88_U231, P1_SUB_88_U81, P1_SUB_88_U86);
  nand ginst6000 (P1_SUB_88_U232, P1_IR_REG_9__SCAN_IN, P1_SUB_88_U28);
  nand ginst6001 (P1_SUB_88_U233, P1_SUB_88_U159, P1_SUB_88_U184);
  nand ginst6002 (P1_SUB_88_U234, P1_IR_REG_5__SCAN_IN, P1_SUB_88_U29);
  nand ginst6003 (P1_SUB_88_U235, P1_SUB_88_U161, P1_SUB_88_U181);
  nand ginst6004 (P1_SUB_88_U236, P1_SUB_88_U163, P1_SUB_88_U228);
  nand ginst6005 (P1_SUB_88_U237, P1_IR_REG_31__SCAN_IN, P1_SUB_88_U164, P1_SUB_88_U205);
  nand ginst6006 (P1_SUB_88_U238, P1_IR_REG_30__SCAN_IN, P1_SUB_88_U33);
  nand ginst6007 (P1_SUB_88_U239, P1_SUB_88_U164, P1_SUB_88_U205);
  and ginst6008 (P1_SUB_88_U24, P1_SUB_88_U188, P1_SUB_88_U30);
  nand ginst6009 (P1_SUB_88_U240, P1_IR_REG_27__SCAN_IN, P1_SUB_88_U203);
  nand ginst6010 (P1_SUB_88_U241, P1_SUB_88_U166, P1_SUB_88_U231);
  nand ginst6011 (P1_SUB_88_U242, P1_IR_REG_25__SCAN_IN, P1_SUB_88_U169);
  nand ginst6012 (P1_SUB_88_U243, P1_SUB_88_U168, P1_SUB_88_U202);
  nand ginst6013 (P1_SUB_88_U244, P1_IR_REG_21__SCAN_IN, P1_SUB_88_U172);
  nand ginst6014 (P1_SUB_88_U245, P1_SUB_88_U171, P1_SUB_88_U199);
  nand ginst6015 (P1_SUB_88_U246, P1_IR_REG_1__SCAN_IN, P1_SUB_88_U175);
  nand ginst6016 (P1_SUB_88_U247, P1_IR_REG_0__SCAN_IN, P1_SUB_88_U174);
  nand ginst6017 (P1_SUB_88_U248, P1_IR_REG_17__SCAN_IN, P1_SUB_88_U34);
  nand ginst6018 (P1_SUB_88_U249, P1_SUB_88_U176, P1_SUB_88_U196);
  and ginst6019 (P1_SUB_88_U25, P1_SUB_88_U183, P1_SUB_88_U186);
  nand ginst6020 (P1_SUB_88_U250, P1_IR_REG_13__SCAN_IN, P1_SUB_88_U35);
  nand ginst6021 (P1_SUB_88_U251, P1_SUB_88_U178, P1_SUB_88_U193);
  and ginst6022 (P1_SUB_88_U26, P1_SUB_88_U185, P1_SUB_88_U28);
  or ginst6023 (P1_SUB_88_U27, P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN);
  nand ginst6024 (P1_SUB_88_U28, P1_SUB_88_U230, P1_SUB_88_U43, P1_SUB_88_U44);
  nand ginst6025 (P1_SUB_88_U29, P1_SUB_88_U230, P1_SUB_88_U45);
  nand ginst6026 (P1_SUB_88_U30, P1_SUB_88_U181, P1_SUB_88_U46);
  not ginst6027 (P1_SUB_88_U31, P1_IR_REG_7__SCAN_IN);
  not ginst6028 (P1_SUB_88_U32, P1_IR_REG_3__SCAN_IN);
  nand ginst6029 (P1_SUB_88_U33, P1_SUB_88_U51, P1_SUB_88_U56);
  nand ginst6030 (P1_SUB_88_U34, P1_SUB_88_U127, P1_SUB_88_U128, P1_SUB_88_U129, P1_SUB_88_U130);
  nand ginst6031 (P1_SUB_88_U35, P1_SUB_88_U156, P1_SUB_88_U184);
  nand ginst6032 (P1_SUB_88_U36, P1_SUB_88_U157, P1_SUB_88_U193);
  not ginst6033 (P1_SUB_88_U37, P1_IR_REG_15__SCAN_IN);
  nand ginst6034 (P1_SUB_88_U38, P1_SUB_88_U158, P1_SUB_88_U184);
  not ginst6035 (P1_SUB_88_U39, P1_IR_REG_11__SCAN_IN);
  nand ginst6036 (P1_SUB_88_U40, P1_SUB_88_U246, P1_SUB_88_U247);
  nand ginst6037 (P1_SUB_88_U41, P1_SUB_88_U236, P1_SUB_88_U237);
  nand ginst6038 (P1_SUB_88_U42, P1_SUB_88_U240, P1_SUB_88_U241);
  nor ginst6039 (P1_SUB_88_U43, P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN);
  nor ginst6040 (P1_SUB_88_U44, P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN);
  nor ginst6041 (P1_SUB_88_U45, P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN);
  nor ginst6042 (P1_SUB_88_U46, P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN);
  nor ginst6043 (P1_SUB_88_U47, P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN);
  nor ginst6044 (P1_SUB_88_U48, P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN);
  nor ginst6045 (P1_SUB_88_U49, P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN, P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN);
  nor ginst6046 (P1_SUB_88_U50, P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN);
  and ginst6047 (P1_SUB_88_U51, P1_SUB_88_U47, P1_SUB_88_U48, P1_SUB_88_U49, P1_SUB_88_U50);
  nor ginst6048 (P1_SUB_88_U52, P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN);
  nor ginst6049 (P1_SUB_88_U53, P1_IR_REG_2__SCAN_IN, P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN);
  nor ginst6050 (P1_SUB_88_U54, P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN);
  nor ginst6051 (P1_SUB_88_U55, P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN);
  and ginst6052 (P1_SUB_88_U56, P1_SUB_88_U52, P1_SUB_88_U53, P1_SUB_88_U54, P1_SUB_88_U55);
  nor ginst6053 (P1_SUB_88_U57, P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN);
  nor ginst6054 (P1_SUB_88_U58, P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN);
  nor ginst6055 (P1_SUB_88_U59, P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN, P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN);
  and ginst6056 (P1_SUB_88_U6, P1_SUB_88_U227, P1_SUB_88_U38);
  nor ginst6057 (P1_SUB_88_U60, P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN);
  and ginst6058 (P1_SUB_88_U61, P1_SUB_88_U57, P1_SUB_88_U58, P1_SUB_88_U59, P1_SUB_88_U60);
  nor ginst6059 (P1_SUB_88_U62, P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN);
  nor ginst6060 (P1_SUB_88_U63, P1_IR_REG_2__SCAN_IN, P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN);
  nor ginst6061 (P1_SUB_88_U64, P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN);
  nor ginst6062 (P1_SUB_88_U65, P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN);
  and ginst6063 (P1_SUB_88_U66, P1_SUB_88_U62, P1_SUB_88_U63, P1_SUB_88_U64, P1_SUB_88_U65);
  nor ginst6064 (P1_SUB_88_U67, P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN);
  nor ginst6065 (P1_SUB_88_U68, P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN);
  nor ginst6066 (P1_SUB_88_U69, P1_IR_REG_1__SCAN_IN, P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN);
  and ginst6067 (P1_SUB_88_U7, P1_SUB_88_U192, P1_SUB_88_U225);
  nor ginst6068 (P1_SUB_88_U70, P1_IR_REG_0__SCAN_IN, P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN);
  and ginst6069 (P1_SUB_88_U71, P1_SUB_88_U67, P1_SUB_88_U68, P1_SUB_88_U69, P1_SUB_88_U70);
  nor ginst6070 (P1_SUB_88_U72, P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN);
  nor ginst6071 (P1_SUB_88_U73, P1_IR_REG_2__SCAN_IN, P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN);
  nor ginst6072 (P1_SUB_88_U74, P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN);
  nor ginst6073 (P1_SUB_88_U75, P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN);
  and ginst6074 (P1_SUB_88_U76, P1_SUB_88_U72, P1_SUB_88_U73, P1_SUB_88_U74, P1_SUB_88_U75);
  nor ginst6075 (P1_SUB_88_U77, P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN);
  nor ginst6076 (P1_SUB_88_U78, P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN);
  nor ginst6077 (P1_SUB_88_U79, P1_IR_REG_1__SCAN_IN, P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN);
  and ginst6078 (P1_SUB_88_U8, P1_SUB_88_U224, P1_SUB_88_U35);
  nor ginst6079 (P1_SUB_88_U80, P1_IR_REG_0__SCAN_IN, P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN);
  and ginst6080 (P1_SUB_88_U81, P1_SUB_88_U77, P1_SUB_88_U78, P1_SUB_88_U79, P1_SUB_88_U80);
  nor ginst6081 (P1_SUB_88_U82, P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN);
  nor ginst6082 (P1_SUB_88_U83, P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN, P1_IR_REG_26__SCAN_IN);
  nor ginst6083 (P1_SUB_88_U84, P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN);
  nor ginst6084 (P1_SUB_88_U85, P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN);
  and ginst6085 (P1_SUB_88_U86, P1_SUB_88_U82, P1_SUB_88_U83, P1_SUB_88_U84, P1_SUB_88_U85);
  nor ginst6086 (P1_SUB_88_U87, P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN);
  nor ginst6087 (P1_SUB_88_U88, P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN);
  nor ginst6088 (P1_SUB_88_U89, P1_IR_REG_1__SCAN_IN, P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN);
  and ginst6089 (P1_SUB_88_U9, P1_SUB_88_U223, P1_SUB_88_U36);
  nor ginst6090 (P1_SUB_88_U90, P1_IR_REG_0__SCAN_IN, P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN);
  and ginst6091 (P1_SUB_88_U91, P1_SUB_88_U87, P1_SUB_88_U88, P1_SUB_88_U89, P1_SUB_88_U90);
  nor ginst6092 (P1_SUB_88_U92, P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN);
  nor ginst6093 (P1_SUB_88_U93, P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN, P1_IR_REG_26__SCAN_IN);
  nor ginst6094 (P1_SUB_88_U94, P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN);
  nor ginst6095 (P1_SUB_88_U95, P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN);
  and ginst6096 (P1_SUB_88_U96, P1_SUB_88_U92, P1_SUB_88_U93, P1_SUB_88_U94, P1_SUB_88_U95);
  nor ginst6097 (P1_SUB_88_U97, P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN);
  nor ginst6098 (P1_SUB_88_U98, P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN);
  nor ginst6099 (P1_SUB_88_U99, P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN);
  and ginst6100 (P1_U3014, P1_U3451, P1_U4002);
  and ginst6101 (P1_U3015, P1_U3449, P1_U3455);
  and ginst6102 (P1_U3016, P1_U3600, P1_U3605);
  and ginst6103 (P1_U3017, P1_U3447, P1_U3448);
  and ginst6104 (P1_U3018, P1_U3447, P1_U5808);
  and ginst6105 (P1_U3019, P1_U3448, P1_U5805);
  and ginst6106 (P1_U3020, P1_U5805, P1_U5808);
  and ginst6107 (P1_U3021, P1_U3425, P1_U5412);
  and ginst6108 (P1_U3022, P1_U3425, P1_U3592);
  and ginst6109 (P1_U3023, P1_U3428, P1_U4043);
  and ginst6110 (P1_U3024, P1_U3048, P1_U5793);
  and ginst6111 (P1_U3025, P1_U4030, P1_U5811);
  and ginst6112 (P1_U3026, P1_U3851, P1_U4015);
  and ginst6113 (P1_U3027, P1_R1352_U6, P1_U3437);
  and ginst6114 (P1_U3028, P1_R1352_U6, P1_U3440);
  and ginst6115 (P1_U3029, P1_STATE_REG_SCAN_IN, P1_U3357);
  and ginst6116 (P1_U3030, P1_U4008, P1_U4031);
  and ginst6117 (P1_U3031, P1_U3426, P1_U4031);
  and ginst6118 (P1_U3032, P1_U4003, P1_U4031);
  and ginst6119 (P1_U3033, P1_U4009, P1_U4031);
  and ginst6120 (P1_U3034, P1_U3449, P1_U4030);
  and ginst6121 (P1_U3035, P1_U4015, P1_U5811);
  and ginst6122 (P1_U3036, P1_U3025, P1_U4031);
  and ginst6123 (P1_U3037, P1_U3449, P1_U4015);
  and ginst6124 (P1_U3038, P1_U4923, P1_U5817);
  and ginst6125 (P1_U3039, P1_U3023, P1_U5817);
  and ginst6126 (P1_U3040, P1_U4923, P1_U5811);
  and ginst6127 (P1_U3041, P1_U3023, P1_U5811);
  and ginst6128 (P1_U3042, P1_U3015, P1_U4923);
  and ginst6129 (P1_U3043, P1_U3015, P1_U3023);
  and ginst6130 (P1_U3044, P1_U3022, P1_U3428);
  and ginst6131 (P1_U3045, P1_U3022, P1_U5159);
  and ginst6132 (P1_U3046, P1_U3016, P1_U3606);
  and ginst6133 (P1_U3047, P1_U3452, P1_U3453);
  and ginst6134 (P1_U3048, P1_U3452, P1_U5799);
  and ginst6135 (P1_U3049, P1_U5796, P1_U5802);
  and ginst6136 (P1_U3050, P1_U3850, P1_U5148);
  and ginst6137 (P1_U3051, P1_U3367, P1_U3419);
  and ginst6138 (P1_U3052, P1_U3422, P1_U3879, P1_U5541);
  nand ginst6139 (P1_U3053, P1_U4679, P1_U4680, P1_U4681, P1_U4682);
  nand ginst6140 (P1_U3054, P1_U4698, P1_U4699, P1_U4700, P1_U4701);
  nand ginst6141 (P1_U3055, P1_U4717, P1_U4718, P1_U4719, P1_U4720);
  nand ginst6142 (P1_U3056, P1_U4756, P1_U4757, P1_U4758);
  nand ginst6143 (P1_U3057, P1_U4660, P1_U4661, P1_U4662, P1_U4663);
  nand ginst6144 (P1_U3058, P1_U4641, P1_U4642, P1_U4643, P1_U4644);
  nand ginst6145 (P1_U3059, P1_U4736, P1_U4737, P1_U4738);
  nand ginst6146 (P1_U3060, P1_U4242, P1_U4243, P1_U4244, P1_U4245);
  nand ginst6147 (P1_U3061, P1_U4584, P1_U4585, P1_U4586, P1_U4587);
  nand ginst6148 (P1_U3062, P1_U4356, P1_U4357, P1_U4358, P1_U4359);
  nand ginst6149 (P1_U3063, P1_U4375, P1_U4376, P1_U4377, P1_U4378);
  nand ginst6150 (P1_U3064, P1_U4223, P1_U4224, P1_U4225, P1_U4226);
  nand ginst6151 (P1_U3065, P1_U4622, P1_U4623, P1_U4624, P1_U4625);
  nand ginst6152 (P1_U3066, P1_U4603, P1_U4604, P1_U4605, P1_U4606);
  nand ginst6153 (P1_U3067, P1_U4261, P1_U4262, P1_U4263, P1_U4264);
  nand ginst6154 (P1_U3068, P1_U4199, P1_U4200, P1_U4201, P1_U4202);
  nand ginst6155 (P1_U3069, P1_U4489, P1_U4490, P1_U4491, P1_U4492);
  nand ginst6156 (P1_U3070, P1_U4299, P1_U4300, P1_U4301, P1_U4302);
  nand ginst6157 (P1_U3071, P1_U4280, P1_U4281, P1_U4282, P1_U4283);
  nand ginst6158 (P1_U3072, P1_U4394, P1_U4395, P1_U4396, P1_U4397);
  nand ginst6159 (P1_U3073, P1_U4470, P1_U4471, P1_U4472, P1_U4473);
  nand ginst6160 (P1_U3074, P1_U4451, P1_U4452, P1_U4453, P1_U4454);
  nand ginst6161 (P1_U3075, P1_U4565, P1_U4566, P1_U4567, P1_U4568);
  nand ginst6162 (P1_U3076, P1_U4546, P1_U4547, P1_U4548, P1_U4549);
  nand ginst6163 (P1_U3077, P1_U4204, P1_U4205, P1_U4206, P1_U4207);
  nand ginst6164 (P1_U3078, P1_U4180, P1_U4181, P1_U4182, P1_U4183);
  nand ginst6165 (P1_U3079, P1_U4432, P1_U4433, P1_U4434, P1_U4435);
  nand ginst6166 (P1_U3080, P1_U4413, P1_U4414, P1_U4415, P1_U4416);
  nand ginst6167 (P1_U3081, P1_U4527, P1_U4528, P1_U4529, P1_U4530);
  nand ginst6168 (P1_U3082, P1_U4508, P1_U4509, P1_U4510, P1_U4511);
  nand ginst6169 (P1_U3083, P1_U4337, P1_U4338, P1_U4339, P1_U4340);
  nand ginst6170 (P1_U3084, P1_U4318, P1_U4319, P1_U4320, P1_U4321);
  nand ginst6171 (P1_U3085, P1_STATE_REG_SCAN_IN, P1_U4930);
  not ginst6172 (P1_U3086, P1_STATE_REG_SCAN_IN);
  nand ginst6173 (P1_U3087, P1_U5666, P1_U5667, P1_U5668);
  nand ginst6174 (P1_U3088, P1_U5669, P1_U5670, P1_U5671);
  nand ginst6175 (P1_U3089, P1_U3929, P1_U5678, P1_U5679);
  nand ginst6176 (P1_U3090, P1_U3930, P1_U5682, P1_U5683);
  nand ginst6177 (P1_U3091, P1_U3931, P1_U5686, P1_U5687);
  nand ginst6178 (P1_U3092, P1_U3932, P1_U5690, P1_U5691);
  nand ginst6179 (P1_U3093, P1_U3933, P1_U5694, P1_U5695);
  nand ginst6180 (P1_U3094, P1_U3934, P1_U5698, P1_U5699);
  nand ginst6181 (P1_U3095, P1_U3935, P1_U5702, P1_U5703);
  nand ginst6182 (P1_U3096, P1_U3936, P1_U5706, P1_U5707);
  nand ginst6183 (P1_U3097, P1_U3937, P1_U5710, P1_U5711);
  nand ginst6184 (P1_U3098, P1_U3938, P1_U5714, P1_U5715);
  nand ginst6185 (P1_U3099, P1_U3940, P1_U5722, P1_U5723);
  nand ginst6186 (P1_U3100, P1_U3941, P1_U5726, P1_U5727);
  nand ginst6187 (P1_U3101, P1_U3942, P1_U5730, P1_U5731);
  nand ginst6188 (P1_U3102, P1_U3943, P1_U5734, P1_U5735);
  nand ginst6189 (P1_U3103, P1_U3944, P1_U5738, P1_U5739);
  nand ginst6190 (P1_U3104, P1_U3945, P1_U5742, P1_U5743);
  nand ginst6191 (P1_U3105, P1_U3946, P1_U5746, P1_U5747);
  nand ginst6192 (P1_U3106, P1_U3947, P1_U5750, P1_U5751);
  nand ginst6193 (P1_U3107, P1_U3948, P1_U5754, P1_U5755);
  nand ginst6194 (P1_U3108, P1_U3949, P1_U5758, P1_U5759);
  nand ginst6195 (P1_U3109, P1_U3922, P1_U5643, P1_U5644);
  nand ginst6196 (P1_U3110, P1_U3923, P1_U5647, P1_U5648);
  nand ginst6197 (P1_U3111, P1_U3924, P1_U5652, P1_U5653);
  nand ginst6198 (P1_U3112, P1_U3925, P1_U5656, P1_U5657);
  nand ginst6199 (P1_U3113, P1_U3926, P1_U5660, P1_U5661);
  nand ginst6200 (P1_U3114, P1_U3927, P1_U5664, P1_U5665);
  nand ginst6201 (P1_U3115, P1_U3928, P1_U5674);
  nand ginst6202 (P1_U3116, P1_U3939, P1_U5718);
  nand ginst6203 (P1_U3117, P1_U3950, P1_U5762);
  nand ginst6204 (P1_U3118, P1_U3951, P1_U5766);
  nand ginst6205 (P1_U3119, P1_U3892, P1_U5563);
  nand ginst6206 (P1_U3120, P1_U3893, P1_U5566);
  nand ginst6207 (P1_U3121, P1_U3896, P1_U5571, P1_U5572);
  nand ginst6208 (P1_U3122, P1_U3897, P1_U5574, P1_U5575);
  nand ginst6209 (P1_U3123, P1_U3898, P1_U5577, P1_U5578);
  nand ginst6210 (P1_U3124, P1_U3899, P1_U5580, P1_U5581);
  nand ginst6211 (P1_U3125, P1_U3900, P1_U5583, P1_U5584);
  nand ginst6212 (P1_U3126, P1_U3901, P1_U5586, P1_U5587);
  nand ginst6213 (P1_U3127, P1_U3902, P1_U5589, P1_U5590);
  nand ginst6214 (P1_U3128, P1_U3903, P1_U5592, P1_U5593);
  nand ginst6215 (P1_U3129, P1_U3904, P1_U5595, P1_U5596);
  nand ginst6216 (P1_U3130, P1_U3905, P1_U5598, P1_U5599);
  nand ginst6217 (P1_U3131, P1_U3908, P1_U5604, P1_U5605);
  nand ginst6218 (P1_U3132, P1_U3909, P1_U5607, P1_U5608);
  nand ginst6219 (P1_U3133, P1_U3910, P1_U5610, P1_U5611);
  nand ginst6220 (P1_U3134, P1_U3911, P1_U5613, P1_U5614);
  nand ginst6221 (P1_U3135, P1_U3912, P1_U5616, P1_U5617);
  nand ginst6222 (P1_U3136, P1_U3913, P1_U5619, P1_U5620);
  nand ginst6223 (P1_U3137, P1_U3914, P1_U5622, P1_U5623);
  nand ginst6224 (P1_U3138, P1_U3915, P1_U5625, P1_U5626);
  nand ginst6225 (P1_U3139, P1_U3916, P1_U5628, P1_U5629);
  nand ginst6226 (P1_U3140, P1_U3917, P1_U5631, P1_U5632);
  nand ginst6227 (P1_U3141, P1_U3880, P1_U5545);
  nand ginst6228 (P1_U3142, P1_U3882, P1_U5548);
  nand ginst6229 (P1_U3143, P1_U3884, P1_U5551);
  nand ginst6230 (P1_U3144, P1_U3886, P1_U5554);
  nand ginst6231 (P1_U3145, P1_U3888, P1_U5557);
  nand ginst6232 (P1_U3146, P1_U3890, P1_U5560);
  nand ginst6233 (P1_U3147, P1_U3894, P1_U5569);
  nand ginst6234 (P1_U3148, P1_U3906, P1_U5602);
  nand ginst6235 (P1_U3149, P1_U3918, P1_U5635);
  nand ginst6236 (P1_U3150, P1_U3920, P1_U5638);
  nand ginst6237 (P1_U3151, P1_U3877, P1_U5537);
  nand ginst6238 (P1_U3152, P1_U3014, P1_U5786);
  nand ginst6239 (P1_U3153, P1_U5491, P1_U5492);
  nand ginst6240 (P1_U3154, P1_U5493, P1_U5494);
  nand ginst6241 (P1_U3155, P1_U5495, P1_U5496);
  nand ginst6242 (P1_U3156, P1_U5497, P1_U5498);
  nand ginst6243 (P1_U3157, P1_U5499, P1_U5500);
  nand ginst6244 (P1_U3158, P1_U5501, P1_U5502);
  nand ginst6245 (P1_U3159, P1_U5503, P1_U5504);
  nand ginst6246 (P1_U3160, P1_U5505, P1_U5506);
  nand ginst6247 (P1_U3161, P1_U5507, P1_U5508);
  nand ginst6248 (P1_U3162, P1_U5511, P1_U5512);
  nand ginst6249 (P1_U3163, P1_U5513, P1_U5514);
  nand ginst6250 (P1_U3164, P1_U5515, P1_U5516);
  nand ginst6251 (P1_U3165, P1_U5517, P1_U5518);
  nand ginst6252 (P1_U3166, P1_U5519, P1_U5520);
  nand ginst6253 (P1_U3167, P1_U5521, P1_U5522);
  nand ginst6254 (P1_U3168, P1_U5523, P1_U5524);
  nand ginst6255 (P1_U3169, P1_U5525, P1_U5526);
  nand ginst6256 (P1_U3170, P1_U5527, P1_U5528);
  nand ginst6257 (P1_U3171, P1_U5529, P1_U5530);
  nand ginst6258 (P1_U3172, P1_U5477, P1_U5478);
  nand ginst6259 (P1_U3173, P1_U5479, P1_U5480);
  nand ginst6260 (P1_U3174, P1_U5481, P1_U5482);
  nand ginst6261 (P1_U3175, P1_U5483, P1_U5484);
  nand ginst6262 (P1_U3176, P1_U5485, P1_U5486);
  nand ginst6263 (P1_U3177, P1_U5487, P1_U5488);
  nand ginst6264 (P1_U3178, P1_U5489, P1_U5490);
  nand ginst6265 (P1_U3179, P1_U5509, P1_U5510);
  nand ginst6266 (P1_U3180, P1_U5531, P1_U5532);
  nand ginst6267 (P1_U3181, P1_U3876, P1_U5534);
  nand ginst6268 (P1_U3182, P1_U5432, P1_U5433);
  nand ginst6269 (P1_U3183, P1_U5434, P1_U5435);
  nand ginst6270 (P1_U3184, P1_U5436, P1_U5437);
  nand ginst6271 (P1_U3185, P1_U5438, P1_U5439);
  nand ginst6272 (P1_U3186, P1_U5440, P1_U5441);
  nand ginst6273 (P1_U3187, P1_U5442, P1_U5443);
  nand ginst6274 (P1_U3188, P1_U5444, P1_U5445);
  nand ginst6275 (P1_U3189, P1_U5446, P1_U5447);
  nand ginst6276 (P1_U3190, P1_U5448, P1_U5449);
  nand ginst6277 (P1_U3191, P1_U5452, P1_U5453);
  nand ginst6278 (P1_U3192, P1_U5454, P1_U5455);
  nand ginst6279 (P1_U3193, P1_U5456, P1_U5457);
  nand ginst6280 (P1_U3194, P1_U5458, P1_U5459);
  nand ginst6281 (P1_U3195, P1_U5460, P1_U5461);
  nand ginst6282 (P1_U3196, P1_U5462, P1_U5463);
  nand ginst6283 (P1_U3197, P1_U5464, P1_U5465);
  nand ginst6284 (P1_U3198, P1_U5466, P1_U5467);
  nand ginst6285 (P1_U3199, P1_U5468, P1_U5469);
  nand ginst6286 (P1_U3200, P1_U5470, P1_U5471);
  nand ginst6287 (P1_U3201, P1_U5418, P1_U5419);
  nand ginst6288 (P1_U3202, P1_U5420, P1_U5421);
  nand ginst6289 (P1_U3203, P1_U5422, P1_U5423);
  nand ginst6290 (P1_U3204, P1_U5424, P1_U5425);
  nand ginst6291 (P1_U3205, P1_U5426, P1_U5427);
  nand ginst6292 (P1_U3206, P1_U5428, P1_U5429);
  nand ginst6293 (P1_U3207, P1_U5430, P1_U5431);
  nand ginst6294 (P1_U3208, P1_U5450, P1_U5451);
  nand ginst6295 (P1_U3209, P1_U5472, P1_U5473);
  nand ginst6296 (P1_U3210, P1_U3875, P1_U5474);
  and ginst6297 (P1_U3211, P1_U3425, P1_U5411);
  nand ginst6298 (P1_U3212, P1_U5409, P1_U6284, P1_U6285);
  nand ginst6299 (P1_U3213, P1_U3872, P1_U5402, P1_U5403, P1_U5404);
  nand ginst6300 (P1_U3214, P1_U5393, P1_U5394, P1_U5395, P1_U5396, P1_U5397);
  nand ginst6301 (P1_U3215, P1_U5384, P1_U5385, P1_U5386, P1_U5387, P1_U5388);
  nand ginst6302 (P1_U3216, P1_U5375, P1_U5376, P1_U5377, P1_U5378, P1_U5379);
  nand ginst6303 (P1_U3217, P1_U3871, P1_U5366, P1_U5367, P1_U5368);
  nand ginst6304 (P1_U3218, P1_U3869, P1_U3870, P1_U5358);
  nand ginst6305 (P1_U3219, P1_U5348, P1_U5349, P1_U5350, P1_U5351, P1_U5352);
  nand ginst6306 (P1_U3220, P1_U5339, P1_U5340, P1_U5341, P1_U5342, P1_U5343);
  nand ginst6307 (P1_U3221, P1_U3868, P1_U5330, P1_U5331, P1_U5332);
  nand ginst6308 (P1_U3222, P1_U3866, P1_U3867, P1_U5322);
  nand ginst6309 (P1_U3223, P1_U5312, P1_U5313, P1_U5314, P1_U5315, P1_U5316);
  nand ginst6310 (P1_U3224, P1_U3865, P1_U5303, P1_U5304, P1_U5305);
  nand ginst6311 (P1_U3225, P1_U5294, P1_U5295, P1_U5296, P1_U5297, P1_U5298);
  nand ginst6312 (P1_U3226, P1_U5285, P1_U5286, P1_U5287, P1_U5288, P1_U5289);
  nand ginst6313 (P1_U3227, P1_U3864, P1_U5276, P1_U5277, P1_U5278);
  nand ginst6314 (P1_U3228, P1_U5267, P1_U5268, P1_U5269, P1_U5270, P1_U5271);
  nand ginst6315 (P1_U3229, P1_U5258, P1_U5259, P1_U5260, P1_U5261, P1_U5262);
  nand ginst6316 (P1_U3230, P1_U3862, P1_U3863, P1_U5250);
  nand ginst6317 (P1_U3231, P1_U3861, P1_U5240, P1_U5241, P1_U5242);
  nand ginst6318 (P1_U3232, P1_U3859, P1_U5233);
  nand ginst6319 (P1_U3233, P1_U5223, P1_U5224, P1_U5225, P1_U5226, P1_U5227);
  nand ginst6320 (P1_U3234, P1_U3857, P1_U5214, P1_U5215, P1_U5216);
  nand ginst6321 (P1_U3235, P1_U5205, P1_U5206, P1_U5207, P1_U5208, P1_U5209);
  nand ginst6322 (P1_U3236, P1_U3856, P1_U5196, P1_U5197, P1_U5198);
  nand ginst6323 (P1_U3237, P1_U3854, P1_U3855, P1_U5188);
  nand ginst6324 (P1_U3238, P1_U5178, P1_U5179, P1_U5180, P1_U5181, P1_U5182);
  nand ginst6325 (P1_U3239, P1_U3853, P1_U5169, P1_U5170, P1_U5171);
  nand ginst6326 (P1_U3240, P1_U5160, P1_U5161, P1_U5162, P1_U5163, P1_U5164);
  nand ginst6327 (P1_U3241, P1_U5149, P1_U5150, P1_U5151, P1_U5152, P1_U5153);
  nand ginst6328 (P1_U3242, P1_U3846, P1_U5137);
  nand ginst6329 (P1_U3243, P1_U3830, P1_U3831, P1_U5123);
  nand ginst6330 (P1_U3244, P1_U3828, P1_U3829, P1_U5113);
  nand ginst6331 (P1_U3245, P1_U3825, P1_U3827, P1_U5103);
  nand ginst6332 (P1_U3246, P1_U3823, P1_U3824, P1_U5093);
  nand ginst6333 (P1_U3247, P1_U3820, P1_U3822, P1_U5083);
  nand ginst6334 (P1_U3248, P1_U3818, P1_U3819, P1_U5073);
  nand ginst6335 (P1_U3249, P1_U3816, P1_U3817, P1_U5063);
  nand ginst6336 (P1_U3250, P1_U3814, P1_U3815, P1_U5053);
  nand ginst6337 (P1_U3251, P1_U3812, P1_U3813, P1_U5043);
  nand ginst6338 (P1_U3252, P1_U3810, P1_U3811, P1_U5033);
  nand ginst6339 (P1_U3253, P1_U3808, P1_U3809, P1_U5023);
  nand ginst6340 (P1_U3254, P1_U3806, P1_U3807, P1_U5013);
  nand ginst6341 (P1_U3255, P1_U3804, P1_U3805, P1_U5003);
  nand ginst6342 (P1_U3256, P1_U3802, P1_U3803, P1_U4993);
  nand ginst6343 (P1_U3257, P1_U3800, P1_U3801, P1_U4983);
  nand ginst6344 (P1_U3258, P1_U3798, P1_U3799, P1_U4973);
  nand ginst6345 (P1_U3259, P1_U3796, P1_U3797, P1_U4963);
  nand ginst6346 (P1_U3260, P1_U3794, P1_U3795, P1_U4953);
  nand ginst6347 (P1_U3261, P1_U3792, P1_U3793, P1_U4943);
  nand ginst6348 (P1_U3262, P1_U3790, P1_U3791, P1_U4933);
  nand ginst6349 (P1_U3263, P1_U3989, P1_U4921, P1_U4922);
  nand ginst6350 (P1_U3264, P1_U3988, P1_U4919, P1_U4920);
  nand ginst6351 (P1_U3265, P1_U3784, P1_U3785, P1_U3985, P1_U4912);
  nand ginst6352 (P1_U3266, P1_U3782, P1_U3783, P1_U3984, P1_U4907);
  nand ginst6353 (P1_U3267, P1_U3780, P1_U3781, P1_U3983, P1_U4902);
  nand ginst6354 (P1_U3268, P1_U3778, P1_U3779, P1_U3982, P1_U4897);
  nand ginst6355 (P1_U3269, P1_U3776, P1_U3777, P1_U3981, P1_U4892);
  nand ginst6356 (P1_U3270, P1_U3774, P1_U3775, P1_U3980, P1_U4887);
  nand ginst6357 (P1_U3271, P1_U3772, P1_U3773, P1_U3979, P1_U4882);
  nand ginst6358 (P1_U3272, P1_U3770, P1_U3771, P1_U3978, P1_U4877);
  nand ginst6359 (P1_U3273, P1_U3768, P1_U3769, P1_U3977, P1_U4872);
  nand ginst6360 (P1_U3274, P1_U3766, P1_U3767, P1_U3976, P1_U4867);
  nand ginst6361 (P1_U3275, P1_U3764, P1_U3765, P1_U3975);
  nand ginst6362 (P1_U3276, P1_U3762, P1_U3763, P1_U3974);
  nand ginst6363 (P1_U3277, P1_U3760, P1_U3761, P1_U3973, P1_U4852);
  nand ginst6364 (P1_U3278, P1_U3758, P1_U3759, P1_U3972, P1_U4847);
  nand ginst6365 (P1_U3279, P1_U3756, P1_U3757, P1_U3971);
  nand ginst6366 (P1_U3280, P1_U3754, P1_U3755, P1_U3970);
  nand ginst6367 (P1_U3281, P1_U3752, P1_U3753, P1_U3969);
  nand ginst6368 (P1_U3282, P1_U3750, P1_U3751, P1_U3968);
  nand ginst6369 (P1_U3283, P1_U3748, P1_U3749, P1_U3967, P1_U4822);
  nand ginst6370 (P1_U3284, P1_U3746, P1_U3747, P1_U3966, P1_U4817);
  nand ginst6371 (P1_U3285, P1_U3744, P1_U3745, P1_U3965);
  nand ginst6372 (P1_U3286, P1_U3742, P1_U3743, P1_U3964);
  nand ginst6373 (P1_U3287, P1_U3740, P1_U3741, P1_U3963);
  nand ginst6374 (P1_U3288, P1_U3738, P1_U3739, P1_U3962);
  nand ginst6375 (P1_U3289, P1_U3736, P1_U3737);
  nand ginst6376 (P1_U3290, P1_U3734, P1_U3735);
  nand ginst6377 (P1_U3291, P1_U3732, P1_U3733);
  nand ginst6378 (P1_U3292, P1_U3730, P1_U3731);
  nand ginst6379 (P1_U3293, P1_U3728, P1_U3729);
  and ginst6380 (P1_U3294, P1_D_REG_31__SCAN_IN, P1_U3953);
  and ginst6381 (P1_U3295, P1_D_REG_30__SCAN_IN, P1_U3953);
  and ginst6382 (P1_U3296, P1_D_REG_29__SCAN_IN, P1_U3953);
  and ginst6383 (P1_U3297, P1_D_REG_28__SCAN_IN, P1_U3953);
  and ginst6384 (P1_U3298, P1_D_REG_27__SCAN_IN, P1_U3953);
  and ginst6385 (P1_U3299, P1_D_REG_26__SCAN_IN, P1_U3953);
  and ginst6386 (P1_U3300, P1_D_REG_25__SCAN_IN, P1_U3953);
  and ginst6387 (P1_U3301, P1_D_REG_24__SCAN_IN, P1_U3953);
  and ginst6388 (P1_U3302, P1_D_REG_23__SCAN_IN, P1_U3953);
  and ginst6389 (P1_U3303, P1_D_REG_22__SCAN_IN, P1_U3953);
  and ginst6390 (P1_U3304, P1_D_REG_21__SCAN_IN, P1_U3953);
  and ginst6391 (P1_U3305, P1_D_REG_20__SCAN_IN, P1_U3953);
  and ginst6392 (P1_U3306, P1_D_REG_19__SCAN_IN, P1_U3953);
  and ginst6393 (P1_U3307, P1_D_REG_18__SCAN_IN, P1_U3953);
  and ginst6394 (P1_U3308, P1_D_REG_17__SCAN_IN, P1_U3953);
  and ginst6395 (P1_U3309, P1_D_REG_16__SCAN_IN, P1_U3953);
  and ginst6396 (P1_U3310, P1_D_REG_15__SCAN_IN, P1_U3953);
  and ginst6397 (P1_U3311, P1_D_REG_14__SCAN_IN, P1_U3953);
  and ginst6398 (P1_U3312, P1_D_REG_13__SCAN_IN, P1_U3953);
  and ginst6399 (P1_U3313, P1_D_REG_12__SCAN_IN, P1_U3953);
  and ginst6400 (P1_U3314, P1_D_REG_11__SCAN_IN, P1_U3953);
  and ginst6401 (P1_U3315, P1_D_REG_10__SCAN_IN, P1_U3953);
  and ginst6402 (P1_U3316, P1_D_REG_9__SCAN_IN, P1_U3953);
  and ginst6403 (P1_U3317, P1_D_REG_8__SCAN_IN, P1_U3953);
  and ginst6404 (P1_U3318, P1_D_REG_7__SCAN_IN, P1_U3953);
  and ginst6405 (P1_U3319, P1_D_REG_6__SCAN_IN, P1_U3953);
  and ginst6406 (P1_U3320, P1_D_REG_5__SCAN_IN, P1_U3953);
  and ginst6407 (P1_U3321, P1_D_REG_4__SCAN_IN, P1_U3953);
  and ginst6408 (P1_U3322, P1_D_REG_3__SCAN_IN, P1_U3953);
  and ginst6409 (P1_U3323, P1_D_REG_2__SCAN_IN, P1_U3953);
  nand ginst6410 (P1_U3324, P1_U4141, P1_U4142, P1_U4143);
  nand ginst6411 (P1_U3325, P1_U4138, P1_U4139, P1_U4140);
  nand ginst6412 (P1_U3326, P1_U4135, P1_U4136, P1_U4137);
  nand ginst6413 (P1_U3327, P1_U4132, P1_U4133, P1_U4134);
  nand ginst6414 (P1_U3328, P1_U4129, P1_U4130, P1_U4131);
  nand ginst6415 (P1_U3329, P1_U4126, P1_U4127, P1_U4128);
  nand ginst6416 (P1_U3330, P1_U4123, P1_U4124, P1_U4125);
  nand ginst6417 (P1_U3331, P1_U4120, P1_U4121, P1_U4122);
  nand ginst6418 (P1_U3332, P1_U4117, P1_U4118, P1_U4119);
  nand ginst6419 (P1_U3333, P1_U4114, P1_U4115, P1_U4116);
  nand ginst6420 (P1_U3334, P1_U4111, P1_U4112, P1_U4113);
  nand ginst6421 (P1_U3335, P1_U4108, P1_U4109, P1_U4110);
  nand ginst6422 (P1_U3336, P1_U4105, P1_U4106, P1_U4107);
  nand ginst6423 (P1_U3337, P1_U4102, P1_U4103, P1_U4104);
  nand ginst6424 (P1_U3338, P1_U4099, P1_U4100, P1_U4101);
  nand ginst6425 (P1_U3339, P1_U4096, P1_U4097, P1_U4098);
  nand ginst6426 (P1_U3340, P1_U4093, P1_U4094, P1_U4095);
  nand ginst6427 (P1_U3341, P1_U4090, P1_U4091, P1_U4092);
  nand ginst6428 (P1_U3342, P1_U4087, P1_U4088, P1_U4089);
  nand ginst6429 (P1_U3343, P1_U4084, P1_U4085, P1_U4086);
  nand ginst6430 (P1_U3344, P1_U4081, P1_U4082, P1_U4083);
  nand ginst6431 (P1_U3345, P1_U4078, P1_U4079, P1_U4080);
  nand ginst6432 (P1_U3346, P1_U4075, P1_U4076, P1_U4077);
  nand ginst6433 (P1_U3347, P1_U4072, P1_U4073, P1_U4074);
  nand ginst6434 (P1_U3348, P1_U4069, P1_U4070, P1_U4071);
  nand ginst6435 (P1_U3349, P1_U4066, P1_U4067, P1_U4068);
  nand ginst6436 (P1_U3350, P1_U4063, P1_U4064, P1_U4065);
  nand ginst6437 (P1_U3351, P1_U4060, P1_U4061, P1_U4062);
  nand ginst6438 (P1_U3352, P1_U4057, P1_U4058, P1_U4059);
  nand ginst6439 (P1_U3353, P1_U4054, P1_U4055, P1_U4056);
  nand ginst6440 (P1_U3354, P1_U4051, P1_U4052, P1_U4053);
  nand ginst6441 (P1_U3355, P1_U4048, P1_U4049, P1_U4050);
  nand ginst6442 (P1_U3356, P1_U3986, P1_U4915, P1_U4916, P1_U4917, P1_U4918);
  nand ginst6443 (P1_U3357, P1_STATE_REG_SCAN_IN, P1_U3952);
  nand ginst6444 (P1_U3358, P1_U3443, P1_U5778);
  not ginst6445 (P1_U3359, P1_B_REG_SCAN_IN);
  nand ginst6446 (P1_U3360, P1_U3443, P1_U5782, P1_U5783);
  nand ginst6447 (P1_U3361, P1_U3048, P1_U3451);
  nand ginst6448 (P1_U3362, P1_U3047, P1_U3451);
  nand ginst6449 (P1_U3363, P1_U3453, P1_U5796);
  nand ginst6450 (P1_U3364, P1_U3451, P1_U4042);
  nand ginst6451 (P1_U3365, P1_U3047, P1_U3450);
  nand ginst6452 (P1_U3366, P1_U3450, P1_U4042);
  nand ginst6453 (P1_U3367, P1_U3049, P1_U3451);
  nand ginst6454 (P1_U3368, P1_U4001, P1_U5799);
  nand ginst6455 (P1_U3369, P1_U5796, P1_U5799);
  nand ginst6456 (P1_U3370, P1_U3450, P1_U4044);
  nand ginst6457 (P1_U3371, P1_U4002, P1_U5793);
  nand ginst6458 (P1_U3372, P1_U3450, P1_U3451);
  nand ginst6459 (P1_U3373, P1_U5793, P1_U5799, P1_U5802);
  nand ginst6460 (P1_U3374, P1_U3049, P1_U5793);
  nand ginst6461 (P1_U3375, P1_U3452, P1_U5802);
  nand ginst6462 (P1_U3376, P1_U3593, P1_U3594, P1_U4190, P1_U4191, P1_U4192);
  not ginst6463 (P1_U3377, P1_REG2_REG_0__SCAN_IN);
  nand ginst6464 (P1_U3378, P1_U3608, P1_U3610, P1_U4209, P1_U4210);
  nand ginst6465 (P1_U3379, P1_U3612, P1_U3614, P1_U4228, P1_U4229);
  nand ginst6466 (P1_U3380, P1_U3616, P1_U3618, P1_U4247, P1_U4248);
  nand ginst6467 (P1_U3381, P1_U3620, P1_U3622, P1_U4266, P1_U4267);
  nand ginst6468 (P1_U3382, P1_U3624, P1_U3626, P1_U4285, P1_U4286);
  nand ginst6469 (P1_U3383, P1_U3628, P1_U3630, P1_U4304, P1_U4305);
  nand ginst6470 (P1_U3384, P1_U3632, P1_U3634, P1_U4323, P1_U4324);
  nand ginst6471 (P1_U3385, P1_U3636, P1_U3638, P1_U4342, P1_U4343);
  nand ginst6472 (P1_U3386, P1_U3640, P1_U3642, P1_U4361, P1_U4362);
  nand ginst6473 (P1_U3387, P1_U3644, P1_U3646, P1_U4380, P1_U4381);
  nand ginst6474 (P1_U3388, P1_U3648, P1_U3650, P1_U4399, P1_U4400);
  nand ginst6475 (P1_U3389, P1_U3652, P1_U3654, P1_U4418, P1_U4419);
  nand ginst6476 (P1_U3390, P1_U3656, P1_U3658, P1_U4437, P1_U4438);
  nand ginst6477 (P1_U3391, P1_U3660, P1_U3662, P1_U4456, P1_U4457);
  nand ginst6478 (P1_U3392, P1_U3664, P1_U3666, P1_U4475, P1_U4476);
  nand ginst6479 (P1_U3393, P1_U3668, P1_U3670, P1_U4494, P1_U4495);
  nand ginst6480 (P1_U3394, P1_U3672, P1_U3674, P1_U4513, P1_U4514);
  nand ginst6481 (P1_U3395, P1_U3676, P1_U3678, P1_U4532, P1_U4533);
  nand ginst6482 (P1_U3396, P1_U3680, P1_U3682, P1_U4551, P1_U4552);
  nand ginst6483 (P1_U3397, P1_U3954, U113);
  nand ginst6484 (P1_U3398, P1_U3684, P1_U3686, P1_U4570, P1_U4571);
  nand ginst6485 (P1_U3399, P1_U3954, U112);
  nand ginst6486 (P1_U3400, P1_U3688, P1_U3690, P1_U4589, P1_U4590);
  nand ginst6487 (P1_U3401, P1_U3954, U111);
  nand ginst6488 (P1_U3402, P1_U3692, P1_U3694, P1_U4608, P1_U4609);
  nand ginst6489 (P1_U3403, P1_U3954, U110);
  nand ginst6490 (P1_U3404, P1_U3696, P1_U3698, P1_U4627, P1_U4628);
  nand ginst6491 (P1_U3405, P1_U3954, U109);
  nand ginst6492 (P1_U3406, P1_U3700, P1_U3702, P1_U4646, P1_U4647);
  nand ginst6493 (P1_U3407, P1_U3954, U108);
  nand ginst6494 (P1_U3408, P1_U3704, P1_U3706, P1_U4665, P1_U4666);
  nand ginst6495 (P1_U3409, P1_U3954, U107);
  nand ginst6496 (P1_U3410, P1_U3708, P1_U3710, P1_U4684, P1_U4685);
  nand ginst6497 (P1_U3411, P1_U3954, U106);
  nand ginst6498 (P1_U3412, P1_U3712, P1_U3714, P1_U4703, P1_U4704);
  nand ginst6499 (P1_U3413, P1_U3954, U105);
  nand ginst6500 (P1_U3414, P1_U3716, P1_U3718, P1_U4722, P1_U4723);
  nand ginst6501 (P1_U3415, P1_U3954, U104);
  nand ginst6502 (P1_U3416, P1_U3721, P1_U3723);
  nand ginst6503 (P1_U3417, P1_U3954, U102);
  nand ginst6504 (P1_U3418, P1_U3954, U101);
  nand ginst6505 (P1_U3419, P1_U4041, P1_U5793);
  nand ginst6506 (P1_U3420, P1_U3022, P1_U4767);
  nand ginst6507 (P1_U3421, P1_U3998, P1_U5799);
  nand ginst6508 (P1_U3422, P1_U3048, P1_U3450);
  nand ginst6509 (P1_U3423, P1_U3047, P1_U5793);
  nand ginst6510 (P1_U3424, P1_U3993, P1_U5799);
  nand ginst6511 (P1_U3425, P1_U3441, P1_U3442, P1_U3443);
  nand ginst6512 (P1_U3426, P1_U4010, P1_U4768);
  nand ginst6513 (P1_U3427, P1_STATE_REG_SCAN_IN, P1_U3444);
  nand ginst6514 (P1_U3428, P1_U3429, P1_U4931);
  nand ginst6515 (P1_U3429, P1_U4145, P1_U5786);
  nand ginst6516 (P1_U3430, P1_STATE_REG_SCAN_IN, P1_U4045);
  nand ginst6517 (P1_U3431, P1_U3014, P1_U3015);
  not ginst6518 (P1_U3432, P1_R1375_U9);
  nand ginst6519 (P1_U3433, P1_U3022, P1_U3426);
  nand ginst6520 (P1_U3434, P1_U3016, P1_U3847);
  nand ginst6521 (P1_U3435, P1_U3852, P1_U5143);
  nand ginst6522 (P1_U3436, P1_U5414, P1_U5415);
  nand ginst6523 (P1_U3437, P1_U3362, P1_U3999);
  nand ginst6524 (P1_U3438, P1_U3051, P1_U5536);
  not ginst6525 (P1_U3439, P1_R1352_U6);
  nand ginst6526 (P1_U3440, P1_U3364, P1_U3423);
  nand ginst6527 (P1_U3441, P1_U5773, P1_U5774);
  nand ginst6528 (P1_U3442, P1_U5776, P1_U5777);
  nand ginst6529 (P1_U3443, P1_U5779, P1_U5780);
  nand ginst6530 (P1_U3444, P1_U5784, P1_U5785);
  nand ginst6531 (P1_U3445, P1_U5787, P1_U5788);
  nand ginst6532 (P1_U3446, P1_U5789, P1_U5790);
  nand ginst6533 (P1_U3447, P1_U5803, P1_U5804);
  nand ginst6534 (P1_U3448, P1_U5806, P1_U5807);
  nand ginst6535 (P1_U3449, P1_U5809, P1_U5810);
  nand ginst6536 (P1_U3450, P1_U5800, P1_U5801);
  nand ginst6537 (P1_U3451, P1_U5791, P1_U5792);
  nand ginst6538 (P1_U3452, P1_U5794, P1_U5795);
  nand ginst6539 (P1_U3453, P1_U5797, P1_U5798);
  nand ginst6540 (P1_U3454, P1_U5812, P1_U5813);
  nand ginst6541 (P1_U3455, P1_U5815, P1_U5816);
  nand ginst6542 (P1_U3456, P1_U5818, P1_U5819);
  nand ginst6543 (P1_U3457, P1_U5826, P1_U5827);
  nand ginst6544 (P1_U3458, P1_U5823, P1_U5824);
  nand ginst6545 (P1_U3459, P1_U5829, P1_U5830);
  nand ginst6546 (P1_U3460, P1_U5831, P1_U5832);
  nand ginst6547 (P1_U3461, P1_U5833, P1_U5834);
  nand ginst6548 (P1_U3462, P1_U5836, P1_U5837);
  nand ginst6549 (P1_U3463, P1_U5838, P1_U5839);
  nand ginst6550 (P1_U3464, P1_U5840, P1_U5841);
  nand ginst6551 (P1_U3465, P1_U5843, P1_U5844);
  nand ginst6552 (P1_U3466, P1_U5845, P1_U5846);
  nand ginst6553 (P1_U3467, P1_U5847, P1_U5848);
  nand ginst6554 (P1_U3468, P1_U5850, P1_U5851);
  nand ginst6555 (P1_U3469, P1_U5852, P1_U5853);
  nand ginst6556 (P1_U3470, P1_U5854, P1_U5855);
  nand ginst6557 (P1_U3471, P1_U5857, P1_U5858);
  nand ginst6558 (P1_U3472, P1_U5859, P1_U5860);
  nand ginst6559 (P1_U3473, P1_U5861, P1_U5862);
  nand ginst6560 (P1_U3474, P1_U5864, P1_U5865);
  nand ginst6561 (P1_U3475, P1_U5866, P1_U5867);
  nand ginst6562 (P1_U3476, P1_U5868, P1_U5869);
  nand ginst6563 (P1_U3477, P1_U5871, P1_U5872);
  nand ginst6564 (P1_U3478, P1_U5873, P1_U5874);
  nand ginst6565 (P1_U3479, P1_U5875, P1_U5876);
  nand ginst6566 (P1_U3480, P1_U5878, P1_U5879);
  nand ginst6567 (P1_U3481, P1_U5880, P1_U5881);
  nand ginst6568 (P1_U3482, P1_U5882, P1_U5883);
  nand ginst6569 (P1_U3483, P1_U5885, P1_U5886);
  nand ginst6570 (P1_U3484, P1_U5887, P1_U5888);
  nand ginst6571 (P1_U3485, P1_U5889, P1_U5890);
  nand ginst6572 (P1_U3486, P1_U5892, P1_U5893);
  nand ginst6573 (P1_U3487, P1_U5894, P1_U5895);
  nand ginst6574 (P1_U3488, P1_U5896, P1_U5897);
  nand ginst6575 (P1_U3489, P1_U5899, P1_U5900);
  nand ginst6576 (P1_U3490, P1_U5901, P1_U5902);
  nand ginst6577 (P1_U3491, P1_U5903, P1_U5904);
  nand ginst6578 (P1_U3492, P1_U5906, P1_U5907);
  nand ginst6579 (P1_U3493, P1_U5908, P1_U5909);
  nand ginst6580 (P1_U3494, P1_U5910, P1_U5911);
  nand ginst6581 (P1_U3495, P1_U5913, P1_U5914);
  nand ginst6582 (P1_U3496, P1_U5915, P1_U5916);
  nand ginst6583 (P1_U3497, P1_U5917, P1_U5918);
  nand ginst6584 (P1_U3498, P1_U5920, P1_U5921);
  nand ginst6585 (P1_U3499, P1_U5922, P1_U5923);
  nand ginst6586 (P1_U3500, P1_U5924, P1_U5925);
  nand ginst6587 (P1_U3501, P1_U5927, P1_U5928);
  nand ginst6588 (P1_U3502, P1_U5929, P1_U5930);
  nand ginst6589 (P1_U3503, P1_U5931, P1_U5932);
  nand ginst6590 (P1_U3504, P1_U5934, P1_U5935);
  nand ginst6591 (P1_U3505, P1_U5936, P1_U5937);
  nand ginst6592 (P1_U3506, P1_U5938, P1_U5939);
  nand ginst6593 (P1_U3507, P1_U5941, P1_U5942);
  nand ginst6594 (P1_U3508, P1_U5943, P1_U5944);
  nand ginst6595 (P1_U3509, P1_U5945, P1_U5946);
  nand ginst6596 (P1_U3510, P1_U5948, P1_U5949);
  nand ginst6597 (P1_U3511, P1_U5950, P1_U5951);
  nand ginst6598 (P1_U3512, P1_U5952, P1_U5953);
  nand ginst6599 (P1_U3513, P1_U5955, P1_U5956);
  nand ginst6600 (P1_U3514, P1_U5957, P1_U5958);
  nand ginst6601 (P1_U3515, P1_U5960, P1_U5961);
  nand ginst6602 (P1_U3516, P1_U5962, P1_U5963);
  nand ginst6603 (P1_U3517, P1_U5964, P1_U5965);
  nand ginst6604 (P1_U3518, P1_U5966, P1_U5967);
  nand ginst6605 (P1_U3519, P1_U5968, P1_U5969);
  nand ginst6606 (P1_U3520, P1_U5970, P1_U5971);
  nand ginst6607 (P1_U3521, P1_U5972, P1_U5973);
  nand ginst6608 (P1_U3522, P1_U5974, P1_U5975);
  nand ginst6609 (P1_U3523, P1_U5976, P1_U5977);
  nand ginst6610 (P1_U3524, P1_U5978, P1_U5979);
  nand ginst6611 (P1_U3525, P1_U5980, P1_U5981);
  nand ginst6612 (P1_U3526, P1_U5982, P1_U5983);
  nand ginst6613 (P1_U3527, P1_U5984, P1_U5985);
  nand ginst6614 (P1_U3528, P1_U5986, P1_U5987);
  nand ginst6615 (P1_U3529, P1_U5988, P1_U5989);
  nand ginst6616 (P1_U3530, P1_U5990, P1_U5991);
  nand ginst6617 (P1_U3531, P1_U5992, P1_U5993);
  nand ginst6618 (P1_U3532, P1_U5994, P1_U5995);
  nand ginst6619 (P1_U3533, P1_U5996, P1_U5997);
  nand ginst6620 (P1_U3534, P1_U5998, P1_U5999);
  nand ginst6621 (P1_U3535, P1_U6000, P1_U6001);
  nand ginst6622 (P1_U3536, P1_U6002, P1_U6003);
  nand ginst6623 (P1_U3537, P1_U6004, P1_U6005);
  nand ginst6624 (P1_U3538, P1_U6006, P1_U6007);
  nand ginst6625 (P1_U3539, P1_U6008, P1_U6009);
  nand ginst6626 (P1_U3540, P1_U6010, P1_U6011);
  nand ginst6627 (P1_U3541, P1_U6012, P1_U6013);
  nand ginst6628 (P1_U3542, P1_U6014, P1_U6015);
  nand ginst6629 (P1_U3543, P1_U6016, P1_U6017);
  nand ginst6630 (P1_U3544, P1_U6018, P1_U6019);
  nand ginst6631 (P1_U3545, P1_U6020, P1_U6021);
  nand ginst6632 (P1_U3546, P1_U6022, P1_U6023);
  nand ginst6633 (P1_U3547, P1_U6024, P1_U6025);
  nand ginst6634 (P1_U3548, P1_U6026, P1_U6027);
  nand ginst6635 (P1_U3549, P1_U6028, P1_U6029);
  nand ginst6636 (P1_U3550, P1_U6030, P1_U6031);
  nand ginst6637 (P1_U3551, P1_U6032, P1_U6033);
  nand ginst6638 (P1_U3552, P1_U6034, P1_U6035);
  nand ginst6639 (P1_U3553, P1_U6036, P1_U6037);
  nand ginst6640 (P1_U3554, P1_U6038, P1_U6039);
  nand ginst6641 (P1_U3555, P1_U6040, P1_U6041);
  nand ginst6642 (P1_U3556, P1_U6042, P1_U6043);
  nand ginst6643 (P1_U3557, P1_U6044, P1_U6045);
  nand ginst6644 (P1_U3558, P1_U6046, P1_U6047);
  nand ginst6645 (P1_U3559, P1_U6048, P1_U6049);
  nand ginst6646 (P1_U3560, P1_U6114, P1_U6115);
  nand ginst6647 (P1_U3561, P1_U6116, P1_U6117);
  nand ginst6648 (P1_U3562, P1_U6118, P1_U6119);
  nand ginst6649 (P1_U3563, P1_U6120, P1_U6121);
  nand ginst6650 (P1_U3564, P1_U6122, P1_U6123);
  nand ginst6651 (P1_U3565, P1_U6124, P1_U6125);
  nand ginst6652 (P1_U3566, P1_U6126, P1_U6127);
  nand ginst6653 (P1_U3567, P1_U6128, P1_U6129);
  nand ginst6654 (P1_U3568, P1_U6130, P1_U6131);
  nand ginst6655 (P1_U3569, P1_U6132, P1_U6133);
  nand ginst6656 (P1_U3570, P1_U6134, P1_U6135);
  nand ginst6657 (P1_U3571, P1_U6136, P1_U6137);
  nand ginst6658 (P1_U3572, P1_U6138, P1_U6139);
  nand ginst6659 (P1_U3573, P1_U6140, P1_U6141);
  nand ginst6660 (P1_U3574, P1_U6142, P1_U6143);
  nand ginst6661 (P1_U3575, P1_U6144, P1_U6145);
  nand ginst6662 (P1_U3576, P1_U6146, P1_U6147);
  nand ginst6663 (P1_U3577, P1_U6148, P1_U6149);
  nand ginst6664 (P1_U3578, P1_U6150, P1_U6151);
  nand ginst6665 (P1_U3579, P1_U6152, P1_U6153);
  nand ginst6666 (P1_U3580, P1_U6154, P1_U6155);
  nand ginst6667 (P1_U3581, P1_U6156, P1_U6157);
  nand ginst6668 (P1_U3582, P1_U6158, P1_U6159);
  nand ginst6669 (P1_U3583, P1_U6160, P1_U6161);
  nand ginst6670 (P1_U3584, P1_U6162, P1_U6163);
  nand ginst6671 (P1_U3585, P1_U6164, P1_U6165);
  nand ginst6672 (P1_U3586, P1_U6166, P1_U6167);
  nand ginst6673 (P1_U3587, P1_U6168, P1_U6169);
  nand ginst6674 (P1_U3588, P1_U6170, P1_U6171);
  nand ginst6675 (P1_U3589, P1_U6172, P1_U6173);
  nand ginst6676 (P1_U3590, P1_U6174, P1_U6175);
  nand ginst6677 (P1_U3591, P1_U6176, P1_U6177);
  and ginst6678 (P1_U3592, P1_STATE_REG_SCAN_IN, P1_U5786);
  and ginst6679 (P1_U3593, P1_U4186, P1_U4187);
  and ginst6680 (P1_U3594, P1_U4188, P1_U4189);
  and ginst6681 (P1_U3595, P1_U4195, P1_U4196);
  and ginst6682 (P1_U3596, P1_U4148, P1_U4149, P1_U4150, P1_U4151);
  and ginst6683 (P1_U3597, P1_U4152, P1_U4153, P1_U4154, P1_U4155);
  and ginst6684 (P1_U3598, P1_U4156, P1_U4157, P1_U4158, P1_U4159);
  and ginst6685 (P1_U3599, P1_U4160, P1_U4161, P1_U4162);
  and ginst6686 (P1_U3600, P1_U3596, P1_U3597, P1_U3598, P1_U3599);
  and ginst6687 (P1_U3601, P1_U4163, P1_U4164, P1_U4165, P1_U4166);
  and ginst6688 (P1_U3602, P1_U4167, P1_U4168, P1_U4169, P1_U4170);
  and ginst6689 (P1_U3603, P1_U4171, P1_U4172, P1_U4173, P1_U4174);
  and ginst6690 (P1_U3604, P1_U4175, P1_U4176, P1_U4177);
  and ginst6691 (P1_U3605, P1_U3601, P1_U3602, P1_U3603, P1_U3604);
  and ginst6692 (P1_U3606, P1_U4179, P1_U5825);
  and ginst6693 (P1_U3607, P1_U3022, P1_U5828);
  and ginst6694 (P1_U3608, P1_U4211, P1_U4212);
  and ginst6695 (P1_U3609, P1_U4213, P1_U4214);
  and ginst6696 (P1_U3610, P1_U3609, P1_U4215, P1_U4216);
  and ginst6697 (P1_U3611, P1_U4218, P1_U4219, P1_U4220, P1_U4221);
  and ginst6698 (P1_U3612, P1_U4230, P1_U4231);
  and ginst6699 (P1_U3613, P1_U4232, P1_U4233);
  and ginst6700 (P1_U3614, P1_U3613, P1_U4234, P1_U4235);
  and ginst6701 (P1_U3615, P1_U4237, P1_U4238, P1_U4239, P1_U4240);
  and ginst6702 (P1_U3616, P1_U4249, P1_U4250);
  and ginst6703 (P1_U3617, P1_U4251, P1_U4252);
  and ginst6704 (P1_U3618, P1_U3617, P1_U4253, P1_U4254);
  and ginst6705 (P1_U3619, P1_U4256, P1_U4257, P1_U4258, P1_U4259);
  and ginst6706 (P1_U3620, P1_U4268, P1_U4269);
  and ginst6707 (P1_U3621, P1_U4270, P1_U4271);
  and ginst6708 (P1_U3622, P1_U3621, P1_U4272, P1_U4273);
  and ginst6709 (P1_U3623, P1_U4275, P1_U4276, P1_U4277, P1_U4278);
  and ginst6710 (P1_U3624, P1_U4287, P1_U4288);
  and ginst6711 (P1_U3625, P1_U4289, P1_U4290);
  and ginst6712 (P1_U3626, P1_U3625, P1_U4291, P1_U4292);
  and ginst6713 (P1_U3627, P1_U4294, P1_U4295, P1_U4296, P1_U4297);
  and ginst6714 (P1_U3628, P1_U4306, P1_U4307);
  and ginst6715 (P1_U3629, P1_U4308, P1_U4309);
  and ginst6716 (P1_U3630, P1_U3629, P1_U4310, P1_U4311);
  and ginst6717 (P1_U3631, P1_U4313, P1_U4314, P1_U4315, P1_U4316);
  and ginst6718 (P1_U3632, P1_U4325, P1_U4326);
  and ginst6719 (P1_U3633, P1_U4327, P1_U4328);
  and ginst6720 (P1_U3634, P1_U3633, P1_U4329, P1_U4330);
  and ginst6721 (P1_U3635, P1_U4332, P1_U4333, P1_U4334, P1_U4335);
  and ginst6722 (P1_U3636, P1_U4344, P1_U4345);
  and ginst6723 (P1_U3637, P1_U4346, P1_U4347);
  and ginst6724 (P1_U3638, P1_U3637, P1_U4348, P1_U4349);
  and ginst6725 (P1_U3639, P1_U4351, P1_U4352, P1_U4353, P1_U4354);
  and ginst6726 (P1_U3640, P1_U4363, P1_U4364);
  and ginst6727 (P1_U3641, P1_U4365, P1_U4366);
  and ginst6728 (P1_U3642, P1_U3641, P1_U4367, P1_U4368);
  and ginst6729 (P1_U3643, P1_U4370, P1_U4371, P1_U4372, P1_U4373);
  and ginst6730 (P1_U3644, P1_U4382, P1_U4383);
  and ginst6731 (P1_U3645, P1_U4384, P1_U4385);
  and ginst6732 (P1_U3646, P1_U3645, P1_U4386, P1_U4387);
  and ginst6733 (P1_U3647, P1_U4389, P1_U4390, P1_U4391, P1_U4392);
  and ginst6734 (P1_U3648, P1_U4401, P1_U4402);
  and ginst6735 (P1_U3649, P1_U4403, P1_U4404);
  and ginst6736 (P1_U3650, P1_U3649, P1_U4405, P1_U4406);
  and ginst6737 (P1_U3651, P1_U4408, P1_U4409, P1_U4410, P1_U4411);
  and ginst6738 (P1_U3652, P1_U4420, P1_U4421);
  and ginst6739 (P1_U3653, P1_U4422, P1_U4423);
  and ginst6740 (P1_U3654, P1_U3653, P1_U4424, P1_U4425);
  and ginst6741 (P1_U3655, P1_U4427, P1_U4428, P1_U4429, P1_U4430);
  and ginst6742 (P1_U3656, P1_U4439, P1_U4440);
  and ginst6743 (P1_U3657, P1_U4441, P1_U4442);
  and ginst6744 (P1_U3658, P1_U3657, P1_U4443, P1_U4444);
  and ginst6745 (P1_U3659, P1_U4446, P1_U4447, P1_U4448, P1_U4449);
  and ginst6746 (P1_U3660, P1_U4458, P1_U4459);
  and ginst6747 (P1_U3661, P1_U4460, P1_U4461);
  and ginst6748 (P1_U3662, P1_U3661, P1_U4462, P1_U4463);
  and ginst6749 (P1_U3663, P1_U4465, P1_U4466, P1_U4467, P1_U4468);
  and ginst6750 (P1_U3664, P1_U4477, P1_U4478);
  and ginst6751 (P1_U3665, P1_U4479, P1_U4480);
  and ginst6752 (P1_U3666, P1_U3665, P1_U4481, P1_U4482);
  and ginst6753 (P1_U3667, P1_U4484, P1_U4485, P1_U4486, P1_U4487);
  and ginst6754 (P1_U3668, P1_U4496, P1_U4497);
  and ginst6755 (P1_U3669, P1_U4498, P1_U4499);
  and ginst6756 (P1_U3670, P1_U3669, P1_U4500, P1_U4501);
  and ginst6757 (P1_U3671, P1_U4503, P1_U4504, P1_U4505, P1_U4506);
  and ginst6758 (P1_U3672, P1_U4515, P1_U4516);
  and ginst6759 (P1_U3673, P1_U4517, P1_U4518);
  and ginst6760 (P1_U3674, P1_U3673, P1_U4519, P1_U4520);
  and ginst6761 (P1_U3675, P1_U4522, P1_U4523, P1_U4524, P1_U4525);
  and ginst6762 (P1_U3676, P1_U4534, P1_U4535);
  and ginst6763 (P1_U3677, P1_U4536, P1_U4537);
  and ginst6764 (P1_U3678, P1_U3677, P1_U4538, P1_U4539);
  and ginst6765 (P1_U3679, P1_U4541, P1_U4542, P1_U4543, P1_U4544);
  and ginst6766 (P1_U3680, P1_U4553, P1_U4554);
  and ginst6767 (P1_U3681, P1_U4555, P1_U4556);
  and ginst6768 (P1_U3682, P1_U3681, P1_U4557, P1_U4558);
  and ginst6769 (P1_U3683, P1_U4560, P1_U4561, P1_U4562, P1_U4563);
  and ginst6770 (P1_U3684, P1_U4572, P1_U4573);
  and ginst6771 (P1_U3685, P1_U4574, P1_U4575);
  and ginst6772 (P1_U3686, P1_U3685, P1_U4576, P1_U4577);
  and ginst6773 (P1_U3687, P1_U4579, P1_U4580, P1_U4581, P1_U4582);
  and ginst6774 (P1_U3688, P1_U4591, P1_U4592);
  and ginst6775 (P1_U3689, P1_U4593, P1_U4594);
  and ginst6776 (P1_U3690, P1_U3689, P1_U4595, P1_U4596);
  and ginst6777 (P1_U3691, P1_U4598, P1_U4599, P1_U4600, P1_U4601);
  and ginst6778 (P1_U3692, P1_U4610, P1_U4611);
  and ginst6779 (P1_U3693, P1_U4612, P1_U4613);
  and ginst6780 (P1_U3694, P1_U3693, P1_U4614, P1_U4615);
  and ginst6781 (P1_U3695, P1_U4617, P1_U4618, P1_U4619, P1_U4620);
  and ginst6782 (P1_U3696, P1_U4629, P1_U4630);
  and ginst6783 (P1_U3697, P1_U4631, P1_U4632);
  and ginst6784 (P1_U3698, P1_U3697, P1_U4633, P1_U4634);
  and ginst6785 (P1_U3699, P1_U4636, P1_U4637, P1_U4638, P1_U4639);
  and ginst6786 (P1_U3700, P1_U4648, P1_U4649);
  and ginst6787 (P1_U3701, P1_U4650, P1_U4651);
  and ginst6788 (P1_U3702, P1_U3701, P1_U4652, P1_U4653);
  and ginst6789 (P1_U3703, P1_U4655, P1_U4656, P1_U4657, P1_U4658);
  and ginst6790 (P1_U3704, P1_U4667, P1_U4668);
  and ginst6791 (P1_U3705, P1_U4669, P1_U4670);
  and ginst6792 (P1_U3706, P1_U3705, P1_U4671, P1_U4672);
  and ginst6793 (P1_U3707, P1_U4674, P1_U4675, P1_U4676, P1_U4677);
  and ginst6794 (P1_U3708, P1_U4686, P1_U4687);
  and ginst6795 (P1_U3709, P1_U4688, P1_U4689);
  and ginst6796 (P1_U3710, P1_U3709, P1_U4690, P1_U4691);
  and ginst6797 (P1_U3711, P1_U4693, P1_U4694, P1_U4695, P1_U4696);
  and ginst6798 (P1_U3712, P1_U4705, P1_U4706);
  and ginst6799 (P1_U3713, P1_U4707, P1_U4708);
  and ginst6800 (P1_U3714, P1_U3713, P1_U4709, P1_U4710);
  and ginst6801 (P1_U3715, P1_U4712, P1_U4713, P1_U4714, P1_U4715);
  and ginst6802 (P1_U3716, P1_U4724, P1_U4725);
  and ginst6803 (P1_U3717, P1_U4726, P1_U4727);
  and ginst6804 (P1_U3718, P1_U3717, P1_U4728, P1_U4729);
  and ginst6805 (P1_U3719, P1_U4731, P1_U4732, P1_U4733, P1_U4734);
  and ginst6806 (P1_U3720, P1_U4030, P1_U4741);
  and ginst6807 (P1_U3721, P1_U4742, P1_U4743, P1_U4744, P1_U4745, P1_U4746);
  and ginst6808 (P1_U3722, P1_U4747, P1_U4748);
  and ginst6809 (P1_U3723, P1_U3722, P1_U4749, P1_U4750);
  and ginst6810 (P1_U3724, P1_U4752, P1_U4753, P1_U4754);
  and ginst6811 (P1_U3725, P1_U4030, P1_U4741);
  and ginst6812 (P1_U3726, P1_U3022, P1_U3457);
  and ginst6813 (P1_U3727, P1_U3458, P1_U4012, P1_U5828);
  and ginst6814 (P1_U3728, P1_U4770, P1_U4771, P1_U4772);
  and ginst6815 (P1_U3729, P1_U3957, P1_U4773, P1_U4774);
  and ginst6816 (P1_U3730, P1_U4775, P1_U4776, P1_U4777);
  and ginst6817 (P1_U3731, P1_U3958, P1_U4778, P1_U4779);
  and ginst6818 (P1_U3732, P1_U4780, P1_U4781, P1_U4782);
  and ginst6819 (P1_U3733, P1_U3959, P1_U4783, P1_U4784);
  and ginst6820 (P1_U3734, P1_U4785, P1_U4786, P1_U4787);
  and ginst6821 (P1_U3735, P1_U3960, P1_U4788, P1_U4789);
  and ginst6822 (P1_U3736, P1_U4790, P1_U4791, P1_U4792);
  and ginst6823 (P1_U3737, P1_U3961, P1_U4793, P1_U4794);
  and ginst6824 (P1_U3738, P1_U4795, P1_U4796, P1_U4797);
  and ginst6825 (P1_U3739, P1_U4798, P1_U4799);
  and ginst6826 (P1_U3740, P1_U4800, P1_U4801, P1_U4802);
  and ginst6827 (P1_U3741, P1_U4803, P1_U4804);
  and ginst6828 (P1_U3742, P1_U4805, P1_U4806, P1_U4807);
  and ginst6829 (P1_U3743, P1_U4808, P1_U4809);
  and ginst6830 (P1_U3744, P1_U4810, P1_U4811, P1_U4812);
  and ginst6831 (P1_U3745, P1_U4813, P1_U4814);
  and ginst6832 (P1_U3746, P1_U4815, P1_U4816);
  and ginst6833 (P1_U3747, P1_U4818, P1_U4819);
  and ginst6834 (P1_U3748, P1_U4820, P1_U4821);
  and ginst6835 (P1_U3749, P1_U4823, P1_U4824);
  and ginst6836 (P1_U3750, P1_U4825, P1_U4826, P1_U4827);
  and ginst6837 (P1_U3751, P1_U4828, P1_U4829);
  and ginst6838 (P1_U3752, P1_U4830, P1_U4831, P1_U4832);
  and ginst6839 (P1_U3753, P1_U4833, P1_U4834);
  and ginst6840 (P1_U3754, P1_U4835, P1_U4836, P1_U4837);
  and ginst6841 (P1_U3755, P1_U4838, P1_U4839);
  and ginst6842 (P1_U3756, P1_U4840, P1_U4841, P1_U4842);
  and ginst6843 (P1_U3757, P1_U4843, P1_U4844);
  and ginst6844 (P1_U3758, P1_U4845, P1_U4846);
  and ginst6845 (P1_U3759, P1_U4848, P1_U4849);
  and ginst6846 (P1_U3760, P1_U4850, P1_U4851);
  and ginst6847 (P1_U3761, P1_U4853, P1_U4854);
  and ginst6848 (P1_U3762, P1_U4855, P1_U4856, P1_U4857);
  and ginst6849 (P1_U3763, P1_U4858, P1_U4859);
  and ginst6850 (P1_U3764, P1_U4860, P1_U4861, P1_U4862);
  and ginst6851 (P1_U3765, P1_U4863, P1_U4864);
  and ginst6852 (P1_U3766, P1_U4865, P1_U4866);
  and ginst6853 (P1_U3767, P1_U4868, P1_U4869);
  and ginst6854 (P1_U3768, P1_U4870, P1_U4871);
  and ginst6855 (P1_U3769, P1_U4873, P1_U4874);
  and ginst6856 (P1_U3770, P1_U4875, P1_U4876);
  and ginst6857 (P1_U3771, P1_U4878, P1_U4879);
  and ginst6858 (P1_U3772, P1_U4880, P1_U4881);
  and ginst6859 (P1_U3773, P1_U4883, P1_U4884);
  and ginst6860 (P1_U3774, P1_U4885, P1_U4886);
  and ginst6861 (P1_U3775, P1_U4888, P1_U4889);
  and ginst6862 (P1_U3776, P1_U4890, P1_U4891);
  and ginst6863 (P1_U3777, P1_U4893, P1_U4894);
  and ginst6864 (P1_U3778, P1_U4895, P1_U4896);
  and ginst6865 (P1_U3779, P1_U4898, P1_U4899);
  and ginst6866 (P1_U3780, P1_U4900, P1_U4901);
  and ginst6867 (P1_U3781, P1_U4903, P1_U4904);
  and ginst6868 (P1_U3782, P1_U4905, P1_U4906);
  and ginst6869 (P1_U3783, P1_U4908, P1_U4909);
  and ginst6870 (P1_U3784, P1_U4910, P1_U4911);
  and ginst6871 (P1_U3785, P1_U4913, P1_U4914);
  and ginst6872 (P1_U3786, P1_U3362, P1_U3364, P1_U3370);
  and ginst6873 (P1_U3787, P1_U3365, P1_U3366, P1_U3422);
  and ginst6874 (P1_U3788, P1_U3361, P1_U4006);
  and ginst6875 (P1_U3789, P1_U3424, P1_U3788);
  and ginst6876 (P1_U3790, P1_U4934, P1_U4935);
  and ginst6877 (P1_U3791, P1_U4936, P1_U4937, P1_U4938);
  and ginst6878 (P1_U3792, P1_U4944, P1_U4945);
  and ginst6879 (P1_U3793, P1_U4946, P1_U4947, P1_U4948);
  and ginst6880 (P1_U3794, P1_U4954, P1_U4955);
  and ginst6881 (P1_U3795, P1_U4956, P1_U4957, P1_U4958);
  and ginst6882 (P1_U3796, P1_U4964, P1_U4965);
  and ginst6883 (P1_U3797, P1_U4966, P1_U4967, P1_U4968);
  and ginst6884 (P1_U3798, P1_U4974, P1_U4975);
  and ginst6885 (P1_U3799, P1_U4976, P1_U4977, P1_U4978);
  and ginst6886 (P1_U3800, P1_U4984, P1_U4985);
  and ginst6887 (P1_U3801, P1_U4986, P1_U4987, P1_U4988);
  and ginst6888 (P1_U3802, P1_U4994, P1_U4995);
  and ginst6889 (P1_U3803, P1_U4996, P1_U4997, P1_U4998);
  and ginst6890 (P1_U3804, P1_U5004, P1_U5005);
  and ginst6891 (P1_U3805, P1_U5006, P1_U5007, P1_U5008);
  and ginst6892 (P1_U3806, P1_U5014, P1_U5015);
  and ginst6893 (P1_U3807, P1_U5016, P1_U5017, P1_U5018);
  and ginst6894 (P1_U3808, P1_U5024, P1_U5025);
  and ginst6895 (P1_U3809, P1_U5026, P1_U5027, P1_U5028);
  and ginst6896 (P1_U3810, P1_U5034, P1_U5035);
  and ginst6897 (P1_U3811, P1_U5036, P1_U5037, P1_U5038);
  and ginst6898 (P1_U3812, P1_U5044, P1_U5045);
  and ginst6899 (P1_U3813, P1_U5046, P1_U5047, P1_U5048);
  and ginst6900 (P1_U3814, P1_U5054, P1_U5055);
  and ginst6901 (P1_U3815, P1_U5056, P1_U5057, P1_U5058);
  and ginst6902 (P1_U3816, P1_U5064, P1_U5065);
  and ginst6903 (P1_U3817, P1_U5066, P1_U5067, P1_U5068);
  and ginst6904 (P1_U3818, P1_U5074, P1_U5075);
  and ginst6905 (P1_U3819, P1_U5076, P1_U5077, P1_U5078);
  and ginst6906 (P1_U3820, P1_U3821, P1_U5084);
  and ginst6907 (P1_U3821, P1_U4040, P1_U5085);
  and ginst6908 (P1_U3822, P1_U5086, P1_U5087, P1_U5088);
  and ginst6909 (P1_U3823, P1_U5094, P1_U5095);
  and ginst6910 (P1_U3824, P1_U5096, P1_U5097, P1_U5098);
  and ginst6911 (P1_U3825, P1_U3826, P1_U5104);
  and ginst6912 (P1_U3826, P1_U4040, P1_U5105);
  and ginst6913 (P1_U3827, P1_U5106, P1_U5107, P1_U5108);
  and ginst6914 (P1_U3828, P1_U5114, P1_U5115);
  and ginst6915 (P1_U3829, P1_U5116, P1_U5117, P1_U5118);
  and ginst6916 (P1_U3830, P1_U5124, P1_U5125);
  and ginst6917 (P1_U3831, P1_U5126, P1_U5127, P1_U5128);
  and ginst6918 (P1_U3832, P1_U6215, P1_U6218, P1_U6221);
  and ginst6919 (P1_U3833, P1_U3832, P1_U3834, P1_U6233);
  and ginst6920 (P1_U3834, P1_U6224, P1_U6227, P1_U6230);
  and ginst6921 (P1_U3835, P1_U6239, P1_U6242, P1_U6245);
  and ginst6922 (P1_U3836, P1_U6248, P1_U6251, P1_U6254);
  and ginst6923 (P1_U3837, P1_U3835, P1_U3836, P1_U6236);
  and ginst6924 (P1_U3838, P1_U6185, P1_U6188, P1_U6191);
  and ginst6925 (P1_U3839, P1_U6194, P1_U6197, P1_U6200, P1_U6203, P1_U6206);
  and ginst6926 (P1_U3840, P1_U6260, P1_U6263, P1_U6266, P1_U6269);
  and ginst6927 (P1_U3841, P1_U6272, P1_U6275);
  and ginst6928 (P1_U3842, P1_U3840, P1_U3841);
  and ginst6929 (P1_U3843, P1_U3833, P1_U3837, P1_U6209, P1_U6212, P1_U6257);
  and ginst6930 (P1_U3844, P1_U3838, P1_U3839, P1_U6182);
  and ginst6931 (P1_U3845, P1_STATE_REG_SCAN_IN, P1_U3429);
  and ginst6932 (P1_U3846, P1_U5136, P1_U5138);
  and ginst6933 (P1_U3847, P1_U3457, P1_U3458);
  and ginst6934 (P1_U3848, P1_U3371, P1_U3996, P1_U3997);
  and ginst6935 (P1_U3849, P1_U3368, P1_U3424);
  and ginst6936 (P1_U3850, P1_U3427, P1_U3430);
  and ginst6937 (P1_U3851, P1_U3022, P1_U5145);
  and ginst6938 (P1_U3852, P1_STATE_REG_SCAN_IN, P1_U3425);
  and ginst6939 (P1_U3853, P1_U5172, P1_U5173);
  and ginst6940 (P1_U3854, P1_U5187, P1_U5189);
  and ginst6941 (P1_U3855, P1_U5190, P1_U5191);
  and ginst6942 (P1_U3856, P1_U5199, P1_U5200);
  and ginst6943 (P1_U3857, P1_U5217, P1_U5218);
  and ginst6944 (P1_U3858, P1_U3078, P1_U4037);
  and ginst6945 (P1_U3859, P1_U3860, P1_U5231, P1_U5232);
  and ginst6946 (P1_U3860, P1_U5234, P1_U5235);
  and ginst6947 (P1_U3861, P1_U5243, P1_U5244);
  and ginst6948 (P1_U3862, P1_U5249, P1_U5251);
  and ginst6949 (P1_U3863, P1_U5252, P1_U5253);
  and ginst6950 (P1_U3864, P1_U5279, P1_U5280);
  and ginst6951 (P1_U3865, P1_U5306, P1_U5307);
  and ginst6952 (P1_U3866, P1_U5321, P1_U5323);
  and ginst6953 (P1_U3867, P1_U5324, P1_U5325);
  and ginst6954 (P1_U3868, P1_U5333, P1_U5334);
  and ginst6955 (P1_U3869, P1_U5357, P1_U5359);
  and ginst6956 (P1_U3870, P1_U5360, P1_U5361);
  and ginst6957 (P1_U3871, P1_U5369, P1_U5370);
  and ginst6958 (P1_U3872, P1_U5405, P1_U5406);
  and ginst6959 (P1_U3873, P1_U5793, P1_U5802);
  and ginst6960 (P1_U3874, P1_U3375, P1_U5410);
  and ginst6961 (P1_U3875, P1_U5475, P1_U5476);
  and ginst6962 (P1_U3876, P1_U5533, P1_U5535);
  and ginst6963 (P1_U3877, P1_U3444, P1_U5538);
  and ginst6964 (P1_U3878, P1_U3374, P1_U3997);
  and ginst6965 (P1_U3879, P1_U3371, P1_U3878);
  and ginst6966 (P1_U3880, P1_U3881, P1_U5546);
  and ginst6967 (P1_U3881, P1_U3444, P1_U5544);
  and ginst6968 (P1_U3882, P1_U3883, P1_U5549);
  and ginst6969 (P1_U3883, P1_U3444, P1_U5547);
  and ginst6970 (P1_U3884, P1_U3885, P1_U5552);
  and ginst6971 (P1_U3885, P1_U3444, P1_U5550);
  and ginst6972 (P1_U3886, P1_U3887, P1_U5555);
  and ginst6973 (P1_U3887, P1_U3444, P1_U5553);
  and ginst6974 (P1_U3888, P1_U3889, P1_U5558);
  and ginst6975 (P1_U3889, P1_U3444, P1_U5556);
  and ginst6976 (P1_U3890, P1_U3891, P1_U5561);
  and ginst6977 (P1_U3891, P1_U3444, P1_U5559);
  and ginst6978 (P1_U3892, P1_U5562, P1_U5564);
  and ginst6979 (P1_U3893, P1_U5565, P1_U5567);
  and ginst6980 (P1_U3894, P1_U3895, P1_U5570);
  and ginst6981 (P1_U3895, P1_U3444, P1_U5568);
  and ginst6982 (P1_U3896, P1_U3444, P1_U5573);
  and ginst6983 (P1_U3897, P1_U3444, P1_U5576);
  and ginst6984 (P1_U3898, P1_U3444, P1_U5579);
  and ginst6985 (P1_U3899, P1_U3444, P1_U5582);
  and ginst6986 (P1_U3900, P1_U3444, P1_U5585);
  and ginst6987 (P1_U3901, P1_U3444, P1_U5588);
  and ginst6988 (P1_U3902, P1_U3444, P1_U5591);
  and ginst6989 (P1_U3903, P1_U3444, P1_U5594);
  and ginst6990 (P1_U3904, P1_U3444, P1_U5597);
  and ginst6991 (P1_U3905, P1_U3444, P1_U5600);
  and ginst6992 (P1_U3906, P1_U3907, P1_U5603);
  and ginst6993 (P1_U3907, P1_U3444, P1_U5601);
  and ginst6994 (P1_U3908, P1_U3444, P1_U5606);
  and ginst6995 (P1_U3909, P1_U3444, P1_U5609);
  and ginst6996 (P1_U3910, P1_U3444, P1_U5612);
  and ginst6997 (P1_U3911, P1_U3444, P1_U5615);
  and ginst6998 (P1_U3912, P1_U3444, P1_U5618);
  and ginst6999 (P1_U3913, P1_U3444, P1_U5621);
  and ginst7000 (P1_U3914, P1_U3444, P1_U5624);
  and ginst7001 (P1_U3915, P1_U3444, P1_U5627);
  and ginst7002 (P1_U3916, P1_U3444, P1_U5630);
  and ginst7003 (P1_U3917, P1_U3444, P1_U5633);
  and ginst7004 (P1_U3918, P1_U3919, P1_U5636);
  and ginst7005 (P1_U3919, P1_U3444, P1_U5634);
  and ginst7006 (P1_U3920, P1_U3921, P1_U5639);
  and ginst7007 (P1_U3921, P1_U3444, P1_U5637);
  and ginst7008 (P1_U3922, P1_U5642, P1_U5645);
  and ginst7009 (P1_U3923, P1_U5646, P1_U5649);
  and ginst7010 (P1_U3924, P1_U5650, P1_U5651);
  and ginst7011 (P1_U3925, P1_U5654, P1_U5655);
  and ginst7012 (P1_U3926, P1_U5658, P1_U5659);
  and ginst7013 (P1_U3927, P1_U5662, P1_U5663);
  and ginst7014 (P1_U3928, P1_U5672, P1_U5673, P1_U5675);
  and ginst7015 (P1_U3929, P1_U5676, P1_U5677);
  and ginst7016 (P1_U3930, P1_U5680, P1_U5681);
  and ginst7017 (P1_U3931, P1_U5684, P1_U5685);
  and ginst7018 (P1_U3932, P1_U5688, P1_U5689);
  and ginst7019 (P1_U3933, P1_U5692, P1_U5693);
  and ginst7020 (P1_U3934, P1_U5696, P1_U5697);
  and ginst7021 (P1_U3935, P1_U5700, P1_U5701);
  and ginst7022 (P1_U3936, P1_U5704, P1_U5705);
  and ginst7023 (P1_U3937, P1_U5708, P1_U5709);
  and ginst7024 (P1_U3938, P1_U5712, P1_U5713);
  and ginst7025 (P1_U3939, P1_U5716, P1_U5717, P1_U5719);
  and ginst7026 (P1_U3940, P1_U5720, P1_U5721);
  and ginst7027 (P1_U3941, P1_U5724, P1_U5725);
  and ginst7028 (P1_U3942, P1_U5728, P1_U5729);
  and ginst7029 (P1_U3943, P1_U5732, P1_U5733);
  and ginst7030 (P1_U3944, P1_U5736, P1_U5737);
  and ginst7031 (P1_U3945, P1_U5740, P1_U5741);
  and ginst7032 (P1_U3946, P1_U5744, P1_U5745);
  and ginst7033 (P1_U3947, P1_U5748, P1_U5749);
  and ginst7034 (P1_U3948, P1_U5752, P1_U5753);
  and ginst7035 (P1_U3949, P1_U5756, P1_U5757);
  and ginst7036 (P1_U3950, P1_U5760, P1_U5761, P1_U5763);
  and ginst7037 (P1_U3951, P1_U5764, P1_U5765);
  not ginst7038 (P1_U3952, P1_IR_REG_31__SCAN_IN);
  nand ginst7039 (P1_U3953, P1_U3022, P1_U3360);
  nand ginst7040 (P1_U3954, P1_U5811, P1_U5817);
  nand ginst7041 (P1_U3955, P1_U3046, P1_U3607);
  nand ginst7042 (P1_U3956, P1_U3046, P1_U3726);
  and ginst7043 (P1_U3957, P1_U6050, P1_U6051);
  and ginst7044 (P1_U3958, P1_U6052, P1_U6053);
  and ginst7045 (P1_U3959, P1_U6054, P1_U6055);
  and ginst7046 (P1_U3960, P1_U6056, P1_U6057);
  and ginst7047 (P1_U3961, P1_U6058, P1_U6059);
  and ginst7048 (P1_U3962, P1_U6060, P1_U6061);
  and ginst7049 (P1_U3963, P1_U6062, P1_U6063);
  and ginst7050 (P1_U3964, P1_U6064, P1_U6065);
  and ginst7051 (P1_U3965, P1_U6066, P1_U6067);
  and ginst7052 (P1_U3966, P1_U6068, P1_U6069);
  and ginst7053 (P1_U3967, P1_U6070, P1_U6071);
  and ginst7054 (P1_U3968, P1_U6072, P1_U6073);
  and ginst7055 (P1_U3969, P1_U6074, P1_U6075);
  and ginst7056 (P1_U3970, P1_U6076, P1_U6077);
  and ginst7057 (P1_U3971, P1_U6078, P1_U6079);
  and ginst7058 (P1_U3972, P1_U6080, P1_U6081);
  and ginst7059 (P1_U3973, P1_U6082, P1_U6083);
  and ginst7060 (P1_U3974, P1_U6084, P1_U6085);
  and ginst7061 (P1_U3975, P1_U6086, P1_U6087);
  and ginst7062 (P1_U3976, P1_U6088, P1_U6089);
  and ginst7063 (P1_U3977, P1_U6090, P1_U6091);
  and ginst7064 (P1_U3978, P1_U6092, P1_U6093);
  and ginst7065 (P1_U3979, P1_U6094, P1_U6095);
  and ginst7066 (P1_U3980, P1_U6096, P1_U6097);
  and ginst7067 (P1_U3981, P1_U6098, P1_U6099);
  and ginst7068 (P1_U3982, P1_U6100, P1_U6101);
  and ginst7069 (P1_U3983, P1_U6102, P1_U6103);
  and ginst7070 (P1_U3984, P1_U6104, P1_U6105);
  and ginst7071 (P1_U3985, P1_U6106, P1_U6107);
  and ginst7072 (P1_U3986, P1_U6108, P1_U6109);
  nand ginst7073 (P1_U3987, P1_U3056, P1_U3725);
  and ginst7074 (P1_U3988, P1_U6110, P1_U6111);
  and ginst7075 (P1_U3989, P1_U6112, P1_U6113);
  and ginst7076 (P1_U3990, P1_U6178, P1_U6179);
  nand ginst7077 (P1_U3991, P1_U3842, P1_U3843, P1_U3844);
  not ginst7078 (P1_U3992, P1_U3371);
  not ginst7079 (P1_U3993, P1_U3374);
  not ginst7080 (P1_U3994, P1_U3364);
  not ginst7081 (P1_U3995, P1_U3423);
  nand ginst7082 (P1_U3996, P1_U4003, P1_U5793);
  nand ginst7083 (P1_U3997, P1_U3451, P1_U4041);
  not ginst7084 (P1_U3998, P1_U3419);
  nand ginst7085 (P1_U3999, P1_U4042, P1_U5793);
  not ginst7086 (P1_U4000, P1_U3362);
  not ginst7087 (P1_U4001, P1_U3367);
  not ginst7088 (P1_U4002, P1_U3370);
  not ginst7089 (P1_U4003, P1_U3422);
  not ginst7090 (P1_U4004, P1_U3366);
  not ginst7091 (P1_U4005, P1_U3365);
  nand ginst7092 (P1_U4006, P1_U3451, P1_U4044);
  not ginst7093 (P1_U4007, P1_U3361);
  not ginst7094 (P1_U4008, P1_U3424);
  not ginst7095 (P1_U4009, P1_U3421);
  nand ginst7096 (P1_U4010, P1_U3453, P1_U3993);
  not ginst7097 (P1_U4011, P1_U3368);
  nand ginst7098 (P1_U4012, P1_U3369, P1_U4030);
  nand ginst7099 (P1_U4013, P1_U3425, P1_U3873);
  not ginst7100 (P1_U4014, P1_U3954);
  not ginst7101 (P1_U4015, P1_U3434);
  not ginst7102 (P1_U4016, P1_U3430);
  not ginst7103 (P1_U4017, P1_U3413);
  not ginst7104 (P1_U4018, P1_U3411);
  not ginst7105 (P1_U4019, P1_U3409);
  not ginst7106 (P1_U4020, P1_U3407);
  not ginst7107 (P1_U4021, P1_U3405);
  not ginst7108 (P1_U4022, P1_U3403);
  not ginst7109 (P1_U4023, P1_U3401);
  not ginst7110 (P1_U4024, P1_U3399);
  not ginst7111 (P1_U4025, P1_U3397);
  not ginst7112 (P1_U4026, P1_U3418);
  not ginst7113 (P1_U4027, P1_U3417);
  not ginst7114 (P1_U4028, P1_U3415);
  not ginst7115 (P1_U4029, P1_U3431);
  not ginst7116 (P1_U4030, P1_U3372);
  not ginst7117 (P1_U4031, P1_U3420);
  not ginst7118 (P1_U4032, P1_U3956);
  not ginst7119 (P1_U4033, P1_U3955);
  not ginst7120 (P1_U4034, P1_U3953);
  not ginst7121 (P1_U4035, P1_U3987);
  not ginst7122 (P1_U4036, P1_U3373);
  not ginst7123 (P1_U4037, P1_U3435);
  not ginst7124 (P1_U4038, P1_U3433);
  nand ginst7125 (P1_U4039, P1_U3022, P1_U4009);
  nand ginst7126 (P1_U4040, P1_U3212, P1_U4016);
  not ginst7127 (P1_U4041, P1_U3375);
  not ginst7128 (P1_U4042, P1_U3363);
  not ginst7129 (P1_U4043, P1_U3427);
  not ginst7130 (P1_U4044, P1_U3369);
  not ginst7131 (P1_U4045, P1_U3429);
  not ginst7132 (P1_U4046, P1_U3358);
  not ginst7133 (P1_U4047, P1_U3357);
  nand ginst7134 (P1_U4048, P1_U3086, U125);
  nand ginst7135 (P1_U4049, P1_IR_REG_0__SCAN_IN, P1_U3029);
  nand ginst7136 (P1_U4050, P1_IR_REG_0__SCAN_IN, P1_U4047);
  nand ginst7137 (P1_U4051, P1_U3086, U114);
  nand ginst7138 (P1_U4052, P1_SUB_88_U40, P1_U3029);
  nand ginst7139 (P1_U4053, P1_IR_REG_1__SCAN_IN, P1_U4047);
  nand ginst7140 (P1_U4054, P1_U3086, U103);
  nand ginst7141 (P1_U4055, P1_SUB_88_U21, P1_U3029);
  nand ginst7142 (P1_U4056, P1_IR_REG_2__SCAN_IN, P1_U4047);
  nand ginst7143 (P1_U4057, P1_U3086, U100);
  nand ginst7144 (P1_U4058, P1_SUB_88_U22, P1_U3029);
  nand ginst7145 (P1_U4059, P1_IR_REG_3__SCAN_IN, P1_U4047);
  nand ginst7146 (P1_U4060, P1_U3086, U99);
  nand ginst7147 (P1_U4061, P1_SUB_88_U23, P1_U3029);
  nand ginst7148 (P1_U4062, P1_IR_REG_4__SCAN_IN, P1_U4047);
  nand ginst7149 (P1_U4063, P1_U3086, U98);
  nand ginst7150 (P1_U4064, P1_SUB_88_U162, P1_U3029);
  nand ginst7151 (P1_U4065, P1_IR_REG_5__SCAN_IN, P1_U4047);
  nand ginst7152 (P1_U4066, P1_U3086, U97);
  nand ginst7153 (P1_U4067, P1_SUB_88_U24, P1_U3029);
  nand ginst7154 (P1_U4068, P1_IR_REG_6__SCAN_IN, P1_U4047);
  nand ginst7155 (P1_U4069, P1_U3086, U96);
  nand ginst7156 (P1_U4070, P1_SUB_88_U25, P1_U3029);
  nand ginst7157 (P1_U4071, P1_IR_REG_7__SCAN_IN, P1_U4047);
  nand ginst7158 (P1_U4072, P1_U3086, U95);
  nand ginst7159 (P1_U4073, P1_SUB_88_U26, P1_U3029);
  nand ginst7160 (P1_U4074, P1_IR_REG_8__SCAN_IN, P1_U4047);
  nand ginst7161 (P1_U4075, P1_U3086, U94);
  nand ginst7162 (P1_U4076, P1_SUB_88_U160, P1_U3029);
  nand ginst7163 (P1_U4077, P1_IR_REG_9__SCAN_IN, P1_U4047);
  nand ginst7164 (P1_U4078, P1_U3086, U124);
  nand ginst7165 (P1_U4079, P1_SUB_88_U6, P1_U3029);
  nand ginst7166 (P1_U4080, P1_IR_REG_10__SCAN_IN, P1_U4047);
  nand ginst7167 (P1_U4081, P1_U3086, U123);
  nand ginst7168 (P1_U4082, P1_SUB_88_U7, P1_U3029);
  nand ginst7169 (P1_U4083, P1_IR_REG_11__SCAN_IN, P1_U4047);
  nand ginst7170 (P1_U4084, P1_U3086, U122);
  nand ginst7171 (P1_U4085, P1_SUB_88_U8, P1_U3029);
  nand ginst7172 (P1_U4086, P1_IR_REG_12__SCAN_IN, P1_U4047);
  nand ginst7173 (P1_U4087, P1_U3086, U121);
  nand ginst7174 (P1_U4088, P1_SUB_88_U179, P1_U3029);
  nand ginst7175 (P1_U4089, P1_IR_REG_13__SCAN_IN, P1_U4047);
  nand ginst7176 (P1_U4090, P1_U3086, U120);
  nand ginst7177 (P1_U4091, P1_SUB_88_U9, P1_U3029);
  nand ginst7178 (P1_U4092, P1_IR_REG_14__SCAN_IN, P1_U4047);
  nand ginst7179 (P1_U4093, P1_U3086, U119);
  nand ginst7180 (P1_U4094, P1_SUB_88_U10, P1_U3029);
  nand ginst7181 (P1_U4095, P1_IR_REG_15__SCAN_IN, P1_U4047);
  nand ginst7182 (P1_U4096, P1_U3086, U118);
  nand ginst7183 (P1_U4097, P1_SUB_88_U11, P1_U3029);
  nand ginst7184 (P1_U4098, P1_IR_REG_16__SCAN_IN, P1_U4047);
  nand ginst7185 (P1_U4099, P1_U3086, U117);
  nand ginst7186 (P1_U4100, P1_SUB_88_U177, P1_U3029);
  nand ginst7187 (P1_U4101, P1_IR_REG_17__SCAN_IN, P1_U4047);
  nand ginst7188 (P1_U4102, P1_U3086, U116);
  nand ginst7189 (P1_U4103, P1_SUB_88_U12, P1_U3029);
  nand ginst7190 (P1_U4104, P1_IR_REG_18__SCAN_IN, P1_U4047);
  nand ginst7191 (P1_U4105, P1_U3086, U115);
  nand ginst7192 (P1_U4106, P1_SUB_88_U13, P1_U3029);
  nand ginst7193 (P1_U4107, P1_IR_REG_19__SCAN_IN, P1_U4047);
  nand ginst7194 (P1_U4108, P1_U3086, U113);
  nand ginst7195 (P1_U4109, P1_SUB_88_U14, P1_U3029);
  nand ginst7196 (P1_U4110, P1_IR_REG_20__SCAN_IN, P1_U4047);
  nand ginst7197 (P1_U4111, P1_U3086, U112);
  nand ginst7198 (P1_U4112, P1_SUB_88_U173, P1_U3029);
  nand ginst7199 (P1_U4113, P1_IR_REG_21__SCAN_IN, P1_U4047);
  nand ginst7200 (P1_U4114, P1_U3086, U111);
  nand ginst7201 (P1_U4115, P1_SUB_88_U15, P1_U3029);
  nand ginst7202 (P1_U4116, P1_IR_REG_22__SCAN_IN, P1_U4047);
  nand ginst7203 (P1_U4117, P1_U3086, U110);
  nand ginst7204 (P1_U4118, P1_SUB_88_U16, P1_U3029);
  nand ginst7205 (P1_U4119, P1_IR_REG_23__SCAN_IN, P1_U4047);
  nand ginst7206 (P1_U4120, P1_U3086, U109);
  nand ginst7207 (P1_U4121, P1_SUB_88_U17, P1_U3029);
  nand ginst7208 (P1_U4122, P1_IR_REG_24__SCAN_IN, P1_U4047);
  nand ginst7209 (P1_U4123, P1_U3086, U108);
  nand ginst7210 (P1_U4124, P1_SUB_88_U170, P1_U3029);
  nand ginst7211 (P1_U4125, P1_IR_REG_25__SCAN_IN, P1_U4047);
  nand ginst7212 (P1_U4126, P1_U3086, U107);
  nand ginst7213 (P1_U4127, P1_SUB_88_U18, P1_U3029);
  nand ginst7214 (P1_U4128, P1_IR_REG_26__SCAN_IN, P1_U4047);
  nand ginst7215 (P1_U4129, P1_U3086, U106);
  nand ginst7216 (P1_U4130, P1_SUB_88_U42, P1_U3029);
  nand ginst7217 (P1_U4131, P1_IR_REG_27__SCAN_IN, P1_U4047);
  nand ginst7218 (P1_U4132, P1_U3086, U105);
  nand ginst7219 (P1_U4133, P1_SUB_88_U19, P1_U3029);
  nand ginst7220 (P1_U4134, P1_IR_REG_28__SCAN_IN, P1_U4047);
  nand ginst7221 (P1_U4135, P1_U3086, U104);
  nand ginst7222 (P1_U4136, P1_SUB_88_U20, P1_U3029);
  nand ginst7223 (P1_U4137, P1_IR_REG_29__SCAN_IN, P1_U4047);
  nand ginst7224 (P1_U4138, P1_U3086, U102);
  nand ginst7225 (P1_U4139, P1_SUB_88_U165, P1_U3029);
  nand ginst7226 (P1_U4140, P1_IR_REG_30__SCAN_IN, P1_U4047);
  nand ginst7227 (P1_U4141, P1_U3086, U101);
  nand ginst7228 (P1_U4142, P1_SUB_88_U41, P1_U3029);
  nand ginst7229 (P1_U4143, P1_IR_REG_31__SCAN_IN, P1_U4047);
  not ginst7230 (P1_U4144, P1_U3360);
  not ginst7231 (P1_U4145, P1_U3425);
  nand ginst7232 (P1_U4146, P1_U3358, P1_U5775);
  nand ginst7233 (P1_U4147, P1_U3358, P1_U5778);
  nand ginst7234 (P1_U4148, P1_D_REG_10__SCAN_IN, P1_U4144);
  nand ginst7235 (P1_U4149, P1_D_REG_11__SCAN_IN, P1_U4144);
  nand ginst7236 (P1_U4150, P1_D_REG_12__SCAN_IN, P1_U4144);
  nand ginst7237 (P1_U4151, P1_D_REG_13__SCAN_IN, P1_U4144);
  nand ginst7238 (P1_U4152, P1_D_REG_14__SCAN_IN, P1_U4144);
  nand ginst7239 (P1_U4153, P1_D_REG_15__SCAN_IN, P1_U4144);
  nand ginst7240 (P1_U4154, P1_D_REG_16__SCAN_IN, P1_U4144);
  nand ginst7241 (P1_U4155, P1_D_REG_17__SCAN_IN, P1_U4144);
  nand ginst7242 (P1_U4156, P1_D_REG_18__SCAN_IN, P1_U4144);
  nand ginst7243 (P1_U4157, P1_D_REG_19__SCAN_IN, P1_U4144);
  nand ginst7244 (P1_U4158, P1_D_REG_20__SCAN_IN, P1_U4144);
  nand ginst7245 (P1_U4159, P1_D_REG_21__SCAN_IN, P1_U4144);
  nand ginst7246 (P1_U4160, P1_D_REG_22__SCAN_IN, P1_U4144);
  nand ginst7247 (P1_U4161, P1_D_REG_23__SCAN_IN, P1_U4144);
  nand ginst7248 (P1_U4162, P1_D_REG_24__SCAN_IN, P1_U4144);
  nand ginst7249 (P1_U4163, P1_D_REG_25__SCAN_IN, P1_U4144);
  nand ginst7250 (P1_U4164, P1_D_REG_26__SCAN_IN, P1_U4144);
  nand ginst7251 (P1_U4165, P1_D_REG_27__SCAN_IN, P1_U4144);
  nand ginst7252 (P1_U4166, P1_D_REG_28__SCAN_IN, P1_U4144);
  nand ginst7253 (P1_U4167, P1_D_REG_29__SCAN_IN, P1_U4144);
  nand ginst7254 (P1_U4168, P1_D_REG_2__SCAN_IN, P1_U4144);
  nand ginst7255 (P1_U4169, P1_D_REG_30__SCAN_IN, P1_U4144);
  nand ginst7256 (P1_U4170, P1_D_REG_31__SCAN_IN, P1_U4144);
  nand ginst7257 (P1_U4171, P1_D_REG_3__SCAN_IN, P1_U4144);
  nand ginst7258 (P1_U4172, P1_D_REG_4__SCAN_IN, P1_U4144);
  nand ginst7259 (P1_U4173, P1_D_REG_5__SCAN_IN, P1_U4144);
  nand ginst7260 (P1_U4174, P1_D_REG_6__SCAN_IN, P1_U4144);
  nand ginst7261 (P1_U4175, P1_D_REG_7__SCAN_IN, P1_U4144);
  nand ginst7262 (P1_U4176, P1_D_REG_8__SCAN_IN, P1_U4144);
  nand ginst7263 (P1_U4177, P1_D_REG_9__SCAN_IN, P1_U4144);
  nand ginst7264 (P1_U4178, P1_U5799, P1_U5802);
  nand ginst7265 (P1_U4179, P1_U3369, P1_U5821, P1_U5822);
  nand ginst7266 (P1_U4180, P1_REG2_REG_1__SCAN_IN, P1_U3018);
  nand ginst7267 (P1_U4181, P1_REG1_REG_1__SCAN_IN, P1_U3019);
  nand ginst7268 (P1_U4182, P1_REG0_REG_1__SCAN_IN, P1_U3020);
  nand ginst7269 (P1_U4183, P1_REG3_REG_1__SCAN_IN, P1_U3017);
  not ginst7270 (P1_U4184, P1_U3078);
  nand ginst7271 (P1_U4185, P1_U3419, P1_U4010);
  nand ginst7272 (P1_U4186, P1_R1150_U21, P1_U4007);
  nand ginst7273 (P1_U4187, P1_R1117_U21, P1_U4000);
  nand ginst7274 (P1_U4188, P1_R1138_U96, P1_U3994);
  nand ginst7275 (P1_U4189, P1_R1192_U21, P1_U4005);
  nand ginst7276 (P1_U4190, P1_R1207_U21, P1_U4004);
  nand ginst7277 (P1_U4191, P1_R1171_U96, P1_U4011);
  nand ginst7278 (P1_U4192, P1_R1240_U96, P1_U3992);
  not ginst7279 (P1_U4193, P1_U3376);
  nand ginst7280 (P1_U4194, P1_U3025, P1_U3078);
  nand ginst7281 (P1_U4195, P1_R1222_U96, P1_U3024);
  nand ginst7282 (P1_U4196, P1_U3456, P1_U4036);
  nand ginst7283 (P1_U4197, P1_U3456, P1_U4185);
  nand ginst7284 (P1_U4198, P1_U3595, P1_U4193, P1_U4194, P1_U4197);
  nand ginst7285 (P1_U4199, P1_REG2_REG_2__SCAN_IN, P1_U3018);
  nand ginst7286 (P1_U4200, P1_REG1_REG_2__SCAN_IN, P1_U3019);
  nand ginst7287 (P1_U4201, P1_REG0_REG_2__SCAN_IN, P1_U3020);
  nand ginst7288 (P1_U4202, P1_REG3_REG_2__SCAN_IN, P1_U3017);
  not ginst7289 (P1_U4203, P1_U3068);
  nand ginst7290 (P1_U4204, P1_REG0_REG_0__SCAN_IN, P1_U3020);
  nand ginst7291 (P1_U4205, P1_REG1_REG_0__SCAN_IN, P1_U3019);
  nand ginst7292 (P1_U4206, P1_REG2_REG_0__SCAN_IN, P1_U3018);
  nand ginst7293 (P1_U4207, P1_REG3_REG_0__SCAN_IN, P1_U3017);
  not ginst7294 (P1_U4208, P1_U3077);
  nand ginst7295 (P1_U4209, P1_U3034, P1_U3077);
  nand ginst7296 (P1_U4210, P1_R1150_U98, P1_U4007);
  nand ginst7297 (P1_U4211, P1_R1117_U98, P1_U4000);
  nand ginst7298 (P1_U4212, P1_R1138_U95, P1_U3994);
  nand ginst7299 (P1_U4213, P1_R1192_U98, P1_U4005);
  nand ginst7300 (P1_U4214, P1_R1207_U98, P1_U4004);
  nand ginst7301 (P1_U4215, P1_R1171_U95, P1_U4011);
  nand ginst7302 (P1_U4216, P1_R1240_U95, P1_U3992);
  not ginst7303 (P1_U4217, P1_U3378);
  nand ginst7304 (P1_U4218, P1_U3025, P1_U3068);
  nand ginst7305 (P1_U4219, P1_R1222_U95, P1_U3024);
  nand ginst7306 (P1_U4220, P1_R1282_U56, P1_U4036);
  nand ginst7307 (P1_U4221, P1_U3461, P1_U4185);
  nand ginst7308 (P1_U4222, P1_U3611, P1_U4217);
  nand ginst7309 (P1_U4223, P1_REG2_REG_3__SCAN_IN, P1_U3018);
  nand ginst7310 (P1_U4224, P1_REG1_REG_3__SCAN_IN, P1_U3019);
  nand ginst7311 (P1_U4225, P1_REG0_REG_3__SCAN_IN, P1_U3020);
  nand ginst7312 (P1_U4226, P1_ADD_99_U4, P1_U3017);
  not ginst7313 (P1_U4227, P1_U3064);
  nand ginst7314 (P1_U4228, P1_U3034, P1_U3078);
  nand ginst7315 (P1_U4229, P1_R1150_U108, P1_U4007);
  nand ginst7316 (P1_U4230, P1_R1117_U108, P1_U4000);
  nand ginst7317 (P1_U4231, P1_R1138_U17, P1_U3994);
  nand ginst7318 (P1_U4232, P1_R1192_U108, P1_U4005);
  nand ginst7319 (P1_U4233, P1_R1207_U108, P1_U4004);
  nand ginst7320 (P1_U4234, P1_R1171_U17, P1_U4011);
  nand ginst7321 (P1_U4235, P1_R1240_U17, P1_U3992);
  not ginst7322 (P1_U4236, P1_U3379);
  nand ginst7323 (P1_U4237, P1_U3025, P1_U3064);
  nand ginst7324 (P1_U4238, P1_R1222_U17, P1_U3024);
  nand ginst7325 (P1_U4239, P1_R1282_U18, P1_U4036);
  nand ginst7326 (P1_U4240, P1_U3464, P1_U4185);
  nand ginst7327 (P1_U4241, P1_U3615, P1_U4236);
  nand ginst7328 (P1_U4242, P1_REG2_REG_4__SCAN_IN, P1_U3018);
  nand ginst7329 (P1_U4243, P1_REG1_REG_4__SCAN_IN, P1_U3019);
  nand ginst7330 (P1_U4244, P1_REG0_REG_4__SCAN_IN, P1_U3020);
  nand ginst7331 (P1_U4245, P1_ADD_99_U59, P1_U3017);
  not ginst7332 (P1_U4246, P1_U3060);
  nand ginst7333 (P1_U4247, P1_U3034, P1_U3068);
  nand ginst7334 (P1_U4248, P1_R1150_U18, P1_U4007);
  nand ginst7335 (P1_U4249, P1_R1117_U18, P1_U4000);
  nand ginst7336 (P1_U4250, P1_R1138_U101, P1_U3994);
  nand ginst7337 (P1_U4251, P1_R1192_U18, P1_U4005);
  nand ginst7338 (P1_U4252, P1_R1207_U18, P1_U4004);
  nand ginst7339 (P1_U4253, P1_R1171_U101, P1_U4011);
  nand ginst7340 (P1_U4254, P1_R1240_U101, P1_U3992);
  not ginst7341 (P1_U4255, P1_U3380);
  nand ginst7342 (P1_U4256, P1_U3025, P1_U3060);
  nand ginst7343 (P1_U4257, P1_R1222_U101, P1_U3024);
  nand ginst7344 (P1_U4258, P1_R1282_U20, P1_U4036);
  nand ginst7345 (P1_U4259, P1_U3467, P1_U4185);
  nand ginst7346 (P1_U4260, P1_U3619, P1_U4255);
  nand ginst7347 (P1_U4261, P1_REG2_REG_5__SCAN_IN, P1_U3018);
  nand ginst7348 (P1_U4262, P1_REG1_REG_5__SCAN_IN, P1_U3019);
  nand ginst7349 (P1_U4263, P1_REG0_REG_5__SCAN_IN, P1_U3020);
  nand ginst7350 (P1_U4264, P1_ADD_99_U58, P1_U3017);
  not ginst7351 (P1_U4265, P1_U3067);
  nand ginst7352 (P1_U4266, P1_U3034, P1_U3064);
  nand ginst7353 (P1_U4267, P1_R1150_U107, P1_U4007);
  nand ginst7354 (P1_U4268, P1_R1117_U107, P1_U4000);
  nand ginst7355 (P1_U4269, P1_R1138_U100, P1_U3994);
  nand ginst7356 (P1_U4270, P1_R1192_U107, P1_U4005);
  nand ginst7357 (P1_U4271, P1_R1207_U107, P1_U4004);
  nand ginst7358 (P1_U4272, P1_R1171_U100, P1_U4011);
  nand ginst7359 (P1_U4273, P1_R1240_U100, P1_U3992);
  not ginst7360 (P1_U4274, P1_U3381);
  nand ginst7361 (P1_U4275, P1_U3025, P1_U3067);
  nand ginst7362 (P1_U4276, P1_R1222_U100, P1_U3024);
  nand ginst7363 (P1_U4277, P1_R1282_U21, P1_U4036);
  nand ginst7364 (P1_U4278, P1_U3470, P1_U4185);
  nand ginst7365 (P1_U4279, P1_U3623, P1_U4274);
  nand ginst7366 (P1_U4280, P1_REG2_REG_6__SCAN_IN, P1_U3018);
  nand ginst7367 (P1_U4281, P1_REG1_REG_6__SCAN_IN, P1_U3019);
  nand ginst7368 (P1_U4282, P1_REG0_REG_6__SCAN_IN, P1_U3020);
  nand ginst7369 (P1_U4283, P1_ADD_99_U57, P1_U3017);
  not ginst7370 (P1_U4284, P1_U3071);
  nand ginst7371 (P1_U4285, P1_U3034, P1_U3060);
  nand ginst7372 (P1_U4286, P1_R1150_U106, P1_U4007);
  nand ginst7373 (P1_U4287, P1_R1117_U106, P1_U4000);
  nand ginst7374 (P1_U4288, P1_R1138_U18, P1_U3994);
  nand ginst7375 (P1_U4289, P1_R1192_U106, P1_U4005);
  nand ginst7376 (P1_U4290, P1_R1207_U106, P1_U4004);
  nand ginst7377 (P1_U4291, P1_R1171_U18, P1_U4011);
  nand ginst7378 (P1_U4292, P1_R1240_U18, P1_U3992);
  not ginst7379 (P1_U4293, P1_U3382);
  nand ginst7380 (P1_U4294, P1_U3025, P1_U3071);
  nand ginst7381 (P1_U4295, P1_R1222_U18, P1_U3024);
  nand ginst7382 (P1_U4296, P1_R1282_U65, P1_U4036);
  nand ginst7383 (P1_U4297, P1_U3473, P1_U4185);
  nand ginst7384 (P1_U4298, P1_U3627, P1_U4293);
  nand ginst7385 (P1_U4299, P1_REG2_REG_7__SCAN_IN, P1_U3018);
  nand ginst7386 (P1_U4300, P1_REG1_REG_7__SCAN_IN, P1_U3019);
  nand ginst7387 (P1_U4301, P1_REG0_REG_7__SCAN_IN, P1_U3020);
  nand ginst7388 (P1_U4302, P1_ADD_99_U56, P1_U3017);
  not ginst7389 (P1_U4303, P1_U3070);
  nand ginst7390 (P1_U4304, P1_U3034, P1_U3067);
  nand ginst7391 (P1_U4305, P1_R1150_U19, P1_U4007);
  nand ginst7392 (P1_U4306, P1_R1117_U19, P1_U4000);
  nand ginst7393 (P1_U4307, P1_R1138_U99, P1_U3994);
  nand ginst7394 (P1_U4308, P1_R1192_U19, P1_U4005);
  nand ginst7395 (P1_U4309, P1_R1207_U19, P1_U4004);
  nand ginst7396 (P1_U4310, P1_R1171_U99, P1_U4011);
  nand ginst7397 (P1_U4311, P1_R1240_U99, P1_U3992);
  not ginst7398 (P1_U4312, P1_U3383);
  nand ginst7399 (P1_U4313, P1_U3025, P1_U3070);
  nand ginst7400 (P1_U4314, P1_R1222_U99, P1_U3024);
  nand ginst7401 (P1_U4315, P1_R1282_U22, P1_U4036);
  nand ginst7402 (P1_U4316, P1_U3476, P1_U4185);
  nand ginst7403 (P1_U4317, P1_U3631, P1_U4312);
  nand ginst7404 (P1_U4318, P1_REG2_REG_8__SCAN_IN, P1_U3018);
  nand ginst7405 (P1_U4319, P1_REG1_REG_8__SCAN_IN, P1_U3019);
  nand ginst7406 (P1_U4320, P1_REG0_REG_8__SCAN_IN, P1_U3020);
  nand ginst7407 (P1_U4321, P1_ADD_99_U55, P1_U3017);
  not ginst7408 (P1_U4322, P1_U3084);
  nand ginst7409 (P1_U4323, P1_U3034, P1_U3071);
  nand ginst7410 (P1_U4324, P1_R1150_U105, P1_U4007);
  nand ginst7411 (P1_U4325, P1_R1117_U105, P1_U4000);
  nand ginst7412 (P1_U4326, P1_R1138_U19, P1_U3994);
  nand ginst7413 (P1_U4327, P1_R1192_U105, P1_U4005);
  nand ginst7414 (P1_U4328, P1_R1207_U105, P1_U4004);
  nand ginst7415 (P1_U4329, P1_R1171_U19, P1_U4011);
  nand ginst7416 (P1_U4330, P1_R1240_U19, P1_U3992);
  not ginst7417 (P1_U4331, P1_U3384);
  nand ginst7418 (P1_U4332, P1_U3025, P1_U3084);
  nand ginst7419 (P1_U4333, P1_R1222_U19, P1_U3024);
  nand ginst7420 (P1_U4334, P1_R1282_U23, P1_U4036);
  nand ginst7421 (P1_U4335, P1_U3479, P1_U4185);
  nand ginst7422 (P1_U4336, P1_U3635, P1_U4331);
  nand ginst7423 (P1_U4337, P1_REG2_REG_9__SCAN_IN, P1_U3018);
  nand ginst7424 (P1_U4338, P1_REG1_REG_9__SCAN_IN, P1_U3019);
  nand ginst7425 (P1_U4339, P1_REG0_REG_9__SCAN_IN, P1_U3020);
  nand ginst7426 (P1_U4340, P1_ADD_99_U54, P1_U3017);
  not ginst7427 (P1_U4341, P1_U3083);
  nand ginst7428 (P1_U4342, P1_U3034, P1_U3070);
  nand ginst7429 (P1_U4343, P1_R1150_U20, P1_U4007);
  nand ginst7430 (P1_U4344, P1_R1117_U20, P1_U4000);
  nand ginst7431 (P1_U4345, P1_R1138_U98, P1_U3994);
  nand ginst7432 (P1_U4346, P1_R1192_U20, P1_U4005);
  nand ginst7433 (P1_U4347, P1_R1207_U20, P1_U4004);
  nand ginst7434 (P1_U4348, P1_R1171_U98, P1_U4011);
  nand ginst7435 (P1_U4349, P1_R1240_U98, P1_U3992);
  not ginst7436 (P1_U4350, P1_U3385);
  nand ginst7437 (P1_U4351, P1_U3025, P1_U3083);
  nand ginst7438 (P1_U4352, P1_R1222_U98, P1_U3024);
  nand ginst7439 (P1_U4353, P1_R1282_U24, P1_U4036);
  nand ginst7440 (P1_U4354, P1_U3482, P1_U4185);
  nand ginst7441 (P1_U4355, P1_U3639, P1_U4350);
  nand ginst7442 (P1_U4356, P1_REG2_REG_10__SCAN_IN, P1_U3018);
  nand ginst7443 (P1_U4357, P1_REG1_REG_10__SCAN_IN, P1_U3019);
  nand ginst7444 (P1_U4358, P1_REG0_REG_10__SCAN_IN, P1_U3020);
  nand ginst7445 (P1_U4359, P1_ADD_99_U78, P1_U3017);
  not ginst7446 (P1_U4360, P1_U3062);
  nand ginst7447 (P1_U4361, P1_U3034, P1_U3084);
  nand ginst7448 (P1_U4362, P1_R1150_U104, P1_U4007);
  nand ginst7449 (P1_U4363, P1_R1117_U104, P1_U4000);
  nand ginst7450 (P1_U4364, P1_R1138_U97, P1_U3994);
  nand ginst7451 (P1_U4365, P1_R1192_U104, P1_U4005);
  nand ginst7452 (P1_U4366, P1_R1207_U104, P1_U4004);
  nand ginst7453 (P1_U4367, P1_R1171_U97, P1_U4011);
  nand ginst7454 (P1_U4368, P1_R1240_U97, P1_U3992);
  not ginst7455 (P1_U4369, P1_U3386);
  nand ginst7456 (P1_U4370, P1_U3025, P1_U3062);
  nand ginst7457 (P1_U4371, P1_R1222_U97, P1_U3024);
  nand ginst7458 (P1_U4372, P1_R1282_U63, P1_U4036);
  nand ginst7459 (P1_U4373, P1_U3485, P1_U4185);
  nand ginst7460 (P1_U4374, P1_U3643, P1_U4369);
  nand ginst7461 (P1_U4375, P1_REG2_REG_11__SCAN_IN, P1_U3018);
  nand ginst7462 (P1_U4376, P1_REG1_REG_11__SCAN_IN, P1_U3019);
  nand ginst7463 (P1_U4377, P1_REG0_REG_11__SCAN_IN, P1_U3020);
  nand ginst7464 (P1_U4378, P1_ADD_99_U77, P1_U3017);
  not ginst7465 (P1_U4379, P1_U3063);
  nand ginst7466 (P1_U4380, P1_U3034, P1_U3083);
  nand ginst7467 (P1_U4381, P1_R1150_U114, P1_U4007);
  nand ginst7468 (P1_U4382, P1_R1117_U114, P1_U4000);
  nand ginst7469 (P1_U4383, P1_R1138_U11, P1_U3994);
  nand ginst7470 (P1_U4384, P1_R1192_U114, P1_U4005);
  nand ginst7471 (P1_U4385, P1_R1207_U114, P1_U4004);
  nand ginst7472 (P1_U4386, P1_R1171_U11, P1_U4011);
  nand ginst7473 (P1_U4387, P1_R1240_U11, P1_U3992);
  not ginst7474 (P1_U4388, P1_U3387);
  nand ginst7475 (P1_U4389, P1_U3025, P1_U3063);
  nand ginst7476 (P1_U4390, P1_R1222_U11, P1_U3024);
  nand ginst7477 (P1_U4391, P1_R1282_U6, P1_U4036);
  nand ginst7478 (P1_U4392, P1_U3488, P1_U4185);
  nand ginst7479 (P1_U4393, P1_U3647, P1_U4388);
  nand ginst7480 (P1_U4394, P1_REG2_REG_12__SCAN_IN, P1_U3018);
  nand ginst7481 (P1_U4395, P1_REG1_REG_12__SCAN_IN, P1_U3019);
  nand ginst7482 (P1_U4396, P1_REG0_REG_12__SCAN_IN, P1_U3020);
  nand ginst7483 (P1_U4397, P1_ADD_99_U76, P1_U3017);
  not ginst7484 (P1_U4398, P1_U3072);
  nand ginst7485 (P1_U4399, P1_U3034, P1_U3062);
  nand ginst7486 (P1_U4400, P1_R1150_U13, P1_U4007);
  nand ginst7487 (P1_U4401, P1_R1117_U13, P1_U4000);
  nand ginst7488 (P1_U4402, P1_R1138_U115, P1_U3994);
  nand ginst7489 (P1_U4403, P1_R1192_U13, P1_U4005);
  nand ginst7490 (P1_U4404, P1_R1207_U13, P1_U4004);
  nand ginst7491 (P1_U4405, P1_R1171_U115, P1_U4011);
  nand ginst7492 (P1_U4406, P1_R1240_U115, P1_U3992);
  not ginst7493 (P1_U4407, P1_U3388);
  nand ginst7494 (P1_U4408, P1_U3025, P1_U3072);
  nand ginst7495 (P1_U4409, P1_R1222_U115, P1_U3024);
  nand ginst7496 (P1_U4410, P1_R1282_U7, P1_U4036);
  nand ginst7497 (P1_U4411, P1_U3491, P1_U4185);
  nand ginst7498 (P1_U4412, P1_U3651, P1_U4407);
  nand ginst7499 (P1_U4413, P1_REG2_REG_13__SCAN_IN, P1_U3018);
  nand ginst7500 (P1_U4414, P1_REG1_REG_13__SCAN_IN, P1_U3019);
  nand ginst7501 (P1_U4415, P1_REG0_REG_13__SCAN_IN, P1_U3020);
  nand ginst7502 (P1_U4416, P1_ADD_99_U75, P1_U3017);
  not ginst7503 (P1_U4417, P1_U3080);
  nand ginst7504 (P1_U4418, P1_U3034, P1_U3063);
  nand ginst7505 (P1_U4419, P1_R1150_U103, P1_U4007);
  nand ginst7506 (P1_U4420, P1_R1117_U103, P1_U4000);
  nand ginst7507 (P1_U4421, P1_R1138_U114, P1_U3994);
  nand ginst7508 (P1_U4422, P1_R1192_U103, P1_U4005);
  nand ginst7509 (P1_U4423, P1_R1207_U103, P1_U4004);
  nand ginst7510 (P1_U4424, P1_R1171_U114, P1_U4011);
  nand ginst7511 (P1_U4425, P1_R1240_U114, P1_U3992);
  not ginst7512 (P1_U4426, P1_U3389);
  nand ginst7513 (P1_U4427, P1_U3025, P1_U3080);
  nand ginst7514 (P1_U4428, P1_R1222_U114, P1_U3024);
  nand ginst7515 (P1_U4429, P1_R1282_U8, P1_U4036);
  nand ginst7516 (P1_U4430, P1_U3494, P1_U4185);
  nand ginst7517 (P1_U4431, P1_U3655, P1_U4426);
  nand ginst7518 (P1_U4432, P1_REG2_REG_14__SCAN_IN, P1_U3018);
  nand ginst7519 (P1_U4433, P1_REG1_REG_14__SCAN_IN, P1_U3019);
  nand ginst7520 (P1_U4434, P1_REG0_REG_14__SCAN_IN, P1_U3020);
  nand ginst7521 (P1_U4435, P1_ADD_99_U74, P1_U3017);
  not ginst7522 (P1_U4436, P1_U3079);
  nand ginst7523 (P1_U4437, P1_U3034, P1_U3072);
  nand ginst7524 (P1_U4438, P1_R1150_U102, P1_U4007);
  nand ginst7525 (P1_U4439, P1_R1117_U102, P1_U4000);
  nand ginst7526 (P1_U4440, P1_R1138_U12, P1_U3994);
  nand ginst7527 (P1_U4441, P1_R1192_U102, P1_U4005);
  nand ginst7528 (P1_U4442, P1_R1207_U102, P1_U4004);
  nand ginst7529 (P1_U4443, P1_R1171_U12, P1_U4011);
  nand ginst7530 (P1_U4444, P1_R1240_U12, P1_U3992);
  not ginst7531 (P1_U4445, P1_U3390);
  nand ginst7532 (P1_U4446, P1_U3025, P1_U3079);
  nand ginst7533 (P1_U4447, P1_R1222_U12, P1_U3024);
  nand ginst7534 (P1_U4448, P1_R1282_U86, P1_U4036);
  nand ginst7535 (P1_U4449, P1_U3497, P1_U4185);
  nand ginst7536 (P1_U4450, P1_U3659, P1_U4445);
  nand ginst7537 (P1_U4451, P1_REG2_REG_15__SCAN_IN, P1_U3018);
  nand ginst7538 (P1_U4452, P1_REG1_REG_15__SCAN_IN, P1_U3019);
  nand ginst7539 (P1_U4453, P1_REG0_REG_15__SCAN_IN, P1_U3020);
  nand ginst7540 (P1_U4454, P1_ADD_99_U73, P1_U3017);
  not ginst7541 (P1_U4455, P1_U3074);
  nand ginst7542 (P1_U4456, P1_U3034, P1_U3080);
  nand ginst7543 (P1_U4457, P1_R1150_U113, P1_U4007);
  nand ginst7544 (P1_U4458, P1_R1117_U113, P1_U4000);
  nand ginst7545 (P1_U4459, P1_R1138_U113, P1_U3994);
  nand ginst7546 (P1_U4460, P1_R1192_U113, P1_U4005);
  nand ginst7547 (P1_U4461, P1_R1207_U113, P1_U4004);
  nand ginst7548 (P1_U4462, P1_R1171_U113, P1_U4011);
  nand ginst7549 (P1_U4463, P1_R1240_U113, P1_U3992);
  not ginst7550 (P1_U4464, P1_U3391);
  nand ginst7551 (P1_U4465, P1_U3025, P1_U3074);
  nand ginst7552 (P1_U4466, P1_R1222_U113, P1_U3024);
  nand ginst7553 (P1_U4467, P1_R1282_U9, P1_U4036);
  nand ginst7554 (P1_U4468, P1_U3500, P1_U4185);
  nand ginst7555 (P1_U4469, P1_U3663, P1_U4464);
  nand ginst7556 (P1_U4470, P1_REG2_REG_16__SCAN_IN, P1_U3018);
  nand ginst7557 (P1_U4471, P1_REG1_REG_16__SCAN_IN, P1_U3019);
  nand ginst7558 (P1_U4472, P1_REG0_REG_16__SCAN_IN, P1_U3020);
  nand ginst7559 (P1_U4473, P1_ADD_99_U72, P1_U3017);
  not ginst7560 (P1_U4474, P1_U3073);
  nand ginst7561 (P1_U4475, P1_U3034, P1_U3079);
  nand ginst7562 (P1_U4476, P1_R1150_U112, P1_U4007);
  nand ginst7563 (P1_U4477, P1_R1117_U112, P1_U4000);
  nand ginst7564 (P1_U4478, P1_R1138_U112, P1_U3994);
  nand ginst7565 (P1_U4479, P1_R1192_U112, P1_U4005);
  nand ginst7566 (P1_U4480, P1_R1207_U112, P1_U4004);
  nand ginst7567 (P1_U4481, P1_R1171_U112, P1_U4011);
  nand ginst7568 (P1_U4482, P1_R1240_U112, P1_U3992);
  not ginst7569 (P1_U4483, P1_U3392);
  nand ginst7570 (P1_U4484, P1_U3025, P1_U3073);
  nand ginst7571 (P1_U4485, P1_R1222_U112, P1_U3024);
  nand ginst7572 (P1_U4486, P1_R1282_U10, P1_U4036);
  nand ginst7573 (P1_U4487, P1_U3503, P1_U4185);
  nand ginst7574 (P1_U4488, P1_U3667, P1_U4483);
  nand ginst7575 (P1_U4489, P1_REG2_REG_17__SCAN_IN, P1_U3018);
  nand ginst7576 (P1_U4490, P1_REG1_REG_17__SCAN_IN, P1_U3019);
  nand ginst7577 (P1_U4491, P1_REG0_REG_17__SCAN_IN, P1_U3020);
  nand ginst7578 (P1_U4492, P1_ADD_99_U71, P1_U3017);
  not ginst7579 (P1_U4493, P1_U3069);
  nand ginst7580 (P1_U4494, P1_U3034, P1_U3074);
  nand ginst7581 (P1_U4495, P1_R1150_U14, P1_U4007);
  nand ginst7582 (P1_U4496, P1_R1117_U14, P1_U4000);
  nand ginst7583 (P1_U4497, P1_R1138_U111, P1_U3994);
  nand ginst7584 (P1_U4498, P1_R1192_U14, P1_U4005);
  nand ginst7585 (P1_U4499, P1_R1207_U14, P1_U4004);
  nand ginst7586 (P1_U4500, P1_R1171_U111, P1_U4011);
  nand ginst7587 (P1_U4501, P1_R1240_U111, P1_U3992);
  not ginst7588 (P1_U4502, P1_U3393);
  nand ginst7589 (P1_U4503, P1_U3025, P1_U3069);
  nand ginst7590 (P1_U4504, P1_R1222_U111, P1_U3024);
  nand ginst7591 (P1_U4505, P1_R1282_U11, P1_U4036);
  nand ginst7592 (P1_U4506, P1_U3506, P1_U4185);
  nand ginst7593 (P1_U4507, P1_U3671, P1_U4502);
  nand ginst7594 (P1_U4508, P1_REG2_REG_18__SCAN_IN, P1_U3018);
  nand ginst7595 (P1_U4509, P1_REG1_REG_18__SCAN_IN, P1_U3019);
  nand ginst7596 (P1_U4510, P1_REG0_REG_18__SCAN_IN, P1_U3020);
  nand ginst7597 (P1_U4511, P1_ADD_99_U70, P1_U3017);
  not ginst7598 (P1_U4512, P1_U3082);
  nand ginst7599 (P1_U4513, P1_U3034, P1_U3073);
  nand ginst7600 (P1_U4514, P1_R1150_U101, P1_U4007);
  nand ginst7601 (P1_U4515, P1_R1117_U101, P1_U4000);
  nand ginst7602 (P1_U4516, P1_R1138_U13, P1_U3994);
  nand ginst7603 (P1_U4517, P1_R1192_U101, P1_U4005);
  nand ginst7604 (P1_U4518, P1_R1207_U101, P1_U4004);
  nand ginst7605 (P1_U4519, P1_R1171_U13, P1_U4011);
  nand ginst7606 (P1_U4520, P1_R1240_U13, P1_U3992);
  not ginst7607 (P1_U4521, P1_U3394);
  nand ginst7608 (P1_U4522, P1_U3025, P1_U3082);
  nand ginst7609 (P1_U4523, P1_R1222_U13, P1_U3024);
  nand ginst7610 (P1_U4524, P1_R1282_U84, P1_U4036);
  nand ginst7611 (P1_U4525, P1_U3509, P1_U4185);
  nand ginst7612 (P1_U4526, P1_U3675, P1_U4521);
  nand ginst7613 (P1_U4527, P1_REG2_REG_19__SCAN_IN, P1_U3018);
  nand ginst7614 (P1_U4528, P1_REG1_REG_19__SCAN_IN, P1_U3019);
  nand ginst7615 (P1_U4529, P1_REG0_REG_19__SCAN_IN, P1_U3020);
  nand ginst7616 (P1_U4530, P1_ADD_99_U69, P1_U3017);
  not ginst7617 (P1_U4531, P1_U3081);
  nand ginst7618 (P1_U4532, P1_U3034, P1_U3069);
  nand ginst7619 (P1_U4533, P1_R1150_U100, P1_U4007);
  nand ginst7620 (P1_U4534, P1_R1117_U100, P1_U4000);
  nand ginst7621 (P1_U4535, P1_R1138_U110, P1_U3994);
  nand ginst7622 (P1_U4536, P1_R1192_U100, P1_U4005);
  nand ginst7623 (P1_U4537, P1_R1207_U100, P1_U4004);
  nand ginst7624 (P1_U4538, P1_R1171_U110, P1_U4011);
  nand ginst7625 (P1_U4539, P1_R1240_U110, P1_U3992);
  not ginst7626 (P1_U4540, P1_U3395);
  nand ginst7627 (P1_U4541, P1_U3025, P1_U3081);
  nand ginst7628 (P1_U4542, P1_R1222_U110, P1_U3024);
  nand ginst7629 (P1_U4543, P1_R1282_U12, P1_U4036);
  nand ginst7630 (P1_U4544, P1_U3512, P1_U4185);
  nand ginst7631 (P1_U4545, P1_U3679, P1_U4540);
  nand ginst7632 (P1_U4546, P1_REG2_REG_20__SCAN_IN, P1_U3018);
  nand ginst7633 (P1_U4547, P1_REG1_REG_20__SCAN_IN, P1_U3019);
  nand ginst7634 (P1_U4548, P1_REG0_REG_20__SCAN_IN, P1_U3020);
  nand ginst7635 (P1_U4549, P1_ADD_99_U68, P1_U3017);
  not ginst7636 (P1_U4550, P1_U3076);
  nand ginst7637 (P1_U4551, P1_U3034, P1_U3082);
  nand ginst7638 (P1_U4552, P1_R1150_U99, P1_U4007);
  nand ginst7639 (P1_U4553, P1_R1117_U99, P1_U4000);
  nand ginst7640 (P1_U4554, P1_R1138_U109, P1_U3994);
  nand ginst7641 (P1_U4555, P1_R1192_U99, P1_U4005);
  nand ginst7642 (P1_U4556, P1_R1207_U99, P1_U4004);
  nand ginst7643 (P1_U4557, P1_R1171_U109, P1_U4011);
  nand ginst7644 (P1_U4558, P1_R1240_U109, P1_U3992);
  not ginst7645 (P1_U4559, P1_U3396);
  nand ginst7646 (P1_U4560, P1_U3025, P1_U3076);
  nand ginst7647 (P1_U4561, P1_R1222_U109, P1_U3024);
  nand ginst7648 (P1_U4562, P1_R1282_U82, P1_U4036);
  nand ginst7649 (P1_U4563, P1_U3514, P1_U4185);
  nand ginst7650 (P1_U4564, P1_U3683, P1_U4559);
  nand ginst7651 (P1_U4565, P1_REG2_REG_21__SCAN_IN, P1_U3018);
  nand ginst7652 (P1_U4566, P1_REG1_REG_21__SCAN_IN, P1_U3019);
  nand ginst7653 (P1_U4567, P1_REG0_REG_21__SCAN_IN, P1_U3020);
  nand ginst7654 (P1_U4568, P1_ADD_99_U67, P1_U3017);
  not ginst7655 (P1_U4569, P1_U3075);
  nand ginst7656 (P1_U4570, P1_U3034, P1_U3081);
  nand ginst7657 (P1_U4571, P1_R1150_U97, P1_U4007);
  nand ginst7658 (P1_U4572, P1_R1117_U97, P1_U4000);
  nand ginst7659 (P1_U4573, P1_R1138_U14, P1_U3994);
  nand ginst7660 (P1_U4574, P1_R1192_U97, P1_U4005);
  nand ginst7661 (P1_U4575, P1_R1207_U97, P1_U4004);
  nand ginst7662 (P1_U4576, P1_R1171_U14, P1_U4011);
  nand ginst7663 (P1_U4577, P1_R1240_U14, P1_U3992);
  not ginst7664 (P1_U4578, P1_U3398);
  nand ginst7665 (P1_U4579, P1_U3025, P1_U3075);
  nand ginst7666 (P1_U4580, P1_R1222_U14, P1_U3024);
  nand ginst7667 (P1_U4581, P1_R1282_U13, P1_U4036);
  nand ginst7668 (P1_U4582, P1_U4025, P1_U4185);
  nand ginst7669 (P1_U4583, P1_U3687, P1_U4578);
  nand ginst7670 (P1_U4584, P1_REG2_REG_22__SCAN_IN, P1_U3018);
  nand ginst7671 (P1_U4585, P1_REG1_REG_22__SCAN_IN, P1_U3019);
  nand ginst7672 (P1_U4586, P1_REG0_REG_22__SCAN_IN, P1_U3020);
  nand ginst7673 (P1_U4587, P1_ADD_99_U66, P1_U3017);
  not ginst7674 (P1_U4588, P1_U3061);
  nand ginst7675 (P1_U4589, P1_U3034, P1_U3076);
  nand ginst7676 (P1_U4590, P1_R1150_U111, P1_U4007);
  nand ginst7677 (P1_U4591, P1_R1117_U111, P1_U4000);
  nand ginst7678 (P1_U4592, P1_R1138_U15, P1_U3994);
  nand ginst7679 (P1_U4593, P1_R1192_U111, P1_U4005);
  nand ginst7680 (P1_U4594, P1_R1207_U111, P1_U4004);
  nand ginst7681 (P1_U4595, P1_R1171_U15, P1_U4011);
  nand ginst7682 (P1_U4596, P1_R1240_U15, P1_U3992);
  not ginst7683 (P1_U4597, P1_U3400);
  nand ginst7684 (P1_U4598, P1_U3025, P1_U3061);
  nand ginst7685 (P1_U4599, P1_R1222_U15, P1_U3024);
  nand ginst7686 (P1_U4600, P1_R1282_U78, P1_U4036);
  nand ginst7687 (P1_U4601, P1_U4024, P1_U4185);
  nand ginst7688 (P1_U4602, P1_U3691, P1_U4597);
  nand ginst7689 (P1_U4603, P1_REG2_REG_23__SCAN_IN, P1_U3018);
  nand ginst7690 (P1_U4604, P1_REG1_REG_23__SCAN_IN, P1_U3019);
  nand ginst7691 (P1_U4605, P1_REG0_REG_23__SCAN_IN, P1_U3020);
  nand ginst7692 (P1_U4606, P1_ADD_99_U65, P1_U3017);
  not ginst7693 (P1_U4607, P1_U3066);
  nand ginst7694 (P1_U4608, P1_U3034, P1_U3075);
  nand ginst7695 (P1_U4609, P1_R1150_U110, P1_U4007);
  nand ginst7696 (P1_U4610, P1_R1117_U110, P1_U4000);
  nand ginst7697 (P1_U4611, P1_R1138_U108, P1_U3994);
  nand ginst7698 (P1_U4612, P1_R1192_U110, P1_U4005);
  nand ginst7699 (P1_U4613, P1_R1207_U110, P1_U4004);
  nand ginst7700 (P1_U4614, P1_R1171_U108, P1_U4011);
  nand ginst7701 (P1_U4615, P1_R1240_U108, P1_U3992);
  not ginst7702 (P1_U4616, P1_U3402);
  nand ginst7703 (P1_U4617, P1_U3025, P1_U3066);
  nand ginst7704 (P1_U4618, P1_R1222_U108, P1_U3024);
  nand ginst7705 (P1_U4619, P1_R1282_U14, P1_U4036);
  nand ginst7706 (P1_U4620, P1_U4023, P1_U4185);
  nand ginst7707 (P1_U4621, P1_U3695, P1_U4616);
  nand ginst7708 (P1_U4622, P1_REG2_REG_24__SCAN_IN, P1_U3018);
  nand ginst7709 (P1_U4623, P1_REG1_REG_24__SCAN_IN, P1_U3019);
  nand ginst7710 (P1_U4624, P1_REG0_REG_24__SCAN_IN, P1_U3020);
  nand ginst7711 (P1_U4625, P1_ADD_99_U64, P1_U3017);
  not ginst7712 (P1_U4626, P1_U3065);
  nand ginst7713 (P1_U4627, P1_U3034, P1_U3061);
  nand ginst7714 (P1_U4628, P1_R1150_U15, P1_U4007);
  nand ginst7715 (P1_U4629, P1_R1117_U15, P1_U4000);
  nand ginst7716 (P1_U4630, P1_R1138_U107, P1_U3994);
  nand ginst7717 (P1_U4631, P1_R1192_U15, P1_U4005);
  nand ginst7718 (P1_U4632, P1_R1207_U15, P1_U4004);
  nand ginst7719 (P1_U4633, P1_R1171_U107, P1_U4011);
  nand ginst7720 (P1_U4634, P1_R1240_U107, P1_U3992);
  not ginst7721 (P1_U4635, P1_U3404);
  nand ginst7722 (P1_U4636, P1_U3025, P1_U3065);
  nand ginst7723 (P1_U4637, P1_R1222_U107, P1_U3024);
  nand ginst7724 (P1_U4638, P1_R1282_U76, P1_U4036);
  nand ginst7725 (P1_U4639, P1_U4022, P1_U4185);
  nand ginst7726 (P1_U4640, P1_U3699, P1_U4635);
  nand ginst7727 (P1_U4641, P1_REG2_REG_25__SCAN_IN, P1_U3018);
  nand ginst7728 (P1_U4642, P1_REG1_REG_25__SCAN_IN, P1_U3019);
  nand ginst7729 (P1_U4643, P1_REG0_REG_25__SCAN_IN, P1_U3020);
  nand ginst7730 (P1_U4644, P1_ADD_99_U63, P1_U3017);
  not ginst7731 (P1_U4645, P1_U3058);
  nand ginst7732 (P1_U4646, P1_U3034, P1_U3066);
  nand ginst7733 (P1_U4647, P1_R1150_U96, P1_U4007);
  nand ginst7734 (P1_U4648, P1_R1117_U96, P1_U4000);
  nand ginst7735 (P1_U4649, P1_R1138_U106, P1_U3994);
  nand ginst7736 (P1_U4650, P1_R1192_U96, P1_U4005);
  nand ginst7737 (P1_U4651, P1_R1207_U96, P1_U4004);
  nand ginst7738 (P1_U4652, P1_R1171_U106, P1_U4011);
  nand ginst7739 (P1_U4653, P1_R1240_U106, P1_U3992);
  not ginst7740 (P1_U4654, P1_U3406);
  nand ginst7741 (P1_U4655, P1_U3025, P1_U3058);
  nand ginst7742 (P1_U4656, P1_R1222_U106, P1_U3024);
  nand ginst7743 (P1_U4657, P1_R1282_U15, P1_U4036);
  nand ginst7744 (P1_U4658, P1_U4021, P1_U4185);
  nand ginst7745 (P1_U4659, P1_U3703, P1_U4654);
  nand ginst7746 (P1_U4660, P1_REG2_REG_26__SCAN_IN, P1_U3018);
  nand ginst7747 (P1_U4661, P1_REG1_REG_26__SCAN_IN, P1_U3019);
  nand ginst7748 (P1_U4662, P1_REG0_REG_26__SCAN_IN, P1_U3020);
  nand ginst7749 (P1_U4663, P1_ADD_99_U62, P1_U3017);
  not ginst7750 (P1_U4664, P1_U3057);
  nand ginst7751 (P1_U4665, P1_U3034, P1_U3065);
  nand ginst7752 (P1_U4666, P1_R1150_U95, P1_U4007);
  nand ginst7753 (P1_U4667, P1_R1117_U95, P1_U4000);
  nand ginst7754 (P1_U4668, P1_R1138_U105, P1_U3994);
  nand ginst7755 (P1_U4669, P1_R1192_U95, P1_U4005);
  nand ginst7756 (P1_U4670, P1_R1207_U95, P1_U4004);
  nand ginst7757 (P1_U4671, P1_R1171_U105, P1_U4011);
  nand ginst7758 (P1_U4672, P1_R1240_U105, P1_U3992);
  not ginst7759 (P1_U4673, P1_U3408);
  nand ginst7760 (P1_U4674, P1_U3025, P1_U3057);
  nand ginst7761 (P1_U4675, P1_R1222_U105, P1_U3024);
  nand ginst7762 (P1_U4676, P1_R1282_U74, P1_U4036);
  nand ginst7763 (P1_U4677, P1_U4020, P1_U4185);
  nand ginst7764 (P1_U4678, P1_U3707, P1_U4673);
  nand ginst7765 (P1_U4679, P1_REG2_REG_27__SCAN_IN, P1_U3018);
  nand ginst7766 (P1_U4680, P1_REG1_REG_27__SCAN_IN, P1_U3019);
  nand ginst7767 (P1_U4681, P1_REG0_REG_27__SCAN_IN, P1_U3020);
  nand ginst7768 (P1_U4682, P1_ADD_99_U61, P1_U3017);
  not ginst7769 (P1_U4683, P1_U3053);
  nand ginst7770 (P1_U4684, P1_U3034, P1_U3058);
  nand ginst7771 (P1_U4685, P1_R1150_U109, P1_U4007);
  nand ginst7772 (P1_U4686, P1_R1117_U109, P1_U4000);
  nand ginst7773 (P1_U4687, P1_R1138_U16, P1_U3994);
  nand ginst7774 (P1_U4688, P1_R1192_U109, P1_U4005);
  nand ginst7775 (P1_U4689, P1_R1207_U109, P1_U4004);
  nand ginst7776 (P1_U4690, P1_R1171_U16, P1_U4011);
  nand ginst7777 (P1_U4691, P1_R1240_U16, P1_U3992);
  not ginst7778 (P1_U4692, P1_U3410);
  nand ginst7779 (P1_U4693, P1_U3025, P1_U3053);
  nand ginst7780 (P1_U4694, P1_R1222_U16, P1_U3024);
  nand ginst7781 (P1_U4695, P1_R1282_U16, P1_U4036);
  nand ginst7782 (P1_U4696, P1_U4019, P1_U4185);
  nand ginst7783 (P1_U4697, P1_U3711, P1_U4692);
  nand ginst7784 (P1_U4698, P1_REG2_REG_28__SCAN_IN, P1_U3018);
  nand ginst7785 (P1_U4699, P1_REG1_REG_28__SCAN_IN, P1_U3019);
  nand ginst7786 (P1_U4700, P1_REG0_REG_28__SCAN_IN, P1_U3020);
  nand ginst7787 (P1_U4701, P1_ADD_99_U60, P1_U3017);
  not ginst7788 (P1_U4702, P1_U3054);
  nand ginst7789 (P1_U4703, P1_U3034, P1_U3057);
  nand ginst7790 (P1_U4704, P1_R1150_U16, P1_U4007);
  nand ginst7791 (P1_U4705, P1_R1117_U16, P1_U4000);
  nand ginst7792 (P1_U4706, P1_R1138_U104, P1_U3994);
  nand ginst7793 (P1_U4707, P1_R1192_U16, P1_U4005);
  nand ginst7794 (P1_U4708, P1_R1207_U16, P1_U4004);
  nand ginst7795 (P1_U4709, P1_R1171_U104, P1_U4011);
  nand ginst7796 (P1_U4710, P1_R1240_U104, P1_U3992);
  not ginst7797 (P1_U4711, P1_U3412);
  nand ginst7798 (P1_U4712, P1_U3025, P1_U3054);
  nand ginst7799 (P1_U4713, P1_R1222_U104, P1_U3024);
  nand ginst7800 (P1_U4714, P1_R1282_U72, P1_U4036);
  nand ginst7801 (P1_U4715, P1_U4018, P1_U4185);
  nand ginst7802 (P1_U4716, P1_U3715, P1_U4711);
  nand ginst7803 (P1_U4717, P1_ADD_99_U5, P1_U3017);
  nand ginst7804 (P1_U4718, P1_REG2_REG_29__SCAN_IN, P1_U3018);
  nand ginst7805 (P1_U4719, P1_REG1_REG_29__SCAN_IN, P1_U3019);
  nand ginst7806 (P1_U4720, P1_REG0_REG_29__SCAN_IN, P1_U3020);
  not ginst7807 (P1_U4721, P1_U3055);
  nand ginst7808 (P1_U4722, P1_U3034, P1_U3053);
  nand ginst7809 (P1_U4723, P1_R1150_U94, P1_U4007);
  nand ginst7810 (P1_U4724, P1_R1117_U94, P1_U4000);
  nand ginst7811 (P1_U4725, P1_R1138_U103, P1_U3994);
  nand ginst7812 (P1_U4726, P1_R1192_U94, P1_U4005);
  nand ginst7813 (P1_U4727, P1_R1207_U94, P1_U4004);
  nand ginst7814 (P1_U4728, P1_R1171_U103, P1_U4011);
  nand ginst7815 (P1_U4729, P1_R1240_U103, P1_U3992);
  not ginst7816 (P1_U4730, P1_U3414);
  nand ginst7817 (P1_U4731, P1_U3025, P1_U3055);
  nand ginst7818 (P1_U4732, P1_R1222_U103, P1_U3024);
  nand ginst7819 (P1_U4733, P1_R1282_U17, P1_U4036);
  nand ginst7820 (P1_U4734, P1_U4017, P1_U4185);
  nand ginst7821 (P1_U4735, P1_U3719, P1_U4730);
  nand ginst7822 (P1_U4736, P1_REG2_REG_30__SCAN_IN, P1_U3018);
  nand ginst7823 (P1_U4737, P1_REG1_REG_30__SCAN_IN, P1_U3019);
  nand ginst7824 (P1_U4738, P1_REG0_REG_30__SCAN_IN, P1_U3020);
  not ginst7825 (P1_U4739, P1_U3059);
  nand ginst7826 (P1_U4740, P1_U3359, P1_U5811);
  nand ginst7827 (P1_U4741, P1_U3954, P1_U4740);
  nand ginst7828 (P1_U4742, P1_U3059, P1_U3720);
  nand ginst7829 (P1_U4743, P1_U3034, P1_U3054);
  nand ginst7830 (P1_U4744, P1_R1150_U17, P1_U4007);
  nand ginst7831 (P1_U4745, P1_R1117_U17, P1_U4000);
  nand ginst7832 (P1_U4746, P1_R1138_U102, P1_U3994);
  nand ginst7833 (P1_U4747, P1_R1192_U17, P1_U4005);
  nand ginst7834 (P1_U4748, P1_R1207_U17, P1_U4004);
  nand ginst7835 (P1_U4749, P1_R1171_U102, P1_U4011);
  nand ginst7836 (P1_U4750, P1_R1240_U102, P1_U3992);
  not ginst7837 (P1_U4751, P1_U3416);
  nand ginst7838 (P1_U4752, P1_R1222_U102, P1_U3024);
  nand ginst7839 (P1_U4753, P1_R1282_U70, P1_U4036);
  nand ginst7840 (P1_U4754, P1_U4028, P1_U4185);
  nand ginst7841 (P1_U4755, P1_U3724, P1_U4751);
  nand ginst7842 (P1_U4756, P1_REG2_REG_31__SCAN_IN, P1_U3018);
  nand ginst7843 (P1_U4757, P1_REG1_REG_31__SCAN_IN, P1_U3019);
  nand ginst7844 (P1_U4758, P1_REG0_REG_31__SCAN_IN, P1_U3020);
  not ginst7845 (P1_U4759, P1_U3056);
  nand ginst7846 (P1_U4760, P1_R1282_U19, P1_U4036);
  nand ginst7847 (P1_U4761, P1_U4027, P1_U4185);
  nand ginst7848 (P1_U4762, P1_U3987, P1_U4760, P1_U4761);
  nand ginst7849 (P1_U4763, P1_R1282_U68, P1_U4036);
  nand ginst7850 (P1_U4764, P1_U4026, P1_U4185);
  nand ginst7851 (P1_U4765, P1_U3987, P1_U4763, P1_U4764);
  nand ginst7852 (P1_U4766, P1_U3016, P1_U3727);
  nand ginst7853 (P1_U4767, P1_U3421, P1_U4766);
  nand ginst7854 (P1_U4768, P1_U3995, P1_U5802);
  not ginst7855 (P1_U4769, P1_U3426);
  nand ginst7856 (P1_U4770, P1_U3036, P1_U3078);
  nand ginst7857 (P1_U4771, P1_REG3_REG_0__SCAN_IN, P1_U3033);
  nand ginst7858 (P1_U4772, P1_R1222_U96, P1_U3032);
  nand ginst7859 (P1_U4773, P1_U3031, P1_U3456);
  nand ginst7860 (P1_U4774, P1_U3030, P1_U3456);
  nand ginst7861 (P1_U4775, P1_U3036, P1_U3068);
  nand ginst7862 (P1_U4776, P1_REG3_REG_1__SCAN_IN, P1_U3033);
  nand ginst7863 (P1_U4777, P1_R1222_U95, P1_U3032);
  nand ginst7864 (P1_U4778, P1_U3031, P1_U3461);
  nand ginst7865 (P1_U4779, P1_R1282_U56, P1_U3030);
  nand ginst7866 (P1_U4780, P1_U3036, P1_U3064);
  nand ginst7867 (P1_U4781, P1_REG3_REG_2__SCAN_IN, P1_U3033);
  nand ginst7868 (P1_U4782, P1_R1222_U17, P1_U3032);
  nand ginst7869 (P1_U4783, P1_U3031, P1_U3464);
  nand ginst7870 (P1_U4784, P1_R1282_U18, P1_U3030);
  nand ginst7871 (P1_U4785, P1_U3036, P1_U3060);
  nand ginst7872 (P1_U4786, P1_ADD_99_U4, P1_U3033);
  nand ginst7873 (P1_U4787, P1_R1222_U101, P1_U3032);
  nand ginst7874 (P1_U4788, P1_U3031, P1_U3467);
  nand ginst7875 (P1_U4789, P1_R1282_U20, P1_U3030);
  nand ginst7876 (P1_U4790, P1_U3036, P1_U3067);
  nand ginst7877 (P1_U4791, P1_ADD_99_U59, P1_U3033);
  nand ginst7878 (P1_U4792, P1_R1222_U100, P1_U3032);
  nand ginst7879 (P1_U4793, P1_U3031, P1_U3470);
  nand ginst7880 (P1_U4794, P1_R1282_U21, P1_U3030);
  nand ginst7881 (P1_U4795, P1_U3036, P1_U3071);
  nand ginst7882 (P1_U4796, P1_ADD_99_U58, P1_U3033);
  nand ginst7883 (P1_U4797, P1_R1222_U18, P1_U3032);
  nand ginst7884 (P1_U4798, P1_U3031, P1_U3473);
  nand ginst7885 (P1_U4799, P1_R1282_U65, P1_U3030);
  nand ginst7886 (P1_U4800, P1_U3036, P1_U3070);
  nand ginst7887 (P1_U4801, P1_ADD_99_U57, P1_U3033);
  nand ginst7888 (P1_U4802, P1_R1222_U99, P1_U3032);
  nand ginst7889 (P1_U4803, P1_U3031, P1_U3476);
  nand ginst7890 (P1_U4804, P1_R1282_U22, P1_U3030);
  nand ginst7891 (P1_U4805, P1_U3036, P1_U3084);
  nand ginst7892 (P1_U4806, P1_ADD_99_U56, P1_U3033);
  nand ginst7893 (P1_U4807, P1_R1222_U19, P1_U3032);
  nand ginst7894 (P1_U4808, P1_U3031, P1_U3479);
  nand ginst7895 (P1_U4809, P1_R1282_U23, P1_U3030);
  nand ginst7896 (P1_U4810, P1_U3036, P1_U3083);
  nand ginst7897 (P1_U4811, P1_ADD_99_U55, P1_U3033);
  nand ginst7898 (P1_U4812, P1_R1222_U98, P1_U3032);
  nand ginst7899 (P1_U4813, P1_U3031, P1_U3482);
  nand ginst7900 (P1_U4814, P1_R1282_U24, P1_U3030);
  nand ginst7901 (P1_U4815, P1_U3036, P1_U3062);
  nand ginst7902 (P1_U4816, P1_ADD_99_U54, P1_U3033);
  nand ginst7903 (P1_U4817, P1_R1222_U97, P1_U3032);
  nand ginst7904 (P1_U4818, P1_U3031, P1_U3485);
  nand ginst7905 (P1_U4819, P1_R1282_U63, P1_U3030);
  nand ginst7906 (P1_U4820, P1_U3036, P1_U3063);
  nand ginst7907 (P1_U4821, P1_ADD_99_U78, P1_U3033);
  nand ginst7908 (P1_U4822, P1_R1222_U11, P1_U3032);
  nand ginst7909 (P1_U4823, P1_U3031, P1_U3488);
  nand ginst7910 (P1_U4824, P1_R1282_U6, P1_U3030);
  nand ginst7911 (P1_U4825, P1_U3036, P1_U3072);
  nand ginst7912 (P1_U4826, P1_ADD_99_U77, P1_U3033);
  nand ginst7913 (P1_U4827, P1_R1222_U115, P1_U3032);
  nand ginst7914 (P1_U4828, P1_U3031, P1_U3491);
  nand ginst7915 (P1_U4829, P1_R1282_U7, P1_U3030);
  nand ginst7916 (P1_U4830, P1_U3036, P1_U3080);
  nand ginst7917 (P1_U4831, P1_ADD_99_U76, P1_U3033);
  nand ginst7918 (P1_U4832, P1_R1222_U114, P1_U3032);
  nand ginst7919 (P1_U4833, P1_U3031, P1_U3494);
  nand ginst7920 (P1_U4834, P1_R1282_U8, P1_U3030);
  nand ginst7921 (P1_U4835, P1_U3036, P1_U3079);
  nand ginst7922 (P1_U4836, P1_ADD_99_U75, P1_U3033);
  nand ginst7923 (P1_U4837, P1_R1222_U12, P1_U3032);
  nand ginst7924 (P1_U4838, P1_U3031, P1_U3497);
  nand ginst7925 (P1_U4839, P1_R1282_U86, P1_U3030);
  nand ginst7926 (P1_U4840, P1_U3036, P1_U3074);
  nand ginst7927 (P1_U4841, P1_ADD_99_U74, P1_U3033);
  nand ginst7928 (P1_U4842, P1_R1222_U113, P1_U3032);
  nand ginst7929 (P1_U4843, P1_U3031, P1_U3500);
  nand ginst7930 (P1_U4844, P1_R1282_U9, P1_U3030);
  nand ginst7931 (P1_U4845, P1_U3036, P1_U3073);
  nand ginst7932 (P1_U4846, P1_ADD_99_U73, P1_U3033);
  nand ginst7933 (P1_U4847, P1_R1222_U112, P1_U3032);
  nand ginst7934 (P1_U4848, P1_U3031, P1_U3503);
  nand ginst7935 (P1_U4849, P1_R1282_U10, P1_U3030);
  nand ginst7936 (P1_U4850, P1_U3036, P1_U3069);
  nand ginst7937 (P1_U4851, P1_ADD_99_U72, P1_U3033);
  nand ginst7938 (P1_U4852, P1_R1222_U111, P1_U3032);
  nand ginst7939 (P1_U4853, P1_U3031, P1_U3506);
  nand ginst7940 (P1_U4854, P1_R1282_U11, P1_U3030);
  nand ginst7941 (P1_U4855, P1_U3036, P1_U3082);
  nand ginst7942 (P1_U4856, P1_ADD_99_U71, P1_U3033);
  nand ginst7943 (P1_U4857, P1_R1222_U13, P1_U3032);
  nand ginst7944 (P1_U4858, P1_U3031, P1_U3509);
  nand ginst7945 (P1_U4859, P1_R1282_U84, P1_U3030);
  nand ginst7946 (P1_U4860, P1_U3036, P1_U3081);
  nand ginst7947 (P1_U4861, P1_ADD_99_U70, P1_U3033);
  nand ginst7948 (P1_U4862, P1_R1222_U110, P1_U3032);
  nand ginst7949 (P1_U4863, P1_U3031, P1_U3512);
  nand ginst7950 (P1_U4864, P1_R1282_U12, P1_U3030);
  nand ginst7951 (P1_U4865, P1_U3036, P1_U3076);
  nand ginst7952 (P1_U4866, P1_ADD_99_U69, P1_U3033);
  nand ginst7953 (P1_U4867, P1_R1222_U109, P1_U3032);
  nand ginst7954 (P1_U4868, P1_U3031, P1_U3514);
  nand ginst7955 (P1_U4869, P1_R1282_U82, P1_U3030);
  nand ginst7956 (P1_U4870, P1_U3036, P1_U3075);
  nand ginst7957 (P1_U4871, P1_ADD_99_U68, P1_U3033);
  nand ginst7958 (P1_U4872, P1_R1222_U14, P1_U3032);
  nand ginst7959 (P1_U4873, P1_U3031, P1_U4025);
  nand ginst7960 (P1_U4874, P1_R1282_U13, P1_U3030);
  nand ginst7961 (P1_U4875, P1_U3036, P1_U3061);
  nand ginst7962 (P1_U4876, P1_ADD_99_U67, P1_U3033);
  nand ginst7963 (P1_U4877, P1_R1222_U15, P1_U3032);
  nand ginst7964 (P1_U4878, P1_U3031, P1_U4024);
  nand ginst7965 (P1_U4879, P1_R1282_U78, P1_U3030);
  nand ginst7966 (P1_U4880, P1_U3036, P1_U3066);
  nand ginst7967 (P1_U4881, P1_ADD_99_U66, P1_U3033);
  nand ginst7968 (P1_U4882, P1_R1222_U108, P1_U3032);
  nand ginst7969 (P1_U4883, P1_U3031, P1_U4023);
  nand ginst7970 (P1_U4884, P1_R1282_U14, P1_U3030);
  nand ginst7971 (P1_U4885, P1_U3036, P1_U3065);
  nand ginst7972 (P1_U4886, P1_ADD_99_U65, P1_U3033);
  nand ginst7973 (P1_U4887, P1_R1222_U107, P1_U3032);
  nand ginst7974 (P1_U4888, P1_U3031, P1_U4022);
  nand ginst7975 (P1_U4889, P1_R1282_U76, P1_U3030);
  nand ginst7976 (P1_U4890, P1_U3036, P1_U3058);
  nand ginst7977 (P1_U4891, P1_ADD_99_U64, P1_U3033);
  nand ginst7978 (P1_U4892, P1_R1222_U106, P1_U3032);
  nand ginst7979 (P1_U4893, P1_U3031, P1_U4021);
  nand ginst7980 (P1_U4894, P1_R1282_U15, P1_U3030);
  nand ginst7981 (P1_U4895, P1_U3036, P1_U3057);
  nand ginst7982 (P1_U4896, P1_ADD_99_U63, P1_U3033);
  nand ginst7983 (P1_U4897, P1_R1222_U105, P1_U3032);
  nand ginst7984 (P1_U4898, P1_U3031, P1_U4020);
  nand ginst7985 (P1_U4899, P1_R1282_U74, P1_U3030);
  nand ginst7986 (P1_U4900, P1_U3036, P1_U3053);
  nand ginst7987 (P1_U4901, P1_ADD_99_U62, P1_U3033);
  nand ginst7988 (P1_U4902, P1_R1222_U16, P1_U3032);
  nand ginst7989 (P1_U4903, P1_U3031, P1_U4019);
  nand ginst7990 (P1_U4904, P1_R1282_U16, P1_U3030);
  nand ginst7991 (P1_U4905, P1_U3036, P1_U3054);
  nand ginst7992 (P1_U4906, P1_ADD_99_U61, P1_U3033);
  nand ginst7993 (P1_U4907, P1_R1222_U104, P1_U3032);
  nand ginst7994 (P1_U4908, P1_U3031, P1_U4018);
  nand ginst7995 (P1_U4909, P1_R1282_U72, P1_U3030);
  nand ginst7996 (P1_U4910, P1_U3036, P1_U3055);
  nand ginst7997 (P1_U4911, P1_ADD_99_U60, P1_U3033);
  nand ginst7998 (P1_U4912, P1_R1222_U103, P1_U3032);
  nand ginst7999 (P1_U4913, P1_U3031, P1_U4017);
  nand ginst8000 (P1_U4914, P1_R1282_U17, P1_U3030);
  nand ginst8001 (P1_U4915, P1_ADD_99_U5, P1_U3033);
  nand ginst8002 (P1_U4916, P1_R1222_U102, P1_U3032);
  nand ginst8003 (P1_U4917, P1_U3031, P1_U4028);
  nand ginst8004 (P1_U4918, P1_R1282_U70, P1_U3030);
  nand ginst8005 (P1_U4919, P1_U3031, P1_U4027);
  nand ginst8006 (P1_U4920, P1_R1282_U19, P1_U3030);
  nand ginst8007 (P1_U4921, P1_U3031, P1_U4026);
  nand ginst8008 (P1_U4922, P1_R1282_U68, P1_U3030);
  nand ginst8009 (P1_U4923, P1_U3421, P1_U3786, P1_U3787, P1_U3789, P1_U4769);
  nand ginst8010 (P1_U4924, P1_R1105_U13, P1_U3042);
  nand ginst8011 (P1_U4925, P1_U3040, P1_U3452);
  nand ginst8012 (P1_U4926, P1_R1162_U13, P1_U3038);
  nand ginst8013 (P1_U4927, P1_U4924, P1_U4925, P1_U4926);
  nand ginst8014 (P1_U4928, P1_U3372, P1_U3425);
  nand ginst8015 (P1_U4929, P1_U4928, P1_U5786);
  nand ginst8016 (P1_U4930, P1_U3954, P1_U4929);
  not ginst8017 (P1_U4931, P1_U3085);
  not ginst8018 (P1_U4932, P1_U3428);
  nand ginst8019 (P1_U4933, P1_U3044, P1_U4927);
  nand ginst8020 (P1_U4934, P1_R1105_U13, P1_U3043);
  nand ginst8021 (P1_U4935, P1_REG3_REG_19__SCAN_IN, P1_U3086);
  nand ginst8022 (P1_U4936, P1_U3041, P1_U3452);
  nand ginst8023 (P1_U4937, P1_R1162_U13, P1_U3039);
  nand ginst8024 (P1_U4938, P1_ADDR_REG_19__SCAN_IN, P1_U4932);
  nand ginst8025 (P1_U4939, P1_R1105_U75, P1_U3042);
  nand ginst8026 (P1_U4940, P1_U3040, P1_U3511);
  nand ginst8027 (P1_U4941, P1_R1162_U75, P1_U3038);
  nand ginst8028 (P1_U4942, P1_U4939, P1_U4940, P1_U4941);
  nand ginst8029 (P1_U4943, P1_U3044, P1_U4942);
  nand ginst8030 (P1_U4944, P1_R1105_U75, P1_U3043);
  nand ginst8031 (P1_U4945, P1_REG3_REG_18__SCAN_IN, P1_U3086);
  nand ginst8032 (P1_U4946, P1_U3041, P1_U3511);
  nand ginst8033 (P1_U4947, P1_R1162_U75, P1_U3039);
  nand ginst8034 (P1_U4948, P1_ADDR_REG_18__SCAN_IN, P1_U4932);
  nand ginst8035 (P1_U4949, P1_R1105_U12, P1_U3042);
  nand ginst8036 (P1_U4950, P1_U3040, P1_U3508);
  nand ginst8037 (P1_U4951, P1_R1162_U12, P1_U3038);
  nand ginst8038 (P1_U4952, P1_U4949, P1_U4950, P1_U4951);
  nand ginst8039 (P1_U4953, P1_U3044, P1_U4952);
  nand ginst8040 (P1_U4954, P1_R1105_U12, P1_U3043);
  nand ginst8041 (P1_U4955, P1_REG3_REG_17__SCAN_IN, P1_U3086);
  nand ginst8042 (P1_U4956, P1_U3041, P1_U3508);
  nand ginst8043 (P1_U4957, P1_R1162_U12, P1_U3039);
  nand ginst8044 (P1_U4958, P1_ADDR_REG_17__SCAN_IN, P1_U4932);
  nand ginst8045 (P1_U4959, P1_R1105_U76, P1_U3042);
  nand ginst8046 (P1_U4960, P1_U3040, P1_U3505);
  nand ginst8047 (P1_U4961, P1_R1162_U76, P1_U3038);
  nand ginst8048 (P1_U4962, P1_U4959, P1_U4960, P1_U4961);
  nand ginst8049 (P1_U4963, P1_U3044, P1_U4962);
  nand ginst8050 (P1_U4964, P1_R1105_U76, P1_U3043);
  nand ginst8051 (P1_U4965, P1_REG3_REG_16__SCAN_IN, P1_U3086);
  nand ginst8052 (P1_U4966, P1_U3041, P1_U3505);
  nand ginst8053 (P1_U4967, P1_R1162_U76, P1_U3039);
  nand ginst8054 (P1_U4968, P1_ADDR_REG_16__SCAN_IN, P1_U4932);
  nand ginst8055 (P1_U4969, P1_R1105_U77, P1_U3042);
  nand ginst8056 (P1_U4970, P1_U3040, P1_U3502);
  nand ginst8057 (P1_U4971, P1_R1162_U77, P1_U3038);
  nand ginst8058 (P1_U4972, P1_U4969, P1_U4970, P1_U4971);
  nand ginst8059 (P1_U4973, P1_U3044, P1_U4972);
  nand ginst8060 (P1_U4974, P1_R1105_U77, P1_U3043);
  nand ginst8061 (P1_U4975, P1_REG3_REG_15__SCAN_IN, P1_U3086);
  nand ginst8062 (P1_U4976, P1_U3041, P1_U3502);
  nand ginst8063 (P1_U4977, P1_R1162_U77, P1_U3039);
  nand ginst8064 (P1_U4978, P1_ADDR_REG_15__SCAN_IN, P1_U4932);
  nand ginst8065 (P1_U4979, P1_R1105_U78, P1_U3042);
  nand ginst8066 (P1_U4980, P1_U3040, P1_U3499);
  nand ginst8067 (P1_U4981, P1_R1162_U78, P1_U3038);
  nand ginst8068 (P1_U4982, P1_U4979, P1_U4980, P1_U4981);
  nand ginst8069 (P1_U4983, P1_U3044, P1_U4982);
  nand ginst8070 (P1_U4984, P1_R1105_U78, P1_U3043);
  nand ginst8071 (P1_U4985, P1_REG3_REG_14__SCAN_IN, P1_U3086);
  nand ginst8072 (P1_U4986, P1_U3041, P1_U3499);
  nand ginst8073 (P1_U4987, P1_R1162_U78, P1_U3039);
  nand ginst8074 (P1_U4988, P1_ADDR_REG_14__SCAN_IN, P1_U4932);
  nand ginst8075 (P1_U4989, P1_R1105_U11, P1_U3042);
  nand ginst8076 (P1_U4990, P1_U3040, P1_U3496);
  nand ginst8077 (P1_U4991, P1_R1162_U11, P1_U3038);
  nand ginst8078 (P1_U4992, P1_U4989, P1_U4990, P1_U4991);
  nand ginst8079 (P1_U4993, P1_U3044, P1_U4992);
  nand ginst8080 (P1_U4994, P1_R1105_U11, P1_U3043);
  nand ginst8081 (P1_U4995, P1_REG3_REG_13__SCAN_IN, P1_U3086);
  nand ginst8082 (P1_U4996, P1_U3041, P1_U3496);
  nand ginst8083 (P1_U4997, P1_R1162_U11, P1_U3039);
  nand ginst8084 (P1_U4998, P1_ADDR_REG_13__SCAN_IN, P1_U4932);
  nand ginst8085 (P1_U4999, P1_R1105_U79, P1_U3042);
  nand ginst8086 (P1_U5000, P1_U3040, P1_U3493);
  nand ginst8087 (P1_U5001, P1_R1162_U79, P1_U3038);
  nand ginst8088 (P1_U5002, P1_U4999, P1_U5000, P1_U5001);
  nand ginst8089 (P1_U5003, P1_U3044, P1_U5002);
  nand ginst8090 (P1_U5004, P1_R1105_U79, P1_U3043);
  nand ginst8091 (P1_U5005, P1_REG3_REG_12__SCAN_IN, P1_U3086);
  nand ginst8092 (P1_U5006, P1_U3041, P1_U3493);
  nand ginst8093 (P1_U5007, P1_R1162_U79, P1_U3039);
  nand ginst8094 (P1_U5008, P1_ADDR_REG_12__SCAN_IN, P1_U4932);
  nand ginst8095 (P1_U5009, P1_R1105_U80, P1_U3042);
  nand ginst8096 (P1_U5010, P1_U3040, P1_U3490);
  nand ginst8097 (P1_U5011, P1_R1162_U80, P1_U3038);
  nand ginst8098 (P1_U5012, P1_U5009, P1_U5010, P1_U5011);
  nand ginst8099 (P1_U5013, P1_U3044, P1_U5012);
  nand ginst8100 (P1_U5014, P1_R1105_U80, P1_U3043);
  nand ginst8101 (P1_U5015, P1_REG3_REG_11__SCAN_IN, P1_U3086);
  nand ginst8102 (P1_U5016, P1_U3041, P1_U3490);
  nand ginst8103 (P1_U5017, P1_R1162_U80, P1_U3039);
  nand ginst8104 (P1_U5018, P1_ADDR_REG_11__SCAN_IN, P1_U4932);
  nand ginst8105 (P1_U5019, P1_R1105_U10, P1_U3042);
  nand ginst8106 (P1_U5020, P1_U3040, P1_U3487);
  nand ginst8107 (P1_U5021, P1_R1162_U10, P1_U3038);
  nand ginst8108 (P1_U5022, P1_U5019, P1_U5020, P1_U5021);
  nand ginst8109 (P1_U5023, P1_U3044, P1_U5022);
  nand ginst8110 (P1_U5024, P1_R1105_U10, P1_U3043);
  nand ginst8111 (P1_U5025, P1_REG3_REG_10__SCAN_IN, P1_U3086);
  nand ginst8112 (P1_U5026, P1_U3041, P1_U3487);
  nand ginst8113 (P1_U5027, P1_R1162_U10, P1_U3039);
  nand ginst8114 (P1_U5028, P1_ADDR_REG_10__SCAN_IN, P1_U4932);
  nand ginst8115 (P1_U5029, P1_R1105_U70, P1_U3042);
  nand ginst8116 (P1_U5030, P1_U3040, P1_U3484);
  nand ginst8117 (P1_U5031, P1_R1162_U70, P1_U3038);
  nand ginst8118 (P1_U5032, P1_U5029, P1_U5030, P1_U5031);
  nand ginst8119 (P1_U5033, P1_U3044, P1_U5032);
  nand ginst8120 (P1_U5034, P1_R1105_U70, P1_U3043);
  nand ginst8121 (P1_U5035, P1_REG3_REG_9__SCAN_IN, P1_U3086);
  nand ginst8122 (P1_U5036, P1_U3041, P1_U3484);
  nand ginst8123 (P1_U5037, P1_R1162_U70, P1_U3039);
  nand ginst8124 (P1_U5038, P1_ADDR_REG_9__SCAN_IN, P1_U4932);
  nand ginst8125 (P1_U5039, P1_R1105_U71, P1_U3042);
  nand ginst8126 (P1_U5040, P1_U3040, P1_U3481);
  nand ginst8127 (P1_U5041, P1_R1162_U71, P1_U3038);
  nand ginst8128 (P1_U5042, P1_U5039, P1_U5040, P1_U5041);
  nand ginst8129 (P1_U5043, P1_U3044, P1_U5042);
  nand ginst8130 (P1_U5044, P1_R1105_U71, P1_U3043);
  nand ginst8131 (P1_U5045, P1_REG3_REG_8__SCAN_IN, P1_U3086);
  nand ginst8132 (P1_U5046, P1_U3041, P1_U3481);
  nand ginst8133 (P1_U5047, P1_R1162_U71, P1_U3039);
  nand ginst8134 (P1_U5048, P1_ADDR_REG_8__SCAN_IN, P1_U4932);
  nand ginst8135 (P1_U5049, P1_R1105_U16, P1_U3042);
  nand ginst8136 (P1_U5050, P1_U3040, P1_U3478);
  nand ginst8137 (P1_U5051, P1_R1162_U16, P1_U3038);
  nand ginst8138 (P1_U5052, P1_U5049, P1_U5050, P1_U5051);
  nand ginst8139 (P1_U5053, P1_U3044, P1_U5052);
  nand ginst8140 (P1_U5054, P1_R1105_U16, P1_U3043);
  nand ginst8141 (P1_U5055, P1_REG3_REG_7__SCAN_IN, P1_U3086);
  nand ginst8142 (P1_U5056, P1_U3041, P1_U3478);
  nand ginst8143 (P1_U5057, P1_R1162_U16, P1_U3039);
  nand ginst8144 (P1_U5058, P1_ADDR_REG_7__SCAN_IN, P1_U4932);
  nand ginst8145 (P1_U5059, P1_R1105_U72, P1_U3042);
  nand ginst8146 (P1_U5060, P1_U3040, P1_U3475);
  nand ginst8147 (P1_U5061, P1_R1162_U72, P1_U3038);
  nand ginst8148 (P1_U5062, P1_U5059, P1_U5060, P1_U5061);
  nand ginst8149 (P1_U5063, P1_U3044, P1_U5062);
  nand ginst8150 (P1_U5064, P1_R1105_U72, P1_U3043);
  nand ginst8151 (P1_U5065, P1_REG3_REG_6__SCAN_IN, P1_U3086);
  nand ginst8152 (P1_U5066, P1_U3041, P1_U3475);
  nand ginst8153 (P1_U5067, P1_R1162_U72, P1_U3039);
  nand ginst8154 (P1_U5068, P1_ADDR_REG_6__SCAN_IN, P1_U4932);
  nand ginst8155 (P1_U5069, P1_R1105_U15, P1_U3042);
  nand ginst8156 (P1_U5070, P1_U3040, P1_U3472);
  nand ginst8157 (P1_U5071, P1_R1162_U15, P1_U3038);
  nand ginst8158 (P1_U5072, P1_U5069, P1_U5070, P1_U5071);
  nand ginst8159 (P1_U5073, P1_U3044, P1_U5072);
  nand ginst8160 (P1_U5074, P1_R1105_U15, P1_U3043);
  nand ginst8161 (P1_U5075, P1_REG3_REG_5__SCAN_IN, P1_U3086);
  nand ginst8162 (P1_U5076, P1_U3041, P1_U3472);
  nand ginst8163 (P1_U5077, P1_R1162_U15, P1_U3039);
  nand ginst8164 (P1_U5078, P1_ADDR_REG_5__SCAN_IN, P1_U4932);
  nand ginst8165 (P1_U5079, P1_R1105_U73, P1_U3042);
  nand ginst8166 (P1_U5080, P1_U3040, P1_U3469);
  nand ginst8167 (P1_U5081, P1_R1162_U73, P1_U3038);
  nand ginst8168 (P1_U5082, P1_U5079, P1_U5080, P1_U5081);
  nand ginst8169 (P1_U5083, P1_U3044, P1_U5082);
  nand ginst8170 (P1_U5084, P1_R1105_U73, P1_U3043);
  nand ginst8171 (P1_U5085, P1_REG3_REG_4__SCAN_IN, P1_U3086);
  nand ginst8172 (P1_U5086, P1_U3041, P1_U3469);
  nand ginst8173 (P1_U5087, P1_R1162_U73, P1_U3039);
  nand ginst8174 (P1_U5088, P1_ADDR_REG_4__SCAN_IN, P1_U4932);
  nand ginst8175 (P1_U5089, P1_R1105_U74, P1_U3042);
  nand ginst8176 (P1_U5090, P1_U3040, P1_U3466);
  nand ginst8177 (P1_U5091, P1_R1162_U74, P1_U3038);
  nand ginst8178 (P1_U5092, P1_U5089, P1_U5090, P1_U5091);
  nand ginst8179 (P1_U5093, P1_U3044, P1_U5092);
  nand ginst8180 (P1_U5094, P1_R1105_U74, P1_U3043);
  nand ginst8181 (P1_U5095, P1_REG3_REG_3__SCAN_IN, P1_U3086);
  nand ginst8182 (P1_U5096, P1_U3041, P1_U3466);
  nand ginst8183 (P1_U5097, P1_R1162_U74, P1_U3039);
  nand ginst8184 (P1_U5098, P1_ADDR_REG_3__SCAN_IN, P1_U4932);
  nand ginst8185 (P1_U5099, P1_R1105_U14, P1_U3042);
  nand ginst8186 (P1_U5100, P1_U3040, P1_U3463);
  nand ginst8187 (P1_U5101, P1_R1162_U14, P1_U3038);
  nand ginst8188 (P1_U5102, P1_U5099, P1_U5100, P1_U5101);
  nand ginst8189 (P1_U5103, P1_U3044, P1_U5102);
  nand ginst8190 (P1_U5104, P1_R1105_U14, P1_U3043);
  nand ginst8191 (P1_U5105, P1_REG3_REG_2__SCAN_IN, P1_U3086);
  nand ginst8192 (P1_U5106, P1_U3041, P1_U3463);
  nand ginst8193 (P1_U5107, P1_R1162_U14, P1_U3039);
  nand ginst8194 (P1_U5108, P1_ADDR_REG_2__SCAN_IN, P1_U4932);
  nand ginst8195 (P1_U5109, P1_R1105_U68, P1_U3042);
  nand ginst8196 (P1_U5110, P1_U3040, P1_U3460);
  nand ginst8197 (P1_U5111, P1_R1162_U68, P1_U3038);
  nand ginst8198 (P1_U5112, P1_U5109, P1_U5110, P1_U5111);
  nand ginst8199 (P1_U5113, P1_U3044, P1_U5112);
  nand ginst8200 (P1_U5114, P1_R1105_U68, P1_U3043);
  nand ginst8201 (P1_U5115, P1_REG3_REG_1__SCAN_IN, P1_U3086);
  nand ginst8202 (P1_U5116, P1_U3041, P1_U3460);
  nand ginst8203 (P1_U5117, P1_R1162_U68, P1_U3039);
  nand ginst8204 (P1_U5118, P1_ADDR_REG_1__SCAN_IN, P1_U4932);
  nand ginst8205 (P1_U5119, P1_R1105_U69, P1_U3042);
  nand ginst8206 (P1_U5120, P1_U3040, P1_U3454);
  nand ginst8207 (P1_U5121, P1_R1162_U69, P1_U3038);
  nand ginst8208 (P1_U5122, P1_U5119, P1_U5120, P1_U5121);
  nand ginst8209 (P1_U5123, P1_U3044, P1_U5122);
  nand ginst8210 (P1_U5124, P1_R1105_U69, P1_U3043);
  nand ginst8211 (P1_U5125, P1_REG3_REG_0__SCAN_IN, P1_U3086);
  nand ginst8212 (P1_U5126, P1_U3041, P1_U3454);
  nand ginst8213 (P1_U5127, P1_R1162_U69, P1_U3039);
  nand ginst8214 (P1_U5128, P1_ADDR_REG_0__SCAN_IN, P1_U4932);
  not ginst8215 (P1_U5129, P1_U3991);
  nand ginst8216 (P1_U5130, P1_U3990, P1_U6276, P1_U6277);
  nand ginst8217 (P1_U5131, P1_U3370, P1_U3373);
  nand ginst8218 (P1_U5132, P1_U3451, P1_U5802);
  nand ginst8219 (P1_U5133, P1_U3422, P1_U5132);
  nand ginst8220 (P1_U5134, P1_U5772, P1_U6278, P1_U6279);
  nand ginst8221 (P1_U5135, P1_U3845, P1_U6280, P1_U6281);
  nand ginst8222 (P1_U5136, P1_U3022, P1_U3432, P1_U4029);
  nand ginst8223 (P1_U5137, P1_U4043, P1_U5134);
  nand ginst8224 (P1_U5138, P1_B_REG_SCAN_IN, P1_U5135);
  nand ginst8225 (P1_U5139, P1_U3037, P1_U3079);
  nand ginst8226 (P1_U5140, P1_U3035, P1_U3073);
  nand ginst8227 (P1_U5141, P1_ADD_99_U73, P1_U3434);
  nand ginst8228 (P1_U5142, P1_U5139, P1_U5140, P1_U5141);
  not ginst8229 (P1_U5143, P1_U3152);
  nand ginst8230 (P1_U5144, P1_U3423, P1_U3999);
  nand ginst8231 (P1_U5145, P1_U3848, P1_U3849, P1_U6282, P1_U6283);
  nand ginst8232 (P1_U5146, P1_U3434, P1_U5145);
  nand ginst8233 (P1_U5147, P1_U4012, P1_U5146);
  nand ginst8234 (P1_U5148, P1_U3022, P1_U5147);
  nand ginst8235 (P1_U5149, P1_U3503, P1_U5770);
  nand ginst8236 (P1_U5150, P1_ADD_99_U73, P1_U5769);
  nand ginst8237 (P1_U5151, P1_R1165_U105, P1_U3026);
  nand ginst8238 (P1_U5152, P1_U4037, P1_U5142);
  nand ginst8239 (P1_U5153, P1_REG3_REG_15__SCAN_IN, P1_U3086);
  nand ginst8240 (P1_U5154, P1_U3037, P1_U3058);
  nand ginst8241 (P1_U5155, P1_U3035, P1_U3053);
  nand ginst8242 (P1_U5156, P1_ADD_99_U62, P1_U3434);
  nand ginst8243 (P1_U5157, P1_U5154, P1_U5155, P1_U5156);
  nand ginst8244 (P1_U5158, P1_U3426, P1_U4015);
  nand ginst8245 (P1_U5159, P1_U3421, P1_U5158);
  nand ginst8246 (P1_U5160, P1_U3045, P1_U4019);
  nand ginst8247 (P1_U5161, P1_ADD_99_U62, P1_U5769);
  nand ginst8248 (P1_U5162, P1_R1165_U12, P1_U3026);
  nand ginst8249 (P1_U5163, P1_U4037, P1_U5157);
  nand ginst8250 (P1_U5164, P1_REG3_REG_26__SCAN_IN, P1_U3086);
  nand ginst8251 (P1_U5165, P1_U3037, P1_U3067);
  nand ginst8252 (P1_U5166, P1_U3035, P1_U3070);
  nand ginst8253 (P1_U5167, P1_ADD_99_U57, P1_U3434);
  nand ginst8254 (P1_U5168, P1_U5165, P1_U5166, P1_U5167);
  nand ginst8255 (P1_U5169, P1_U3476, P1_U5770);
  nand ginst8256 (P1_U5170, P1_ADD_99_U57, P1_U5769);
  nand ginst8257 (P1_U5171, P1_R1165_U90, P1_U3026);
  nand ginst8258 (P1_U5172, P1_U4037, P1_U5168);
  nand ginst8259 (P1_U5173, P1_REG3_REG_6__SCAN_IN, P1_U3086);
  nand ginst8260 (P1_U5174, P1_U3037, P1_U3069);
  nand ginst8261 (P1_U5175, P1_U3035, P1_U3081);
  nand ginst8262 (P1_U5176, P1_ADD_99_U70, P1_U3434);
  nand ginst8263 (P1_U5177, P1_U5174, P1_U5175, P1_U5176);
  nand ginst8264 (P1_U5178, P1_U3512, P1_U5770);
  nand ginst8265 (P1_U5179, P1_ADD_99_U70, P1_U5769);
  nand ginst8266 (P1_U5180, P1_R1165_U103, P1_U3026);
  nand ginst8267 (P1_U5181, P1_U4037, P1_U5177);
  nand ginst8268 (P1_U5182, P1_REG3_REG_18__SCAN_IN, P1_U3086);
  nand ginst8269 (P1_U5183, P1_U3037, P1_U3078);
  nand ginst8270 (P1_U5184, P1_U3035, P1_U3064);
  nand ginst8271 (P1_U5185, P1_REG3_REG_2__SCAN_IN, P1_U3434);
  nand ginst8272 (P1_U5186, P1_U5183, P1_U5184, P1_U5185);
  nand ginst8273 (P1_U5187, P1_U3464, P1_U5770);
  nand ginst8274 (P1_U5188, P1_REG3_REG_2__SCAN_IN, P1_U5769);
  nand ginst8275 (P1_U5189, P1_R1165_U93, P1_U3026);
  nand ginst8276 (P1_U5190, P1_U4037, P1_U5186);
  nand ginst8277 (P1_U5191, P1_REG3_REG_2__SCAN_IN, P1_U3086);
  nand ginst8278 (P1_U5192, P1_U3037, P1_U3062);
  nand ginst8279 (P1_U5193, P1_U3035, P1_U3072);
  nand ginst8280 (P1_U5194, P1_ADD_99_U77, P1_U3434);
  nand ginst8281 (P1_U5195, P1_U5192, P1_U5193, P1_U5194);
  nand ginst8282 (P1_U5196, P1_U3491, P1_U5770);
  nand ginst8283 (P1_U5197, P1_ADD_99_U77, P1_U5769);
  nand ginst8284 (P1_U5198, P1_R1165_U108, P1_U3026);
  nand ginst8285 (P1_U5199, P1_U4037, P1_U5195);
  nand ginst8286 (P1_U5200, P1_REG3_REG_11__SCAN_IN, P1_U3086);
  nand ginst8287 (P1_U5201, P1_U3037, P1_U3075);
  nand ginst8288 (P1_U5202, P1_U3035, P1_U3066);
  nand ginst8289 (P1_U5203, P1_ADD_99_U66, P1_U3434);
  nand ginst8290 (P1_U5204, P1_U5201, P1_U5202, P1_U5203);
  nand ginst8291 (P1_U5205, P1_U3045, P1_U4023);
  nand ginst8292 (P1_U5206, P1_ADD_99_U66, P1_U5769);
  nand ginst8293 (P1_U5207, P1_R1165_U99, P1_U3026);
  nand ginst8294 (P1_U5208, P1_U4037, P1_U5204);
  nand ginst8295 (P1_U5209, P1_REG3_REG_22__SCAN_IN, P1_U3086);
  nand ginst8296 (P1_U5210, P1_U3037, P1_U3072);
  nand ginst8297 (P1_U5211, P1_U3035, P1_U3079);
  nand ginst8298 (P1_U5212, P1_ADD_99_U75, P1_U3434);
  nand ginst8299 (P1_U5213, P1_U5210, P1_U5211, P1_U5212);
  nand ginst8300 (P1_U5214, P1_U3497, P1_U5770);
  nand ginst8301 (P1_U5215, P1_ADD_99_U75, P1_U5769);
  nand ginst8302 (P1_U5216, P1_R1165_U9, P1_U3026);
  nand ginst8303 (P1_U5217, P1_U4037, P1_U5213);
  nand ginst8304 (P1_U5218, P1_REG3_REG_13__SCAN_IN, P1_U3086);
  nand ginst8305 (P1_U5219, P1_U3037, P1_U3081);
  nand ginst8306 (P1_U5220, P1_U3035, P1_U3075);
  nand ginst8307 (P1_U5221, P1_ADD_99_U68, P1_U3434);
  nand ginst8308 (P1_U5222, P1_U5219, P1_U5220, P1_U5221);
  nand ginst8309 (P1_U5223, P1_U3045, P1_U4025);
  nand ginst8310 (P1_U5224, P1_ADD_99_U68, P1_U5769);
  nand ginst8311 (P1_U5225, P1_R1165_U100, P1_U3026);
  nand ginst8312 (P1_U5226, P1_U4037, P1_U5222);
  nand ginst8313 (P1_U5227, P1_REG3_REG_20__SCAN_IN, P1_U3086);
  nand ginst8314 (P1_U5228, P1_U3433, P1_U3435);
  nand ginst8315 (P1_U5229, P1_U3434, P1_U5228);
  nand ginst8316 (P1_U5230, P1_U3050, P1_U5229);
  nand ginst8317 (P1_U5231, P1_U3035, P1_U3858);
  nand ginst8318 (P1_U5232, P1_U3456, P1_U5770);
  nand ginst8319 (P1_U5233, P1_REG3_REG_0__SCAN_IN, P1_U5230);
  nand ginst8320 (P1_U5234, P1_R1165_U87, P1_U3026);
  nand ginst8321 (P1_U5235, P1_REG3_REG_0__SCAN_IN, P1_U3086);
  nand ginst8322 (P1_U5236, P1_U3037, P1_U3084);
  nand ginst8323 (P1_U5237, P1_U3035, P1_U3062);
  nand ginst8324 (P1_U5238, P1_ADD_99_U54, P1_U3434);
  nand ginst8325 (P1_U5239, P1_U5236, P1_U5237, P1_U5238);
  nand ginst8326 (P1_U5240, P1_U3485, P1_U5770);
  nand ginst8327 (P1_U5241, P1_ADD_99_U54, P1_U5769);
  nand ginst8328 (P1_U5242, P1_R1165_U88, P1_U3026);
  nand ginst8329 (P1_U5243, P1_U4037, P1_U5239);
  nand ginst8330 (P1_U5244, P1_REG3_REG_9__SCAN_IN, P1_U3086);
  nand ginst8331 (P1_U5245, P1_U3037, P1_U3064);
  nand ginst8332 (P1_U5246, P1_U3035, P1_U3067);
  nand ginst8333 (P1_U5247, P1_ADD_99_U59, P1_U3434);
  nand ginst8334 (P1_U5248, P1_U5245, P1_U5246, P1_U5247);
  nand ginst8335 (P1_U5249, P1_U3470, P1_U5770);
  nand ginst8336 (P1_U5250, P1_ADD_99_U59, P1_U5769);
  nand ginst8337 (P1_U5251, P1_R1165_U92, P1_U3026);
  nand ginst8338 (P1_U5252, P1_U4037, P1_U5248);
  nand ginst8339 (P1_U5253, P1_REG3_REG_4__SCAN_IN, P1_U3086);
  nand ginst8340 (P1_U5254, P1_U3037, P1_U3066);
  nand ginst8341 (P1_U5255, P1_U3035, P1_U3058);
  nand ginst8342 (P1_U5256, P1_ADD_99_U64, P1_U3434);
  nand ginst8343 (P1_U5257, P1_U5254, P1_U5255, P1_U5256);
  nand ginst8344 (P1_U5258, P1_U3045, P1_U4021);
  nand ginst8345 (P1_U5259, P1_ADD_99_U64, P1_U5769);
  nand ginst8346 (P1_U5260, P1_R1165_U97, P1_U3026);
  nand ginst8347 (P1_U5261, P1_U4037, P1_U5257);
  nand ginst8348 (P1_U5262, P1_REG3_REG_24__SCAN_IN, P1_U3086);
  nand ginst8349 (P1_U5263, P1_U3037, P1_U3073);
  nand ginst8350 (P1_U5264, P1_U3035, P1_U3082);
  nand ginst8351 (P1_U5265, P1_ADD_99_U71, P1_U3434);
  nand ginst8352 (P1_U5266, P1_U5263, P1_U5264, P1_U5265);
  nand ginst8353 (P1_U5267, P1_U3509, P1_U5770);
  nand ginst8354 (P1_U5268, P1_ADD_99_U71, P1_U5769);
  nand ginst8355 (P1_U5269, P1_R1165_U10, P1_U3026);
  nand ginst8356 (P1_U5270, P1_U4037, P1_U5266);
  nand ginst8357 (P1_U5271, P1_REG3_REG_17__SCAN_IN, P1_U3086);
  nand ginst8358 (P1_U5272, P1_U3037, P1_U3060);
  nand ginst8359 (P1_U5273, P1_U3035, P1_U3071);
  nand ginst8360 (P1_U5274, P1_ADD_99_U58, P1_U3434);
  nand ginst8361 (P1_U5275, P1_U5272, P1_U5273, P1_U5274);
  nand ginst8362 (P1_U5276, P1_U3473, P1_U5770);
  nand ginst8363 (P1_U5277, P1_ADD_99_U58, P1_U5769);
  nand ginst8364 (P1_U5278, P1_R1165_U91, P1_U3026);
  nand ginst8365 (P1_U5279, P1_U4037, P1_U5275);
  nand ginst8366 (P1_U5280, P1_REG3_REG_5__SCAN_IN, P1_U3086);
  nand ginst8367 (P1_U5281, P1_U3037, P1_U3074);
  nand ginst8368 (P1_U5282, P1_U3035, P1_U3069);
  nand ginst8369 (P1_U5283, P1_ADD_99_U72, P1_U3434);
  nand ginst8370 (P1_U5284, P1_U5281, P1_U5282, P1_U5283);
  nand ginst8371 (P1_U5285, P1_U3506, P1_U5770);
  nand ginst8372 (P1_U5286, P1_ADD_99_U72, P1_U5769);
  nand ginst8373 (P1_U5287, P1_R1165_U104, P1_U3026);
  nand ginst8374 (P1_U5288, P1_U4037, P1_U5284);
  nand ginst8375 (P1_U5289, P1_REG3_REG_16__SCAN_IN, P1_U3086);
  nand ginst8376 (P1_U5290, P1_U3037, P1_U3065);
  nand ginst8377 (P1_U5291, P1_U3035, P1_U3057);
  nand ginst8378 (P1_U5292, P1_ADD_99_U63, P1_U3434);
  nand ginst8379 (P1_U5293, P1_U5290, P1_U5291, P1_U5292);
  nand ginst8380 (P1_U5294, P1_U3045, P1_U4020);
  nand ginst8381 (P1_U5295, P1_ADD_99_U63, P1_U5769);
  nand ginst8382 (P1_U5296, P1_R1165_U96, P1_U3026);
  nand ginst8383 (P1_U5297, P1_U4037, P1_U5293);
  nand ginst8384 (P1_U5298, P1_REG3_REG_25__SCAN_IN, P1_U3086);
  nand ginst8385 (P1_U5299, P1_U3037, P1_U3063);
  nand ginst8386 (P1_U5300, P1_U3035, P1_U3080);
  nand ginst8387 (P1_U5301, P1_ADD_99_U76, P1_U3434);
  nand ginst8388 (P1_U5302, P1_U5299, P1_U5300, P1_U5301);
  nand ginst8389 (P1_U5303, P1_U3494, P1_U5770);
  nand ginst8390 (P1_U5304, P1_ADD_99_U76, P1_U5769);
  nand ginst8391 (P1_U5305, P1_R1165_U107, P1_U3026);
  nand ginst8392 (P1_U5306, P1_U4037, P1_U5302);
  nand ginst8393 (P1_U5307, P1_REG3_REG_12__SCAN_IN, P1_U3086);
  nand ginst8394 (P1_U5308, P1_U3037, P1_U3076);
  nand ginst8395 (P1_U5309, P1_U3035, P1_U3061);
  nand ginst8396 (P1_U5310, P1_ADD_99_U67, P1_U3434);
  nand ginst8397 (P1_U5311, P1_U5308, P1_U5309, P1_U5310);
  nand ginst8398 (P1_U5312, P1_U3045, P1_U4024);
  nand ginst8399 (P1_U5313, P1_ADD_99_U67, P1_U5769);
  nand ginst8400 (P1_U5314, P1_R1165_U11, P1_U3026);
  nand ginst8401 (P1_U5315, P1_U4037, P1_U5311);
  nand ginst8402 (P1_U5316, P1_REG3_REG_21__SCAN_IN, P1_U3086);
  nand ginst8403 (P1_U5317, P1_U3037, P1_U3077);
  nand ginst8404 (P1_U5318, P1_U3035, P1_U3068);
  nand ginst8405 (P1_U5319, P1_REG3_REG_1__SCAN_IN, P1_U3434);
  nand ginst8406 (P1_U5320, P1_U5317, P1_U5318, P1_U5319);
  nand ginst8407 (P1_U5321, P1_U3461, P1_U5770);
  nand ginst8408 (P1_U5322, P1_REG3_REG_1__SCAN_IN, P1_U5769);
  nand ginst8409 (P1_U5323, P1_R1165_U101, P1_U3026);
  nand ginst8410 (P1_U5324, P1_U4037, P1_U5320);
  nand ginst8411 (P1_U5325, P1_REG3_REG_1__SCAN_IN, P1_U3086);
  nand ginst8412 (P1_U5326, P1_U3037, P1_U3070);
  nand ginst8413 (P1_U5327, P1_U3035, P1_U3083);
  nand ginst8414 (P1_U5328, P1_ADD_99_U55, P1_U3434);
  nand ginst8415 (P1_U5329, P1_U5326, P1_U5327, P1_U5328);
  nand ginst8416 (P1_U5330, P1_U3482, P1_U5770);
  nand ginst8417 (P1_U5331, P1_ADD_99_U55, P1_U5769);
  nand ginst8418 (P1_U5332, P1_R1165_U89, P1_U3026);
  nand ginst8419 (P1_U5333, P1_U4037, P1_U5329);
  nand ginst8420 (P1_U5334, P1_REG3_REG_8__SCAN_IN, P1_U3086);
  nand ginst8421 (P1_U5335, P1_U3037, P1_U3053);
  nand ginst8422 (P1_U5336, P1_U3035, P1_U3055);
  nand ginst8423 (P1_U5337, P1_ADD_99_U60, P1_U3434);
  nand ginst8424 (P1_U5338, P1_U5335, P1_U5336, P1_U5337);
  nand ginst8425 (P1_U5339, P1_U3045, P1_U4017);
  nand ginst8426 (P1_U5340, P1_ADD_99_U60, P1_U5769);
  nand ginst8427 (P1_U5341, P1_R1165_U94, P1_U3026);
  nand ginst8428 (P1_U5342, P1_U4037, P1_U5338);
  nand ginst8429 (P1_U5343, P1_REG3_REG_28__SCAN_IN, P1_U3086);
  nand ginst8430 (P1_U5344, P1_U3037, P1_U3082);
  nand ginst8431 (P1_U5345, P1_U3035, P1_U3076);
  nand ginst8432 (P1_U5346, P1_ADD_99_U69, P1_U3434);
  nand ginst8433 (P1_U5347, P1_U5344, P1_U5345, P1_U5346);
  nand ginst8434 (P1_U5348, P1_U3514, P1_U5770);
  nand ginst8435 (P1_U5349, P1_ADD_99_U69, P1_U5769);
  nand ginst8436 (P1_U5350, P1_R1165_U102, P1_U3026);
  nand ginst8437 (P1_U5351, P1_U4037, P1_U5347);
  nand ginst8438 (P1_U5352, P1_REG3_REG_19__SCAN_IN, P1_U3086);
  nand ginst8439 (P1_U5353, P1_U3037, P1_U3068);
  nand ginst8440 (P1_U5354, P1_U3035, P1_U3060);
  nand ginst8441 (P1_U5355, P1_ADD_99_U4, P1_U3434);
  nand ginst8442 (P1_U5356, P1_U5353, P1_U5354, P1_U5355);
  nand ginst8443 (P1_U5357, P1_U3467, P1_U5770);
  nand ginst8444 (P1_U5358, P1_ADD_99_U4, P1_U5769);
  nand ginst8445 (P1_U5359, P1_R1165_U13, P1_U3026);
  nand ginst8446 (P1_U5360, P1_U4037, P1_U5356);
  nand ginst8447 (P1_U5361, P1_REG3_REG_3__SCAN_IN, P1_U3086);
  nand ginst8448 (P1_U5362, P1_U3037, P1_U3083);
  nand ginst8449 (P1_U5363, P1_U3035, P1_U3063);
  nand ginst8450 (P1_U5364, P1_ADD_99_U78, P1_U3434);
  nand ginst8451 (P1_U5365, P1_U5362, P1_U5363, P1_U5364);
  nand ginst8452 (P1_U5366, P1_U3488, P1_U5770);
  nand ginst8453 (P1_U5367, P1_ADD_99_U78, P1_U5769);
  nand ginst8454 (P1_U5368, P1_R1165_U109, P1_U3026);
  nand ginst8455 (P1_U5369, P1_U4037, P1_U5365);
  nand ginst8456 (P1_U5370, P1_REG3_REG_10__SCAN_IN, P1_U3086);
  nand ginst8457 (P1_U5371, P1_U3037, P1_U3061);
  nand ginst8458 (P1_U5372, P1_U3035, P1_U3065);
  nand ginst8459 (P1_U5373, P1_ADD_99_U65, P1_U3434);
  nand ginst8460 (P1_U5374, P1_U5371, P1_U5372, P1_U5373);
  nand ginst8461 (P1_U5375, P1_U3045, P1_U4022);
  nand ginst8462 (P1_U5376, P1_ADD_99_U65, P1_U5769);
  nand ginst8463 (P1_U5377, P1_R1165_U98, P1_U3026);
  nand ginst8464 (P1_U5378, P1_U4037, P1_U5374);
  nand ginst8465 (P1_U5379, P1_REG3_REG_23__SCAN_IN, P1_U3086);
  nand ginst8466 (P1_U5380, P1_U3037, P1_U3080);
  nand ginst8467 (P1_U5381, P1_U3035, P1_U3074);
  nand ginst8468 (P1_U5382, P1_ADD_99_U74, P1_U3434);
  nand ginst8469 (P1_U5383, P1_U5380, P1_U5381, P1_U5382);
  nand ginst8470 (P1_U5384, P1_U3500, P1_U5770);
  nand ginst8471 (P1_U5385, P1_ADD_99_U74, P1_U5769);
  nand ginst8472 (P1_U5386, P1_R1165_U106, P1_U3026);
  nand ginst8473 (P1_U5387, P1_U4037, P1_U5383);
  nand ginst8474 (P1_U5388, P1_REG3_REG_14__SCAN_IN, P1_U3086);
  nand ginst8475 (P1_U5389, P1_U3037, P1_U3057);
  nand ginst8476 (P1_U5390, P1_U3035, P1_U3054);
  nand ginst8477 (P1_U5391, P1_ADD_99_U61, P1_U3434);
  nand ginst8478 (P1_U5392, P1_U5389, P1_U5390, P1_U5391);
  nand ginst8479 (P1_U5393, P1_U3045, P1_U4018);
  nand ginst8480 (P1_U5394, P1_ADD_99_U61, P1_U5769);
  nand ginst8481 (P1_U5395, P1_R1165_U95, P1_U3026);
  nand ginst8482 (P1_U5396, P1_U4037, P1_U5392);
  nand ginst8483 (P1_U5397, P1_REG3_REG_27__SCAN_IN, P1_U3086);
  nand ginst8484 (P1_U5398, P1_U3037, P1_U3071);
  nand ginst8485 (P1_U5399, P1_U3035, P1_U3084);
  nand ginst8486 (P1_U5400, P1_ADD_99_U56, P1_U3434);
  nand ginst8487 (P1_U5401, P1_U5398, P1_U5399, P1_U5400);
  nand ginst8488 (P1_U5402, P1_U3479, P1_U5770);
  nand ginst8489 (P1_U5403, P1_ADD_99_U56, P1_U5769);
  nand ginst8490 (P1_U5404, P1_R1165_U14, P1_U3026);
  nand ginst8491 (P1_U5405, P1_U4037, P1_U5401);
  nand ginst8492 (P1_U5406, P1_REG3_REG_7__SCAN_IN, P1_U3086);
  nand ginst8493 (P1_U5407, P1_U3377, P1_U3455);
  nand ginst8494 (P1_U5408, P1_U3449, P1_U5407);
  nand ginst8495 (P1_U5409, P1_R1165_U87, P1_U3449, P1_U5817);
  nand ginst8496 (P1_U5410, P1_U3450, P1_U3453);
  nand ginst8497 (P1_U5411, P1_U3874, P1_U4013);
  nand ginst8498 (P1_U5412, P1_U3370, P1_U3422);
  nand ginst8499 (P1_U5413, P1_U3363, P1_U3365, P1_U4006);
  nand ginst8500 (P1_U5414, P1_U3425, P1_U4041);
  nand ginst8501 (P1_U5415, P1_U3425, P1_U5413);
  not ginst8502 (P1_U5416, P1_U3436);
  nand ginst8503 (P1_U5417, P1_U4013, P1_U5416);
  nand ginst8504 (P1_U5418, P1_U3485, P1_U5417);
  nand ginst8505 (P1_U5419, P1_U3021, P1_U3083);
  nand ginst8506 (P1_U5420, P1_U3482, P1_U5417);
  nand ginst8507 (P1_U5421, P1_U3021, P1_U3084);
  nand ginst8508 (P1_U5422, P1_U3479, P1_U5417);
  nand ginst8509 (P1_U5423, P1_U3021, P1_U3070);
  nand ginst8510 (P1_U5424, P1_U3476, P1_U5417);
  nand ginst8511 (P1_U5425, P1_U3021, P1_U3071);
  nand ginst8512 (P1_U5426, P1_U3473, P1_U5417);
  nand ginst8513 (P1_U5427, P1_U3021, P1_U3067);
  nand ginst8514 (P1_U5428, P1_U3470, P1_U5417);
  nand ginst8515 (P1_U5429, P1_U3021, P1_U3060);
  nand ginst8516 (P1_U5430, P1_U3467, P1_U5417);
  nand ginst8517 (P1_U5431, P1_U3021, P1_U3064);
  nand ginst8518 (P1_U5432, P1_U4017, P1_U5417);
  nand ginst8519 (P1_U5433, P1_U3021, P1_U3054);
  nand ginst8520 (P1_U5434, P1_U4018, P1_U5417);
  nand ginst8521 (P1_U5435, P1_U3021, P1_U3053);
  nand ginst8522 (P1_U5436, P1_U4019, P1_U5417);
  nand ginst8523 (P1_U5437, P1_U3021, P1_U3057);
  nand ginst8524 (P1_U5438, P1_U4020, P1_U5417);
  nand ginst8525 (P1_U5439, P1_U3021, P1_U3058);
  nand ginst8526 (P1_U5440, P1_U4021, P1_U5417);
  nand ginst8527 (P1_U5441, P1_U3021, P1_U3065);
  nand ginst8528 (P1_U5442, P1_U4022, P1_U5417);
  nand ginst8529 (P1_U5443, P1_U3021, P1_U3066);
  nand ginst8530 (P1_U5444, P1_U4023, P1_U5417);
  nand ginst8531 (P1_U5445, P1_U3021, P1_U3061);
  nand ginst8532 (P1_U5446, P1_U4024, P1_U5417);
  nand ginst8533 (P1_U5447, P1_U3021, P1_U3075);
  nand ginst8534 (P1_U5448, P1_U4025, P1_U5417);
  nand ginst8535 (P1_U5449, P1_U3021, P1_U3076);
  nand ginst8536 (P1_U5450, P1_U3464, P1_U5417);
  nand ginst8537 (P1_U5451, P1_U3021, P1_U3068);
  nand ginst8538 (P1_U5452, P1_U3514, P1_U5417);
  nand ginst8539 (P1_U5453, P1_U3021, P1_U3081);
  nand ginst8540 (P1_U5454, P1_U3512, P1_U5417);
  nand ginst8541 (P1_U5455, P1_U3021, P1_U3082);
  nand ginst8542 (P1_U5456, P1_U3509, P1_U5417);
  nand ginst8543 (P1_U5457, P1_U3021, P1_U3069);
  nand ginst8544 (P1_U5458, P1_U3506, P1_U5417);
  nand ginst8545 (P1_U5459, P1_U3021, P1_U3073);
  nand ginst8546 (P1_U5460, P1_U3503, P1_U5417);
  nand ginst8547 (P1_U5461, P1_U3021, P1_U3074);
  nand ginst8548 (P1_U5462, P1_U3500, P1_U5417);
  nand ginst8549 (P1_U5463, P1_U3021, P1_U3079);
  nand ginst8550 (P1_U5464, P1_U3497, P1_U5417);
  nand ginst8551 (P1_U5465, P1_U3021, P1_U3080);
  nand ginst8552 (P1_U5466, P1_U3494, P1_U5417);
  nand ginst8553 (P1_U5467, P1_U3021, P1_U3072);
  nand ginst8554 (P1_U5468, P1_U3491, P1_U5417);
  nand ginst8555 (P1_U5469, P1_U3021, P1_U3063);
  nand ginst8556 (P1_U5470, P1_U3488, P1_U5417);
  nand ginst8557 (P1_U5471, P1_U3021, P1_U3062);
  nand ginst8558 (P1_U5472, P1_U3461, P1_U5417);
  nand ginst8559 (P1_U5473, P1_U3021, P1_U3078);
  nand ginst8560 (P1_U5474, P1_U3456, P1_U5417);
  nand ginst8561 (P1_U5475, P1_U3021, P1_U3077);
  nand ginst8562 (P1_U5476, P1_REG1_REG_0__SCAN_IN, P1_U4145);
  nand ginst8563 (P1_U5477, P1_U3021, P1_U3485);
  nand ginst8564 (P1_U5478, P1_U3083, P1_U3436);
  nand ginst8565 (P1_U5479, P1_U3021, P1_U3482);
  nand ginst8566 (P1_U5480, P1_U3084, P1_U3436);
  nand ginst8567 (P1_U5481, P1_U3021, P1_U3479);
  nand ginst8568 (P1_U5482, P1_U3070, P1_U3436);
  nand ginst8569 (P1_U5483, P1_U3021, P1_U3476);
  nand ginst8570 (P1_U5484, P1_U3071, P1_U3436);
  nand ginst8571 (P1_U5485, P1_U3021, P1_U3473);
  nand ginst8572 (P1_U5486, P1_U3067, P1_U3436);
  nand ginst8573 (P1_U5487, P1_U3021, P1_U3470);
  nand ginst8574 (P1_U5488, P1_U3060, P1_U3436);
  nand ginst8575 (P1_U5489, P1_U3021, P1_U3467);
  nand ginst8576 (P1_U5490, P1_U3064, P1_U3436);
  nand ginst8577 (P1_U5491, P1_U3021, P1_U4017);
  nand ginst8578 (P1_U5492, P1_U3054, P1_U3436);
  nand ginst8579 (P1_U5493, P1_U3021, P1_U4018);
  nand ginst8580 (P1_U5494, P1_U3053, P1_U3436);
  nand ginst8581 (P1_U5495, P1_U3021, P1_U4019);
  nand ginst8582 (P1_U5496, P1_U3057, P1_U3436);
  nand ginst8583 (P1_U5497, P1_U3021, P1_U4020);
  nand ginst8584 (P1_U5498, P1_U3058, P1_U3436);
  nand ginst8585 (P1_U5499, P1_U3021, P1_U4021);
  nand ginst8586 (P1_U5500, P1_U3065, P1_U3436);
  nand ginst8587 (P1_U5501, P1_U3021, P1_U4022);
  nand ginst8588 (P1_U5502, P1_U3066, P1_U3436);
  nand ginst8589 (P1_U5503, P1_U3021, P1_U4023);
  nand ginst8590 (P1_U5504, P1_U3061, P1_U3436);
  nand ginst8591 (P1_U5505, P1_U3021, P1_U4024);
  nand ginst8592 (P1_U5506, P1_U3075, P1_U3436);
  nand ginst8593 (P1_U5507, P1_U3021, P1_U4025);
  nand ginst8594 (P1_U5508, P1_U3076, P1_U3436);
  nand ginst8595 (P1_U5509, P1_U3021, P1_U3464);
  nand ginst8596 (P1_U5510, P1_U3068, P1_U3436);
  nand ginst8597 (P1_U5511, P1_U3021, P1_U3514);
  nand ginst8598 (P1_U5512, P1_U3081, P1_U3436);
  nand ginst8599 (P1_U5513, P1_U3021, P1_U3512);
  nand ginst8600 (P1_U5514, P1_U3082, P1_U3436);
  nand ginst8601 (P1_U5515, P1_U3021, P1_U3509);
  nand ginst8602 (P1_U5516, P1_U3069, P1_U3436);
  nand ginst8603 (P1_U5517, P1_U3021, P1_U3506);
  nand ginst8604 (P1_U5518, P1_U3073, P1_U3436);
  nand ginst8605 (P1_U5519, P1_U3021, P1_U3503);
  nand ginst8606 (P1_U5520, P1_U3074, P1_U3436);
  nand ginst8607 (P1_U5521, P1_U3021, P1_U3500);
  nand ginst8608 (P1_U5522, P1_U3079, P1_U3436);
  nand ginst8609 (P1_U5523, P1_U3021, P1_U3497);
  nand ginst8610 (P1_U5524, P1_U3080, P1_U3436);
  nand ginst8611 (P1_U5525, P1_U3021, P1_U3494);
  nand ginst8612 (P1_U5526, P1_U3072, P1_U3436);
  nand ginst8613 (P1_U5527, P1_U3021, P1_U3491);
  nand ginst8614 (P1_U5528, P1_U3063, P1_U3436);
  nand ginst8615 (P1_U5529, P1_U3021, P1_U3488);
  nand ginst8616 (P1_U5530, P1_U3062, P1_U3436);
  nand ginst8617 (P1_U5531, P1_U3021, P1_U3461);
  nand ginst8618 (P1_U5532, P1_U3078, P1_U3436);
  nand ginst8619 (P1_U5533, P1_U3021, P1_U3456);
  nand ginst8620 (P1_U5534, P1_U3077, P1_U3436);
  nand ginst8621 (P1_U5535, P1_U3454, P1_U4145);
  not ginst8622 (P1_U5536, P1_U3437);
  not ginst8623 (P1_U5537, P1_U3438);
  nand ginst8624 (P1_U5538, P1_U3450, P1_U5799);
  nand ginst8625 (P1_U5539, P1_U3437, P1_U3439);
  nand ginst8626 (P1_U5540, P1_U3051, P1_U5539);
  nand ginst8627 (P1_U5541, P1_U3014, P1_U3444);
  not ginst8628 (P1_U5542, P1_U3440);
  nand ginst8629 (P1_U5543, P1_U3052, P1_U5542);
  nand ginst8630 (P1_U5544, P1_U3027, P1_U3083);
  nand ginst8631 (P1_U5545, P1_U3485, P1_U5543);
  nand ginst8632 (P1_U5546, P1_U3083, P1_U5540);
  nand ginst8633 (P1_U5547, P1_U3027, P1_U3084);
  nand ginst8634 (P1_U5548, P1_U3482, P1_U5543);
  nand ginst8635 (P1_U5549, P1_U3084, P1_U5540);
  nand ginst8636 (P1_U5550, P1_U3027, P1_U3070);
  nand ginst8637 (P1_U5551, P1_U3479, P1_U5543);
  nand ginst8638 (P1_U5552, P1_U3070, P1_U5540);
  nand ginst8639 (P1_U5553, P1_U3027, P1_U3071);
  nand ginst8640 (P1_U5554, P1_U3476, P1_U5543);
  nand ginst8641 (P1_U5555, P1_U3071, P1_U5540);
  nand ginst8642 (P1_U5556, P1_U3027, P1_U3067);
  nand ginst8643 (P1_U5557, P1_U3473, P1_U5543);
  nand ginst8644 (P1_U5558, P1_U3067, P1_U5540);
  nand ginst8645 (P1_U5559, P1_U3027, P1_U3060);
  nand ginst8646 (P1_U5560, P1_U3470, P1_U5543);
  nand ginst8647 (P1_U5561, P1_U3060, P1_U5540);
  nand ginst8648 (P1_U5562, P1_R1309_U8, P1_U3027);
  nand ginst8649 (P1_U5563, P1_U4026, P1_U5543);
  nand ginst8650 (P1_U5564, P1_U3056, P1_U5540);
  nand ginst8651 (P1_U5565, P1_R1309_U6, P1_U3027);
  nand ginst8652 (P1_U5566, P1_U4027, P1_U5543);
  nand ginst8653 (P1_U5567, P1_U3059, P1_U5540);
  nand ginst8654 (P1_U5568, P1_U3027, P1_U3064);
  nand ginst8655 (P1_U5569, P1_U3467, P1_U5543);
  nand ginst8656 (P1_U5570, P1_U3064, P1_U5540);
  nand ginst8657 (P1_U5571, P1_U3027, P1_U3055);
  nand ginst8658 (P1_U5572, P1_U4028, P1_U5543);
  nand ginst8659 (P1_U5573, P1_U3055, P1_U5540);
  nand ginst8660 (P1_U5574, P1_U3027, P1_U3054);
  nand ginst8661 (P1_U5575, P1_U4017, P1_U5543);
  nand ginst8662 (P1_U5576, P1_U3054, P1_U5540);
  nand ginst8663 (P1_U5577, P1_U3027, P1_U3053);
  nand ginst8664 (P1_U5578, P1_U4018, P1_U5543);
  nand ginst8665 (P1_U5579, P1_U3053, P1_U5540);
  nand ginst8666 (P1_U5580, P1_U3027, P1_U3057);
  nand ginst8667 (P1_U5581, P1_U4019, P1_U5543);
  nand ginst8668 (P1_U5582, P1_U3057, P1_U5540);
  nand ginst8669 (P1_U5583, P1_U3027, P1_U3058);
  nand ginst8670 (P1_U5584, P1_U4020, P1_U5543);
  nand ginst8671 (P1_U5585, P1_U3058, P1_U5540);
  nand ginst8672 (P1_U5586, P1_U3027, P1_U3065);
  nand ginst8673 (P1_U5587, P1_U4021, P1_U5543);
  nand ginst8674 (P1_U5588, P1_U3065, P1_U5540);
  nand ginst8675 (P1_U5589, P1_U3027, P1_U3066);
  nand ginst8676 (P1_U5590, P1_U4022, P1_U5543);
  nand ginst8677 (P1_U5591, P1_U3066, P1_U5540);
  nand ginst8678 (P1_U5592, P1_U3027, P1_U3061);
  nand ginst8679 (P1_U5593, P1_U4023, P1_U5543);
  nand ginst8680 (P1_U5594, P1_U3061, P1_U5540);
  nand ginst8681 (P1_U5595, P1_U3027, P1_U3075);
  nand ginst8682 (P1_U5596, P1_U4024, P1_U5543);
  nand ginst8683 (P1_U5597, P1_U3075, P1_U5540);
  nand ginst8684 (P1_U5598, P1_U3027, P1_U3076);
  nand ginst8685 (P1_U5599, P1_U4025, P1_U5543);
  nand ginst8686 (P1_U5600, P1_U3076, P1_U5540);
  nand ginst8687 (P1_U5601, P1_U3027, P1_U3068);
  nand ginst8688 (P1_U5602, P1_U3464, P1_U5543);
  nand ginst8689 (P1_U5603, P1_U3068, P1_U5540);
  nand ginst8690 (P1_U5604, P1_U3027, P1_U3081);
  nand ginst8691 (P1_U5605, P1_U3514, P1_U5543);
  nand ginst8692 (P1_U5606, P1_U3081, P1_U5540);
  nand ginst8693 (P1_U5607, P1_U3027, P1_U3082);
  nand ginst8694 (P1_U5608, P1_U3512, P1_U5543);
  nand ginst8695 (P1_U5609, P1_U3082, P1_U5540);
  nand ginst8696 (P1_U5610, P1_U3027, P1_U3069);
  nand ginst8697 (P1_U5611, P1_U3509, P1_U5543);
  nand ginst8698 (P1_U5612, P1_U3069, P1_U5540);
  nand ginst8699 (P1_U5613, P1_U3027, P1_U3073);
  nand ginst8700 (P1_U5614, P1_U3506, P1_U5543);
  nand ginst8701 (P1_U5615, P1_U3073, P1_U5540);
  nand ginst8702 (P1_U5616, P1_U3027, P1_U3074);
  nand ginst8703 (P1_U5617, P1_U3503, P1_U5543);
  nand ginst8704 (P1_U5618, P1_U3074, P1_U5540);
  nand ginst8705 (P1_U5619, P1_U3027, P1_U3079);
  nand ginst8706 (P1_U5620, P1_U3500, P1_U5543);
  nand ginst8707 (P1_U5621, P1_U3079, P1_U5540);
  nand ginst8708 (P1_U5622, P1_U3027, P1_U3080);
  nand ginst8709 (P1_U5623, P1_U3497, P1_U5543);
  nand ginst8710 (P1_U5624, P1_U3080, P1_U5540);
  nand ginst8711 (P1_U5625, P1_U3027, P1_U3072);
  nand ginst8712 (P1_U5626, P1_U3494, P1_U5543);
  nand ginst8713 (P1_U5627, P1_U3072, P1_U5540);
  nand ginst8714 (P1_U5628, P1_U3027, P1_U3063);
  nand ginst8715 (P1_U5629, P1_U3491, P1_U5543);
  nand ginst8716 (P1_U5630, P1_U3063, P1_U5540);
  nand ginst8717 (P1_U5631, P1_U3027, P1_U3062);
  nand ginst8718 (P1_U5632, P1_U3488, P1_U5543);
  nand ginst8719 (P1_U5633, P1_U3062, P1_U5540);
  nand ginst8720 (P1_U5634, P1_U3027, P1_U3078);
  nand ginst8721 (P1_U5635, P1_U3461, P1_U5543);
  nand ginst8722 (P1_U5636, P1_U3078, P1_U5540);
  nand ginst8723 (P1_U5637, P1_U3027, P1_U3077);
  nand ginst8724 (P1_U5638, P1_U3456, P1_U5543);
  nand ginst8725 (P1_U5639, P1_U3077, P1_U5540);
  nand ginst8726 (P1_U5640, P1_U3439, P1_U3440);
  nand ginst8727 (P1_U5641, P1_U3052, P1_U5640);
  nand ginst8728 (P1_U5642, P1_U3028, P1_U3083);
  nand ginst8729 (P1_U5643, P1_U3438, P1_U3485);
  nand ginst8730 (P1_U5644, P1_U3083, P1_U5641);
  nand ginst8731 (P1_U5645, P1_U3084, P1_U5786);
  nand ginst8732 (P1_U5646, P1_U3028, P1_U3084);
  nand ginst8733 (P1_U5647, P1_U3438, P1_U3482);
  nand ginst8734 (P1_U5648, P1_U3084, P1_U5641);
  nand ginst8735 (P1_U5649, P1_U3070, P1_U5786);
  nand ginst8736 (P1_U5650, P1_U3028, P1_U3070);
  nand ginst8737 (P1_U5651, P1_U3438, P1_U3479);
  nand ginst8738 (P1_U5652, P1_U3070, P1_U5641);
  nand ginst8739 (P1_U5653, P1_U3071, P1_U5786);
  nand ginst8740 (P1_U5654, P1_U3028, P1_U3071);
  nand ginst8741 (P1_U5655, P1_U3438, P1_U3476);
  nand ginst8742 (P1_U5656, P1_U3071, P1_U5641);
  nand ginst8743 (P1_U5657, P1_U3067, P1_U5786);
  nand ginst8744 (P1_U5658, P1_U3028, P1_U3067);
  nand ginst8745 (P1_U5659, P1_U3438, P1_U3473);
  nand ginst8746 (P1_U5660, P1_U3067, P1_U5641);
  nand ginst8747 (P1_U5661, P1_U3060, P1_U5786);
  nand ginst8748 (P1_U5662, P1_U3028, P1_U3060);
  nand ginst8749 (P1_U5663, P1_U3438, P1_U3470);
  nand ginst8750 (P1_U5664, P1_U3060, P1_U5641);
  nand ginst8751 (P1_U5665, P1_U3064, P1_U5786);
  nand ginst8752 (P1_U5666, P1_R1309_U8, P1_U3028);
  nand ginst8753 (P1_U5667, P1_U3438, P1_U4026);
  nand ginst8754 (P1_U5668, P1_U3056, P1_U5641);
  nand ginst8755 (P1_U5669, P1_R1309_U6, P1_U3028);
  nand ginst8756 (P1_U5670, P1_U3438, P1_U4027);
  nand ginst8757 (P1_U5671, P1_U3059, P1_U5641);
  nand ginst8758 (P1_U5672, P1_U3028, P1_U3064);
  nand ginst8759 (P1_U5673, P1_U3438, P1_U3467);
  nand ginst8760 (P1_U5674, P1_U3064, P1_U5641);
  nand ginst8761 (P1_U5675, P1_U3068, P1_U5786);
  nand ginst8762 (P1_U5676, P1_U3028, P1_U3055);
  nand ginst8763 (P1_U5677, P1_U3438, P1_U4028);
  nand ginst8764 (P1_U5678, P1_U3055, P1_U5641);
  nand ginst8765 (P1_U5679, P1_U3054, P1_U5786);
  nand ginst8766 (P1_U5680, P1_U3028, P1_U3054);
  nand ginst8767 (P1_U5681, P1_U3438, P1_U4017);
  nand ginst8768 (P1_U5682, P1_U3054, P1_U5641);
  nand ginst8769 (P1_U5683, P1_U3053, P1_U5786);
  nand ginst8770 (P1_U5684, P1_U3028, P1_U3053);
  nand ginst8771 (P1_U5685, P1_U3438, P1_U4018);
  nand ginst8772 (P1_U5686, P1_U3053, P1_U5641);
  nand ginst8773 (P1_U5687, P1_U3057, P1_U5786);
  nand ginst8774 (P1_U5688, P1_U3028, P1_U3057);
  nand ginst8775 (P1_U5689, P1_U3438, P1_U4019);
  nand ginst8776 (P1_U5690, P1_U3057, P1_U5641);
  nand ginst8777 (P1_U5691, P1_U3058, P1_U5786);
  nand ginst8778 (P1_U5692, P1_U3028, P1_U3058);
  nand ginst8779 (P1_U5693, P1_U3438, P1_U4020);
  nand ginst8780 (P1_U5694, P1_U3058, P1_U5641);
  nand ginst8781 (P1_U5695, P1_U3065, P1_U5786);
  nand ginst8782 (P1_U5696, P1_U3028, P1_U3065);
  nand ginst8783 (P1_U5697, P1_U3438, P1_U4021);
  nand ginst8784 (P1_U5698, P1_U3065, P1_U5641);
  nand ginst8785 (P1_U5699, P1_U3066, P1_U5786);
  nand ginst8786 (P1_U5700, P1_U3028, P1_U3066);
  nand ginst8787 (P1_U5701, P1_U3438, P1_U4022);
  nand ginst8788 (P1_U5702, P1_U3066, P1_U5641);
  nand ginst8789 (P1_U5703, P1_U3061, P1_U5786);
  nand ginst8790 (P1_U5704, P1_U3028, P1_U3061);
  nand ginst8791 (P1_U5705, P1_U3438, P1_U4023);
  nand ginst8792 (P1_U5706, P1_U3061, P1_U5641);
  nand ginst8793 (P1_U5707, P1_U3075, P1_U5786);
  nand ginst8794 (P1_U5708, P1_U3028, P1_U3075);
  nand ginst8795 (P1_U5709, P1_U3438, P1_U4024);
  nand ginst8796 (P1_U5710, P1_U3075, P1_U5641);
  nand ginst8797 (P1_U5711, P1_U3076, P1_U5786);
  nand ginst8798 (P1_U5712, P1_U3028, P1_U3076);
  nand ginst8799 (P1_U5713, P1_U3438, P1_U4025);
  nand ginst8800 (P1_U5714, P1_U3076, P1_U5641);
  nand ginst8801 (P1_U5715, P1_U3081, P1_U5786);
  nand ginst8802 (P1_U5716, P1_U3028, P1_U3068);
  nand ginst8803 (P1_U5717, P1_U3438, P1_U3464);
  nand ginst8804 (P1_U5718, P1_U3068, P1_U5641);
  nand ginst8805 (P1_U5719, P1_U3078, P1_U5786);
  nand ginst8806 (P1_U5720, P1_U3028, P1_U3081);
  nand ginst8807 (P1_U5721, P1_U3438, P1_U3514);
  nand ginst8808 (P1_U5722, P1_U3081, P1_U5641);
  nand ginst8809 (P1_U5723, P1_U3082, P1_U5786);
  nand ginst8810 (P1_U5724, P1_U3028, P1_U3082);
  nand ginst8811 (P1_U5725, P1_U3438, P1_U3512);
  nand ginst8812 (P1_U5726, P1_U3082, P1_U5641);
  nand ginst8813 (P1_U5727, P1_U3069, P1_U5786);
  nand ginst8814 (P1_U5728, P1_U3028, P1_U3069);
  nand ginst8815 (P1_U5729, P1_U3438, P1_U3509);
  nand ginst8816 (P1_U5730, P1_U3069, P1_U5641);
  nand ginst8817 (P1_U5731, P1_U3073, P1_U5786);
  nand ginst8818 (P1_U5732, P1_U3028, P1_U3073);
  nand ginst8819 (P1_U5733, P1_U3438, P1_U3506);
  nand ginst8820 (P1_U5734, P1_U3073, P1_U5641);
  nand ginst8821 (P1_U5735, P1_U3074, P1_U5786);
  nand ginst8822 (P1_U5736, P1_U3028, P1_U3074);
  nand ginst8823 (P1_U5737, P1_U3438, P1_U3503);
  nand ginst8824 (P1_U5738, P1_U3074, P1_U5641);
  nand ginst8825 (P1_U5739, P1_U3079, P1_U5786);
  nand ginst8826 (P1_U5740, P1_U3028, P1_U3079);
  nand ginst8827 (P1_U5741, P1_U3438, P1_U3500);
  nand ginst8828 (P1_U5742, P1_U3079, P1_U5641);
  nand ginst8829 (P1_U5743, P1_U3080, P1_U5786);
  nand ginst8830 (P1_U5744, P1_U3028, P1_U3080);
  nand ginst8831 (P1_U5745, P1_U3438, P1_U3497);
  nand ginst8832 (P1_U5746, P1_U3080, P1_U5641);
  nand ginst8833 (P1_U5747, P1_U3072, P1_U5786);
  nand ginst8834 (P1_U5748, P1_U3028, P1_U3072);
  nand ginst8835 (P1_U5749, P1_U3438, P1_U3494);
  nand ginst8836 (P1_U5750, P1_U3072, P1_U5641);
  nand ginst8837 (P1_U5751, P1_U3063, P1_U5786);
  nand ginst8838 (P1_U5752, P1_U3028, P1_U3063);
  nand ginst8839 (P1_U5753, P1_U3438, P1_U3491);
  nand ginst8840 (P1_U5754, P1_U3063, P1_U5641);
  nand ginst8841 (P1_U5755, P1_U3062, P1_U5786);
  nand ginst8842 (P1_U5756, P1_U3028, P1_U3062);
  nand ginst8843 (P1_U5757, P1_U3438, P1_U3488);
  nand ginst8844 (P1_U5758, P1_U3062, P1_U5641);
  nand ginst8845 (P1_U5759, P1_U3083, P1_U5786);
  nand ginst8846 (P1_U5760, P1_U3028, P1_U3078);
  nand ginst8847 (P1_U5761, P1_U3438, P1_U3461);
  nand ginst8848 (P1_U5762, P1_U3078, P1_U5641);
  nand ginst8849 (P1_U5763, P1_U3077, P1_U5786);
  nand ginst8850 (P1_U5764, P1_U3028, P1_U3077);
  nand ginst8851 (P1_U5765, P1_U3438, P1_U3456);
  nand ginst8852 (P1_U5766, P1_U3077, P1_U5641);
  nand ginst8853 (P1_U5767, P1_U3434, P1_U4038);
  nand ginst8854 (P1_U5768, P1_U4015, P1_U4038);
  nand ginst8855 (P1_U5769, P1_U3050, P1_U5767);
  nand ginst8856 (P1_U5770, P1_U4039, P1_U5768);
  nand ginst8857 (P1_U5771, P1_U5775, P1_U5781);
  nand ginst8858 (P1_U5772, P1_R1375_U9, P1_U5131);
  nand ginst8859 (P1_U5773, P1_IR_REG_24__SCAN_IN, P1_U3952);
  nand ginst8860 (P1_U5774, P1_IR_REG_31__SCAN_IN, P1_SUB_88_U17);
  not ginst8861 (P1_U5775, P1_U3441);
  nand ginst8862 (P1_U5776, P1_IR_REG_25__SCAN_IN, P1_U3952);
  nand ginst8863 (P1_U5777, P1_IR_REG_31__SCAN_IN, P1_SUB_88_U170);
  not ginst8864 (P1_U5778, P1_U3442);
  nand ginst8865 (P1_U5779, P1_IR_REG_26__SCAN_IN, P1_U3952);
  nand ginst8866 (P1_U5780, P1_IR_REG_31__SCAN_IN, P1_SUB_88_U18);
  not ginst8867 (P1_U5781, P1_U3443);
  nand ginst8868 (P1_U5782, P1_U3359, P1_U3441);
  nand ginst8869 (P1_U5783, P1_B_REG_SCAN_IN, P1_U4046, P1_U5775);
  nand ginst8870 (P1_U5784, P1_IR_REG_23__SCAN_IN, P1_U3952);
  nand ginst8871 (P1_U5785, P1_IR_REG_31__SCAN_IN, P1_SUB_88_U16);
  not ginst8872 (P1_U5786, P1_U3444);
  nand ginst8873 (P1_U5787, P1_D_REG_0__SCAN_IN, P1_U3953);
  nand ginst8874 (P1_U5788, P1_U4034, P1_U4146);
  nand ginst8875 (P1_U5789, P1_D_REG_1__SCAN_IN, P1_U3953);
  nand ginst8876 (P1_U5790, P1_U4034, P1_U4147);
  nand ginst8877 (P1_U5791, P1_IR_REG_22__SCAN_IN, P1_U3952);
  nand ginst8878 (P1_U5792, P1_IR_REG_31__SCAN_IN, P1_SUB_88_U15);
  not ginst8879 (P1_U5793, P1_U3451);
  nand ginst8880 (P1_U5794, P1_IR_REG_19__SCAN_IN, P1_U3952);
  nand ginst8881 (P1_U5795, P1_IR_REG_31__SCAN_IN, P1_SUB_88_U13);
  not ginst8882 (P1_U5796, P1_U3452);
  nand ginst8883 (P1_U5797, P1_IR_REG_20__SCAN_IN, P1_U3952);
  nand ginst8884 (P1_U5798, P1_IR_REG_31__SCAN_IN, P1_SUB_88_U14);
  not ginst8885 (P1_U5799, P1_U3453);
  nand ginst8886 (P1_U5800, P1_IR_REG_21__SCAN_IN, P1_U3952);
  nand ginst8887 (P1_U5801, P1_IR_REG_31__SCAN_IN, P1_SUB_88_U173);
  not ginst8888 (P1_U5802, P1_U3450);
  nand ginst8889 (P1_U5803, P1_IR_REG_30__SCAN_IN, P1_U3952);
  nand ginst8890 (P1_U5804, P1_IR_REG_31__SCAN_IN, P1_SUB_88_U165);
  not ginst8891 (P1_U5805, P1_U3447);
  nand ginst8892 (P1_U5806, P1_IR_REG_29__SCAN_IN, P1_U3952);
  nand ginst8893 (P1_U5807, P1_IR_REG_31__SCAN_IN, P1_SUB_88_U20);
  not ginst8894 (P1_U5808, P1_U3448);
  nand ginst8895 (P1_U5809, P1_IR_REG_28__SCAN_IN, P1_U3952);
  nand ginst8896 (P1_U5810, P1_IR_REG_31__SCAN_IN, P1_SUB_88_U19);
  not ginst8897 (P1_U5811, P1_U3449);
  nand ginst8898 (P1_U5812, P1_IR_REG_0__SCAN_IN, P1_U3952);
  nand ginst8899 (P1_U5813, P1_IR_REG_0__SCAN_IN, P1_IR_REG_31__SCAN_IN);
  not ginst8900 (P1_U5814, P1_U3454);
  nand ginst8901 (P1_U5815, P1_IR_REG_27__SCAN_IN, P1_U3952);
  nand ginst8902 (P1_U5816, P1_IR_REG_31__SCAN_IN, P1_SUB_88_U42);
  not ginst8903 (P1_U5817, P1_U3455);
  nand ginst8904 (P1_U5818, P1_U3954, U125);
  nand ginst8905 (P1_U5819, P1_U3454, P1_U4014);
  not ginst8906 (P1_U5820, P1_U3456);
  nand ginst8907 (P1_U5821, P1_U3451, P1_U5802);
  nand ginst8908 (P1_U5822, P1_U4178, P1_U5793);
  nand ginst8909 (P1_U5823, P1_D_REG_1__SCAN_IN, P1_U4144);
  nand ginst8910 (P1_U5824, P1_U3360, P1_U4147);
  not ginst8911 (P1_U5825, P1_U3458);
  nand ginst8912 (P1_U5826, P1_U3360, P1_U5771);
  nand ginst8913 (P1_U5827, P1_D_REG_0__SCAN_IN, P1_U4144);
  not ginst8914 (P1_U5828, P1_U3457);
  nand ginst8915 (P1_U5829, P1_REG0_REG_0__SCAN_IN, P1_U3955);
  nand ginst8916 (P1_U5830, P1_U4033, P1_U4198);
  nand ginst8917 (P1_U5831, P1_IR_REG_1__SCAN_IN, P1_U3952);
  nand ginst8918 (P1_U5832, P1_IR_REG_31__SCAN_IN, P1_SUB_88_U40);
  nand ginst8919 (P1_U5833, P1_U3954, U114);
  nand ginst8920 (P1_U5834, P1_U3460, P1_U4014);
  not ginst8921 (P1_U5835, P1_U3461);
  nand ginst8922 (P1_U5836, P1_REG0_REG_1__SCAN_IN, P1_U3955);
  nand ginst8923 (P1_U5837, P1_U4033, P1_U4222);
  nand ginst8924 (P1_U5838, P1_IR_REG_2__SCAN_IN, P1_U3952);
  nand ginst8925 (P1_U5839, P1_IR_REG_31__SCAN_IN, P1_SUB_88_U21);
  nand ginst8926 (P1_U5840, P1_U3954, U103);
  nand ginst8927 (P1_U5841, P1_U3463, P1_U4014);
  not ginst8928 (P1_U5842, P1_U3464);
  nand ginst8929 (P1_U5843, P1_REG0_REG_2__SCAN_IN, P1_U3955);
  nand ginst8930 (P1_U5844, P1_U4033, P1_U4241);
  nand ginst8931 (P1_U5845, P1_IR_REG_3__SCAN_IN, P1_U3952);
  nand ginst8932 (P1_U5846, P1_IR_REG_31__SCAN_IN, P1_SUB_88_U22);
  nand ginst8933 (P1_U5847, P1_U3954, U100);
  nand ginst8934 (P1_U5848, P1_U3466, P1_U4014);
  not ginst8935 (P1_U5849, P1_U3467);
  nand ginst8936 (P1_U5850, P1_REG0_REG_3__SCAN_IN, P1_U3955);
  nand ginst8937 (P1_U5851, P1_U4033, P1_U4260);
  nand ginst8938 (P1_U5852, P1_IR_REG_4__SCAN_IN, P1_U3952);
  nand ginst8939 (P1_U5853, P1_IR_REG_31__SCAN_IN, P1_SUB_88_U23);
  nand ginst8940 (P1_U5854, P1_U3954, U99);
  nand ginst8941 (P1_U5855, P1_U3469, P1_U4014);
  not ginst8942 (P1_U5856, P1_U3470);
  nand ginst8943 (P1_U5857, P1_REG0_REG_4__SCAN_IN, P1_U3955);
  nand ginst8944 (P1_U5858, P1_U4033, P1_U4279);
  nand ginst8945 (P1_U5859, P1_IR_REG_5__SCAN_IN, P1_U3952);
  nand ginst8946 (P1_U5860, P1_IR_REG_31__SCAN_IN, P1_SUB_88_U162);
  nand ginst8947 (P1_U5861, P1_U3954, U98);
  nand ginst8948 (P1_U5862, P1_U3472, P1_U4014);
  not ginst8949 (P1_U5863, P1_U3473);
  nand ginst8950 (P1_U5864, P1_REG0_REG_5__SCAN_IN, P1_U3955);
  nand ginst8951 (P1_U5865, P1_U4033, P1_U4298);
  nand ginst8952 (P1_U5866, P1_IR_REG_6__SCAN_IN, P1_U3952);
  nand ginst8953 (P1_U5867, P1_IR_REG_31__SCAN_IN, P1_SUB_88_U24);
  nand ginst8954 (P1_U5868, P1_U3954, U97);
  nand ginst8955 (P1_U5869, P1_U3475, P1_U4014);
  not ginst8956 (P1_U5870, P1_U3476);
  nand ginst8957 (P1_U5871, P1_REG0_REG_6__SCAN_IN, P1_U3955);
  nand ginst8958 (P1_U5872, P1_U4033, P1_U4317);
  nand ginst8959 (P1_U5873, P1_IR_REG_7__SCAN_IN, P1_U3952);
  nand ginst8960 (P1_U5874, P1_IR_REG_31__SCAN_IN, P1_SUB_88_U25);
  nand ginst8961 (P1_U5875, P1_U3954, U96);
  nand ginst8962 (P1_U5876, P1_U3478, P1_U4014);
  not ginst8963 (P1_U5877, P1_U3479);
  nand ginst8964 (P1_U5878, P1_REG0_REG_7__SCAN_IN, P1_U3955);
  nand ginst8965 (P1_U5879, P1_U4033, P1_U4336);
  nand ginst8966 (P1_U5880, P1_IR_REG_8__SCAN_IN, P1_U3952);
  nand ginst8967 (P1_U5881, P1_IR_REG_31__SCAN_IN, P1_SUB_88_U26);
  nand ginst8968 (P1_U5882, P1_U3954, U95);
  nand ginst8969 (P1_U5883, P1_U3481, P1_U4014);
  not ginst8970 (P1_U5884, P1_U3482);
  nand ginst8971 (P1_U5885, P1_REG0_REG_8__SCAN_IN, P1_U3955);
  nand ginst8972 (P1_U5886, P1_U4033, P1_U4355);
  nand ginst8973 (P1_U5887, P1_IR_REG_9__SCAN_IN, P1_U3952);
  nand ginst8974 (P1_U5888, P1_IR_REG_31__SCAN_IN, P1_SUB_88_U160);
  nand ginst8975 (P1_U5889, P1_U3954, U94);
  nand ginst8976 (P1_U5890, P1_U3484, P1_U4014);
  not ginst8977 (P1_U5891, P1_U3485);
  nand ginst8978 (P1_U5892, P1_REG0_REG_9__SCAN_IN, P1_U3955);
  nand ginst8979 (P1_U5893, P1_U4033, P1_U4374);
  nand ginst8980 (P1_U5894, P1_IR_REG_10__SCAN_IN, P1_U3952);
  nand ginst8981 (P1_U5895, P1_IR_REG_31__SCAN_IN, P1_SUB_88_U6);
  nand ginst8982 (P1_U5896, P1_U3954, U124);
  nand ginst8983 (P1_U5897, P1_U3487, P1_U4014);
  not ginst8984 (P1_U5898, P1_U3488);
  nand ginst8985 (P1_U5899, P1_REG0_REG_10__SCAN_IN, P1_U3955);
  nand ginst8986 (P1_U5900, P1_U4033, P1_U4393);
  nand ginst8987 (P1_U5901, P1_IR_REG_11__SCAN_IN, P1_U3952);
  nand ginst8988 (P1_U5902, P1_IR_REG_31__SCAN_IN, P1_SUB_88_U7);
  nand ginst8989 (P1_U5903, P1_U3954, U123);
  nand ginst8990 (P1_U5904, P1_U3490, P1_U4014);
  not ginst8991 (P1_U5905, P1_U3491);
  nand ginst8992 (P1_U5906, P1_REG0_REG_11__SCAN_IN, P1_U3955);
  nand ginst8993 (P1_U5907, P1_U4033, P1_U4412);
  nand ginst8994 (P1_U5908, P1_IR_REG_12__SCAN_IN, P1_U3952);
  nand ginst8995 (P1_U5909, P1_IR_REG_31__SCAN_IN, P1_SUB_88_U8);
  nand ginst8996 (P1_U5910, P1_U3954, U122);
  nand ginst8997 (P1_U5911, P1_U3493, P1_U4014);
  not ginst8998 (P1_U5912, P1_U3494);
  nand ginst8999 (P1_U5913, P1_REG0_REG_12__SCAN_IN, P1_U3955);
  nand ginst9000 (P1_U5914, P1_U4033, P1_U4431);
  nand ginst9001 (P1_U5915, P1_IR_REG_13__SCAN_IN, P1_U3952);
  nand ginst9002 (P1_U5916, P1_IR_REG_31__SCAN_IN, P1_SUB_88_U179);
  nand ginst9003 (P1_U5917, P1_U3954, U121);
  nand ginst9004 (P1_U5918, P1_U3496, P1_U4014);
  not ginst9005 (P1_U5919, P1_U3497);
  nand ginst9006 (P1_U5920, P1_REG0_REG_13__SCAN_IN, P1_U3955);
  nand ginst9007 (P1_U5921, P1_U4033, P1_U4450);
  nand ginst9008 (P1_U5922, P1_IR_REG_14__SCAN_IN, P1_U3952);
  nand ginst9009 (P1_U5923, P1_IR_REG_31__SCAN_IN, P1_SUB_88_U9);
  nand ginst9010 (P1_U5924, P1_U3954, U120);
  nand ginst9011 (P1_U5925, P1_U3499, P1_U4014);
  not ginst9012 (P1_U5926, P1_U3500);
  nand ginst9013 (P1_U5927, P1_REG0_REG_14__SCAN_IN, P1_U3955);
  nand ginst9014 (P1_U5928, P1_U4033, P1_U4469);
  nand ginst9015 (P1_U5929, P1_IR_REG_15__SCAN_IN, P1_U3952);
  nand ginst9016 (P1_U5930, P1_IR_REG_31__SCAN_IN, P1_SUB_88_U10);
  nand ginst9017 (P1_U5931, P1_U3954, U119);
  nand ginst9018 (P1_U5932, P1_U3502, P1_U4014);
  not ginst9019 (P1_U5933, P1_U3503);
  nand ginst9020 (P1_U5934, P1_REG0_REG_15__SCAN_IN, P1_U3955);
  nand ginst9021 (P1_U5935, P1_U4033, P1_U4488);
  nand ginst9022 (P1_U5936, P1_IR_REG_16__SCAN_IN, P1_U3952);
  nand ginst9023 (P1_U5937, P1_IR_REG_31__SCAN_IN, P1_SUB_88_U11);
  nand ginst9024 (P1_U5938, P1_U3954, U118);
  nand ginst9025 (P1_U5939, P1_U3505, P1_U4014);
  not ginst9026 (P1_U5940, P1_U3506);
  nand ginst9027 (P1_U5941, P1_REG0_REG_16__SCAN_IN, P1_U3955);
  nand ginst9028 (P1_U5942, P1_U4033, P1_U4507);
  nand ginst9029 (P1_U5943, P1_IR_REG_17__SCAN_IN, P1_U3952);
  nand ginst9030 (P1_U5944, P1_IR_REG_31__SCAN_IN, P1_SUB_88_U177);
  nand ginst9031 (P1_U5945, P1_U3954, U117);
  nand ginst9032 (P1_U5946, P1_U3508, P1_U4014);
  not ginst9033 (P1_U5947, P1_U3509);
  nand ginst9034 (P1_U5948, P1_REG0_REG_17__SCAN_IN, P1_U3955);
  nand ginst9035 (P1_U5949, P1_U4033, P1_U4526);
  nand ginst9036 (P1_U5950, P1_IR_REG_18__SCAN_IN, P1_U3952);
  nand ginst9037 (P1_U5951, P1_IR_REG_31__SCAN_IN, P1_SUB_88_U12);
  nand ginst9038 (P1_U5952, P1_U3954, U116);
  nand ginst9039 (P1_U5953, P1_U3511, P1_U4014);
  not ginst9040 (P1_U5954, P1_U3512);
  nand ginst9041 (P1_U5955, P1_REG0_REG_18__SCAN_IN, P1_U3955);
  nand ginst9042 (P1_U5956, P1_U4033, P1_U4545);
  nand ginst9043 (P1_U5957, P1_U3954, U115);
  nand ginst9044 (P1_U5958, P1_U3452, P1_U4014);
  not ginst9045 (P1_U5959, P1_U3514);
  nand ginst9046 (P1_U5960, P1_REG0_REG_19__SCAN_IN, P1_U3955);
  nand ginst9047 (P1_U5961, P1_U4033, P1_U4564);
  nand ginst9048 (P1_U5962, P1_REG0_REG_20__SCAN_IN, P1_U3955);
  nand ginst9049 (P1_U5963, P1_U4033, P1_U4583);
  nand ginst9050 (P1_U5964, P1_REG0_REG_21__SCAN_IN, P1_U3955);
  nand ginst9051 (P1_U5965, P1_U4033, P1_U4602);
  nand ginst9052 (P1_U5966, P1_REG0_REG_22__SCAN_IN, P1_U3955);
  nand ginst9053 (P1_U5967, P1_U4033, P1_U4621);
  nand ginst9054 (P1_U5968, P1_REG0_REG_23__SCAN_IN, P1_U3955);
  nand ginst9055 (P1_U5969, P1_U4033, P1_U4640);
  nand ginst9056 (P1_U5970, P1_REG0_REG_24__SCAN_IN, P1_U3955);
  nand ginst9057 (P1_U5971, P1_U4033, P1_U4659);
  nand ginst9058 (P1_U5972, P1_REG0_REG_25__SCAN_IN, P1_U3955);
  nand ginst9059 (P1_U5973, P1_U4033, P1_U4678);
  nand ginst9060 (P1_U5974, P1_REG0_REG_26__SCAN_IN, P1_U3955);
  nand ginst9061 (P1_U5975, P1_U4033, P1_U4697);
  nand ginst9062 (P1_U5976, P1_REG0_REG_27__SCAN_IN, P1_U3955);
  nand ginst9063 (P1_U5977, P1_U4033, P1_U4716);
  nand ginst9064 (P1_U5978, P1_REG0_REG_28__SCAN_IN, P1_U3955);
  nand ginst9065 (P1_U5979, P1_U4033, P1_U4735);
  nand ginst9066 (P1_U5980, P1_REG0_REG_29__SCAN_IN, P1_U3955);
  nand ginst9067 (P1_U5981, P1_U4033, P1_U4755);
  nand ginst9068 (P1_U5982, P1_REG0_REG_30__SCAN_IN, P1_U3955);
  nand ginst9069 (P1_U5983, P1_U4033, P1_U4762);
  nand ginst9070 (P1_U5984, P1_REG0_REG_31__SCAN_IN, P1_U3955);
  nand ginst9071 (P1_U5985, P1_U4033, P1_U4765);
  nand ginst9072 (P1_U5986, P1_REG1_REG_0__SCAN_IN, P1_U3956);
  nand ginst9073 (P1_U5987, P1_U4032, P1_U4198);
  nand ginst9074 (P1_U5988, P1_REG1_REG_1__SCAN_IN, P1_U3956);
  nand ginst9075 (P1_U5989, P1_U4032, P1_U4222);
  nand ginst9076 (P1_U5990, P1_REG1_REG_2__SCAN_IN, P1_U3956);
  nand ginst9077 (P1_U5991, P1_U4032, P1_U4241);
  nand ginst9078 (P1_U5992, P1_REG1_REG_3__SCAN_IN, P1_U3956);
  nand ginst9079 (P1_U5993, P1_U4032, P1_U4260);
  nand ginst9080 (P1_U5994, P1_REG1_REG_4__SCAN_IN, P1_U3956);
  nand ginst9081 (P1_U5995, P1_U4032, P1_U4279);
  nand ginst9082 (P1_U5996, P1_REG1_REG_5__SCAN_IN, P1_U3956);
  nand ginst9083 (P1_U5997, P1_U4032, P1_U4298);
  nand ginst9084 (P1_U5998, P1_REG1_REG_6__SCAN_IN, P1_U3956);
  nand ginst9085 (P1_U5999, P1_U4032, P1_U4317);
  nand ginst9086 (P1_U6000, P1_REG1_REG_7__SCAN_IN, P1_U3956);
  nand ginst9087 (P1_U6001, P1_U4032, P1_U4336);
  nand ginst9088 (P1_U6002, P1_REG1_REG_8__SCAN_IN, P1_U3956);
  nand ginst9089 (P1_U6003, P1_U4032, P1_U4355);
  nand ginst9090 (P1_U6004, P1_REG1_REG_9__SCAN_IN, P1_U3956);
  nand ginst9091 (P1_U6005, P1_U4032, P1_U4374);
  nand ginst9092 (P1_U6006, P1_REG1_REG_10__SCAN_IN, P1_U3956);
  nand ginst9093 (P1_U6007, P1_U4032, P1_U4393);
  nand ginst9094 (P1_U6008, P1_REG1_REG_11__SCAN_IN, P1_U3956);
  nand ginst9095 (P1_U6009, P1_U4032, P1_U4412);
  nand ginst9096 (P1_U6010, P1_REG1_REG_12__SCAN_IN, P1_U3956);
  nand ginst9097 (P1_U6011, P1_U4032, P1_U4431);
  nand ginst9098 (P1_U6012, P1_REG1_REG_13__SCAN_IN, P1_U3956);
  nand ginst9099 (P1_U6013, P1_U4032, P1_U4450);
  nand ginst9100 (P1_U6014, P1_REG1_REG_14__SCAN_IN, P1_U3956);
  nand ginst9101 (P1_U6015, P1_U4032, P1_U4469);
  nand ginst9102 (P1_U6016, P1_REG1_REG_15__SCAN_IN, P1_U3956);
  nand ginst9103 (P1_U6017, P1_U4032, P1_U4488);
  nand ginst9104 (P1_U6018, P1_REG1_REG_16__SCAN_IN, P1_U3956);
  nand ginst9105 (P1_U6019, P1_U4032, P1_U4507);
  nand ginst9106 (P1_U6020, P1_REG1_REG_17__SCAN_IN, P1_U3956);
  nand ginst9107 (P1_U6021, P1_U4032, P1_U4526);
  nand ginst9108 (P1_U6022, P1_REG1_REG_18__SCAN_IN, P1_U3956);
  nand ginst9109 (P1_U6023, P1_U4032, P1_U4545);
  nand ginst9110 (P1_U6024, P1_REG1_REG_19__SCAN_IN, P1_U3956);
  nand ginst9111 (P1_U6025, P1_U4032, P1_U4564);
  nand ginst9112 (P1_U6026, P1_REG1_REG_20__SCAN_IN, P1_U3956);
  nand ginst9113 (P1_U6027, P1_U4032, P1_U4583);
  nand ginst9114 (P1_U6028, P1_REG1_REG_21__SCAN_IN, P1_U3956);
  nand ginst9115 (P1_U6029, P1_U4032, P1_U4602);
  nand ginst9116 (P1_U6030, P1_REG1_REG_22__SCAN_IN, P1_U3956);
  nand ginst9117 (P1_U6031, P1_U4032, P1_U4621);
  nand ginst9118 (P1_U6032, P1_REG1_REG_23__SCAN_IN, P1_U3956);
  nand ginst9119 (P1_U6033, P1_U4032, P1_U4640);
  nand ginst9120 (P1_U6034, P1_REG1_REG_24__SCAN_IN, P1_U3956);
  nand ginst9121 (P1_U6035, P1_U4032, P1_U4659);
  nand ginst9122 (P1_U6036, P1_REG1_REG_25__SCAN_IN, P1_U3956);
  nand ginst9123 (P1_U6037, P1_U4032, P1_U4678);
  nand ginst9124 (P1_U6038, P1_REG1_REG_26__SCAN_IN, P1_U3956);
  nand ginst9125 (P1_U6039, P1_U4032, P1_U4697);
  nand ginst9126 (P1_U6040, P1_REG1_REG_27__SCAN_IN, P1_U3956);
  nand ginst9127 (P1_U6041, P1_U4032, P1_U4716);
  nand ginst9128 (P1_U6042, P1_REG1_REG_28__SCAN_IN, P1_U3956);
  nand ginst9129 (P1_U6043, P1_U4032, P1_U4735);
  nand ginst9130 (P1_U6044, P1_REG1_REG_29__SCAN_IN, P1_U3956);
  nand ginst9131 (P1_U6045, P1_U4032, P1_U4755);
  nand ginst9132 (P1_U6046, P1_REG1_REG_30__SCAN_IN, P1_U3956);
  nand ginst9133 (P1_U6047, P1_U4032, P1_U4762);
  nand ginst9134 (P1_U6048, P1_REG1_REG_31__SCAN_IN, P1_U3956);
  nand ginst9135 (P1_U6049, P1_U4032, P1_U4765);
  nand ginst9136 (P1_U6050, P1_REG2_REG_0__SCAN_IN, P1_U3420);
  nand ginst9137 (P1_U6051, P1_U3376, P1_U4031);
  nand ginst9138 (P1_U6052, P1_REG2_REG_1__SCAN_IN, P1_U3420);
  nand ginst9139 (P1_U6053, P1_U3378, P1_U4031);
  nand ginst9140 (P1_U6054, P1_REG2_REG_2__SCAN_IN, P1_U3420);
  nand ginst9141 (P1_U6055, P1_U3379, P1_U4031);
  nand ginst9142 (P1_U6056, P1_REG2_REG_3__SCAN_IN, P1_U3420);
  nand ginst9143 (P1_U6057, P1_U3380, P1_U4031);
  nand ginst9144 (P1_U6058, P1_REG2_REG_4__SCAN_IN, P1_U3420);
  nand ginst9145 (P1_U6059, P1_U3381, P1_U4031);
  nand ginst9146 (P1_U6060, P1_REG2_REG_5__SCAN_IN, P1_U3420);
  nand ginst9147 (P1_U6061, P1_U3382, P1_U4031);
  nand ginst9148 (P1_U6062, P1_REG2_REG_6__SCAN_IN, P1_U3420);
  nand ginst9149 (P1_U6063, P1_U3383, P1_U4031);
  nand ginst9150 (P1_U6064, P1_REG2_REG_7__SCAN_IN, P1_U3420);
  nand ginst9151 (P1_U6065, P1_U3384, P1_U4031);
  nand ginst9152 (P1_U6066, P1_REG2_REG_8__SCAN_IN, P1_U3420);
  nand ginst9153 (P1_U6067, P1_U3385, P1_U4031);
  nand ginst9154 (P1_U6068, P1_REG2_REG_9__SCAN_IN, P1_U3420);
  nand ginst9155 (P1_U6069, P1_U3386, P1_U4031);
  nand ginst9156 (P1_U6070, P1_REG2_REG_10__SCAN_IN, P1_U3420);
  nand ginst9157 (P1_U6071, P1_U3387, P1_U4031);
  nand ginst9158 (P1_U6072, P1_REG2_REG_11__SCAN_IN, P1_U3420);
  nand ginst9159 (P1_U6073, P1_U3388, P1_U4031);
  nand ginst9160 (P1_U6074, P1_REG2_REG_12__SCAN_IN, P1_U3420);
  nand ginst9161 (P1_U6075, P1_U3389, P1_U4031);
  nand ginst9162 (P1_U6076, P1_REG2_REG_13__SCAN_IN, P1_U3420);
  nand ginst9163 (P1_U6077, P1_U3390, P1_U4031);
  nand ginst9164 (P1_U6078, P1_REG2_REG_14__SCAN_IN, P1_U3420);
  nand ginst9165 (P1_U6079, P1_U3391, P1_U4031);
  nand ginst9166 (P1_U6080, P1_REG2_REG_15__SCAN_IN, P1_U3420);
  nand ginst9167 (P1_U6081, P1_U3392, P1_U4031);
  nand ginst9168 (P1_U6082, P1_REG2_REG_16__SCAN_IN, P1_U3420);
  nand ginst9169 (P1_U6083, P1_U3393, P1_U4031);
  nand ginst9170 (P1_U6084, P1_REG2_REG_17__SCAN_IN, P1_U3420);
  nand ginst9171 (P1_U6085, P1_U3394, P1_U4031);
  nand ginst9172 (P1_U6086, P1_REG2_REG_18__SCAN_IN, P1_U3420);
  nand ginst9173 (P1_U6087, P1_U3395, P1_U4031);
  nand ginst9174 (P1_U6088, P1_REG2_REG_19__SCAN_IN, P1_U3420);
  nand ginst9175 (P1_U6089, P1_U3396, P1_U4031);
  nand ginst9176 (P1_U6090, P1_REG2_REG_20__SCAN_IN, P1_U3420);
  nand ginst9177 (P1_U6091, P1_U3398, P1_U4031);
  nand ginst9178 (P1_U6092, P1_REG2_REG_21__SCAN_IN, P1_U3420);
  nand ginst9179 (P1_U6093, P1_U3400, P1_U4031);
  nand ginst9180 (P1_U6094, P1_REG2_REG_22__SCAN_IN, P1_U3420);
  nand ginst9181 (P1_U6095, P1_U3402, P1_U4031);
  nand ginst9182 (P1_U6096, P1_REG2_REG_23__SCAN_IN, P1_U3420);
  nand ginst9183 (P1_U6097, P1_U3404, P1_U4031);
  nand ginst9184 (P1_U6098, P1_REG2_REG_24__SCAN_IN, P1_U3420);
  nand ginst9185 (P1_U6099, P1_U3406, P1_U4031);
  nand ginst9186 (P1_U6100, P1_REG2_REG_25__SCAN_IN, P1_U3420);
  nand ginst9187 (P1_U6101, P1_U3408, P1_U4031);
  nand ginst9188 (P1_U6102, P1_REG2_REG_26__SCAN_IN, P1_U3420);
  nand ginst9189 (P1_U6103, P1_U3410, P1_U4031);
  nand ginst9190 (P1_U6104, P1_REG2_REG_27__SCAN_IN, P1_U3420);
  nand ginst9191 (P1_U6105, P1_U3412, P1_U4031);
  nand ginst9192 (P1_U6106, P1_REG2_REG_28__SCAN_IN, P1_U3420);
  nand ginst9193 (P1_U6107, P1_U3414, P1_U4031);
  nand ginst9194 (P1_U6108, P1_REG2_REG_29__SCAN_IN, P1_U3420);
  nand ginst9195 (P1_U6109, P1_U3416, P1_U4031);
  nand ginst9196 (P1_U6110, P1_REG2_REG_30__SCAN_IN, P1_U3420);
  nand ginst9197 (P1_U6111, P1_U4031, P1_U4035);
  nand ginst9198 (P1_U6112, P1_REG2_REG_31__SCAN_IN, P1_U3420);
  nand ginst9199 (P1_U6113, P1_U4031, P1_U4035);
  nand ginst9200 (P1_U6114, P1_DATAO_REG_0__SCAN_IN, P1_U3430);
  nand ginst9201 (P1_U6115, P1_U3077, P1_U4016);
  nand ginst9202 (P1_U6116, P1_DATAO_REG_1__SCAN_IN, P1_U3430);
  nand ginst9203 (P1_U6117, P1_U3078, P1_U4016);
  nand ginst9204 (P1_U6118, P1_DATAO_REG_2__SCAN_IN, P1_U3430);
  nand ginst9205 (P1_U6119, P1_U3068, P1_U4016);
  nand ginst9206 (P1_U6120, P1_DATAO_REG_3__SCAN_IN, P1_U3430);
  nand ginst9207 (P1_U6121, P1_U3064, P1_U4016);
  nand ginst9208 (P1_U6122, P1_DATAO_REG_4__SCAN_IN, P1_U3430);
  nand ginst9209 (P1_U6123, P1_U3060, P1_U4016);
  nand ginst9210 (P1_U6124, P1_DATAO_REG_5__SCAN_IN, P1_U3430);
  nand ginst9211 (P1_U6125, P1_U3067, P1_U4016);
  nand ginst9212 (P1_U6126, P1_DATAO_REG_6__SCAN_IN, P1_U3430);
  nand ginst9213 (P1_U6127, P1_U3071, P1_U4016);
  nand ginst9214 (P1_U6128, P1_DATAO_REG_7__SCAN_IN, P1_U3430);
  nand ginst9215 (P1_U6129, P1_U3070, P1_U4016);
  nand ginst9216 (P1_U6130, P1_DATAO_REG_8__SCAN_IN, P1_U3430);
  nand ginst9217 (P1_U6131, P1_U3084, P1_U4016);
  nand ginst9218 (P1_U6132, P1_DATAO_REG_9__SCAN_IN, P1_U3430);
  nand ginst9219 (P1_U6133, P1_U3083, P1_U4016);
  nand ginst9220 (P1_U6134, P1_DATAO_REG_10__SCAN_IN, P1_U3430);
  nand ginst9221 (P1_U6135, P1_U3062, P1_U4016);
  nand ginst9222 (P1_U6136, P1_DATAO_REG_11__SCAN_IN, P1_U3430);
  nand ginst9223 (P1_U6137, P1_U3063, P1_U4016);
  nand ginst9224 (P1_U6138, P1_DATAO_REG_12__SCAN_IN, P1_U3430);
  nand ginst9225 (P1_U6139, P1_U3072, P1_U4016);
  nand ginst9226 (P1_U6140, P1_DATAO_REG_13__SCAN_IN, P1_U3430);
  nand ginst9227 (P1_U6141, P1_U3080, P1_U4016);
  nand ginst9228 (P1_U6142, P1_DATAO_REG_14__SCAN_IN, P1_U3430);
  nand ginst9229 (P1_U6143, P1_U3079, P1_U4016);
  nand ginst9230 (P1_U6144, P1_DATAO_REG_15__SCAN_IN, P1_U3430);
  nand ginst9231 (P1_U6145, P1_U3074, P1_U4016);
  nand ginst9232 (P1_U6146, P1_DATAO_REG_16__SCAN_IN, P1_U3430);
  nand ginst9233 (P1_U6147, P1_U3073, P1_U4016);
  nand ginst9234 (P1_U6148, P1_DATAO_REG_17__SCAN_IN, P1_U3430);
  nand ginst9235 (P1_U6149, P1_U3069, P1_U4016);
  nand ginst9236 (P1_U6150, P1_DATAO_REG_18__SCAN_IN, P1_U3430);
  nand ginst9237 (P1_U6151, P1_U3082, P1_U4016);
  nand ginst9238 (P1_U6152, P1_DATAO_REG_19__SCAN_IN, P1_U3430);
  nand ginst9239 (P1_U6153, P1_U3081, P1_U4016);
  nand ginst9240 (P1_U6154, P1_DATAO_REG_20__SCAN_IN, P1_U3430);
  nand ginst9241 (P1_U6155, P1_U3076, P1_U4016);
  nand ginst9242 (P1_U6156, P1_DATAO_REG_21__SCAN_IN, P1_U3430);
  nand ginst9243 (P1_U6157, P1_U3075, P1_U4016);
  nand ginst9244 (P1_U6158, P1_DATAO_REG_22__SCAN_IN, P1_U3430);
  nand ginst9245 (P1_U6159, P1_U3061, P1_U4016);
  nand ginst9246 (P1_U6160, P1_DATAO_REG_23__SCAN_IN, P1_U3430);
  nand ginst9247 (P1_U6161, P1_U3066, P1_U4016);
  nand ginst9248 (P1_U6162, P1_DATAO_REG_24__SCAN_IN, P1_U3430);
  nand ginst9249 (P1_U6163, P1_U3065, P1_U4016);
  nand ginst9250 (P1_U6164, P1_DATAO_REG_25__SCAN_IN, P1_U3430);
  nand ginst9251 (P1_U6165, P1_U3058, P1_U4016);
  nand ginst9252 (P1_U6166, P1_DATAO_REG_26__SCAN_IN, P1_U3430);
  nand ginst9253 (P1_U6167, P1_U3057, P1_U4016);
  nand ginst9254 (P1_U6168, P1_DATAO_REG_27__SCAN_IN, P1_U3430);
  nand ginst9255 (P1_U6169, P1_U3053, P1_U4016);
  nand ginst9256 (P1_U6170, P1_DATAO_REG_28__SCAN_IN, P1_U3430);
  nand ginst9257 (P1_U6171, P1_U3054, P1_U4016);
  nand ginst9258 (P1_U6172, P1_DATAO_REG_29__SCAN_IN, P1_U3430);
  nand ginst9259 (P1_U6173, P1_U3055, P1_U4016);
  nand ginst9260 (P1_U6174, P1_DATAO_REG_30__SCAN_IN, P1_U3430);
  nand ginst9261 (P1_U6175, P1_U3059, P1_U4016);
  nand ginst9262 (P1_U6176, P1_DATAO_REG_31__SCAN_IN, P1_U3430);
  nand ginst9263 (P1_U6177, P1_U3056, P1_U4016);
  nand ginst9264 (P1_U6178, P1_U3432, P1_U3450, P1_U5793);
  nand ginst9265 (P1_U6179, P1_R1375_U9, P1_U4030);
  nand ginst9266 (P1_U6180, P1_U3054, P1_U4017);
  nand ginst9267 (P1_U6181, P1_U3413, P1_U4702);
  nand ginst9268 (P1_U6182, P1_U6180, P1_U6181);
  nand ginst9269 (P1_U6183, P1_U3056, P1_U4026);
  nand ginst9270 (P1_U6184, P1_U3418, P1_U4759);
  nand ginst9271 (P1_U6185, P1_U6183, P1_U6184);
  nand ginst9272 (P1_U6186, P1_U3076, P1_U4025);
  nand ginst9273 (P1_U6187, P1_U3397, P1_U4550);
  nand ginst9274 (P1_U6188, P1_U6186, P1_U6187);
  nand ginst9275 (P1_U6189, P1_U3059, P1_U4027);
  nand ginst9276 (P1_U6190, P1_U3417, P1_U4739);
  nand ginst9277 (P1_U6191, P1_U6189, P1_U6190);
  nand ginst9278 (P1_U6192, P1_U4531, P1_U5959);
  nand ginst9279 (P1_U6193, P1_U3081, P1_U3514);
  nand ginst9280 (P1_U6194, P1_U6192, P1_U6193);
  nand ginst9281 (P1_U6195, P1_U4379, P1_U5905);
  nand ginst9282 (P1_U6196, P1_U3063, P1_U3491);
  nand ginst9283 (P1_U6197, P1_U6195, P1_U6196);
  nand ginst9284 (P1_U6198, P1_U4246, P1_U5856);
  nand ginst9285 (P1_U6199, P1_U3060, P1_U3470);
  nand ginst9286 (P1_U6200, P1_U6198, P1_U6199);
  nand ginst9287 (P1_U6201, P1_U4360, P1_U5898);
  nand ginst9288 (P1_U6202, P1_U3062, P1_U3488);
  nand ginst9289 (P1_U6203, P1_U6201, P1_U6202);
  nand ginst9290 (P1_U6204, P1_U3055, P1_U4028);
  nand ginst9291 (P1_U6205, P1_U3415, P1_U4721);
  nand ginst9292 (P1_U6206, P1_U6204, P1_U6205);
  nand ginst9293 (P1_U6207, P1_U3053, P1_U4018);
  nand ginst9294 (P1_U6208, P1_U3411, P1_U4683);
  nand ginst9295 (P1_U6209, P1_U6207, P1_U6208);
  nand ginst9296 (P1_U6210, P1_U4493, P1_U5947);
  nand ginst9297 (P1_U6211, P1_U3069, P1_U3509);
  nand ginst9298 (P1_U6212, P1_U6210, P1_U6211);
  nand ginst9299 (P1_U6213, P1_U4322, P1_U5884);
  nand ginst9300 (P1_U6214, P1_U3084, P1_U3482);
  nand ginst9301 (P1_U6215, P1_U6213, P1_U6214);
  nand ginst9302 (P1_U6216, P1_U4341, P1_U5891);
  nand ginst9303 (P1_U6217, P1_U3083, P1_U3485);
  nand ginst9304 (P1_U6218, P1_U6216, P1_U6217);
  nand ginst9305 (P1_U6219, P1_U4417, P1_U5919);
  nand ginst9306 (P1_U6220, P1_U3080, P1_U3497);
  nand ginst9307 (P1_U6221, P1_U6219, P1_U6220);
  nand ginst9308 (P1_U6222, P1_U4436, P1_U5926);
  nand ginst9309 (P1_U6223, P1_U3079, P1_U3500);
  nand ginst9310 (P1_U6224, P1_U6222, P1_U6223);
  nand ginst9311 (P1_U6225, P1_U4208, P1_U5820);
  nand ginst9312 (P1_U6226, P1_U3077, P1_U3456);
  nand ginst9313 (P1_U6227, P1_U6225, P1_U6226);
  nand ginst9314 (P1_U6228, P1_U4184, P1_U5835);
  nand ginst9315 (P1_U6229, P1_U3078, P1_U3461);
  nand ginst9316 (P1_U6230, P1_U6228, P1_U6229);
  nand ginst9317 (P1_U6231, P1_U4455, P1_U5933);
  nand ginst9318 (P1_U6232, P1_U3074, P1_U3503);
  nand ginst9319 (P1_U6233, P1_U6231, P1_U6232);
  nand ginst9320 (P1_U6234, P1_U4474, P1_U5940);
  nand ginst9321 (P1_U6235, P1_U3073, P1_U3506);
  nand ginst9322 (P1_U6236, P1_U6234, P1_U6235);
  nand ginst9323 (P1_U6237, P1_U4284, P1_U5870);
  nand ginst9324 (P1_U6238, P1_U3071, P1_U3476);
  nand ginst9325 (P1_U6239, P1_U6237, P1_U6238);
  nand ginst9326 (P1_U6240, P1_U4303, P1_U5877);
  nand ginst9327 (P1_U6241, P1_U3070, P1_U3479);
  nand ginst9328 (P1_U6242, P1_U6240, P1_U6241);
  nand ginst9329 (P1_U6243, P1_U4398, P1_U5912);
  nand ginst9330 (P1_U6244, P1_U3072, P1_U3494);
  nand ginst9331 (P1_U6245, P1_U6243, P1_U6244);
  nand ginst9332 (P1_U6246, P1_U4203, P1_U5842);
  nand ginst9333 (P1_U6247, P1_U3068, P1_U3464);
  nand ginst9334 (P1_U6248, P1_U6246, P1_U6247);
  nand ginst9335 (P1_U6249, P1_U4227, P1_U5849);
  nand ginst9336 (P1_U6250, P1_U3064, P1_U3467);
  nand ginst9337 (P1_U6251, P1_U6249, P1_U6250);
  nand ginst9338 (P1_U6252, P1_U4265, P1_U5863);
  nand ginst9339 (P1_U6253, P1_U3067, P1_U3473);
  nand ginst9340 (P1_U6254, P1_U6252, P1_U6253);
  nand ginst9341 (P1_U6255, P1_U4512, P1_U5954);
  nand ginst9342 (P1_U6256, P1_U3082, P1_U3512);
  nand ginst9343 (P1_U6257, P1_U6255, P1_U6256);
  nand ginst9344 (P1_U6258, P1_U3065, P1_U4021);
  nand ginst9345 (P1_U6259, P1_U3405, P1_U4626);
  nand ginst9346 (P1_U6260, P1_U6258, P1_U6259);
  nand ginst9347 (P1_U6261, P1_U3066, P1_U4022);
  nand ginst9348 (P1_U6262, P1_U3403, P1_U4607);
  nand ginst9349 (P1_U6263, P1_U6261, P1_U6262);
  nand ginst9350 (P1_U6264, P1_U3075, P1_U4024);
  nand ginst9351 (P1_U6265, P1_U3399, P1_U4569);
  nand ginst9352 (P1_U6266, P1_U6264, P1_U6265);
  nand ginst9353 (P1_U6267, P1_U3061, P1_U4023);
  nand ginst9354 (P1_U6268, P1_U3401, P1_U4588);
  nand ginst9355 (P1_U6269, P1_U6267, P1_U6268);
  nand ginst9356 (P1_U6270, P1_U3058, P1_U4020);
  nand ginst9357 (P1_U6271, P1_U3407, P1_U4645);
  nand ginst9358 (P1_U6272, P1_U6270, P1_U6271);
  nand ginst9359 (P1_U6273, P1_U3057, P1_U4019);
  nand ginst9360 (P1_U6274, P1_U3409, P1_U4664);
  nand ginst9361 (P1_U6275, P1_U6273, P1_U6274);
  nand ginst9362 (P1_U6276, P1_U3991, P1_U4041);
  nand ginst9363 (P1_U6277, P1_U3049, P1_U5129);
  nand ginst9364 (P1_U6278, P1_U3432, P1_U5133, P1_U5799);
  nand ginst9365 (P1_U6279, P1_U3453, P1_U5130);
  nand ginst9366 (P1_U6280, P1_U3431, P1_U5786);
  nand ginst9367 (P1_U6281, P1_U3444, P1_U3451);
  nand ginst9368 (P1_U6282, P1_U3450, P1_U5144);
  nand ginst9369 (P1_U6283, P1_U3994, P1_U5802);
  nand ginst9370 (P1_U6284, P1_U3454, P1_U5408);
  nand ginst9371 (P1_U6285, P1_REG2_REG_0__SCAN_IN, P1_U3015, P1_U5814);
  not ginst9372 (P2_ADD_1119_U10, P2_REG3_REG_6__SCAN_IN);
  not ginst9373 (P2_ADD_1119_U100, P2_ADD_1119_U35);
  not ginst9374 (P2_ADD_1119_U101, P2_ADD_1119_U37);
  not ginst9375 (P2_ADD_1119_U102, P2_ADD_1119_U39);
  not ginst9376 (P2_ADD_1119_U103, P2_ADD_1119_U41);
  not ginst9377 (P2_ADD_1119_U104, P2_ADD_1119_U43);
  not ginst9378 (P2_ADD_1119_U105, P2_ADD_1119_U45);
  not ginst9379 (P2_ADD_1119_U106, P2_ADD_1119_U47);
  not ginst9380 (P2_ADD_1119_U107, P2_ADD_1119_U82);
  nand ginst9381 (P2_ADD_1119_U108, P2_REG3_REG_9__SCAN_IN, P2_ADD_1119_U79);
  nand ginst9382 (P2_ADD_1119_U109, P2_ADD_1119_U13, P2_ADD_1119_U88);
  nand ginst9383 (P2_ADD_1119_U11, P2_ADD_1119_U75, P2_ADD_1119_U85);
  nand ginst9384 (P2_ADD_1119_U110, P2_REG3_REG_8__SCAN_IN, P2_ADD_1119_U11);
  nand ginst9385 (P2_ADD_1119_U111, P2_ADD_1119_U12, P2_ADD_1119_U87);
  nand ginst9386 (P2_ADD_1119_U112, P2_REG3_REG_7__SCAN_IN, P2_ADD_1119_U80);
  nand ginst9387 (P2_ADD_1119_U113, P2_ADD_1119_U86, P2_ADD_1119_U9);
  nand ginst9388 (P2_ADD_1119_U114, P2_REG3_REG_6__SCAN_IN, P2_ADD_1119_U8);
  nand ginst9389 (P2_ADD_1119_U115, P2_ADD_1119_U10, P2_ADD_1119_U85);
  nand ginst9390 (P2_ADD_1119_U116, P2_REG3_REG_5__SCAN_IN, P2_ADD_1119_U81);
  nand ginst9391 (P2_ADD_1119_U117, P2_ADD_1119_U6, P2_ADD_1119_U84);
  nand ginst9392 (P2_ADD_1119_U118, P2_REG3_REG_4__SCAN_IN, P2_ADD_1119_U4);
  nand ginst9393 (P2_ADD_1119_U119, P2_REG3_REG_3__SCAN_IN, P2_ADD_1119_U7);
  not ginst9394 (P2_ADD_1119_U12, P2_REG3_REG_8__SCAN_IN);
  nand ginst9395 (P2_ADD_1119_U120, P2_REG3_REG_28__SCAN_IN, P2_ADD_1119_U82);
  nand ginst9396 (P2_ADD_1119_U121, P2_ADD_1119_U107, P2_ADD_1119_U48);
  nand ginst9397 (P2_ADD_1119_U122, P2_REG3_REG_27__SCAN_IN, P2_ADD_1119_U47);
  nand ginst9398 (P2_ADD_1119_U123, P2_ADD_1119_U106, P2_ADD_1119_U49);
  nand ginst9399 (P2_ADD_1119_U124, P2_REG3_REG_26__SCAN_IN, P2_ADD_1119_U45);
  nand ginst9400 (P2_ADD_1119_U125, P2_ADD_1119_U105, P2_ADD_1119_U46);
  nand ginst9401 (P2_ADD_1119_U126, P2_REG3_REG_25__SCAN_IN, P2_ADD_1119_U43);
  nand ginst9402 (P2_ADD_1119_U127, P2_ADD_1119_U104, P2_ADD_1119_U44);
  nand ginst9403 (P2_ADD_1119_U128, P2_REG3_REG_24__SCAN_IN, P2_ADD_1119_U41);
  nand ginst9404 (P2_ADD_1119_U129, P2_ADD_1119_U103, P2_ADD_1119_U42);
  not ginst9405 (P2_ADD_1119_U13, P2_REG3_REG_9__SCAN_IN);
  nand ginst9406 (P2_ADD_1119_U130, P2_REG3_REG_23__SCAN_IN, P2_ADD_1119_U39);
  nand ginst9407 (P2_ADD_1119_U131, P2_ADD_1119_U102, P2_ADD_1119_U40);
  nand ginst9408 (P2_ADD_1119_U132, P2_REG3_REG_22__SCAN_IN, P2_ADD_1119_U37);
  nand ginst9409 (P2_ADD_1119_U133, P2_ADD_1119_U101, P2_ADD_1119_U38);
  nand ginst9410 (P2_ADD_1119_U134, P2_REG3_REG_21__SCAN_IN, P2_ADD_1119_U35);
  nand ginst9411 (P2_ADD_1119_U135, P2_ADD_1119_U100, P2_ADD_1119_U36);
  nand ginst9412 (P2_ADD_1119_U136, P2_REG3_REG_20__SCAN_IN, P2_ADD_1119_U33);
  nand ginst9413 (P2_ADD_1119_U137, P2_ADD_1119_U34, P2_ADD_1119_U99);
  nand ginst9414 (P2_ADD_1119_U138, P2_REG3_REG_19__SCAN_IN, P2_ADD_1119_U31);
  nand ginst9415 (P2_ADD_1119_U139, P2_ADD_1119_U32, P2_ADD_1119_U98);
  nand ginst9416 (P2_ADD_1119_U14, P2_ADD_1119_U76, P2_ADD_1119_U87);
  nand ginst9417 (P2_ADD_1119_U140, P2_REG3_REG_18__SCAN_IN, P2_ADD_1119_U29);
  nand ginst9418 (P2_ADD_1119_U141, P2_ADD_1119_U30, P2_ADD_1119_U97);
  nand ginst9419 (P2_ADD_1119_U142, P2_REG3_REG_17__SCAN_IN, P2_ADD_1119_U27);
  nand ginst9420 (P2_ADD_1119_U143, P2_ADD_1119_U28, P2_ADD_1119_U96);
  nand ginst9421 (P2_ADD_1119_U144, P2_REG3_REG_16__SCAN_IN, P2_ADD_1119_U25);
  nand ginst9422 (P2_ADD_1119_U145, P2_ADD_1119_U26, P2_ADD_1119_U95);
  nand ginst9423 (P2_ADD_1119_U146, P2_REG3_REG_15__SCAN_IN, P2_ADD_1119_U23);
  nand ginst9424 (P2_ADD_1119_U147, P2_ADD_1119_U24, P2_ADD_1119_U94);
  nand ginst9425 (P2_ADD_1119_U148, P2_REG3_REG_14__SCAN_IN, P2_ADD_1119_U21);
  nand ginst9426 (P2_ADD_1119_U149, P2_ADD_1119_U22, P2_ADD_1119_U93);
  not ginst9427 (P2_ADD_1119_U15, P2_REG3_REG_11__SCAN_IN);
  nand ginst9428 (P2_ADD_1119_U150, P2_REG3_REG_13__SCAN_IN, P2_ADD_1119_U19);
  nand ginst9429 (P2_ADD_1119_U151, P2_ADD_1119_U20, P2_ADD_1119_U92);
  nand ginst9430 (P2_ADD_1119_U152, P2_REG3_REG_12__SCAN_IN, P2_ADD_1119_U17);
  nand ginst9431 (P2_ADD_1119_U153, P2_ADD_1119_U18, P2_ADD_1119_U91);
  nand ginst9432 (P2_ADD_1119_U154, P2_REG3_REG_11__SCAN_IN, P2_ADD_1119_U83);
  nand ginst9433 (P2_ADD_1119_U155, P2_ADD_1119_U15, P2_ADD_1119_U90);
  nand ginst9434 (P2_ADD_1119_U156, P2_REG3_REG_10__SCAN_IN, P2_ADD_1119_U14);
  nand ginst9435 (P2_ADD_1119_U157, P2_ADD_1119_U16, P2_ADD_1119_U89);
  not ginst9436 (P2_ADD_1119_U16, P2_REG3_REG_10__SCAN_IN);
  nand ginst9437 (P2_ADD_1119_U17, P2_ADD_1119_U77, P2_ADD_1119_U89);
  not ginst9438 (P2_ADD_1119_U18, P2_REG3_REG_12__SCAN_IN);
  nand ginst9439 (P2_ADD_1119_U19, P2_REG3_REG_12__SCAN_IN, P2_ADD_1119_U91);
  not ginst9440 (P2_ADD_1119_U20, P2_REG3_REG_13__SCAN_IN);
  nand ginst9441 (P2_ADD_1119_U21, P2_REG3_REG_13__SCAN_IN, P2_ADD_1119_U92);
  not ginst9442 (P2_ADD_1119_U22, P2_REG3_REG_14__SCAN_IN);
  nand ginst9443 (P2_ADD_1119_U23, P2_REG3_REG_14__SCAN_IN, P2_ADD_1119_U93);
  not ginst9444 (P2_ADD_1119_U24, P2_REG3_REG_15__SCAN_IN);
  nand ginst9445 (P2_ADD_1119_U25, P2_REG3_REG_15__SCAN_IN, P2_ADD_1119_U94);
  not ginst9446 (P2_ADD_1119_U26, P2_REG3_REG_16__SCAN_IN);
  nand ginst9447 (P2_ADD_1119_U27, P2_REG3_REG_16__SCAN_IN, P2_ADD_1119_U95);
  not ginst9448 (P2_ADD_1119_U28, P2_REG3_REG_17__SCAN_IN);
  nand ginst9449 (P2_ADD_1119_U29, P2_REG3_REG_17__SCAN_IN, P2_ADD_1119_U96);
  not ginst9450 (P2_ADD_1119_U30, P2_REG3_REG_18__SCAN_IN);
  nand ginst9451 (P2_ADD_1119_U31, P2_REG3_REG_18__SCAN_IN, P2_ADD_1119_U97);
  not ginst9452 (P2_ADD_1119_U32, P2_REG3_REG_19__SCAN_IN);
  nand ginst9453 (P2_ADD_1119_U33, P2_REG3_REG_19__SCAN_IN, P2_ADD_1119_U98);
  not ginst9454 (P2_ADD_1119_U34, P2_REG3_REG_20__SCAN_IN);
  nand ginst9455 (P2_ADD_1119_U35, P2_REG3_REG_20__SCAN_IN, P2_ADD_1119_U99);
  not ginst9456 (P2_ADD_1119_U36, P2_REG3_REG_21__SCAN_IN);
  nand ginst9457 (P2_ADD_1119_U37, P2_REG3_REG_21__SCAN_IN, P2_ADD_1119_U100);
  not ginst9458 (P2_ADD_1119_U38, P2_REG3_REG_22__SCAN_IN);
  nand ginst9459 (P2_ADD_1119_U39, P2_REG3_REG_22__SCAN_IN, P2_ADD_1119_U101);
  not ginst9460 (P2_ADD_1119_U4, P2_REG3_REG_3__SCAN_IN);
  not ginst9461 (P2_ADD_1119_U40, P2_REG3_REG_23__SCAN_IN);
  nand ginst9462 (P2_ADD_1119_U41, P2_REG3_REG_23__SCAN_IN, P2_ADD_1119_U102);
  not ginst9463 (P2_ADD_1119_U42, P2_REG3_REG_24__SCAN_IN);
  nand ginst9464 (P2_ADD_1119_U43, P2_REG3_REG_24__SCAN_IN, P2_ADD_1119_U103);
  not ginst9465 (P2_ADD_1119_U44, P2_REG3_REG_25__SCAN_IN);
  nand ginst9466 (P2_ADD_1119_U45, P2_REG3_REG_25__SCAN_IN, P2_ADD_1119_U104);
  not ginst9467 (P2_ADD_1119_U46, P2_REG3_REG_26__SCAN_IN);
  nand ginst9468 (P2_ADD_1119_U47, P2_REG3_REG_26__SCAN_IN, P2_ADD_1119_U105);
  not ginst9469 (P2_ADD_1119_U48, P2_REG3_REG_28__SCAN_IN);
  not ginst9470 (P2_ADD_1119_U49, P2_REG3_REG_27__SCAN_IN);
  and ginst9471 (P2_ADD_1119_U5, P2_ADD_1119_U106, P2_ADD_1119_U78);
  nand ginst9472 (P2_ADD_1119_U50, P2_ADD_1119_U108, P2_ADD_1119_U109);
  nand ginst9473 (P2_ADD_1119_U51, P2_ADD_1119_U110, P2_ADD_1119_U111);
  nand ginst9474 (P2_ADD_1119_U52, P2_ADD_1119_U112, P2_ADD_1119_U113);
  nand ginst9475 (P2_ADD_1119_U53, P2_ADD_1119_U114, P2_ADD_1119_U115);
  nand ginst9476 (P2_ADD_1119_U54, P2_ADD_1119_U116, P2_ADD_1119_U117);
  nand ginst9477 (P2_ADD_1119_U55, P2_ADD_1119_U118, P2_ADD_1119_U119);
  nand ginst9478 (P2_ADD_1119_U56, P2_ADD_1119_U120, P2_ADD_1119_U121);
  nand ginst9479 (P2_ADD_1119_U57, P2_ADD_1119_U122, P2_ADD_1119_U123);
  nand ginst9480 (P2_ADD_1119_U58, P2_ADD_1119_U124, P2_ADD_1119_U125);
  nand ginst9481 (P2_ADD_1119_U59, P2_ADD_1119_U126, P2_ADD_1119_U127);
  not ginst9482 (P2_ADD_1119_U6, P2_REG3_REG_5__SCAN_IN);
  nand ginst9483 (P2_ADD_1119_U60, P2_ADD_1119_U128, P2_ADD_1119_U129);
  nand ginst9484 (P2_ADD_1119_U61, P2_ADD_1119_U130, P2_ADD_1119_U131);
  nand ginst9485 (P2_ADD_1119_U62, P2_ADD_1119_U132, P2_ADD_1119_U133);
  nand ginst9486 (P2_ADD_1119_U63, P2_ADD_1119_U134, P2_ADD_1119_U135);
  nand ginst9487 (P2_ADD_1119_U64, P2_ADD_1119_U136, P2_ADD_1119_U137);
  nand ginst9488 (P2_ADD_1119_U65, P2_ADD_1119_U138, P2_ADD_1119_U139);
  nand ginst9489 (P2_ADD_1119_U66, P2_ADD_1119_U140, P2_ADD_1119_U141);
  nand ginst9490 (P2_ADD_1119_U67, P2_ADD_1119_U142, P2_ADD_1119_U143);
  nand ginst9491 (P2_ADD_1119_U68, P2_ADD_1119_U144, P2_ADD_1119_U145);
  nand ginst9492 (P2_ADD_1119_U69, P2_ADD_1119_U146, P2_ADD_1119_U147);
  not ginst9493 (P2_ADD_1119_U7, P2_REG3_REG_4__SCAN_IN);
  nand ginst9494 (P2_ADD_1119_U70, P2_ADD_1119_U148, P2_ADD_1119_U149);
  nand ginst9495 (P2_ADD_1119_U71, P2_ADD_1119_U150, P2_ADD_1119_U151);
  nand ginst9496 (P2_ADD_1119_U72, P2_ADD_1119_U152, P2_ADD_1119_U153);
  nand ginst9497 (P2_ADD_1119_U73, P2_ADD_1119_U154, P2_ADD_1119_U155);
  nand ginst9498 (P2_ADD_1119_U74, P2_ADD_1119_U156, P2_ADD_1119_U157);
  and ginst9499 (P2_ADD_1119_U75, P2_REG3_REG_6__SCAN_IN, P2_REG3_REG_7__SCAN_IN);
  and ginst9500 (P2_ADD_1119_U76, P2_REG3_REG_9__SCAN_IN, P2_REG3_REG_8__SCAN_IN);
  and ginst9501 (P2_ADD_1119_U77, P2_REG3_REG_11__SCAN_IN, P2_REG3_REG_10__SCAN_IN);
  and ginst9502 (P2_ADD_1119_U78, P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_27__SCAN_IN);
  nand ginst9503 (P2_ADD_1119_U79, P2_REG3_REG_8__SCAN_IN, P2_ADD_1119_U87);
  nand ginst9504 (P2_ADD_1119_U8, P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_5__SCAN_IN, P2_REG3_REG_3__SCAN_IN);
  nand ginst9505 (P2_ADD_1119_U80, P2_REG3_REG_6__SCAN_IN, P2_ADD_1119_U85);
  nand ginst9506 (P2_ADD_1119_U81, P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_3__SCAN_IN);
  nand ginst9507 (P2_ADD_1119_U82, P2_REG3_REG_27__SCAN_IN, P2_ADD_1119_U106);
  nand ginst9508 (P2_ADD_1119_U83, P2_REG3_REG_10__SCAN_IN, P2_ADD_1119_U89);
  not ginst9509 (P2_ADD_1119_U84, P2_ADD_1119_U81);
  not ginst9510 (P2_ADD_1119_U85, P2_ADD_1119_U8);
  not ginst9511 (P2_ADD_1119_U86, P2_ADD_1119_U80);
  not ginst9512 (P2_ADD_1119_U87, P2_ADD_1119_U11);
  not ginst9513 (P2_ADD_1119_U88, P2_ADD_1119_U79);
  not ginst9514 (P2_ADD_1119_U89, P2_ADD_1119_U14);
  not ginst9515 (P2_ADD_1119_U9, P2_REG3_REG_7__SCAN_IN);
  not ginst9516 (P2_ADD_1119_U90, P2_ADD_1119_U83);
  not ginst9517 (P2_ADD_1119_U91, P2_ADD_1119_U17);
  not ginst9518 (P2_ADD_1119_U92, P2_ADD_1119_U19);
  not ginst9519 (P2_ADD_1119_U93, P2_ADD_1119_U21);
  not ginst9520 (P2_ADD_1119_U94, P2_ADD_1119_U23);
  not ginst9521 (P2_ADD_1119_U95, P2_ADD_1119_U25);
  not ginst9522 (P2_ADD_1119_U96, P2_ADD_1119_U27);
  not ginst9523 (P2_ADD_1119_U97, P2_ADD_1119_U29);
  not ginst9524 (P2_ADD_1119_U98, P2_ADD_1119_U31);
  not ginst9525 (P2_ADD_1119_U99, P2_ADD_1119_U33);
  and ginst9526 (P2_R1113_U10, P2_R1113_U182, P2_R1113_U282);
  nand ginst9527 (P2_R1113_U100, P2_R1113_U449, P2_R1113_U450);
  nand ginst9528 (P2_R1113_U101, P2_R1113_U465, P2_R1113_U466);
  nand ginst9529 (P2_R1113_U102, P2_R1113_U470, P2_R1113_U471);
  nand ginst9530 (P2_R1113_U103, P2_R1113_U355, P2_R1113_U356);
  nand ginst9531 (P2_R1113_U104, P2_R1113_U364, P2_R1113_U365);
  nand ginst9532 (P2_R1113_U105, P2_R1113_U371, P2_R1113_U372);
  nand ginst9533 (P2_R1113_U106, P2_R1113_U375, P2_R1113_U376);
  nand ginst9534 (P2_R1113_U107, P2_R1113_U384, P2_R1113_U385);
  nand ginst9535 (P2_R1113_U108, P2_R1113_U403, P2_R1113_U404);
  nand ginst9536 (P2_R1113_U109, P2_R1113_U420, P2_R1113_U421);
  and ginst9537 (P2_R1113_U11, P2_R1113_U283, P2_R1113_U284);
  nand ginst9538 (P2_R1113_U110, P2_R1113_U424, P2_R1113_U425);
  nand ginst9539 (P2_R1113_U111, P2_R1113_U456, P2_R1113_U457);
  nand ginst9540 (P2_R1113_U112, P2_R1113_U460, P2_R1113_U461);
  nand ginst9541 (P2_R1113_U113, P2_R1113_U477, P2_R1113_U478);
  and ginst9542 (P2_R1113_U114, P2_R1113_U184, P2_R1113_U194);
  and ginst9543 (P2_R1113_U115, P2_R1113_U197, P2_R1113_U198);
  and ginst9544 (P2_R1113_U116, P2_R1113_U185, P2_R1113_U200, P2_R1113_U205);
  and ginst9545 (P2_R1113_U117, P2_R1113_U186, P2_R1113_U210);
  and ginst9546 (P2_R1113_U118, P2_R1113_U213, P2_R1113_U214);
  and ginst9547 (P2_R1113_U119, P2_R1113_U357, P2_R1113_U358, P2_R1113_U38);
  nand ginst9548 (P2_R1113_U12, P2_R1113_U344, P2_R1113_U347);
  and ginst9549 (P2_R1113_U120, P2_R1113_U186, P2_R1113_U361);
  and ginst9550 (P2_R1113_U121, P2_R1113_U229, P2_R1113_U6);
  and ginst9551 (P2_R1113_U122, P2_R1113_U185, P2_R1113_U368);
  and ginst9552 (P2_R1113_U123, P2_R1113_U28, P2_R1113_U377, P2_R1113_U378);
  and ginst9553 (P2_R1113_U124, P2_R1113_U184, P2_R1113_U381);
  and ginst9554 (P2_R1113_U125, P2_R1113_U180, P2_R1113_U216, P2_R1113_U239);
  and ginst9555 (P2_R1113_U126, P2_R1113_U261, P2_R1113_U8);
  and ginst9556 (P2_R1113_U127, P2_R1113_U10, P2_R1113_U287);
  and ginst9557 (P2_R1113_U128, P2_R1113_U303, P2_R1113_U304);
  and ginst9558 (P2_R1113_U129, P2_R1113_U311, P2_R1113_U386, P2_R1113_U387);
  nand ginst9559 (P2_R1113_U13, P2_R1113_U333, P2_R1113_U336);
  and ginst9560 (P2_R1113_U130, P2_R1113_U308, P2_R1113_U390);
  nand ginst9561 (P2_R1113_U131, P2_R1113_U391, P2_R1113_U392);
  and ginst9562 (P2_R1113_U132, P2_R1113_U396, P2_R1113_U397, P2_R1113_U83);
  and ginst9563 (P2_R1113_U133, P2_R1113_U183, P2_R1113_U400);
  nand ginst9564 (P2_R1113_U134, P2_R1113_U405, P2_R1113_U406);
  nand ginst9565 (P2_R1113_U135, P2_R1113_U410, P2_R1113_U411);
  and ginst9566 (P2_R1113_U136, P2_R1113_U11, P2_R1113_U324);
  and ginst9567 (P2_R1113_U137, P2_R1113_U182, P2_R1113_U417);
  nand ginst9568 (P2_R1113_U138, P2_R1113_U426, P2_R1113_U427);
  nand ginst9569 (P2_R1113_U139, P2_R1113_U431, P2_R1113_U432);
  nand ginst9570 (P2_R1113_U14, P2_R1113_U322, P2_R1113_U325);
  nand ginst9571 (P2_R1113_U140, P2_R1113_U436, P2_R1113_U437);
  nand ginst9572 (P2_R1113_U141, P2_R1113_U441, P2_R1113_U442);
  nand ginst9573 (P2_R1113_U142, P2_R1113_U446, P2_R1113_U447);
  and ginst9574 (P2_R1113_U143, P2_R1113_U335, P2_R1113_U9);
  and ginst9575 (P2_R1113_U144, P2_R1113_U181, P2_R1113_U453);
  nand ginst9576 (P2_R1113_U145, P2_R1113_U462, P2_R1113_U463);
  nand ginst9577 (P2_R1113_U146, P2_R1113_U467, P2_R1113_U468);
  and ginst9578 (P2_R1113_U147, P2_R1113_U346, P2_R1113_U7);
  and ginst9579 (P2_R1113_U148, P2_R1113_U180, P2_R1113_U474);
  and ginst9580 (P2_R1113_U149, P2_R1113_U353, P2_R1113_U354);
  nand ginst9581 (P2_R1113_U15, P2_R1113_U314, P2_R1113_U316);
  nand ginst9582 (P2_R1113_U150, P2_R1113_U118, P2_R1113_U211);
  and ginst9583 (P2_R1113_U151, P2_R1113_U362, P2_R1113_U363);
  and ginst9584 (P2_R1113_U152, P2_R1113_U369, P2_R1113_U370);
  and ginst9585 (P2_R1113_U153, P2_R1113_U373, P2_R1113_U374);
  nand ginst9586 (P2_R1113_U154, P2_R1113_U115, P2_R1113_U195);
  and ginst9587 (P2_R1113_U155, P2_R1113_U382, P2_R1113_U383);
  not ginst9588 (P2_R1113_U156, P2_U3960);
  not ginst9589 (P2_R1113_U157, P2_U3057);
  and ginst9590 (P2_R1113_U158, P2_R1113_U401, P2_R1113_U402);
  nand ginst9591 (P2_R1113_U159, P2_R1113_U293, P2_R1113_U294);
  nand ginst9592 (P2_R1113_U16, P2_R1113_U312, P2_R1113_U352);
  nand ginst9593 (P2_R1113_U160, P2_R1113_U289, P2_R1113_U290);
  and ginst9594 (P2_R1113_U161, P2_R1113_U418, P2_R1113_U419);
  and ginst9595 (P2_R1113_U162, P2_R1113_U422, P2_R1113_U423);
  nand ginst9596 (P2_R1113_U163, P2_R1113_U279, P2_R1113_U280);
  nand ginst9597 (P2_R1113_U164, P2_R1113_U275, P2_R1113_U276);
  not ginst9598 (P2_R1113_U165, P2_U3432);
  nand ginst9599 (P2_R1113_U166, P2_R1113_U92, P2_U3427);
  nand ginst9600 (P2_R1113_U167, P2_R1113_U271, P2_R1113_U272);
  not ginst9601 (P2_R1113_U168, P2_U3483);
  nand ginst9602 (P2_R1113_U169, P2_R1113_U263, P2_R1113_U264);
  nand ginst9603 (P2_R1113_U17, P2_R1113_U235, P2_R1113_U237);
  and ginst9604 (P2_R1113_U170, P2_R1113_U454, P2_R1113_U455);
  and ginst9605 (P2_R1113_U171, P2_R1113_U458, P2_R1113_U459);
  nand ginst9606 (P2_R1113_U172, P2_R1113_U253, P2_R1113_U254);
  nand ginst9607 (P2_R1113_U173, P2_R1113_U249, P2_R1113_U250);
  nand ginst9608 (P2_R1113_U174, P2_R1113_U245, P2_R1113_U246);
  and ginst9609 (P2_R1113_U175, P2_R1113_U475, P2_R1113_U476);
  nand ginst9610 (P2_R1113_U176, P2_R1113_U165, P2_R1113_U166);
  not ginst9611 (P2_R1113_U177, P2_R1113_U83);
  not ginst9612 (P2_R1113_U178, P2_R1113_U28);
  not ginst9613 (P2_R1113_U179, P2_R1113_U38);
  nand ginst9614 (P2_R1113_U18, P2_R1113_U227, P2_R1113_U230);
  nand ginst9615 (P2_R1113_U180, P2_R1113_U49, P2_U3459);
  nand ginst9616 (P2_R1113_U181, P2_R1113_U59, P2_U3474);
  nand ginst9617 (P2_R1113_U182, P2_R1113_U74, P2_U3955);
  nand ginst9618 (P2_R1113_U183, P2_R1113_U82, P2_U3951);
  nand ginst9619 (P2_R1113_U184, P2_R1113_U27, P2_U3435);
  nand ginst9620 (P2_R1113_U185, P2_R1113_U33, P2_U3444);
  nand ginst9621 (P2_R1113_U186, P2_R1113_U37, P2_U3450);
  not ginst9622 (P2_R1113_U187, P2_R1113_U61);
  not ginst9623 (P2_R1113_U188, P2_R1113_U76);
  not ginst9624 (P2_R1113_U189, P2_R1113_U35);
  nand ginst9625 (P2_R1113_U19, P2_R1113_U219, P2_R1113_U221);
  not ginst9626 (P2_R1113_U190, P2_R1113_U50);
  not ginst9627 (P2_R1113_U191, P2_R1113_U166);
  nand ginst9628 (P2_R1113_U192, P2_R1113_U166, P2_U3080);
  not ginst9629 (P2_R1113_U193, P2_R1113_U44);
  nand ginst9630 (P2_R1113_U194, P2_R1113_U29, P2_U3438);
  nand ginst9631 (P2_R1113_U195, P2_R1113_U114, P2_R1113_U44);
  nand ginst9632 (P2_R1113_U196, P2_R1113_U28, P2_R1113_U29);
  nand ginst9633 (P2_R1113_U197, P2_R1113_U196, P2_R1113_U26);
  nand ginst9634 (P2_R1113_U198, P2_R1113_U178, P2_U3066);
  not ginst9635 (P2_R1113_U199, P2_R1113_U154);
  nand ginst9636 (P2_R1113_U20, P2_R1113_U166, P2_R1113_U350);
  nand ginst9637 (P2_R1113_U200, P2_R1113_U32, P2_U3447);
  nand ginst9638 (P2_R1113_U201, P2_R1113_U30, P2_U3073);
  nand ginst9639 (P2_R1113_U202, P2_R1113_U22, P2_U3069);
  nand ginst9640 (P2_R1113_U203, P2_R1113_U185, P2_R1113_U189);
  nand ginst9641 (P2_R1113_U204, P2_R1113_U203, P2_R1113_U6);
  nand ginst9642 (P2_R1113_U205, P2_R1113_U34, P2_U3441);
  nand ginst9643 (P2_R1113_U206, P2_R1113_U32, P2_U3447);
  nand ginst9644 (P2_R1113_U207, P2_R1113_U116, P2_R1113_U154);
  nand ginst9645 (P2_R1113_U208, P2_R1113_U204, P2_R1113_U206);
  not ginst9646 (P2_R1113_U209, P2_R1113_U42);
  not ginst9647 (P2_R1113_U21, P2_U3450);
  nand ginst9648 (P2_R1113_U210, P2_R1113_U39, P2_U3453);
  nand ginst9649 (P2_R1113_U211, P2_R1113_U117, P2_R1113_U42);
  nand ginst9650 (P2_R1113_U212, P2_R1113_U38, P2_R1113_U39);
  nand ginst9651 (P2_R1113_U213, P2_R1113_U212, P2_R1113_U36);
  nand ginst9652 (P2_R1113_U214, P2_R1113_U179, P2_U3086);
  not ginst9653 (P2_R1113_U215, P2_R1113_U150);
  nand ginst9654 (P2_R1113_U216, P2_R1113_U41, P2_U3456);
  nand ginst9655 (P2_R1113_U217, P2_R1113_U216, P2_R1113_U50);
  nand ginst9656 (P2_R1113_U218, P2_R1113_U209, P2_R1113_U38);
  nand ginst9657 (P2_R1113_U219, P2_R1113_U120, P2_R1113_U218);
  not ginst9658 (P2_R1113_U22, P2_U3444);
  nand ginst9659 (P2_R1113_U220, P2_R1113_U186, P2_R1113_U42);
  nand ginst9660 (P2_R1113_U221, P2_R1113_U119, P2_R1113_U220);
  nand ginst9661 (P2_R1113_U222, P2_R1113_U186, P2_R1113_U38);
  nand ginst9662 (P2_R1113_U223, P2_R1113_U154, P2_R1113_U205);
  not ginst9663 (P2_R1113_U224, P2_R1113_U43);
  nand ginst9664 (P2_R1113_U225, P2_R1113_U22, P2_U3069);
  nand ginst9665 (P2_R1113_U226, P2_R1113_U224, P2_R1113_U225);
  nand ginst9666 (P2_R1113_U227, P2_R1113_U122, P2_R1113_U226);
  nand ginst9667 (P2_R1113_U228, P2_R1113_U185, P2_R1113_U43);
  nand ginst9668 (P2_R1113_U229, P2_R1113_U32, P2_U3447);
  not ginst9669 (P2_R1113_U23, P2_U3435);
  nand ginst9670 (P2_R1113_U230, P2_R1113_U121, P2_R1113_U228);
  nand ginst9671 (P2_R1113_U231, P2_R1113_U22, P2_U3069);
  nand ginst9672 (P2_R1113_U232, P2_R1113_U185, P2_R1113_U231);
  nand ginst9673 (P2_R1113_U233, P2_R1113_U205, P2_R1113_U35);
  nand ginst9674 (P2_R1113_U234, P2_R1113_U193, P2_R1113_U28);
  nand ginst9675 (P2_R1113_U235, P2_R1113_U124, P2_R1113_U234);
  nand ginst9676 (P2_R1113_U236, P2_R1113_U184, P2_R1113_U44);
  nand ginst9677 (P2_R1113_U237, P2_R1113_U123, P2_R1113_U236);
  nand ginst9678 (P2_R1113_U238, P2_R1113_U184, P2_R1113_U28);
  nand ginst9679 (P2_R1113_U239, P2_R1113_U48, P2_U3462);
  not ginst9680 (P2_R1113_U24, P2_U3427);
  nand ginst9681 (P2_R1113_U240, P2_R1113_U47, P2_U3065);
  nand ginst9682 (P2_R1113_U241, P2_R1113_U46, P2_U3064);
  nand ginst9683 (P2_R1113_U242, P2_R1113_U180, P2_R1113_U190);
  nand ginst9684 (P2_R1113_U243, P2_R1113_U242, P2_R1113_U7);
  nand ginst9685 (P2_R1113_U244, P2_R1113_U48, P2_U3462);
  nand ginst9686 (P2_R1113_U245, P2_R1113_U125, P2_R1113_U150);
  nand ginst9687 (P2_R1113_U246, P2_R1113_U243, P2_R1113_U244);
  not ginst9688 (P2_R1113_U247, P2_R1113_U174);
  nand ginst9689 (P2_R1113_U248, P2_R1113_U52, P2_U3465);
  nand ginst9690 (P2_R1113_U249, P2_R1113_U174, P2_R1113_U248);
  not ginst9691 (P2_R1113_U25, P2_U3080);
  nand ginst9692 (P2_R1113_U250, P2_R1113_U51, P2_U3074);
  not ginst9693 (P2_R1113_U251, P2_R1113_U173);
  nand ginst9694 (P2_R1113_U252, P2_R1113_U54, P2_U3468);
  nand ginst9695 (P2_R1113_U253, P2_R1113_U173, P2_R1113_U252);
  nand ginst9696 (P2_R1113_U254, P2_R1113_U53, P2_U3082);
  not ginst9697 (P2_R1113_U255, P2_R1113_U172);
  nand ginst9698 (P2_R1113_U256, P2_R1113_U58, P2_U3477);
  nand ginst9699 (P2_R1113_U257, P2_R1113_U55, P2_U3075);
  nand ginst9700 (P2_R1113_U258, P2_R1113_U56, P2_U3076);
  nand ginst9701 (P2_R1113_U259, P2_R1113_U187, P2_R1113_U8);
  not ginst9702 (P2_R1113_U26, P2_U3438);
  nand ginst9703 (P2_R1113_U260, P2_R1113_U259, P2_R1113_U9);
  nand ginst9704 (P2_R1113_U261, P2_R1113_U60, P2_U3471);
  nand ginst9705 (P2_R1113_U262, P2_R1113_U58, P2_U3477);
  nand ginst9706 (P2_R1113_U263, P2_R1113_U126, P2_R1113_U172);
  nand ginst9707 (P2_R1113_U264, P2_R1113_U260, P2_R1113_U262);
  not ginst9708 (P2_R1113_U265, P2_R1113_U169);
  nand ginst9709 (P2_R1113_U266, P2_R1113_U63, P2_U3480);
  nand ginst9710 (P2_R1113_U267, P2_R1113_U169, P2_R1113_U266);
  nand ginst9711 (P2_R1113_U268, P2_R1113_U62, P2_U3071);
  not ginst9712 (P2_R1113_U269, P2_R1113_U64);
  not ginst9713 (P2_R1113_U27, P2_U3070);
  nand ginst9714 (P2_R1113_U270, P2_R1113_U269, P2_R1113_U65);
  nand ginst9715 (P2_R1113_U271, P2_R1113_U168, P2_R1113_U270);
  nand ginst9716 (P2_R1113_U272, P2_R1113_U64, P2_U3084);
  not ginst9717 (P2_R1113_U273, P2_R1113_U167);
  nand ginst9718 (P2_R1113_U274, P2_R1113_U67, P2_U3485);
  nand ginst9719 (P2_R1113_U275, P2_R1113_U167, P2_R1113_U274);
  nand ginst9720 (P2_R1113_U276, P2_R1113_U66, P2_U3083);
  not ginst9721 (P2_R1113_U277, P2_R1113_U164);
  nand ginst9722 (P2_R1113_U278, P2_R1113_U69, P2_U3957);
  nand ginst9723 (P2_R1113_U279, P2_R1113_U164, P2_R1113_U278);
  nand ginst9724 (P2_R1113_U28, P2_R1113_U23, P2_U3070);
  nand ginst9725 (P2_R1113_U280, P2_R1113_U68, P2_U3078);
  not ginst9726 (P2_R1113_U281, P2_R1113_U163);
  nand ginst9727 (P2_R1113_U282, P2_R1113_U73, P2_U3954);
  nand ginst9728 (P2_R1113_U283, P2_R1113_U70, P2_U3068);
  nand ginst9729 (P2_R1113_U284, P2_R1113_U71, P2_U3063);
  nand ginst9730 (P2_R1113_U285, P2_R1113_U10, P2_R1113_U188);
  nand ginst9731 (P2_R1113_U286, P2_R1113_U11, P2_R1113_U285);
  nand ginst9732 (P2_R1113_U287, P2_R1113_U75, P2_U3956);
  nand ginst9733 (P2_R1113_U288, P2_R1113_U73, P2_U3954);
  nand ginst9734 (P2_R1113_U289, P2_R1113_U127, P2_R1113_U163);
  not ginst9735 (P2_R1113_U29, P2_U3066);
  nand ginst9736 (P2_R1113_U290, P2_R1113_U286, P2_R1113_U288);
  not ginst9737 (P2_R1113_U291, P2_R1113_U160);
  nand ginst9738 (P2_R1113_U292, P2_R1113_U78, P2_U3953);
  nand ginst9739 (P2_R1113_U293, P2_R1113_U160, P2_R1113_U292);
  nand ginst9740 (P2_R1113_U294, P2_R1113_U77, P2_U3067);
  not ginst9741 (P2_R1113_U295, P2_R1113_U159);
  nand ginst9742 (P2_R1113_U296, P2_R1113_U80, P2_U3952);
  nand ginst9743 (P2_R1113_U297, P2_R1113_U159, P2_R1113_U296);
  nand ginst9744 (P2_R1113_U298, P2_R1113_U79, P2_U3060);
  not ginst9745 (P2_R1113_U299, P2_R1113_U88);
  not ginst9746 (P2_R1113_U30, P2_U3447);
  nand ginst9747 (P2_R1113_U300, P2_R1113_U84, P2_U3950);
  nand ginst9748 (P2_R1113_U301, P2_R1113_U183, P2_R1113_U300, P2_R1113_U88);
  nand ginst9749 (P2_R1113_U302, P2_R1113_U83, P2_R1113_U84);
  nand ginst9750 (P2_R1113_U303, P2_R1113_U302, P2_R1113_U81);
  nand ginst9751 (P2_R1113_U304, P2_R1113_U177, P2_U3055);
  not ginst9752 (P2_R1113_U305, P2_R1113_U87);
  nand ginst9753 (P2_R1113_U306, P2_R1113_U85, P2_U3056);
  nand ginst9754 (P2_R1113_U307, P2_R1113_U305, P2_R1113_U306);
  nand ginst9755 (P2_R1113_U308, P2_R1113_U86, P2_U3949);
  nand ginst9756 (P2_R1113_U309, P2_R1113_U86, P2_U3949);
  not ginst9757 (P2_R1113_U31, P2_U3441);
  nand ginst9758 (P2_R1113_U310, P2_R1113_U309, P2_R1113_U87);
  nand ginst9759 (P2_R1113_U311, P2_R1113_U85, P2_U3056);
  nand ginst9760 (P2_R1113_U312, P2_R1113_U129, P2_R1113_U310);
  nand ginst9761 (P2_R1113_U313, P2_R1113_U299, P2_R1113_U83);
  nand ginst9762 (P2_R1113_U314, P2_R1113_U133, P2_R1113_U313);
  nand ginst9763 (P2_R1113_U315, P2_R1113_U183, P2_R1113_U88);
  nand ginst9764 (P2_R1113_U316, P2_R1113_U132, P2_R1113_U315);
  nand ginst9765 (P2_R1113_U317, P2_R1113_U183, P2_R1113_U83);
  nand ginst9766 (P2_R1113_U318, P2_R1113_U163, P2_R1113_U287);
  not ginst9767 (P2_R1113_U319, P2_R1113_U89);
  not ginst9768 (P2_R1113_U32, P2_U3073);
  nand ginst9769 (P2_R1113_U320, P2_R1113_U71, P2_U3063);
  nand ginst9770 (P2_R1113_U321, P2_R1113_U319, P2_R1113_U320);
  nand ginst9771 (P2_R1113_U322, P2_R1113_U137, P2_R1113_U321);
  nand ginst9772 (P2_R1113_U323, P2_R1113_U182, P2_R1113_U89);
  nand ginst9773 (P2_R1113_U324, P2_R1113_U73, P2_U3954);
  nand ginst9774 (P2_R1113_U325, P2_R1113_U136, P2_R1113_U323);
  nand ginst9775 (P2_R1113_U326, P2_R1113_U71, P2_U3063);
  nand ginst9776 (P2_R1113_U327, P2_R1113_U182, P2_R1113_U326);
  nand ginst9777 (P2_R1113_U328, P2_R1113_U287, P2_R1113_U76);
  nand ginst9778 (P2_R1113_U329, P2_R1113_U172, P2_R1113_U261);
  not ginst9779 (P2_R1113_U33, P2_U3069);
  not ginst9780 (P2_R1113_U330, P2_R1113_U90);
  nand ginst9781 (P2_R1113_U331, P2_R1113_U56, P2_U3076);
  nand ginst9782 (P2_R1113_U332, P2_R1113_U330, P2_R1113_U331);
  nand ginst9783 (P2_R1113_U333, P2_R1113_U144, P2_R1113_U332);
  nand ginst9784 (P2_R1113_U334, P2_R1113_U181, P2_R1113_U90);
  nand ginst9785 (P2_R1113_U335, P2_R1113_U58, P2_U3477);
  nand ginst9786 (P2_R1113_U336, P2_R1113_U143, P2_R1113_U334);
  nand ginst9787 (P2_R1113_U337, P2_R1113_U56, P2_U3076);
  nand ginst9788 (P2_R1113_U338, P2_R1113_U181, P2_R1113_U337);
  nand ginst9789 (P2_R1113_U339, P2_R1113_U261, P2_R1113_U61);
  not ginst9790 (P2_R1113_U34, P2_U3062);
  nand ginst9791 (P2_R1113_U340, P2_R1113_U150, P2_R1113_U216);
  not ginst9792 (P2_R1113_U341, P2_R1113_U91);
  nand ginst9793 (P2_R1113_U342, P2_R1113_U46, P2_U3064);
  nand ginst9794 (P2_R1113_U343, P2_R1113_U341, P2_R1113_U342);
  nand ginst9795 (P2_R1113_U344, P2_R1113_U148, P2_R1113_U343);
  nand ginst9796 (P2_R1113_U345, P2_R1113_U180, P2_R1113_U91);
  nand ginst9797 (P2_R1113_U346, P2_R1113_U48, P2_U3462);
  nand ginst9798 (P2_R1113_U347, P2_R1113_U147, P2_R1113_U345);
  nand ginst9799 (P2_R1113_U348, P2_R1113_U46, P2_U3064);
  nand ginst9800 (P2_R1113_U349, P2_R1113_U180, P2_R1113_U348);
  nand ginst9801 (P2_R1113_U35, P2_R1113_U31, P2_U3062);
  nand ginst9802 (P2_R1113_U350, P2_R1113_U24, P2_U3079);
  nand ginst9803 (P2_R1113_U351, P2_R1113_U165, P2_U3080);
  nand ginst9804 (P2_R1113_U352, P2_R1113_U130, P2_R1113_U307);
  nand ginst9805 (P2_R1113_U353, P2_R1113_U41, P2_U3456);
  nand ginst9806 (P2_R1113_U354, P2_R1113_U40, P2_U3085);
  nand ginst9807 (P2_R1113_U355, P2_R1113_U150, P2_R1113_U217);
  nand ginst9808 (P2_R1113_U356, P2_R1113_U149, P2_R1113_U215);
  nand ginst9809 (P2_R1113_U357, P2_R1113_U39, P2_U3453);
  nand ginst9810 (P2_R1113_U358, P2_R1113_U36, P2_U3086);
  nand ginst9811 (P2_R1113_U359, P2_R1113_U39, P2_U3453);
  not ginst9812 (P2_R1113_U36, P2_U3453);
  nand ginst9813 (P2_R1113_U360, P2_R1113_U36, P2_U3086);
  nand ginst9814 (P2_R1113_U361, P2_R1113_U359, P2_R1113_U360);
  nand ginst9815 (P2_R1113_U362, P2_R1113_U37, P2_U3450);
  nand ginst9816 (P2_R1113_U363, P2_R1113_U21, P2_U3072);
  nand ginst9817 (P2_R1113_U364, P2_R1113_U222, P2_R1113_U42);
  nand ginst9818 (P2_R1113_U365, P2_R1113_U151, P2_R1113_U209);
  nand ginst9819 (P2_R1113_U366, P2_R1113_U32, P2_U3447);
  nand ginst9820 (P2_R1113_U367, P2_R1113_U30, P2_U3073);
  nand ginst9821 (P2_R1113_U368, P2_R1113_U366, P2_R1113_U367);
  nand ginst9822 (P2_R1113_U369, P2_R1113_U33, P2_U3444);
  not ginst9823 (P2_R1113_U37, P2_U3072);
  nand ginst9824 (P2_R1113_U370, P2_R1113_U22, P2_U3069);
  nand ginst9825 (P2_R1113_U371, P2_R1113_U232, P2_R1113_U43);
  nand ginst9826 (P2_R1113_U372, P2_R1113_U152, P2_R1113_U224);
  nand ginst9827 (P2_R1113_U373, P2_R1113_U34, P2_U3441);
  nand ginst9828 (P2_R1113_U374, P2_R1113_U31, P2_U3062);
  nand ginst9829 (P2_R1113_U375, P2_R1113_U154, P2_R1113_U233);
  nand ginst9830 (P2_R1113_U376, P2_R1113_U153, P2_R1113_U199);
  nand ginst9831 (P2_R1113_U377, P2_R1113_U29, P2_U3438);
  nand ginst9832 (P2_R1113_U378, P2_R1113_U26, P2_U3066);
  nand ginst9833 (P2_R1113_U379, P2_R1113_U29, P2_U3438);
  nand ginst9834 (P2_R1113_U38, P2_R1113_U21, P2_U3072);
  nand ginst9835 (P2_R1113_U380, P2_R1113_U26, P2_U3066);
  nand ginst9836 (P2_R1113_U381, P2_R1113_U379, P2_R1113_U380);
  nand ginst9837 (P2_R1113_U382, P2_R1113_U27, P2_U3435);
  nand ginst9838 (P2_R1113_U383, P2_R1113_U23, P2_U3070);
  nand ginst9839 (P2_R1113_U384, P2_R1113_U238, P2_R1113_U44);
  nand ginst9840 (P2_R1113_U385, P2_R1113_U155, P2_R1113_U193);
  nand ginst9841 (P2_R1113_U386, P2_R1113_U157, P2_U3960);
  nand ginst9842 (P2_R1113_U387, P2_R1113_U156, P2_U3057);
  nand ginst9843 (P2_R1113_U388, P2_R1113_U157, P2_U3960);
  nand ginst9844 (P2_R1113_U389, P2_R1113_U156, P2_U3057);
  not ginst9845 (P2_R1113_U39, P2_U3086);
  nand ginst9846 (P2_R1113_U390, P2_R1113_U388, P2_R1113_U389);
  nand ginst9847 (P2_R1113_U391, P2_R1113_U86, P2_U3949);
  nand ginst9848 (P2_R1113_U392, P2_R1113_U85, P2_U3056);
  not ginst9849 (P2_R1113_U393, P2_R1113_U131);
  nand ginst9850 (P2_R1113_U394, P2_R1113_U305, P2_R1113_U393);
  nand ginst9851 (P2_R1113_U395, P2_R1113_U131, P2_R1113_U87);
  nand ginst9852 (P2_R1113_U396, P2_R1113_U84, P2_U3950);
  nand ginst9853 (P2_R1113_U397, P2_R1113_U81, P2_U3055);
  nand ginst9854 (P2_R1113_U398, P2_R1113_U84, P2_U3950);
  nand ginst9855 (P2_R1113_U399, P2_R1113_U81, P2_U3055);
  not ginst9856 (P2_R1113_U40, P2_U3456);
  nand ginst9857 (P2_R1113_U400, P2_R1113_U398, P2_R1113_U399);
  nand ginst9858 (P2_R1113_U401, P2_R1113_U82, P2_U3951);
  nand ginst9859 (P2_R1113_U402, P2_R1113_U45, P2_U3059);
  nand ginst9860 (P2_R1113_U403, P2_R1113_U317, P2_R1113_U88);
  nand ginst9861 (P2_R1113_U404, P2_R1113_U158, P2_R1113_U299);
  nand ginst9862 (P2_R1113_U405, P2_R1113_U80, P2_U3952);
  nand ginst9863 (P2_R1113_U406, P2_R1113_U79, P2_U3060);
  not ginst9864 (P2_R1113_U407, P2_R1113_U134);
  nand ginst9865 (P2_R1113_U408, P2_R1113_U295, P2_R1113_U407);
  nand ginst9866 (P2_R1113_U409, P2_R1113_U134, P2_R1113_U159);
  not ginst9867 (P2_R1113_U41, P2_U3085);
  nand ginst9868 (P2_R1113_U410, P2_R1113_U78, P2_U3953);
  nand ginst9869 (P2_R1113_U411, P2_R1113_U77, P2_U3067);
  not ginst9870 (P2_R1113_U412, P2_R1113_U135);
  nand ginst9871 (P2_R1113_U413, P2_R1113_U291, P2_R1113_U412);
  nand ginst9872 (P2_R1113_U414, P2_R1113_U135, P2_R1113_U160);
  nand ginst9873 (P2_R1113_U415, P2_R1113_U73, P2_U3954);
  nand ginst9874 (P2_R1113_U416, P2_R1113_U70, P2_U3068);
  nand ginst9875 (P2_R1113_U417, P2_R1113_U415, P2_R1113_U416);
  nand ginst9876 (P2_R1113_U418, P2_R1113_U74, P2_U3955);
  nand ginst9877 (P2_R1113_U419, P2_R1113_U71, P2_U3063);
  nand ginst9878 (P2_R1113_U42, P2_R1113_U207, P2_R1113_U208);
  nand ginst9879 (P2_R1113_U420, P2_R1113_U327, P2_R1113_U89);
  nand ginst9880 (P2_R1113_U421, P2_R1113_U161, P2_R1113_U319);
  nand ginst9881 (P2_R1113_U422, P2_R1113_U75, P2_U3956);
  nand ginst9882 (P2_R1113_U423, P2_R1113_U72, P2_U3077);
  nand ginst9883 (P2_R1113_U424, P2_R1113_U163, P2_R1113_U328);
  nand ginst9884 (P2_R1113_U425, P2_R1113_U162, P2_R1113_U281);
  nand ginst9885 (P2_R1113_U426, P2_R1113_U69, P2_U3957);
  nand ginst9886 (P2_R1113_U427, P2_R1113_U68, P2_U3078);
  not ginst9887 (P2_R1113_U428, P2_R1113_U138);
  nand ginst9888 (P2_R1113_U429, P2_R1113_U277, P2_R1113_U428);
  nand ginst9889 (P2_R1113_U43, P2_R1113_U223, P2_R1113_U35);
  nand ginst9890 (P2_R1113_U430, P2_R1113_U138, P2_R1113_U164);
  nand ginst9891 (P2_R1113_U431, P2_R1113_U25, P2_U3432);
  nand ginst9892 (P2_R1113_U432, P2_R1113_U165, P2_U3080);
  not ginst9893 (P2_R1113_U433, P2_R1113_U139);
  nand ginst9894 (P2_R1113_U434, P2_R1113_U191, P2_R1113_U433);
  nand ginst9895 (P2_R1113_U435, P2_R1113_U139, P2_R1113_U166);
  nand ginst9896 (P2_R1113_U436, P2_R1113_U67, P2_U3485);
  nand ginst9897 (P2_R1113_U437, P2_R1113_U66, P2_U3083);
  not ginst9898 (P2_R1113_U438, P2_R1113_U140);
  nand ginst9899 (P2_R1113_U439, P2_R1113_U273, P2_R1113_U438);
  nand ginst9900 (P2_R1113_U44, P2_R1113_U176, P2_R1113_U192, P2_R1113_U351);
  nand ginst9901 (P2_R1113_U440, P2_R1113_U140, P2_R1113_U167);
  nand ginst9902 (P2_R1113_U441, P2_R1113_U65, P2_U3483);
  nand ginst9903 (P2_R1113_U442, P2_R1113_U168, P2_U3084);
  not ginst9904 (P2_R1113_U443, P2_R1113_U141);
  nand ginst9905 (P2_R1113_U444, P2_R1113_U269, P2_R1113_U443);
  nand ginst9906 (P2_R1113_U445, P2_R1113_U141, P2_R1113_U64);
  nand ginst9907 (P2_R1113_U446, P2_R1113_U63, P2_U3480);
  nand ginst9908 (P2_R1113_U447, P2_R1113_U62, P2_U3071);
  not ginst9909 (P2_R1113_U448, P2_R1113_U142);
  nand ginst9910 (P2_R1113_U449, P2_R1113_U265, P2_R1113_U448);
  not ginst9911 (P2_R1113_U45, P2_U3951);
  nand ginst9912 (P2_R1113_U450, P2_R1113_U142, P2_R1113_U169);
  nand ginst9913 (P2_R1113_U451, P2_R1113_U58, P2_U3477);
  nand ginst9914 (P2_R1113_U452, P2_R1113_U55, P2_U3075);
  nand ginst9915 (P2_R1113_U453, P2_R1113_U451, P2_R1113_U452);
  nand ginst9916 (P2_R1113_U454, P2_R1113_U59, P2_U3474);
  nand ginst9917 (P2_R1113_U455, P2_R1113_U56, P2_U3076);
  nand ginst9918 (P2_R1113_U456, P2_R1113_U338, P2_R1113_U90);
  nand ginst9919 (P2_R1113_U457, P2_R1113_U170, P2_R1113_U330);
  nand ginst9920 (P2_R1113_U458, P2_R1113_U60, P2_U3471);
  nand ginst9921 (P2_R1113_U459, P2_R1113_U57, P2_U3081);
  not ginst9922 (P2_R1113_U46, P2_U3459);
  nand ginst9923 (P2_R1113_U460, P2_R1113_U172, P2_R1113_U339);
  nand ginst9924 (P2_R1113_U461, P2_R1113_U171, P2_R1113_U255);
  nand ginst9925 (P2_R1113_U462, P2_R1113_U54, P2_U3468);
  nand ginst9926 (P2_R1113_U463, P2_R1113_U53, P2_U3082);
  not ginst9927 (P2_R1113_U464, P2_R1113_U145);
  nand ginst9928 (P2_R1113_U465, P2_R1113_U251, P2_R1113_U464);
  nand ginst9929 (P2_R1113_U466, P2_R1113_U145, P2_R1113_U173);
  nand ginst9930 (P2_R1113_U467, P2_R1113_U52, P2_U3465);
  nand ginst9931 (P2_R1113_U468, P2_R1113_U51, P2_U3074);
  not ginst9932 (P2_R1113_U469, P2_R1113_U146);
  not ginst9933 (P2_R1113_U47, P2_U3462);
  nand ginst9934 (P2_R1113_U470, P2_R1113_U247, P2_R1113_U469);
  nand ginst9935 (P2_R1113_U471, P2_R1113_U146, P2_R1113_U174);
  nand ginst9936 (P2_R1113_U472, P2_R1113_U48, P2_U3462);
  nand ginst9937 (P2_R1113_U473, P2_R1113_U47, P2_U3065);
  nand ginst9938 (P2_R1113_U474, P2_R1113_U472, P2_R1113_U473);
  nand ginst9939 (P2_R1113_U475, P2_R1113_U49, P2_U3459);
  nand ginst9940 (P2_R1113_U476, P2_R1113_U46, P2_U3064);
  nand ginst9941 (P2_R1113_U477, P2_R1113_U349, P2_R1113_U91);
  nand ginst9942 (P2_R1113_U478, P2_R1113_U175, P2_R1113_U341);
  not ginst9943 (P2_R1113_U48, P2_U3065);
  not ginst9944 (P2_R1113_U49, P2_U3064);
  nand ginst9945 (P2_R1113_U50, P2_R1113_U40, P2_U3085);
  not ginst9946 (P2_R1113_U51, P2_U3465);
  not ginst9947 (P2_R1113_U52, P2_U3074);
  not ginst9948 (P2_R1113_U53, P2_U3468);
  not ginst9949 (P2_R1113_U54, P2_U3082);
  not ginst9950 (P2_R1113_U55, P2_U3477);
  not ginst9951 (P2_R1113_U56, P2_U3474);
  not ginst9952 (P2_R1113_U57, P2_U3471);
  not ginst9953 (P2_R1113_U58, P2_U3075);
  not ginst9954 (P2_R1113_U59, P2_U3076);
  and ginst9955 (P2_R1113_U6, P2_R1113_U201, P2_R1113_U202);
  not ginst9956 (P2_R1113_U60, P2_U3081);
  nand ginst9957 (P2_R1113_U61, P2_R1113_U57, P2_U3081);
  not ginst9958 (P2_R1113_U62, P2_U3480);
  not ginst9959 (P2_R1113_U63, P2_U3071);
  nand ginst9960 (P2_R1113_U64, P2_R1113_U267, P2_R1113_U268);
  not ginst9961 (P2_R1113_U65, P2_U3084);
  not ginst9962 (P2_R1113_U66, P2_U3485);
  not ginst9963 (P2_R1113_U67, P2_U3083);
  not ginst9964 (P2_R1113_U68, P2_U3957);
  not ginst9965 (P2_R1113_U69, P2_U3078);
  and ginst9966 (P2_R1113_U7, P2_R1113_U240, P2_R1113_U241);
  not ginst9967 (P2_R1113_U70, P2_U3954);
  not ginst9968 (P2_R1113_U71, P2_U3955);
  not ginst9969 (P2_R1113_U72, P2_U3956);
  not ginst9970 (P2_R1113_U73, P2_U3068);
  not ginst9971 (P2_R1113_U74, P2_U3063);
  not ginst9972 (P2_R1113_U75, P2_U3077);
  nand ginst9973 (P2_R1113_U76, P2_R1113_U72, P2_U3077);
  not ginst9974 (P2_R1113_U77, P2_U3953);
  not ginst9975 (P2_R1113_U78, P2_U3067);
  not ginst9976 (P2_R1113_U79, P2_U3952);
  and ginst9977 (P2_R1113_U8, P2_R1113_U181, P2_R1113_U256);
  not ginst9978 (P2_R1113_U80, P2_U3060);
  not ginst9979 (P2_R1113_U81, P2_U3950);
  not ginst9980 (P2_R1113_U82, P2_U3059);
  nand ginst9981 (P2_R1113_U83, P2_R1113_U45, P2_U3059);
  not ginst9982 (P2_R1113_U84, P2_U3055);
  not ginst9983 (P2_R1113_U85, P2_U3949);
  not ginst9984 (P2_R1113_U86, P2_U3056);
  nand ginst9985 (P2_R1113_U87, P2_R1113_U128, P2_R1113_U301);
  nand ginst9986 (P2_R1113_U88, P2_R1113_U297, P2_R1113_U298);
  nand ginst9987 (P2_R1113_U89, P2_R1113_U318, P2_R1113_U76);
  and ginst9988 (P2_R1113_U9, P2_R1113_U257, P2_R1113_U258);
  nand ginst9989 (P2_R1113_U90, P2_R1113_U329, P2_R1113_U61);
  nand ginst9990 (P2_R1113_U91, P2_R1113_U340, P2_R1113_U50);
  not ginst9991 (P2_R1113_U92, P2_U3079);
  nand ginst9992 (P2_R1113_U93, P2_R1113_U394, P2_R1113_U395);
  nand ginst9993 (P2_R1113_U94, P2_R1113_U408, P2_R1113_U409);
  nand ginst9994 (P2_R1113_U95, P2_R1113_U413, P2_R1113_U414);
  nand ginst9995 (P2_R1113_U96, P2_R1113_U429, P2_R1113_U430);
  nand ginst9996 (P2_R1113_U97, P2_R1113_U434, P2_R1113_U435);
  nand ginst9997 (P2_R1113_U98, P2_R1113_U439, P2_R1113_U440);
  nand ginst9998 (P2_R1113_U99, P2_R1113_U444, P2_R1113_U445);
  and ginst9999 (P2_R1131_U10, P2_R1131_U348, P2_R1131_U351);
  nand ginst10000 (P2_R1131_U100, P2_R1131_U398, P2_R1131_U399);
  nand ginst10001 (P2_R1131_U101, P2_R1131_U407, P2_R1131_U408);
  nand ginst10002 (P2_R1131_U102, P2_R1131_U414, P2_R1131_U415);
  nand ginst10003 (P2_R1131_U103, P2_R1131_U421, P2_R1131_U422);
  nand ginst10004 (P2_R1131_U104, P2_R1131_U428, P2_R1131_U429);
  nand ginst10005 (P2_R1131_U105, P2_R1131_U433, P2_R1131_U434);
  nand ginst10006 (P2_R1131_U106, P2_R1131_U440, P2_R1131_U441);
  nand ginst10007 (P2_R1131_U107, P2_R1131_U447, P2_R1131_U448);
  nand ginst10008 (P2_R1131_U108, P2_R1131_U461, P2_R1131_U462);
  nand ginst10009 (P2_R1131_U109, P2_R1131_U466, P2_R1131_U467);
  and ginst10010 (P2_R1131_U11, P2_R1131_U341, P2_R1131_U344);
  nand ginst10011 (P2_R1131_U110, P2_R1131_U473, P2_R1131_U474);
  nand ginst10012 (P2_R1131_U111, P2_R1131_U480, P2_R1131_U481);
  nand ginst10013 (P2_R1131_U112, P2_R1131_U487, P2_R1131_U488);
  nand ginst10014 (P2_R1131_U113, P2_R1131_U494, P2_R1131_U495);
  nand ginst10015 (P2_R1131_U114, P2_R1131_U499, P2_R1131_U500);
  and ginst10016 (P2_R1131_U115, P2_R1131_U187, P2_R1131_U189);
  and ginst10017 (P2_R1131_U116, P2_R1131_U180, P2_R1131_U4);
  and ginst10018 (P2_R1131_U117, P2_R1131_U192, P2_R1131_U194);
  and ginst10019 (P2_R1131_U118, P2_R1131_U200, P2_R1131_U201);
  and ginst10020 (P2_R1131_U119, P2_R1131_U22, P2_R1131_U381, P2_R1131_U382);
  and ginst10021 (P2_R1131_U12, P2_R1131_U332, P2_R1131_U335);
  and ginst10022 (P2_R1131_U120, P2_R1131_U212, P2_R1131_U5);
  and ginst10023 (P2_R1131_U121, P2_R1131_U180, P2_R1131_U181);
  and ginst10024 (P2_R1131_U122, P2_R1131_U218, P2_R1131_U220);
  and ginst10025 (P2_R1131_U123, P2_R1131_U34, P2_R1131_U388, P2_R1131_U389);
  and ginst10026 (P2_R1131_U124, P2_R1131_U226, P2_R1131_U4);
  and ginst10027 (P2_R1131_U125, P2_R1131_U181, P2_R1131_U234);
  and ginst10028 (P2_R1131_U126, P2_R1131_U204, P2_R1131_U6);
  and ginst10029 (P2_R1131_U127, P2_R1131_U171, P2_R1131_U239);
  and ginst10030 (P2_R1131_U128, P2_R1131_U250, P2_R1131_U7);
  and ginst10031 (P2_R1131_U129, P2_R1131_U172, P2_R1131_U248);
  and ginst10032 (P2_R1131_U13, P2_R1131_U323, P2_R1131_U326);
  and ginst10033 (P2_R1131_U130, P2_R1131_U267, P2_R1131_U268);
  and ginst10034 (P2_R1131_U131, P2_R1131_U282, P2_R1131_U9);
  and ginst10035 (P2_R1131_U132, P2_R1131_U280, P2_R1131_U285);
  and ginst10036 (P2_R1131_U133, P2_R1131_U298, P2_R1131_U301);
  and ginst10037 (P2_R1131_U134, P2_R1131_U302, P2_R1131_U368);
  and ginst10038 (P2_R1131_U135, P2_R1131_U160, P2_R1131_U278);
  and ginst10039 (P2_R1131_U136, P2_R1131_U454, P2_R1131_U455, P2_R1131_U80);
  and ginst10040 (P2_R1131_U137, P2_R1131_U325, P2_R1131_U9);
  and ginst10041 (P2_R1131_U138, P2_R1131_U468, P2_R1131_U469, P2_R1131_U59);
  and ginst10042 (P2_R1131_U139, P2_R1131_U334, P2_R1131_U8);
  and ginst10043 (P2_R1131_U14, P2_R1131_U318, P2_R1131_U320);
  and ginst10044 (P2_R1131_U140, P2_R1131_U172, P2_R1131_U489, P2_R1131_U490);
  and ginst10045 (P2_R1131_U141, P2_R1131_U343, P2_R1131_U7);
  and ginst10046 (P2_R1131_U142, P2_R1131_U171, P2_R1131_U501, P2_R1131_U502);
  and ginst10047 (P2_R1131_U143, P2_R1131_U350, P2_R1131_U6);
  nand ginst10048 (P2_R1131_U144, P2_R1131_U118, P2_R1131_U202);
  nand ginst10049 (P2_R1131_U145, P2_R1131_U217, P2_R1131_U229);
  not ginst10050 (P2_R1131_U146, P2_U3057);
  not ginst10051 (P2_R1131_U147, P2_U3960);
  and ginst10052 (P2_R1131_U148, P2_R1131_U402, P2_R1131_U403);
  nand ginst10053 (P2_R1131_U149, P2_R1131_U169, P2_R1131_U304, P2_R1131_U364);
  and ginst10054 (P2_R1131_U15, P2_R1131_U310, P2_R1131_U313);
  and ginst10055 (P2_R1131_U150, P2_R1131_U409, P2_R1131_U410);
  nand ginst10056 (P2_R1131_U151, P2_R1131_U134, P2_R1131_U369, P2_R1131_U370);
  and ginst10057 (P2_R1131_U152, P2_R1131_U416, P2_R1131_U417);
  nand ginst10058 (P2_R1131_U153, P2_R1131_U299, P2_R1131_U365, P2_R1131_U86);
  and ginst10059 (P2_R1131_U154, P2_R1131_U423, P2_R1131_U424);
  nand ginst10060 (P2_R1131_U155, P2_R1131_U292, P2_R1131_U293);
  and ginst10061 (P2_R1131_U156, P2_R1131_U435, P2_R1131_U436);
  nand ginst10062 (P2_R1131_U157, P2_R1131_U288, P2_R1131_U289);
  and ginst10063 (P2_R1131_U158, P2_R1131_U442, P2_R1131_U443);
  nand ginst10064 (P2_R1131_U159, P2_R1131_U132, P2_R1131_U284);
  and ginst10065 (P2_R1131_U16, P2_R1131_U232, P2_R1131_U235);
  and ginst10066 (P2_R1131_U160, P2_R1131_U449, P2_R1131_U450);
  nand ginst10067 (P2_R1131_U161, P2_R1131_U327, P2_R1131_U43);
  nand ginst10068 (P2_R1131_U162, P2_R1131_U130, P2_R1131_U269);
  and ginst10069 (P2_R1131_U163, P2_R1131_U475, P2_R1131_U476);
  nand ginst10070 (P2_R1131_U164, P2_R1131_U256, P2_R1131_U257);
  and ginst10071 (P2_R1131_U165, P2_R1131_U482, P2_R1131_U483);
  nand ginst10072 (P2_R1131_U166, P2_R1131_U252, P2_R1131_U253);
  nand ginst10073 (P2_R1131_U167, P2_R1131_U242, P2_R1131_U243);
  nand ginst10074 (P2_R1131_U168, P2_R1131_U366, P2_R1131_U367);
  nand ginst10075 (P2_R1131_U169, P2_R1131_U151, P2_U3056);
  and ginst10076 (P2_R1131_U17, P2_R1131_U224, P2_R1131_U227);
  not ginst10077 (P2_R1131_U170, P2_R1131_U34);
  nand ginst10078 (P2_R1131_U171, P2_U3085, P2_U3456);
  nand ginst10079 (P2_R1131_U172, P2_U3074, P2_U3465);
  nand ginst10080 (P2_R1131_U173, P2_U3060, P2_U3952);
  not ginst10081 (P2_R1131_U174, P2_R1131_U68);
  not ginst10082 (P2_R1131_U175, P2_R1131_U77);
  nand ginst10083 (P2_R1131_U176, P2_U3067, P2_U3953);
  not ginst10084 (P2_R1131_U177, P2_R1131_U61);
  or ginst10085 (P2_R1131_U178, P2_U3069, P2_U3444);
  or ginst10086 (P2_R1131_U179, P2_U3062, P2_U3441);
  and ginst10087 (P2_R1131_U18, P2_R1131_U210, P2_R1131_U213);
  or ginst10088 (P2_R1131_U180, P2_U3066, P2_U3438);
  or ginst10089 (P2_R1131_U181, P2_U3070, P2_U3435);
  not ginst10090 (P2_R1131_U182, P2_R1131_U31);
  or ginst10091 (P2_R1131_U183, P2_U3080, P2_U3432);
  not ginst10092 (P2_R1131_U184, P2_R1131_U42);
  not ginst10093 (P2_R1131_U185, P2_R1131_U43);
  nand ginst10094 (P2_R1131_U186, P2_R1131_U42, P2_R1131_U43);
  nand ginst10095 (P2_R1131_U187, P2_U3070, P2_U3435);
  nand ginst10096 (P2_R1131_U188, P2_R1131_U181, P2_R1131_U186);
  nand ginst10097 (P2_R1131_U189, P2_U3066, P2_U3438);
  not ginst10098 (P2_R1131_U19, P2_U3447);
  nand ginst10099 (P2_R1131_U190, P2_R1131_U115, P2_R1131_U188);
  nand ginst10100 (P2_R1131_U191, P2_R1131_U34, P2_R1131_U35);
  nand ginst10101 (P2_R1131_U192, P2_R1131_U191, P2_U3069);
  nand ginst10102 (P2_R1131_U193, P2_R1131_U116, P2_R1131_U190);
  nand ginst10103 (P2_R1131_U194, P2_R1131_U170, P2_U3444);
  not ginst10104 (P2_R1131_U195, P2_R1131_U41);
  or ginst10105 (P2_R1131_U196, P2_U3072, P2_U3450);
  or ginst10106 (P2_R1131_U197, P2_U3073, P2_U3447);
  not ginst10107 (P2_R1131_U198, P2_R1131_U22);
  nand ginst10108 (P2_R1131_U199, P2_R1131_U22, P2_R1131_U23);
  not ginst10109 (P2_R1131_U20, P2_U3073);
  nand ginst10110 (P2_R1131_U200, P2_R1131_U199, P2_U3072);
  nand ginst10111 (P2_R1131_U201, P2_R1131_U198, P2_U3450);
  nand ginst10112 (P2_R1131_U202, P2_R1131_U41, P2_R1131_U5);
  not ginst10113 (P2_R1131_U203, P2_R1131_U144);
  or ginst10114 (P2_R1131_U204, P2_U3086, P2_U3453);
  nand ginst10115 (P2_R1131_U205, P2_R1131_U144, P2_R1131_U204);
  not ginst10116 (P2_R1131_U206, P2_R1131_U40);
  or ginst10117 (P2_R1131_U207, P2_U3085, P2_U3456);
  or ginst10118 (P2_R1131_U208, P2_U3073, P2_U3447);
  nand ginst10119 (P2_R1131_U209, P2_R1131_U208, P2_R1131_U41);
  not ginst10120 (P2_R1131_U21, P2_U3072);
  nand ginst10121 (P2_R1131_U210, P2_R1131_U119, P2_R1131_U209);
  nand ginst10122 (P2_R1131_U211, P2_R1131_U195, P2_R1131_U22);
  nand ginst10123 (P2_R1131_U212, P2_U3072, P2_U3450);
  nand ginst10124 (P2_R1131_U213, P2_R1131_U120, P2_R1131_U211);
  or ginst10125 (P2_R1131_U214, P2_U3073, P2_U3447);
  nand ginst10126 (P2_R1131_U215, P2_R1131_U181, P2_R1131_U185);
  nand ginst10127 (P2_R1131_U216, P2_U3070, P2_U3435);
  not ginst10128 (P2_R1131_U217, P2_R1131_U45);
  nand ginst10129 (P2_R1131_U218, P2_R1131_U121, P2_R1131_U184);
  nand ginst10130 (P2_R1131_U219, P2_R1131_U180, P2_R1131_U45);
  nand ginst10131 (P2_R1131_U22, P2_U3073, P2_U3447);
  nand ginst10132 (P2_R1131_U220, P2_U3066, P2_U3438);
  not ginst10133 (P2_R1131_U221, P2_R1131_U44);
  or ginst10134 (P2_R1131_U222, P2_U3062, P2_U3441);
  nand ginst10135 (P2_R1131_U223, P2_R1131_U222, P2_R1131_U44);
  nand ginst10136 (P2_R1131_U224, P2_R1131_U123, P2_R1131_U223);
  nand ginst10137 (P2_R1131_U225, P2_R1131_U221, P2_R1131_U34);
  nand ginst10138 (P2_R1131_U226, P2_U3069, P2_U3444);
  nand ginst10139 (P2_R1131_U227, P2_R1131_U124, P2_R1131_U225);
  or ginst10140 (P2_R1131_U228, P2_U3062, P2_U3441);
  nand ginst10141 (P2_R1131_U229, P2_R1131_U181, P2_R1131_U184);
  not ginst10142 (P2_R1131_U23, P2_U3450);
  not ginst10143 (P2_R1131_U230, P2_R1131_U145);
  nand ginst10144 (P2_R1131_U231, P2_U3066, P2_U3438);
  nand ginst10145 (P2_R1131_U232, P2_R1131_U400, P2_R1131_U401, P2_R1131_U42, P2_R1131_U43);
  nand ginst10146 (P2_R1131_U233, P2_R1131_U42, P2_R1131_U43);
  nand ginst10147 (P2_R1131_U234, P2_U3070, P2_U3435);
  nand ginst10148 (P2_R1131_U235, P2_R1131_U125, P2_R1131_U233);
  or ginst10149 (P2_R1131_U236, P2_U3085, P2_U3456);
  or ginst10150 (P2_R1131_U237, P2_U3064, P2_U3459);
  nand ginst10151 (P2_R1131_U238, P2_R1131_U177, P2_R1131_U6);
  nand ginst10152 (P2_R1131_U239, P2_U3064, P2_U3459);
  not ginst10153 (P2_R1131_U24, P2_U3441);
  nand ginst10154 (P2_R1131_U240, P2_R1131_U127, P2_R1131_U238);
  or ginst10155 (P2_R1131_U241, P2_U3064, P2_U3459);
  nand ginst10156 (P2_R1131_U242, P2_R1131_U126, P2_R1131_U144);
  nand ginst10157 (P2_R1131_U243, P2_R1131_U240, P2_R1131_U241);
  not ginst10158 (P2_R1131_U244, P2_R1131_U167);
  or ginst10159 (P2_R1131_U245, P2_U3082, P2_U3468);
  or ginst10160 (P2_R1131_U246, P2_U3074, P2_U3465);
  nand ginst10161 (P2_R1131_U247, P2_R1131_U174, P2_R1131_U7);
  nand ginst10162 (P2_R1131_U248, P2_U3082, P2_U3468);
  nand ginst10163 (P2_R1131_U249, P2_R1131_U129, P2_R1131_U247);
  not ginst10164 (P2_R1131_U25, P2_U3062);
  or ginst10165 (P2_R1131_U250, P2_U3065, P2_U3462);
  or ginst10166 (P2_R1131_U251, P2_U3082, P2_U3468);
  nand ginst10167 (P2_R1131_U252, P2_R1131_U128, P2_R1131_U167);
  nand ginst10168 (P2_R1131_U253, P2_R1131_U249, P2_R1131_U251);
  not ginst10169 (P2_R1131_U254, P2_R1131_U166);
  or ginst10170 (P2_R1131_U255, P2_U3081, P2_U3471);
  nand ginst10171 (P2_R1131_U256, P2_R1131_U166, P2_R1131_U255);
  nand ginst10172 (P2_R1131_U257, P2_U3081, P2_U3471);
  not ginst10173 (P2_R1131_U258, P2_R1131_U164);
  or ginst10174 (P2_R1131_U259, P2_U3076, P2_U3474);
  not ginst10175 (P2_R1131_U26, P2_U3069);
  nand ginst10176 (P2_R1131_U260, P2_R1131_U164, P2_R1131_U259);
  nand ginst10177 (P2_R1131_U261, P2_U3076, P2_U3474);
  not ginst10178 (P2_R1131_U262, P2_R1131_U92);
  or ginst10179 (P2_R1131_U263, P2_U3071, P2_U3480);
  or ginst10180 (P2_R1131_U264, P2_U3075, P2_U3477);
  not ginst10181 (P2_R1131_U265, P2_R1131_U59);
  nand ginst10182 (P2_R1131_U266, P2_R1131_U59, P2_R1131_U60);
  nand ginst10183 (P2_R1131_U267, P2_R1131_U266, P2_U3071);
  nand ginst10184 (P2_R1131_U268, P2_R1131_U265, P2_U3480);
  nand ginst10185 (P2_R1131_U269, P2_R1131_U8, P2_R1131_U92);
  not ginst10186 (P2_R1131_U27, P2_U3435);
  not ginst10187 (P2_R1131_U270, P2_R1131_U162);
  or ginst10188 (P2_R1131_U271, P2_U3078, P2_U3957);
  or ginst10189 (P2_R1131_U272, P2_U3083, P2_U3485);
  or ginst10190 (P2_R1131_U273, P2_U3077, P2_U3956);
  not ginst10191 (P2_R1131_U274, P2_R1131_U80);
  nand ginst10192 (P2_R1131_U275, P2_R1131_U274, P2_U3957);
  nand ginst10193 (P2_R1131_U276, P2_R1131_U275, P2_R1131_U90);
  nand ginst10194 (P2_R1131_U277, P2_R1131_U80, P2_R1131_U81);
  nand ginst10195 (P2_R1131_U278, P2_R1131_U276, P2_R1131_U277);
  nand ginst10196 (P2_R1131_U279, P2_R1131_U175, P2_R1131_U9);
  not ginst10197 (P2_R1131_U28, P2_U3070);
  nand ginst10198 (P2_R1131_U280, P2_U3077, P2_U3956);
  nand ginst10199 (P2_R1131_U281, P2_R1131_U278, P2_R1131_U279);
  or ginst10200 (P2_R1131_U282, P2_U3084, P2_U3483);
  or ginst10201 (P2_R1131_U283, P2_U3077, P2_U3956);
  nand ginst10202 (P2_R1131_U284, P2_R1131_U131, P2_R1131_U162, P2_R1131_U273);
  nand ginst10203 (P2_R1131_U285, P2_R1131_U281, P2_R1131_U283);
  not ginst10204 (P2_R1131_U286, P2_R1131_U159);
  or ginst10205 (P2_R1131_U287, P2_U3063, P2_U3955);
  nand ginst10206 (P2_R1131_U288, P2_R1131_U159, P2_R1131_U287);
  nand ginst10207 (P2_R1131_U289, P2_U3063, P2_U3955);
  not ginst10208 (P2_R1131_U29, P2_U3427);
  not ginst10209 (P2_R1131_U290, P2_R1131_U157);
  or ginst10210 (P2_R1131_U291, P2_U3068, P2_U3954);
  nand ginst10211 (P2_R1131_U292, P2_R1131_U157, P2_R1131_U291);
  nand ginst10212 (P2_R1131_U293, P2_U3068, P2_U3954);
  not ginst10213 (P2_R1131_U294, P2_R1131_U155);
  or ginst10214 (P2_R1131_U295, P2_U3060, P2_U3952);
  nand ginst10215 (P2_R1131_U296, P2_R1131_U173, P2_R1131_U176);
  not ginst10216 (P2_R1131_U297, P2_R1131_U86);
  or ginst10217 (P2_R1131_U298, P2_U3067, P2_U3953);
  nand ginst10218 (P2_R1131_U299, P2_R1131_U155, P2_R1131_U168, P2_R1131_U298);
  not ginst10219 (P2_R1131_U30, P2_U3079);
  not ginst10220 (P2_R1131_U300, P2_R1131_U153);
  or ginst10221 (P2_R1131_U301, P2_U3055, P2_U3950);
  nand ginst10222 (P2_R1131_U302, P2_U3055, P2_U3950);
  not ginst10223 (P2_R1131_U303, P2_R1131_U151);
  nand ginst10224 (P2_R1131_U304, P2_R1131_U151, P2_U3949);
  not ginst10225 (P2_R1131_U305, P2_R1131_U149);
  nand ginst10226 (P2_R1131_U306, P2_R1131_U155, P2_R1131_U298);
  not ginst10227 (P2_R1131_U307, P2_R1131_U89);
  or ginst10228 (P2_R1131_U308, P2_U3060, P2_U3952);
  nand ginst10229 (P2_R1131_U309, P2_R1131_U308, P2_R1131_U89);
  nand ginst10230 (P2_R1131_U31, P2_U3079, P2_U3427);
  nand ginst10231 (P2_R1131_U310, P2_R1131_U154, P2_R1131_U173, P2_R1131_U309);
  nand ginst10232 (P2_R1131_U311, P2_R1131_U173, P2_R1131_U307);
  nand ginst10233 (P2_R1131_U312, P2_U3059, P2_U3951);
  nand ginst10234 (P2_R1131_U313, P2_R1131_U168, P2_R1131_U311, P2_R1131_U312);
  or ginst10235 (P2_R1131_U314, P2_U3060, P2_U3952);
  nand ginst10236 (P2_R1131_U315, P2_R1131_U162, P2_R1131_U282);
  not ginst10237 (P2_R1131_U316, P2_R1131_U91);
  nand ginst10238 (P2_R1131_U317, P2_R1131_U9, P2_R1131_U91);
  nand ginst10239 (P2_R1131_U318, P2_R1131_U135, P2_R1131_U317);
  nand ginst10240 (P2_R1131_U319, P2_R1131_U278, P2_R1131_U317);
  not ginst10241 (P2_R1131_U32, P2_U3438);
  nand ginst10242 (P2_R1131_U320, P2_R1131_U319, P2_R1131_U453);
  or ginst10243 (P2_R1131_U321, P2_U3083, P2_U3485);
  nand ginst10244 (P2_R1131_U322, P2_R1131_U321, P2_R1131_U91);
  nand ginst10245 (P2_R1131_U323, P2_R1131_U136, P2_R1131_U322);
  nand ginst10246 (P2_R1131_U324, P2_R1131_U316, P2_R1131_U80);
  nand ginst10247 (P2_R1131_U325, P2_U3078, P2_U3957);
  nand ginst10248 (P2_R1131_U326, P2_R1131_U137, P2_R1131_U324);
  or ginst10249 (P2_R1131_U327, P2_U3080, P2_U3432);
  not ginst10250 (P2_R1131_U328, P2_R1131_U161);
  or ginst10251 (P2_R1131_U329, P2_U3083, P2_U3485);
  not ginst10252 (P2_R1131_U33, P2_U3066);
  or ginst10253 (P2_R1131_U330, P2_U3075, P2_U3477);
  nand ginst10254 (P2_R1131_U331, P2_R1131_U330, P2_R1131_U92);
  nand ginst10255 (P2_R1131_U332, P2_R1131_U138, P2_R1131_U331);
  nand ginst10256 (P2_R1131_U333, P2_R1131_U262, P2_R1131_U59);
  nand ginst10257 (P2_R1131_U334, P2_U3071, P2_U3480);
  nand ginst10258 (P2_R1131_U335, P2_R1131_U139, P2_R1131_U333);
  or ginst10259 (P2_R1131_U336, P2_U3075, P2_U3477);
  nand ginst10260 (P2_R1131_U337, P2_R1131_U167, P2_R1131_U250);
  not ginst10261 (P2_R1131_U338, P2_R1131_U93);
  or ginst10262 (P2_R1131_U339, P2_U3074, P2_U3465);
  nand ginst10263 (P2_R1131_U34, P2_U3062, P2_U3441);
  nand ginst10264 (P2_R1131_U340, P2_R1131_U339, P2_R1131_U93);
  nand ginst10265 (P2_R1131_U341, P2_R1131_U140, P2_R1131_U340);
  nand ginst10266 (P2_R1131_U342, P2_R1131_U172, P2_R1131_U338);
  nand ginst10267 (P2_R1131_U343, P2_U3082, P2_U3468);
  nand ginst10268 (P2_R1131_U344, P2_R1131_U141, P2_R1131_U342);
  or ginst10269 (P2_R1131_U345, P2_U3074, P2_U3465);
  or ginst10270 (P2_R1131_U346, P2_U3085, P2_U3456);
  nand ginst10271 (P2_R1131_U347, P2_R1131_U346, P2_R1131_U40);
  nand ginst10272 (P2_R1131_U348, P2_R1131_U142, P2_R1131_U347);
  nand ginst10273 (P2_R1131_U349, P2_R1131_U171, P2_R1131_U206);
  not ginst10274 (P2_R1131_U35, P2_U3444);
  nand ginst10275 (P2_R1131_U350, P2_U3064, P2_U3459);
  nand ginst10276 (P2_R1131_U351, P2_R1131_U143, P2_R1131_U349);
  nand ginst10277 (P2_R1131_U352, P2_R1131_U171, P2_R1131_U207);
  nand ginst10278 (P2_R1131_U353, P2_R1131_U204, P2_R1131_U61);
  nand ginst10279 (P2_R1131_U354, P2_R1131_U214, P2_R1131_U22);
  nand ginst10280 (P2_R1131_U355, P2_R1131_U228, P2_R1131_U34);
  nand ginst10281 (P2_R1131_U356, P2_R1131_U180, P2_R1131_U231);
  nand ginst10282 (P2_R1131_U357, P2_R1131_U173, P2_R1131_U314);
  nand ginst10283 (P2_R1131_U358, P2_R1131_U176, P2_R1131_U298);
  nand ginst10284 (P2_R1131_U359, P2_R1131_U329, P2_R1131_U80);
  not ginst10285 (P2_R1131_U36, P2_U3453);
  nand ginst10286 (P2_R1131_U360, P2_R1131_U282, P2_R1131_U77);
  nand ginst10287 (P2_R1131_U361, P2_R1131_U336, P2_R1131_U59);
  nand ginst10288 (P2_R1131_U362, P2_R1131_U172, P2_R1131_U345);
  nand ginst10289 (P2_R1131_U363, P2_R1131_U250, P2_R1131_U68);
  nand ginst10290 (P2_R1131_U364, P2_U3056, P2_U3949);
  nand ginst10291 (P2_R1131_U365, P2_R1131_U168, P2_R1131_U296);
  nand ginst10292 (P2_R1131_U366, P2_R1131_U295, P2_U3059);
  nand ginst10293 (P2_R1131_U367, P2_R1131_U295, P2_U3951);
  nand ginst10294 (P2_R1131_U368, P2_R1131_U168, P2_R1131_U296, P2_R1131_U301);
  nand ginst10295 (P2_R1131_U369, P2_R1131_U133, P2_R1131_U155, P2_R1131_U168);
  not ginst10296 (P2_R1131_U37, P2_U3086);
  nand ginst10297 (P2_R1131_U370, P2_R1131_U297, P2_R1131_U301);
  nand ginst10298 (P2_R1131_U371, P2_R1131_U39, P2_U3085);
  nand ginst10299 (P2_R1131_U372, P2_R1131_U38, P2_U3456);
  nand ginst10300 (P2_R1131_U373, P2_R1131_U371, P2_R1131_U372);
  nand ginst10301 (P2_R1131_U374, P2_R1131_U352, P2_R1131_U40);
  nand ginst10302 (P2_R1131_U375, P2_R1131_U206, P2_R1131_U373);
  nand ginst10303 (P2_R1131_U376, P2_R1131_U36, P2_U3086);
  nand ginst10304 (P2_R1131_U377, P2_R1131_U37, P2_U3453);
  nand ginst10305 (P2_R1131_U378, P2_R1131_U376, P2_R1131_U377);
  nand ginst10306 (P2_R1131_U379, P2_R1131_U144, P2_R1131_U353);
  not ginst10307 (P2_R1131_U38, P2_U3085);
  nand ginst10308 (P2_R1131_U380, P2_R1131_U203, P2_R1131_U378);
  nand ginst10309 (P2_R1131_U381, P2_R1131_U23, P2_U3072);
  nand ginst10310 (P2_R1131_U382, P2_R1131_U21, P2_U3450);
  nand ginst10311 (P2_R1131_U383, P2_R1131_U19, P2_U3073);
  nand ginst10312 (P2_R1131_U384, P2_R1131_U20, P2_U3447);
  nand ginst10313 (P2_R1131_U385, P2_R1131_U383, P2_R1131_U384);
  nand ginst10314 (P2_R1131_U386, P2_R1131_U354, P2_R1131_U41);
  nand ginst10315 (P2_R1131_U387, P2_R1131_U195, P2_R1131_U385);
  nand ginst10316 (P2_R1131_U388, P2_R1131_U35, P2_U3069);
  nand ginst10317 (P2_R1131_U389, P2_R1131_U26, P2_U3444);
  not ginst10318 (P2_R1131_U39, P2_U3456);
  nand ginst10319 (P2_R1131_U390, P2_R1131_U24, P2_U3062);
  nand ginst10320 (P2_R1131_U391, P2_R1131_U25, P2_U3441);
  nand ginst10321 (P2_R1131_U392, P2_R1131_U390, P2_R1131_U391);
  nand ginst10322 (P2_R1131_U393, P2_R1131_U355, P2_R1131_U44);
  nand ginst10323 (P2_R1131_U394, P2_R1131_U221, P2_R1131_U392);
  nand ginst10324 (P2_R1131_U395, P2_R1131_U32, P2_U3066);
  nand ginst10325 (P2_R1131_U396, P2_R1131_U33, P2_U3438);
  nand ginst10326 (P2_R1131_U397, P2_R1131_U395, P2_R1131_U396);
  nand ginst10327 (P2_R1131_U398, P2_R1131_U145, P2_R1131_U356);
  nand ginst10328 (P2_R1131_U399, P2_R1131_U230, P2_R1131_U397);
  and ginst10329 (P2_R1131_U4, P2_R1131_U178, P2_R1131_U179);
  nand ginst10330 (P2_R1131_U40, P2_R1131_U205, P2_R1131_U61);
  nand ginst10331 (P2_R1131_U400, P2_R1131_U27, P2_U3070);
  nand ginst10332 (P2_R1131_U401, P2_R1131_U28, P2_U3435);
  nand ginst10333 (P2_R1131_U402, P2_R1131_U147, P2_U3057);
  nand ginst10334 (P2_R1131_U403, P2_R1131_U146, P2_U3960);
  nand ginst10335 (P2_R1131_U404, P2_R1131_U147, P2_U3057);
  nand ginst10336 (P2_R1131_U405, P2_R1131_U146, P2_U3960);
  nand ginst10337 (P2_R1131_U406, P2_R1131_U404, P2_R1131_U405);
  nand ginst10338 (P2_R1131_U407, P2_R1131_U148, P2_R1131_U149);
  nand ginst10339 (P2_R1131_U408, P2_R1131_U305, P2_R1131_U406);
  nand ginst10340 (P2_R1131_U409, P2_R1131_U88, P2_U3056);
  nand ginst10341 (P2_R1131_U41, P2_R1131_U117, P2_R1131_U193);
  nand ginst10342 (P2_R1131_U410, P2_R1131_U87, P2_U3949);
  nand ginst10343 (P2_R1131_U411, P2_R1131_U88, P2_U3056);
  nand ginst10344 (P2_R1131_U412, P2_R1131_U87, P2_U3949);
  nand ginst10345 (P2_R1131_U413, P2_R1131_U411, P2_R1131_U412);
  nand ginst10346 (P2_R1131_U414, P2_R1131_U150, P2_R1131_U151);
  nand ginst10347 (P2_R1131_U415, P2_R1131_U303, P2_R1131_U413);
  nand ginst10348 (P2_R1131_U416, P2_R1131_U46, P2_U3055);
  nand ginst10349 (P2_R1131_U417, P2_R1131_U47, P2_U3950);
  nand ginst10350 (P2_R1131_U418, P2_R1131_U46, P2_U3055);
  nand ginst10351 (P2_R1131_U419, P2_R1131_U47, P2_U3950);
  nand ginst10352 (P2_R1131_U42, P2_R1131_U182, P2_R1131_U183);
  nand ginst10353 (P2_R1131_U420, P2_R1131_U418, P2_R1131_U419);
  nand ginst10354 (P2_R1131_U421, P2_R1131_U152, P2_R1131_U153);
  nand ginst10355 (P2_R1131_U422, P2_R1131_U300, P2_R1131_U420);
  nand ginst10356 (P2_R1131_U423, P2_R1131_U49, P2_U3059);
  nand ginst10357 (P2_R1131_U424, P2_R1131_U48, P2_U3951);
  nand ginst10358 (P2_R1131_U425, P2_R1131_U50, P2_U3060);
  nand ginst10359 (P2_R1131_U426, P2_R1131_U51, P2_U3952);
  nand ginst10360 (P2_R1131_U427, P2_R1131_U425, P2_R1131_U426);
  nand ginst10361 (P2_R1131_U428, P2_R1131_U357, P2_R1131_U89);
  nand ginst10362 (P2_R1131_U429, P2_R1131_U307, P2_R1131_U427);
  nand ginst10363 (P2_R1131_U43, P2_U3080, P2_U3432);
  nand ginst10364 (P2_R1131_U430, P2_R1131_U52, P2_U3067);
  nand ginst10365 (P2_R1131_U431, P2_R1131_U53, P2_U3953);
  nand ginst10366 (P2_R1131_U432, P2_R1131_U430, P2_R1131_U431);
  nand ginst10367 (P2_R1131_U433, P2_R1131_U155, P2_R1131_U358);
  nand ginst10368 (P2_R1131_U434, P2_R1131_U294, P2_R1131_U432);
  nand ginst10369 (P2_R1131_U435, P2_R1131_U84, P2_U3068);
  nand ginst10370 (P2_R1131_U436, P2_R1131_U85, P2_U3954);
  nand ginst10371 (P2_R1131_U437, P2_R1131_U84, P2_U3068);
  nand ginst10372 (P2_R1131_U438, P2_R1131_U85, P2_U3954);
  nand ginst10373 (P2_R1131_U439, P2_R1131_U437, P2_R1131_U438);
  nand ginst10374 (P2_R1131_U44, P2_R1131_U122, P2_R1131_U219);
  nand ginst10375 (P2_R1131_U440, P2_R1131_U156, P2_R1131_U157);
  nand ginst10376 (P2_R1131_U441, P2_R1131_U290, P2_R1131_U439);
  nand ginst10377 (P2_R1131_U442, P2_R1131_U82, P2_U3063);
  nand ginst10378 (P2_R1131_U443, P2_R1131_U83, P2_U3955);
  nand ginst10379 (P2_R1131_U444, P2_R1131_U82, P2_U3063);
  nand ginst10380 (P2_R1131_U445, P2_R1131_U83, P2_U3955);
  nand ginst10381 (P2_R1131_U446, P2_R1131_U444, P2_R1131_U445);
  nand ginst10382 (P2_R1131_U447, P2_R1131_U158, P2_R1131_U159);
  nand ginst10383 (P2_R1131_U448, P2_R1131_U286, P2_R1131_U446);
  nand ginst10384 (P2_R1131_U449, P2_R1131_U54, P2_U3077);
  nand ginst10385 (P2_R1131_U45, P2_R1131_U215, P2_R1131_U216);
  nand ginst10386 (P2_R1131_U450, P2_R1131_U55, P2_U3956);
  nand ginst10387 (P2_R1131_U451, P2_R1131_U54, P2_U3077);
  nand ginst10388 (P2_R1131_U452, P2_R1131_U55, P2_U3956);
  nand ginst10389 (P2_R1131_U453, P2_R1131_U451, P2_R1131_U452);
  nand ginst10390 (P2_R1131_U454, P2_R1131_U81, P2_U3078);
  nand ginst10391 (P2_R1131_U455, P2_R1131_U90, P2_U3957);
  nand ginst10392 (P2_R1131_U456, P2_R1131_U161, P2_R1131_U182);
  nand ginst10393 (P2_R1131_U457, P2_R1131_U31, P2_R1131_U328);
  nand ginst10394 (P2_R1131_U458, P2_R1131_U78, P2_U3083);
  nand ginst10395 (P2_R1131_U459, P2_R1131_U79, P2_U3485);
  not ginst10396 (P2_R1131_U46, P2_U3950);
  nand ginst10397 (P2_R1131_U460, P2_R1131_U458, P2_R1131_U459);
  nand ginst10398 (P2_R1131_U461, P2_R1131_U359, P2_R1131_U91);
  nand ginst10399 (P2_R1131_U462, P2_R1131_U316, P2_R1131_U460);
  nand ginst10400 (P2_R1131_U463, P2_R1131_U75, P2_U3084);
  nand ginst10401 (P2_R1131_U464, P2_R1131_U76, P2_U3483);
  nand ginst10402 (P2_R1131_U465, P2_R1131_U463, P2_R1131_U464);
  nand ginst10403 (P2_R1131_U466, P2_R1131_U162, P2_R1131_U360);
  nand ginst10404 (P2_R1131_U467, P2_R1131_U270, P2_R1131_U465);
  nand ginst10405 (P2_R1131_U468, P2_R1131_U60, P2_U3071);
  nand ginst10406 (P2_R1131_U469, P2_R1131_U58, P2_U3480);
  not ginst10407 (P2_R1131_U47, P2_U3055);
  nand ginst10408 (P2_R1131_U470, P2_R1131_U56, P2_U3075);
  nand ginst10409 (P2_R1131_U471, P2_R1131_U57, P2_U3477);
  nand ginst10410 (P2_R1131_U472, P2_R1131_U470, P2_R1131_U471);
  nand ginst10411 (P2_R1131_U473, P2_R1131_U361, P2_R1131_U92);
  nand ginst10412 (P2_R1131_U474, P2_R1131_U262, P2_R1131_U472);
  nand ginst10413 (P2_R1131_U475, P2_R1131_U73, P2_U3076);
  nand ginst10414 (P2_R1131_U476, P2_R1131_U74, P2_U3474);
  nand ginst10415 (P2_R1131_U477, P2_R1131_U73, P2_U3076);
  nand ginst10416 (P2_R1131_U478, P2_R1131_U74, P2_U3474);
  nand ginst10417 (P2_R1131_U479, P2_R1131_U477, P2_R1131_U478);
  not ginst10418 (P2_R1131_U48, P2_U3059);
  nand ginst10419 (P2_R1131_U480, P2_R1131_U163, P2_R1131_U164);
  nand ginst10420 (P2_R1131_U481, P2_R1131_U258, P2_R1131_U479);
  nand ginst10421 (P2_R1131_U482, P2_R1131_U71, P2_U3081);
  nand ginst10422 (P2_R1131_U483, P2_R1131_U72, P2_U3471);
  nand ginst10423 (P2_R1131_U484, P2_R1131_U71, P2_U3081);
  nand ginst10424 (P2_R1131_U485, P2_R1131_U72, P2_U3471);
  nand ginst10425 (P2_R1131_U486, P2_R1131_U484, P2_R1131_U485);
  nand ginst10426 (P2_R1131_U487, P2_R1131_U165, P2_R1131_U166);
  nand ginst10427 (P2_R1131_U488, P2_R1131_U254, P2_R1131_U486);
  nand ginst10428 (P2_R1131_U489, P2_R1131_U69, P2_U3082);
  not ginst10429 (P2_R1131_U49, P2_U3951);
  nand ginst10430 (P2_R1131_U490, P2_R1131_U70, P2_U3468);
  nand ginst10431 (P2_R1131_U491, P2_R1131_U64, P2_U3074);
  nand ginst10432 (P2_R1131_U492, P2_R1131_U65, P2_U3465);
  nand ginst10433 (P2_R1131_U493, P2_R1131_U491, P2_R1131_U492);
  nand ginst10434 (P2_R1131_U494, P2_R1131_U362, P2_R1131_U93);
  nand ginst10435 (P2_R1131_U495, P2_R1131_U338, P2_R1131_U493);
  nand ginst10436 (P2_R1131_U496, P2_R1131_U66, P2_U3065);
  nand ginst10437 (P2_R1131_U497, P2_R1131_U67, P2_U3462);
  nand ginst10438 (P2_R1131_U498, P2_R1131_U496, P2_R1131_U497);
  nand ginst10439 (P2_R1131_U499, P2_R1131_U167, P2_R1131_U363);
  and ginst10440 (P2_R1131_U5, P2_R1131_U196, P2_R1131_U197);
  not ginst10441 (P2_R1131_U50, P2_U3952);
  nand ginst10442 (P2_R1131_U500, P2_R1131_U244, P2_R1131_U498);
  nand ginst10443 (P2_R1131_U501, P2_R1131_U62, P2_U3064);
  nand ginst10444 (P2_R1131_U502, P2_R1131_U63, P2_U3459);
  nand ginst10445 (P2_R1131_U503, P2_R1131_U29, P2_U3079);
  nand ginst10446 (P2_R1131_U504, P2_R1131_U30, P2_U3427);
  not ginst10447 (P2_R1131_U51, P2_U3060);
  not ginst10448 (P2_R1131_U52, P2_U3953);
  not ginst10449 (P2_R1131_U53, P2_U3067);
  not ginst10450 (P2_R1131_U54, P2_U3956);
  not ginst10451 (P2_R1131_U55, P2_U3077);
  not ginst10452 (P2_R1131_U56, P2_U3477);
  not ginst10453 (P2_R1131_U57, P2_U3075);
  not ginst10454 (P2_R1131_U58, P2_U3071);
  nand ginst10455 (P2_R1131_U59, P2_U3075, P2_U3477);
  and ginst10456 (P2_R1131_U6, P2_R1131_U236, P2_R1131_U237);
  not ginst10457 (P2_R1131_U60, P2_U3480);
  nand ginst10458 (P2_R1131_U61, P2_U3086, P2_U3453);
  not ginst10459 (P2_R1131_U62, P2_U3459);
  not ginst10460 (P2_R1131_U63, P2_U3064);
  not ginst10461 (P2_R1131_U64, P2_U3465);
  not ginst10462 (P2_R1131_U65, P2_U3074);
  not ginst10463 (P2_R1131_U66, P2_U3462);
  not ginst10464 (P2_R1131_U67, P2_U3065);
  nand ginst10465 (P2_R1131_U68, P2_U3065, P2_U3462);
  not ginst10466 (P2_R1131_U69, P2_U3468);
  and ginst10467 (P2_R1131_U7, P2_R1131_U245, P2_R1131_U246);
  not ginst10468 (P2_R1131_U70, P2_U3082);
  not ginst10469 (P2_R1131_U71, P2_U3471);
  not ginst10470 (P2_R1131_U72, P2_U3081);
  not ginst10471 (P2_R1131_U73, P2_U3474);
  not ginst10472 (P2_R1131_U74, P2_U3076);
  not ginst10473 (P2_R1131_U75, P2_U3483);
  not ginst10474 (P2_R1131_U76, P2_U3084);
  nand ginst10475 (P2_R1131_U77, P2_U3084, P2_U3483);
  not ginst10476 (P2_R1131_U78, P2_U3485);
  not ginst10477 (P2_R1131_U79, P2_U3083);
  and ginst10478 (P2_R1131_U8, P2_R1131_U263, P2_R1131_U264);
  nand ginst10479 (P2_R1131_U80, P2_U3083, P2_U3485);
  not ginst10480 (P2_R1131_U81, P2_U3957);
  not ginst10481 (P2_R1131_U82, P2_U3955);
  not ginst10482 (P2_R1131_U83, P2_U3063);
  not ginst10483 (P2_R1131_U84, P2_U3954);
  not ginst10484 (P2_R1131_U85, P2_U3068);
  nand ginst10485 (P2_R1131_U86, P2_U3059, P2_U3951);
  not ginst10486 (P2_R1131_U87, P2_U3056);
  not ginst10487 (P2_R1131_U88, P2_U3949);
  nand ginst10488 (P2_R1131_U89, P2_R1131_U176, P2_R1131_U306);
  and ginst10489 (P2_R1131_U9, P2_R1131_U271, P2_R1131_U272);
  not ginst10490 (P2_R1131_U90, P2_U3078);
  nand ginst10491 (P2_R1131_U91, P2_R1131_U315, P2_R1131_U77);
  nand ginst10492 (P2_R1131_U92, P2_R1131_U260, P2_R1131_U261);
  nand ginst10493 (P2_R1131_U93, P2_R1131_U337, P2_R1131_U68);
  nand ginst10494 (P2_R1131_U94, P2_R1131_U456, P2_R1131_U457);
  nand ginst10495 (P2_R1131_U95, P2_R1131_U503, P2_R1131_U504);
  nand ginst10496 (P2_R1131_U96, P2_R1131_U374, P2_R1131_U375);
  nand ginst10497 (P2_R1131_U97, P2_R1131_U379, P2_R1131_U380);
  nand ginst10498 (P2_R1131_U98, P2_R1131_U386, P2_R1131_U387);
  nand ginst10499 (P2_R1131_U99, P2_R1131_U393, P2_R1131_U394);
  and ginst10500 (P2_R1146_U10, P2_R1146_U182, P2_R1146_U282);
  nand ginst10501 (P2_R1146_U100, P2_R1146_U449, P2_R1146_U450);
  nand ginst10502 (P2_R1146_U101, P2_R1146_U465, P2_R1146_U466);
  nand ginst10503 (P2_R1146_U102, P2_R1146_U470, P2_R1146_U471);
  nand ginst10504 (P2_R1146_U103, P2_R1146_U355, P2_R1146_U356);
  nand ginst10505 (P2_R1146_U104, P2_R1146_U364, P2_R1146_U365);
  nand ginst10506 (P2_R1146_U105, P2_R1146_U371, P2_R1146_U372);
  nand ginst10507 (P2_R1146_U106, P2_R1146_U375, P2_R1146_U376);
  nand ginst10508 (P2_R1146_U107, P2_R1146_U384, P2_R1146_U385);
  nand ginst10509 (P2_R1146_U108, P2_R1146_U403, P2_R1146_U404);
  nand ginst10510 (P2_R1146_U109, P2_R1146_U420, P2_R1146_U421);
  and ginst10511 (P2_R1146_U11, P2_R1146_U283, P2_R1146_U284);
  nand ginst10512 (P2_R1146_U110, P2_R1146_U424, P2_R1146_U425);
  nand ginst10513 (P2_R1146_U111, P2_R1146_U456, P2_R1146_U457);
  nand ginst10514 (P2_R1146_U112, P2_R1146_U460, P2_R1146_U461);
  nand ginst10515 (P2_R1146_U113, P2_R1146_U477, P2_R1146_U478);
  and ginst10516 (P2_R1146_U114, P2_R1146_U184, P2_R1146_U194);
  and ginst10517 (P2_R1146_U115, P2_R1146_U197, P2_R1146_U198);
  and ginst10518 (P2_R1146_U116, P2_R1146_U185, P2_R1146_U200, P2_R1146_U205);
  and ginst10519 (P2_R1146_U117, P2_R1146_U186, P2_R1146_U210);
  and ginst10520 (P2_R1146_U118, P2_R1146_U213, P2_R1146_U214);
  and ginst10521 (P2_R1146_U119, P2_R1146_U357, P2_R1146_U358, P2_R1146_U38);
  nand ginst10522 (P2_R1146_U12, P2_R1146_U344, P2_R1146_U347);
  and ginst10523 (P2_R1146_U120, P2_R1146_U186, P2_R1146_U361);
  and ginst10524 (P2_R1146_U121, P2_R1146_U229, P2_R1146_U6);
  and ginst10525 (P2_R1146_U122, P2_R1146_U185, P2_R1146_U368);
  and ginst10526 (P2_R1146_U123, P2_R1146_U28, P2_R1146_U377, P2_R1146_U378);
  and ginst10527 (P2_R1146_U124, P2_R1146_U184, P2_R1146_U381);
  and ginst10528 (P2_R1146_U125, P2_R1146_U180, P2_R1146_U216, P2_R1146_U239);
  and ginst10529 (P2_R1146_U126, P2_R1146_U261, P2_R1146_U8);
  and ginst10530 (P2_R1146_U127, P2_R1146_U10, P2_R1146_U287);
  and ginst10531 (P2_R1146_U128, P2_R1146_U303, P2_R1146_U304);
  and ginst10532 (P2_R1146_U129, P2_R1146_U311, P2_R1146_U386, P2_R1146_U387);
  nand ginst10533 (P2_R1146_U13, P2_R1146_U333, P2_R1146_U336);
  and ginst10534 (P2_R1146_U130, P2_R1146_U308, P2_R1146_U390);
  nand ginst10535 (P2_R1146_U131, P2_R1146_U391, P2_R1146_U392);
  and ginst10536 (P2_R1146_U132, P2_R1146_U396, P2_R1146_U397, P2_R1146_U83);
  and ginst10537 (P2_R1146_U133, P2_R1146_U183, P2_R1146_U400);
  nand ginst10538 (P2_R1146_U134, P2_R1146_U405, P2_R1146_U406);
  nand ginst10539 (P2_R1146_U135, P2_R1146_U410, P2_R1146_U411);
  and ginst10540 (P2_R1146_U136, P2_R1146_U11, P2_R1146_U324);
  and ginst10541 (P2_R1146_U137, P2_R1146_U182, P2_R1146_U417);
  nand ginst10542 (P2_R1146_U138, P2_R1146_U426, P2_R1146_U427);
  nand ginst10543 (P2_R1146_U139, P2_R1146_U431, P2_R1146_U432);
  nand ginst10544 (P2_R1146_U14, P2_R1146_U322, P2_R1146_U325);
  nand ginst10545 (P2_R1146_U140, P2_R1146_U436, P2_R1146_U437);
  nand ginst10546 (P2_R1146_U141, P2_R1146_U441, P2_R1146_U442);
  nand ginst10547 (P2_R1146_U142, P2_R1146_U446, P2_R1146_U447);
  and ginst10548 (P2_R1146_U143, P2_R1146_U335, P2_R1146_U9);
  and ginst10549 (P2_R1146_U144, P2_R1146_U181, P2_R1146_U453);
  nand ginst10550 (P2_R1146_U145, P2_R1146_U462, P2_R1146_U463);
  nand ginst10551 (P2_R1146_U146, P2_R1146_U467, P2_R1146_U468);
  and ginst10552 (P2_R1146_U147, P2_R1146_U346, P2_R1146_U7);
  and ginst10553 (P2_R1146_U148, P2_R1146_U180, P2_R1146_U474);
  and ginst10554 (P2_R1146_U149, P2_R1146_U353, P2_R1146_U354);
  nand ginst10555 (P2_R1146_U15, P2_R1146_U314, P2_R1146_U316);
  nand ginst10556 (P2_R1146_U150, P2_R1146_U118, P2_R1146_U211);
  and ginst10557 (P2_R1146_U151, P2_R1146_U362, P2_R1146_U363);
  and ginst10558 (P2_R1146_U152, P2_R1146_U369, P2_R1146_U370);
  and ginst10559 (P2_R1146_U153, P2_R1146_U373, P2_R1146_U374);
  nand ginst10560 (P2_R1146_U154, P2_R1146_U115, P2_R1146_U195);
  and ginst10561 (P2_R1146_U155, P2_R1146_U382, P2_R1146_U383);
  not ginst10562 (P2_R1146_U156, P2_U3960);
  not ginst10563 (P2_R1146_U157, P2_U3057);
  and ginst10564 (P2_R1146_U158, P2_R1146_U401, P2_R1146_U402);
  nand ginst10565 (P2_R1146_U159, P2_R1146_U293, P2_R1146_U294);
  nand ginst10566 (P2_R1146_U16, P2_R1146_U312, P2_R1146_U352);
  nand ginst10567 (P2_R1146_U160, P2_R1146_U289, P2_R1146_U290);
  and ginst10568 (P2_R1146_U161, P2_R1146_U418, P2_R1146_U419);
  and ginst10569 (P2_R1146_U162, P2_R1146_U422, P2_R1146_U423);
  nand ginst10570 (P2_R1146_U163, P2_R1146_U279, P2_R1146_U280);
  nand ginst10571 (P2_R1146_U164, P2_R1146_U275, P2_R1146_U276);
  not ginst10572 (P2_R1146_U165, P2_U3432);
  nand ginst10573 (P2_R1146_U166, P2_R1146_U92, P2_U3427);
  nand ginst10574 (P2_R1146_U167, P2_R1146_U271, P2_R1146_U272);
  not ginst10575 (P2_R1146_U168, P2_U3483);
  nand ginst10576 (P2_R1146_U169, P2_R1146_U263, P2_R1146_U264);
  nand ginst10577 (P2_R1146_U17, P2_R1146_U235, P2_R1146_U237);
  and ginst10578 (P2_R1146_U170, P2_R1146_U454, P2_R1146_U455);
  and ginst10579 (P2_R1146_U171, P2_R1146_U458, P2_R1146_U459);
  nand ginst10580 (P2_R1146_U172, P2_R1146_U253, P2_R1146_U254);
  nand ginst10581 (P2_R1146_U173, P2_R1146_U249, P2_R1146_U250);
  nand ginst10582 (P2_R1146_U174, P2_R1146_U245, P2_R1146_U246);
  and ginst10583 (P2_R1146_U175, P2_R1146_U475, P2_R1146_U476);
  nand ginst10584 (P2_R1146_U176, P2_R1146_U165, P2_R1146_U166);
  not ginst10585 (P2_R1146_U177, P2_R1146_U83);
  not ginst10586 (P2_R1146_U178, P2_R1146_U28);
  not ginst10587 (P2_R1146_U179, P2_R1146_U38);
  nand ginst10588 (P2_R1146_U18, P2_R1146_U227, P2_R1146_U230);
  nand ginst10589 (P2_R1146_U180, P2_R1146_U49, P2_U3459);
  nand ginst10590 (P2_R1146_U181, P2_R1146_U59, P2_U3474);
  nand ginst10591 (P2_R1146_U182, P2_R1146_U74, P2_U3955);
  nand ginst10592 (P2_R1146_U183, P2_R1146_U82, P2_U3951);
  nand ginst10593 (P2_R1146_U184, P2_R1146_U27, P2_U3435);
  nand ginst10594 (P2_R1146_U185, P2_R1146_U33, P2_U3444);
  nand ginst10595 (P2_R1146_U186, P2_R1146_U37, P2_U3450);
  not ginst10596 (P2_R1146_U187, P2_R1146_U61);
  not ginst10597 (P2_R1146_U188, P2_R1146_U76);
  not ginst10598 (P2_R1146_U189, P2_R1146_U35);
  nand ginst10599 (P2_R1146_U19, P2_R1146_U219, P2_R1146_U221);
  not ginst10600 (P2_R1146_U190, P2_R1146_U50);
  not ginst10601 (P2_R1146_U191, P2_R1146_U166);
  nand ginst10602 (P2_R1146_U192, P2_R1146_U166, P2_U3080);
  not ginst10603 (P2_R1146_U193, P2_R1146_U44);
  nand ginst10604 (P2_R1146_U194, P2_R1146_U29, P2_U3438);
  nand ginst10605 (P2_R1146_U195, P2_R1146_U114, P2_R1146_U44);
  nand ginst10606 (P2_R1146_U196, P2_R1146_U28, P2_R1146_U29);
  nand ginst10607 (P2_R1146_U197, P2_R1146_U196, P2_R1146_U26);
  nand ginst10608 (P2_R1146_U198, P2_R1146_U178, P2_U3066);
  not ginst10609 (P2_R1146_U199, P2_R1146_U154);
  nand ginst10610 (P2_R1146_U20, P2_R1146_U166, P2_R1146_U350);
  nand ginst10611 (P2_R1146_U200, P2_R1146_U32, P2_U3447);
  nand ginst10612 (P2_R1146_U201, P2_R1146_U30, P2_U3073);
  nand ginst10613 (P2_R1146_U202, P2_R1146_U22, P2_U3069);
  nand ginst10614 (P2_R1146_U203, P2_R1146_U185, P2_R1146_U189);
  nand ginst10615 (P2_R1146_U204, P2_R1146_U203, P2_R1146_U6);
  nand ginst10616 (P2_R1146_U205, P2_R1146_U34, P2_U3441);
  nand ginst10617 (P2_R1146_U206, P2_R1146_U32, P2_U3447);
  nand ginst10618 (P2_R1146_U207, P2_R1146_U116, P2_R1146_U154);
  nand ginst10619 (P2_R1146_U208, P2_R1146_U204, P2_R1146_U206);
  not ginst10620 (P2_R1146_U209, P2_R1146_U42);
  not ginst10621 (P2_R1146_U21, P2_U3450);
  nand ginst10622 (P2_R1146_U210, P2_R1146_U39, P2_U3453);
  nand ginst10623 (P2_R1146_U211, P2_R1146_U117, P2_R1146_U42);
  nand ginst10624 (P2_R1146_U212, P2_R1146_U38, P2_R1146_U39);
  nand ginst10625 (P2_R1146_U213, P2_R1146_U212, P2_R1146_U36);
  nand ginst10626 (P2_R1146_U214, P2_R1146_U179, P2_U3086);
  not ginst10627 (P2_R1146_U215, P2_R1146_U150);
  nand ginst10628 (P2_R1146_U216, P2_R1146_U41, P2_U3456);
  nand ginst10629 (P2_R1146_U217, P2_R1146_U216, P2_R1146_U50);
  nand ginst10630 (P2_R1146_U218, P2_R1146_U209, P2_R1146_U38);
  nand ginst10631 (P2_R1146_U219, P2_R1146_U120, P2_R1146_U218);
  not ginst10632 (P2_R1146_U22, P2_U3444);
  nand ginst10633 (P2_R1146_U220, P2_R1146_U186, P2_R1146_U42);
  nand ginst10634 (P2_R1146_U221, P2_R1146_U119, P2_R1146_U220);
  nand ginst10635 (P2_R1146_U222, P2_R1146_U186, P2_R1146_U38);
  nand ginst10636 (P2_R1146_U223, P2_R1146_U154, P2_R1146_U205);
  not ginst10637 (P2_R1146_U224, P2_R1146_U43);
  nand ginst10638 (P2_R1146_U225, P2_R1146_U22, P2_U3069);
  nand ginst10639 (P2_R1146_U226, P2_R1146_U224, P2_R1146_U225);
  nand ginst10640 (P2_R1146_U227, P2_R1146_U122, P2_R1146_U226);
  nand ginst10641 (P2_R1146_U228, P2_R1146_U185, P2_R1146_U43);
  nand ginst10642 (P2_R1146_U229, P2_R1146_U32, P2_U3447);
  not ginst10643 (P2_R1146_U23, P2_U3435);
  nand ginst10644 (P2_R1146_U230, P2_R1146_U121, P2_R1146_U228);
  nand ginst10645 (P2_R1146_U231, P2_R1146_U22, P2_U3069);
  nand ginst10646 (P2_R1146_U232, P2_R1146_U185, P2_R1146_U231);
  nand ginst10647 (P2_R1146_U233, P2_R1146_U205, P2_R1146_U35);
  nand ginst10648 (P2_R1146_U234, P2_R1146_U193, P2_R1146_U28);
  nand ginst10649 (P2_R1146_U235, P2_R1146_U124, P2_R1146_U234);
  nand ginst10650 (P2_R1146_U236, P2_R1146_U184, P2_R1146_U44);
  nand ginst10651 (P2_R1146_U237, P2_R1146_U123, P2_R1146_U236);
  nand ginst10652 (P2_R1146_U238, P2_R1146_U184, P2_R1146_U28);
  nand ginst10653 (P2_R1146_U239, P2_R1146_U48, P2_U3462);
  not ginst10654 (P2_R1146_U24, P2_U3427);
  nand ginst10655 (P2_R1146_U240, P2_R1146_U47, P2_U3065);
  nand ginst10656 (P2_R1146_U241, P2_R1146_U46, P2_U3064);
  nand ginst10657 (P2_R1146_U242, P2_R1146_U180, P2_R1146_U190);
  nand ginst10658 (P2_R1146_U243, P2_R1146_U242, P2_R1146_U7);
  nand ginst10659 (P2_R1146_U244, P2_R1146_U48, P2_U3462);
  nand ginst10660 (P2_R1146_U245, P2_R1146_U125, P2_R1146_U150);
  nand ginst10661 (P2_R1146_U246, P2_R1146_U243, P2_R1146_U244);
  not ginst10662 (P2_R1146_U247, P2_R1146_U174);
  nand ginst10663 (P2_R1146_U248, P2_R1146_U52, P2_U3465);
  nand ginst10664 (P2_R1146_U249, P2_R1146_U174, P2_R1146_U248);
  not ginst10665 (P2_R1146_U25, P2_U3080);
  nand ginst10666 (P2_R1146_U250, P2_R1146_U51, P2_U3074);
  not ginst10667 (P2_R1146_U251, P2_R1146_U173);
  nand ginst10668 (P2_R1146_U252, P2_R1146_U54, P2_U3468);
  nand ginst10669 (P2_R1146_U253, P2_R1146_U173, P2_R1146_U252);
  nand ginst10670 (P2_R1146_U254, P2_R1146_U53, P2_U3082);
  not ginst10671 (P2_R1146_U255, P2_R1146_U172);
  nand ginst10672 (P2_R1146_U256, P2_R1146_U58, P2_U3477);
  nand ginst10673 (P2_R1146_U257, P2_R1146_U55, P2_U3075);
  nand ginst10674 (P2_R1146_U258, P2_R1146_U56, P2_U3076);
  nand ginst10675 (P2_R1146_U259, P2_R1146_U187, P2_R1146_U8);
  not ginst10676 (P2_R1146_U26, P2_U3438);
  nand ginst10677 (P2_R1146_U260, P2_R1146_U259, P2_R1146_U9);
  nand ginst10678 (P2_R1146_U261, P2_R1146_U60, P2_U3471);
  nand ginst10679 (P2_R1146_U262, P2_R1146_U58, P2_U3477);
  nand ginst10680 (P2_R1146_U263, P2_R1146_U126, P2_R1146_U172);
  nand ginst10681 (P2_R1146_U264, P2_R1146_U260, P2_R1146_U262);
  not ginst10682 (P2_R1146_U265, P2_R1146_U169);
  nand ginst10683 (P2_R1146_U266, P2_R1146_U63, P2_U3480);
  nand ginst10684 (P2_R1146_U267, P2_R1146_U169, P2_R1146_U266);
  nand ginst10685 (P2_R1146_U268, P2_R1146_U62, P2_U3071);
  not ginst10686 (P2_R1146_U269, P2_R1146_U64);
  not ginst10687 (P2_R1146_U27, P2_U3070);
  nand ginst10688 (P2_R1146_U270, P2_R1146_U269, P2_R1146_U65);
  nand ginst10689 (P2_R1146_U271, P2_R1146_U168, P2_R1146_U270);
  nand ginst10690 (P2_R1146_U272, P2_R1146_U64, P2_U3084);
  not ginst10691 (P2_R1146_U273, P2_R1146_U167);
  nand ginst10692 (P2_R1146_U274, P2_R1146_U67, P2_U3485);
  nand ginst10693 (P2_R1146_U275, P2_R1146_U167, P2_R1146_U274);
  nand ginst10694 (P2_R1146_U276, P2_R1146_U66, P2_U3083);
  not ginst10695 (P2_R1146_U277, P2_R1146_U164);
  nand ginst10696 (P2_R1146_U278, P2_R1146_U69, P2_U3957);
  nand ginst10697 (P2_R1146_U279, P2_R1146_U164, P2_R1146_U278);
  nand ginst10698 (P2_R1146_U28, P2_R1146_U23, P2_U3070);
  nand ginst10699 (P2_R1146_U280, P2_R1146_U68, P2_U3078);
  not ginst10700 (P2_R1146_U281, P2_R1146_U163);
  nand ginst10701 (P2_R1146_U282, P2_R1146_U73, P2_U3954);
  nand ginst10702 (P2_R1146_U283, P2_R1146_U70, P2_U3068);
  nand ginst10703 (P2_R1146_U284, P2_R1146_U71, P2_U3063);
  nand ginst10704 (P2_R1146_U285, P2_R1146_U10, P2_R1146_U188);
  nand ginst10705 (P2_R1146_U286, P2_R1146_U11, P2_R1146_U285);
  nand ginst10706 (P2_R1146_U287, P2_R1146_U75, P2_U3956);
  nand ginst10707 (P2_R1146_U288, P2_R1146_U73, P2_U3954);
  nand ginst10708 (P2_R1146_U289, P2_R1146_U127, P2_R1146_U163);
  not ginst10709 (P2_R1146_U29, P2_U3066);
  nand ginst10710 (P2_R1146_U290, P2_R1146_U286, P2_R1146_U288);
  not ginst10711 (P2_R1146_U291, P2_R1146_U160);
  nand ginst10712 (P2_R1146_U292, P2_R1146_U78, P2_U3953);
  nand ginst10713 (P2_R1146_U293, P2_R1146_U160, P2_R1146_U292);
  nand ginst10714 (P2_R1146_U294, P2_R1146_U77, P2_U3067);
  not ginst10715 (P2_R1146_U295, P2_R1146_U159);
  nand ginst10716 (P2_R1146_U296, P2_R1146_U80, P2_U3952);
  nand ginst10717 (P2_R1146_U297, P2_R1146_U159, P2_R1146_U296);
  nand ginst10718 (P2_R1146_U298, P2_R1146_U79, P2_U3060);
  not ginst10719 (P2_R1146_U299, P2_R1146_U88);
  not ginst10720 (P2_R1146_U30, P2_U3447);
  nand ginst10721 (P2_R1146_U300, P2_R1146_U84, P2_U3950);
  nand ginst10722 (P2_R1146_U301, P2_R1146_U183, P2_R1146_U300, P2_R1146_U88);
  nand ginst10723 (P2_R1146_U302, P2_R1146_U83, P2_R1146_U84);
  nand ginst10724 (P2_R1146_U303, P2_R1146_U302, P2_R1146_U81);
  nand ginst10725 (P2_R1146_U304, P2_R1146_U177, P2_U3055);
  not ginst10726 (P2_R1146_U305, P2_R1146_U87);
  nand ginst10727 (P2_R1146_U306, P2_R1146_U85, P2_U3056);
  nand ginst10728 (P2_R1146_U307, P2_R1146_U305, P2_R1146_U306);
  nand ginst10729 (P2_R1146_U308, P2_R1146_U86, P2_U3949);
  nand ginst10730 (P2_R1146_U309, P2_R1146_U86, P2_U3949);
  not ginst10731 (P2_R1146_U31, P2_U3441);
  nand ginst10732 (P2_R1146_U310, P2_R1146_U309, P2_R1146_U87);
  nand ginst10733 (P2_R1146_U311, P2_R1146_U85, P2_U3056);
  nand ginst10734 (P2_R1146_U312, P2_R1146_U129, P2_R1146_U310);
  nand ginst10735 (P2_R1146_U313, P2_R1146_U299, P2_R1146_U83);
  nand ginst10736 (P2_R1146_U314, P2_R1146_U133, P2_R1146_U313);
  nand ginst10737 (P2_R1146_U315, P2_R1146_U183, P2_R1146_U88);
  nand ginst10738 (P2_R1146_U316, P2_R1146_U132, P2_R1146_U315);
  nand ginst10739 (P2_R1146_U317, P2_R1146_U183, P2_R1146_U83);
  nand ginst10740 (P2_R1146_U318, P2_R1146_U163, P2_R1146_U287);
  not ginst10741 (P2_R1146_U319, P2_R1146_U89);
  not ginst10742 (P2_R1146_U32, P2_U3073);
  nand ginst10743 (P2_R1146_U320, P2_R1146_U71, P2_U3063);
  nand ginst10744 (P2_R1146_U321, P2_R1146_U319, P2_R1146_U320);
  nand ginst10745 (P2_R1146_U322, P2_R1146_U137, P2_R1146_U321);
  nand ginst10746 (P2_R1146_U323, P2_R1146_U182, P2_R1146_U89);
  nand ginst10747 (P2_R1146_U324, P2_R1146_U73, P2_U3954);
  nand ginst10748 (P2_R1146_U325, P2_R1146_U136, P2_R1146_U323);
  nand ginst10749 (P2_R1146_U326, P2_R1146_U71, P2_U3063);
  nand ginst10750 (P2_R1146_U327, P2_R1146_U182, P2_R1146_U326);
  nand ginst10751 (P2_R1146_U328, P2_R1146_U287, P2_R1146_U76);
  nand ginst10752 (P2_R1146_U329, P2_R1146_U172, P2_R1146_U261);
  not ginst10753 (P2_R1146_U33, P2_U3069);
  not ginst10754 (P2_R1146_U330, P2_R1146_U90);
  nand ginst10755 (P2_R1146_U331, P2_R1146_U56, P2_U3076);
  nand ginst10756 (P2_R1146_U332, P2_R1146_U330, P2_R1146_U331);
  nand ginst10757 (P2_R1146_U333, P2_R1146_U144, P2_R1146_U332);
  nand ginst10758 (P2_R1146_U334, P2_R1146_U181, P2_R1146_U90);
  nand ginst10759 (P2_R1146_U335, P2_R1146_U58, P2_U3477);
  nand ginst10760 (P2_R1146_U336, P2_R1146_U143, P2_R1146_U334);
  nand ginst10761 (P2_R1146_U337, P2_R1146_U56, P2_U3076);
  nand ginst10762 (P2_R1146_U338, P2_R1146_U181, P2_R1146_U337);
  nand ginst10763 (P2_R1146_U339, P2_R1146_U261, P2_R1146_U61);
  not ginst10764 (P2_R1146_U34, P2_U3062);
  nand ginst10765 (P2_R1146_U340, P2_R1146_U150, P2_R1146_U216);
  not ginst10766 (P2_R1146_U341, P2_R1146_U91);
  nand ginst10767 (P2_R1146_U342, P2_R1146_U46, P2_U3064);
  nand ginst10768 (P2_R1146_U343, P2_R1146_U341, P2_R1146_U342);
  nand ginst10769 (P2_R1146_U344, P2_R1146_U148, P2_R1146_U343);
  nand ginst10770 (P2_R1146_U345, P2_R1146_U180, P2_R1146_U91);
  nand ginst10771 (P2_R1146_U346, P2_R1146_U48, P2_U3462);
  nand ginst10772 (P2_R1146_U347, P2_R1146_U147, P2_R1146_U345);
  nand ginst10773 (P2_R1146_U348, P2_R1146_U46, P2_U3064);
  nand ginst10774 (P2_R1146_U349, P2_R1146_U180, P2_R1146_U348);
  nand ginst10775 (P2_R1146_U35, P2_R1146_U31, P2_U3062);
  nand ginst10776 (P2_R1146_U350, P2_R1146_U24, P2_U3079);
  nand ginst10777 (P2_R1146_U351, P2_R1146_U165, P2_U3080);
  nand ginst10778 (P2_R1146_U352, P2_R1146_U130, P2_R1146_U307);
  nand ginst10779 (P2_R1146_U353, P2_R1146_U41, P2_U3456);
  nand ginst10780 (P2_R1146_U354, P2_R1146_U40, P2_U3085);
  nand ginst10781 (P2_R1146_U355, P2_R1146_U150, P2_R1146_U217);
  nand ginst10782 (P2_R1146_U356, P2_R1146_U149, P2_R1146_U215);
  nand ginst10783 (P2_R1146_U357, P2_R1146_U39, P2_U3453);
  nand ginst10784 (P2_R1146_U358, P2_R1146_U36, P2_U3086);
  nand ginst10785 (P2_R1146_U359, P2_R1146_U39, P2_U3453);
  not ginst10786 (P2_R1146_U36, P2_U3453);
  nand ginst10787 (P2_R1146_U360, P2_R1146_U36, P2_U3086);
  nand ginst10788 (P2_R1146_U361, P2_R1146_U359, P2_R1146_U360);
  nand ginst10789 (P2_R1146_U362, P2_R1146_U37, P2_U3450);
  nand ginst10790 (P2_R1146_U363, P2_R1146_U21, P2_U3072);
  nand ginst10791 (P2_R1146_U364, P2_R1146_U222, P2_R1146_U42);
  nand ginst10792 (P2_R1146_U365, P2_R1146_U151, P2_R1146_U209);
  nand ginst10793 (P2_R1146_U366, P2_R1146_U32, P2_U3447);
  nand ginst10794 (P2_R1146_U367, P2_R1146_U30, P2_U3073);
  nand ginst10795 (P2_R1146_U368, P2_R1146_U366, P2_R1146_U367);
  nand ginst10796 (P2_R1146_U369, P2_R1146_U33, P2_U3444);
  not ginst10797 (P2_R1146_U37, P2_U3072);
  nand ginst10798 (P2_R1146_U370, P2_R1146_U22, P2_U3069);
  nand ginst10799 (P2_R1146_U371, P2_R1146_U232, P2_R1146_U43);
  nand ginst10800 (P2_R1146_U372, P2_R1146_U152, P2_R1146_U224);
  nand ginst10801 (P2_R1146_U373, P2_R1146_U34, P2_U3441);
  nand ginst10802 (P2_R1146_U374, P2_R1146_U31, P2_U3062);
  nand ginst10803 (P2_R1146_U375, P2_R1146_U154, P2_R1146_U233);
  nand ginst10804 (P2_R1146_U376, P2_R1146_U153, P2_R1146_U199);
  nand ginst10805 (P2_R1146_U377, P2_R1146_U29, P2_U3438);
  nand ginst10806 (P2_R1146_U378, P2_R1146_U26, P2_U3066);
  nand ginst10807 (P2_R1146_U379, P2_R1146_U29, P2_U3438);
  nand ginst10808 (P2_R1146_U38, P2_R1146_U21, P2_U3072);
  nand ginst10809 (P2_R1146_U380, P2_R1146_U26, P2_U3066);
  nand ginst10810 (P2_R1146_U381, P2_R1146_U379, P2_R1146_U380);
  nand ginst10811 (P2_R1146_U382, P2_R1146_U27, P2_U3435);
  nand ginst10812 (P2_R1146_U383, P2_R1146_U23, P2_U3070);
  nand ginst10813 (P2_R1146_U384, P2_R1146_U238, P2_R1146_U44);
  nand ginst10814 (P2_R1146_U385, P2_R1146_U155, P2_R1146_U193);
  nand ginst10815 (P2_R1146_U386, P2_R1146_U157, P2_U3960);
  nand ginst10816 (P2_R1146_U387, P2_R1146_U156, P2_U3057);
  nand ginst10817 (P2_R1146_U388, P2_R1146_U157, P2_U3960);
  nand ginst10818 (P2_R1146_U389, P2_R1146_U156, P2_U3057);
  not ginst10819 (P2_R1146_U39, P2_U3086);
  nand ginst10820 (P2_R1146_U390, P2_R1146_U388, P2_R1146_U389);
  nand ginst10821 (P2_R1146_U391, P2_R1146_U86, P2_U3949);
  nand ginst10822 (P2_R1146_U392, P2_R1146_U85, P2_U3056);
  not ginst10823 (P2_R1146_U393, P2_R1146_U131);
  nand ginst10824 (P2_R1146_U394, P2_R1146_U305, P2_R1146_U393);
  nand ginst10825 (P2_R1146_U395, P2_R1146_U131, P2_R1146_U87);
  nand ginst10826 (P2_R1146_U396, P2_R1146_U84, P2_U3950);
  nand ginst10827 (P2_R1146_U397, P2_R1146_U81, P2_U3055);
  nand ginst10828 (P2_R1146_U398, P2_R1146_U84, P2_U3950);
  nand ginst10829 (P2_R1146_U399, P2_R1146_U81, P2_U3055);
  not ginst10830 (P2_R1146_U40, P2_U3456);
  nand ginst10831 (P2_R1146_U400, P2_R1146_U398, P2_R1146_U399);
  nand ginst10832 (P2_R1146_U401, P2_R1146_U82, P2_U3951);
  nand ginst10833 (P2_R1146_U402, P2_R1146_U45, P2_U3059);
  nand ginst10834 (P2_R1146_U403, P2_R1146_U317, P2_R1146_U88);
  nand ginst10835 (P2_R1146_U404, P2_R1146_U158, P2_R1146_U299);
  nand ginst10836 (P2_R1146_U405, P2_R1146_U80, P2_U3952);
  nand ginst10837 (P2_R1146_U406, P2_R1146_U79, P2_U3060);
  not ginst10838 (P2_R1146_U407, P2_R1146_U134);
  nand ginst10839 (P2_R1146_U408, P2_R1146_U295, P2_R1146_U407);
  nand ginst10840 (P2_R1146_U409, P2_R1146_U134, P2_R1146_U159);
  not ginst10841 (P2_R1146_U41, P2_U3085);
  nand ginst10842 (P2_R1146_U410, P2_R1146_U78, P2_U3953);
  nand ginst10843 (P2_R1146_U411, P2_R1146_U77, P2_U3067);
  not ginst10844 (P2_R1146_U412, P2_R1146_U135);
  nand ginst10845 (P2_R1146_U413, P2_R1146_U291, P2_R1146_U412);
  nand ginst10846 (P2_R1146_U414, P2_R1146_U135, P2_R1146_U160);
  nand ginst10847 (P2_R1146_U415, P2_R1146_U73, P2_U3954);
  nand ginst10848 (P2_R1146_U416, P2_R1146_U70, P2_U3068);
  nand ginst10849 (P2_R1146_U417, P2_R1146_U415, P2_R1146_U416);
  nand ginst10850 (P2_R1146_U418, P2_R1146_U74, P2_U3955);
  nand ginst10851 (P2_R1146_U419, P2_R1146_U71, P2_U3063);
  nand ginst10852 (P2_R1146_U42, P2_R1146_U207, P2_R1146_U208);
  nand ginst10853 (P2_R1146_U420, P2_R1146_U327, P2_R1146_U89);
  nand ginst10854 (P2_R1146_U421, P2_R1146_U161, P2_R1146_U319);
  nand ginst10855 (P2_R1146_U422, P2_R1146_U75, P2_U3956);
  nand ginst10856 (P2_R1146_U423, P2_R1146_U72, P2_U3077);
  nand ginst10857 (P2_R1146_U424, P2_R1146_U163, P2_R1146_U328);
  nand ginst10858 (P2_R1146_U425, P2_R1146_U162, P2_R1146_U281);
  nand ginst10859 (P2_R1146_U426, P2_R1146_U69, P2_U3957);
  nand ginst10860 (P2_R1146_U427, P2_R1146_U68, P2_U3078);
  not ginst10861 (P2_R1146_U428, P2_R1146_U138);
  nand ginst10862 (P2_R1146_U429, P2_R1146_U277, P2_R1146_U428);
  nand ginst10863 (P2_R1146_U43, P2_R1146_U223, P2_R1146_U35);
  nand ginst10864 (P2_R1146_U430, P2_R1146_U138, P2_R1146_U164);
  nand ginst10865 (P2_R1146_U431, P2_R1146_U25, P2_U3432);
  nand ginst10866 (P2_R1146_U432, P2_R1146_U165, P2_U3080);
  not ginst10867 (P2_R1146_U433, P2_R1146_U139);
  nand ginst10868 (P2_R1146_U434, P2_R1146_U191, P2_R1146_U433);
  nand ginst10869 (P2_R1146_U435, P2_R1146_U139, P2_R1146_U166);
  nand ginst10870 (P2_R1146_U436, P2_R1146_U67, P2_U3485);
  nand ginst10871 (P2_R1146_U437, P2_R1146_U66, P2_U3083);
  not ginst10872 (P2_R1146_U438, P2_R1146_U140);
  nand ginst10873 (P2_R1146_U439, P2_R1146_U273, P2_R1146_U438);
  nand ginst10874 (P2_R1146_U44, P2_R1146_U176, P2_R1146_U192, P2_R1146_U351);
  nand ginst10875 (P2_R1146_U440, P2_R1146_U140, P2_R1146_U167);
  nand ginst10876 (P2_R1146_U441, P2_R1146_U65, P2_U3483);
  nand ginst10877 (P2_R1146_U442, P2_R1146_U168, P2_U3084);
  not ginst10878 (P2_R1146_U443, P2_R1146_U141);
  nand ginst10879 (P2_R1146_U444, P2_R1146_U269, P2_R1146_U443);
  nand ginst10880 (P2_R1146_U445, P2_R1146_U141, P2_R1146_U64);
  nand ginst10881 (P2_R1146_U446, P2_R1146_U63, P2_U3480);
  nand ginst10882 (P2_R1146_U447, P2_R1146_U62, P2_U3071);
  not ginst10883 (P2_R1146_U448, P2_R1146_U142);
  nand ginst10884 (P2_R1146_U449, P2_R1146_U265, P2_R1146_U448);
  not ginst10885 (P2_R1146_U45, P2_U3951);
  nand ginst10886 (P2_R1146_U450, P2_R1146_U142, P2_R1146_U169);
  nand ginst10887 (P2_R1146_U451, P2_R1146_U58, P2_U3477);
  nand ginst10888 (P2_R1146_U452, P2_R1146_U55, P2_U3075);
  nand ginst10889 (P2_R1146_U453, P2_R1146_U451, P2_R1146_U452);
  nand ginst10890 (P2_R1146_U454, P2_R1146_U59, P2_U3474);
  nand ginst10891 (P2_R1146_U455, P2_R1146_U56, P2_U3076);
  nand ginst10892 (P2_R1146_U456, P2_R1146_U338, P2_R1146_U90);
  nand ginst10893 (P2_R1146_U457, P2_R1146_U170, P2_R1146_U330);
  nand ginst10894 (P2_R1146_U458, P2_R1146_U60, P2_U3471);
  nand ginst10895 (P2_R1146_U459, P2_R1146_U57, P2_U3081);
  not ginst10896 (P2_R1146_U46, P2_U3459);
  nand ginst10897 (P2_R1146_U460, P2_R1146_U172, P2_R1146_U339);
  nand ginst10898 (P2_R1146_U461, P2_R1146_U171, P2_R1146_U255);
  nand ginst10899 (P2_R1146_U462, P2_R1146_U54, P2_U3468);
  nand ginst10900 (P2_R1146_U463, P2_R1146_U53, P2_U3082);
  not ginst10901 (P2_R1146_U464, P2_R1146_U145);
  nand ginst10902 (P2_R1146_U465, P2_R1146_U251, P2_R1146_U464);
  nand ginst10903 (P2_R1146_U466, P2_R1146_U145, P2_R1146_U173);
  nand ginst10904 (P2_R1146_U467, P2_R1146_U52, P2_U3465);
  nand ginst10905 (P2_R1146_U468, P2_R1146_U51, P2_U3074);
  not ginst10906 (P2_R1146_U469, P2_R1146_U146);
  not ginst10907 (P2_R1146_U47, P2_U3462);
  nand ginst10908 (P2_R1146_U470, P2_R1146_U247, P2_R1146_U469);
  nand ginst10909 (P2_R1146_U471, P2_R1146_U146, P2_R1146_U174);
  nand ginst10910 (P2_R1146_U472, P2_R1146_U48, P2_U3462);
  nand ginst10911 (P2_R1146_U473, P2_R1146_U47, P2_U3065);
  nand ginst10912 (P2_R1146_U474, P2_R1146_U472, P2_R1146_U473);
  nand ginst10913 (P2_R1146_U475, P2_R1146_U49, P2_U3459);
  nand ginst10914 (P2_R1146_U476, P2_R1146_U46, P2_U3064);
  nand ginst10915 (P2_R1146_U477, P2_R1146_U349, P2_R1146_U91);
  nand ginst10916 (P2_R1146_U478, P2_R1146_U175, P2_R1146_U341);
  not ginst10917 (P2_R1146_U48, P2_U3065);
  not ginst10918 (P2_R1146_U49, P2_U3064);
  nand ginst10919 (P2_R1146_U50, P2_R1146_U40, P2_U3085);
  not ginst10920 (P2_R1146_U51, P2_U3465);
  not ginst10921 (P2_R1146_U52, P2_U3074);
  not ginst10922 (P2_R1146_U53, P2_U3468);
  not ginst10923 (P2_R1146_U54, P2_U3082);
  not ginst10924 (P2_R1146_U55, P2_U3477);
  not ginst10925 (P2_R1146_U56, P2_U3474);
  not ginst10926 (P2_R1146_U57, P2_U3471);
  not ginst10927 (P2_R1146_U58, P2_U3075);
  not ginst10928 (P2_R1146_U59, P2_U3076);
  and ginst10929 (P2_R1146_U6, P2_R1146_U201, P2_R1146_U202);
  not ginst10930 (P2_R1146_U60, P2_U3081);
  nand ginst10931 (P2_R1146_U61, P2_R1146_U57, P2_U3081);
  not ginst10932 (P2_R1146_U62, P2_U3480);
  not ginst10933 (P2_R1146_U63, P2_U3071);
  nand ginst10934 (P2_R1146_U64, P2_R1146_U267, P2_R1146_U268);
  not ginst10935 (P2_R1146_U65, P2_U3084);
  not ginst10936 (P2_R1146_U66, P2_U3485);
  not ginst10937 (P2_R1146_U67, P2_U3083);
  not ginst10938 (P2_R1146_U68, P2_U3957);
  not ginst10939 (P2_R1146_U69, P2_U3078);
  and ginst10940 (P2_R1146_U7, P2_R1146_U240, P2_R1146_U241);
  not ginst10941 (P2_R1146_U70, P2_U3954);
  not ginst10942 (P2_R1146_U71, P2_U3955);
  not ginst10943 (P2_R1146_U72, P2_U3956);
  not ginst10944 (P2_R1146_U73, P2_U3068);
  not ginst10945 (P2_R1146_U74, P2_U3063);
  not ginst10946 (P2_R1146_U75, P2_U3077);
  nand ginst10947 (P2_R1146_U76, P2_R1146_U72, P2_U3077);
  not ginst10948 (P2_R1146_U77, P2_U3953);
  not ginst10949 (P2_R1146_U78, P2_U3067);
  not ginst10950 (P2_R1146_U79, P2_U3952);
  and ginst10951 (P2_R1146_U8, P2_R1146_U181, P2_R1146_U256);
  not ginst10952 (P2_R1146_U80, P2_U3060);
  not ginst10953 (P2_R1146_U81, P2_U3950);
  not ginst10954 (P2_R1146_U82, P2_U3059);
  nand ginst10955 (P2_R1146_U83, P2_R1146_U45, P2_U3059);
  not ginst10956 (P2_R1146_U84, P2_U3055);
  not ginst10957 (P2_R1146_U85, P2_U3949);
  not ginst10958 (P2_R1146_U86, P2_U3056);
  nand ginst10959 (P2_R1146_U87, P2_R1146_U128, P2_R1146_U301);
  nand ginst10960 (P2_R1146_U88, P2_R1146_U297, P2_R1146_U298);
  nand ginst10961 (P2_R1146_U89, P2_R1146_U318, P2_R1146_U76);
  and ginst10962 (P2_R1146_U9, P2_R1146_U257, P2_R1146_U258);
  nand ginst10963 (P2_R1146_U90, P2_R1146_U329, P2_R1146_U61);
  nand ginst10964 (P2_R1146_U91, P2_R1146_U340, P2_R1146_U50);
  not ginst10965 (P2_R1146_U92, P2_U3079);
  nand ginst10966 (P2_R1146_U93, P2_R1146_U394, P2_R1146_U395);
  nand ginst10967 (P2_R1146_U94, P2_R1146_U408, P2_R1146_U409);
  nand ginst10968 (P2_R1146_U95, P2_R1146_U413, P2_R1146_U414);
  nand ginst10969 (P2_R1146_U96, P2_R1146_U429, P2_R1146_U430);
  nand ginst10970 (P2_R1146_U97, P2_R1146_U434, P2_R1146_U435);
  nand ginst10971 (P2_R1146_U98, P2_R1146_U439, P2_R1146_U440);
  nand ginst10972 (P2_R1146_U99, P2_R1146_U444, P2_R1146_U445);
  and ginst10973 (P2_R1164_U10, P2_R1164_U348, P2_R1164_U351);
  nand ginst10974 (P2_R1164_U100, P2_R1164_U398, P2_R1164_U399);
  nand ginst10975 (P2_R1164_U101, P2_R1164_U407, P2_R1164_U408);
  nand ginst10976 (P2_R1164_U102, P2_R1164_U414, P2_R1164_U415);
  nand ginst10977 (P2_R1164_U103, P2_R1164_U421, P2_R1164_U422);
  nand ginst10978 (P2_R1164_U104, P2_R1164_U428, P2_R1164_U429);
  nand ginst10979 (P2_R1164_U105, P2_R1164_U433, P2_R1164_U434);
  nand ginst10980 (P2_R1164_U106, P2_R1164_U440, P2_R1164_U441);
  nand ginst10981 (P2_R1164_U107, P2_R1164_U447, P2_R1164_U448);
  nand ginst10982 (P2_R1164_U108, P2_R1164_U461, P2_R1164_U462);
  nand ginst10983 (P2_R1164_U109, P2_R1164_U466, P2_R1164_U467);
  and ginst10984 (P2_R1164_U11, P2_R1164_U341, P2_R1164_U344);
  nand ginst10985 (P2_R1164_U110, P2_R1164_U473, P2_R1164_U474);
  nand ginst10986 (P2_R1164_U111, P2_R1164_U480, P2_R1164_U481);
  nand ginst10987 (P2_R1164_U112, P2_R1164_U487, P2_R1164_U488);
  nand ginst10988 (P2_R1164_U113, P2_R1164_U494, P2_R1164_U495);
  nand ginst10989 (P2_R1164_U114, P2_R1164_U499, P2_R1164_U500);
  and ginst10990 (P2_R1164_U115, P2_R1164_U187, P2_R1164_U189);
  and ginst10991 (P2_R1164_U116, P2_R1164_U180, P2_R1164_U4);
  and ginst10992 (P2_R1164_U117, P2_R1164_U192, P2_R1164_U194);
  and ginst10993 (P2_R1164_U118, P2_R1164_U200, P2_R1164_U201);
  and ginst10994 (P2_R1164_U119, P2_R1164_U22, P2_R1164_U381, P2_R1164_U382);
  and ginst10995 (P2_R1164_U12, P2_R1164_U332, P2_R1164_U335);
  and ginst10996 (P2_R1164_U120, P2_R1164_U212, P2_R1164_U5);
  and ginst10997 (P2_R1164_U121, P2_R1164_U180, P2_R1164_U181);
  and ginst10998 (P2_R1164_U122, P2_R1164_U218, P2_R1164_U220);
  and ginst10999 (P2_R1164_U123, P2_R1164_U34, P2_R1164_U388, P2_R1164_U389);
  and ginst11000 (P2_R1164_U124, P2_R1164_U226, P2_R1164_U4);
  and ginst11001 (P2_R1164_U125, P2_R1164_U181, P2_R1164_U234);
  and ginst11002 (P2_R1164_U126, P2_R1164_U204, P2_R1164_U6);
  and ginst11003 (P2_R1164_U127, P2_R1164_U171, P2_R1164_U239);
  and ginst11004 (P2_R1164_U128, P2_R1164_U250, P2_R1164_U7);
  and ginst11005 (P2_R1164_U129, P2_R1164_U172, P2_R1164_U248);
  and ginst11006 (P2_R1164_U13, P2_R1164_U323, P2_R1164_U326);
  and ginst11007 (P2_R1164_U130, P2_R1164_U267, P2_R1164_U268);
  and ginst11008 (P2_R1164_U131, P2_R1164_U282, P2_R1164_U9);
  and ginst11009 (P2_R1164_U132, P2_R1164_U280, P2_R1164_U285);
  and ginst11010 (P2_R1164_U133, P2_R1164_U298, P2_R1164_U301);
  and ginst11011 (P2_R1164_U134, P2_R1164_U302, P2_R1164_U368);
  and ginst11012 (P2_R1164_U135, P2_R1164_U160, P2_R1164_U278);
  and ginst11013 (P2_R1164_U136, P2_R1164_U454, P2_R1164_U455, P2_R1164_U80);
  and ginst11014 (P2_R1164_U137, P2_R1164_U325, P2_R1164_U9);
  and ginst11015 (P2_R1164_U138, P2_R1164_U468, P2_R1164_U469, P2_R1164_U59);
  and ginst11016 (P2_R1164_U139, P2_R1164_U334, P2_R1164_U8);
  and ginst11017 (P2_R1164_U14, P2_R1164_U318, P2_R1164_U320);
  and ginst11018 (P2_R1164_U140, P2_R1164_U172, P2_R1164_U489, P2_R1164_U490);
  and ginst11019 (P2_R1164_U141, P2_R1164_U343, P2_R1164_U7);
  and ginst11020 (P2_R1164_U142, P2_R1164_U171, P2_R1164_U501, P2_R1164_U502);
  and ginst11021 (P2_R1164_U143, P2_R1164_U350, P2_R1164_U6);
  nand ginst11022 (P2_R1164_U144, P2_R1164_U118, P2_R1164_U202);
  nand ginst11023 (P2_R1164_U145, P2_R1164_U217, P2_R1164_U229);
  not ginst11024 (P2_R1164_U146, P2_U3057);
  not ginst11025 (P2_R1164_U147, P2_U3960);
  and ginst11026 (P2_R1164_U148, P2_R1164_U402, P2_R1164_U403);
  nand ginst11027 (P2_R1164_U149, P2_R1164_U169, P2_R1164_U304, P2_R1164_U364);
  and ginst11028 (P2_R1164_U15, P2_R1164_U310, P2_R1164_U313);
  and ginst11029 (P2_R1164_U150, P2_R1164_U409, P2_R1164_U410);
  nand ginst11030 (P2_R1164_U151, P2_R1164_U134, P2_R1164_U369, P2_R1164_U370);
  and ginst11031 (P2_R1164_U152, P2_R1164_U416, P2_R1164_U417);
  nand ginst11032 (P2_R1164_U153, P2_R1164_U299, P2_R1164_U365, P2_R1164_U86);
  and ginst11033 (P2_R1164_U154, P2_R1164_U423, P2_R1164_U424);
  nand ginst11034 (P2_R1164_U155, P2_R1164_U292, P2_R1164_U293);
  and ginst11035 (P2_R1164_U156, P2_R1164_U435, P2_R1164_U436);
  nand ginst11036 (P2_R1164_U157, P2_R1164_U288, P2_R1164_U289);
  and ginst11037 (P2_R1164_U158, P2_R1164_U442, P2_R1164_U443);
  nand ginst11038 (P2_R1164_U159, P2_R1164_U132, P2_R1164_U284);
  and ginst11039 (P2_R1164_U16, P2_R1164_U232, P2_R1164_U235);
  and ginst11040 (P2_R1164_U160, P2_R1164_U449, P2_R1164_U450);
  nand ginst11041 (P2_R1164_U161, P2_R1164_U327, P2_R1164_U43);
  nand ginst11042 (P2_R1164_U162, P2_R1164_U130, P2_R1164_U269);
  and ginst11043 (P2_R1164_U163, P2_R1164_U475, P2_R1164_U476);
  nand ginst11044 (P2_R1164_U164, P2_R1164_U256, P2_R1164_U257);
  and ginst11045 (P2_R1164_U165, P2_R1164_U482, P2_R1164_U483);
  nand ginst11046 (P2_R1164_U166, P2_R1164_U252, P2_R1164_U253);
  nand ginst11047 (P2_R1164_U167, P2_R1164_U242, P2_R1164_U243);
  nand ginst11048 (P2_R1164_U168, P2_R1164_U366, P2_R1164_U367);
  nand ginst11049 (P2_R1164_U169, P2_R1164_U151, P2_U3056);
  and ginst11050 (P2_R1164_U17, P2_R1164_U224, P2_R1164_U227);
  not ginst11051 (P2_R1164_U170, P2_R1164_U34);
  nand ginst11052 (P2_R1164_U171, P2_U3085, P2_U3456);
  nand ginst11053 (P2_R1164_U172, P2_U3074, P2_U3465);
  nand ginst11054 (P2_R1164_U173, P2_U3060, P2_U3952);
  not ginst11055 (P2_R1164_U174, P2_R1164_U68);
  not ginst11056 (P2_R1164_U175, P2_R1164_U77);
  nand ginst11057 (P2_R1164_U176, P2_U3067, P2_U3953);
  not ginst11058 (P2_R1164_U177, P2_R1164_U61);
  or ginst11059 (P2_R1164_U178, P2_U3069, P2_U3444);
  or ginst11060 (P2_R1164_U179, P2_U3062, P2_U3441);
  and ginst11061 (P2_R1164_U18, P2_R1164_U210, P2_R1164_U213);
  or ginst11062 (P2_R1164_U180, P2_U3066, P2_U3438);
  or ginst11063 (P2_R1164_U181, P2_U3070, P2_U3435);
  not ginst11064 (P2_R1164_U182, P2_R1164_U31);
  or ginst11065 (P2_R1164_U183, P2_U3080, P2_U3432);
  not ginst11066 (P2_R1164_U184, P2_R1164_U42);
  not ginst11067 (P2_R1164_U185, P2_R1164_U43);
  nand ginst11068 (P2_R1164_U186, P2_R1164_U42, P2_R1164_U43);
  nand ginst11069 (P2_R1164_U187, P2_U3070, P2_U3435);
  nand ginst11070 (P2_R1164_U188, P2_R1164_U181, P2_R1164_U186);
  nand ginst11071 (P2_R1164_U189, P2_U3066, P2_U3438);
  not ginst11072 (P2_R1164_U19, P2_U3447);
  nand ginst11073 (P2_R1164_U190, P2_R1164_U115, P2_R1164_U188);
  nand ginst11074 (P2_R1164_U191, P2_R1164_U34, P2_R1164_U35);
  nand ginst11075 (P2_R1164_U192, P2_R1164_U191, P2_U3069);
  nand ginst11076 (P2_R1164_U193, P2_R1164_U116, P2_R1164_U190);
  nand ginst11077 (P2_R1164_U194, P2_R1164_U170, P2_U3444);
  not ginst11078 (P2_R1164_U195, P2_R1164_U41);
  or ginst11079 (P2_R1164_U196, P2_U3072, P2_U3450);
  or ginst11080 (P2_R1164_U197, P2_U3073, P2_U3447);
  not ginst11081 (P2_R1164_U198, P2_R1164_U22);
  nand ginst11082 (P2_R1164_U199, P2_R1164_U22, P2_R1164_U23);
  not ginst11083 (P2_R1164_U20, P2_U3073);
  nand ginst11084 (P2_R1164_U200, P2_R1164_U199, P2_U3072);
  nand ginst11085 (P2_R1164_U201, P2_R1164_U198, P2_U3450);
  nand ginst11086 (P2_R1164_U202, P2_R1164_U41, P2_R1164_U5);
  not ginst11087 (P2_R1164_U203, P2_R1164_U144);
  or ginst11088 (P2_R1164_U204, P2_U3086, P2_U3453);
  nand ginst11089 (P2_R1164_U205, P2_R1164_U144, P2_R1164_U204);
  not ginst11090 (P2_R1164_U206, P2_R1164_U40);
  or ginst11091 (P2_R1164_U207, P2_U3085, P2_U3456);
  or ginst11092 (P2_R1164_U208, P2_U3073, P2_U3447);
  nand ginst11093 (P2_R1164_U209, P2_R1164_U208, P2_R1164_U41);
  not ginst11094 (P2_R1164_U21, P2_U3072);
  nand ginst11095 (P2_R1164_U210, P2_R1164_U119, P2_R1164_U209);
  nand ginst11096 (P2_R1164_U211, P2_R1164_U195, P2_R1164_U22);
  nand ginst11097 (P2_R1164_U212, P2_U3072, P2_U3450);
  nand ginst11098 (P2_R1164_U213, P2_R1164_U120, P2_R1164_U211);
  or ginst11099 (P2_R1164_U214, P2_U3073, P2_U3447);
  nand ginst11100 (P2_R1164_U215, P2_R1164_U181, P2_R1164_U185);
  nand ginst11101 (P2_R1164_U216, P2_U3070, P2_U3435);
  not ginst11102 (P2_R1164_U217, P2_R1164_U45);
  nand ginst11103 (P2_R1164_U218, P2_R1164_U121, P2_R1164_U184);
  nand ginst11104 (P2_R1164_U219, P2_R1164_U180, P2_R1164_U45);
  nand ginst11105 (P2_R1164_U22, P2_U3073, P2_U3447);
  nand ginst11106 (P2_R1164_U220, P2_U3066, P2_U3438);
  not ginst11107 (P2_R1164_U221, P2_R1164_U44);
  or ginst11108 (P2_R1164_U222, P2_U3062, P2_U3441);
  nand ginst11109 (P2_R1164_U223, P2_R1164_U222, P2_R1164_U44);
  nand ginst11110 (P2_R1164_U224, P2_R1164_U123, P2_R1164_U223);
  nand ginst11111 (P2_R1164_U225, P2_R1164_U221, P2_R1164_U34);
  nand ginst11112 (P2_R1164_U226, P2_U3069, P2_U3444);
  nand ginst11113 (P2_R1164_U227, P2_R1164_U124, P2_R1164_U225);
  or ginst11114 (P2_R1164_U228, P2_U3062, P2_U3441);
  nand ginst11115 (P2_R1164_U229, P2_R1164_U181, P2_R1164_U184);
  not ginst11116 (P2_R1164_U23, P2_U3450);
  not ginst11117 (P2_R1164_U230, P2_R1164_U145);
  nand ginst11118 (P2_R1164_U231, P2_U3066, P2_U3438);
  nand ginst11119 (P2_R1164_U232, P2_R1164_U400, P2_R1164_U401, P2_R1164_U42, P2_R1164_U43);
  nand ginst11120 (P2_R1164_U233, P2_R1164_U42, P2_R1164_U43);
  nand ginst11121 (P2_R1164_U234, P2_U3070, P2_U3435);
  nand ginst11122 (P2_R1164_U235, P2_R1164_U125, P2_R1164_U233);
  or ginst11123 (P2_R1164_U236, P2_U3085, P2_U3456);
  or ginst11124 (P2_R1164_U237, P2_U3064, P2_U3459);
  nand ginst11125 (P2_R1164_U238, P2_R1164_U177, P2_R1164_U6);
  nand ginst11126 (P2_R1164_U239, P2_U3064, P2_U3459);
  not ginst11127 (P2_R1164_U24, P2_U3441);
  nand ginst11128 (P2_R1164_U240, P2_R1164_U127, P2_R1164_U238);
  or ginst11129 (P2_R1164_U241, P2_U3064, P2_U3459);
  nand ginst11130 (P2_R1164_U242, P2_R1164_U126, P2_R1164_U144);
  nand ginst11131 (P2_R1164_U243, P2_R1164_U240, P2_R1164_U241);
  not ginst11132 (P2_R1164_U244, P2_R1164_U167);
  or ginst11133 (P2_R1164_U245, P2_U3082, P2_U3468);
  or ginst11134 (P2_R1164_U246, P2_U3074, P2_U3465);
  nand ginst11135 (P2_R1164_U247, P2_R1164_U174, P2_R1164_U7);
  nand ginst11136 (P2_R1164_U248, P2_U3082, P2_U3468);
  nand ginst11137 (P2_R1164_U249, P2_R1164_U129, P2_R1164_U247);
  not ginst11138 (P2_R1164_U25, P2_U3062);
  or ginst11139 (P2_R1164_U250, P2_U3065, P2_U3462);
  or ginst11140 (P2_R1164_U251, P2_U3082, P2_U3468);
  nand ginst11141 (P2_R1164_U252, P2_R1164_U128, P2_R1164_U167);
  nand ginst11142 (P2_R1164_U253, P2_R1164_U249, P2_R1164_U251);
  not ginst11143 (P2_R1164_U254, P2_R1164_U166);
  or ginst11144 (P2_R1164_U255, P2_U3081, P2_U3471);
  nand ginst11145 (P2_R1164_U256, P2_R1164_U166, P2_R1164_U255);
  nand ginst11146 (P2_R1164_U257, P2_U3081, P2_U3471);
  not ginst11147 (P2_R1164_U258, P2_R1164_U164);
  or ginst11148 (P2_R1164_U259, P2_U3076, P2_U3474);
  not ginst11149 (P2_R1164_U26, P2_U3069);
  nand ginst11150 (P2_R1164_U260, P2_R1164_U164, P2_R1164_U259);
  nand ginst11151 (P2_R1164_U261, P2_U3076, P2_U3474);
  not ginst11152 (P2_R1164_U262, P2_R1164_U92);
  or ginst11153 (P2_R1164_U263, P2_U3071, P2_U3480);
  or ginst11154 (P2_R1164_U264, P2_U3075, P2_U3477);
  not ginst11155 (P2_R1164_U265, P2_R1164_U59);
  nand ginst11156 (P2_R1164_U266, P2_R1164_U59, P2_R1164_U60);
  nand ginst11157 (P2_R1164_U267, P2_R1164_U266, P2_U3071);
  nand ginst11158 (P2_R1164_U268, P2_R1164_U265, P2_U3480);
  nand ginst11159 (P2_R1164_U269, P2_R1164_U8, P2_R1164_U92);
  not ginst11160 (P2_R1164_U27, P2_U3435);
  not ginst11161 (P2_R1164_U270, P2_R1164_U162);
  or ginst11162 (P2_R1164_U271, P2_U3078, P2_U3957);
  or ginst11163 (P2_R1164_U272, P2_U3083, P2_U3485);
  or ginst11164 (P2_R1164_U273, P2_U3077, P2_U3956);
  not ginst11165 (P2_R1164_U274, P2_R1164_U80);
  nand ginst11166 (P2_R1164_U275, P2_R1164_U274, P2_U3957);
  nand ginst11167 (P2_R1164_U276, P2_R1164_U275, P2_R1164_U90);
  nand ginst11168 (P2_R1164_U277, P2_R1164_U80, P2_R1164_U81);
  nand ginst11169 (P2_R1164_U278, P2_R1164_U276, P2_R1164_U277);
  nand ginst11170 (P2_R1164_U279, P2_R1164_U175, P2_R1164_U9);
  not ginst11171 (P2_R1164_U28, P2_U3070);
  nand ginst11172 (P2_R1164_U280, P2_U3077, P2_U3956);
  nand ginst11173 (P2_R1164_U281, P2_R1164_U278, P2_R1164_U279);
  or ginst11174 (P2_R1164_U282, P2_U3084, P2_U3483);
  or ginst11175 (P2_R1164_U283, P2_U3077, P2_U3956);
  nand ginst11176 (P2_R1164_U284, P2_R1164_U131, P2_R1164_U162, P2_R1164_U273);
  nand ginst11177 (P2_R1164_U285, P2_R1164_U281, P2_R1164_U283);
  not ginst11178 (P2_R1164_U286, P2_R1164_U159);
  or ginst11179 (P2_R1164_U287, P2_U3063, P2_U3955);
  nand ginst11180 (P2_R1164_U288, P2_R1164_U159, P2_R1164_U287);
  nand ginst11181 (P2_R1164_U289, P2_U3063, P2_U3955);
  not ginst11182 (P2_R1164_U29, P2_U3427);
  not ginst11183 (P2_R1164_U290, P2_R1164_U157);
  or ginst11184 (P2_R1164_U291, P2_U3068, P2_U3954);
  nand ginst11185 (P2_R1164_U292, P2_R1164_U157, P2_R1164_U291);
  nand ginst11186 (P2_R1164_U293, P2_U3068, P2_U3954);
  not ginst11187 (P2_R1164_U294, P2_R1164_U155);
  or ginst11188 (P2_R1164_U295, P2_U3060, P2_U3952);
  nand ginst11189 (P2_R1164_U296, P2_R1164_U173, P2_R1164_U176);
  not ginst11190 (P2_R1164_U297, P2_R1164_U86);
  or ginst11191 (P2_R1164_U298, P2_U3067, P2_U3953);
  nand ginst11192 (P2_R1164_U299, P2_R1164_U155, P2_R1164_U168, P2_R1164_U298);
  not ginst11193 (P2_R1164_U30, P2_U3079);
  not ginst11194 (P2_R1164_U300, P2_R1164_U153);
  or ginst11195 (P2_R1164_U301, P2_U3055, P2_U3950);
  nand ginst11196 (P2_R1164_U302, P2_U3055, P2_U3950);
  not ginst11197 (P2_R1164_U303, P2_R1164_U151);
  nand ginst11198 (P2_R1164_U304, P2_R1164_U151, P2_U3949);
  not ginst11199 (P2_R1164_U305, P2_R1164_U149);
  nand ginst11200 (P2_R1164_U306, P2_R1164_U155, P2_R1164_U298);
  not ginst11201 (P2_R1164_U307, P2_R1164_U89);
  or ginst11202 (P2_R1164_U308, P2_U3060, P2_U3952);
  nand ginst11203 (P2_R1164_U309, P2_R1164_U308, P2_R1164_U89);
  nand ginst11204 (P2_R1164_U31, P2_U3079, P2_U3427);
  nand ginst11205 (P2_R1164_U310, P2_R1164_U154, P2_R1164_U173, P2_R1164_U309);
  nand ginst11206 (P2_R1164_U311, P2_R1164_U173, P2_R1164_U307);
  nand ginst11207 (P2_R1164_U312, P2_U3059, P2_U3951);
  nand ginst11208 (P2_R1164_U313, P2_R1164_U168, P2_R1164_U311, P2_R1164_U312);
  or ginst11209 (P2_R1164_U314, P2_U3060, P2_U3952);
  nand ginst11210 (P2_R1164_U315, P2_R1164_U162, P2_R1164_U282);
  not ginst11211 (P2_R1164_U316, P2_R1164_U91);
  nand ginst11212 (P2_R1164_U317, P2_R1164_U9, P2_R1164_U91);
  nand ginst11213 (P2_R1164_U318, P2_R1164_U135, P2_R1164_U317);
  nand ginst11214 (P2_R1164_U319, P2_R1164_U278, P2_R1164_U317);
  not ginst11215 (P2_R1164_U32, P2_U3438);
  nand ginst11216 (P2_R1164_U320, P2_R1164_U319, P2_R1164_U453);
  or ginst11217 (P2_R1164_U321, P2_U3083, P2_U3485);
  nand ginst11218 (P2_R1164_U322, P2_R1164_U321, P2_R1164_U91);
  nand ginst11219 (P2_R1164_U323, P2_R1164_U136, P2_R1164_U322);
  nand ginst11220 (P2_R1164_U324, P2_R1164_U316, P2_R1164_U80);
  nand ginst11221 (P2_R1164_U325, P2_U3078, P2_U3957);
  nand ginst11222 (P2_R1164_U326, P2_R1164_U137, P2_R1164_U324);
  or ginst11223 (P2_R1164_U327, P2_U3080, P2_U3432);
  not ginst11224 (P2_R1164_U328, P2_R1164_U161);
  or ginst11225 (P2_R1164_U329, P2_U3083, P2_U3485);
  not ginst11226 (P2_R1164_U33, P2_U3066);
  or ginst11227 (P2_R1164_U330, P2_U3075, P2_U3477);
  nand ginst11228 (P2_R1164_U331, P2_R1164_U330, P2_R1164_U92);
  nand ginst11229 (P2_R1164_U332, P2_R1164_U138, P2_R1164_U331);
  nand ginst11230 (P2_R1164_U333, P2_R1164_U262, P2_R1164_U59);
  nand ginst11231 (P2_R1164_U334, P2_U3071, P2_U3480);
  nand ginst11232 (P2_R1164_U335, P2_R1164_U139, P2_R1164_U333);
  or ginst11233 (P2_R1164_U336, P2_U3075, P2_U3477);
  nand ginst11234 (P2_R1164_U337, P2_R1164_U167, P2_R1164_U250);
  not ginst11235 (P2_R1164_U338, P2_R1164_U93);
  or ginst11236 (P2_R1164_U339, P2_U3074, P2_U3465);
  nand ginst11237 (P2_R1164_U34, P2_U3062, P2_U3441);
  nand ginst11238 (P2_R1164_U340, P2_R1164_U339, P2_R1164_U93);
  nand ginst11239 (P2_R1164_U341, P2_R1164_U140, P2_R1164_U340);
  nand ginst11240 (P2_R1164_U342, P2_R1164_U172, P2_R1164_U338);
  nand ginst11241 (P2_R1164_U343, P2_U3082, P2_U3468);
  nand ginst11242 (P2_R1164_U344, P2_R1164_U141, P2_R1164_U342);
  or ginst11243 (P2_R1164_U345, P2_U3074, P2_U3465);
  or ginst11244 (P2_R1164_U346, P2_U3085, P2_U3456);
  nand ginst11245 (P2_R1164_U347, P2_R1164_U346, P2_R1164_U40);
  nand ginst11246 (P2_R1164_U348, P2_R1164_U142, P2_R1164_U347);
  nand ginst11247 (P2_R1164_U349, P2_R1164_U171, P2_R1164_U206);
  not ginst11248 (P2_R1164_U35, P2_U3444);
  nand ginst11249 (P2_R1164_U350, P2_U3064, P2_U3459);
  nand ginst11250 (P2_R1164_U351, P2_R1164_U143, P2_R1164_U349);
  nand ginst11251 (P2_R1164_U352, P2_R1164_U171, P2_R1164_U207);
  nand ginst11252 (P2_R1164_U353, P2_R1164_U204, P2_R1164_U61);
  nand ginst11253 (P2_R1164_U354, P2_R1164_U214, P2_R1164_U22);
  nand ginst11254 (P2_R1164_U355, P2_R1164_U228, P2_R1164_U34);
  nand ginst11255 (P2_R1164_U356, P2_R1164_U180, P2_R1164_U231);
  nand ginst11256 (P2_R1164_U357, P2_R1164_U173, P2_R1164_U314);
  nand ginst11257 (P2_R1164_U358, P2_R1164_U176, P2_R1164_U298);
  nand ginst11258 (P2_R1164_U359, P2_R1164_U329, P2_R1164_U80);
  not ginst11259 (P2_R1164_U36, P2_U3453);
  nand ginst11260 (P2_R1164_U360, P2_R1164_U282, P2_R1164_U77);
  nand ginst11261 (P2_R1164_U361, P2_R1164_U336, P2_R1164_U59);
  nand ginst11262 (P2_R1164_U362, P2_R1164_U172, P2_R1164_U345);
  nand ginst11263 (P2_R1164_U363, P2_R1164_U250, P2_R1164_U68);
  nand ginst11264 (P2_R1164_U364, P2_U3056, P2_U3949);
  nand ginst11265 (P2_R1164_U365, P2_R1164_U168, P2_R1164_U296);
  nand ginst11266 (P2_R1164_U366, P2_R1164_U295, P2_U3059);
  nand ginst11267 (P2_R1164_U367, P2_R1164_U295, P2_U3951);
  nand ginst11268 (P2_R1164_U368, P2_R1164_U168, P2_R1164_U296, P2_R1164_U301);
  nand ginst11269 (P2_R1164_U369, P2_R1164_U133, P2_R1164_U155, P2_R1164_U168);
  not ginst11270 (P2_R1164_U37, P2_U3086);
  nand ginst11271 (P2_R1164_U370, P2_R1164_U297, P2_R1164_U301);
  nand ginst11272 (P2_R1164_U371, P2_R1164_U39, P2_U3085);
  nand ginst11273 (P2_R1164_U372, P2_R1164_U38, P2_U3456);
  nand ginst11274 (P2_R1164_U373, P2_R1164_U371, P2_R1164_U372);
  nand ginst11275 (P2_R1164_U374, P2_R1164_U352, P2_R1164_U40);
  nand ginst11276 (P2_R1164_U375, P2_R1164_U206, P2_R1164_U373);
  nand ginst11277 (P2_R1164_U376, P2_R1164_U36, P2_U3086);
  nand ginst11278 (P2_R1164_U377, P2_R1164_U37, P2_U3453);
  nand ginst11279 (P2_R1164_U378, P2_R1164_U376, P2_R1164_U377);
  nand ginst11280 (P2_R1164_U379, P2_R1164_U144, P2_R1164_U353);
  not ginst11281 (P2_R1164_U38, P2_U3085);
  nand ginst11282 (P2_R1164_U380, P2_R1164_U203, P2_R1164_U378);
  nand ginst11283 (P2_R1164_U381, P2_R1164_U23, P2_U3072);
  nand ginst11284 (P2_R1164_U382, P2_R1164_U21, P2_U3450);
  nand ginst11285 (P2_R1164_U383, P2_R1164_U19, P2_U3073);
  nand ginst11286 (P2_R1164_U384, P2_R1164_U20, P2_U3447);
  nand ginst11287 (P2_R1164_U385, P2_R1164_U383, P2_R1164_U384);
  nand ginst11288 (P2_R1164_U386, P2_R1164_U354, P2_R1164_U41);
  nand ginst11289 (P2_R1164_U387, P2_R1164_U195, P2_R1164_U385);
  nand ginst11290 (P2_R1164_U388, P2_R1164_U35, P2_U3069);
  nand ginst11291 (P2_R1164_U389, P2_R1164_U26, P2_U3444);
  not ginst11292 (P2_R1164_U39, P2_U3456);
  nand ginst11293 (P2_R1164_U390, P2_R1164_U24, P2_U3062);
  nand ginst11294 (P2_R1164_U391, P2_R1164_U25, P2_U3441);
  nand ginst11295 (P2_R1164_U392, P2_R1164_U390, P2_R1164_U391);
  nand ginst11296 (P2_R1164_U393, P2_R1164_U355, P2_R1164_U44);
  nand ginst11297 (P2_R1164_U394, P2_R1164_U221, P2_R1164_U392);
  nand ginst11298 (P2_R1164_U395, P2_R1164_U32, P2_U3066);
  nand ginst11299 (P2_R1164_U396, P2_R1164_U33, P2_U3438);
  nand ginst11300 (P2_R1164_U397, P2_R1164_U395, P2_R1164_U396);
  nand ginst11301 (P2_R1164_U398, P2_R1164_U145, P2_R1164_U356);
  nand ginst11302 (P2_R1164_U399, P2_R1164_U230, P2_R1164_U397);
  and ginst11303 (P2_R1164_U4, P2_R1164_U178, P2_R1164_U179);
  nand ginst11304 (P2_R1164_U40, P2_R1164_U205, P2_R1164_U61);
  nand ginst11305 (P2_R1164_U400, P2_R1164_U27, P2_U3070);
  nand ginst11306 (P2_R1164_U401, P2_R1164_U28, P2_U3435);
  nand ginst11307 (P2_R1164_U402, P2_R1164_U147, P2_U3057);
  nand ginst11308 (P2_R1164_U403, P2_R1164_U146, P2_U3960);
  nand ginst11309 (P2_R1164_U404, P2_R1164_U147, P2_U3057);
  nand ginst11310 (P2_R1164_U405, P2_R1164_U146, P2_U3960);
  nand ginst11311 (P2_R1164_U406, P2_R1164_U404, P2_R1164_U405);
  nand ginst11312 (P2_R1164_U407, P2_R1164_U148, P2_R1164_U149);
  nand ginst11313 (P2_R1164_U408, P2_R1164_U305, P2_R1164_U406);
  nand ginst11314 (P2_R1164_U409, P2_R1164_U88, P2_U3056);
  nand ginst11315 (P2_R1164_U41, P2_R1164_U117, P2_R1164_U193);
  nand ginst11316 (P2_R1164_U410, P2_R1164_U87, P2_U3949);
  nand ginst11317 (P2_R1164_U411, P2_R1164_U88, P2_U3056);
  nand ginst11318 (P2_R1164_U412, P2_R1164_U87, P2_U3949);
  nand ginst11319 (P2_R1164_U413, P2_R1164_U411, P2_R1164_U412);
  nand ginst11320 (P2_R1164_U414, P2_R1164_U150, P2_R1164_U151);
  nand ginst11321 (P2_R1164_U415, P2_R1164_U303, P2_R1164_U413);
  nand ginst11322 (P2_R1164_U416, P2_R1164_U46, P2_U3055);
  nand ginst11323 (P2_R1164_U417, P2_R1164_U47, P2_U3950);
  nand ginst11324 (P2_R1164_U418, P2_R1164_U46, P2_U3055);
  nand ginst11325 (P2_R1164_U419, P2_R1164_U47, P2_U3950);
  nand ginst11326 (P2_R1164_U42, P2_R1164_U182, P2_R1164_U183);
  nand ginst11327 (P2_R1164_U420, P2_R1164_U418, P2_R1164_U419);
  nand ginst11328 (P2_R1164_U421, P2_R1164_U152, P2_R1164_U153);
  nand ginst11329 (P2_R1164_U422, P2_R1164_U300, P2_R1164_U420);
  nand ginst11330 (P2_R1164_U423, P2_R1164_U49, P2_U3059);
  nand ginst11331 (P2_R1164_U424, P2_R1164_U48, P2_U3951);
  nand ginst11332 (P2_R1164_U425, P2_R1164_U50, P2_U3060);
  nand ginst11333 (P2_R1164_U426, P2_R1164_U51, P2_U3952);
  nand ginst11334 (P2_R1164_U427, P2_R1164_U425, P2_R1164_U426);
  nand ginst11335 (P2_R1164_U428, P2_R1164_U357, P2_R1164_U89);
  nand ginst11336 (P2_R1164_U429, P2_R1164_U307, P2_R1164_U427);
  nand ginst11337 (P2_R1164_U43, P2_U3080, P2_U3432);
  nand ginst11338 (P2_R1164_U430, P2_R1164_U52, P2_U3067);
  nand ginst11339 (P2_R1164_U431, P2_R1164_U53, P2_U3953);
  nand ginst11340 (P2_R1164_U432, P2_R1164_U430, P2_R1164_U431);
  nand ginst11341 (P2_R1164_U433, P2_R1164_U155, P2_R1164_U358);
  nand ginst11342 (P2_R1164_U434, P2_R1164_U294, P2_R1164_U432);
  nand ginst11343 (P2_R1164_U435, P2_R1164_U84, P2_U3068);
  nand ginst11344 (P2_R1164_U436, P2_R1164_U85, P2_U3954);
  nand ginst11345 (P2_R1164_U437, P2_R1164_U84, P2_U3068);
  nand ginst11346 (P2_R1164_U438, P2_R1164_U85, P2_U3954);
  nand ginst11347 (P2_R1164_U439, P2_R1164_U437, P2_R1164_U438);
  nand ginst11348 (P2_R1164_U44, P2_R1164_U122, P2_R1164_U219);
  nand ginst11349 (P2_R1164_U440, P2_R1164_U156, P2_R1164_U157);
  nand ginst11350 (P2_R1164_U441, P2_R1164_U290, P2_R1164_U439);
  nand ginst11351 (P2_R1164_U442, P2_R1164_U82, P2_U3063);
  nand ginst11352 (P2_R1164_U443, P2_R1164_U83, P2_U3955);
  nand ginst11353 (P2_R1164_U444, P2_R1164_U82, P2_U3063);
  nand ginst11354 (P2_R1164_U445, P2_R1164_U83, P2_U3955);
  nand ginst11355 (P2_R1164_U446, P2_R1164_U444, P2_R1164_U445);
  nand ginst11356 (P2_R1164_U447, P2_R1164_U158, P2_R1164_U159);
  nand ginst11357 (P2_R1164_U448, P2_R1164_U286, P2_R1164_U446);
  nand ginst11358 (P2_R1164_U449, P2_R1164_U54, P2_U3077);
  nand ginst11359 (P2_R1164_U45, P2_R1164_U215, P2_R1164_U216);
  nand ginst11360 (P2_R1164_U450, P2_R1164_U55, P2_U3956);
  nand ginst11361 (P2_R1164_U451, P2_R1164_U54, P2_U3077);
  nand ginst11362 (P2_R1164_U452, P2_R1164_U55, P2_U3956);
  nand ginst11363 (P2_R1164_U453, P2_R1164_U451, P2_R1164_U452);
  nand ginst11364 (P2_R1164_U454, P2_R1164_U81, P2_U3078);
  nand ginst11365 (P2_R1164_U455, P2_R1164_U90, P2_U3957);
  nand ginst11366 (P2_R1164_U456, P2_R1164_U161, P2_R1164_U182);
  nand ginst11367 (P2_R1164_U457, P2_R1164_U31, P2_R1164_U328);
  nand ginst11368 (P2_R1164_U458, P2_R1164_U78, P2_U3083);
  nand ginst11369 (P2_R1164_U459, P2_R1164_U79, P2_U3485);
  not ginst11370 (P2_R1164_U46, P2_U3950);
  nand ginst11371 (P2_R1164_U460, P2_R1164_U458, P2_R1164_U459);
  nand ginst11372 (P2_R1164_U461, P2_R1164_U359, P2_R1164_U91);
  nand ginst11373 (P2_R1164_U462, P2_R1164_U316, P2_R1164_U460);
  nand ginst11374 (P2_R1164_U463, P2_R1164_U75, P2_U3084);
  nand ginst11375 (P2_R1164_U464, P2_R1164_U76, P2_U3483);
  nand ginst11376 (P2_R1164_U465, P2_R1164_U463, P2_R1164_U464);
  nand ginst11377 (P2_R1164_U466, P2_R1164_U162, P2_R1164_U360);
  nand ginst11378 (P2_R1164_U467, P2_R1164_U270, P2_R1164_U465);
  nand ginst11379 (P2_R1164_U468, P2_R1164_U60, P2_U3071);
  nand ginst11380 (P2_R1164_U469, P2_R1164_U58, P2_U3480);
  not ginst11381 (P2_R1164_U47, P2_U3055);
  nand ginst11382 (P2_R1164_U470, P2_R1164_U56, P2_U3075);
  nand ginst11383 (P2_R1164_U471, P2_R1164_U57, P2_U3477);
  nand ginst11384 (P2_R1164_U472, P2_R1164_U470, P2_R1164_U471);
  nand ginst11385 (P2_R1164_U473, P2_R1164_U361, P2_R1164_U92);
  nand ginst11386 (P2_R1164_U474, P2_R1164_U262, P2_R1164_U472);
  nand ginst11387 (P2_R1164_U475, P2_R1164_U73, P2_U3076);
  nand ginst11388 (P2_R1164_U476, P2_R1164_U74, P2_U3474);
  nand ginst11389 (P2_R1164_U477, P2_R1164_U73, P2_U3076);
  nand ginst11390 (P2_R1164_U478, P2_R1164_U74, P2_U3474);
  nand ginst11391 (P2_R1164_U479, P2_R1164_U477, P2_R1164_U478);
  not ginst11392 (P2_R1164_U48, P2_U3059);
  nand ginst11393 (P2_R1164_U480, P2_R1164_U163, P2_R1164_U164);
  nand ginst11394 (P2_R1164_U481, P2_R1164_U258, P2_R1164_U479);
  nand ginst11395 (P2_R1164_U482, P2_R1164_U71, P2_U3081);
  nand ginst11396 (P2_R1164_U483, P2_R1164_U72, P2_U3471);
  nand ginst11397 (P2_R1164_U484, P2_R1164_U71, P2_U3081);
  nand ginst11398 (P2_R1164_U485, P2_R1164_U72, P2_U3471);
  nand ginst11399 (P2_R1164_U486, P2_R1164_U484, P2_R1164_U485);
  nand ginst11400 (P2_R1164_U487, P2_R1164_U165, P2_R1164_U166);
  nand ginst11401 (P2_R1164_U488, P2_R1164_U254, P2_R1164_U486);
  nand ginst11402 (P2_R1164_U489, P2_R1164_U69, P2_U3082);
  not ginst11403 (P2_R1164_U49, P2_U3951);
  nand ginst11404 (P2_R1164_U490, P2_R1164_U70, P2_U3468);
  nand ginst11405 (P2_R1164_U491, P2_R1164_U64, P2_U3074);
  nand ginst11406 (P2_R1164_U492, P2_R1164_U65, P2_U3465);
  nand ginst11407 (P2_R1164_U493, P2_R1164_U491, P2_R1164_U492);
  nand ginst11408 (P2_R1164_U494, P2_R1164_U362, P2_R1164_U93);
  nand ginst11409 (P2_R1164_U495, P2_R1164_U338, P2_R1164_U493);
  nand ginst11410 (P2_R1164_U496, P2_R1164_U66, P2_U3065);
  nand ginst11411 (P2_R1164_U497, P2_R1164_U67, P2_U3462);
  nand ginst11412 (P2_R1164_U498, P2_R1164_U496, P2_R1164_U497);
  nand ginst11413 (P2_R1164_U499, P2_R1164_U167, P2_R1164_U363);
  and ginst11414 (P2_R1164_U5, P2_R1164_U196, P2_R1164_U197);
  not ginst11415 (P2_R1164_U50, P2_U3952);
  nand ginst11416 (P2_R1164_U500, P2_R1164_U244, P2_R1164_U498);
  nand ginst11417 (P2_R1164_U501, P2_R1164_U62, P2_U3064);
  nand ginst11418 (P2_R1164_U502, P2_R1164_U63, P2_U3459);
  nand ginst11419 (P2_R1164_U503, P2_R1164_U29, P2_U3079);
  nand ginst11420 (P2_R1164_U504, P2_R1164_U30, P2_U3427);
  not ginst11421 (P2_R1164_U51, P2_U3060);
  not ginst11422 (P2_R1164_U52, P2_U3953);
  not ginst11423 (P2_R1164_U53, P2_U3067);
  not ginst11424 (P2_R1164_U54, P2_U3956);
  not ginst11425 (P2_R1164_U55, P2_U3077);
  not ginst11426 (P2_R1164_U56, P2_U3477);
  not ginst11427 (P2_R1164_U57, P2_U3075);
  not ginst11428 (P2_R1164_U58, P2_U3071);
  nand ginst11429 (P2_R1164_U59, P2_U3075, P2_U3477);
  and ginst11430 (P2_R1164_U6, P2_R1164_U236, P2_R1164_U237);
  not ginst11431 (P2_R1164_U60, P2_U3480);
  nand ginst11432 (P2_R1164_U61, P2_U3086, P2_U3453);
  not ginst11433 (P2_R1164_U62, P2_U3459);
  not ginst11434 (P2_R1164_U63, P2_U3064);
  not ginst11435 (P2_R1164_U64, P2_U3465);
  not ginst11436 (P2_R1164_U65, P2_U3074);
  not ginst11437 (P2_R1164_U66, P2_U3462);
  not ginst11438 (P2_R1164_U67, P2_U3065);
  nand ginst11439 (P2_R1164_U68, P2_U3065, P2_U3462);
  not ginst11440 (P2_R1164_U69, P2_U3468);
  and ginst11441 (P2_R1164_U7, P2_R1164_U245, P2_R1164_U246);
  not ginst11442 (P2_R1164_U70, P2_U3082);
  not ginst11443 (P2_R1164_U71, P2_U3471);
  not ginst11444 (P2_R1164_U72, P2_U3081);
  not ginst11445 (P2_R1164_U73, P2_U3474);
  not ginst11446 (P2_R1164_U74, P2_U3076);
  not ginst11447 (P2_R1164_U75, P2_U3483);
  not ginst11448 (P2_R1164_U76, P2_U3084);
  nand ginst11449 (P2_R1164_U77, P2_U3084, P2_U3483);
  not ginst11450 (P2_R1164_U78, P2_U3485);
  not ginst11451 (P2_R1164_U79, P2_U3083);
  and ginst11452 (P2_R1164_U8, P2_R1164_U263, P2_R1164_U264);
  nand ginst11453 (P2_R1164_U80, P2_U3083, P2_U3485);
  not ginst11454 (P2_R1164_U81, P2_U3957);
  not ginst11455 (P2_R1164_U82, P2_U3955);
  not ginst11456 (P2_R1164_U83, P2_U3063);
  not ginst11457 (P2_R1164_U84, P2_U3954);
  not ginst11458 (P2_R1164_U85, P2_U3068);
  nand ginst11459 (P2_R1164_U86, P2_U3059, P2_U3951);
  not ginst11460 (P2_R1164_U87, P2_U3056);
  not ginst11461 (P2_R1164_U88, P2_U3949);
  nand ginst11462 (P2_R1164_U89, P2_R1164_U176, P2_R1164_U306);
  and ginst11463 (P2_R1164_U9, P2_R1164_U271, P2_R1164_U272);
  not ginst11464 (P2_R1164_U90, P2_U3078);
  nand ginst11465 (P2_R1164_U91, P2_R1164_U315, P2_R1164_U77);
  nand ginst11466 (P2_R1164_U92, P2_R1164_U260, P2_R1164_U261);
  nand ginst11467 (P2_R1164_U93, P2_R1164_U337, P2_R1164_U68);
  nand ginst11468 (P2_R1164_U94, P2_R1164_U456, P2_R1164_U457);
  nand ginst11469 (P2_R1164_U95, P2_R1164_U503, P2_R1164_U504);
  nand ginst11470 (P2_R1164_U96, P2_R1164_U374, P2_R1164_U375);
  nand ginst11471 (P2_R1164_U97, P2_R1164_U379, P2_R1164_U380);
  nand ginst11472 (P2_R1164_U98, P2_R1164_U386, P2_R1164_U387);
  nand ginst11473 (P2_R1164_U99, P2_R1164_U393, P2_R1164_U394);
  and ginst11474 (P2_R1170_U10, P2_R1170_U215, P2_R1170_U218);
  not ginst11475 (P2_R1170_U100, P2_R1170_U40);
  not ginst11476 (P2_R1170_U101, P2_R1170_U41);
  nand ginst11477 (P2_R1170_U102, P2_R1170_U40, P2_R1170_U41);
  nand ginst11478 (P2_R1170_U103, P2_REG2_REG_2__SCAN_IN, P2_R1170_U96, P2_U3434);
  nand ginst11479 (P2_R1170_U104, P2_R1170_U102, P2_R1170_U5);
  nand ginst11480 (P2_R1170_U105, P2_REG2_REG_3__SCAN_IN, P2_U3437);
  nand ginst11481 (P2_R1170_U106, P2_R1170_U103, P2_R1170_U104, P2_R1170_U105);
  nand ginst11482 (P2_R1170_U107, P2_R1170_U32, P2_R1170_U33);
  nand ginst11483 (P2_R1170_U108, P2_R1170_U107, P2_U3443);
  nand ginst11484 (P2_R1170_U109, P2_R1170_U106, P2_R1170_U4);
  and ginst11485 (P2_R1170_U11, P2_R1170_U208, P2_R1170_U211);
  nand ginst11486 (P2_R1170_U110, P2_REG2_REG_5__SCAN_IN, P2_R1170_U89);
  not ginst11487 (P2_R1170_U111, P2_R1170_U39);
  or ginst11488 (P2_R1170_U112, P2_REG2_REG_7__SCAN_IN, P2_U3449);
  or ginst11489 (P2_R1170_U113, P2_REG2_REG_6__SCAN_IN, P2_U3446);
  not ginst11490 (P2_R1170_U114, P2_R1170_U20);
  nand ginst11491 (P2_R1170_U115, P2_R1170_U20, P2_R1170_U21);
  nand ginst11492 (P2_R1170_U116, P2_R1170_U115, P2_U3449);
  nand ginst11493 (P2_R1170_U117, P2_REG2_REG_7__SCAN_IN, P2_R1170_U114);
  nand ginst11494 (P2_R1170_U118, P2_R1170_U39, P2_R1170_U6);
  not ginst11495 (P2_R1170_U119, P2_R1170_U81);
  and ginst11496 (P2_R1170_U12, P2_R1170_U199, P2_R1170_U202);
  or ginst11497 (P2_R1170_U120, P2_REG2_REG_8__SCAN_IN, P2_U3452);
  nand ginst11498 (P2_R1170_U121, P2_R1170_U120, P2_R1170_U81);
  not ginst11499 (P2_R1170_U122, P2_R1170_U38);
  or ginst11500 (P2_R1170_U123, P2_REG2_REG_9__SCAN_IN, P2_U3455);
  or ginst11501 (P2_R1170_U124, P2_REG2_REG_6__SCAN_IN, P2_U3446);
  nand ginst11502 (P2_R1170_U125, P2_R1170_U124, P2_R1170_U39);
  nand ginst11503 (P2_R1170_U126, P2_R1170_U125, P2_R1170_U20, P2_R1170_U237, P2_R1170_U238);
  nand ginst11504 (P2_R1170_U127, P2_R1170_U111, P2_R1170_U20);
  nand ginst11505 (P2_R1170_U128, P2_REG2_REG_7__SCAN_IN, P2_U3449);
  nand ginst11506 (P2_R1170_U129, P2_R1170_U127, P2_R1170_U128, P2_R1170_U6);
  and ginst11507 (P2_R1170_U13, P2_R1170_U192, P2_R1170_U196);
  or ginst11508 (P2_R1170_U130, P2_REG2_REG_6__SCAN_IN, P2_U3446);
  nand ginst11509 (P2_R1170_U131, P2_R1170_U101, P2_R1170_U97);
  nand ginst11510 (P2_R1170_U132, P2_REG2_REG_2__SCAN_IN, P2_U3434);
  not ginst11511 (P2_R1170_U133, P2_R1170_U43);
  nand ginst11512 (P2_R1170_U134, P2_R1170_U100, P2_R1170_U5);
  nand ginst11513 (P2_R1170_U135, P2_R1170_U43, P2_R1170_U96);
  nand ginst11514 (P2_R1170_U136, P2_REG2_REG_3__SCAN_IN, P2_U3437);
  not ginst11515 (P2_R1170_U137, P2_R1170_U42);
  or ginst11516 (P2_R1170_U138, P2_REG2_REG_4__SCAN_IN, P2_U3440);
  nand ginst11517 (P2_R1170_U139, P2_R1170_U138, P2_R1170_U42);
  and ginst11518 (P2_R1170_U14, P2_R1170_U148, P2_R1170_U151);
  nand ginst11519 (P2_R1170_U140, P2_R1170_U139, P2_R1170_U244, P2_R1170_U245, P2_R1170_U32);
  nand ginst11520 (P2_R1170_U141, P2_R1170_U137, P2_R1170_U32);
  nand ginst11521 (P2_R1170_U142, P2_REG2_REG_5__SCAN_IN, P2_U3443);
  nand ginst11522 (P2_R1170_U143, P2_R1170_U141, P2_R1170_U142, P2_R1170_U4);
  or ginst11523 (P2_R1170_U144, P2_REG2_REG_4__SCAN_IN, P2_U3440);
  nand ginst11524 (P2_R1170_U145, P2_R1170_U100, P2_R1170_U97);
  not ginst11525 (P2_R1170_U146, P2_R1170_U82);
  nand ginst11526 (P2_R1170_U147, P2_REG2_REG_3__SCAN_IN, P2_U3437);
  nand ginst11527 (P2_R1170_U148, P2_R1170_U256, P2_R1170_U257, P2_R1170_U40, P2_R1170_U41);
  nand ginst11528 (P2_R1170_U149, P2_R1170_U40, P2_R1170_U41);
  and ginst11529 (P2_R1170_U15, P2_R1170_U140, P2_R1170_U143);
  nand ginst11530 (P2_R1170_U150, P2_REG2_REG_2__SCAN_IN, P2_U3434);
  nand ginst11531 (P2_R1170_U151, P2_R1170_U149, P2_R1170_U150, P2_R1170_U97);
  or ginst11532 (P2_R1170_U152, P2_REG2_REG_1__SCAN_IN, P2_U3431);
  not ginst11533 (P2_R1170_U153, P2_R1170_U83);
  or ginst11534 (P2_R1170_U154, P2_REG2_REG_9__SCAN_IN, P2_U3455);
  or ginst11535 (P2_R1170_U155, P2_REG2_REG_10__SCAN_IN, P2_U3458);
  nand ginst11536 (P2_R1170_U156, P2_R1170_U7, P2_R1170_U93);
  nand ginst11537 (P2_R1170_U157, P2_REG2_REG_10__SCAN_IN, P2_U3458);
  nand ginst11538 (P2_R1170_U158, P2_R1170_U156, P2_R1170_U157, P2_R1170_U90);
  or ginst11539 (P2_R1170_U159, P2_REG2_REG_10__SCAN_IN, P2_U3458);
  and ginst11540 (P2_R1170_U16, P2_R1170_U126, P2_R1170_U129);
  nand ginst11541 (P2_R1170_U160, P2_R1170_U120, P2_R1170_U7, P2_R1170_U81);
  nand ginst11542 (P2_R1170_U161, P2_R1170_U158, P2_R1170_U159);
  not ginst11543 (P2_R1170_U162, P2_R1170_U88);
  or ginst11544 (P2_R1170_U163, P2_REG2_REG_13__SCAN_IN, P2_U3467);
  or ginst11545 (P2_R1170_U164, P2_REG2_REG_12__SCAN_IN, P2_U3464);
  nand ginst11546 (P2_R1170_U165, P2_R1170_U8, P2_R1170_U92);
  nand ginst11547 (P2_R1170_U166, P2_REG2_REG_13__SCAN_IN, P2_U3467);
  nand ginst11548 (P2_R1170_U167, P2_R1170_U165, P2_R1170_U166, P2_R1170_U91);
  or ginst11549 (P2_R1170_U168, P2_REG2_REG_11__SCAN_IN, P2_U3461);
  or ginst11550 (P2_R1170_U169, P2_REG2_REG_13__SCAN_IN, P2_U3467);
  not ginst11551 (P2_R1170_U17, P2_REG2_REG_6__SCAN_IN);
  nand ginst11552 (P2_R1170_U170, P2_R1170_U168, P2_R1170_U8, P2_R1170_U88);
  nand ginst11553 (P2_R1170_U171, P2_R1170_U167, P2_R1170_U169);
  not ginst11554 (P2_R1170_U172, P2_R1170_U87);
  or ginst11555 (P2_R1170_U173, P2_REG2_REG_14__SCAN_IN, P2_U3470);
  nand ginst11556 (P2_R1170_U174, P2_R1170_U173, P2_R1170_U87);
  nand ginst11557 (P2_R1170_U175, P2_REG2_REG_14__SCAN_IN, P2_U3470);
  not ginst11558 (P2_R1170_U176, P2_R1170_U86);
  or ginst11559 (P2_R1170_U177, P2_REG2_REG_15__SCAN_IN, P2_U3473);
  nand ginst11560 (P2_R1170_U178, P2_R1170_U177, P2_R1170_U86);
  nand ginst11561 (P2_R1170_U179, P2_REG2_REG_15__SCAN_IN, P2_U3473);
  not ginst11562 (P2_R1170_U18, P2_U3446);
  not ginst11563 (P2_R1170_U180, P2_R1170_U66);
  or ginst11564 (P2_R1170_U181, P2_REG2_REG_17__SCAN_IN, P2_U3479);
  or ginst11565 (P2_R1170_U182, P2_REG2_REG_16__SCAN_IN, P2_U3476);
  not ginst11566 (P2_R1170_U183, P2_R1170_U47);
  nand ginst11567 (P2_R1170_U184, P2_R1170_U47, P2_R1170_U48);
  nand ginst11568 (P2_R1170_U185, P2_R1170_U184, P2_U3479);
  nand ginst11569 (P2_R1170_U186, P2_REG2_REG_17__SCAN_IN, P2_R1170_U183);
  nand ginst11570 (P2_R1170_U187, P2_R1170_U66, P2_R1170_U9);
  not ginst11571 (P2_R1170_U188, P2_R1170_U65);
  or ginst11572 (P2_R1170_U189, P2_REG2_REG_18__SCAN_IN, P2_U3482);
  not ginst11573 (P2_R1170_U19, P2_U3449);
  nand ginst11574 (P2_R1170_U190, P2_R1170_U189, P2_R1170_U65);
  nand ginst11575 (P2_R1170_U191, P2_REG2_REG_18__SCAN_IN, P2_U3482);
  nand ginst11576 (P2_R1170_U192, P2_R1170_U190, P2_R1170_U191, P2_R1170_U260, P2_R1170_U261);
  nand ginst11577 (P2_R1170_U193, P2_REG2_REG_18__SCAN_IN, P2_U3482);
  nand ginst11578 (P2_R1170_U194, P2_R1170_U188, P2_R1170_U193);
  or ginst11579 (P2_R1170_U195, P2_REG2_REG_18__SCAN_IN, P2_U3482);
  nand ginst11580 (P2_R1170_U196, P2_R1170_U194, P2_R1170_U195, P2_R1170_U264);
  or ginst11581 (P2_R1170_U197, P2_REG2_REG_16__SCAN_IN, P2_U3476);
  nand ginst11582 (P2_R1170_U198, P2_R1170_U197, P2_R1170_U66);
  nand ginst11583 (P2_R1170_U199, P2_R1170_U198, P2_R1170_U272, P2_R1170_U273, P2_R1170_U47);
  nand ginst11584 (P2_R1170_U20, P2_REG2_REG_6__SCAN_IN, P2_U3446);
  nand ginst11585 (P2_R1170_U200, P2_R1170_U180, P2_R1170_U47);
  nand ginst11586 (P2_R1170_U201, P2_REG2_REG_17__SCAN_IN, P2_U3479);
  nand ginst11587 (P2_R1170_U202, P2_R1170_U200, P2_R1170_U201, P2_R1170_U9);
  or ginst11588 (P2_R1170_U203, P2_REG2_REG_16__SCAN_IN, P2_U3476);
  nand ginst11589 (P2_R1170_U204, P2_R1170_U168, P2_R1170_U88);
  not ginst11590 (P2_R1170_U205, P2_R1170_U67);
  or ginst11591 (P2_R1170_U206, P2_REG2_REG_12__SCAN_IN, P2_U3464);
  nand ginst11592 (P2_R1170_U207, P2_R1170_U206, P2_R1170_U67);
  nand ginst11593 (P2_R1170_U208, P2_R1170_U207, P2_R1170_U293, P2_R1170_U294, P2_R1170_U91);
  nand ginst11594 (P2_R1170_U209, P2_R1170_U205, P2_R1170_U91);
  not ginst11595 (P2_R1170_U21, P2_REG2_REG_7__SCAN_IN);
  nand ginst11596 (P2_R1170_U210, P2_REG2_REG_13__SCAN_IN, P2_U3467);
  nand ginst11597 (P2_R1170_U211, P2_R1170_U209, P2_R1170_U210, P2_R1170_U8);
  or ginst11598 (P2_R1170_U212, P2_REG2_REG_12__SCAN_IN, P2_U3464);
  or ginst11599 (P2_R1170_U213, P2_REG2_REG_9__SCAN_IN, P2_U3455);
  nand ginst11600 (P2_R1170_U214, P2_R1170_U213, P2_R1170_U38);
  nand ginst11601 (P2_R1170_U215, P2_R1170_U214, P2_R1170_U305, P2_R1170_U306, P2_R1170_U90);
  nand ginst11602 (P2_R1170_U216, P2_R1170_U122, P2_R1170_U90);
  nand ginst11603 (P2_R1170_U217, P2_REG2_REG_10__SCAN_IN, P2_U3458);
  nand ginst11604 (P2_R1170_U218, P2_R1170_U216, P2_R1170_U217, P2_R1170_U7);
  nand ginst11605 (P2_R1170_U219, P2_R1170_U123, P2_R1170_U90);
  not ginst11606 (P2_R1170_U22, P2_REG2_REG_4__SCAN_IN);
  nand ginst11607 (P2_R1170_U220, P2_R1170_U120, P2_R1170_U49);
  nand ginst11608 (P2_R1170_U221, P2_R1170_U130, P2_R1170_U20);
  nand ginst11609 (P2_R1170_U222, P2_R1170_U144, P2_R1170_U32);
  nand ginst11610 (P2_R1170_U223, P2_R1170_U147, P2_R1170_U96);
  nand ginst11611 (P2_R1170_U224, P2_R1170_U203, P2_R1170_U47);
  nand ginst11612 (P2_R1170_U225, P2_R1170_U212, P2_R1170_U91);
  nand ginst11613 (P2_R1170_U226, P2_R1170_U168, P2_R1170_U56);
  nand ginst11614 (P2_R1170_U227, P2_R1170_U37, P2_U3455);
  nand ginst11615 (P2_R1170_U228, P2_REG2_REG_9__SCAN_IN, P2_R1170_U36);
  nand ginst11616 (P2_R1170_U229, P2_R1170_U227, P2_R1170_U228);
  not ginst11617 (P2_R1170_U23, P2_U3440);
  nand ginst11618 (P2_R1170_U230, P2_R1170_U219, P2_R1170_U38);
  nand ginst11619 (P2_R1170_U231, P2_R1170_U122, P2_R1170_U229);
  nand ginst11620 (P2_R1170_U232, P2_R1170_U34, P2_U3452);
  nand ginst11621 (P2_R1170_U233, P2_REG2_REG_8__SCAN_IN, P2_R1170_U35);
  nand ginst11622 (P2_R1170_U234, P2_R1170_U232, P2_R1170_U233);
  nand ginst11623 (P2_R1170_U235, P2_R1170_U220, P2_R1170_U81);
  nand ginst11624 (P2_R1170_U236, P2_R1170_U119, P2_R1170_U234);
  nand ginst11625 (P2_R1170_U237, P2_R1170_U21, P2_U3449);
  nand ginst11626 (P2_R1170_U238, P2_REG2_REG_7__SCAN_IN, P2_R1170_U19);
  nand ginst11627 (P2_R1170_U239, P2_R1170_U17, P2_U3446);
  not ginst11628 (P2_R1170_U24, P2_U3443);
  nand ginst11629 (P2_R1170_U240, P2_REG2_REG_6__SCAN_IN, P2_R1170_U18);
  nand ginst11630 (P2_R1170_U241, P2_R1170_U239, P2_R1170_U240);
  nand ginst11631 (P2_R1170_U242, P2_R1170_U221, P2_R1170_U39);
  nand ginst11632 (P2_R1170_U243, P2_R1170_U111, P2_R1170_U241);
  nand ginst11633 (P2_R1170_U244, P2_R1170_U33, P2_U3443);
  nand ginst11634 (P2_R1170_U245, P2_REG2_REG_5__SCAN_IN, P2_R1170_U24);
  nand ginst11635 (P2_R1170_U246, P2_R1170_U22, P2_U3440);
  nand ginst11636 (P2_R1170_U247, P2_REG2_REG_4__SCAN_IN, P2_R1170_U23);
  nand ginst11637 (P2_R1170_U248, P2_R1170_U246, P2_R1170_U247);
  nand ginst11638 (P2_R1170_U249, P2_R1170_U222, P2_R1170_U42);
  not ginst11639 (P2_R1170_U25, P2_REG2_REG_2__SCAN_IN);
  nand ginst11640 (P2_R1170_U250, P2_R1170_U137, P2_R1170_U248);
  nand ginst11641 (P2_R1170_U251, P2_R1170_U30, P2_U3437);
  nand ginst11642 (P2_R1170_U252, P2_REG2_REG_3__SCAN_IN, P2_R1170_U31);
  nand ginst11643 (P2_R1170_U253, P2_R1170_U251, P2_R1170_U252);
  nand ginst11644 (P2_R1170_U254, P2_R1170_U223, P2_R1170_U82);
  nand ginst11645 (P2_R1170_U255, P2_R1170_U146, P2_R1170_U253);
  nand ginst11646 (P2_R1170_U256, P2_R1170_U25, P2_U3434);
  nand ginst11647 (P2_R1170_U257, P2_REG2_REG_2__SCAN_IN, P2_R1170_U26);
  nand ginst11648 (P2_R1170_U258, P2_R1170_U83, P2_R1170_U98);
  nand ginst11649 (P2_R1170_U259, P2_R1170_U153, P2_R1170_U29);
  not ginst11650 (P2_R1170_U26, P2_U3434);
  nand ginst11651 (P2_R1170_U260, P2_R1170_U85, P2_U3424);
  nand ginst11652 (P2_R1170_U261, P2_REG2_REG_19__SCAN_IN, P2_R1170_U84);
  nand ginst11653 (P2_R1170_U262, P2_R1170_U85, P2_U3424);
  nand ginst11654 (P2_R1170_U263, P2_REG2_REG_19__SCAN_IN, P2_R1170_U84);
  nand ginst11655 (P2_R1170_U264, P2_R1170_U262, P2_R1170_U263);
  nand ginst11656 (P2_R1170_U265, P2_R1170_U63, P2_U3482);
  nand ginst11657 (P2_R1170_U266, P2_REG2_REG_18__SCAN_IN, P2_R1170_U64);
  nand ginst11658 (P2_R1170_U267, P2_R1170_U63, P2_U3482);
  nand ginst11659 (P2_R1170_U268, P2_REG2_REG_18__SCAN_IN, P2_R1170_U64);
  nand ginst11660 (P2_R1170_U269, P2_R1170_U267, P2_R1170_U268);
  not ginst11661 (P2_R1170_U27, P2_REG2_REG_0__SCAN_IN);
  nand ginst11662 (P2_R1170_U270, P2_R1170_U265, P2_R1170_U266, P2_R1170_U65);
  nand ginst11663 (P2_R1170_U271, P2_R1170_U188, P2_R1170_U269);
  nand ginst11664 (P2_R1170_U272, P2_R1170_U48, P2_U3479);
  nand ginst11665 (P2_R1170_U273, P2_REG2_REG_17__SCAN_IN, P2_R1170_U46);
  nand ginst11666 (P2_R1170_U274, P2_R1170_U44, P2_U3476);
  nand ginst11667 (P2_R1170_U275, P2_REG2_REG_16__SCAN_IN, P2_R1170_U45);
  nand ginst11668 (P2_R1170_U276, P2_R1170_U274, P2_R1170_U275);
  nand ginst11669 (P2_R1170_U277, P2_R1170_U224, P2_R1170_U66);
  nand ginst11670 (P2_R1170_U278, P2_R1170_U180, P2_R1170_U276);
  nand ginst11671 (P2_R1170_U279, P2_R1170_U61, P2_U3473);
  not ginst11672 (P2_R1170_U28, P2_U3425);
  nand ginst11673 (P2_R1170_U280, P2_REG2_REG_15__SCAN_IN, P2_R1170_U62);
  nand ginst11674 (P2_R1170_U281, P2_R1170_U61, P2_U3473);
  nand ginst11675 (P2_R1170_U282, P2_REG2_REG_15__SCAN_IN, P2_R1170_U62);
  nand ginst11676 (P2_R1170_U283, P2_R1170_U281, P2_R1170_U282);
  nand ginst11677 (P2_R1170_U284, P2_R1170_U279, P2_R1170_U280, P2_R1170_U86);
  nand ginst11678 (P2_R1170_U285, P2_R1170_U176, P2_R1170_U283);
  nand ginst11679 (P2_R1170_U286, P2_R1170_U59, P2_U3470);
  nand ginst11680 (P2_R1170_U287, P2_REG2_REG_14__SCAN_IN, P2_R1170_U60);
  nand ginst11681 (P2_R1170_U288, P2_R1170_U59, P2_U3470);
  nand ginst11682 (P2_R1170_U289, P2_REG2_REG_14__SCAN_IN, P2_R1170_U60);
  nand ginst11683 (P2_R1170_U29, P2_REG2_REG_0__SCAN_IN, P2_U3425);
  nand ginst11684 (P2_R1170_U290, P2_R1170_U288, P2_R1170_U289);
  nand ginst11685 (P2_R1170_U291, P2_R1170_U286, P2_R1170_U287, P2_R1170_U87);
  nand ginst11686 (P2_R1170_U292, P2_R1170_U172, P2_R1170_U290);
  nand ginst11687 (P2_R1170_U293, P2_R1170_U57, P2_U3467);
  nand ginst11688 (P2_R1170_U294, P2_REG2_REG_13__SCAN_IN, P2_R1170_U58);
  nand ginst11689 (P2_R1170_U295, P2_R1170_U52, P2_U3464);
  nand ginst11690 (P2_R1170_U296, P2_REG2_REG_12__SCAN_IN, P2_R1170_U53);
  nand ginst11691 (P2_R1170_U297, P2_R1170_U295, P2_R1170_U296);
  nand ginst11692 (P2_R1170_U298, P2_R1170_U225, P2_R1170_U67);
  nand ginst11693 (P2_R1170_U299, P2_R1170_U205, P2_R1170_U297);
  not ginst11694 (P2_R1170_U30, P2_REG2_REG_3__SCAN_IN);
  nand ginst11695 (P2_R1170_U300, P2_R1170_U54, P2_U3461);
  nand ginst11696 (P2_R1170_U301, P2_REG2_REG_11__SCAN_IN, P2_R1170_U55);
  nand ginst11697 (P2_R1170_U302, P2_R1170_U300, P2_R1170_U301);
  nand ginst11698 (P2_R1170_U303, P2_R1170_U226, P2_R1170_U88);
  nand ginst11699 (P2_R1170_U304, P2_R1170_U162, P2_R1170_U302);
  nand ginst11700 (P2_R1170_U305, P2_R1170_U50, P2_U3458);
  nand ginst11701 (P2_R1170_U306, P2_REG2_REG_10__SCAN_IN, P2_R1170_U51);
  nand ginst11702 (P2_R1170_U307, P2_R1170_U27, P2_U3425);
  nand ginst11703 (P2_R1170_U308, P2_REG2_REG_0__SCAN_IN, P2_R1170_U28);
  not ginst11704 (P2_R1170_U31, P2_U3437);
  nand ginst11705 (P2_R1170_U32, P2_REG2_REG_4__SCAN_IN, P2_U3440);
  not ginst11706 (P2_R1170_U33, P2_REG2_REG_5__SCAN_IN);
  not ginst11707 (P2_R1170_U34, P2_REG2_REG_8__SCAN_IN);
  not ginst11708 (P2_R1170_U35, P2_U3452);
  not ginst11709 (P2_R1170_U36, P2_U3455);
  not ginst11710 (P2_R1170_U37, P2_REG2_REG_9__SCAN_IN);
  nand ginst11711 (P2_R1170_U38, P2_R1170_U121, P2_R1170_U49);
  nand ginst11712 (P2_R1170_U39, P2_R1170_U108, P2_R1170_U109, P2_R1170_U110);
  and ginst11713 (P2_R1170_U4, P2_R1170_U94, P2_R1170_U95);
  nand ginst11714 (P2_R1170_U40, P2_R1170_U98, P2_R1170_U99);
  nand ginst11715 (P2_R1170_U41, P2_REG2_REG_1__SCAN_IN, P2_U3431);
  nand ginst11716 (P2_R1170_U42, P2_R1170_U134, P2_R1170_U135, P2_R1170_U136);
  nand ginst11717 (P2_R1170_U43, P2_R1170_U131, P2_R1170_U132);
  not ginst11718 (P2_R1170_U44, P2_REG2_REG_16__SCAN_IN);
  not ginst11719 (P2_R1170_U45, P2_U3476);
  not ginst11720 (P2_R1170_U46, P2_U3479);
  nand ginst11721 (P2_R1170_U47, P2_REG2_REG_16__SCAN_IN, P2_U3476);
  not ginst11722 (P2_R1170_U48, P2_REG2_REG_17__SCAN_IN);
  nand ginst11723 (P2_R1170_U49, P2_REG2_REG_8__SCAN_IN, P2_U3452);
  and ginst11724 (P2_R1170_U5, P2_R1170_U96, P2_R1170_U97);
  not ginst11725 (P2_R1170_U50, P2_REG2_REG_10__SCAN_IN);
  not ginst11726 (P2_R1170_U51, P2_U3458);
  not ginst11727 (P2_R1170_U52, P2_REG2_REG_12__SCAN_IN);
  not ginst11728 (P2_R1170_U53, P2_U3464);
  not ginst11729 (P2_R1170_U54, P2_REG2_REG_11__SCAN_IN);
  not ginst11730 (P2_R1170_U55, P2_U3461);
  nand ginst11731 (P2_R1170_U56, P2_REG2_REG_11__SCAN_IN, P2_U3461);
  not ginst11732 (P2_R1170_U57, P2_REG2_REG_13__SCAN_IN);
  not ginst11733 (P2_R1170_U58, P2_U3467);
  not ginst11734 (P2_R1170_U59, P2_REG2_REG_14__SCAN_IN);
  and ginst11735 (P2_R1170_U6, P2_R1170_U112, P2_R1170_U113);
  not ginst11736 (P2_R1170_U60, P2_U3470);
  not ginst11737 (P2_R1170_U61, P2_REG2_REG_15__SCAN_IN);
  not ginst11738 (P2_R1170_U62, P2_U3473);
  not ginst11739 (P2_R1170_U63, P2_REG2_REG_18__SCAN_IN);
  not ginst11740 (P2_R1170_U64, P2_U3482);
  nand ginst11741 (P2_R1170_U65, P2_R1170_U185, P2_R1170_U186, P2_R1170_U187);
  nand ginst11742 (P2_R1170_U66, P2_R1170_U178, P2_R1170_U179);
  nand ginst11743 (P2_R1170_U67, P2_R1170_U204, P2_R1170_U56);
  nand ginst11744 (P2_R1170_U68, P2_R1170_U258, P2_R1170_U259);
  nand ginst11745 (P2_R1170_U69, P2_R1170_U307, P2_R1170_U308);
  and ginst11746 (P2_R1170_U7, P2_R1170_U154, P2_R1170_U155);
  nand ginst11747 (P2_R1170_U70, P2_R1170_U230, P2_R1170_U231);
  nand ginst11748 (P2_R1170_U71, P2_R1170_U235, P2_R1170_U236);
  nand ginst11749 (P2_R1170_U72, P2_R1170_U242, P2_R1170_U243);
  nand ginst11750 (P2_R1170_U73, P2_R1170_U249, P2_R1170_U250);
  nand ginst11751 (P2_R1170_U74, P2_R1170_U254, P2_R1170_U255);
  nand ginst11752 (P2_R1170_U75, P2_R1170_U270, P2_R1170_U271);
  nand ginst11753 (P2_R1170_U76, P2_R1170_U277, P2_R1170_U278);
  nand ginst11754 (P2_R1170_U77, P2_R1170_U284, P2_R1170_U285);
  nand ginst11755 (P2_R1170_U78, P2_R1170_U291, P2_R1170_U292);
  nand ginst11756 (P2_R1170_U79, P2_R1170_U298, P2_R1170_U299);
  and ginst11757 (P2_R1170_U8, P2_R1170_U163, P2_R1170_U164);
  nand ginst11758 (P2_R1170_U80, P2_R1170_U303, P2_R1170_U304);
  nand ginst11759 (P2_R1170_U81, P2_R1170_U116, P2_R1170_U117, P2_R1170_U118);
  nand ginst11760 (P2_R1170_U82, P2_R1170_U133, P2_R1170_U145);
  nand ginst11761 (P2_R1170_U83, P2_R1170_U152, P2_R1170_U41);
  not ginst11762 (P2_R1170_U84, P2_U3424);
  not ginst11763 (P2_R1170_U85, P2_REG2_REG_19__SCAN_IN);
  nand ginst11764 (P2_R1170_U86, P2_R1170_U174, P2_R1170_U175);
  nand ginst11765 (P2_R1170_U87, P2_R1170_U170, P2_R1170_U171);
  nand ginst11766 (P2_R1170_U88, P2_R1170_U160, P2_R1170_U161);
  not ginst11767 (P2_R1170_U89, P2_R1170_U32);
  and ginst11768 (P2_R1170_U9, P2_R1170_U181, P2_R1170_U182);
  nand ginst11769 (P2_R1170_U90, P2_REG2_REG_9__SCAN_IN, P2_U3455);
  nand ginst11770 (P2_R1170_U91, P2_REG2_REG_12__SCAN_IN, P2_U3464);
  not ginst11771 (P2_R1170_U92, P2_R1170_U56);
  not ginst11772 (P2_R1170_U93, P2_R1170_U49);
  or ginst11773 (P2_R1170_U94, P2_REG2_REG_5__SCAN_IN, P2_U3443);
  or ginst11774 (P2_R1170_U95, P2_REG2_REG_4__SCAN_IN, P2_U3440);
  or ginst11775 (P2_R1170_U96, P2_REG2_REG_3__SCAN_IN, P2_U3437);
  or ginst11776 (P2_R1170_U97, P2_REG2_REG_2__SCAN_IN, P2_U3434);
  not ginst11777 (P2_R1170_U98, P2_R1170_U29);
  or ginst11778 (P2_R1170_U99, P2_REG2_REG_1__SCAN_IN, P2_U3431);
  and ginst11779 (P2_R1176_U10, P2_R1176_U229, P2_R1176_U5);
  nand ginst11780 (P2_R1176_U100, P2_R1176_U518, P2_R1176_U519);
  nand ginst11781 (P2_R1176_U101, P2_R1176_U525, P2_R1176_U526);
  nand ginst11782 (P2_R1176_U102, P2_R1176_U532, P2_R1176_U533);
  nand ginst11783 (P2_R1176_U103, P2_R1176_U537, P2_R1176_U538);
  nand ginst11784 (P2_R1176_U104, P2_R1176_U544, P2_R1176_U545);
  nand ginst11785 (P2_R1176_U105, P2_R1176_U551, P2_R1176_U552);
  nand ginst11786 (P2_R1176_U106, P2_R1176_U558, P2_R1176_U559);
  nand ginst11787 (P2_R1176_U107, P2_R1176_U565, P2_R1176_U566);
  nand ginst11788 (P2_R1176_U108, P2_R1176_U570, P2_R1176_U571);
  nand ginst11789 (P2_R1176_U109, P2_R1176_U577, P2_R1176_U578);
  and ginst11790 (P2_R1176_U11, P2_R1176_U259, P2_R1176_U9);
  nand ginst11791 (P2_R1176_U110, P2_R1176_U584, P2_R1176_U585);
  nand ginst11792 (P2_R1176_U111, P2_R1176_U591, P2_R1176_U592);
  nand ginst11793 (P2_R1176_U112, P2_R1176_U598, P2_R1176_U599);
  nand ginst11794 (P2_R1176_U113, P2_R1176_U605, P2_R1176_U606);
  nand ginst11795 (P2_R1176_U114, P2_R1176_U610, P2_R1176_U611);
  nand ginst11796 (P2_R1176_U115, P2_R1176_U617, P2_R1176_U618);
  and ginst11797 (P2_R1176_U116, P2_R1176_U223, P2_R1176_U224);
  and ginst11798 (P2_R1176_U117, P2_R1176_U10, P2_R1176_U240);
  and ginst11799 (P2_R1176_U118, P2_R1176_U241, P2_R1176_U372);
  and ginst11800 (P2_R1176_U119, P2_R1176_U29, P2_R1176_U430, P2_R1176_U431);
  and ginst11801 (P2_R1176_U12, P2_R1176_U527, P2_R1176_U528);
  and ginst11802 (P2_R1176_U120, P2_R1176_U247, P2_R1176_U5);
  and ginst11803 (P2_R1176_U121, P2_R1176_U22, P2_R1176_U451, P2_R1176_U452);
  and ginst11804 (P2_R1176_U122, P2_R1176_U254, P2_R1176_U4);
  and ginst11805 (P2_R1176_U123, P2_R1176_U11, P2_R1176_U272);
  and ginst11806 (P2_R1176_U124, P2_R1176_U207, P2_R1176_U266);
  and ginst11807 (P2_R1176_U125, P2_R1176_U273, P2_R1176_U380);
  and ginst11808 (P2_R1176_U126, P2_R1176_U283, P2_R1176_U284);
  and ginst11809 (P2_R1176_U127, P2_R1176_U296, P2_R1176_U8);
  and ginst11810 (P2_R1176_U128, P2_R1176_U208, P2_R1176_U294);
  and ginst11811 (P2_R1176_U129, P2_R1176_U203, P2_R1176_U312);
  and ginst11812 (P2_R1176_U13, P2_R1176_U348, P2_R1176_U351);
  and ginst11813 (P2_R1176_U130, P2_R1176_U318, P2_R1176_U383);
  and ginst11814 (P2_R1176_U131, P2_R1176_U310, P2_R1176_U320);
  and ginst11815 (P2_R1176_U132, P2_R1176_U312, P2_R1176_U320);
  and ginst11816 (P2_R1176_U133, P2_R1176_U319, P2_R1176_U381);
  nand ginst11817 (P2_R1176_U134, P2_R1176_U512, P2_R1176_U513);
  and ginst11818 (P2_R1176_U135, P2_R1176_U38, P2_R1176_U508);
  and ginst11819 (P2_R1176_U136, P2_R1176_U209, P2_R1176_U212);
  and ginst11820 (P2_R1176_U137, P2_R1176_U203, P2_R1176_U325);
  and ginst11821 (P2_R1176_U138, P2_R1176_U12, P2_R1176_U209);
  and ginst11822 (P2_R1176_U139, P2_R1176_U208, P2_R1176_U553, P2_R1176_U554);
  and ginst11823 (P2_R1176_U14, P2_R1176_U339, P2_R1176_U342);
  and ginst11824 (P2_R1176_U140, P2_R1176_U334, P2_R1176_U8);
  and ginst11825 (P2_R1176_U141, P2_R1176_U42, P2_R1176_U579, P2_R1176_U580);
  and ginst11826 (P2_R1176_U142, P2_R1176_U341, P2_R1176_U7);
  and ginst11827 (P2_R1176_U143, P2_R1176_U207, P2_R1176_U600, P2_R1176_U601);
  and ginst11828 (P2_R1176_U144, P2_R1176_U350, P2_R1176_U6);
  nand ginst11829 (P2_R1176_U145, P2_R1176_U619, P2_R1176_U620);
  not ginst11830 (P2_R1176_U146, P2_U3456);
  and ginst11831 (P2_R1176_U147, P2_R1176_U389, P2_R1176_U390);
  not ginst11832 (P2_R1176_U148, P2_U3441);
  not ginst11833 (P2_R1176_U149, P2_U3432);
  and ginst11834 (P2_R1176_U15, P2_R1176_U332, P2_R1176_U335);
  not ginst11835 (P2_R1176_U150, P2_U3427);
  not ginst11836 (P2_R1176_U151, P2_U3438);
  not ginst11837 (P2_R1176_U152, P2_U3435);
  not ginst11838 (P2_R1176_U153, P2_U3444);
  not ginst11839 (P2_R1176_U154, P2_U3450);
  not ginst11840 (P2_R1176_U155, P2_U3447);
  not ginst11841 (P2_R1176_U156, P2_U3453);
  nand ginst11842 (P2_R1176_U157, P2_R1176_U118, P2_R1176_U371);
  and ginst11843 (P2_R1176_U158, P2_R1176_U423, P2_R1176_U424);
  nand ginst11844 (P2_R1176_U159, P2_R1176_U368, P2_R1176_U370);
  and ginst11845 (P2_R1176_U16, P2_R1176_U323, P2_R1176_U326, P2_R1176_U385);
  and ginst11846 (P2_R1176_U160, P2_R1176_U437, P2_R1176_U438);
  nand ginst11847 (P2_R1176_U161, P2_R1176_U205, P2_R1176_U227, P2_R1176_U362);
  and ginst11848 (P2_R1176_U162, P2_R1176_U444, P2_R1176_U445);
  nand ginst11849 (P2_R1176_U163, P2_R1176_U116, P2_R1176_U225);
  not ginst11850 (P2_R1176_U164, P2_U3950);
  not ginst11851 (P2_R1176_U165, P2_U3951);
  not ginst11852 (P2_R1176_U166, P2_U3459);
  not ginst11853 (P2_R1176_U167, P2_U3462);
  not ginst11854 (P2_R1176_U168, P2_U3468);
  not ginst11855 (P2_R1176_U169, P2_U3465);
  and ginst11856 (P2_R1176_U17, P2_R1176_U252, P2_R1176_U255);
  not ginst11857 (P2_R1176_U170, P2_U3471);
  not ginst11858 (P2_R1176_U171, P2_U3474);
  not ginst11859 (P2_R1176_U172, P2_U3480);
  not ginst11860 (P2_R1176_U173, P2_U3477);
  not ginst11861 (P2_R1176_U174, P2_U3483);
  not ginst11862 (P2_R1176_U175, P2_U3956);
  not ginst11863 (P2_R1176_U176, P2_U3957);
  not ginst11864 (P2_R1176_U177, P2_U3485);
  not ginst11865 (P2_R1176_U178, P2_U3955);
  not ginst11866 (P2_R1176_U179, P2_U3954);
  and ginst11867 (P2_R1176_U18, P2_R1176_U245, P2_R1176_U248);
  not ginst11868 (P2_R1176_U180, P2_U3952);
  not ginst11869 (P2_R1176_U181, P2_U3953);
  not ginst11870 (P2_R1176_U182, P2_U3949);
  not ginst11871 (P2_R1176_U183, P2_U3155);
  and ginst11872 (P2_R1176_U184, P2_R1176_U520, P2_R1176_U521);
  nand ginst11873 (P2_R1176_U185, P2_R1176_U314, P2_R1176_U315);
  nand ginst11874 (P2_R1176_U186, P2_R1176_U306, P2_R1176_U307);
  and ginst11875 (P2_R1176_U187, P2_R1176_U539, P2_R1176_U540);
  nand ginst11876 (P2_R1176_U188, P2_R1176_U302, P2_R1176_U303);
  and ginst11877 (P2_R1176_U189, P2_R1176_U546, P2_R1176_U547);
  not ginst11878 (P2_R1176_U19, P2_U3184);
  nand ginst11879 (P2_R1176_U190, P2_R1176_U298, P2_R1176_U299);
  and ginst11880 (P2_R1176_U191, P2_R1176_U560, P2_R1176_U561);
  nand ginst11881 (P2_R1176_U192, P2_R1176_U214, P2_R1176_U26);
  nand ginst11882 (P2_R1176_U193, P2_R1176_U288, P2_R1176_U289);
  and ginst11883 (P2_R1176_U194, P2_R1176_U572, P2_R1176_U573);
  nand ginst11884 (P2_R1176_U195, P2_R1176_U126, P2_R1176_U285);
  and ginst11885 (P2_R1176_U196, P2_R1176_U586, P2_R1176_U587);
  nand ginst11886 (P2_R1176_U197, P2_R1176_U125, P2_R1176_U379);
  and ginst11887 (P2_R1176_U198, P2_R1176_U593, P2_R1176_U594);
  nand ginst11888 (P2_R1176_U199, P2_R1176_U373, P2_R1176_U378);
  not ginst11889 (P2_R1176_U20, P2_U3175);
  nand ginst11890 (P2_R1176_U200, P2_R1176_U260, P2_R1176_U50);
  and ginst11891 (P2_R1176_U201, P2_R1176_U612, P2_R1176_U613);
  nand ginst11892 (P2_R1176_U202, P2_R1176_U204, P2_R1176_U257, P2_R1176_U363);
  nand ginst11893 (P2_R1176_U203, P2_R1176_U376, P2_R1176_U377);
  nand ginst11894 (P2_R1176_U204, P2_R1176_U157, P2_R1176_U64);
  nand ginst11895 (P2_R1176_U205, P2_R1176_U163, P2_R1176_U70);
  not ginst11896 (P2_R1176_U206, P2_R1176_U22);
  nand ginst11897 (P2_R1176_U207, P2_R1176_U84, P2_U3171);
  nand ginst11898 (P2_R1176_U208, P2_R1176_U89, P2_U3163);
  nand ginst11899 (P2_R1176_U209, P2_R1176_U75, P2_U3158);
  not ginst11900 (P2_R1176_U21, P2_U3181);
  not ginst11901 (P2_R1176_U210, P2_R1176_U47);
  not ginst11902 (P2_R1176_U211, P2_R1176_U55);
  nand ginst11903 (P2_R1176_U212, P2_R1176_U76, P2_U3159);
  nand ginst11904 (P2_R1176_U213, P2_R1176_U19, P2_R1176_U402);
  nand ginst11905 (P2_R1176_U214, P2_R1176_U213, P2_U3183);
  not ginst11906 (P2_R1176_U215, P2_R1176_U26);
  not ginst11907 (P2_R1176_U216, P2_R1176_U192);
  nand ginst11908 (P2_R1176_U217, P2_R1176_U24, P2_R1176_U399);
  nand ginst11909 (P2_R1176_U218, P2_R1176_U68, P2_U3182);
  not ginst11910 (P2_R1176_U219, P2_R1176_U36);
  nand ginst11911 (P2_R1176_U22, P2_R1176_U66, P2_U3181);
  nand ginst11912 (P2_R1176_U220, P2_R1176_U23, P2_R1176_U405);
  nand ginst11913 (P2_R1176_U221, P2_R1176_U21, P2_R1176_U408);
  nand ginst11914 (P2_R1176_U222, P2_R1176_U22, P2_R1176_U23);
  nand ginst11915 (P2_R1176_U223, P2_R1176_U222, P2_R1176_U67);
  nand ginst11916 (P2_R1176_U224, P2_R1176_U206, P2_U3180);
  nand ginst11917 (P2_R1176_U225, P2_R1176_U36, P2_R1176_U4);
  not ginst11918 (P2_R1176_U226, P2_R1176_U163);
  nand ginst11919 (P2_R1176_U227, P2_R1176_U163, P2_U3179);
  not ginst11920 (P2_R1176_U228, P2_R1176_U161);
  nand ginst11921 (P2_R1176_U229, P2_R1176_U31, P2_R1176_U411);
  not ginst11922 (P2_R1176_U23, P2_U3180);
  nand ginst11923 (P2_R1176_U230, P2_R1176_U161, P2_R1176_U229);
  not ginst11924 (P2_R1176_U231, P2_R1176_U32);
  not ginst11925 (P2_R1176_U232, P2_R1176_U35);
  nand ginst11926 (P2_R1176_U233, P2_R1176_U30, P2_R1176_U414);
  nand ginst11927 (P2_R1176_U234, P2_R1176_U28, P2_R1176_U417);
  not ginst11928 (P2_R1176_U235, P2_R1176_U29);
  nand ginst11929 (P2_R1176_U236, P2_R1176_U29, P2_R1176_U30);
  nand ginst11930 (P2_R1176_U237, P2_R1176_U236, P2_R1176_U72);
  nand ginst11931 (P2_R1176_U238, P2_R1176_U235, P2_U3176);
  not ginst11932 (P2_R1176_U239, P2_R1176_U159);
  not ginst11933 (P2_R1176_U24, P2_U3182);
  nand ginst11934 (P2_R1176_U240, P2_R1176_U20, P2_R1176_U420);
  nand ginst11935 (P2_R1176_U241, P2_R1176_U65, P2_U3175);
  not ginst11936 (P2_R1176_U242, P2_R1176_U157);
  nand ginst11937 (P2_R1176_U243, P2_R1176_U28, P2_R1176_U417);
  nand ginst11938 (P2_R1176_U244, P2_R1176_U243, P2_R1176_U35);
  nand ginst11939 (P2_R1176_U245, P2_R1176_U119, P2_R1176_U244);
  nand ginst11940 (P2_R1176_U246, P2_R1176_U232, P2_R1176_U29);
  nand ginst11941 (P2_R1176_U247, P2_R1176_U72, P2_U3176);
  nand ginst11942 (P2_R1176_U248, P2_R1176_U120, P2_R1176_U246);
  nand ginst11943 (P2_R1176_U249, P2_R1176_U28, P2_R1176_U417);
  not ginst11944 (P2_R1176_U25, P2_U3183);
  nand ginst11945 (P2_R1176_U250, P2_R1176_U21, P2_R1176_U408);
  nand ginst11946 (P2_R1176_U251, P2_R1176_U250, P2_R1176_U36);
  nand ginst11947 (P2_R1176_U252, P2_R1176_U121, P2_R1176_U251);
  nand ginst11948 (P2_R1176_U253, P2_R1176_U219, P2_R1176_U22);
  nand ginst11949 (P2_R1176_U254, P2_R1176_U67, P2_U3180);
  nand ginst11950 (P2_R1176_U255, P2_R1176_U122, P2_R1176_U253);
  nand ginst11951 (P2_R1176_U256, P2_R1176_U21, P2_R1176_U408);
  nand ginst11952 (P2_R1176_U257, P2_R1176_U157, P2_U3174);
  not ginst11953 (P2_R1176_U258, P2_R1176_U202);
  nand ginst11954 (P2_R1176_U259, P2_R1176_U466, P2_R1176_U49);
  nand ginst11955 (P2_R1176_U26, P2_R1176_U69, P2_U3184);
  nand ginst11956 (P2_R1176_U260, P2_R1176_U202, P2_R1176_U259);
  not ginst11957 (P2_R1176_U261, P2_R1176_U50);
  not ginst11958 (P2_R1176_U262, P2_R1176_U200);
  nand ginst11959 (P2_R1176_U263, P2_R1176_U472, P2_R1176_U48);
  nand ginst11960 (P2_R1176_U264, P2_R1176_U45, P2_R1176_U475);
  nand ginst11961 (P2_R1176_U265, P2_R1176_U210, P2_R1176_U6);
  nand ginst11962 (P2_R1176_U266, P2_R1176_U83, P2_U3170);
  nand ginst11963 (P2_R1176_U267, P2_R1176_U124, P2_R1176_U265);
  nand ginst11964 (P2_R1176_U268, P2_R1176_U46, P2_R1176_U469);
  nand ginst11965 (P2_R1176_U269, P2_R1176_U472, P2_R1176_U48);
  not ginst11966 (P2_R1176_U27, P2_U3179);
  nand ginst11967 (P2_R1176_U270, P2_R1176_U267, P2_R1176_U269);
  not ginst11968 (P2_R1176_U271, P2_R1176_U199);
  nand ginst11969 (P2_R1176_U272, P2_R1176_U44, P2_R1176_U478);
  nand ginst11970 (P2_R1176_U273, P2_R1176_U80, P2_U3169);
  not ginst11971 (P2_R1176_U274, P2_R1176_U197);
  nand ginst11972 (P2_R1176_U275, P2_R1176_U481, P2_R1176_U51);
  nand ginst11973 (P2_R1176_U276, P2_R1176_U197, P2_R1176_U275);
  nand ginst11974 (P2_R1176_U277, P2_R1176_U85, P2_U3168);
  not ginst11975 (P2_R1176_U278, P2_R1176_U61);
  nand ginst11976 (P2_R1176_U279, P2_R1176_U43, P2_R1176_U484);
  not ginst11977 (P2_R1176_U28, P2_U3177);
  nand ginst11978 (P2_R1176_U280, P2_R1176_U41, P2_R1176_U487);
  not ginst11979 (P2_R1176_U281, P2_R1176_U42);
  nand ginst11980 (P2_R1176_U282, P2_R1176_U42, P2_R1176_U43);
  nand ginst11981 (P2_R1176_U283, P2_R1176_U282, P2_R1176_U79);
  nand ginst11982 (P2_R1176_U284, P2_R1176_U281, P2_U3166);
  nand ginst11983 (P2_R1176_U285, P2_R1176_U61, P2_R1176_U7);
  not ginst11984 (P2_R1176_U286, P2_R1176_U195);
  nand ginst11985 (P2_R1176_U287, P2_R1176_U490, P2_R1176_U52);
  nand ginst11986 (P2_R1176_U288, P2_R1176_U195, P2_R1176_U287);
  nand ginst11987 (P2_R1176_U289, P2_R1176_U86, P2_U3165);
  nand ginst11988 (P2_R1176_U29, P2_R1176_U73, P2_U3177);
  not ginst11989 (P2_R1176_U290, P2_R1176_U193);
  nand ginst11990 (P2_R1176_U291, P2_R1176_U493, P2_R1176_U56);
  nand ginst11991 (P2_R1176_U292, P2_R1176_U496, P2_R1176_U53);
  nand ginst11992 (P2_R1176_U293, P2_R1176_U211, P2_R1176_U8);
  nand ginst11993 (P2_R1176_U294, P2_R1176_U88, P2_U3162);
  nand ginst11994 (P2_R1176_U295, P2_R1176_U128, P2_R1176_U293);
  nand ginst11995 (P2_R1176_U296, P2_R1176_U499, P2_R1176_U54);
  nand ginst11996 (P2_R1176_U297, P2_R1176_U493, P2_R1176_U56);
  nand ginst11997 (P2_R1176_U298, P2_R1176_U127, P2_R1176_U193);
  nand ginst11998 (P2_R1176_U299, P2_R1176_U295, P2_R1176_U297);
  not ginst11999 (P2_R1176_U30, P2_U3176);
  not ginst12000 (P2_R1176_U300, P2_R1176_U190);
  nand ginst12001 (P2_R1176_U301, P2_R1176_U502, P2_R1176_U57);
  nand ginst12002 (P2_R1176_U302, P2_R1176_U190, P2_R1176_U301);
  nand ginst12003 (P2_R1176_U303, P2_R1176_U90, P2_U3161);
  not ginst12004 (P2_R1176_U304, P2_R1176_U188);
  nand ginst12005 (P2_R1176_U305, P2_R1176_U505, P2_R1176_U58);
  nand ginst12006 (P2_R1176_U306, P2_R1176_U188, P2_R1176_U305);
  nand ginst12007 (P2_R1176_U307, P2_R1176_U91, P2_U3160);
  not ginst12008 (P2_R1176_U308, P2_R1176_U186);
  nand ginst12009 (P2_R1176_U309, P2_R1176_U38, P2_R1176_U508);
  not ginst12010 (P2_R1176_U31, P2_U3178);
  nand ginst12011 (P2_R1176_U310, P2_R1176_U209, P2_R1176_U212, P2_R1176_U311);
  nand ginst12012 (P2_R1176_U311, P2_R1176_U77, P2_U3157);
  nand ginst12013 (P2_R1176_U312, P2_R1176_U39, P2_R1176_U511);
  nand ginst12014 (P2_R1176_U313, P2_R1176_U40, P2_R1176_U463);
  nand ginst12015 (P2_R1176_U314, P2_R1176_U129, P2_R1176_U186);
  nand ginst12016 (P2_R1176_U315, P2_R1176_U310, P2_R1176_U375);
  not ginst12017 (P2_R1176_U316, P2_R1176_U185);
  nand ginst12018 (P2_R1176_U317, P2_R1176_U37, P2_R1176_U460);
  nand ginst12019 (P2_R1176_U318, P2_R1176_U74, P2_U3156);
  nand ginst12020 (P2_R1176_U319, P2_R1176_U74, P2_U3156);
  nand ginst12021 (P2_R1176_U32, P2_R1176_U71, P2_U3178);
  nand ginst12022 (P2_R1176_U320, P2_R1176_U37, P2_R1176_U460);
  nand ginst12023 (P2_R1176_U321, P2_R1176_U186, P2_R1176_U312);
  not ginst12024 (P2_R1176_U322, P2_R1176_U59);
  nand ginst12025 (P2_R1176_U323, P2_R1176_U12, P2_R1176_U135);
  nand ginst12026 (P2_R1176_U324, P2_R1176_U136, P2_R1176_U321);
  nand ginst12027 (P2_R1176_U325, P2_R1176_U77, P2_U3157);
  nand ginst12028 (P2_R1176_U326, P2_R1176_U137, P2_R1176_U324);
  nand ginst12029 (P2_R1176_U327, P2_R1176_U38, P2_R1176_U508);
  nand ginst12030 (P2_R1176_U328, P2_R1176_U193, P2_R1176_U296);
  not ginst12031 (P2_R1176_U329, P2_R1176_U60);
  not ginst12032 (P2_R1176_U33, P2_U3174);
  nand ginst12033 (P2_R1176_U330, P2_R1176_U496, P2_R1176_U53);
  nand ginst12034 (P2_R1176_U331, P2_R1176_U330, P2_R1176_U60);
  nand ginst12035 (P2_R1176_U332, P2_R1176_U139, P2_R1176_U331);
  nand ginst12036 (P2_R1176_U333, P2_R1176_U208, P2_R1176_U329);
  nand ginst12037 (P2_R1176_U334, P2_R1176_U88, P2_U3162);
  nand ginst12038 (P2_R1176_U335, P2_R1176_U140, P2_R1176_U333);
  nand ginst12039 (P2_R1176_U336, P2_R1176_U496, P2_R1176_U53);
  nand ginst12040 (P2_R1176_U337, P2_R1176_U41, P2_R1176_U487);
  nand ginst12041 (P2_R1176_U338, P2_R1176_U337, P2_R1176_U61);
  nand ginst12042 (P2_R1176_U339, P2_R1176_U141, P2_R1176_U338);
  nand ginst12043 (P2_R1176_U34, P2_R1176_U237, P2_R1176_U238, P2_R1176_U369);
  nand ginst12044 (P2_R1176_U340, P2_R1176_U278, P2_R1176_U42);
  nand ginst12045 (P2_R1176_U341, P2_R1176_U79, P2_U3166);
  nand ginst12046 (P2_R1176_U342, P2_R1176_U142, P2_R1176_U340);
  nand ginst12047 (P2_R1176_U343, P2_R1176_U41, P2_R1176_U487);
  nand ginst12048 (P2_R1176_U344, P2_R1176_U200, P2_R1176_U268);
  not ginst12049 (P2_R1176_U345, P2_R1176_U63);
  nand ginst12050 (P2_R1176_U346, P2_R1176_U45, P2_R1176_U475);
  nand ginst12051 (P2_R1176_U347, P2_R1176_U346, P2_R1176_U63);
  nand ginst12052 (P2_R1176_U348, P2_R1176_U143, P2_R1176_U347);
  nand ginst12053 (P2_R1176_U349, P2_R1176_U207, P2_R1176_U345);
  nand ginst12054 (P2_R1176_U35, P2_R1176_U230, P2_R1176_U32);
  nand ginst12055 (P2_R1176_U350, P2_R1176_U83, P2_U3170);
  nand ginst12056 (P2_R1176_U351, P2_R1176_U144, P2_R1176_U349);
  nand ginst12057 (P2_R1176_U352, P2_R1176_U45, P2_R1176_U475);
  nand ginst12058 (P2_R1176_U353, P2_R1176_U249, P2_R1176_U29);
  nand ginst12059 (P2_R1176_U354, P2_R1176_U22, P2_R1176_U256);
  nand ginst12060 (P2_R1176_U355, P2_R1176_U209, P2_R1176_U327);
  nand ginst12061 (P2_R1176_U356, P2_R1176_U212, P2_R1176_U312);
  nand ginst12062 (P2_R1176_U357, P2_R1176_U208, P2_R1176_U336);
  nand ginst12063 (P2_R1176_U358, P2_R1176_U296, P2_R1176_U55);
  nand ginst12064 (P2_R1176_U359, P2_R1176_U343, P2_R1176_U42);
  nand ginst12065 (P2_R1176_U36, P2_R1176_U218, P2_R1176_U365, P2_R1176_U366);
  nand ginst12066 (P2_R1176_U360, P2_R1176_U207, P2_R1176_U352);
  nand ginst12067 (P2_R1176_U361, P2_R1176_U268, P2_R1176_U47);
  nand ginst12068 (P2_R1176_U362, P2_R1176_U70, P2_U3179);
  nand ginst12069 (P2_R1176_U363, P2_R1176_U64, P2_U3174);
  nand ginst12070 (P2_R1176_U364, P2_R1176_U130, P2_R1176_U311, P2_R1176_U314);
  nand ginst12071 (P2_R1176_U365, P2_R1176_U213, P2_R1176_U367, P2_U3183);
  nand ginst12072 (P2_R1176_U366, P2_R1176_U215, P2_R1176_U217);
  nand ginst12073 (P2_R1176_U367, P2_R1176_U24, P2_R1176_U399);
  nand ginst12074 (P2_R1176_U368, P2_R1176_U10, P2_R1176_U161);
  nand ginst12075 (P2_R1176_U369, P2_R1176_U231, P2_R1176_U5);
  not ginst12076 (P2_R1176_U37, P2_U3156);
  not ginst12077 (P2_R1176_U370, P2_R1176_U34);
  nand ginst12078 (P2_R1176_U371, P2_R1176_U117, P2_R1176_U161);
  nand ginst12079 (P2_R1176_U372, P2_R1176_U240, P2_R1176_U34);
  nand ginst12080 (P2_R1176_U373, P2_R1176_U11, P2_R1176_U202);
  nand ginst12081 (P2_R1176_U374, P2_R1176_U261, P2_R1176_U9);
  nand ginst12082 (P2_R1176_U375, P2_R1176_U311, P2_R1176_U376, P2_R1176_U377);
  nand ginst12083 (P2_R1176_U376, P2_R1176_U309, P2_R1176_U77);
  nand ginst12084 (P2_R1176_U377, P2_R1176_U309, P2_U3157);
  not ginst12085 (P2_R1176_U378, P2_R1176_U62);
  nand ginst12086 (P2_R1176_U379, P2_R1176_U123, P2_R1176_U202);
  not ginst12087 (P2_R1176_U38, P2_U3158);
  nand ginst12088 (P2_R1176_U380, P2_R1176_U272, P2_R1176_U62);
  nand ginst12089 (P2_R1176_U381, P2_R1176_U131, P2_R1176_U375);
  nand ginst12090 (P2_R1176_U382, P2_R1176_U132, P2_R1176_U186, P2_R1176_U203);
  nand ginst12091 (P2_R1176_U383, P2_R1176_U309, P2_R1176_U313, P2_R1176_U384);
  nand ginst12092 (P2_R1176_U384, P2_R1176_U209, P2_R1176_U212);
  nand ginst12093 (P2_R1176_U385, P2_R1176_U138, P2_R1176_U322);
  nand ginst12094 (P2_R1176_U386, P2_R1176_U146, P2_U3184);
  nand ginst12095 (P2_R1176_U387, P2_R1176_U19, P2_U3456);
  not ginst12096 (P2_R1176_U388, P2_R1176_U64);
  nand ginst12097 (P2_R1176_U389, P2_R1176_U388, P2_U3174);
  not ginst12098 (P2_R1176_U39, P2_U3159);
  nand ginst12099 (P2_R1176_U390, P2_R1176_U33, P2_R1176_U64);
  nand ginst12100 (P2_R1176_U391, P2_R1176_U388, P2_U3174);
  nand ginst12101 (P2_R1176_U392, P2_R1176_U33, P2_R1176_U64);
  nand ginst12102 (P2_R1176_U393, P2_R1176_U391, P2_R1176_U392);
  nand ginst12103 (P2_R1176_U394, P2_R1176_U148, P2_U3184);
  nand ginst12104 (P2_R1176_U395, P2_R1176_U19, P2_U3441);
  not ginst12105 (P2_R1176_U396, P2_R1176_U70);
  nand ginst12106 (P2_R1176_U397, P2_R1176_U149, P2_U3184);
  nand ginst12107 (P2_R1176_U398, P2_R1176_U19, P2_U3432);
  not ginst12108 (P2_R1176_U399, P2_R1176_U68);
  and ginst12109 (P2_R1176_U4, P2_R1176_U220, P2_R1176_U221);
  not ginst12110 (P2_R1176_U40, P2_U3157);
  nand ginst12111 (P2_R1176_U400, P2_R1176_U150, P2_U3184);
  nand ginst12112 (P2_R1176_U401, P2_R1176_U19, P2_U3427);
  not ginst12113 (P2_R1176_U402, P2_R1176_U69);
  nand ginst12114 (P2_R1176_U403, P2_R1176_U151, P2_U3184);
  nand ginst12115 (P2_R1176_U404, P2_R1176_U19, P2_U3438);
  not ginst12116 (P2_R1176_U405, P2_R1176_U67);
  nand ginst12117 (P2_R1176_U406, P2_R1176_U152, P2_U3184);
  nand ginst12118 (P2_R1176_U407, P2_R1176_U19, P2_U3435);
  not ginst12119 (P2_R1176_U408, P2_R1176_U66);
  nand ginst12120 (P2_R1176_U409, P2_R1176_U153, P2_U3184);
  not ginst12121 (P2_R1176_U41, P2_U3167);
  nand ginst12122 (P2_R1176_U410, P2_R1176_U19, P2_U3444);
  not ginst12123 (P2_R1176_U411, P2_R1176_U71);
  nand ginst12124 (P2_R1176_U412, P2_R1176_U154, P2_U3184);
  nand ginst12125 (P2_R1176_U413, P2_R1176_U19, P2_U3450);
  not ginst12126 (P2_R1176_U414, P2_R1176_U72);
  nand ginst12127 (P2_R1176_U415, P2_R1176_U155, P2_U3184);
  nand ginst12128 (P2_R1176_U416, P2_R1176_U19, P2_U3447);
  not ginst12129 (P2_R1176_U417, P2_R1176_U73);
  nand ginst12130 (P2_R1176_U418, P2_R1176_U156, P2_U3184);
  nand ginst12131 (P2_R1176_U419, P2_R1176_U19, P2_U3453);
  nand ginst12132 (P2_R1176_U42, P2_R1176_U78, P2_U3167);
  not ginst12133 (P2_R1176_U420, P2_R1176_U65);
  nand ginst12134 (P2_R1176_U421, P2_R1176_U147, P2_R1176_U157);
  nand ginst12135 (P2_R1176_U422, P2_R1176_U242, P2_R1176_U393);
  nand ginst12136 (P2_R1176_U423, P2_R1176_U420, P2_U3175);
  nand ginst12137 (P2_R1176_U424, P2_R1176_U20, P2_R1176_U65);
  nand ginst12138 (P2_R1176_U425, P2_R1176_U420, P2_U3175);
  nand ginst12139 (P2_R1176_U426, P2_R1176_U20, P2_R1176_U65);
  nand ginst12140 (P2_R1176_U427, P2_R1176_U425, P2_R1176_U426);
  nand ginst12141 (P2_R1176_U428, P2_R1176_U158, P2_R1176_U159);
  nand ginst12142 (P2_R1176_U429, P2_R1176_U239, P2_R1176_U427);
  not ginst12143 (P2_R1176_U43, P2_U3166);
  nand ginst12144 (P2_R1176_U430, P2_R1176_U414, P2_U3176);
  nand ginst12145 (P2_R1176_U431, P2_R1176_U30, P2_R1176_U72);
  nand ginst12146 (P2_R1176_U432, P2_R1176_U417, P2_U3177);
  nand ginst12147 (P2_R1176_U433, P2_R1176_U28, P2_R1176_U73);
  nand ginst12148 (P2_R1176_U434, P2_R1176_U432, P2_R1176_U433);
  nand ginst12149 (P2_R1176_U435, P2_R1176_U35, P2_R1176_U353);
  nand ginst12150 (P2_R1176_U436, P2_R1176_U232, P2_R1176_U434);
  nand ginst12151 (P2_R1176_U437, P2_R1176_U411, P2_U3178);
  nand ginst12152 (P2_R1176_U438, P2_R1176_U31, P2_R1176_U71);
  nand ginst12153 (P2_R1176_U439, P2_R1176_U411, P2_U3178);
  not ginst12154 (P2_R1176_U44, P2_U3169);
  nand ginst12155 (P2_R1176_U440, P2_R1176_U31, P2_R1176_U71);
  nand ginst12156 (P2_R1176_U441, P2_R1176_U439, P2_R1176_U440);
  nand ginst12157 (P2_R1176_U442, P2_R1176_U160, P2_R1176_U161);
  nand ginst12158 (P2_R1176_U443, P2_R1176_U228, P2_R1176_U441);
  nand ginst12159 (P2_R1176_U444, P2_R1176_U396, P2_U3179);
  nand ginst12160 (P2_R1176_U445, P2_R1176_U27, P2_R1176_U70);
  nand ginst12161 (P2_R1176_U446, P2_R1176_U396, P2_U3179);
  nand ginst12162 (P2_R1176_U447, P2_R1176_U27, P2_R1176_U70);
  nand ginst12163 (P2_R1176_U448, P2_R1176_U446, P2_R1176_U447);
  nand ginst12164 (P2_R1176_U449, P2_R1176_U162, P2_R1176_U163);
  not ginst12165 (P2_R1176_U45, P2_U3171);
  nand ginst12166 (P2_R1176_U450, P2_R1176_U226, P2_R1176_U448);
  nand ginst12167 (P2_R1176_U451, P2_R1176_U405, P2_U3180);
  nand ginst12168 (P2_R1176_U452, P2_R1176_U23, P2_R1176_U67);
  nand ginst12169 (P2_R1176_U453, P2_R1176_U408, P2_U3181);
  nand ginst12170 (P2_R1176_U454, P2_R1176_U21, P2_R1176_U66);
  nand ginst12171 (P2_R1176_U455, P2_R1176_U453, P2_R1176_U454);
  nand ginst12172 (P2_R1176_U456, P2_R1176_U354, P2_R1176_U36);
  nand ginst12173 (P2_R1176_U457, P2_R1176_U219, P2_R1176_U455);
  nand ginst12174 (P2_R1176_U458, P2_R1176_U164, P2_U3184);
  nand ginst12175 (P2_R1176_U459, P2_R1176_U19, P2_U3950);
  not ginst12176 (P2_R1176_U46, P2_U3172);
  not ginst12177 (P2_R1176_U460, P2_R1176_U74);
  nand ginst12178 (P2_R1176_U461, P2_R1176_U165, P2_U3184);
  nand ginst12179 (P2_R1176_U462, P2_R1176_U19, P2_U3951);
  not ginst12180 (P2_R1176_U463, P2_R1176_U77);
  nand ginst12181 (P2_R1176_U464, P2_R1176_U166, P2_U3184);
  nand ginst12182 (P2_R1176_U465, P2_R1176_U19, P2_U3459);
  not ginst12183 (P2_R1176_U466, P2_R1176_U81);
  nand ginst12184 (P2_R1176_U467, P2_R1176_U167, P2_U3184);
  nand ginst12185 (P2_R1176_U468, P2_R1176_U19, P2_U3462);
  not ginst12186 (P2_R1176_U469, P2_R1176_U82);
  nand ginst12187 (P2_R1176_U47, P2_R1176_U82, P2_U3172);
  nand ginst12188 (P2_R1176_U470, P2_R1176_U168, P2_U3184);
  nand ginst12189 (P2_R1176_U471, P2_R1176_U19, P2_U3468);
  not ginst12190 (P2_R1176_U472, P2_R1176_U83);
  nand ginst12191 (P2_R1176_U473, P2_R1176_U169, P2_U3184);
  nand ginst12192 (P2_R1176_U474, P2_R1176_U19, P2_U3465);
  not ginst12193 (P2_R1176_U475, P2_R1176_U84);
  nand ginst12194 (P2_R1176_U476, P2_R1176_U170, P2_U3184);
  nand ginst12195 (P2_R1176_U477, P2_R1176_U19, P2_U3471);
  not ginst12196 (P2_R1176_U478, P2_R1176_U80);
  nand ginst12197 (P2_R1176_U479, P2_R1176_U171, P2_U3184);
  not ginst12198 (P2_R1176_U48, P2_U3170);
  nand ginst12199 (P2_R1176_U480, P2_R1176_U19, P2_U3474);
  not ginst12200 (P2_R1176_U481, P2_R1176_U85);
  nand ginst12201 (P2_R1176_U482, P2_R1176_U172, P2_U3184);
  nand ginst12202 (P2_R1176_U483, P2_R1176_U19, P2_U3480);
  not ginst12203 (P2_R1176_U484, P2_R1176_U79);
  nand ginst12204 (P2_R1176_U485, P2_R1176_U173, P2_U3184);
  nand ginst12205 (P2_R1176_U486, P2_R1176_U19, P2_U3477);
  not ginst12206 (P2_R1176_U487, P2_R1176_U78);
  nand ginst12207 (P2_R1176_U488, P2_R1176_U174, P2_U3184);
  nand ginst12208 (P2_R1176_U489, P2_R1176_U19, P2_U3483);
  not ginst12209 (P2_R1176_U49, P2_U3173);
  not ginst12210 (P2_R1176_U490, P2_R1176_U86);
  nand ginst12211 (P2_R1176_U491, P2_R1176_U175, P2_U3184);
  nand ginst12212 (P2_R1176_U492, P2_R1176_U19, P2_U3956);
  not ginst12213 (P2_R1176_U493, P2_R1176_U88);
  nand ginst12214 (P2_R1176_U494, P2_R1176_U176, P2_U3184);
  nand ginst12215 (P2_R1176_U495, P2_R1176_U19, P2_U3957);
  not ginst12216 (P2_R1176_U496, P2_R1176_U89);
  nand ginst12217 (P2_R1176_U497, P2_R1176_U177, P2_U3184);
  nand ginst12218 (P2_R1176_U498, P2_R1176_U19, P2_U3485);
  not ginst12219 (P2_R1176_U499, P2_R1176_U87);
  and ginst12220 (P2_R1176_U5, P2_R1176_U233, P2_R1176_U234);
  nand ginst12221 (P2_R1176_U50, P2_R1176_U81, P2_U3173);
  nand ginst12222 (P2_R1176_U500, P2_R1176_U178, P2_U3184);
  nand ginst12223 (P2_R1176_U501, P2_R1176_U19, P2_U3955);
  not ginst12224 (P2_R1176_U502, P2_R1176_U90);
  nand ginst12225 (P2_R1176_U503, P2_R1176_U179, P2_U3184);
  nand ginst12226 (P2_R1176_U504, P2_R1176_U19, P2_U3954);
  not ginst12227 (P2_R1176_U505, P2_R1176_U91);
  nand ginst12228 (P2_R1176_U506, P2_R1176_U180, P2_U3184);
  nand ginst12229 (P2_R1176_U507, P2_R1176_U19, P2_U3952);
  not ginst12230 (P2_R1176_U508, P2_R1176_U75);
  nand ginst12231 (P2_R1176_U509, P2_R1176_U181, P2_U3184);
  not ginst12232 (P2_R1176_U51, P2_U3168);
  nand ginst12233 (P2_R1176_U510, P2_R1176_U19, P2_U3953);
  not ginst12234 (P2_R1176_U511, P2_R1176_U76);
  nand ginst12235 (P2_R1176_U512, P2_R1176_U182, P2_U3184);
  nand ginst12236 (P2_R1176_U513, P2_R1176_U19, P2_U3949);
  not ginst12237 (P2_R1176_U514, P2_R1176_U134);
  nand ginst12238 (P2_R1176_U515, P2_R1176_U514, P2_U3155);
  nand ginst12239 (P2_R1176_U516, P2_R1176_U134, P2_R1176_U183);
  not ginst12240 (P2_R1176_U517, P2_R1176_U92);
  nand ginst12241 (P2_R1176_U518, P2_R1176_U317, P2_R1176_U364, P2_R1176_U517);
  nand ginst12242 (P2_R1176_U519, P2_R1176_U133, P2_R1176_U382, P2_R1176_U92);
  not ginst12243 (P2_R1176_U52, P2_U3165);
  nand ginst12244 (P2_R1176_U520, P2_R1176_U460, P2_U3156);
  nand ginst12245 (P2_R1176_U521, P2_R1176_U37, P2_R1176_U74);
  nand ginst12246 (P2_R1176_U522, P2_R1176_U460, P2_U3156);
  nand ginst12247 (P2_R1176_U523, P2_R1176_U37, P2_R1176_U74);
  nand ginst12248 (P2_R1176_U524, P2_R1176_U522, P2_R1176_U523);
  nand ginst12249 (P2_R1176_U525, P2_R1176_U184, P2_R1176_U185);
  nand ginst12250 (P2_R1176_U526, P2_R1176_U316, P2_R1176_U524);
  nand ginst12251 (P2_R1176_U527, P2_R1176_U463, P2_U3157);
  nand ginst12252 (P2_R1176_U528, P2_R1176_U40, P2_R1176_U77);
  nand ginst12253 (P2_R1176_U529, P2_R1176_U508, P2_U3158);
  not ginst12254 (P2_R1176_U53, P2_U3163);
  nand ginst12255 (P2_R1176_U530, P2_R1176_U38, P2_R1176_U75);
  nand ginst12256 (P2_R1176_U531, P2_R1176_U529, P2_R1176_U530);
  nand ginst12257 (P2_R1176_U532, P2_R1176_U355, P2_R1176_U59);
  nand ginst12258 (P2_R1176_U533, P2_R1176_U322, P2_R1176_U531);
  nand ginst12259 (P2_R1176_U534, P2_R1176_U511, P2_U3159);
  nand ginst12260 (P2_R1176_U535, P2_R1176_U39, P2_R1176_U76);
  nand ginst12261 (P2_R1176_U536, P2_R1176_U534, P2_R1176_U535);
  nand ginst12262 (P2_R1176_U537, P2_R1176_U186, P2_R1176_U356);
  nand ginst12263 (P2_R1176_U538, P2_R1176_U308, P2_R1176_U536);
  nand ginst12264 (P2_R1176_U539, P2_R1176_U505, P2_U3160);
  not ginst12265 (P2_R1176_U54, P2_U3164);
  nand ginst12266 (P2_R1176_U540, P2_R1176_U58, P2_R1176_U91);
  nand ginst12267 (P2_R1176_U541, P2_R1176_U505, P2_U3160);
  nand ginst12268 (P2_R1176_U542, P2_R1176_U58, P2_R1176_U91);
  nand ginst12269 (P2_R1176_U543, P2_R1176_U541, P2_R1176_U542);
  nand ginst12270 (P2_R1176_U544, P2_R1176_U187, P2_R1176_U188);
  nand ginst12271 (P2_R1176_U545, P2_R1176_U304, P2_R1176_U543);
  nand ginst12272 (P2_R1176_U546, P2_R1176_U502, P2_U3161);
  nand ginst12273 (P2_R1176_U547, P2_R1176_U57, P2_R1176_U90);
  nand ginst12274 (P2_R1176_U548, P2_R1176_U502, P2_U3161);
  nand ginst12275 (P2_R1176_U549, P2_R1176_U57, P2_R1176_U90);
  nand ginst12276 (P2_R1176_U55, P2_R1176_U87, P2_U3164);
  nand ginst12277 (P2_R1176_U550, P2_R1176_U548, P2_R1176_U549);
  nand ginst12278 (P2_R1176_U551, P2_R1176_U189, P2_R1176_U190);
  nand ginst12279 (P2_R1176_U552, P2_R1176_U300, P2_R1176_U550);
  nand ginst12280 (P2_R1176_U553, P2_R1176_U493, P2_U3162);
  nand ginst12281 (P2_R1176_U554, P2_R1176_U56, P2_R1176_U88);
  nand ginst12282 (P2_R1176_U555, P2_R1176_U496, P2_U3163);
  nand ginst12283 (P2_R1176_U556, P2_R1176_U53, P2_R1176_U89);
  nand ginst12284 (P2_R1176_U557, P2_R1176_U555, P2_R1176_U556);
  nand ginst12285 (P2_R1176_U558, P2_R1176_U357, P2_R1176_U60);
  nand ginst12286 (P2_R1176_U559, P2_R1176_U329, P2_R1176_U557);
  not ginst12287 (P2_R1176_U56, P2_U3162);
  nand ginst12288 (P2_R1176_U560, P2_R1176_U399, P2_U3182);
  nand ginst12289 (P2_R1176_U561, P2_R1176_U24, P2_R1176_U68);
  nand ginst12290 (P2_R1176_U562, P2_R1176_U399, P2_U3182);
  nand ginst12291 (P2_R1176_U563, P2_R1176_U24, P2_R1176_U68);
  nand ginst12292 (P2_R1176_U564, P2_R1176_U562, P2_R1176_U563);
  nand ginst12293 (P2_R1176_U565, P2_R1176_U191, P2_R1176_U192);
  nand ginst12294 (P2_R1176_U566, P2_R1176_U216, P2_R1176_U564);
  nand ginst12295 (P2_R1176_U567, P2_R1176_U499, P2_U3164);
  nand ginst12296 (P2_R1176_U568, P2_R1176_U54, P2_R1176_U87);
  nand ginst12297 (P2_R1176_U569, P2_R1176_U567, P2_R1176_U568);
  not ginst12298 (P2_R1176_U57, P2_U3161);
  nand ginst12299 (P2_R1176_U570, P2_R1176_U193, P2_R1176_U358);
  nand ginst12300 (P2_R1176_U571, P2_R1176_U290, P2_R1176_U569);
  nand ginst12301 (P2_R1176_U572, P2_R1176_U490, P2_U3165);
  nand ginst12302 (P2_R1176_U573, P2_R1176_U52, P2_R1176_U86);
  nand ginst12303 (P2_R1176_U574, P2_R1176_U490, P2_U3165);
  nand ginst12304 (P2_R1176_U575, P2_R1176_U52, P2_R1176_U86);
  nand ginst12305 (P2_R1176_U576, P2_R1176_U574, P2_R1176_U575);
  nand ginst12306 (P2_R1176_U577, P2_R1176_U194, P2_R1176_U195);
  nand ginst12307 (P2_R1176_U578, P2_R1176_U286, P2_R1176_U576);
  nand ginst12308 (P2_R1176_U579, P2_R1176_U484, P2_U3166);
  not ginst12309 (P2_R1176_U58, P2_U3160);
  nand ginst12310 (P2_R1176_U580, P2_R1176_U43, P2_R1176_U79);
  nand ginst12311 (P2_R1176_U581, P2_R1176_U487, P2_U3167);
  nand ginst12312 (P2_R1176_U582, P2_R1176_U41, P2_R1176_U78);
  nand ginst12313 (P2_R1176_U583, P2_R1176_U581, P2_R1176_U582);
  nand ginst12314 (P2_R1176_U584, P2_R1176_U359, P2_R1176_U61);
  nand ginst12315 (P2_R1176_U585, P2_R1176_U278, P2_R1176_U583);
  nand ginst12316 (P2_R1176_U586, P2_R1176_U481, P2_U3168);
  nand ginst12317 (P2_R1176_U587, P2_R1176_U51, P2_R1176_U85);
  nand ginst12318 (P2_R1176_U588, P2_R1176_U481, P2_U3168);
  nand ginst12319 (P2_R1176_U589, P2_R1176_U51, P2_R1176_U85);
  nand ginst12320 (P2_R1176_U59, P2_R1176_U212, P2_R1176_U321);
  nand ginst12321 (P2_R1176_U590, P2_R1176_U588, P2_R1176_U589);
  nand ginst12322 (P2_R1176_U591, P2_R1176_U196, P2_R1176_U197);
  nand ginst12323 (P2_R1176_U592, P2_R1176_U274, P2_R1176_U590);
  nand ginst12324 (P2_R1176_U593, P2_R1176_U478, P2_U3169);
  nand ginst12325 (P2_R1176_U594, P2_R1176_U44, P2_R1176_U80);
  nand ginst12326 (P2_R1176_U595, P2_R1176_U478, P2_U3169);
  nand ginst12327 (P2_R1176_U596, P2_R1176_U44, P2_R1176_U80);
  nand ginst12328 (P2_R1176_U597, P2_R1176_U595, P2_R1176_U596);
  nand ginst12329 (P2_R1176_U598, P2_R1176_U198, P2_R1176_U199);
  nand ginst12330 (P2_R1176_U599, P2_R1176_U271, P2_R1176_U597);
  and ginst12331 (P2_R1176_U6, P2_R1176_U263, P2_R1176_U264);
  nand ginst12332 (P2_R1176_U60, P2_R1176_U328, P2_R1176_U55);
  nand ginst12333 (P2_R1176_U600, P2_R1176_U472, P2_U3170);
  nand ginst12334 (P2_R1176_U601, P2_R1176_U48, P2_R1176_U83);
  nand ginst12335 (P2_R1176_U602, P2_R1176_U475, P2_U3171);
  nand ginst12336 (P2_R1176_U603, P2_R1176_U45, P2_R1176_U84);
  nand ginst12337 (P2_R1176_U604, P2_R1176_U602, P2_R1176_U603);
  nand ginst12338 (P2_R1176_U605, P2_R1176_U360, P2_R1176_U63);
  nand ginst12339 (P2_R1176_U606, P2_R1176_U345, P2_R1176_U604);
  nand ginst12340 (P2_R1176_U607, P2_R1176_U469, P2_U3172);
  nand ginst12341 (P2_R1176_U608, P2_R1176_U46, P2_R1176_U82);
  nand ginst12342 (P2_R1176_U609, P2_R1176_U607, P2_R1176_U608);
  nand ginst12343 (P2_R1176_U61, P2_R1176_U276, P2_R1176_U277);
  nand ginst12344 (P2_R1176_U610, P2_R1176_U200, P2_R1176_U361);
  nand ginst12345 (P2_R1176_U611, P2_R1176_U262, P2_R1176_U609);
  nand ginst12346 (P2_R1176_U612, P2_R1176_U466, P2_U3173);
  nand ginst12347 (P2_R1176_U613, P2_R1176_U49, P2_R1176_U81);
  nand ginst12348 (P2_R1176_U614, P2_R1176_U466, P2_U3173);
  nand ginst12349 (P2_R1176_U615, P2_R1176_U49, P2_R1176_U81);
  nand ginst12350 (P2_R1176_U616, P2_R1176_U614, P2_R1176_U615);
  nand ginst12351 (P2_R1176_U617, P2_R1176_U201, P2_R1176_U202);
  nand ginst12352 (P2_R1176_U618, P2_R1176_U258, P2_R1176_U616);
  nand ginst12353 (P2_R1176_U619, P2_R1176_U19, P2_R1176_U69);
  nand ginst12354 (P2_R1176_U62, P2_R1176_U270, P2_R1176_U374);
  nand ginst12355 (P2_R1176_U620, P2_R1176_U402, P2_U3184);
  not ginst12356 (P2_R1176_U621, P2_R1176_U145);
  nand ginst12357 (P2_R1176_U622, P2_R1176_U621, P2_U3183);
  nand ginst12358 (P2_R1176_U623, P2_R1176_U145, P2_R1176_U25);
  nand ginst12359 (P2_R1176_U63, P2_R1176_U344, P2_R1176_U47);
  nand ginst12360 (P2_R1176_U64, P2_R1176_U386, P2_R1176_U387);
  nand ginst12361 (P2_R1176_U65, P2_R1176_U418, P2_R1176_U419);
  nand ginst12362 (P2_R1176_U66, P2_R1176_U406, P2_R1176_U407);
  nand ginst12363 (P2_R1176_U67, P2_R1176_U403, P2_R1176_U404);
  nand ginst12364 (P2_R1176_U68, P2_R1176_U397, P2_R1176_U398);
  nand ginst12365 (P2_R1176_U69, P2_R1176_U400, P2_R1176_U401);
  and ginst12366 (P2_R1176_U7, P2_R1176_U279, P2_R1176_U280);
  nand ginst12367 (P2_R1176_U70, P2_R1176_U394, P2_R1176_U395);
  nand ginst12368 (P2_R1176_U71, P2_R1176_U409, P2_R1176_U410);
  nand ginst12369 (P2_R1176_U72, P2_R1176_U412, P2_R1176_U413);
  nand ginst12370 (P2_R1176_U73, P2_R1176_U415, P2_R1176_U416);
  nand ginst12371 (P2_R1176_U74, P2_R1176_U458, P2_R1176_U459);
  nand ginst12372 (P2_R1176_U75, P2_R1176_U506, P2_R1176_U507);
  nand ginst12373 (P2_R1176_U76, P2_R1176_U509, P2_R1176_U510);
  nand ginst12374 (P2_R1176_U77, P2_R1176_U461, P2_R1176_U462);
  nand ginst12375 (P2_R1176_U78, P2_R1176_U485, P2_R1176_U486);
  nand ginst12376 (P2_R1176_U79, P2_R1176_U482, P2_R1176_U483);
  and ginst12377 (P2_R1176_U8, P2_R1176_U291, P2_R1176_U292);
  nand ginst12378 (P2_R1176_U80, P2_R1176_U476, P2_R1176_U477);
  nand ginst12379 (P2_R1176_U81, P2_R1176_U464, P2_R1176_U465);
  nand ginst12380 (P2_R1176_U82, P2_R1176_U467, P2_R1176_U468);
  nand ginst12381 (P2_R1176_U83, P2_R1176_U470, P2_R1176_U471);
  nand ginst12382 (P2_R1176_U84, P2_R1176_U473, P2_R1176_U474);
  nand ginst12383 (P2_R1176_U85, P2_R1176_U479, P2_R1176_U480);
  nand ginst12384 (P2_R1176_U86, P2_R1176_U488, P2_R1176_U489);
  nand ginst12385 (P2_R1176_U87, P2_R1176_U497, P2_R1176_U498);
  nand ginst12386 (P2_R1176_U88, P2_R1176_U491, P2_R1176_U492);
  nand ginst12387 (P2_R1176_U89, P2_R1176_U494, P2_R1176_U495);
  and ginst12388 (P2_R1176_U9, P2_R1176_U268, P2_R1176_U6);
  nand ginst12389 (P2_R1176_U90, P2_R1176_U500, P2_R1176_U501);
  nand ginst12390 (P2_R1176_U91, P2_R1176_U503, P2_R1176_U504);
  nand ginst12391 (P2_R1176_U92, P2_R1176_U515, P2_R1176_U516);
  nand ginst12392 (P2_R1176_U93, P2_R1176_U622, P2_R1176_U623);
  nand ginst12393 (P2_R1176_U94, P2_R1176_U421, P2_R1176_U422);
  nand ginst12394 (P2_R1176_U95, P2_R1176_U428, P2_R1176_U429);
  nand ginst12395 (P2_R1176_U96, P2_R1176_U435, P2_R1176_U436);
  nand ginst12396 (P2_R1176_U97, P2_R1176_U442, P2_R1176_U443);
  nand ginst12397 (P2_R1176_U98, P2_R1176_U449, P2_R1176_U450);
  nand ginst12398 (P2_R1176_U99, P2_R1176_U456, P2_R1176_U457);
  and ginst12399 (P2_R1179_U10, P2_R1179_U182, P2_R1179_U282);
  nand ginst12400 (P2_R1179_U100, P2_R1179_U449, P2_R1179_U450);
  nand ginst12401 (P2_R1179_U101, P2_R1179_U465, P2_R1179_U466);
  nand ginst12402 (P2_R1179_U102, P2_R1179_U470, P2_R1179_U471);
  nand ginst12403 (P2_R1179_U103, P2_R1179_U355, P2_R1179_U356);
  nand ginst12404 (P2_R1179_U104, P2_R1179_U364, P2_R1179_U365);
  nand ginst12405 (P2_R1179_U105, P2_R1179_U371, P2_R1179_U372);
  nand ginst12406 (P2_R1179_U106, P2_R1179_U375, P2_R1179_U376);
  nand ginst12407 (P2_R1179_U107, P2_R1179_U384, P2_R1179_U385);
  nand ginst12408 (P2_R1179_U108, P2_R1179_U403, P2_R1179_U404);
  nand ginst12409 (P2_R1179_U109, P2_R1179_U420, P2_R1179_U421);
  and ginst12410 (P2_R1179_U11, P2_R1179_U283, P2_R1179_U284);
  nand ginst12411 (P2_R1179_U110, P2_R1179_U424, P2_R1179_U425);
  nand ginst12412 (P2_R1179_U111, P2_R1179_U456, P2_R1179_U457);
  nand ginst12413 (P2_R1179_U112, P2_R1179_U460, P2_R1179_U461);
  nand ginst12414 (P2_R1179_U113, P2_R1179_U477, P2_R1179_U478);
  and ginst12415 (P2_R1179_U114, P2_R1179_U184, P2_R1179_U194);
  and ginst12416 (P2_R1179_U115, P2_R1179_U197, P2_R1179_U198);
  and ginst12417 (P2_R1179_U116, P2_R1179_U185, P2_R1179_U200, P2_R1179_U205);
  and ginst12418 (P2_R1179_U117, P2_R1179_U186, P2_R1179_U210);
  and ginst12419 (P2_R1179_U118, P2_R1179_U213, P2_R1179_U214);
  and ginst12420 (P2_R1179_U119, P2_R1179_U357, P2_R1179_U358, P2_R1179_U38);
  nand ginst12421 (P2_R1179_U12, P2_R1179_U344, P2_R1179_U347);
  and ginst12422 (P2_R1179_U120, P2_R1179_U186, P2_R1179_U361);
  and ginst12423 (P2_R1179_U121, P2_R1179_U229, P2_R1179_U6);
  and ginst12424 (P2_R1179_U122, P2_R1179_U185, P2_R1179_U368);
  and ginst12425 (P2_R1179_U123, P2_R1179_U28, P2_R1179_U377, P2_R1179_U378);
  and ginst12426 (P2_R1179_U124, P2_R1179_U184, P2_R1179_U381);
  and ginst12427 (P2_R1179_U125, P2_R1179_U180, P2_R1179_U216, P2_R1179_U239);
  and ginst12428 (P2_R1179_U126, P2_R1179_U261, P2_R1179_U8);
  and ginst12429 (P2_R1179_U127, P2_R1179_U10, P2_R1179_U287);
  and ginst12430 (P2_R1179_U128, P2_R1179_U303, P2_R1179_U304);
  and ginst12431 (P2_R1179_U129, P2_R1179_U311, P2_R1179_U386, P2_R1179_U387);
  nand ginst12432 (P2_R1179_U13, P2_R1179_U333, P2_R1179_U336);
  and ginst12433 (P2_R1179_U130, P2_R1179_U308, P2_R1179_U390);
  nand ginst12434 (P2_R1179_U131, P2_R1179_U391, P2_R1179_U392);
  and ginst12435 (P2_R1179_U132, P2_R1179_U396, P2_R1179_U397, P2_R1179_U83);
  and ginst12436 (P2_R1179_U133, P2_R1179_U183, P2_R1179_U400);
  nand ginst12437 (P2_R1179_U134, P2_R1179_U405, P2_R1179_U406);
  nand ginst12438 (P2_R1179_U135, P2_R1179_U410, P2_R1179_U411);
  and ginst12439 (P2_R1179_U136, P2_R1179_U11, P2_R1179_U324);
  and ginst12440 (P2_R1179_U137, P2_R1179_U182, P2_R1179_U417);
  nand ginst12441 (P2_R1179_U138, P2_R1179_U426, P2_R1179_U427);
  nand ginst12442 (P2_R1179_U139, P2_R1179_U431, P2_R1179_U432);
  nand ginst12443 (P2_R1179_U14, P2_R1179_U322, P2_R1179_U325);
  nand ginst12444 (P2_R1179_U140, P2_R1179_U436, P2_R1179_U437);
  nand ginst12445 (P2_R1179_U141, P2_R1179_U441, P2_R1179_U442);
  nand ginst12446 (P2_R1179_U142, P2_R1179_U446, P2_R1179_U447);
  and ginst12447 (P2_R1179_U143, P2_R1179_U335, P2_R1179_U9);
  and ginst12448 (P2_R1179_U144, P2_R1179_U181, P2_R1179_U453);
  nand ginst12449 (P2_R1179_U145, P2_R1179_U462, P2_R1179_U463);
  nand ginst12450 (P2_R1179_U146, P2_R1179_U467, P2_R1179_U468);
  and ginst12451 (P2_R1179_U147, P2_R1179_U346, P2_R1179_U7);
  and ginst12452 (P2_R1179_U148, P2_R1179_U180, P2_R1179_U474);
  and ginst12453 (P2_R1179_U149, P2_R1179_U353, P2_R1179_U354);
  nand ginst12454 (P2_R1179_U15, P2_R1179_U314, P2_R1179_U316);
  nand ginst12455 (P2_R1179_U150, P2_R1179_U118, P2_R1179_U211);
  and ginst12456 (P2_R1179_U151, P2_R1179_U362, P2_R1179_U363);
  and ginst12457 (P2_R1179_U152, P2_R1179_U369, P2_R1179_U370);
  and ginst12458 (P2_R1179_U153, P2_R1179_U373, P2_R1179_U374);
  nand ginst12459 (P2_R1179_U154, P2_R1179_U115, P2_R1179_U195);
  and ginst12460 (P2_R1179_U155, P2_R1179_U382, P2_R1179_U383);
  not ginst12461 (P2_R1179_U156, P2_U3960);
  not ginst12462 (P2_R1179_U157, P2_U3057);
  and ginst12463 (P2_R1179_U158, P2_R1179_U401, P2_R1179_U402);
  nand ginst12464 (P2_R1179_U159, P2_R1179_U293, P2_R1179_U294);
  nand ginst12465 (P2_R1179_U16, P2_R1179_U312, P2_R1179_U352);
  nand ginst12466 (P2_R1179_U160, P2_R1179_U289, P2_R1179_U290);
  and ginst12467 (P2_R1179_U161, P2_R1179_U418, P2_R1179_U419);
  and ginst12468 (P2_R1179_U162, P2_R1179_U422, P2_R1179_U423);
  nand ginst12469 (P2_R1179_U163, P2_R1179_U279, P2_R1179_U280);
  nand ginst12470 (P2_R1179_U164, P2_R1179_U275, P2_R1179_U276);
  not ginst12471 (P2_R1179_U165, P2_U3432);
  nand ginst12472 (P2_R1179_U166, P2_R1179_U92, P2_U3427);
  nand ginst12473 (P2_R1179_U167, P2_R1179_U271, P2_R1179_U272);
  not ginst12474 (P2_R1179_U168, P2_U3483);
  nand ginst12475 (P2_R1179_U169, P2_R1179_U263, P2_R1179_U264);
  nand ginst12476 (P2_R1179_U17, P2_R1179_U235, P2_R1179_U237);
  and ginst12477 (P2_R1179_U170, P2_R1179_U454, P2_R1179_U455);
  and ginst12478 (P2_R1179_U171, P2_R1179_U458, P2_R1179_U459);
  nand ginst12479 (P2_R1179_U172, P2_R1179_U253, P2_R1179_U254);
  nand ginst12480 (P2_R1179_U173, P2_R1179_U249, P2_R1179_U250);
  nand ginst12481 (P2_R1179_U174, P2_R1179_U245, P2_R1179_U246);
  and ginst12482 (P2_R1179_U175, P2_R1179_U475, P2_R1179_U476);
  nand ginst12483 (P2_R1179_U176, P2_R1179_U165, P2_R1179_U166);
  not ginst12484 (P2_R1179_U177, P2_R1179_U83);
  not ginst12485 (P2_R1179_U178, P2_R1179_U28);
  not ginst12486 (P2_R1179_U179, P2_R1179_U38);
  nand ginst12487 (P2_R1179_U18, P2_R1179_U227, P2_R1179_U230);
  nand ginst12488 (P2_R1179_U180, P2_R1179_U49, P2_U3459);
  nand ginst12489 (P2_R1179_U181, P2_R1179_U59, P2_U3474);
  nand ginst12490 (P2_R1179_U182, P2_R1179_U74, P2_U3955);
  nand ginst12491 (P2_R1179_U183, P2_R1179_U82, P2_U3951);
  nand ginst12492 (P2_R1179_U184, P2_R1179_U27, P2_U3435);
  nand ginst12493 (P2_R1179_U185, P2_R1179_U33, P2_U3444);
  nand ginst12494 (P2_R1179_U186, P2_R1179_U37, P2_U3450);
  not ginst12495 (P2_R1179_U187, P2_R1179_U61);
  not ginst12496 (P2_R1179_U188, P2_R1179_U76);
  not ginst12497 (P2_R1179_U189, P2_R1179_U35);
  nand ginst12498 (P2_R1179_U19, P2_R1179_U219, P2_R1179_U221);
  not ginst12499 (P2_R1179_U190, P2_R1179_U50);
  not ginst12500 (P2_R1179_U191, P2_R1179_U166);
  nand ginst12501 (P2_R1179_U192, P2_R1179_U166, P2_U3080);
  not ginst12502 (P2_R1179_U193, P2_R1179_U44);
  nand ginst12503 (P2_R1179_U194, P2_R1179_U29, P2_U3438);
  nand ginst12504 (P2_R1179_U195, P2_R1179_U114, P2_R1179_U44);
  nand ginst12505 (P2_R1179_U196, P2_R1179_U28, P2_R1179_U29);
  nand ginst12506 (P2_R1179_U197, P2_R1179_U196, P2_R1179_U26);
  nand ginst12507 (P2_R1179_U198, P2_R1179_U178, P2_U3066);
  not ginst12508 (P2_R1179_U199, P2_R1179_U154);
  nand ginst12509 (P2_R1179_U20, P2_R1179_U166, P2_R1179_U350);
  nand ginst12510 (P2_R1179_U200, P2_R1179_U32, P2_U3447);
  nand ginst12511 (P2_R1179_U201, P2_R1179_U30, P2_U3073);
  nand ginst12512 (P2_R1179_U202, P2_R1179_U22, P2_U3069);
  nand ginst12513 (P2_R1179_U203, P2_R1179_U185, P2_R1179_U189);
  nand ginst12514 (P2_R1179_U204, P2_R1179_U203, P2_R1179_U6);
  nand ginst12515 (P2_R1179_U205, P2_R1179_U34, P2_U3441);
  nand ginst12516 (P2_R1179_U206, P2_R1179_U32, P2_U3447);
  nand ginst12517 (P2_R1179_U207, P2_R1179_U116, P2_R1179_U154);
  nand ginst12518 (P2_R1179_U208, P2_R1179_U204, P2_R1179_U206);
  not ginst12519 (P2_R1179_U209, P2_R1179_U42);
  not ginst12520 (P2_R1179_U21, P2_U3450);
  nand ginst12521 (P2_R1179_U210, P2_R1179_U39, P2_U3453);
  nand ginst12522 (P2_R1179_U211, P2_R1179_U117, P2_R1179_U42);
  nand ginst12523 (P2_R1179_U212, P2_R1179_U38, P2_R1179_U39);
  nand ginst12524 (P2_R1179_U213, P2_R1179_U212, P2_R1179_U36);
  nand ginst12525 (P2_R1179_U214, P2_R1179_U179, P2_U3086);
  not ginst12526 (P2_R1179_U215, P2_R1179_U150);
  nand ginst12527 (P2_R1179_U216, P2_R1179_U41, P2_U3456);
  nand ginst12528 (P2_R1179_U217, P2_R1179_U216, P2_R1179_U50);
  nand ginst12529 (P2_R1179_U218, P2_R1179_U209, P2_R1179_U38);
  nand ginst12530 (P2_R1179_U219, P2_R1179_U120, P2_R1179_U218);
  not ginst12531 (P2_R1179_U22, P2_U3444);
  nand ginst12532 (P2_R1179_U220, P2_R1179_U186, P2_R1179_U42);
  nand ginst12533 (P2_R1179_U221, P2_R1179_U119, P2_R1179_U220);
  nand ginst12534 (P2_R1179_U222, P2_R1179_U186, P2_R1179_U38);
  nand ginst12535 (P2_R1179_U223, P2_R1179_U154, P2_R1179_U205);
  not ginst12536 (P2_R1179_U224, P2_R1179_U43);
  nand ginst12537 (P2_R1179_U225, P2_R1179_U22, P2_U3069);
  nand ginst12538 (P2_R1179_U226, P2_R1179_U224, P2_R1179_U225);
  nand ginst12539 (P2_R1179_U227, P2_R1179_U122, P2_R1179_U226);
  nand ginst12540 (P2_R1179_U228, P2_R1179_U185, P2_R1179_U43);
  nand ginst12541 (P2_R1179_U229, P2_R1179_U32, P2_U3447);
  not ginst12542 (P2_R1179_U23, P2_U3435);
  nand ginst12543 (P2_R1179_U230, P2_R1179_U121, P2_R1179_U228);
  nand ginst12544 (P2_R1179_U231, P2_R1179_U22, P2_U3069);
  nand ginst12545 (P2_R1179_U232, P2_R1179_U185, P2_R1179_U231);
  nand ginst12546 (P2_R1179_U233, P2_R1179_U205, P2_R1179_U35);
  nand ginst12547 (P2_R1179_U234, P2_R1179_U193, P2_R1179_U28);
  nand ginst12548 (P2_R1179_U235, P2_R1179_U124, P2_R1179_U234);
  nand ginst12549 (P2_R1179_U236, P2_R1179_U184, P2_R1179_U44);
  nand ginst12550 (P2_R1179_U237, P2_R1179_U123, P2_R1179_U236);
  nand ginst12551 (P2_R1179_U238, P2_R1179_U184, P2_R1179_U28);
  nand ginst12552 (P2_R1179_U239, P2_R1179_U48, P2_U3462);
  not ginst12553 (P2_R1179_U24, P2_U3427);
  nand ginst12554 (P2_R1179_U240, P2_R1179_U47, P2_U3065);
  nand ginst12555 (P2_R1179_U241, P2_R1179_U46, P2_U3064);
  nand ginst12556 (P2_R1179_U242, P2_R1179_U180, P2_R1179_U190);
  nand ginst12557 (P2_R1179_U243, P2_R1179_U242, P2_R1179_U7);
  nand ginst12558 (P2_R1179_U244, P2_R1179_U48, P2_U3462);
  nand ginst12559 (P2_R1179_U245, P2_R1179_U125, P2_R1179_U150);
  nand ginst12560 (P2_R1179_U246, P2_R1179_U243, P2_R1179_U244);
  not ginst12561 (P2_R1179_U247, P2_R1179_U174);
  nand ginst12562 (P2_R1179_U248, P2_R1179_U52, P2_U3465);
  nand ginst12563 (P2_R1179_U249, P2_R1179_U174, P2_R1179_U248);
  not ginst12564 (P2_R1179_U25, P2_U3080);
  nand ginst12565 (P2_R1179_U250, P2_R1179_U51, P2_U3074);
  not ginst12566 (P2_R1179_U251, P2_R1179_U173);
  nand ginst12567 (P2_R1179_U252, P2_R1179_U54, P2_U3468);
  nand ginst12568 (P2_R1179_U253, P2_R1179_U173, P2_R1179_U252);
  nand ginst12569 (P2_R1179_U254, P2_R1179_U53, P2_U3082);
  not ginst12570 (P2_R1179_U255, P2_R1179_U172);
  nand ginst12571 (P2_R1179_U256, P2_R1179_U58, P2_U3477);
  nand ginst12572 (P2_R1179_U257, P2_R1179_U55, P2_U3075);
  nand ginst12573 (P2_R1179_U258, P2_R1179_U56, P2_U3076);
  nand ginst12574 (P2_R1179_U259, P2_R1179_U187, P2_R1179_U8);
  not ginst12575 (P2_R1179_U26, P2_U3438);
  nand ginst12576 (P2_R1179_U260, P2_R1179_U259, P2_R1179_U9);
  nand ginst12577 (P2_R1179_U261, P2_R1179_U60, P2_U3471);
  nand ginst12578 (P2_R1179_U262, P2_R1179_U58, P2_U3477);
  nand ginst12579 (P2_R1179_U263, P2_R1179_U126, P2_R1179_U172);
  nand ginst12580 (P2_R1179_U264, P2_R1179_U260, P2_R1179_U262);
  not ginst12581 (P2_R1179_U265, P2_R1179_U169);
  nand ginst12582 (P2_R1179_U266, P2_R1179_U63, P2_U3480);
  nand ginst12583 (P2_R1179_U267, P2_R1179_U169, P2_R1179_U266);
  nand ginst12584 (P2_R1179_U268, P2_R1179_U62, P2_U3071);
  not ginst12585 (P2_R1179_U269, P2_R1179_U64);
  not ginst12586 (P2_R1179_U27, P2_U3070);
  nand ginst12587 (P2_R1179_U270, P2_R1179_U269, P2_R1179_U65);
  nand ginst12588 (P2_R1179_U271, P2_R1179_U168, P2_R1179_U270);
  nand ginst12589 (P2_R1179_U272, P2_R1179_U64, P2_U3084);
  not ginst12590 (P2_R1179_U273, P2_R1179_U167);
  nand ginst12591 (P2_R1179_U274, P2_R1179_U67, P2_U3485);
  nand ginst12592 (P2_R1179_U275, P2_R1179_U167, P2_R1179_U274);
  nand ginst12593 (P2_R1179_U276, P2_R1179_U66, P2_U3083);
  not ginst12594 (P2_R1179_U277, P2_R1179_U164);
  nand ginst12595 (P2_R1179_U278, P2_R1179_U69, P2_U3957);
  nand ginst12596 (P2_R1179_U279, P2_R1179_U164, P2_R1179_U278);
  nand ginst12597 (P2_R1179_U28, P2_R1179_U23, P2_U3070);
  nand ginst12598 (P2_R1179_U280, P2_R1179_U68, P2_U3078);
  not ginst12599 (P2_R1179_U281, P2_R1179_U163);
  nand ginst12600 (P2_R1179_U282, P2_R1179_U73, P2_U3954);
  nand ginst12601 (P2_R1179_U283, P2_R1179_U70, P2_U3068);
  nand ginst12602 (P2_R1179_U284, P2_R1179_U71, P2_U3063);
  nand ginst12603 (P2_R1179_U285, P2_R1179_U10, P2_R1179_U188);
  nand ginst12604 (P2_R1179_U286, P2_R1179_U11, P2_R1179_U285);
  nand ginst12605 (P2_R1179_U287, P2_R1179_U75, P2_U3956);
  nand ginst12606 (P2_R1179_U288, P2_R1179_U73, P2_U3954);
  nand ginst12607 (P2_R1179_U289, P2_R1179_U127, P2_R1179_U163);
  not ginst12608 (P2_R1179_U29, P2_U3066);
  nand ginst12609 (P2_R1179_U290, P2_R1179_U286, P2_R1179_U288);
  not ginst12610 (P2_R1179_U291, P2_R1179_U160);
  nand ginst12611 (P2_R1179_U292, P2_R1179_U78, P2_U3953);
  nand ginst12612 (P2_R1179_U293, P2_R1179_U160, P2_R1179_U292);
  nand ginst12613 (P2_R1179_U294, P2_R1179_U77, P2_U3067);
  not ginst12614 (P2_R1179_U295, P2_R1179_U159);
  nand ginst12615 (P2_R1179_U296, P2_R1179_U80, P2_U3952);
  nand ginst12616 (P2_R1179_U297, P2_R1179_U159, P2_R1179_U296);
  nand ginst12617 (P2_R1179_U298, P2_R1179_U79, P2_U3060);
  not ginst12618 (P2_R1179_U299, P2_R1179_U88);
  not ginst12619 (P2_R1179_U30, P2_U3447);
  nand ginst12620 (P2_R1179_U300, P2_R1179_U84, P2_U3950);
  nand ginst12621 (P2_R1179_U301, P2_R1179_U183, P2_R1179_U300, P2_R1179_U88);
  nand ginst12622 (P2_R1179_U302, P2_R1179_U83, P2_R1179_U84);
  nand ginst12623 (P2_R1179_U303, P2_R1179_U302, P2_R1179_U81);
  nand ginst12624 (P2_R1179_U304, P2_R1179_U177, P2_U3055);
  not ginst12625 (P2_R1179_U305, P2_R1179_U87);
  nand ginst12626 (P2_R1179_U306, P2_R1179_U85, P2_U3056);
  nand ginst12627 (P2_R1179_U307, P2_R1179_U305, P2_R1179_U306);
  nand ginst12628 (P2_R1179_U308, P2_R1179_U86, P2_U3949);
  nand ginst12629 (P2_R1179_U309, P2_R1179_U86, P2_U3949);
  not ginst12630 (P2_R1179_U31, P2_U3441);
  nand ginst12631 (P2_R1179_U310, P2_R1179_U309, P2_R1179_U87);
  nand ginst12632 (P2_R1179_U311, P2_R1179_U85, P2_U3056);
  nand ginst12633 (P2_R1179_U312, P2_R1179_U129, P2_R1179_U310);
  nand ginst12634 (P2_R1179_U313, P2_R1179_U299, P2_R1179_U83);
  nand ginst12635 (P2_R1179_U314, P2_R1179_U133, P2_R1179_U313);
  nand ginst12636 (P2_R1179_U315, P2_R1179_U183, P2_R1179_U88);
  nand ginst12637 (P2_R1179_U316, P2_R1179_U132, P2_R1179_U315);
  nand ginst12638 (P2_R1179_U317, P2_R1179_U183, P2_R1179_U83);
  nand ginst12639 (P2_R1179_U318, P2_R1179_U163, P2_R1179_U287);
  not ginst12640 (P2_R1179_U319, P2_R1179_U89);
  not ginst12641 (P2_R1179_U32, P2_U3073);
  nand ginst12642 (P2_R1179_U320, P2_R1179_U71, P2_U3063);
  nand ginst12643 (P2_R1179_U321, P2_R1179_U319, P2_R1179_U320);
  nand ginst12644 (P2_R1179_U322, P2_R1179_U137, P2_R1179_U321);
  nand ginst12645 (P2_R1179_U323, P2_R1179_U182, P2_R1179_U89);
  nand ginst12646 (P2_R1179_U324, P2_R1179_U73, P2_U3954);
  nand ginst12647 (P2_R1179_U325, P2_R1179_U136, P2_R1179_U323);
  nand ginst12648 (P2_R1179_U326, P2_R1179_U71, P2_U3063);
  nand ginst12649 (P2_R1179_U327, P2_R1179_U182, P2_R1179_U326);
  nand ginst12650 (P2_R1179_U328, P2_R1179_U287, P2_R1179_U76);
  nand ginst12651 (P2_R1179_U329, P2_R1179_U172, P2_R1179_U261);
  not ginst12652 (P2_R1179_U33, P2_U3069);
  not ginst12653 (P2_R1179_U330, P2_R1179_U90);
  nand ginst12654 (P2_R1179_U331, P2_R1179_U56, P2_U3076);
  nand ginst12655 (P2_R1179_U332, P2_R1179_U330, P2_R1179_U331);
  nand ginst12656 (P2_R1179_U333, P2_R1179_U144, P2_R1179_U332);
  nand ginst12657 (P2_R1179_U334, P2_R1179_U181, P2_R1179_U90);
  nand ginst12658 (P2_R1179_U335, P2_R1179_U58, P2_U3477);
  nand ginst12659 (P2_R1179_U336, P2_R1179_U143, P2_R1179_U334);
  nand ginst12660 (P2_R1179_U337, P2_R1179_U56, P2_U3076);
  nand ginst12661 (P2_R1179_U338, P2_R1179_U181, P2_R1179_U337);
  nand ginst12662 (P2_R1179_U339, P2_R1179_U261, P2_R1179_U61);
  not ginst12663 (P2_R1179_U34, P2_U3062);
  nand ginst12664 (P2_R1179_U340, P2_R1179_U150, P2_R1179_U216);
  not ginst12665 (P2_R1179_U341, P2_R1179_U91);
  nand ginst12666 (P2_R1179_U342, P2_R1179_U46, P2_U3064);
  nand ginst12667 (P2_R1179_U343, P2_R1179_U341, P2_R1179_U342);
  nand ginst12668 (P2_R1179_U344, P2_R1179_U148, P2_R1179_U343);
  nand ginst12669 (P2_R1179_U345, P2_R1179_U180, P2_R1179_U91);
  nand ginst12670 (P2_R1179_U346, P2_R1179_U48, P2_U3462);
  nand ginst12671 (P2_R1179_U347, P2_R1179_U147, P2_R1179_U345);
  nand ginst12672 (P2_R1179_U348, P2_R1179_U46, P2_U3064);
  nand ginst12673 (P2_R1179_U349, P2_R1179_U180, P2_R1179_U348);
  nand ginst12674 (P2_R1179_U35, P2_R1179_U31, P2_U3062);
  nand ginst12675 (P2_R1179_U350, P2_R1179_U24, P2_U3079);
  nand ginst12676 (P2_R1179_U351, P2_R1179_U165, P2_U3080);
  nand ginst12677 (P2_R1179_U352, P2_R1179_U130, P2_R1179_U307);
  nand ginst12678 (P2_R1179_U353, P2_R1179_U41, P2_U3456);
  nand ginst12679 (P2_R1179_U354, P2_R1179_U40, P2_U3085);
  nand ginst12680 (P2_R1179_U355, P2_R1179_U150, P2_R1179_U217);
  nand ginst12681 (P2_R1179_U356, P2_R1179_U149, P2_R1179_U215);
  nand ginst12682 (P2_R1179_U357, P2_R1179_U39, P2_U3453);
  nand ginst12683 (P2_R1179_U358, P2_R1179_U36, P2_U3086);
  nand ginst12684 (P2_R1179_U359, P2_R1179_U39, P2_U3453);
  not ginst12685 (P2_R1179_U36, P2_U3453);
  nand ginst12686 (P2_R1179_U360, P2_R1179_U36, P2_U3086);
  nand ginst12687 (P2_R1179_U361, P2_R1179_U359, P2_R1179_U360);
  nand ginst12688 (P2_R1179_U362, P2_R1179_U37, P2_U3450);
  nand ginst12689 (P2_R1179_U363, P2_R1179_U21, P2_U3072);
  nand ginst12690 (P2_R1179_U364, P2_R1179_U222, P2_R1179_U42);
  nand ginst12691 (P2_R1179_U365, P2_R1179_U151, P2_R1179_U209);
  nand ginst12692 (P2_R1179_U366, P2_R1179_U32, P2_U3447);
  nand ginst12693 (P2_R1179_U367, P2_R1179_U30, P2_U3073);
  nand ginst12694 (P2_R1179_U368, P2_R1179_U366, P2_R1179_U367);
  nand ginst12695 (P2_R1179_U369, P2_R1179_U33, P2_U3444);
  not ginst12696 (P2_R1179_U37, P2_U3072);
  nand ginst12697 (P2_R1179_U370, P2_R1179_U22, P2_U3069);
  nand ginst12698 (P2_R1179_U371, P2_R1179_U232, P2_R1179_U43);
  nand ginst12699 (P2_R1179_U372, P2_R1179_U152, P2_R1179_U224);
  nand ginst12700 (P2_R1179_U373, P2_R1179_U34, P2_U3441);
  nand ginst12701 (P2_R1179_U374, P2_R1179_U31, P2_U3062);
  nand ginst12702 (P2_R1179_U375, P2_R1179_U154, P2_R1179_U233);
  nand ginst12703 (P2_R1179_U376, P2_R1179_U153, P2_R1179_U199);
  nand ginst12704 (P2_R1179_U377, P2_R1179_U29, P2_U3438);
  nand ginst12705 (P2_R1179_U378, P2_R1179_U26, P2_U3066);
  nand ginst12706 (P2_R1179_U379, P2_R1179_U29, P2_U3438);
  nand ginst12707 (P2_R1179_U38, P2_R1179_U21, P2_U3072);
  nand ginst12708 (P2_R1179_U380, P2_R1179_U26, P2_U3066);
  nand ginst12709 (P2_R1179_U381, P2_R1179_U379, P2_R1179_U380);
  nand ginst12710 (P2_R1179_U382, P2_R1179_U27, P2_U3435);
  nand ginst12711 (P2_R1179_U383, P2_R1179_U23, P2_U3070);
  nand ginst12712 (P2_R1179_U384, P2_R1179_U238, P2_R1179_U44);
  nand ginst12713 (P2_R1179_U385, P2_R1179_U155, P2_R1179_U193);
  nand ginst12714 (P2_R1179_U386, P2_R1179_U157, P2_U3960);
  nand ginst12715 (P2_R1179_U387, P2_R1179_U156, P2_U3057);
  nand ginst12716 (P2_R1179_U388, P2_R1179_U157, P2_U3960);
  nand ginst12717 (P2_R1179_U389, P2_R1179_U156, P2_U3057);
  not ginst12718 (P2_R1179_U39, P2_U3086);
  nand ginst12719 (P2_R1179_U390, P2_R1179_U388, P2_R1179_U389);
  nand ginst12720 (P2_R1179_U391, P2_R1179_U86, P2_U3949);
  nand ginst12721 (P2_R1179_U392, P2_R1179_U85, P2_U3056);
  not ginst12722 (P2_R1179_U393, P2_R1179_U131);
  nand ginst12723 (P2_R1179_U394, P2_R1179_U305, P2_R1179_U393);
  nand ginst12724 (P2_R1179_U395, P2_R1179_U131, P2_R1179_U87);
  nand ginst12725 (P2_R1179_U396, P2_R1179_U84, P2_U3950);
  nand ginst12726 (P2_R1179_U397, P2_R1179_U81, P2_U3055);
  nand ginst12727 (P2_R1179_U398, P2_R1179_U84, P2_U3950);
  nand ginst12728 (P2_R1179_U399, P2_R1179_U81, P2_U3055);
  not ginst12729 (P2_R1179_U40, P2_U3456);
  nand ginst12730 (P2_R1179_U400, P2_R1179_U398, P2_R1179_U399);
  nand ginst12731 (P2_R1179_U401, P2_R1179_U82, P2_U3951);
  nand ginst12732 (P2_R1179_U402, P2_R1179_U45, P2_U3059);
  nand ginst12733 (P2_R1179_U403, P2_R1179_U317, P2_R1179_U88);
  nand ginst12734 (P2_R1179_U404, P2_R1179_U158, P2_R1179_U299);
  nand ginst12735 (P2_R1179_U405, P2_R1179_U80, P2_U3952);
  nand ginst12736 (P2_R1179_U406, P2_R1179_U79, P2_U3060);
  not ginst12737 (P2_R1179_U407, P2_R1179_U134);
  nand ginst12738 (P2_R1179_U408, P2_R1179_U295, P2_R1179_U407);
  nand ginst12739 (P2_R1179_U409, P2_R1179_U134, P2_R1179_U159);
  not ginst12740 (P2_R1179_U41, P2_U3085);
  nand ginst12741 (P2_R1179_U410, P2_R1179_U78, P2_U3953);
  nand ginst12742 (P2_R1179_U411, P2_R1179_U77, P2_U3067);
  not ginst12743 (P2_R1179_U412, P2_R1179_U135);
  nand ginst12744 (P2_R1179_U413, P2_R1179_U291, P2_R1179_U412);
  nand ginst12745 (P2_R1179_U414, P2_R1179_U135, P2_R1179_U160);
  nand ginst12746 (P2_R1179_U415, P2_R1179_U73, P2_U3954);
  nand ginst12747 (P2_R1179_U416, P2_R1179_U70, P2_U3068);
  nand ginst12748 (P2_R1179_U417, P2_R1179_U415, P2_R1179_U416);
  nand ginst12749 (P2_R1179_U418, P2_R1179_U74, P2_U3955);
  nand ginst12750 (P2_R1179_U419, P2_R1179_U71, P2_U3063);
  nand ginst12751 (P2_R1179_U42, P2_R1179_U207, P2_R1179_U208);
  nand ginst12752 (P2_R1179_U420, P2_R1179_U327, P2_R1179_U89);
  nand ginst12753 (P2_R1179_U421, P2_R1179_U161, P2_R1179_U319);
  nand ginst12754 (P2_R1179_U422, P2_R1179_U75, P2_U3956);
  nand ginst12755 (P2_R1179_U423, P2_R1179_U72, P2_U3077);
  nand ginst12756 (P2_R1179_U424, P2_R1179_U163, P2_R1179_U328);
  nand ginst12757 (P2_R1179_U425, P2_R1179_U162, P2_R1179_U281);
  nand ginst12758 (P2_R1179_U426, P2_R1179_U69, P2_U3957);
  nand ginst12759 (P2_R1179_U427, P2_R1179_U68, P2_U3078);
  not ginst12760 (P2_R1179_U428, P2_R1179_U138);
  nand ginst12761 (P2_R1179_U429, P2_R1179_U277, P2_R1179_U428);
  nand ginst12762 (P2_R1179_U43, P2_R1179_U223, P2_R1179_U35);
  nand ginst12763 (P2_R1179_U430, P2_R1179_U138, P2_R1179_U164);
  nand ginst12764 (P2_R1179_U431, P2_R1179_U25, P2_U3432);
  nand ginst12765 (P2_R1179_U432, P2_R1179_U165, P2_U3080);
  not ginst12766 (P2_R1179_U433, P2_R1179_U139);
  nand ginst12767 (P2_R1179_U434, P2_R1179_U191, P2_R1179_U433);
  nand ginst12768 (P2_R1179_U435, P2_R1179_U139, P2_R1179_U166);
  nand ginst12769 (P2_R1179_U436, P2_R1179_U67, P2_U3485);
  nand ginst12770 (P2_R1179_U437, P2_R1179_U66, P2_U3083);
  not ginst12771 (P2_R1179_U438, P2_R1179_U140);
  nand ginst12772 (P2_R1179_U439, P2_R1179_U273, P2_R1179_U438);
  nand ginst12773 (P2_R1179_U44, P2_R1179_U176, P2_R1179_U192, P2_R1179_U351);
  nand ginst12774 (P2_R1179_U440, P2_R1179_U140, P2_R1179_U167);
  nand ginst12775 (P2_R1179_U441, P2_R1179_U65, P2_U3483);
  nand ginst12776 (P2_R1179_U442, P2_R1179_U168, P2_U3084);
  not ginst12777 (P2_R1179_U443, P2_R1179_U141);
  nand ginst12778 (P2_R1179_U444, P2_R1179_U269, P2_R1179_U443);
  nand ginst12779 (P2_R1179_U445, P2_R1179_U141, P2_R1179_U64);
  nand ginst12780 (P2_R1179_U446, P2_R1179_U63, P2_U3480);
  nand ginst12781 (P2_R1179_U447, P2_R1179_U62, P2_U3071);
  not ginst12782 (P2_R1179_U448, P2_R1179_U142);
  nand ginst12783 (P2_R1179_U449, P2_R1179_U265, P2_R1179_U448);
  not ginst12784 (P2_R1179_U45, P2_U3951);
  nand ginst12785 (P2_R1179_U450, P2_R1179_U142, P2_R1179_U169);
  nand ginst12786 (P2_R1179_U451, P2_R1179_U58, P2_U3477);
  nand ginst12787 (P2_R1179_U452, P2_R1179_U55, P2_U3075);
  nand ginst12788 (P2_R1179_U453, P2_R1179_U451, P2_R1179_U452);
  nand ginst12789 (P2_R1179_U454, P2_R1179_U59, P2_U3474);
  nand ginst12790 (P2_R1179_U455, P2_R1179_U56, P2_U3076);
  nand ginst12791 (P2_R1179_U456, P2_R1179_U338, P2_R1179_U90);
  nand ginst12792 (P2_R1179_U457, P2_R1179_U170, P2_R1179_U330);
  nand ginst12793 (P2_R1179_U458, P2_R1179_U60, P2_U3471);
  nand ginst12794 (P2_R1179_U459, P2_R1179_U57, P2_U3081);
  not ginst12795 (P2_R1179_U46, P2_U3459);
  nand ginst12796 (P2_R1179_U460, P2_R1179_U172, P2_R1179_U339);
  nand ginst12797 (P2_R1179_U461, P2_R1179_U171, P2_R1179_U255);
  nand ginst12798 (P2_R1179_U462, P2_R1179_U54, P2_U3468);
  nand ginst12799 (P2_R1179_U463, P2_R1179_U53, P2_U3082);
  not ginst12800 (P2_R1179_U464, P2_R1179_U145);
  nand ginst12801 (P2_R1179_U465, P2_R1179_U251, P2_R1179_U464);
  nand ginst12802 (P2_R1179_U466, P2_R1179_U145, P2_R1179_U173);
  nand ginst12803 (P2_R1179_U467, P2_R1179_U52, P2_U3465);
  nand ginst12804 (P2_R1179_U468, P2_R1179_U51, P2_U3074);
  not ginst12805 (P2_R1179_U469, P2_R1179_U146);
  not ginst12806 (P2_R1179_U47, P2_U3462);
  nand ginst12807 (P2_R1179_U470, P2_R1179_U247, P2_R1179_U469);
  nand ginst12808 (P2_R1179_U471, P2_R1179_U146, P2_R1179_U174);
  nand ginst12809 (P2_R1179_U472, P2_R1179_U48, P2_U3462);
  nand ginst12810 (P2_R1179_U473, P2_R1179_U47, P2_U3065);
  nand ginst12811 (P2_R1179_U474, P2_R1179_U472, P2_R1179_U473);
  nand ginst12812 (P2_R1179_U475, P2_R1179_U49, P2_U3459);
  nand ginst12813 (P2_R1179_U476, P2_R1179_U46, P2_U3064);
  nand ginst12814 (P2_R1179_U477, P2_R1179_U349, P2_R1179_U91);
  nand ginst12815 (P2_R1179_U478, P2_R1179_U175, P2_R1179_U341);
  not ginst12816 (P2_R1179_U48, P2_U3065);
  not ginst12817 (P2_R1179_U49, P2_U3064);
  nand ginst12818 (P2_R1179_U50, P2_R1179_U40, P2_U3085);
  not ginst12819 (P2_R1179_U51, P2_U3465);
  not ginst12820 (P2_R1179_U52, P2_U3074);
  not ginst12821 (P2_R1179_U53, P2_U3468);
  not ginst12822 (P2_R1179_U54, P2_U3082);
  not ginst12823 (P2_R1179_U55, P2_U3477);
  not ginst12824 (P2_R1179_U56, P2_U3474);
  not ginst12825 (P2_R1179_U57, P2_U3471);
  not ginst12826 (P2_R1179_U58, P2_U3075);
  not ginst12827 (P2_R1179_U59, P2_U3076);
  and ginst12828 (P2_R1179_U6, P2_R1179_U201, P2_R1179_U202);
  not ginst12829 (P2_R1179_U60, P2_U3081);
  nand ginst12830 (P2_R1179_U61, P2_R1179_U57, P2_U3081);
  not ginst12831 (P2_R1179_U62, P2_U3480);
  not ginst12832 (P2_R1179_U63, P2_U3071);
  nand ginst12833 (P2_R1179_U64, P2_R1179_U267, P2_R1179_U268);
  not ginst12834 (P2_R1179_U65, P2_U3084);
  not ginst12835 (P2_R1179_U66, P2_U3485);
  not ginst12836 (P2_R1179_U67, P2_U3083);
  not ginst12837 (P2_R1179_U68, P2_U3957);
  not ginst12838 (P2_R1179_U69, P2_U3078);
  and ginst12839 (P2_R1179_U7, P2_R1179_U240, P2_R1179_U241);
  not ginst12840 (P2_R1179_U70, P2_U3954);
  not ginst12841 (P2_R1179_U71, P2_U3955);
  not ginst12842 (P2_R1179_U72, P2_U3956);
  not ginst12843 (P2_R1179_U73, P2_U3068);
  not ginst12844 (P2_R1179_U74, P2_U3063);
  not ginst12845 (P2_R1179_U75, P2_U3077);
  nand ginst12846 (P2_R1179_U76, P2_R1179_U72, P2_U3077);
  not ginst12847 (P2_R1179_U77, P2_U3953);
  not ginst12848 (P2_R1179_U78, P2_U3067);
  not ginst12849 (P2_R1179_U79, P2_U3952);
  and ginst12850 (P2_R1179_U8, P2_R1179_U181, P2_R1179_U256);
  not ginst12851 (P2_R1179_U80, P2_U3060);
  not ginst12852 (P2_R1179_U81, P2_U3950);
  not ginst12853 (P2_R1179_U82, P2_U3059);
  nand ginst12854 (P2_R1179_U83, P2_R1179_U45, P2_U3059);
  not ginst12855 (P2_R1179_U84, P2_U3055);
  not ginst12856 (P2_R1179_U85, P2_U3949);
  not ginst12857 (P2_R1179_U86, P2_U3056);
  nand ginst12858 (P2_R1179_U87, P2_R1179_U128, P2_R1179_U301);
  nand ginst12859 (P2_R1179_U88, P2_R1179_U297, P2_R1179_U298);
  nand ginst12860 (P2_R1179_U89, P2_R1179_U318, P2_R1179_U76);
  and ginst12861 (P2_R1179_U9, P2_R1179_U257, P2_R1179_U258);
  nand ginst12862 (P2_R1179_U90, P2_R1179_U329, P2_R1179_U61);
  nand ginst12863 (P2_R1179_U91, P2_R1179_U340, P2_R1179_U50);
  not ginst12864 (P2_R1179_U92, P2_U3079);
  nand ginst12865 (P2_R1179_U93, P2_R1179_U394, P2_R1179_U395);
  nand ginst12866 (P2_R1179_U94, P2_R1179_U408, P2_R1179_U409);
  nand ginst12867 (P2_R1179_U95, P2_R1179_U413, P2_R1179_U414);
  nand ginst12868 (P2_R1179_U96, P2_R1179_U429, P2_R1179_U430);
  nand ginst12869 (P2_R1179_U97, P2_R1179_U434, P2_R1179_U435);
  nand ginst12870 (P2_R1179_U98, P2_R1179_U439, P2_R1179_U440);
  nand ginst12871 (P2_R1179_U99, P2_R1179_U444, P2_R1179_U445);
  and ginst12872 (P2_R1203_U10, P2_R1203_U182, P2_R1203_U282);
  nand ginst12873 (P2_R1203_U100, P2_R1203_U449, P2_R1203_U450);
  nand ginst12874 (P2_R1203_U101, P2_R1203_U465, P2_R1203_U466);
  nand ginst12875 (P2_R1203_U102, P2_R1203_U470, P2_R1203_U471);
  nand ginst12876 (P2_R1203_U103, P2_R1203_U355, P2_R1203_U356);
  nand ginst12877 (P2_R1203_U104, P2_R1203_U364, P2_R1203_U365);
  nand ginst12878 (P2_R1203_U105, P2_R1203_U371, P2_R1203_U372);
  nand ginst12879 (P2_R1203_U106, P2_R1203_U375, P2_R1203_U376);
  nand ginst12880 (P2_R1203_U107, P2_R1203_U384, P2_R1203_U385);
  nand ginst12881 (P2_R1203_U108, P2_R1203_U403, P2_R1203_U404);
  nand ginst12882 (P2_R1203_U109, P2_R1203_U420, P2_R1203_U421);
  and ginst12883 (P2_R1203_U11, P2_R1203_U283, P2_R1203_U284);
  nand ginst12884 (P2_R1203_U110, P2_R1203_U424, P2_R1203_U425);
  nand ginst12885 (P2_R1203_U111, P2_R1203_U456, P2_R1203_U457);
  nand ginst12886 (P2_R1203_U112, P2_R1203_U460, P2_R1203_U461);
  nand ginst12887 (P2_R1203_U113, P2_R1203_U477, P2_R1203_U478);
  and ginst12888 (P2_R1203_U114, P2_R1203_U184, P2_R1203_U194);
  and ginst12889 (P2_R1203_U115, P2_R1203_U197, P2_R1203_U198);
  and ginst12890 (P2_R1203_U116, P2_R1203_U185, P2_R1203_U200, P2_R1203_U205);
  and ginst12891 (P2_R1203_U117, P2_R1203_U186, P2_R1203_U210);
  and ginst12892 (P2_R1203_U118, P2_R1203_U213, P2_R1203_U214);
  and ginst12893 (P2_R1203_U119, P2_R1203_U357, P2_R1203_U358, P2_R1203_U38);
  nand ginst12894 (P2_R1203_U12, P2_R1203_U344, P2_R1203_U347);
  and ginst12895 (P2_R1203_U120, P2_R1203_U186, P2_R1203_U361);
  and ginst12896 (P2_R1203_U121, P2_R1203_U229, P2_R1203_U6);
  and ginst12897 (P2_R1203_U122, P2_R1203_U185, P2_R1203_U368);
  and ginst12898 (P2_R1203_U123, P2_R1203_U28, P2_R1203_U377, P2_R1203_U378);
  and ginst12899 (P2_R1203_U124, P2_R1203_U184, P2_R1203_U381);
  and ginst12900 (P2_R1203_U125, P2_R1203_U180, P2_R1203_U216, P2_R1203_U239);
  and ginst12901 (P2_R1203_U126, P2_R1203_U261, P2_R1203_U8);
  and ginst12902 (P2_R1203_U127, P2_R1203_U10, P2_R1203_U287);
  and ginst12903 (P2_R1203_U128, P2_R1203_U303, P2_R1203_U304);
  and ginst12904 (P2_R1203_U129, P2_R1203_U311, P2_R1203_U386, P2_R1203_U387);
  nand ginst12905 (P2_R1203_U13, P2_R1203_U333, P2_R1203_U336);
  and ginst12906 (P2_R1203_U130, P2_R1203_U308, P2_R1203_U390);
  nand ginst12907 (P2_R1203_U131, P2_R1203_U391, P2_R1203_U392);
  and ginst12908 (P2_R1203_U132, P2_R1203_U396, P2_R1203_U397, P2_R1203_U83);
  and ginst12909 (P2_R1203_U133, P2_R1203_U183, P2_R1203_U400);
  nand ginst12910 (P2_R1203_U134, P2_R1203_U405, P2_R1203_U406);
  nand ginst12911 (P2_R1203_U135, P2_R1203_U410, P2_R1203_U411);
  and ginst12912 (P2_R1203_U136, P2_R1203_U11, P2_R1203_U324);
  and ginst12913 (P2_R1203_U137, P2_R1203_U182, P2_R1203_U417);
  nand ginst12914 (P2_R1203_U138, P2_R1203_U426, P2_R1203_U427);
  nand ginst12915 (P2_R1203_U139, P2_R1203_U431, P2_R1203_U432);
  nand ginst12916 (P2_R1203_U14, P2_R1203_U322, P2_R1203_U325);
  nand ginst12917 (P2_R1203_U140, P2_R1203_U436, P2_R1203_U437);
  nand ginst12918 (P2_R1203_U141, P2_R1203_U441, P2_R1203_U442);
  nand ginst12919 (P2_R1203_U142, P2_R1203_U446, P2_R1203_U447);
  and ginst12920 (P2_R1203_U143, P2_R1203_U335, P2_R1203_U9);
  and ginst12921 (P2_R1203_U144, P2_R1203_U181, P2_R1203_U453);
  nand ginst12922 (P2_R1203_U145, P2_R1203_U462, P2_R1203_U463);
  nand ginst12923 (P2_R1203_U146, P2_R1203_U467, P2_R1203_U468);
  and ginst12924 (P2_R1203_U147, P2_R1203_U346, P2_R1203_U7);
  and ginst12925 (P2_R1203_U148, P2_R1203_U180, P2_R1203_U474);
  and ginst12926 (P2_R1203_U149, P2_R1203_U353, P2_R1203_U354);
  nand ginst12927 (P2_R1203_U15, P2_R1203_U314, P2_R1203_U316);
  nand ginst12928 (P2_R1203_U150, P2_R1203_U118, P2_R1203_U211);
  and ginst12929 (P2_R1203_U151, P2_R1203_U362, P2_R1203_U363);
  and ginst12930 (P2_R1203_U152, P2_R1203_U369, P2_R1203_U370);
  and ginst12931 (P2_R1203_U153, P2_R1203_U373, P2_R1203_U374);
  nand ginst12932 (P2_R1203_U154, P2_R1203_U115, P2_R1203_U195);
  and ginst12933 (P2_R1203_U155, P2_R1203_U382, P2_R1203_U383);
  not ginst12934 (P2_R1203_U156, P2_U3960);
  not ginst12935 (P2_R1203_U157, P2_U3057);
  and ginst12936 (P2_R1203_U158, P2_R1203_U401, P2_R1203_U402);
  nand ginst12937 (P2_R1203_U159, P2_R1203_U293, P2_R1203_U294);
  nand ginst12938 (P2_R1203_U16, P2_R1203_U312, P2_R1203_U352);
  nand ginst12939 (P2_R1203_U160, P2_R1203_U289, P2_R1203_U290);
  and ginst12940 (P2_R1203_U161, P2_R1203_U418, P2_R1203_U419);
  and ginst12941 (P2_R1203_U162, P2_R1203_U422, P2_R1203_U423);
  nand ginst12942 (P2_R1203_U163, P2_R1203_U279, P2_R1203_U280);
  nand ginst12943 (P2_R1203_U164, P2_R1203_U275, P2_R1203_U276);
  not ginst12944 (P2_R1203_U165, P2_U3432);
  nand ginst12945 (P2_R1203_U166, P2_R1203_U92, P2_U3427);
  nand ginst12946 (P2_R1203_U167, P2_R1203_U271, P2_R1203_U272);
  not ginst12947 (P2_R1203_U168, P2_U3483);
  nand ginst12948 (P2_R1203_U169, P2_R1203_U263, P2_R1203_U264);
  nand ginst12949 (P2_R1203_U17, P2_R1203_U235, P2_R1203_U237);
  and ginst12950 (P2_R1203_U170, P2_R1203_U454, P2_R1203_U455);
  and ginst12951 (P2_R1203_U171, P2_R1203_U458, P2_R1203_U459);
  nand ginst12952 (P2_R1203_U172, P2_R1203_U253, P2_R1203_U254);
  nand ginst12953 (P2_R1203_U173, P2_R1203_U249, P2_R1203_U250);
  nand ginst12954 (P2_R1203_U174, P2_R1203_U245, P2_R1203_U246);
  and ginst12955 (P2_R1203_U175, P2_R1203_U475, P2_R1203_U476);
  nand ginst12956 (P2_R1203_U176, P2_R1203_U165, P2_R1203_U166);
  not ginst12957 (P2_R1203_U177, P2_R1203_U83);
  not ginst12958 (P2_R1203_U178, P2_R1203_U28);
  not ginst12959 (P2_R1203_U179, P2_R1203_U38);
  nand ginst12960 (P2_R1203_U18, P2_R1203_U227, P2_R1203_U230);
  nand ginst12961 (P2_R1203_U180, P2_R1203_U49, P2_U3459);
  nand ginst12962 (P2_R1203_U181, P2_R1203_U59, P2_U3474);
  nand ginst12963 (P2_R1203_U182, P2_R1203_U74, P2_U3955);
  nand ginst12964 (P2_R1203_U183, P2_R1203_U82, P2_U3951);
  nand ginst12965 (P2_R1203_U184, P2_R1203_U27, P2_U3435);
  nand ginst12966 (P2_R1203_U185, P2_R1203_U33, P2_U3444);
  nand ginst12967 (P2_R1203_U186, P2_R1203_U37, P2_U3450);
  not ginst12968 (P2_R1203_U187, P2_R1203_U61);
  not ginst12969 (P2_R1203_U188, P2_R1203_U76);
  not ginst12970 (P2_R1203_U189, P2_R1203_U35);
  nand ginst12971 (P2_R1203_U19, P2_R1203_U219, P2_R1203_U221);
  not ginst12972 (P2_R1203_U190, P2_R1203_U50);
  not ginst12973 (P2_R1203_U191, P2_R1203_U166);
  nand ginst12974 (P2_R1203_U192, P2_R1203_U166, P2_U3080);
  not ginst12975 (P2_R1203_U193, P2_R1203_U44);
  nand ginst12976 (P2_R1203_U194, P2_R1203_U29, P2_U3438);
  nand ginst12977 (P2_R1203_U195, P2_R1203_U114, P2_R1203_U44);
  nand ginst12978 (P2_R1203_U196, P2_R1203_U28, P2_R1203_U29);
  nand ginst12979 (P2_R1203_U197, P2_R1203_U196, P2_R1203_U26);
  nand ginst12980 (P2_R1203_U198, P2_R1203_U178, P2_U3066);
  not ginst12981 (P2_R1203_U199, P2_R1203_U154);
  nand ginst12982 (P2_R1203_U20, P2_R1203_U166, P2_R1203_U350);
  nand ginst12983 (P2_R1203_U200, P2_R1203_U32, P2_U3447);
  nand ginst12984 (P2_R1203_U201, P2_R1203_U30, P2_U3073);
  nand ginst12985 (P2_R1203_U202, P2_R1203_U22, P2_U3069);
  nand ginst12986 (P2_R1203_U203, P2_R1203_U185, P2_R1203_U189);
  nand ginst12987 (P2_R1203_U204, P2_R1203_U203, P2_R1203_U6);
  nand ginst12988 (P2_R1203_U205, P2_R1203_U34, P2_U3441);
  nand ginst12989 (P2_R1203_U206, P2_R1203_U32, P2_U3447);
  nand ginst12990 (P2_R1203_U207, P2_R1203_U116, P2_R1203_U154);
  nand ginst12991 (P2_R1203_U208, P2_R1203_U204, P2_R1203_U206);
  not ginst12992 (P2_R1203_U209, P2_R1203_U42);
  not ginst12993 (P2_R1203_U21, P2_U3450);
  nand ginst12994 (P2_R1203_U210, P2_R1203_U39, P2_U3453);
  nand ginst12995 (P2_R1203_U211, P2_R1203_U117, P2_R1203_U42);
  nand ginst12996 (P2_R1203_U212, P2_R1203_U38, P2_R1203_U39);
  nand ginst12997 (P2_R1203_U213, P2_R1203_U212, P2_R1203_U36);
  nand ginst12998 (P2_R1203_U214, P2_R1203_U179, P2_U3086);
  not ginst12999 (P2_R1203_U215, P2_R1203_U150);
  nand ginst13000 (P2_R1203_U216, P2_R1203_U41, P2_U3456);
  nand ginst13001 (P2_R1203_U217, P2_R1203_U216, P2_R1203_U50);
  nand ginst13002 (P2_R1203_U218, P2_R1203_U209, P2_R1203_U38);
  nand ginst13003 (P2_R1203_U219, P2_R1203_U120, P2_R1203_U218);
  not ginst13004 (P2_R1203_U22, P2_U3444);
  nand ginst13005 (P2_R1203_U220, P2_R1203_U186, P2_R1203_U42);
  nand ginst13006 (P2_R1203_U221, P2_R1203_U119, P2_R1203_U220);
  nand ginst13007 (P2_R1203_U222, P2_R1203_U186, P2_R1203_U38);
  nand ginst13008 (P2_R1203_U223, P2_R1203_U154, P2_R1203_U205);
  not ginst13009 (P2_R1203_U224, P2_R1203_U43);
  nand ginst13010 (P2_R1203_U225, P2_R1203_U22, P2_U3069);
  nand ginst13011 (P2_R1203_U226, P2_R1203_U224, P2_R1203_U225);
  nand ginst13012 (P2_R1203_U227, P2_R1203_U122, P2_R1203_U226);
  nand ginst13013 (P2_R1203_U228, P2_R1203_U185, P2_R1203_U43);
  nand ginst13014 (P2_R1203_U229, P2_R1203_U32, P2_U3447);
  not ginst13015 (P2_R1203_U23, P2_U3435);
  nand ginst13016 (P2_R1203_U230, P2_R1203_U121, P2_R1203_U228);
  nand ginst13017 (P2_R1203_U231, P2_R1203_U22, P2_U3069);
  nand ginst13018 (P2_R1203_U232, P2_R1203_U185, P2_R1203_U231);
  nand ginst13019 (P2_R1203_U233, P2_R1203_U205, P2_R1203_U35);
  nand ginst13020 (P2_R1203_U234, P2_R1203_U193, P2_R1203_U28);
  nand ginst13021 (P2_R1203_U235, P2_R1203_U124, P2_R1203_U234);
  nand ginst13022 (P2_R1203_U236, P2_R1203_U184, P2_R1203_U44);
  nand ginst13023 (P2_R1203_U237, P2_R1203_U123, P2_R1203_U236);
  nand ginst13024 (P2_R1203_U238, P2_R1203_U184, P2_R1203_U28);
  nand ginst13025 (P2_R1203_U239, P2_R1203_U48, P2_U3462);
  not ginst13026 (P2_R1203_U24, P2_U3427);
  nand ginst13027 (P2_R1203_U240, P2_R1203_U47, P2_U3065);
  nand ginst13028 (P2_R1203_U241, P2_R1203_U46, P2_U3064);
  nand ginst13029 (P2_R1203_U242, P2_R1203_U180, P2_R1203_U190);
  nand ginst13030 (P2_R1203_U243, P2_R1203_U242, P2_R1203_U7);
  nand ginst13031 (P2_R1203_U244, P2_R1203_U48, P2_U3462);
  nand ginst13032 (P2_R1203_U245, P2_R1203_U125, P2_R1203_U150);
  nand ginst13033 (P2_R1203_U246, P2_R1203_U243, P2_R1203_U244);
  not ginst13034 (P2_R1203_U247, P2_R1203_U174);
  nand ginst13035 (P2_R1203_U248, P2_R1203_U52, P2_U3465);
  nand ginst13036 (P2_R1203_U249, P2_R1203_U174, P2_R1203_U248);
  not ginst13037 (P2_R1203_U25, P2_U3080);
  nand ginst13038 (P2_R1203_U250, P2_R1203_U51, P2_U3074);
  not ginst13039 (P2_R1203_U251, P2_R1203_U173);
  nand ginst13040 (P2_R1203_U252, P2_R1203_U54, P2_U3468);
  nand ginst13041 (P2_R1203_U253, P2_R1203_U173, P2_R1203_U252);
  nand ginst13042 (P2_R1203_U254, P2_R1203_U53, P2_U3082);
  not ginst13043 (P2_R1203_U255, P2_R1203_U172);
  nand ginst13044 (P2_R1203_U256, P2_R1203_U58, P2_U3477);
  nand ginst13045 (P2_R1203_U257, P2_R1203_U55, P2_U3075);
  nand ginst13046 (P2_R1203_U258, P2_R1203_U56, P2_U3076);
  nand ginst13047 (P2_R1203_U259, P2_R1203_U187, P2_R1203_U8);
  not ginst13048 (P2_R1203_U26, P2_U3438);
  nand ginst13049 (P2_R1203_U260, P2_R1203_U259, P2_R1203_U9);
  nand ginst13050 (P2_R1203_U261, P2_R1203_U60, P2_U3471);
  nand ginst13051 (P2_R1203_U262, P2_R1203_U58, P2_U3477);
  nand ginst13052 (P2_R1203_U263, P2_R1203_U126, P2_R1203_U172);
  nand ginst13053 (P2_R1203_U264, P2_R1203_U260, P2_R1203_U262);
  not ginst13054 (P2_R1203_U265, P2_R1203_U169);
  nand ginst13055 (P2_R1203_U266, P2_R1203_U63, P2_U3480);
  nand ginst13056 (P2_R1203_U267, P2_R1203_U169, P2_R1203_U266);
  nand ginst13057 (P2_R1203_U268, P2_R1203_U62, P2_U3071);
  not ginst13058 (P2_R1203_U269, P2_R1203_U64);
  not ginst13059 (P2_R1203_U27, P2_U3070);
  nand ginst13060 (P2_R1203_U270, P2_R1203_U269, P2_R1203_U65);
  nand ginst13061 (P2_R1203_U271, P2_R1203_U168, P2_R1203_U270);
  nand ginst13062 (P2_R1203_U272, P2_R1203_U64, P2_U3084);
  not ginst13063 (P2_R1203_U273, P2_R1203_U167);
  nand ginst13064 (P2_R1203_U274, P2_R1203_U67, P2_U3485);
  nand ginst13065 (P2_R1203_U275, P2_R1203_U167, P2_R1203_U274);
  nand ginst13066 (P2_R1203_U276, P2_R1203_U66, P2_U3083);
  not ginst13067 (P2_R1203_U277, P2_R1203_U164);
  nand ginst13068 (P2_R1203_U278, P2_R1203_U69, P2_U3957);
  nand ginst13069 (P2_R1203_U279, P2_R1203_U164, P2_R1203_U278);
  nand ginst13070 (P2_R1203_U28, P2_R1203_U23, P2_U3070);
  nand ginst13071 (P2_R1203_U280, P2_R1203_U68, P2_U3078);
  not ginst13072 (P2_R1203_U281, P2_R1203_U163);
  nand ginst13073 (P2_R1203_U282, P2_R1203_U73, P2_U3954);
  nand ginst13074 (P2_R1203_U283, P2_R1203_U70, P2_U3068);
  nand ginst13075 (P2_R1203_U284, P2_R1203_U71, P2_U3063);
  nand ginst13076 (P2_R1203_U285, P2_R1203_U10, P2_R1203_U188);
  nand ginst13077 (P2_R1203_U286, P2_R1203_U11, P2_R1203_U285);
  nand ginst13078 (P2_R1203_U287, P2_R1203_U75, P2_U3956);
  nand ginst13079 (P2_R1203_U288, P2_R1203_U73, P2_U3954);
  nand ginst13080 (P2_R1203_U289, P2_R1203_U127, P2_R1203_U163);
  not ginst13081 (P2_R1203_U29, P2_U3066);
  nand ginst13082 (P2_R1203_U290, P2_R1203_U286, P2_R1203_U288);
  not ginst13083 (P2_R1203_U291, P2_R1203_U160);
  nand ginst13084 (P2_R1203_U292, P2_R1203_U78, P2_U3953);
  nand ginst13085 (P2_R1203_U293, P2_R1203_U160, P2_R1203_U292);
  nand ginst13086 (P2_R1203_U294, P2_R1203_U77, P2_U3067);
  not ginst13087 (P2_R1203_U295, P2_R1203_U159);
  nand ginst13088 (P2_R1203_U296, P2_R1203_U80, P2_U3952);
  nand ginst13089 (P2_R1203_U297, P2_R1203_U159, P2_R1203_U296);
  nand ginst13090 (P2_R1203_U298, P2_R1203_U79, P2_U3060);
  not ginst13091 (P2_R1203_U299, P2_R1203_U88);
  not ginst13092 (P2_R1203_U30, P2_U3447);
  nand ginst13093 (P2_R1203_U300, P2_R1203_U84, P2_U3950);
  nand ginst13094 (P2_R1203_U301, P2_R1203_U183, P2_R1203_U300, P2_R1203_U88);
  nand ginst13095 (P2_R1203_U302, P2_R1203_U83, P2_R1203_U84);
  nand ginst13096 (P2_R1203_U303, P2_R1203_U302, P2_R1203_U81);
  nand ginst13097 (P2_R1203_U304, P2_R1203_U177, P2_U3055);
  not ginst13098 (P2_R1203_U305, P2_R1203_U87);
  nand ginst13099 (P2_R1203_U306, P2_R1203_U85, P2_U3056);
  nand ginst13100 (P2_R1203_U307, P2_R1203_U305, P2_R1203_U306);
  nand ginst13101 (P2_R1203_U308, P2_R1203_U86, P2_U3949);
  nand ginst13102 (P2_R1203_U309, P2_R1203_U86, P2_U3949);
  not ginst13103 (P2_R1203_U31, P2_U3441);
  nand ginst13104 (P2_R1203_U310, P2_R1203_U309, P2_R1203_U87);
  nand ginst13105 (P2_R1203_U311, P2_R1203_U85, P2_U3056);
  nand ginst13106 (P2_R1203_U312, P2_R1203_U129, P2_R1203_U310);
  nand ginst13107 (P2_R1203_U313, P2_R1203_U299, P2_R1203_U83);
  nand ginst13108 (P2_R1203_U314, P2_R1203_U133, P2_R1203_U313);
  nand ginst13109 (P2_R1203_U315, P2_R1203_U183, P2_R1203_U88);
  nand ginst13110 (P2_R1203_U316, P2_R1203_U132, P2_R1203_U315);
  nand ginst13111 (P2_R1203_U317, P2_R1203_U183, P2_R1203_U83);
  nand ginst13112 (P2_R1203_U318, P2_R1203_U163, P2_R1203_U287);
  not ginst13113 (P2_R1203_U319, P2_R1203_U89);
  not ginst13114 (P2_R1203_U32, P2_U3073);
  nand ginst13115 (P2_R1203_U320, P2_R1203_U71, P2_U3063);
  nand ginst13116 (P2_R1203_U321, P2_R1203_U319, P2_R1203_U320);
  nand ginst13117 (P2_R1203_U322, P2_R1203_U137, P2_R1203_U321);
  nand ginst13118 (P2_R1203_U323, P2_R1203_U182, P2_R1203_U89);
  nand ginst13119 (P2_R1203_U324, P2_R1203_U73, P2_U3954);
  nand ginst13120 (P2_R1203_U325, P2_R1203_U136, P2_R1203_U323);
  nand ginst13121 (P2_R1203_U326, P2_R1203_U71, P2_U3063);
  nand ginst13122 (P2_R1203_U327, P2_R1203_U182, P2_R1203_U326);
  nand ginst13123 (P2_R1203_U328, P2_R1203_U287, P2_R1203_U76);
  nand ginst13124 (P2_R1203_U329, P2_R1203_U172, P2_R1203_U261);
  not ginst13125 (P2_R1203_U33, P2_U3069);
  not ginst13126 (P2_R1203_U330, P2_R1203_U90);
  nand ginst13127 (P2_R1203_U331, P2_R1203_U56, P2_U3076);
  nand ginst13128 (P2_R1203_U332, P2_R1203_U330, P2_R1203_U331);
  nand ginst13129 (P2_R1203_U333, P2_R1203_U144, P2_R1203_U332);
  nand ginst13130 (P2_R1203_U334, P2_R1203_U181, P2_R1203_U90);
  nand ginst13131 (P2_R1203_U335, P2_R1203_U58, P2_U3477);
  nand ginst13132 (P2_R1203_U336, P2_R1203_U143, P2_R1203_U334);
  nand ginst13133 (P2_R1203_U337, P2_R1203_U56, P2_U3076);
  nand ginst13134 (P2_R1203_U338, P2_R1203_U181, P2_R1203_U337);
  nand ginst13135 (P2_R1203_U339, P2_R1203_U261, P2_R1203_U61);
  not ginst13136 (P2_R1203_U34, P2_U3062);
  nand ginst13137 (P2_R1203_U340, P2_R1203_U150, P2_R1203_U216);
  not ginst13138 (P2_R1203_U341, P2_R1203_U91);
  nand ginst13139 (P2_R1203_U342, P2_R1203_U46, P2_U3064);
  nand ginst13140 (P2_R1203_U343, P2_R1203_U341, P2_R1203_U342);
  nand ginst13141 (P2_R1203_U344, P2_R1203_U148, P2_R1203_U343);
  nand ginst13142 (P2_R1203_U345, P2_R1203_U180, P2_R1203_U91);
  nand ginst13143 (P2_R1203_U346, P2_R1203_U48, P2_U3462);
  nand ginst13144 (P2_R1203_U347, P2_R1203_U147, P2_R1203_U345);
  nand ginst13145 (P2_R1203_U348, P2_R1203_U46, P2_U3064);
  nand ginst13146 (P2_R1203_U349, P2_R1203_U180, P2_R1203_U348);
  nand ginst13147 (P2_R1203_U35, P2_R1203_U31, P2_U3062);
  nand ginst13148 (P2_R1203_U350, P2_R1203_U24, P2_U3079);
  nand ginst13149 (P2_R1203_U351, P2_R1203_U165, P2_U3080);
  nand ginst13150 (P2_R1203_U352, P2_R1203_U130, P2_R1203_U307);
  nand ginst13151 (P2_R1203_U353, P2_R1203_U41, P2_U3456);
  nand ginst13152 (P2_R1203_U354, P2_R1203_U40, P2_U3085);
  nand ginst13153 (P2_R1203_U355, P2_R1203_U150, P2_R1203_U217);
  nand ginst13154 (P2_R1203_U356, P2_R1203_U149, P2_R1203_U215);
  nand ginst13155 (P2_R1203_U357, P2_R1203_U39, P2_U3453);
  nand ginst13156 (P2_R1203_U358, P2_R1203_U36, P2_U3086);
  nand ginst13157 (P2_R1203_U359, P2_R1203_U39, P2_U3453);
  not ginst13158 (P2_R1203_U36, P2_U3453);
  nand ginst13159 (P2_R1203_U360, P2_R1203_U36, P2_U3086);
  nand ginst13160 (P2_R1203_U361, P2_R1203_U359, P2_R1203_U360);
  nand ginst13161 (P2_R1203_U362, P2_R1203_U37, P2_U3450);
  nand ginst13162 (P2_R1203_U363, P2_R1203_U21, P2_U3072);
  nand ginst13163 (P2_R1203_U364, P2_R1203_U222, P2_R1203_U42);
  nand ginst13164 (P2_R1203_U365, P2_R1203_U151, P2_R1203_U209);
  nand ginst13165 (P2_R1203_U366, P2_R1203_U32, P2_U3447);
  nand ginst13166 (P2_R1203_U367, P2_R1203_U30, P2_U3073);
  nand ginst13167 (P2_R1203_U368, P2_R1203_U366, P2_R1203_U367);
  nand ginst13168 (P2_R1203_U369, P2_R1203_U33, P2_U3444);
  not ginst13169 (P2_R1203_U37, P2_U3072);
  nand ginst13170 (P2_R1203_U370, P2_R1203_U22, P2_U3069);
  nand ginst13171 (P2_R1203_U371, P2_R1203_U232, P2_R1203_U43);
  nand ginst13172 (P2_R1203_U372, P2_R1203_U152, P2_R1203_U224);
  nand ginst13173 (P2_R1203_U373, P2_R1203_U34, P2_U3441);
  nand ginst13174 (P2_R1203_U374, P2_R1203_U31, P2_U3062);
  nand ginst13175 (P2_R1203_U375, P2_R1203_U154, P2_R1203_U233);
  nand ginst13176 (P2_R1203_U376, P2_R1203_U153, P2_R1203_U199);
  nand ginst13177 (P2_R1203_U377, P2_R1203_U29, P2_U3438);
  nand ginst13178 (P2_R1203_U378, P2_R1203_U26, P2_U3066);
  nand ginst13179 (P2_R1203_U379, P2_R1203_U29, P2_U3438);
  nand ginst13180 (P2_R1203_U38, P2_R1203_U21, P2_U3072);
  nand ginst13181 (P2_R1203_U380, P2_R1203_U26, P2_U3066);
  nand ginst13182 (P2_R1203_U381, P2_R1203_U379, P2_R1203_U380);
  nand ginst13183 (P2_R1203_U382, P2_R1203_U27, P2_U3435);
  nand ginst13184 (P2_R1203_U383, P2_R1203_U23, P2_U3070);
  nand ginst13185 (P2_R1203_U384, P2_R1203_U238, P2_R1203_U44);
  nand ginst13186 (P2_R1203_U385, P2_R1203_U155, P2_R1203_U193);
  nand ginst13187 (P2_R1203_U386, P2_R1203_U157, P2_U3960);
  nand ginst13188 (P2_R1203_U387, P2_R1203_U156, P2_U3057);
  nand ginst13189 (P2_R1203_U388, P2_R1203_U157, P2_U3960);
  nand ginst13190 (P2_R1203_U389, P2_R1203_U156, P2_U3057);
  not ginst13191 (P2_R1203_U39, P2_U3086);
  nand ginst13192 (P2_R1203_U390, P2_R1203_U388, P2_R1203_U389);
  nand ginst13193 (P2_R1203_U391, P2_R1203_U86, P2_U3949);
  nand ginst13194 (P2_R1203_U392, P2_R1203_U85, P2_U3056);
  not ginst13195 (P2_R1203_U393, P2_R1203_U131);
  nand ginst13196 (P2_R1203_U394, P2_R1203_U305, P2_R1203_U393);
  nand ginst13197 (P2_R1203_U395, P2_R1203_U131, P2_R1203_U87);
  nand ginst13198 (P2_R1203_U396, P2_R1203_U84, P2_U3950);
  nand ginst13199 (P2_R1203_U397, P2_R1203_U81, P2_U3055);
  nand ginst13200 (P2_R1203_U398, P2_R1203_U84, P2_U3950);
  nand ginst13201 (P2_R1203_U399, P2_R1203_U81, P2_U3055);
  not ginst13202 (P2_R1203_U40, P2_U3456);
  nand ginst13203 (P2_R1203_U400, P2_R1203_U398, P2_R1203_U399);
  nand ginst13204 (P2_R1203_U401, P2_R1203_U82, P2_U3951);
  nand ginst13205 (P2_R1203_U402, P2_R1203_U45, P2_U3059);
  nand ginst13206 (P2_R1203_U403, P2_R1203_U317, P2_R1203_U88);
  nand ginst13207 (P2_R1203_U404, P2_R1203_U158, P2_R1203_U299);
  nand ginst13208 (P2_R1203_U405, P2_R1203_U80, P2_U3952);
  nand ginst13209 (P2_R1203_U406, P2_R1203_U79, P2_U3060);
  not ginst13210 (P2_R1203_U407, P2_R1203_U134);
  nand ginst13211 (P2_R1203_U408, P2_R1203_U295, P2_R1203_U407);
  nand ginst13212 (P2_R1203_U409, P2_R1203_U134, P2_R1203_U159);
  not ginst13213 (P2_R1203_U41, P2_U3085);
  nand ginst13214 (P2_R1203_U410, P2_R1203_U78, P2_U3953);
  nand ginst13215 (P2_R1203_U411, P2_R1203_U77, P2_U3067);
  not ginst13216 (P2_R1203_U412, P2_R1203_U135);
  nand ginst13217 (P2_R1203_U413, P2_R1203_U291, P2_R1203_U412);
  nand ginst13218 (P2_R1203_U414, P2_R1203_U135, P2_R1203_U160);
  nand ginst13219 (P2_R1203_U415, P2_R1203_U73, P2_U3954);
  nand ginst13220 (P2_R1203_U416, P2_R1203_U70, P2_U3068);
  nand ginst13221 (P2_R1203_U417, P2_R1203_U415, P2_R1203_U416);
  nand ginst13222 (P2_R1203_U418, P2_R1203_U74, P2_U3955);
  nand ginst13223 (P2_R1203_U419, P2_R1203_U71, P2_U3063);
  nand ginst13224 (P2_R1203_U42, P2_R1203_U207, P2_R1203_U208);
  nand ginst13225 (P2_R1203_U420, P2_R1203_U327, P2_R1203_U89);
  nand ginst13226 (P2_R1203_U421, P2_R1203_U161, P2_R1203_U319);
  nand ginst13227 (P2_R1203_U422, P2_R1203_U75, P2_U3956);
  nand ginst13228 (P2_R1203_U423, P2_R1203_U72, P2_U3077);
  nand ginst13229 (P2_R1203_U424, P2_R1203_U163, P2_R1203_U328);
  nand ginst13230 (P2_R1203_U425, P2_R1203_U162, P2_R1203_U281);
  nand ginst13231 (P2_R1203_U426, P2_R1203_U69, P2_U3957);
  nand ginst13232 (P2_R1203_U427, P2_R1203_U68, P2_U3078);
  not ginst13233 (P2_R1203_U428, P2_R1203_U138);
  nand ginst13234 (P2_R1203_U429, P2_R1203_U277, P2_R1203_U428);
  nand ginst13235 (P2_R1203_U43, P2_R1203_U223, P2_R1203_U35);
  nand ginst13236 (P2_R1203_U430, P2_R1203_U138, P2_R1203_U164);
  nand ginst13237 (P2_R1203_U431, P2_R1203_U25, P2_U3432);
  nand ginst13238 (P2_R1203_U432, P2_R1203_U165, P2_U3080);
  not ginst13239 (P2_R1203_U433, P2_R1203_U139);
  nand ginst13240 (P2_R1203_U434, P2_R1203_U191, P2_R1203_U433);
  nand ginst13241 (P2_R1203_U435, P2_R1203_U139, P2_R1203_U166);
  nand ginst13242 (P2_R1203_U436, P2_R1203_U67, P2_U3485);
  nand ginst13243 (P2_R1203_U437, P2_R1203_U66, P2_U3083);
  not ginst13244 (P2_R1203_U438, P2_R1203_U140);
  nand ginst13245 (P2_R1203_U439, P2_R1203_U273, P2_R1203_U438);
  nand ginst13246 (P2_R1203_U44, P2_R1203_U176, P2_R1203_U192, P2_R1203_U351);
  nand ginst13247 (P2_R1203_U440, P2_R1203_U140, P2_R1203_U167);
  nand ginst13248 (P2_R1203_U441, P2_R1203_U65, P2_U3483);
  nand ginst13249 (P2_R1203_U442, P2_R1203_U168, P2_U3084);
  not ginst13250 (P2_R1203_U443, P2_R1203_U141);
  nand ginst13251 (P2_R1203_U444, P2_R1203_U269, P2_R1203_U443);
  nand ginst13252 (P2_R1203_U445, P2_R1203_U141, P2_R1203_U64);
  nand ginst13253 (P2_R1203_U446, P2_R1203_U63, P2_U3480);
  nand ginst13254 (P2_R1203_U447, P2_R1203_U62, P2_U3071);
  not ginst13255 (P2_R1203_U448, P2_R1203_U142);
  nand ginst13256 (P2_R1203_U449, P2_R1203_U265, P2_R1203_U448);
  not ginst13257 (P2_R1203_U45, P2_U3951);
  nand ginst13258 (P2_R1203_U450, P2_R1203_U142, P2_R1203_U169);
  nand ginst13259 (P2_R1203_U451, P2_R1203_U58, P2_U3477);
  nand ginst13260 (P2_R1203_U452, P2_R1203_U55, P2_U3075);
  nand ginst13261 (P2_R1203_U453, P2_R1203_U451, P2_R1203_U452);
  nand ginst13262 (P2_R1203_U454, P2_R1203_U59, P2_U3474);
  nand ginst13263 (P2_R1203_U455, P2_R1203_U56, P2_U3076);
  nand ginst13264 (P2_R1203_U456, P2_R1203_U338, P2_R1203_U90);
  nand ginst13265 (P2_R1203_U457, P2_R1203_U170, P2_R1203_U330);
  nand ginst13266 (P2_R1203_U458, P2_R1203_U60, P2_U3471);
  nand ginst13267 (P2_R1203_U459, P2_R1203_U57, P2_U3081);
  not ginst13268 (P2_R1203_U46, P2_U3459);
  nand ginst13269 (P2_R1203_U460, P2_R1203_U172, P2_R1203_U339);
  nand ginst13270 (P2_R1203_U461, P2_R1203_U171, P2_R1203_U255);
  nand ginst13271 (P2_R1203_U462, P2_R1203_U54, P2_U3468);
  nand ginst13272 (P2_R1203_U463, P2_R1203_U53, P2_U3082);
  not ginst13273 (P2_R1203_U464, P2_R1203_U145);
  nand ginst13274 (P2_R1203_U465, P2_R1203_U251, P2_R1203_U464);
  nand ginst13275 (P2_R1203_U466, P2_R1203_U145, P2_R1203_U173);
  nand ginst13276 (P2_R1203_U467, P2_R1203_U52, P2_U3465);
  nand ginst13277 (P2_R1203_U468, P2_R1203_U51, P2_U3074);
  not ginst13278 (P2_R1203_U469, P2_R1203_U146);
  not ginst13279 (P2_R1203_U47, P2_U3462);
  nand ginst13280 (P2_R1203_U470, P2_R1203_U247, P2_R1203_U469);
  nand ginst13281 (P2_R1203_U471, P2_R1203_U146, P2_R1203_U174);
  nand ginst13282 (P2_R1203_U472, P2_R1203_U48, P2_U3462);
  nand ginst13283 (P2_R1203_U473, P2_R1203_U47, P2_U3065);
  nand ginst13284 (P2_R1203_U474, P2_R1203_U472, P2_R1203_U473);
  nand ginst13285 (P2_R1203_U475, P2_R1203_U49, P2_U3459);
  nand ginst13286 (P2_R1203_U476, P2_R1203_U46, P2_U3064);
  nand ginst13287 (P2_R1203_U477, P2_R1203_U349, P2_R1203_U91);
  nand ginst13288 (P2_R1203_U478, P2_R1203_U175, P2_R1203_U341);
  not ginst13289 (P2_R1203_U48, P2_U3065);
  not ginst13290 (P2_R1203_U49, P2_U3064);
  nand ginst13291 (P2_R1203_U50, P2_R1203_U40, P2_U3085);
  not ginst13292 (P2_R1203_U51, P2_U3465);
  not ginst13293 (P2_R1203_U52, P2_U3074);
  not ginst13294 (P2_R1203_U53, P2_U3468);
  not ginst13295 (P2_R1203_U54, P2_U3082);
  not ginst13296 (P2_R1203_U55, P2_U3477);
  not ginst13297 (P2_R1203_U56, P2_U3474);
  not ginst13298 (P2_R1203_U57, P2_U3471);
  not ginst13299 (P2_R1203_U58, P2_U3075);
  not ginst13300 (P2_R1203_U59, P2_U3076);
  and ginst13301 (P2_R1203_U6, P2_R1203_U201, P2_R1203_U202);
  not ginst13302 (P2_R1203_U60, P2_U3081);
  nand ginst13303 (P2_R1203_U61, P2_R1203_U57, P2_U3081);
  not ginst13304 (P2_R1203_U62, P2_U3480);
  not ginst13305 (P2_R1203_U63, P2_U3071);
  nand ginst13306 (P2_R1203_U64, P2_R1203_U267, P2_R1203_U268);
  not ginst13307 (P2_R1203_U65, P2_U3084);
  not ginst13308 (P2_R1203_U66, P2_U3485);
  not ginst13309 (P2_R1203_U67, P2_U3083);
  not ginst13310 (P2_R1203_U68, P2_U3957);
  not ginst13311 (P2_R1203_U69, P2_U3078);
  and ginst13312 (P2_R1203_U7, P2_R1203_U240, P2_R1203_U241);
  not ginst13313 (P2_R1203_U70, P2_U3954);
  not ginst13314 (P2_R1203_U71, P2_U3955);
  not ginst13315 (P2_R1203_U72, P2_U3956);
  not ginst13316 (P2_R1203_U73, P2_U3068);
  not ginst13317 (P2_R1203_U74, P2_U3063);
  not ginst13318 (P2_R1203_U75, P2_U3077);
  nand ginst13319 (P2_R1203_U76, P2_R1203_U72, P2_U3077);
  not ginst13320 (P2_R1203_U77, P2_U3953);
  not ginst13321 (P2_R1203_U78, P2_U3067);
  not ginst13322 (P2_R1203_U79, P2_U3952);
  and ginst13323 (P2_R1203_U8, P2_R1203_U181, P2_R1203_U256);
  not ginst13324 (P2_R1203_U80, P2_U3060);
  not ginst13325 (P2_R1203_U81, P2_U3950);
  not ginst13326 (P2_R1203_U82, P2_U3059);
  nand ginst13327 (P2_R1203_U83, P2_R1203_U45, P2_U3059);
  not ginst13328 (P2_R1203_U84, P2_U3055);
  not ginst13329 (P2_R1203_U85, P2_U3949);
  not ginst13330 (P2_R1203_U86, P2_U3056);
  nand ginst13331 (P2_R1203_U87, P2_R1203_U128, P2_R1203_U301);
  nand ginst13332 (P2_R1203_U88, P2_R1203_U297, P2_R1203_U298);
  nand ginst13333 (P2_R1203_U89, P2_R1203_U318, P2_R1203_U76);
  and ginst13334 (P2_R1203_U9, P2_R1203_U257, P2_R1203_U258);
  nand ginst13335 (P2_R1203_U90, P2_R1203_U329, P2_R1203_U61);
  nand ginst13336 (P2_R1203_U91, P2_R1203_U340, P2_R1203_U50);
  not ginst13337 (P2_R1203_U92, P2_U3079);
  nand ginst13338 (P2_R1203_U93, P2_R1203_U394, P2_R1203_U395);
  nand ginst13339 (P2_R1203_U94, P2_R1203_U408, P2_R1203_U409);
  nand ginst13340 (P2_R1203_U95, P2_R1203_U413, P2_R1203_U414);
  nand ginst13341 (P2_R1203_U96, P2_R1203_U429, P2_R1203_U430);
  nand ginst13342 (P2_R1203_U97, P2_R1203_U434, P2_R1203_U435);
  nand ginst13343 (P2_R1203_U98, P2_R1203_U439, P2_R1203_U440);
  nand ginst13344 (P2_R1203_U99, P2_R1203_U444, P2_R1203_U445);
  and ginst13345 (P2_R1209_U10, P2_R1209_U215, P2_R1209_U218);
  not ginst13346 (P2_R1209_U100, P2_R1209_U40);
  not ginst13347 (P2_R1209_U101, P2_R1209_U41);
  nand ginst13348 (P2_R1209_U102, P2_R1209_U40, P2_R1209_U41);
  nand ginst13349 (P2_R1209_U103, P2_REG1_REG_2__SCAN_IN, P2_R1209_U96, P2_U3434);
  nand ginst13350 (P2_R1209_U104, P2_R1209_U102, P2_R1209_U5);
  nand ginst13351 (P2_R1209_U105, P2_REG1_REG_3__SCAN_IN, P2_U3437);
  nand ginst13352 (P2_R1209_U106, P2_R1209_U103, P2_R1209_U104, P2_R1209_U105);
  nand ginst13353 (P2_R1209_U107, P2_R1209_U32, P2_R1209_U33);
  nand ginst13354 (P2_R1209_U108, P2_R1209_U107, P2_U3443);
  nand ginst13355 (P2_R1209_U109, P2_R1209_U106, P2_R1209_U4);
  and ginst13356 (P2_R1209_U11, P2_R1209_U208, P2_R1209_U211);
  nand ginst13357 (P2_R1209_U110, P2_REG1_REG_5__SCAN_IN, P2_R1209_U89);
  not ginst13358 (P2_R1209_U111, P2_R1209_U39);
  or ginst13359 (P2_R1209_U112, P2_REG1_REG_7__SCAN_IN, P2_U3449);
  or ginst13360 (P2_R1209_U113, P2_REG1_REG_6__SCAN_IN, P2_U3446);
  not ginst13361 (P2_R1209_U114, P2_R1209_U20);
  nand ginst13362 (P2_R1209_U115, P2_R1209_U20, P2_R1209_U21);
  nand ginst13363 (P2_R1209_U116, P2_R1209_U115, P2_U3449);
  nand ginst13364 (P2_R1209_U117, P2_REG1_REG_7__SCAN_IN, P2_R1209_U114);
  nand ginst13365 (P2_R1209_U118, P2_R1209_U39, P2_R1209_U6);
  not ginst13366 (P2_R1209_U119, P2_R1209_U81);
  and ginst13367 (P2_R1209_U12, P2_R1209_U199, P2_R1209_U202);
  or ginst13368 (P2_R1209_U120, P2_REG1_REG_8__SCAN_IN, P2_U3452);
  nand ginst13369 (P2_R1209_U121, P2_R1209_U120, P2_R1209_U81);
  not ginst13370 (P2_R1209_U122, P2_R1209_U38);
  or ginst13371 (P2_R1209_U123, P2_REG1_REG_9__SCAN_IN, P2_U3455);
  or ginst13372 (P2_R1209_U124, P2_REG1_REG_6__SCAN_IN, P2_U3446);
  nand ginst13373 (P2_R1209_U125, P2_R1209_U124, P2_R1209_U39);
  nand ginst13374 (P2_R1209_U126, P2_R1209_U125, P2_R1209_U20, P2_R1209_U237, P2_R1209_U238);
  nand ginst13375 (P2_R1209_U127, P2_R1209_U111, P2_R1209_U20);
  nand ginst13376 (P2_R1209_U128, P2_REG1_REG_7__SCAN_IN, P2_U3449);
  nand ginst13377 (P2_R1209_U129, P2_R1209_U127, P2_R1209_U128, P2_R1209_U6);
  and ginst13378 (P2_R1209_U13, P2_R1209_U192, P2_R1209_U196);
  or ginst13379 (P2_R1209_U130, P2_REG1_REG_6__SCAN_IN, P2_U3446);
  nand ginst13380 (P2_R1209_U131, P2_R1209_U101, P2_R1209_U97);
  nand ginst13381 (P2_R1209_U132, P2_REG1_REG_2__SCAN_IN, P2_U3434);
  not ginst13382 (P2_R1209_U133, P2_R1209_U43);
  nand ginst13383 (P2_R1209_U134, P2_R1209_U100, P2_R1209_U5);
  nand ginst13384 (P2_R1209_U135, P2_R1209_U43, P2_R1209_U96);
  nand ginst13385 (P2_R1209_U136, P2_REG1_REG_3__SCAN_IN, P2_U3437);
  not ginst13386 (P2_R1209_U137, P2_R1209_U42);
  or ginst13387 (P2_R1209_U138, P2_REG1_REG_4__SCAN_IN, P2_U3440);
  nand ginst13388 (P2_R1209_U139, P2_R1209_U138, P2_R1209_U42);
  and ginst13389 (P2_R1209_U14, P2_R1209_U148, P2_R1209_U151);
  nand ginst13390 (P2_R1209_U140, P2_R1209_U139, P2_R1209_U244, P2_R1209_U245, P2_R1209_U32);
  nand ginst13391 (P2_R1209_U141, P2_R1209_U137, P2_R1209_U32);
  nand ginst13392 (P2_R1209_U142, P2_REG1_REG_5__SCAN_IN, P2_U3443);
  nand ginst13393 (P2_R1209_U143, P2_R1209_U141, P2_R1209_U142, P2_R1209_U4);
  or ginst13394 (P2_R1209_U144, P2_REG1_REG_4__SCAN_IN, P2_U3440);
  nand ginst13395 (P2_R1209_U145, P2_R1209_U100, P2_R1209_U97);
  not ginst13396 (P2_R1209_U146, P2_R1209_U82);
  nand ginst13397 (P2_R1209_U147, P2_REG1_REG_3__SCAN_IN, P2_U3437);
  nand ginst13398 (P2_R1209_U148, P2_R1209_U256, P2_R1209_U257, P2_R1209_U40, P2_R1209_U41);
  nand ginst13399 (P2_R1209_U149, P2_R1209_U40, P2_R1209_U41);
  and ginst13400 (P2_R1209_U15, P2_R1209_U140, P2_R1209_U143);
  nand ginst13401 (P2_R1209_U150, P2_REG1_REG_2__SCAN_IN, P2_U3434);
  nand ginst13402 (P2_R1209_U151, P2_R1209_U149, P2_R1209_U150, P2_R1209_U97);
  or ginst13403 (P2_R1209_U152, P2_REG1_REG_1__SCAN_IN, P2_U3431);
  not ginst13404 (P2_R1209_U153, P2_R1209_U83);
  or ginst13405 (P2_R1209_U154, P2_REG1_REG_9__SCAN_IN, P2_U3455);
  or ginst13406 (P2_R1209_U155, P2_REG1_REG_10__SCAN_IN, P2_U3458);
  nand ginst13407 (P2_R1209_U156, P2_R1209_U7, P2_R1209_U93);
  nand ginst13408 (P2_R1209_U157, P2_REG1_REG_10__SCAN_IN, P2_U3458);
  nand ginst13409 (P2_R1209_U158, P2_R1209_U156, P2_R1209_U157, P2_R1209_U90);
  or ginst13410 (P2_R1209_U159, P2_REG1_REG_10__SCAN_IN, P2_U3458);
  and ginst13411 (P2_R1209_U16, P2_R1209_U126, P2_R1209_U129);
  nand ginst13412 (P2_R1209_U160, P2_R1209_U120, P2_R1209_U7, P2_R1209_U81);
  nand ginst13413 (P2_R1209_U161, P2_R1209_U158, P2_R1209_U159);
  not ginst13414 (P2_R1209_U162, P2_R1209_U88);
  or ginst13415 (P2_R1209_U163, P2_REG1_REG_13__SCAN_IN, P2_U3467);
  or ginst13416 (P2_R1209_U164, P2_REG1_REG_12__SCAN_IN, P2_U3464);
  nand ginst13417 (P2_R1209_U165, P2_R1209_U8, P2_R1209_U92);
  nand ginst13418 (P2_R1209_U166, P2_REG1_REG_13__SCAN_IN, P2_U3467);
  nand ginst13419 (P2_R1209_U167, P2_R1209_U165, P2_R1209_U166, P2_R1209_U91);
  or ginst13420 (P2_R1209_U168, P2_REG1_REG_11__SCAN_IN, P2_U3461);
  or ginst13421 (P2_R1209_U169, P2_REG1_REG_13__SCAN_IN, P2_U3467);
  not ginst13422 (P2_R1209_U17, P2_REG1_REG_6__SCAN_IN);
  nand ginst13423 (P2_R1209_U170, P2_R1209_U168, P2_R1209_U8, P2_R1209_U88);
  nand ginst13424 (P2_R1209_U171, P2_R1209_U167, P2_R1209_U169);
  not ginst13425 (P2_R1209_U172, P2_R1209_U87);
  or ginst13426 (P2_R1209_U173, P2_REG1_REG_14__SCAN_IN, P2_U3470);
  nand ginst13427 (P2_R1209_U174, P2_R1209_U173, P2_R1209_U87);
  nand ginst13428 (P2_R1209_U175, P2_REG1_REG_14__SCAN_IN, P2_U3470);
  not ginst13429 (P2_R1209_U176, P2_R1209_U86);
  or ginst13430 (P2_R1209_U177, P2_REG1_REG_15__SCAN_IN, P2_U3473);
  nand ginst13431 (P2_R1209_U178, P2_R1209_U177, P2_R1209_U86);
  nand ginst13432 (P2_R1209_U179, P2_REG1_REG_15__SCAN_IN, P2_U3473);
  not ginst13433 (P2_R1209_U18, P2_U3446);
  not ginst13434 (P2_R1209_U180, P2_R1209_U66);
  or ginst13435 (P2_R1209_U181, P2_REG1_REG_17__SCAN_IN, P2_U3479);
  or ginst13436 (P2_R1209_U182, P2_REG1_REG_16__SCAN_IN, P2_U3476);
  not ginst13437 (P2_R1209_U183, P2_R1209_U47);
  nand ginst13438 (P2_R1209_U184, P2_R1209_U47, P2_R1209_U48);
  nand ginst13439 (P2_R1209_U185, P2_R1209_U184, P2_U3479);
  nand ginst13440 (P2_R1209_U186, P2_REG1_REG_17__SCAN_IN, P2_R1209_U183);
  nand ginst13441 (P2_R1209_U187, P2_R1209_U66, P2_R1209_U9);
  not ginst13442 (P2_R1209_U188, P2_R1209_U65);
  or ginst13443 (P2_R1209_U189, P2_REG1_REG_18__SCAN_IN, P2_U3482);
  not ginst13444 (P2_R1209_U19, P2_U3449);
  nand ginst13445 (P2_R1209_U190, P2_R1209_U189, P2_R1209_U65);
  nand ginst13446 (P2_R1209_U191, P2_REG1_REG_18__SCAN_IN, P2_U3482);
  nand ginst13447 (P2_R1209_U192, P2_R1209_U190, P2_R1209_U191, P2_R1209_U260, P2_R1209_U261);
  nand ginst13448 (P2_R1209_U193, P2_REG1_REG_18__SCAN_IN, P2_U3482);
  nand ginst13449 (P2_R1209_U194, P2_R1209_U188, P2_R1209_U193);
  or ginst13450 (P2_R1209_U195, P2_REG1_REG_18__SCAN_IN, P2_U3482);
  nand ginst13451 (P2_R1209_U196, P2_R1209_U194, P2_R1209_U195, P2_R1209_U264);
  or ginst13452 (P2_R1209_U197, P2_REG1_REG_16__SCAN_IN, P2_U3476);
  nand ginst13453 (P2_R1209_U198, P2_R1209_U197, P2_R1209_U66);
  nand ginst13454 (P2_R1209_U199, P2_R1209_U198, P2_R1209_U272, P2_R1209_U273, P2_R1209_U47);
  nand ginst13455 (P2_R1209_U20, P2_REG1_REG_6__SCAN_IN, P2_U3446);
  nand ginst13456 (P2_R1209_U200, P2_R1209_U180, P2_R1209_U47);
  nand ginst13457 (P2_R1209_U201, P2_REG1_REG_17__SCAN_IN, P2_U3479);
  nand ginst13458 (P2_R1209_U202, P2_R1209_U200, P2_R1209_U201, P2_R1209_U9);
  or ginst13459 (P2_R1209_U203, P2_REG1_REG_16__SCAN_IN, P2_U3476);
  nand ginst13460 (P2_R1209_U204, P2_R1209_U168, P2_R1209_U88);
  not ginst13461 (P2_R1209_U205, P2_R1209_U67);
  or ginst13462 (P2_R1209_U206, P2_REG1_REG_12__SCAN_IN, P2_U3464);
  nand ginst13463 (P2_R1209_U207, P2_R1209_U206, P2_R1209_U67);
  nand ginst13464 (P2_R1209_U208, P2_R1209_U207, P2_R1209_U293, P2_R1209_U294, P2_R1209_U91);
  nand ginst13465 (P2_R1209_U209, P2_R1209_U205, P2_R1209_U91);
  not ginst13466 (P2_R1209_U21, P2_REG1_REG_7__SCAN_IN);
  nand ginst13467 (P2_R1209_U210, P2_REG1_REG_13__SCAN_IN, P2_U3467);
  nand ginst13468 (P2_R1209_U211, P2_R1209_U209, P2_R1209_U210, P2_R1209_U8);
  or ginst13469 (P2_R1209_U212, P2_REG1_REG_12__SCAN_IN, P2_U3464);
  or ginst13470 (P2_R1209_U213, P2_REG1_REG_9__SCAN_IN, P2_U3455);
  nand ginst13471 (P2_R1209_U214, P2_R1209_U213, P2_R1209_U38);
  nand ginst13472 (P2_R1209_U215, P2_R1209_U214, P2_R1209_U305, P2_R1209_U306, P2_R1209_U90);
  nand ginst13473 (P2_R1209_U216, P2_R1209_U122, P2_R1209_U90);
  nand ginst13474 (P2_R1209_U217, P2_REG1_REG_10__SCAN_IN, P2_U3458);
  nand ginst13475 (P2_R1209_U218, P2_R1209_U216, P2_R1209_U217, P2_R1209_U7);
  nand ginst13476 (P2_R1209_U219, P2_R1209_U123, P2_R1209_U90);
  not ginst13477 (P2_R1209_U22, P2_REG1_REG_4__SCAN_IN);
  nand ginst13478 (P2_R1209_U220, P2_R1209_U120, P2_R1209_U49);
  nand ginst13479 (P2_R1209_U221, P2_R1209_U130, P2_R1209_U20);
  nand ginst13480 (P2_R1209_U222, P2_R1209_U144, P2_R1209_U32);
  nand ginst13481 (P2_R1209_U223, P2_R1209_U147, P2_R1209_U96);
  nand ginst13482 (P2_R1209_U224, P2_R1209_U203, P2_R1209_U47);
  nand ginst13483 (P2_R1209_U225, P2_R1209_U212, P2_R1209_U91);
  nand ginst13484 (P2_R1209_U226, P2_R1209_U168, P2_R1209_U56);
  nand ginst13485 (P2_R1209_U227, P2_R1209_U37, P2_U3455);
  nand ginst13486 (P2_R1209_U228, P2_REG1_REG_9__SCAN_IN, P2_R1209_U36);
  nand ginst13487 (P2_R1209_U229, P2_R1209_U227, P2_R1209_U228);
  not ginst13488 (P2_R1209_U23, P2_U3440);
  nand ginst13489 (P2_R1209_U230, P2_R1209_U219, P2_R1209_U38);
  nand ginst13490 (P2_R1209_U231, P2_R1209_U122, P2_R1209_U229);
  nand ginst13491 (P2_R1209_U232, P2_R1209_U34, P2_U3452);
  nand ginst13492 (P2_R1209_U233, P2_REG1_REG_8__SCAN_IN, P2_R1209_U35);
  nand ginst13493 (P2_R1209_U234, P2_R1209_U232, P2_R1209_U233);
  nand ginst13494 (P2_R1209_U235, P2_R1209_U220, P2_R1209_U81);
  nand ginst13495 (P2_R1209_U236, P2_R1209_U119, P2_R1209_U234);
  nand ginst13496 (P2_R1209_U237, P2_R1209_U21, P2_U3449);
  nand ginst13497 (P2_R1209_U238, P2_REG1_REG_7__SCAN_IN, P2_R1209_U19);
  nand ginst13498 (P2_R1209_U239, P2_R1209_U17, P2_U3446);
  not ginst13499 (P2_R1209_U24, P2_U3443);
  nand ginst13500 (P2_R1209_U240, P2_REG1_REG_6__SCAN_IN, P2_R1209_U18);
  nand ginst13501 (P2_R1209_U241, P2_R1209_U239, P2_R1209_U240);
  nand ginst13502 (P2_R1209_U242, P2_R1209_U221, P2_R1209_U39);
  nand ginst13503 (P2_R1209_U243, P2_R1209_U111, P2_R1209_U241);
  nand ginst13504 (P2_R1209_U244, P2_R1209_U33, P2_U3443);
  nand ginst13505 (P2_R1209_U245, P2_REG1_REG_5__SCAN_IN, P2_R1209_U24);
  nand ginst13506 (P2_R1209_U246, P2_R1209_U22, P2_U3440);
  nand ginst13507 (P2_R1209_U247, P2_REG1_REG_4__SCAN_IN, P2_R1209_U23);
  nand ginst13508 (P2_R1209_U248, P2_R1209_U246, P2_R1209_U247);
  nand ginst13509 (P2_R1209_U249, P2_R1209_U222, P2_R1209_U42);
  not ginst13510 (P2_R1209_U25, P2_REG1_REG_2__SCAN_IN);
  nand ginst13511 (P2_R1209_U250, P2_R1209_U137, P2_R1209_U248);
  nand ginst13512 (P2_R1209_U251, P2_R1209_U30, P2_U3437);
  nand ginst13513 (P2_R1209_U252, P2_REG1_REG_3__SCAN_IN, P2_R1209_U31);
  nand ginst13514 (P2_R1209_U253, P2_R1209_U251, P2_R1209_U252);
  nand ginst13515 (P2_R1209_U254, P2_R1209_U223, P2_R1209_U82);
  nand ginst13516 (P2_R1209_U255, P2_R1209_U146, P2_R1209_U253);
  nand ginst13517 (P2_R1209_U256, P2_R1209_U25, P2_U3434);
  nand ginst13518 (P2_R1209_U257, P2_REG1_REG_2__SCAN_IN, P2_R1209_U26);
  nand ginst13519 (P2_R1209_U258, P2_R1209_U83, P2_R1209_U98);
  nand ginst13520 (P2_R1209_U259, P2_R1209_U153, P2_R1209_U29);
  not ginst13521 (P2_R1209_U26, P2_U3434);
  nand ginst13522 (P2_R1209_U260, P2_R1209_U85, P2_U3424);
  nand ginst13523 (P2_R1209_U261, P2_REG1_REG_19__SCAN_IN, P2_R1209_U84);
  nand ginst13524 (P2_R1209_U262, P2_R1209_U85, P2_U3424);
  nand ginst13525 (P2_R1209_U263, P2_REG1_REG_19__SCAN_IN, P2_R1209_U84);
  nand ginst13526 (P2_R1209_U264, P2_R1209_U262, P2_R1209_U263);
  nand ginst13527 (P2_R1209_U265, P2_R1209_U63, P2_U3482);
  nand ginst13528 (P2_R1209_U266, P2_REG1_REG_18__SCAN_IN, P2_R1209_U64);
  nand ginst13529 (P2_R1209_U267, P2_R1209_U63, P2_U3482);
  nand ginst13530 (P2_R1209_U268, P2_REG1_REG_18__SCAN_IN, P2_R1209_U64);
  nand ginst13531 (P2_R1209_U269, P2_R1209_U267, P2_R1209_U268);
  not ginst13532 (P2_R1209_U27, P2_REG1_REG_0__SCAN_IN);
  nand ginst13533 (P2_R1209_U270, P2_R1209_U265, P2_R1209_U266, P2_R1209_U65);
  nand ginst13534 (P2_R1209_U271, P2_R1209_U188, P2_R1209_U269);
  nand ginst13535 (P2_R1209_U272, P2_R1209_U48, P2_U3479);
  nand ginst13536 (P2_R1209_U273, P2_REG1_REG_17__SCAN_IN, P2_R1209_U46);
  nand ginst13537 (P2_R1209_U274, P2_R1209_U44, P2_U3476);
  nand ginst13538 (P2_R1209_U275, P2_REG1_REG_16__SCAN_IN, P2_R1209_U45);
  nand ginst13539 (P2_R1209_U276, P2_R1209_U274, P2_R1209_U275);
  nand ginst13540 (P2_R1209_U277, P2_R1209_U224, P2_R1209_U66);
  nand ginst13541 (P2_R1209_U278, P2_R1209_U180, P2_R1209_U276);
  nand ginst13542 (P2_R1209_U279, P2_R1209_U61, P2_U3473);
  not ginst13543 (P2_R1209_U28, P2_U3425);
  nand ginst13544 (P2_R1209_U280, P2_REG1_REG_15__SCAN_IN, P2_R1209_U62);
  nand ginst13545 (P2_R1209_U281, P2_R1209_U61, P2_U3473);
  nand ginst13546 (P2_R1209_U282, P2_REG1_REG_15__SCAN_IN, P2_R1209_U62);
  nand ginst13547 (P2_R1209_U283, P2_R1209_U281, P2_R1209_U282);
  nand ginst13548 (P2_R1209_U284, P2_R1209_U279, P2_R1209_U280, P2_R1209_U86);
  nand ginst13549 (P2_R1209_U285, P2_R1209_U176, P2_R1209_U283);
  nand ginst13550 (P2_R1209_U286, P2_R1209_U59, P2_U3470);
  nand ginst13551 (P2_R1209_U287, P2_REG1_REG_14__SCAN_IN, P2_R1209_U60);
  nand ginst13552 (P2_R1209_U288, P2_R1209_U59, P2_U3470);
  nand ginst13553 (P2_R1209_U289, P2_REG1_REG_14__SCAN_IN, P2_R1209_U60);
  nand ginst13554 (P2_R1209_U29, P2_REG1_REG_0__SCAN_IN, P2_U3425);
  nand ginst13555 (P2_R1209_U290, P2_R1209_U288, P2_R1209_U289);
  nand ginst13556 (P2_R1209_U291, P2_R1209_U286, P2_R1209_U287, P2_R1209_U87);
  nand ginst13557 (P2_R1209_U292, P2_R1209_U172, P2_R1209_U290);
  nand ginst13558 (P2_R1209_U293, P2_R1209_U57, P2_U3467);
  nand ginst13559 (P2_R1209_U294, P2_REG1_REG_13__SCAN_IN, P2_R1209_U58);
  nand ginst13560 (P2_R1209_U295, P2_R1209_U52, P2_U3464);
  nand ginst13561 (P2_R1209_U296, P2_REG1_REG_12__SCAN_IN, P2_R1209_U53);
  nand ginst13562 (P2_R1209_U297, P2_R1209_U295, P2_R1209_U296);
  nand ginst13563 (P2_R1209_U298, P2_R1209_U225, P2_R1209_U67);
  nand ginst13564 (P2_R1209_U299, P2_R1209_U205, P2_R1209_U297);
  not ginst13565 (P2_R1209_U30, P2_REG1_REG_3__SCAN_IN);
  nand ginst13566 (P2_R1209_U300, P2_R1209_U54, P2_U3461);
  nand ginst13567 (P2_R1209_U301, P2_REG1_REG_11__SCAN_IN, P2_R1209_U55);
  nand ginst13568 (P2_R1209_U302, P2_R1209_U300, P2_R1209_U301);
  nand ginst13569 (P2_R1209_U303, P2_R1209_U226, P2_R1209_U88);
  nand ginst13570 (P2_R1209_U304, P2_R1209_U162, P2_R1209_U302);
  nand ginst13571 (P2_R1209_U305, P2_R1209_U50, P2_U3458);
  nand ginst13572 (P2_R1209_U306, P2_REG1_REG_10__SCAN_IN, P2_R1209_U51);
  nand ginst13573 (P2_R1209_U307, P2_R1209_U27, P2_U3425);
  nand ginst13574 (P2_R1209_U308, P2_REG1_REG_0__SCAN_IN, P2_R1209_U28);
  not ginst13575 (P2_R1209_U31, P2_U3437);
  nand ginst13576 (P2_R1209_U32, P2_REG1_REG_4__SCAN_IN, P2_U3440);
  not ginst13577 (P2_R1209_U33, P2_REG1_REG_5__SCAN_IN);
  not ginst13578 (P2_R1209_U34, P2_REG1_REG_8__SCAN_IN);
  not ginst13579 (P2_R1209_U35, P2_U3452);
  not ginst13580 (P2_R1209_U36, P2_U3455);
  not ginst13581 (P2_R1209_U37, P2_REG1_REG_9__SCAN_IN);
  nand ginst13582 (P2_R1209_U38, P2_R1209_U121, P2_R1209_U49);
  nand ginst13583 (P2_R1209_U39, P2_R1209_U108, P2_R1209_U109, P2_R1209_U110);
  and ginst13584 (P2_R1209_U4, P2_R1209_U94, P2_R1209_U95);
  nand ginst13585 (P2_R1209_U40, P2_R1209_U98, P2_R1209_U99);
  nand ginst13586 (P2_R1209_U41, P2_REG1_REG_1__SCAN_IN, P2_U3431);
  nand ginst13587 (P2_R1209_U42, P2_R1209_U134, P2_R1209_U135, P2_R1209_U136);
  nand ginst13588 (P2_R1209_U43, P2_R1209_U131, P2_R1209_U132);
  not ginst13589 (P2_R1209_U44, P2_REG1_REG_16__SCAN_IN);
  not ginst13590 (P2_R1209_U45, P2_U3476);
  not ginst13591 (P2_R1209_U46, P2_U3479);
  nand ginst13592 (P2_R1209_U47, P2_REG1_REG_16__SCAN_IN, P2_U3476);
  not ginst13593 (P2_R1209_U48, P2_REG1_REG_17__SCAN_IN);
  nand ginst13594 (P2_R1209_U49, P2_REG1_REG_8__SCAN_IN, P2_U3452);
  and ginst13595 (P2_R1209_U5, P2_R1209_U96, P2_R1209_U97);
  not ginst13596 (P2_R1209_U50, P2_REG1_REG_10__SCAN_IN);
  not ginst13597 (P2_R1209_U51, P2_U3458);
  not ginst13598 (P2_R1209_U52, P2_REG1_REG_12__SCAN_IN);
  not ginst13599 (P2_R1209_U53, P2_U3464);
  not ginst13600 (P2_R1209_U54, P2_REG1_REG_11__SCAN_IN);
  not ginst13601 (P2_R1209_U55, P2_U3461);
  nand ginst13602 (P2_R1209_U56, P2_REG1_REG_11__SCAN_IN, P2_U3461);
  not ginst13603 (P2_R1209_U57, P2_REG1_REG_13__SCAN_IN);
  not ginst13604 (P2_R1209_U58, P2_U3467);
  not ginst13605 (P2_R1209_U59, P2_REG1_REG_14__SCAN_IN);
  and ginst13606 (P2_R1209_U6, P2_R1209_U112, P2_R1209_U113);
  not ginst13607 (P2_R1209_U60, P2_U3470);
  not ginst13608 (P2_R1209_U61, P2_REG1_REG_15__SCAN_IN);
  not ginst13609 (P2_R1209_U62, P2_U3473);
  not ginst13610 (P2_R1209_U63, P2_REG1_REG_18__SCAN_IN);
  not ginst13611 (P2_R1209_U64, P2_U3482);
  nand ginst13612 (P2_R1209_U65, P2_R1209_U185, P2_R1209_U186, P2_R1209_U187);
  nand ginst13613 (P2_R1209_U66, P2_R1209_U178, P2_R1209_U179);
  nand ginst13614 (P2_R1209_U67, P2_R1209_U204, P2_R1209_U56);
  nand ginst13615 (P2_R1209_U68, P2_R1209_U258, P2_R1209_U259);
  nand ginst13616 (P2_R1209_U69, P2_R1209_U307, P2_R1209_U308);
  and ginst13617 (P2_R1209_U7, P2_R1209_U154, P2_R1209_U155);
  nand ginst13618 (P2_R1209_U70, P2_R1209_U230, P2_R1209_U231);
  nand ginst13619 (P2_R1209_U71, P2_R1209_U235, P2_R1209_U236);
  nand ginst13620 (P2_R1209_U72, P2_R1209_U242, P2_R1209_U243);
  nand ginst13621 (P2_R1209_U73, P2_R1209_U249, P2_R1209_U250);
  nand ginst13622 (P2_R1209_U74, P2_R1209_U254, P2_R1209_U255);
  nand ginst13623 (P2_R1209_U75, P2_R1209_U270, P2_R1209_U271);
  nand ginst13624 (P2_R1209_U76, P2_R1209_U277, P2_R1209_U278);
  nand ginst13625 (P2_R1209_U77, P2_R1209_U284, P2_R1209_U285);
  nand ginst13626 (P2_R1209_U78, P2_R1209_U291, P2_R1209_U292);
  nand ginst13627 (P2_R1209_U79, P2_R1209_U298, P2_R1209_U299);
  and ginst13628 (P2_R1209_U8, P2_R1209_U163, P2_R1209_U164);
  nand ginst13629 (P2_R1209_U80, P2_R1209_U303, P2_R1209_U304);
  nand ginst13630 (P2_R1209_U81, P2_R1209_U116, P2_R1209_U117, P2_R1209_U118);
  nand ginst13631 (P2_R1209_U82, P2_R1209_U133, P2_R1209_U145);
  nand ginst13632 (P2_R1209_U83, P2_R1209_U152, P2_R1209_U41);
  not ginst13633 (P2_R1209_U84, P2_U3424);
  not ginst13634 (P2_R1209_U85, P2_REG1_REG_19__SCAN_IN);
  nand ginst13635 (P2_R1209_U86, P2_R1209_U174, P2_R1209_U175);
  nand ginst13636 (P2_R1209_U87, P2_R1209_U170, P2_R1209_U171);
  nand ginst13637 (P2_R1209_U88, P2_R1209_U160, P2_R1209_U161);
  not ginst13638 (P2_R1209_U89, P2_R1209_U32);
  and ginst13639 (P2_R1209_U9, P2_R1209_U181, P2_R1209_U182);
  nand ginst13640 (P2_R1209_U90, P2_REG1_REG_9__SCAN_IN, P2_U3455);
  nand ginst13641 (P2_R1209_U91, P2_REG1_REG_12__SCAN_IN, P2_U3464);
  not ginst13642 (P2_R1209_U92, P2_R1209_U56);
  not ginst13643 (P2_R1209_U93, P2_R1209_U49);
  or ginst13644 (P2_R1209_U94, P2_REG1_REG_5__SCAN_IN, P2_U3443);
  or ginst13645 (P2_R1209_U95, P2_REG1_REG_4__SCAN_IN, P2_U3440);
  or ginst13646 (P2_R1209_U96, P2_REG1_REG_3__SCAN_IN, P2_U3437);
  or ginst13647 (P2_R1209_U97, P2_REG1_REG_2__SCAN_IN, P2_U3434);
  not ginst13648 (P2_R1209_U98, P2_R1209_U29);
  or ginst13649 (P2_R1209_U99, P2_REG1_REG_1__SCAN_IN, P2_U3431);
  and ginst13650 (P2_R1215_U10, P2_R1215_U271, P2_R1215_U272);
  nand ginst13651 (P2_R1215_U100, P2_R1215_U393, P2_R1215_U394);
  nand ginst13652 (P2_R1215_U101, P2_R1215_U398, P2_R1215_U399);
  nand ginst13653 (P2_R1215_U102, P2_R1215_U407, P2_R1215_U408);
  nand ginst13654 (P2_R1215_U103, P2_R1215_U414, P2_R1215_U415);
  nand ginst13655 (P2_R1215_U104, P2_R1215_U421, P2_R1215_U422);
  nand ginst13656 (P2_R1215_U105, P2_R1215_U428, P2_R1215_U429);
  nand ginst13657 (P2_R1215_U106, P2_R1215_U433, P2_R1215_U434);
  nand ginst13658 (P2_R1215_U107, P2_R1215_U440, P2_R1215_U441);
  nand ginst13659 (P2_R1215_U108, P2_R1215_U447, P2_R1215_U448);
  nand ginst13660 (P2_R1215_U109, P2_R1215_U461, P2_R1215_U462);
  and ginst13661 (P2_R1215_U11, P2_R1215_U348, P2_R1215_U351);
  nand ginst13662 (P2_R1215_U110, P2_R1215_U466, P2_R1215_U467);
  nand ginst13663 (P2_R1215_U111, P2_R1215_U473, P2_R1215_U474);
  nand ginst13664 (P2_R1215_U112, P2_R1215_U480, P2_R1215_U481);
  nand ginst13665 (P2_R1215_U113, P2_R1215_U487, P2_R1215_U488);
  nand ginst13666 (P2_R1215_U114, P2_R1215_U494, P2_R1215_U495);
  nand ginst13667 (P2_R1215_U115, P2_R1215_U499, P2_R1215_U500);
  and ginst13668 (P2_R1215_U116, P2_U3070, P2_U3435);
  and ginst13669 (P2_R1215_U117, P2_R1215_U187, P2_R1215_U189);
  and ginst13670 (P2_R1215_U118, P2_R1215_U192, P2_R1215_U194);
  and ginst13671 (P2_R1215_U119, P2_R1215_U200, P2_R1215_U201);
  and ginst13672 (P2_R1215_U12, P2_R1215_U341, P2_R1215_U344);
  and ginst13673 (P2_R1215_U120, P2_R1215_U23, P2_R1215_U381, P2_R1215_U382);
  and ginst13674 (P2_R1215_U121, P2_R1215_U212, P2_R1215_U6);
  and ginst13675 (P2_R1215_U122, P2_R1215_U218, P2_R1215_U220);
  and ginst13676 (P2_R1215_U123, P2_R1215_U35, P2_R1215_U388, P2_R1215_U389);
  and ginst13677 (P2_R1215_U124, P2_R1215_U226, P2_R1215_U4);
  and ginst13678 (P2_R1215_U125, P2_R1215_U181, P2_R1215_U234);
  and ginst13679 (P2_R1215_U126, P2_R1215_U204, P2_R1215_U7);
  and ginst13680 (P2_R1215_U127, P2_R1215_U171, P2_R1215_U239);
  and ginst13681 (P2_R1215_U128, P2_R1215_U250, P2_R1215_U8);
  and ginst13682 (P2_R1215_U129, P2_R1215_U172, P2_R1215_U248);
  and ginst13683 (P2_R1215_U13, P2_R1215_U332, P2_R1215_U335);
  and ginst13684 (P2_R1215_U130, P2_R1215_U267, P2_R1215_U268);
  and ginst13685 (P2_R1215_U131, P2_R1215_U10, P2_R1215_U282);
  and ginst13686 (P2_R1215_U132, P2_R1215_U280, P2_R1215_U285);
  and ginst13687 (P2_R1215_U133, P2_R1215_U298, P2_R1215_U301);
  and ginst13688 (P2_R1215_U134, P2_R1215_U302, P2_R1215_U368);
  and ginst13689 (P2_R1215_U135, P2_R1215_U160, P2_R1215_U278);
  and ginst13690 (P2_R1215_U136, P2_R1215_U454, P2_R1215_U455, P2_R1215_U81);
  and ginst13691 (P2_R1215_U137, P2_R1215_U10, P2_R1215_U325);
  and ginst13692 (P2_R1215_U138, P2_R1215_U468, P2_R1215_U469, P2_R1215_U60);
  and ginst13693 (P2_R1215_U139, P2_R1215_U334, P2_R1215_U9);
  and ginst13694 (P2_R1215_U14, P2_R1215_U323, P2_R1215_U326);
  and ginst13695 (P2_R1215_U140, P2_R1215_U172, P2_R1215_U489, P2_R1215_U490);
  and ginst13696 (P2_R1215_U141, P2_R1215_U343, P2_R1215_U8);
  and ginst13697 (P2_R1215_U142, P2_R1215_U171, P2_R1215_U501, P2_R1215_U502);
  and ginst13698 (P2_R1215_U143, P2_R1215_U350, P2_R1215_U7);
  nand ginst13699 (P2_R1215_U144, P2_R1215_U119, P2_R1215_U202);
  nand ginst13700 (P2_R1215_U145, P2_R1215_U217, P2_R1215_U229);
  not ginst13701 (P2_R1215_U146, P2_U3057);
  not ginst13702 (P2_R1215_U147, P2_U3960);
  and ginst13703 (P2_R1215_U148, P2_R1215_U402, P2_R1215_U403);
  nand ginst13704 (P2_R1215_U149, P2_R1215_U169, P2_R1215_U304, P2_R1215_U364);
  and ginst13705 (P2_R1215_U15, P2_R1215_U318, P2_R1215_U320);
  and ginst13706 (P2_R1215_U150, P2_R1215_U409, P2_R1215_U410);
  nand ginst13707 (P2_R1215_U151, P2_R1215_U134, P2_R1215_U369, P2_R1215_U370);
  and ginst13708 (P2_R1215_U152, P2_R1215_U416, P2_R1215_U417);
  nand ginst13709 (P2_R1215_U153, P2_R1215_U299, P2_R1215_U365, P2_R1215_U87);
  and ginst13710 (P2_R1215_U154, P2_R1215_U423, P2_R1215_U424);
  nand ginst13711 (P2_R1215_U155, P2_R1215_U292, P2_R1215_U293);
  and ginst13712 (P2_R1215_U156, P2_R1215_U435, P2_R1215_U436);
  nand ginst13713 (P2_R1215_U157, P2_R1215_U288, P2_R1215_U289);
  and ginst13714 (P2_R1215_U158, P2_R1215_U442, P2_R1215_U443);
  nand ginst13715 (P2_R1215_U159, P2_R1215_U132, P2_R1215_U284);
  and ginst13716 (P2_R1215_U16, P2_R1215_U310, P2_R1215_U313);
  and ginst13717 (P2_R1215_U160, P2_R1215_U449, P2_R1215_U450);
  nand ginst13718 (P2_R1215_U161, P2_R1215_U327, P2_R1215_U44);
  nand ginst13719 (P2_R1215_U162, P2_R1215_U130, P2_R1215_U269);
  and ginst13720 (P2_R1215_U163, P2_R1215_U475, P2_R1215_U476);
  nand ginst13721 (P2_R1215_U164, P2_R1215_U256, P2_R1215_U257);
  and ginst13722 (P2_R1215_U165, P2_R1215_U482, P2_R1215_U483);
  nand ginst13723 (P2_R1215_U166, P2_R1215_U252, P2_R1215_U253);
  nand ginst13724 (P2_R1215_U167, P2_R1215_U242, P2_R1215_U243);
  nand ginst13725 (P2_R1215_U168, P2_R1215_U366, P2_R1215_U367);
  nand ginst13726 (P2_R1215_U169, P2_R1215_U151, P2_U3056);
  and ginst13727 (P2_R1215_U17, P2_R1215_U232, P2_R1215_U235);
  not ginst13728 (P2_R1215_U170, P2_R1215_U35);
  nand ginst13729 (P2_R1215_U171, P2_U3085, P2_U3456);
  nand ginst13730 (P2_R1215_U172, P2_U3074, P2_U3465);
  nand ginst13731 (P2_R1215_U173, P2_U3060, P2_U3952);
  not ginst13732 (P2_R1215_U174, P2_R1215_U69);
  not ginst13733 (P2_R1215_U175, P2_R1215_U78);
  nand ginst13734 (P2_R1215_U176, P2_U3067, P2_U3953);
  not ginst13735 (P2_R1215_U177, P2_R1215_U62);
  or ginst13736 (P2_R1215_U178, P2_U3069, P2_U3444);
  or ginst13737 (P2_R1215_U179, P2_U3062, P2_U3441);
  and ginst13738 (P2_R1215_U18, P2_R1215_U224, P2_R1215_U227);
  or ginst13739 (P2_R1215_U180, P2_U3066, P2_U3438);
  or ginst13740 (P2_R1215_U181, P2_U3070, P2_U3435);
  not ginst13741 (P2_R1215_U182, P2_R1215_U32);
  or ginst13742 (P2_R1215_U183, P2_U3080, P2_U3432);
  not ginst13743 (P2_R1215_U184, P2_R1215_U43);
  not ginst13744 (P2_R1215_U185, P2_R1215_U44);
  nand ginst13745 (P2_R1215_U186, P2_R1215_U43, P2_R1215_U44);
  nand ginst13746 (P2_R1215_U187, P2_R1215_U116, P2_R1215_U180);
  nand ginst13747 (P2_R1215_U188, P2_R1215_U186, P2_R1215_U5);
  nand ginst13748 (P2_R1215_U189, P2_U3066, P2_U3438);
  and ginst13749 (P2_R1215_U19, P2_R1215_U210, P2_R1215_U213);
  nand ginst13750 (P2_R1215_U190, P2_R1215_U117, P2_R1215_U188);
  nand ginst13751 (P2_R1215_U191, P2_R1215_U35, P2_R1215_U36);
  nand ginst13752 (P2_R1215_U192, P2_R1215_U191, P2_U3069);
  nand ginst13753 (P2_R1215_U193, P2_R1215_U190, P2_R1215_U4);
  nand ginst13754 (P2_R1215_U194, P2_R1215_U170, P2_U3444);
  not ginst13755 (P2_R1215_U195, P2_R1215_U42);
  or ginst13756 (P2_R1215_U196, P2_U3072, P2_U3450);
  or ginst13757 (P2_R1215_U197, P2_U3073, P2_U3447);
  not ginst13758 (P2_R1215_U198, P2_R1215_U23);
  nand ginst13759 (P2_R1215_U199, P2_R1215_U23, P2_R1215_U24);
  not ginst13760 (P2_R1215_U20, P2_U3447);
  nand ginst13761 (P2_R1215_U200, P2_R1215_U199, P2_U3072);
  nand ginst13762 (P2_R1215_U201, P2_R1215_U198, P2_U3450);
  nand ginst13763 (P2_R1215_U202, P2_R1215_U42, P2_R1215_U6);
  not ginst13764 (P2_R1215_U203, P2_R1215_U144);
  or ginst13765 (P2_R1215_U204, P2_U3086, P2_U3453);
  nand ginst13766 (P2_R1215_U205, P2_R1215_U144, P2_R1215_U204);
  not ginst13767 (P2_R1215_U206, P2_R1215_U41);
  or ginst13768 (P2_R1215_U207, P2_U3085, P2_U3456);
  or ginst13769 (P2_R1215_U208, P2_U3073, P2_U3447);
  nand ginst13770 (P2_R1215_U209, P2_R1215_U208, P2_R1215_U42);
  not ginst13771 (P2_R1215_U21, P2_U3073);
  nand ginst13772 (P2_R1215_U210, P2_R1215_U120, P2_R1215_U209);
  nand ginst13773 (P2_R1215_U211, P2_R1215_U195, P2_R1215_U23);
  nand ginst13774 (P2_R1215_U212, P2_U3072, P2_U3450);
  nand ginst13775 (P2_R1215_U213, P2_R1215_U121, P2_R1215_U211);
  or ginst13776 (P2_R1215_U214, P2_U3073, P2_U3447);
  nand ginst13777 (P2_R1215_U215, P2_R1215_U181, P2_R1215_U185);
  nand ginst13778 (P2_R1215_U216, P2_U3070, P2_U3435);
  not ginst13779 (P2_R1215_U217, P2_R1215_U46);
  nand ginst13780 (P2_R1215_U218, P2_R1215_U184, P2_R1215_U5);
  nand ginst13781 (P2_R1215_U219, P2_R1215_U180, P2_R1215_U46);
  not ginst13782 (P2_R1215_U22, P2_U3072);
  nand ginst13783 (P2_R1215_U220, P2_U3066, P2_U3438);
  not ginst13784 (P2_R1215_U221, P2_R1215_U45);
  or ginst13785 (P2_R1215_U222, P2_U3062, P2_U3441);
  nand ginst13786 (P2_R1215_U223, P2_R1215_U222, P2_R1215_U45);
  nand ginst13787 (P2_R1215_U224, P2_R1215_U123, P2_R1215_U223);
  nand ginst13788 (P2_R1215_U225, P2_R1215_U221, P2_R1215_U35);
  nand ginst13789 (P2_R1215_U226, P2_U3069, P2_U3444);
  nand ginst13790 (P2_R1215_U227, P2_R1215_U124, P2_R1215_U225);
  or ginst13791 (P2_R1215_U228, P2_U3062, P2_U3441);
  nand ginst13792 (P2_R1215_U229, P2_R1215_U181, P2_R1215_U184);
  nand ginst13793 (P2_R1215_U23, P2_U3073, P2_U3447);
  not ginst13794 (P2_R1215_U230, P2_R1215_U145);
  nand ginst13795 (P2_R1215_U231, P2_U3066, P2_U3438);
  nand ginst13796 (P2_R1215_U232, P2_R1215_U400, P2_R1215_U401, P2_R1215_U43, P2_R1215_U44);
  nand ginst13797 (P2_R1215_U233, P2_R1215_U43, P2_R1215_U44);
  nand ginst13798 (P2_R1215_U234, P2_U3070, P2_U3435);
  nand ginst13799 (P2_R1215_U235, P2_R1215_U125, P2_R1215_U233);
  or ginst13800 (P2_R1215_U236, P2_U3085, P2_U3456);
  or ginst13801 (P2_R1215_U237, P2_U3064, P2_U3459);
  nand ginst13802 (P2_R1215_U238, P2_R1215_U177, P2_R1215_U7);
  nand ginst13803 (P2_R1215_U239, P2_U3064, P2_U3459);
  not ginst13804 (P2_R1215_U24, P2_U3450);
  nand ginst13805 (P2_R1215_U240, P2_R1215_U127, P2_R1215_U238);
  or ginst13806 (P2_R1215_U241, P2_U3064, P2_U3459);
  nand ginst13807 (P2_R1215_U242, P2_R1215_U126, P2_R1215_U144);
  nand ginst13808 (P2_R1215_U243, P2_R1215_U240, P2_R1215_U241);
  not ginst13809 (P2_R1215_U244, P2_R1215_U167);
  or ginst13810 (P2_R1215_U245, P2_U3082, P2_U3468);
  or ginst13811 (P2_R1215_U246, P2_U3074, P2_U3465);
  nand ginst13812 (P2_R1215_U247, P2_R1215_U174, P2_R1215_U8);
  nand ginst13813 (P2_R1215_U248, P2_U3082, P2_U3468);
  nand ginst13814 (P2_R1215_U249, P2_R1215_U129, P2_R1215_U247);
  not ginst13815 (P2_R1215_U25, P2_U3441);
  or ginst13816 (P2_R1215_U250, P2_U3065, P2_U3462);
  or ginst13817 (P2_R1215_U251, P2_U3082, P2_U3468);
  nand ginst13818 (P2_R1215_U252, P2_R1215_U128, P2_R1215_U167);
  nand ginst13819 (P2_R1215_U253, P2_R1215_U249, P2_R1215_U251);
  not ginst13820 (P2_R1215_U254, P2_R1215_U166);
  or ginst13821 (P2_R1215_U255, P2_U3081, P2_U3471);
  nand ginst13822 (P2_R1215_U256, P2_R1215_U166, P2_R1215_U255);
  nand ginst13823 (P2_R1215_U257, P2_U3081, P2_U3471);
  not ginst13824 (P2_R1215_U258, P2_R1215_U164);
  or ginst13825 (P2_R1215_U259, P2_U3076, P2_U3474);
  not ginst13826 (P2_R1215_U26, P2_U3062);
  nand ginst13827 (P2_R1215_U260, P2_R1215_U164, P2_R1215_U259);
  nand ginst13828 (P2_R1215_U261, P2_U3076, P2_U3474);
  not ginst13829 (P2_R1215_U262, P2_R1215_U93);
  or ginst13830 (P2_R1215_U263, P2_U3071, P2_U3480);
  or ginst13831 (P2_R1215_U264, P2_U3075, P2_U3477);
  not ginst13832 (P2_R1215_U265, P2_R1215_U60);
  nand ginst13833 (P2_R1215_U266, P2_R1215_U60, P2_R1215_U61);
  nand ginst13834 (P2_R1215_U267, P2_R1215_U266, P2_U3071);
  nand ginst13835 (P2_R1215_U268, P2_R1215_U265, P2_U3480);
  nand ginst13836 (P2_R1215_U269, P2_R1215_U9, P2_R1215_U93);
  not ginst13837 (P2_R1215_U27, P2_U3069);
  not ginst13838 (P2_R1215_U270, P2_R1215_U162);
  or ginst13839 (P2_R1215_U271, P2_U3078, P2_U3957);
  or ginst13840 (P2_R1215_U272, P2_U3083, P2_U3485);
  or ginst13841 (P2_R1215_U273, P2_U3077, P2_U3956);
  not ginst13842 (P2_R1215_U274, P2_R1215_U81);
  nand ginst13843 (P2_R1215_U275, P2_R1215_U274, P2_U3957);
  nand ginst13844 (P2_R1215_U276, P2_R1215_U275, P2_R1215_U91);
  nand ginst13845 (P2_R1215_U277, P2_R1215_U81, P2_R1215_U82);
  nand ginst13846 (P2_R1215_U278, P2_R1215_U276, P2_R1215_U277);
  nand ginst13847 (P2_R1215_U279, P2_R1215_U10, P2_R1215_U175);
  not ginst13848 (P2_R1215_U28, P2_U3435);
  nand ginst13849 (P2_R1215_U280, P2_U3077, P2_U3956);
  nand ginst13850 (P2_R1215_U281, P2_R1215_U278, P2_R1215_U279);
  or ginst13851 (P2_R1215_U282, P2_U3084, P2_U3483);
  or ginst13852 (P2_R1215_U283, P2_U3077, P2_U3956);
  nand ginst13853 (P2_R1215_U284, P2_R1215_U131, P2_R1215_U162, P2_R1215_U273);
  nand ginst13854 (P2_R1215_U285, P2_R1215_U281, P2_R1215_U283);
  not ginst13855 (P2_R1215_U286, P2_R1215_U159);
  or ginst13856 (P2_R1215_U287, P2_U3063, P2_U3955);
  nand ginst13857 (P2_R1215_U288, P2_R1215_U159, P2_R1215_U287);
  nand ginst13858 (P2_R1215_U289, P2_U3063, P2_U3955);
  not ginst13859 (P2_R1215_U29, P2_U3070);
  not ginst13860 (P2_R1215_U290, P2_R1215_U157);
  or ginst13861 (P2_R1215_U291, P2_U3068, P2_U3954);
  nand ginst13862 (P2_R1215_U292, P2_R1215_U157, P2_R1215_U291);
  nand ginst13863 (P2_R1215_U293, P2_U3068, P2_U3954);
  not ginst13864 (P2_R1215_U294, P2_R1215_U155);
  or ginst13865 (P2_R1215_U295, P2_U3060, P2_U3952);
  nand ginst13866 (P2_R1215_U296, P2_R1215_U173, P2_R1215_U176);
  not ginst13867 (P2_R1215_U297, P2_R1215_U87);
  or ginst13868 (P2_R1215_U298, P2_U3067, P2_U3953);
  nand ginst13869 (P2_R1215_U299, P2_R1215_U155, P2_R1215_U168, P2_R1215_U298);
  not ginst13870 (P2_R1215_U30, P2_U3427);
  not ginst13871 (P2_R1215_U300, P2_R1215_U153);
  or ginst13872 (P2_R1215_U301, P2_U3055, P2_U3950);
  nand ginst13873 (P2_R1215_U302, P2_U3055, P2_U3950);
  not ginst13874 (P2_R1215_U303, P2_R1215_U151);
  nand ginst13875 (P2_R1215_U304, P2_R1215_U151, P2_U3949);
  not ginst13876 (P2_R1215_U305, P2_R1215_U149);
  nand ginst13877 (P2_R1215_U306, P2_R1215_U155, P2_R1215_U298);
  not ginst13878 (P2_R1215_U307, P2_R1215_U90);
  or ginst13879 (P2_R1215_U308, P2_U3060, P2_U3952);
  nand ginst13880 (P2_R1215_U309, P2_R1215_U308, P2_R1215_U90);
  not ginst13881 (P2_R1215_U31, P2_U3079);
  nand ginst13882 (P2_R1215_U310, P2_R1215_U154, P2_R1215_U173, P2_R1215_U309);
  nand ginst13883 (P2_R1215_U311, P2_R1215_U173, P2_R1215_U307);
  nand ginst13884 (P2_R1215_U312, P2_U3059, P2_U3951);
  nand ginst13885 (P2_R1215_U313, P2_R1215_U168, P2_R1215_U311, P2_R1215_U312);
  or ginst13886 (P2_R1215_U314, P2_U3060, P2_U3952);
  nand ginst13887 (P2_R1215_U315, P2_R1215_U162, P2_R1215_U282);
  not ginst13888 (P2_R1215_U316, P2_R1215_U92);
  nand ginst13889 (P2_R1215_U317, P2_R1215_U10, P2_R1215_U92);
  nand ginst13890 (P2_R1215_U318, P2_R1215_U135, P2_R1215_U317);
  nand ginst13891 (P2_R1215_U319, P2_R1215_U278, P2_R1215_U317);
  nand ginst13892 (P2_R1215_U32, P2_U3079, P2_U3427);
  nand ginst13893 (P2_R1215_U320, P2_R1215_U319, P2_R1215_U453);
  or ginst13894 (P2_R1215_U321, P2_U3083, P2_U3485);
  nand ginst13895 (P2_R1215_U322, P2_R1215_U321, P2_R1215_U92);
  nand ginst13896 (P2_R1215_U323, P2_R1215_U136, P2_R1215_U322);
  nand ginst13897 (P2_R1215_U324, P2_R1215_U316, P2_R1215_U81);
  nand ginst13898 (P2_R1215_U325, P2_U3078, P2_U3957);
  nand ginst13899 (P2_R1215_U326, P2_R1215_U137, P2_R1215_U324);
  or ginst13900 (P2_R1215_U327, P2_U3080, P2_U3432);
  not ginst13901 (P2_R1215_U328, P2_R1215_U161);
  or ginst13902 (P2_R1215_U329, P2_U3083, P2_U3485);
  not ginst13903 (P2_R1215_U33, P2_U3438);
  or ginst13904 (P2_R1215_U330, P2_U3075, P2_U3477);
  nand ginst13905 (P2_R1215_U331, P2_R1215_U330, P2_R1215_U93);
  nand ginst13906 (P2_R1215_U332, P2_R1215_U138, P2_R1215_U331);
  nand ginst13907 (P2_R1215_U333, P2_R1215_U262, P2_R1215_U60);
  nand ginst13908 (P2_R1215_U334, P2_U3071, P2_U3480);
  nand ginst13909 (P2_R1215_U335, P2_R1215_U139, P2_R1215_U333);
  or ginst13910 (P2_R1215_U336, P2_U3075, P2_U3477);
  nand ginst13911 (P2_R1215_U337, P2_R1215_U167, P2_R1215_U250);
  not ginst13912 (P2_R1215_U338, P2_R1215_U94);
  or ginst13913 (P2_R1215_U339, P2_U3074, P2_U3465);
  not ginst13914 (P2_R1215_U34, P2_U3066);
  nand ginst13915 (P2_R1215_U340, P2_R1215_U339, P2_R1215_U94);
  nand ginst13916 (P2_R1215_U341, P2_R1215_U140, P2_R1215_U340);
  nand ginst13917 (P2_R1215_U342, P2_R1215_U172, P2_R1215_U338);
  nand ginst13918 (P2_R1215_U343, P2_U3082, P2_U3468);
  nand ginst13919 (P2_R1215_U344, P2_R1215_U141, P2_R1215_U342);
  or ginst13920 (P2_R1215_U345, P2_U3074, P2_U3465);
  or ginst13921 (P2_R1215_U346, P2_U3085, P2_U3456);
  nand ginst13922 (P2_R1215_U347, P2_R1215_U346, P2_R1215_U41);
  nand ginst13923 (P2_R1215_U348, P2_R1215_U142, P2_R1215_U347);
  nand ginst13924 (P2_R1215_U349, P2_R1215_U171, P2_R1215_U206);
  nand ginst13925 (P2_R1215_U35, P2_U3062, P2_U3441);
  nand ginst13926 (P2_R1215_U350, P2_U3064, P2_U3459);
  nand ginst13927 (P2_R1215_U351, P2_R1215_U143, P2_R1215_U349);
  nand ginst13928 (P2_R1215_U352, P2_R1215_U171, P2_R1215_U207);
  nand ginst13929 (P2_R1215_U353, P2_R1215_U204, P2_R1215_U62);
  nand ginst13930 (P2_R1215_U354, P2_R1215_U214, P2_R1215_U23);
  nand ginst13931 (P2_R1215_U355, P2_R1215_U228, P2_R1215_U35);
  nand ginst13932 (P2_R1215_U356, P2_R1215_U180, P2_R1215_U231);
  nand ginst13933 (P2_R1215_U357, P2_R1215_U173, P2_R1215_U314);
  nand ginst13934 (P2_R1215_U358, P2_R1215_U176, P2_R1215_U298);
  nand ginst13935 (P2_R1215_U359, P2_R1215_U329, P2_R1215_U81);
  not ginst13936 (P2_R1215_U36, P2_U3444);
  nand ginst13937 (P2_R1215_U360, P2_R1215_U282, P2_R1215_U78);
  nand ginst13938 (P2_R1215_U361, P2_R1215_U336, P2_R1215_U60);
  nand ginst13939 (P2_R1215_U362, P2_R1215_U172, P2_R1215_U345);
  nand ginst13940 (P2_R1215_U363, P2_R1215_U250, P2_R1215_U69);
  nand ginst13941 (P2_R1215_U364, P2_U3056, P2_U3949);
  nand ginst13942 (P2_R1215_U365, P2_R1215_U168, P2_R1215_U296);
  nand ginst13943 (P2_R1215_U366, P2_R1215_U295, P2_U3059);
  nand ginst13944 (P2_R1215_U367, P2_R1215_U295, P2_U3951);
  nand ginst13945 (P2_R1215_U368, P2_R1215_U168, P2_R1215_U296, P2_R1215_U301);
  nand ginst13946 (P2_R1215_U369, P2_R1215_U133, P2_R1215_U155, P2_R1215_U168);
  not ginst13947 (P2_R1215_U37, P2_U3453);
  nand ginst13948 (P2_R1215_U370, P2_R1215_U297, P2_R1215_U301);
  nand ginst13949 (P2_R1215_U371, P2_R1215_U40, P2_U3085);
  nand ginst13950 (P2_R1215_U372, P2_R1215_U39, P2_U3456);
  nand ginst13951 (P2_R1215_U373, P2_R1215_U371, P2_R1215_U372);
  nand ginst13952 (P2_R1215_U374, P2_R1215_U352, P2_R1215_U41);
  nand ginst13953 (P2_R1215_U375, P2_R1215_U206, P2_R1215_U373);
  nand ginst13954 (P2_R1215_U376, P2_R1215_U37, P2_U3086);
  nand ginst13955 (P2_R1215_U377, P2_R1215_U38, P2_U3453);
  nand ginst13956 (P2_R1215_U378, P2_R1215_U376, P2_R1215_U377);
  nand ginst13957 (P2_R1215_U379, P2_R1215_U144, P2_R1215_U353);
  not ginst13958 (P2_R1215_U38, P2_U3086);
  nand ginst13959 (P2_R1215_U380, P2_R1215_U203, P2_R1215_U378);
  nand ginst13960 (P2_R1215_U381, P2_R1215_U24, P2_U3072);
  nand ginst13961 (P2_R1215_U382, P2_R1215_U22, P2_U3450);
  nand ginst13962 (P2_R1215_U383, P2_R1215_U20, P2_U3073);
  nand ginst13963 (P2_R1215_U384, P2_R1215_U21, P2_U3447);
  nand ginst13964 (P2_R1215_U385, P2_R1215_U383, P2_R1215_U384);
  nand ginst13965 (P2_R1215_U386, P2_R1215_U354, P2_R1215_U42);
  nand ginst13966 (P2_R1215_U387, P2_R1215_U195, P2_R1215_U385);
  nand ginst13967 (P2_R1215_U388, P2_R1215_U36, P2_U3069);
  nand ginst13968 (P2_R1215_U389, P2_R1215_U27, P2_U3444);
  not ginst13969 (P2_R1215_U39, P2_U3085);
  nand ginst13970 (P2_R1215_U390, P2_R1215_U25, P2_U3062);
  nand ginst13971 (P2_R1215_U391, P2_R1215_U26, P2_U3441);
  nand ginst13972 (P2_R1215_U392, P2_R1215_U390, P2_R1215_U391);
  nand ginst13973 (P2_R1215_U393, P2_R1215_U355, P2_R1215_U45);
  nand ginst13974 (P2_R1215_U394, P2_R1215_U221, P2_R1215_U392);
  nand ginst13975 (P2_R1215_U395, P2_R1215_U33, P2_U3066);
  nand ginst13976 (P2_R1215_U396, P2_R1215_U34, P2_U3438);
  nand ginst13977 (P2_R1215_U397, P2_R1215_U395, P2_R1215_U396);
  nand ginst13978 (P2_R1215_U398, P2_R1215_U145, P2_R1215_U356);
  nand ginst13979 (P2_R1215_U399, P2_R1215_U230, P2_R1215_U397);
  and ginst13980 (P2_R1215_U4, P2_R1215_U178, P2_R1215_U179);
  not ginst13981 (P2_R1215_U40, P2_U3456);
  nand ginst13982 (P2_R1215_U400, P2_R1215_U28, P2_U3070);
  nand ginst13983 (P2_R1215_U401, P2_R1215_U29, P2_U3435);
  nand ginst13984 (P2_R1215_U402, P2_R1215_U147, P2_U3057);
  nand ginst13985 (P2_R1215_U403, P2_R1215_U146, P2_U3960);
  nand ginst13986 (P2_R1215_U404, P2_R1215_U147, P2_U3057);
  nand ginst13987 (P2_R1215_U405, P2_R1215_U146, P2_U3960);
  nand ginst13988 (P2_R1215_U406, P2_R1215_U404, P2_R1215_U405);
  nand ginst13989 (P2_R1215_U407, P2_R1215_U148, P2_R1215_U149);
  nand ginst13990 (P2_R1215_U408, P2_R1215_U305, P2_R1215_U406);
  nand ginst13991 (P2_R1215_U409, P2_R1215_U89, P2_U3056);
  nand ginst13992 (P2_R1215_U41, P2_R1215_U205, P2_R1215_U62);
  nand ginst13993 (P2_R1215_U410, P2_R1215_U88, P2_U3949);
  nand ginst13994 (P2_R1215_U411, P2_R1215_U89, P2_U3056);
  nand ginst13995 (P2_R1215_U412, P2_R1215_U88, P2_U3949);
  nand ginst13996 (P2_R1215_U413, P2_R1215_U411, P2_R1215_U412);
  nand ginst13997 (P2_R1215_U414, P2_R1215_U150, P2_R1215_U151);
  nand ginst13998 (P2_R1215_U415, P2_R1215_U303, P2_R1215_U413);
  nand ginst13999 (P2_R1215_U416, P2_R1215_U47, P2_U3055);
  nand ginst14000 (P2_R1215_U417, P2_R1215_U48, P2_U3950);
  nand ginst14001 (P2_R1215_U418, P2_R1215_U47, P2_U3055);
  nand ginst14002 (P2_R1215_U419, P2_R1215_U48, P2_U3950);
  nand ginst14003 (P2_R1215_U42, P2_R1215_U118, P2_R1215_U193);
  nand ginst14004 (P2_R1215_U420, P2_R1215_U418, P2_R1215_U419);
  nand ginst14005 (P2_R1215_U421, P2_R1215_U152, P2_R1215_U153);
  nand ginst14006 (P2_R1215_U422, P2_R1215_U300, P2_R1215_U420);
  nand ginst14007 (P2_R1215_U423, P2_R1215_U50, P2_U3059);
  nand ginst14008 (P2_R1215_U424, P2_R1215_U49, P2_U3951);
  nand ginst14009 (P2_R1215_U425, P2_R1215_U51, P2_U3060);
  nand ginst14010 (P2_R1215_U426, P2_R1215_U52, P2_U3952);
  nand ginst14011 (P2_R1215_U427, P2_R1215_U425, P2_R1215_U426);
  nand ginst14012 (P2_R1215_U428, P2_R1215_U357, P2_R1215_U90);
  nand ginst14013 (P2_R1215_U429, P2_R1215_U307, P2_R1215_U427);
  nand ginst14014 (P2_R1215_U43, P2_R1215_U182, P2_R1215_U183);
  nand ginst14015 (P2_R1215_U430, P2_R1215_U53, P2_U3067);
  nand ginst14016 (P2_R1215_U431, P2_R1215_U54, P2_U3953);
  nand ginst14017 (P2_R1215_U432, P2_R1215_U430, P2_R1215_U431);
  nand ginst14018 (P2_R1215_U433, P2_R1215_U155, P2_R1215_U358);
  nand ginst14019 (P2_R1215_U434, P2_R1215_U294, P2_R1215_U432);
  nand ginst14020 (P2_R1215_U435, P2_R1215_U85, P2_U3068);
  nand ginst14021 (P2_R1215_U436, P2_R1215_U86, P2_U3954);
  nand ginst14022 (P2_R1215_U437, P2_R1215_U85, P2_U3068);
  nand ginst14023 (P2_R1215_U438, P2_R1215_U86, P2_U3954);
  nand ginst14024 (P2_R1215_U439, P2_R1215_U437, P2_R1215_U438);
  nand ginst14025 (P2_R1215_U44, P2_U3080, P2_U3432);
  nand ginst14026 (P2_R1215_U440, P2_R1215_U156, P2_R1215_U157);
  nand ginst14027 (P2_R1215_U441, P2_R1215_U290, P2_R1215_U439);
  nand ginst14028 (P2_R1215_U442, P2_R1215_U83, P2_U3063);
  nand ginst14029 (P2_R1215_U443, P2_R1215_U84, P2_U3955);
  nand ginst14030 (P2_R1215_U444, P2_R1215_U83, P2_U3063);
  nand ginst14031 (P2_R1215_U445, P2_R1215_U84, P2_U3955);
  nand ginst14032 (P2_R1215_U446, P2_R1215_U444, P2_R1215_U445);
  nand ginst14033 (P2_R1215_U447, P2_R1215_U158, P2_R1215_U159);
  nand ginst14034 (P2_R1215_U448, P2_R1215_U286, P2_R1215_U446);
  nand ginst14035 (P2_R1215_U449, P2_R1215_U55, P2_U3077);
  nand ginst14036 (P2_R1215_U45, P2_R1215_U122, P2_R1215_U219);
  nand ginst14037 (P2_R1215_U450, P2_R1215_U56, P2_U3956);
  nand ginst14038 (P2_R1215_U451, P2_R1215_U55, P2_U3077);
  nand ginst14039 (P2_R1215_U452, P2_R1215_U56, P2_U3956);
  nand ginst14040 (P2_R1215_U453, P2_R1215_U451, P2_R1215_U452);
  nand ginst14041 (P2_R1215_U454, P2_R1215_U82, P2_U3078);
  nand ginst14042 (P2_R1215_U455, P2_R1215_U91, P2_U3957);
  nand ginst14043 (P2_R1215_U456, P2_R1215_U161, P2_R1215_U182);
  nand ginst14044 (P2_R1215_U457, P2_R1215_U32, P2_R1215_U328);
  nand ginst14045 (P2_R1215_U458, P2_R1215_U79, P2_U3083);
  nand ginst14046 (P2_R1215_U459, P2_R1215_U80, P2_U3485);
  nand ginst14047 (P2_R1215_U46, P2_R1215_U215, P2_R1215_U216);
  nand ginst14048 (P2_R1215_U460, P2_R1215_U458, P2_R1215_U459);
  nand ginst14049 (P2_R1215_U461, P2_R1215_U359, P2_R1215_U92);
  nand ginst14050 (P2_R1215_U462, P2_R1215_U316, P2_R1215_U460);
  nand ginst14051 (P2_R1215_U463, P2_R1215_U76, P2_U3084);
  nand ginst14052 (P2_R1215_U464, P2_R1215_U77, P2_U3483);
  nand ginst14053 (P2_R1215_U465, P2_R1215_U463, P2_R1215_U464);
  nand ginst14054 (P2_R1215_U466, P2_R1215_U162, P2_R1215_U360);
  nand ginst14055 (P2_R1215_U467, P2_R1215_U270, P2_R1215_U465);
  nand ginst14056 (P2_R1215_U468, P2_R1215_U61, P2_U3071);
  nand ginst14057 (P2_R1215_U469, P2_R1215_U59, P2_U3480);
  not ginst14058 (P2_R1215_U47, P2_U3950);
  nand ginst14059 (P2_R1215_U470, P2_R1215_U57, P2_U3075);
  nand ginst14060 (P2_R1215_U471, P2_R1215_U58, P2_U3477);
  nand ginst14061 (P2_R1215_U472, P2_R1215_U470, P2_R1215_U471);
  nand ginst14062 (P2_R1215_U473, P2_R1215_U361, P2_R1215_U93);
  nand ginst14063 (P2_R1215_U474, P2_R1215_U262, P2_R1215_U472);
  nand ginst14064 (P2_R1215_U475, P2_R1215_U74, P2_U3076);
  nand ginst14065 (P2_R1215_U476, P2_R1215_U75, P2_U3474);
  nand ginst14066 (P2_R1215_U477, P2_R1215_U74, P2_U3076);
  nand ginst14067 (P2_R1215_U478, P2_R1215_U75, P2_U3474);
  nand ginst14068 (P2_R1215_U479, P2_R1215_U477, P2_R1215_U478);
  not ginst14069 (P2_R1215_U48, P2_U3055);
  nand ginst14070 (P2_R1215_U480, P2_R1215_U163, P2_R1215_U164);
  nand ginst14071 (P2_R1215_U481, P2_R1215_U258, P2_R1215_U479);
  nand ginst14072 (P2_R1215_U482, P2_R1215_U72, P2_U3081);
  nand ginst14073 (P2_R1215_U483, P2_R1215_U73, P2_U3471);
  nand ginst14074 (P2_R1215_U484, P2_R1215_U72, P2_U3081);
  nand ginst14075 (P2_R1215_U485, P2_R1215_U73, P2_U3471);
  nand ginst14076 (P2_R1215_U486, P2_R1215_U484, P2_R1215_U485);
  nand ginst14077 (P2_R1215_U487, P2_R1215_U165, P2_R1215_U166);
  nand ginst14078 (P2_R1215_U488, P2_R1215_U254, P2_R1215_U486);
  nand ginst14079 (P2_R1215_U489, P2_R1215_U70, P2_U3082);
  not ginst14080 (P2_R1215_U49, P2_U3059);
  nand ginst14081 (P2_R1215_U490, P2_R1215_U71, P2_U3468);
  nand ginst14082 (P2_R1215_U491, P2_R1215_U65, P2_U3074);
  nand ginst14083 (P2_R1215_U492, P2_R1215_U66, P2_U3465);
  nand ginst14084 (P2_R1215_U493, P2_R1215_U491, P2_R1215_U492);
  nand ginst14085 (P2_R1215_U494, P2_R1215_U362, P2_R1215_U94);
  nand ginst14086 (P2_R1215_U495, P2_R1215_U338, P2_R1215_U493);
  nand ginst14087 (P2_R1215_U496, P2_R1215_U67, P2_U3065);
  nand ginst14088 (P2_R1215_U497, P2_R1215_U68, P2_U3462);
  nand ginst14089 (P2_R1215_U498, P2_R1215_U496, P2_R1215_U497);
  nand ginst14090 (P2_R1215_U499, P2_R1215_U167, P2_R1215_U363);
  and ginst14091 (P2_R1215_U5, P2_R1215_U180, P2_R1215_U181);
  not ginst14092 (P2_R1215_U50, P2_U3951);
  nand ginst14093 (P2_R1215_U500, P2_R1215_U244, P2_R1215_U498);
  nand ginst14094 (P2_R1215_U501, P2_R1215_U63, P2_U3064);
  nand ginst14095 (P2_R1215_U502, P2_R1215_U64, P2_U3459);
  nand ginst14096 (P2_R1215_U503, P2_R1215_U30, P2_U3079);
  nand ginst14097 (P2_R1215_U504, P2_R1215_U31, P2_U3427);
  not ginst14098 (P2_R1215_U51, P2_U3952);
  not ginst14099 (P2_R1215_U52, P2_U3060);
  not ginst14100 (P2_R1215_U53, P2_U3953);
  not ginst14101 (P2_R1215_U54, P2_U3067);
  not ginst14102 (P2_R1215_U55, P2_U3956);
  not ginst14103 (P2_R1215_U56, P2_U3077);
  not ginst14104 (P2_R1215_U57, P2_U3477);
  not ginst14105 (P2_R1215_U58, P2_U3075);
  not ginst14106 (P2_R1215_U59, P2_U3071);
  and ginst14107 (P2_R1215_U6, P2_R1215_U196, P2_R1215_U197);
  nand ginst14108 (P2_R1215_U60, P2_U3075, P2_U3477);
  not ginst14109 (P2_R1215_U61, P2_U3480);
  nand ginst14110 (P2_R1215_U62, P2_U3086, P2_U3453);
  not ginst14111 (P2_R1215_U63, P2_U3459);
  not ginst14112 (P2_R1215_U64, P2_U3064);
  not ginst14113 (P2_R1215_U65, P2_U3465);
  not ginst14114 (P2_R1215_U66, P2_U3074);
  not ginst14115 (P2_R1215_U67, P2_U3462);
  not ginst14116 (P2_R1215_U68, P2_U3065);
  nand ginst14117 (P2_R1215_U69, P2_U3065, P2_U3462);
  and ginst14118 (P2_R1215_U7, P2_R1215_U236, P2_R1215_U237);
  not ginst14119 (P2_R1215_U70, P2_U3468);
  not ginst14120 (P2_R1215_U71, P2_U3082);
  not ginst14121 (P2_R1215_U72, P2_U3471);
  not ginst14122 (P2_R1215_U73, P2_U3081);
  not ginst14123 (P2_R1215_U74, P2_U3474);
  not ginst14124 (P2_R1215_U75, P2_U3076);
  not ginst14125 (P2_R1215_U76, P2_U3483);
  not ginst14126 (P2_R1215_U77, P2_U3084);
  nand ginst14127 (P2_R1215_U78, P2_U3084, P2_U3483);
  not ginst14128 (P2_R1215_U79, P2_U3485);
  and ginst14129 (P2_R1215_U8, P2_R1215_U245, P2_R1215_U246);
  not ginst14130 (P2_R1215_U80, P2_U3083);
  nand ginst14131 (P2_R1215_U81, P2_U3083, P2_U3485);
  not ginst14132 (P2_R1215_U82, P2_U3957);
  not ginst14133 (P2_R1215_U83, P2_U3955);
  not ginst14134 (P2_R1215_U84, P2_U3063);
  not ginst14135 (P2_R1215_U85, P2_U3954);
  not ginst14136 (P2_R1215_U86, P2_U3068);
  nand ginst14137 (P2_R1215_U87, P2_U3059, P2_U3951);
  not ginst14138 (P2_R1215_U88, P2_U3056);
  not ginst14139 (P2_R1215_U89, P2_U3949);
  and ginst14140 (P2_R1215_U9, P2_R1215_U263, P2_R1215_U264);
  nand ginst14141 (P2_R1215_U90, P2_R1215_U176, P2_R1215_U306);
  not ginst14142 (P2_R1215_U91, P2_U3078);
  nand ginst14143 (P2_R1215_U92, P2_R1215_U315, P2_R1215_U78);
  nand ginst14144 (P2_R1215_U93, P2_R1215_U260, P2_R1215_U261);
  nand ginst14145 (P2_R1215_U94, P2_R1215_U337, P2_R1215_U69);
  nand ginst14146 (P2_R1215_U95, P2_R1215_U456, P2_R1215_U457);
  nand ginst14147 (P2_R1215_U96, P2_R1215_U503, P2_R1215_U504);
  nand ginst14148 (P2_R1215_U97, P2_R1215_U374, P2_R1215_U375);
  nand ginst14149 (P2_R1215_U98, P2_R1215_U379, P2_R1215_U380);
  nand ginst14150 (P2_R1215_U99, P2_R1215_U386, P2_R1215_U387);
  and ginst14151 (P2_R1233_U10, P2_R1233_U348, P2_R1233_U351);
  nand ginst14152 (P2_R1233_U100, P2_R1233_U398, P2_R1233_U399);
  nand ginst14153 (P2_R1233_U101, P2_R1233_U407, P2_R1233_U408);
  nand ginst14154 (P2_R1233_U102, P2_R1233_U414, P2_R1233_U415);
  nand ginst14155 (P2_R1233_U103, P2_R1233_U421, P2_R1233_U422);
  nand ginst14156 (P2_R1233_U104, P2_R1233_U428, P2_R1233_U429);
  nand ginst14157 (P2_R1233_U105, P2_R1233_U433, P2_R1233_U434);
  nand ginst14158 (P2_R1233_U106, P2_R1233_U440, P2_R1233_U441);
  nand ginst14159 (P2_R1233_U107, P2_R1233_U447, P2_R1233_U448);
  nand ginst14160 (P2_R1233_U108, P2_R1233_U461, P2_R1233_U462);
  nand ginst14161 (P2_R1233_U109, P2_R1233_U466, P2_R1233_U467);
  and ginst14162 (P2_R1233_U11, P2_R1233_U341, P2_R1233_U344);
  nand ginst14163 (P2_R1233_U110, P2_R1233_U473, P2_R1233_U474);
  nand ginst14164 (P2_R1233_U111, P2_R1233_U480, P2_R1233_U481);
  nand ginst14165 (P2_R1233_U112, P2_R1233_U487, P2_R1233_U488);
  nand ginst14166 (P2_R1233_U113, P2_R1233_U494, P2_R1233_U495);
  nand ginst14167 (P2_R1233_U114, P2_R1233_U499, P2_R1233_U500);
  and ginst14168 (P2_R1233_U115, P2_R1233_U187, P2_R1233_U189);
  and ginst14169 (P2_R1233_U116, P2_R1233_U180, P2_R1233_U4);
  and ginst14170 (P2_R1233_U117, P2_R1233_U192, P2_R1233_U194);
  and ginst14171 (P2_R1233_U118, P2_R1233_U200, P2_R1233_U201);
  and ginst14172 (P2_R1233_U119, P2_R1233_U22, P2_R1233_U381, P2_R1233_U382);
  and ginst14173 (P2_R1233_U12, P2_R1233_U332, P2_R1233_U335);
  and ginst14174 (P2_R1233_U120, P2_R1233_U212, P2_R1233_U5);
  and ginst14175 (P2_R1233_U121, P2_R1233_U180, P2_R1233_U181);
  and ginst14176 (P2_R1233_U122, P2_R1233_U218, P2_R1233_U220);
  and ginst14177 (P2_R1233_U123, P2_R1233_U34, P2_R1233_U388, P2_R1233_U389);
  and ginst14178 (P2_R1233_U124, P2_R1233_U226, P2_R1233_U4);
  and ginst14179 (P2_R1233_U125, P2_R1233_U181, P2_R1233_U234);
  and ginst14180 (P2_R1233_U126, P2_R1233_U204, P2_R1233_U6);
  and ginst14181 (P2_R1233_U127, P2_R1233_U171, P2_R1233_U239);
  and ginst14182 (P2_R1233_U128, P2_R1233_U250, P2_R1233_U7);
  and ginst14183 (P2_R1233_U129, P2_R1233_U172, P2_R1233_U248);
  and ginst14184 (P2_R1233_U13, P2_R1233_U323, P2_R1233_U326);
  and ginst14185 (P2_R1233_U130, P2_R1233_U267, P2_R1233_U268);
  and ginst14186 (P2_R1233_U131, P2_R1233_U282, P2_R1233_U9);
  and ginst14187 (P2_R1233_U132, P2_R1233_U280, P2_R1233_U285);
  and ginst14188 (P2_R1233_U133, P2_R1233_U298, P2_R1233_U301);
  and ginst14189 (P2_R1233_U134, P2_R1233_U302, P2_R1233_U368);
  and ginst14190 (P2_R1233_U135, P2_R1233_U160, P2_R1233_U278);
  and ginst14191 (P2_R1233_U136, P2_R1233_U454, P2_R1233_U455, P2_R1233_U80);
  and ginst14192 (P2_R1233_U137, P2_R1233_U325, P2_R1233_U9);
  and ginst14193 (P2_R1233_U138, P2_R1233_U468, P2_R1233_U469, P2_R1233_U59);
  and ginst14194 (P2_R1233_U139, P2_R1233_U334, P2_R1233_U8);
  and ginst14195 (P2_R1233_U14, P2_R1233_U318, P2_R1233_U320);
  and ginst14196 (P2_R1233_U140, P2_R1233_U172, P2_R1233_U489, P2_R1233_U490);
  and ginst14197 (P2_R1233_U141, P2_R1233_U343, P2_R1233_U7);
  and ginst14198 (P2_R1233_U142, P2_R1233_U171, P2_R1233_U501, P2_R1233_U502);
  and ginst14199 (P2_R1233_U143, P2_R1233_U350, P2_R1233_U6);
  nand ginst14200 (P2_R1233_U144, P2_R1233_U118, P2_R1233_U202);
  nand ginst14201 (P2_R1233_U145, P2_R1233_U217, P2_R1233_U229);
  not ginst14202 (P2_R1233_U146, P2_U3057);
  not ginst14203 (P2_R1233_U147, P2_U3960);
  and ginst14204 (P2_R1233_U148, P2_R1233_U402, P2_R1233_U403);
  nand ginst14205 (P2_R1233_U149, P2_R1233_U169, P2_R1233_U304, P2_R1233_U364);
  and ginst14206 (P2_R1233_U15, P2_R1233_U310, P2_R1233_U313);
  and ginst14207 (P2_R1233_U150, P2_R1233_U409, P2_R1233_U410);
  nand ginst14208 (P2_R1233_U151, P2_R1233_U134, P2_R1233_U369, P2_R1233_U370);
  and ginst14209 (P2_R1233_U152, P2_R1233_U416, P2_R1233_U417);
  nand ginst14210 (P2_R1233_U153, P2_R1233_U299, P2_R1233_U365, P2_R1233_U86);
  and ginst14211 (P2_R1233_U154, P2_R1233_U423, P2_R1233_U424);
  nand ginst14212 (P2_R1233_U155, P2_R1233_U292, P2_R1233_U293);
  and ginst14213 (P2_R1233_U156, P2_R1233_U435, P2_R1233_U436);
  nand ginst14214 (P2_R1233_U157, P2_R1233_U288, P2_R1233_U289);
  and ginst14215 (P2_R1233_U158, P2_R1233_U442, P2_R1233_U443);
  nand ginst14216 (P2_R1233_U159, P2_R1233_U132, P2_R1233_U284);
  and ginst14217 (P2_R1233_U16, P2_R1233_U232, P2_R1233_U235);
  and ginst14218 (P2_R1233_U160, P2_R1233_U449, P2_R1233_U450);
  nand ginst14219 (P2_R1233_U161, P2_R1233_U327, P2_R1233_U43);
  nand ginst14220 (P2_R1233_U162, P2_R1233_U130, P2_R1233_U269);
  and ginst14221 (P2_R1233_U163, P2_R1233_U475, P2_R1233_U476);
  nand ginst14222 (P2_R1233_U164, P2_R1233_U256, P2_R1233_U257);
  and ginst14223 (P2_R1233_U165, P2_R1233_U482, P2_R1233_U483);
  nand ginst14224 (P2_R1233_U166, P2_R1233_U252, P2_R1233_U253);
  nand ginst14225 (P2_R1233_U167, P2_R1233_U242, P2_R1233_U243);
  nand ginst14226 (P2_R1233_U168, P2_R1233_U366, P2_R1233_U367);
  nand ginst14227 (P2_R1233_U169, P2_R1233_U151, P2_U3056);
  and ginst14228 (P2_R1233_U17, P2_R1233_U224, P2_R1233_U227);
  not ginst14229 (P2_R1233_U170, P2_R1233_U34);
  nand ginst14230 (P2_R1233_U171, P2_U3085, P2_U3456);
  nand ginst14231 (P2_R1233_U172, P2_U3074, P2_U3465);
  nand ginst14232 (P2_R1233_U173, P2_U3060, P2_U3952);
  not ginst14233 (P2_R1233_U174, P2_R1233_U68);
  not ginst14234 (P2_R1233_U175, P2_R1233_U77);
  nand ginst14235 (P2_R1233_U176, P2_U3067, P2_U3953);
  not ginst14236 (P2_R1233_U177, P2_R1233_U61);
  or ginst14237 (P2_R1233_U178, P2_U3069, P2_U3444);
  or ginst14238 (P2_R1233_U179, P2_U3062, P2_U3441);
  and ginst14239 (P2_R1233_U18, P2_R1233_U210, P2_R1233_U213);
  or ginst14240 (P2_R1233_U180, P2_U3066, P2_U3438);
  or ginst14241 (P2_R1233_U181, P2_U3070, P2_U3435);
  not ginst14242 (P2_R1233_U182, P2_R1233_U31);
  or ginst14243 (P2_R1233_U183, P2_U3080, P2_U3432);
  not ginst14244 (P2_R1233_U184, P2_R1233_U42);
  not ginst14245 (P2_R1233_U185, P2_R1233_U43);
  nand ginst14246 (P2_R1233_U186, P2_R1233_U42, P2_R1233_U43);
  nand ginst14247 (P2_R1233_U187, P2_U3070, P2_U3435);
  nand ginst14248 (P2_R1233_U188, P2_R1233_U181, P2_R1233_U186);
  nand ginst14249 (P2_R1233_U189, P2_U3066, P2_U3438);
  not ginst14250 (P2_R1233_U19, P2_U3447);
  nand ginst14251 (P2_R1233_U190, P2_R1233_U115, P2_R1233_U188);
  nand ginst14252 (P2_R1233_U191, P2_R1233_U34, P2_R1233_U35);
  nand ginst14253 (P2_R1233_U192, P2_R1233_U191, P2_U3069);
  nand ginst14254 (P2_R1233_U193, P2_R1233_U116, P2_R1233_U190);
  nand ginst14255 (P2_R1233_U194, P2_R1233_U170, P2_U3444);
  not ginst14256 (P2_R1233_U195, P2_R1233_U41);
  or ginst14257 (P2_R1233_U196, P2_U3072, P2_U3450);
  or ginst14258 (P2_R1233_U197, P2_U3073, P2_U3447);
  not ginst14259 (P2_R1233_U198, P2_R1233_U22);
  nand ginst14260 (P2_R1233_U199, P2_R1233_U22, P2_R1233_U23);
  not ginst14261 (P2_R1233_U20, P2_U3073);
  nand ginst14262 (P2_R1233_U200, P2_R1233_U199, P2_U3072);
  nand ginst14263 (P2_R1233_U201, P2_R1233_U198, P2_U3450);
  nand ginst14264 (P2_R1233_U202, P2_R1233_U41, P2_R1233_U5);
  not ginst14265 (P2_R1233_U203, P2_R1233_U144);
  or ginst14266 (P2_R1233_U204, P2_U3086, P2_U3453);
  nand ginst14267 (P2_R1233_U205, P2_R1233_U144, P2_R1233_U204);
  not ginst14268 (P2_R1233_U206, P2_R1233_U40);
  or ginst14269 (P2_R1233_U207, P2_U3085, P2_U3456);
  or ginst14270 (P2_R1233_U208, P2_U3073, P2_U3447);
  nand ginst14271 (P2_R1233_U209, P2_R1233_U208, P2_R1233_U41);
  not ginst14272 (P2_R1233_U21, P2_U3072);
  nand ginst14273 (P2_R1233_U210, P2_R1233_U119, P2_R1233_U209);
  nand ginst14274 (P2_R1233_U211, P2_R1233_U195, P2_R1233_U22);
  nand ginst14275 (P2_R1233_U212, P2_U3072, P2_U3450);
  nand ginst14276 (P2_R1233_U213, P2_R1233_U120, P2_R1233_U211);
  or ginst14277 (P2_R1233_U214, P2_U3073, P2_U3447);
  nand ginst14278 (P2_R1233_U215, P2_R1233_U181, P2_R1233_U185);
  nand ginst14279 (P2_R1233_U216, P2_U3070, P2_U3435);
  not ginst14280 (P2_R1233_U217, P2_R1233_U45);
  nand ginst14281 (P2_R1233_U218, P2_R1233_U121, P2_R1233_U184);
  nand ginst14282 (P2_R1233_U219, P2_R1233_U180, P2_R1233_U45);
  nand ginst14283 (P2_R1233_U22, P2_U3073, P2_U3447);
  nand ginst14284 (P2_R1233_U220, P2_U3066, P2_U3438);
  not ginst14285 (P2_R1233_U221, P2_R1233_U44);
  or ginst14286 (P2_R1233_U222, P2_U3062, P2_U3441);
  nand ginst14287 (P2_R1233_U223, P2_R1233_U222, P2_R1233_U44);
  nand ginst14288 (P2_R1233_U224, P2_R1233_U123, P2_R1233_U223);
  nand ginst14289 (P2_R1233_U225, P2_R1233_U221, P2_R1233_U34);
  nand ginst14290 (P2_R1233_U226, P2_U3069, P2_U3444);
  nand ginst14291 (P2_R1233_U227, P2_R1233_U124, P2_R1233_U225);
  or ginst14292 (P2_R1233_U228, P2_U3062, P2_U3441);
  nand ginst14293 (P2_R1233_U229, P2_R1233_U181, P2_R1233_U184);
  not ginst14294 (P2_R1233_U23, P2_U3450);
  not ginst14295 (P2_R1233_U230, P2_R1233_U145);
  nand ginst14296 (P2_R1233_U231, P2_U3066, P2_U3438);
  nand ginst14297 (P2_R1233_U232, P2_R1233_U400, P2_R1233_U401, P2_R1233_U42, P2_R1233_U43);
  nand ginst14298 (P2_R1233_U233, P2_R1233_U42, P2_R1233_U43);
  nand ginst14299 (P2_R1233_U234, P2_U3070, P2_U3435);
  nand ginst14300 (P2_R1233_U235, P2_R1233_U125, P2_R1233_U233);
  or ginst14301 (P2_R1233_U236, P2_U3085, P2_U3456);
  or ginst14302 (P2_R1233_U237, P2_U3064, P2_U3459);
  nand ginst14303 (P2_R1233_U238, P2_R1233_U177, P2_R1233_U6);
  nand ginst14304 (P2_R1233_U239, P2_U3064, P2_U3459);
  not ginst14305 (P2_R1233_U24, P2_U3441);
  nand ginst14306 (P2_R1233_U240, P2_R1233_U127, P2_R1233_U238);
  or ginst14307 (P2_R1233_U241, P2_U3064, P2_U3459);
  nand ginst14308 (P2_R1233_U242, P2_R1233_U126, P2_R1233_U144);
  nand ginst14309 (P2_R1233_U243, P2_R1233_U240, P2_R1233_U241);
  not ginst14310 (P2_R1233_U244, P2_R1233_U167);
  or ginst14311 (P2_R1233_U245, P2_U3082, P2_U3468);
  or ginst14312 (P2_R1233_U246, P2_U3074, P2_U3465);
  nand ginst14313 (P2_R1233_U247, P2_R1233_U174, P2_R1233_U7);
  nand ginst14314 (P2_R1233_U248, P2_U3082, P2_U3468);
  nand ginst14315 (P2_R1233_U249, P2_R1233_U129, P2_R1233_U247);
  not ginst14316 (P2_R1233_U25, P2_U3062);
  or ginst14317 (P2_R1233_U250, P2_U3065, P2_U3462);
  or ginst14318 (P2_R1233_U251, P2_U3082, P2_U3468);
  nand ginst14319 (P2_R1233_U252, P2_R1233_U128, P2_R1233_U167);
  nand ginst14320 (P2_R1233_U253, P2_R1233_U249, P2_R1233_U251);
  not ginst14321 (P2_R1233_U254, P2_R1233_U166);
  or ginst14322 (P2_R1233_U255, P2_U3081, P2_U3471);
  nand ginst14323 (P2_R1233_U256, P2_R1233_U166, P2_R1233_U255);
  nand ginst14324 (P2_R1233_U257, P2_U3081, P2_U3471);
  not ginst14325 (P2_R1233_U258, P2_R1233_U164);
  or ginst14326 (P2_R1233_U259, P2_U3076, P2_U3474);
  not ginst14327 (P2_R1233_U26, P2_U3069);
  nand ginst14328 (P2_R1233_U260, P2_R1233_U164, P2_R1233_U259);
  nand ginst14329 (P2_R1233_U261, P2_U3076, P2_U3474);
  not ginst14330 (P2_R1233_U262, P2_R1233_U92);
  or ginst14331 (P2_R1233_U263, P2_U3071, P2_U3480);
  or ginst14332 (P2_R1233_U264, P2_U3075, P2_U3477);
  not ginst14333 (P2_R1233_U265, P2_R1233_U59);
  nand ginst14334 (P2_R1233_U266, P2_R1233_U59, P2_R1233_U60);
  nand ginst14335 (P2_R1233_U267, P2_R1233_U266, P2_U3071);
  nand ginst14336 (P2_R1233_U268, P2_R1233_U265, P2_U3480);
  nand ginst14337 (P2_R1233_U269, P2_R1233_U8, P2_R1233_U92);
  not ginst14338 (P2_R1233_U27, P2_U3435);
  not ginst14339 (P2_R1233_U270, P2_R1233_U162);
  or ginst14340 (P2_R1233_U271, P2_U3078, P2_U3957);
  or ginst14341 (P2_R1233_U272, P2_U3083, P2_U3485);
  or ginst14342 (P2_R1233_U273, P2_U3077, P2_U3956);
  not ginst14343 (P2_R1233_U274, P2_R1233_U80);
  nand ginst14344 (P2_R1233_U275, P2_R1233_U274, P2_U3957);
  nand ginst14345 (P2_R1233_U276, P2_R1233_U275, P2_R1233_U90);
  nand ginst14346 (P2_R1233_U277, P2_R1233_U80, P2_R1233_U81);
  nand ginst14347 (P2_R1233_U278, P2_R1233_U276, P2_R1233_U277);
  nand ginst14348 (P2_R1233_U279, P2_R1233_U175, P2_R1233_U9);
  not ginst14349 (P2_R1233_U28, P2_U3070);
  nand ginst14350 (P2_R1233_U280, P2_U3077, P2_U3956);
  nand ginst14351 (P2_R1233_U281, P2_R1233_U278, P2_R1233_U279);
  or ginst14352 (P2_R1233_U282, P2_U3084, P2_U3483);
  or ginst14353 (P2_R1233_U283, P2_U3077, P2_U3956);
  nand ginst14354 (P2_R1233_U284, P2_R1233_U131, P2_R1233_U162, P2_R1233_U273);
  nand ginst14355 (P2_R1233_U285, P2_R1233_U281, P2_R1233_U283);
  not ginst14356 (P2_R1233_U286, P2_R1233_U159);
  or ginst14357 (P2_R1233_U287, P2_U3063, P2_U3955);
  nand ginst14358 (P2_R1233_U288, P2_R1233_U159, P2_R1233_U287);
  nand ginst14359 (P2_R1233_U289, P2_U3063, P2_U3955);
  not ginst14360 (P2_R1233_U29, P2_U3427);
  not ginst14361 (P2_R1233_U290, P2_R1233_U157);
  or ginst14362 (P2_R1233_U291, P2_U3068, P2_U3954);
  nand ginst14363 (P2_R1233_U292, P2_R1233_U157, P2_R1233_U291);
  nand ginst14364 (P2_R1233_U293, P2_U3068, P2_U3954);
  not ginst14365 (P2_R1233_U294, P2_R1233_U155);
  or ginst14366 (P2_R1233_U295, P2_U3060, P2_U3952);
  nand ginst14367 (P2_R1233_U296, P2_R1233_U173, P2_R1233_U176);
  not ginst14368 (P2_R1233_U297, P2_R1233_U86);
  or ginst14369 (P2_R1233_U298, P2_U3067, P2_U3953);
  nand ginst14370 (P2_R1233_U299, P2_R1233_U155, P2_R1233_U168, P2_R1233_U298);
  not ginst14371 (P2_R1233_U30, P2_U3079);
  not ginst14372 (P2_R1233_U300, P2_R1233_U153);
  or ginst14373 (P2_R1233_U301, P2_U3055, P2_U3950);
  nand ginst14374 (P2_R1233_U302, P2_U3055, P2_U3950);
  not ginst14375 (P2_R1233_U303, P2_R1233_U151);
  nand ginst14376 (P2_R1233_U304, P2_R1233_U151, P2_U3949);
  not ginst14377 (P2_R1233_U305, P2_R1233_U149);
  nand ginst14378 (P2_R1233_U306, P2_R1233_U155, P2_R1233_U298);
  not ginst14379 (P2_R1233_U307, P2_R1233_U89);
  or ginst14380 (P2_R1233_U308, P2_U3060, P2_U3952);
  nand ginst14381 (P2_R1233_U309, P2_R1233_U308, P2_R1233_U89);
  nand ginst14382 (P2_R1233_U31, P2_U3079, P2_U3427);
  nand ginst14383 (P2_R1233_U310, P2_R1233_U154, P2_R1233_U173, P2_R1233_U309);
  nand ginst14384 (P2_R1233_U311, P2_R1233_U173, P2_R1233_U307);
  nand ginst14385 (P2_R1233_U312, P2_U3059, P2_U3951);
  nand ginst14386 (P2_R1233_U313, P2_R1233_U168, P2_R1233_U311, P2_R1233_U312);
  or ginst14387 (P2_R1233_U314, P2_U3060, P2_U3952);
  nand ginst14388 (P2_R1233_U315, P2_R1233_U162, P2_R1233_U282);
  not ginst14389 (P2_R1233_U316, P2_R1233_U91);
  nand ginst14390 (P2_R1233_U317, P2_R1233_U9, P2_R1233_U91);
  nand ginst14391 (P2_R1233_U318, P2_R1233_U135, P2_R1233_U317);
  nand ginst14392 (P2_R1233_U319, P2_R1233_U278, P2_R1233_U317);
  not ginst14393 (P2_R1233_U32, P2_U3438);
  nand ginst14394 (P2_R1233_U320, P2_R1233_U319, P2_R1233_U453);
  or ginst14395 (P2_R1233_U321, P2_U3083, P2_U3485);
  nand ginst14396 (P2_R1233_U322, P2_R1233_U321, P2_R1233_U91);
  nand ginst14397 (P2_R1233_U323, P2_R1233_U136, P2_R1233_U322);
  nand ginst14398 (P2_R1233_U324, P2_R1233_U316, P2_R1233_U80);
  nand ginst14399 (P2_R1233_U325, P2_U3078, P2_U3957);
  nand ginst14400 (P2_R1233_U326, P2_R1233_U137, P2_R1233_U324);
  or ginst14401 (P2_R1233_U327, P2_U3080, P2_U3432);
  not ginst14402 (P2_R1233_U328, P2_R1233_U161);
  or ginst14403 (P2_R1233_U329, P2_U3083, P2_U3485);
  not ginst14404 (P2_R1233_U33, P2_U3066);
  or ginst14405 (P2_R1233_U330, P2_U3075, P2_U3477);
  nand ginst14406 (P2_R1233_U331, P2_R1233_U330, P2_R1233_U92);
  nand ginst14407 (P2_R1233_U332, P2_R1233_U138, P2_R1233_U331);
  nand ginst14408 (P2_R1233_U333, P2_R1233_U262, P2_R1233_U59);
  nand ginst14409 (P2_R1233_U334, P2_U3071, P2_U3480);
  nand ginst14410 (P2_R1233_U335, P2_R1233_U139, P2_R1233_U333);
  or ginst14411 (P2_R1233_U336, P2_U3075, P2_U3477);
  nand ginst14412 (P2_R1233_U337, P2_R1233_U167, P2_R1233_U250);
  not ginst14413 (P2_R1233_U338, P2_R1233_U93);
  or ginst14414 (P2_R1233_U339, P2_U3074, P2_U3465);
  nand ginst14415 (P2_R1233_U34, P2_U3062, P2_U3441);
  nand ginst14416 (P2_R1233_U340, P2_R1233_U339, P2_R1233_U93);
  nand ginst14417 (P2_R1233_U341, P2_R1233_U140, P2_R1233_U340);
  nand ginst14418 (P2_R1233_U342, P2_R1233_U172, P2_R1233_U338);
  nand ginst14419 (P2_R1233_U343, P2_U3082, P2_U3468);
  nand ginst14420 (P2_R1233_U344, P2_R1233_U141, P2_R1233_U342);
  or ginst14421 (P2_R1233_U345, P2_U3074, P2_U3465);
  or ginst14422 (P2_R1233_U346, P2_U3085, P2_U3456);
  nand ginst14423 (P2_R1233_U347, P2_R1233_U346, P2_R1233_U40);
  nand ginst14424 (P2_R1233_U348, P2_R1233_U142, P2_R1233_U347);
  nand ginst14425 (P2_R1233_U349, P2_R1233_U171, P2_R1233_U206);
  not ginst14426 (P2_R1233_U35, P2_U3444);
  nand ginst14427 (P2_R1233_U350, P2_U3064, P2_U3459);
  nand ginst14428 (P2_R1233_U351, P2_R1233_U143, P2_R1233_U349);
  nand ginst14429 (P2_R1233_U352, P2_R1233_U171, P2_R1233_U207);
  nand ginst14430 (P2_R1233_U353, P2_R1233_U204, P2_R1233_U61);
  nand ginst14431 (P2_R1233_U354, P2_R1233_U214, P2_R1233_U22);
  nand ginst14432 (P2_R1233_U355, P2_R1233_U228, P2_R1233_U34);
  nand ginst14433 (P2_R1233_U356, P2_R1233_U180, P2_R1233_U231);
  nand ginst14434 (P2_R1233_U357, P2_R1233_U173, P2_R1233_U314);
  nand ginst14435 (P2_R1233_U358, P2_R1233_U176, P2_R1233_U298);
  nand ginst14436 (P2_R1233_U359, P2_R1233_U329, P2_R1233_U80);
  not ginst14437 (P2_R1233_U36, P2_U3453);
  nand ginst14438 (P2_R1233_U360, P2_R1233_U282, P2_R1233_U77);
  nand ginst14439 (P2_R1233_U361, P2_R1233_U336, P2_R1233_U59);
  nand ginst14440 (P2_R1233_U362, P2_R1233_U172, P2_R1233_U345);
  nand ginst14441 (P2_R1233_U363, P2_R1233_U250, P2_R1233_U68);
  nand ginst14442 (P2_R1233_U364, P2_U3056, P2_U3949);
  nand ginst14443 (P2_R1233_U365, P2_R1233_U168, P2_R1233_U296);
  nand ginst14444 (P2_R1233_U366, P2_R1233_U295, P2_U3059);
  nand ginst14445 (P2_R1233_U367, P2_R1233_U295, P2_U3951);
  nand ginst14446 (P2_R1233_U368, P2_R1233_U168, P2_R1233_U296, P2_R1233_U301);
  nand ginst14447 (P2_R1233_U369, P2_R1233_U133, P2_R1233_U155, P2_R1233_U168);
  not ginst14448 (P2_R1233_U37, P2_U3086);
  nand ginst14449 (P2_R1233_U370, P2_R1233_U297, P2_R1233_U301);
  nand ginst14450 (P2_R1233_U371, P2_R1233_U39, P2_U3085);
  nand ginst14451 (P2_R1233_U372, P2_R1233_U38, P2_U3456);
  nand ginst14452 (P2_R1233_U373, P2_R1233_U371, P2_R1233_U372);
  nand ginst14453 (P2_R1233_U374, P2_R1233_U352, P2_R1233_U40);
  nand ginst14454 (P2_R1233_U375, P2_R1233_U206, P2_R1233_U373);
  nand ginst14455 (P2_R1233_U376, P2_R1233_U36, P2_U3086);
  nand ginst14456 (P2_R1233_U377, P2_R1233_U37, P2_U3453);
  nand ginst14457 (P2_R1233_U378, P2_R1233_U376, P2_R1233_U377);
  nand ginst14458 (P2_R1233_U379, P2_R1233_U144, P2_R1233_U353);
  not ginst14459 (P2_R1233_U38, P2_U3085);
  nand ginst14460 (P2_R1233_U380, P2_R1233_U203, P2_R1233_U378);
  nand ginst14461 (P2_R1233_U381, P2_R1233_U23, P2_U3072);
  nand ginst14462 (P2_R1233_U382, P2_R1233_U21, P2_U3450);
  nand ginst14463 (P2_R1233_U383, P2_R1233_U19, P2_U3073);
  nand ginst14464 (P2_R1233_U384, P2_R1233_U20, P2_U3447);
  nand ginst14465 (P2_R1233_U385, P2_R1233_U383, P2_R1233_U384);
  nand ginst14466 (P2_R1233_U386, P2_R1233_U354, P2_R1233_U41);
  nand ginst14467 (P2_R1233_U387, P2_R1233_U195, P2_R1233_U385);
  nand ginst14468 (P2_R1233_U388, P2_R1233_U35, P2_U3069);
  nand ginst14469 (P2_R1233_U389, P2_R1233_U26, P2_U3444);
  not ginst14470 (P2_R1233_U39, P2_U3456);
  nand ginst14471 (P2_R1233_U390, P2_R1233_U24, P2_U3062);
  nand ginst14472 (P2_R1233_U391, P2_R1233_U25, P2_U3441);
  nand ginst14473 (P2_R1233_U392, P2_R1233_U390, P2_R1233_U391);
  nand ginst14474 (P2_R1233_U393, P2_R1233_U355, P2_R1233_U44);
  nand ginst14475 (P2_R1233_U394, P2_R1233_U221, P2_R1233_U392);
  nand ginst14476 (P2_R1233_U395, P2_R1233_U32, P2_U3066);
  nand ginst14477 (P2_R1233_U396, P2_R1233_U33, P2_U3438);
  nand ginst14478 (P2_R1233_U397, P2_R1233_U395, P2_R1233_U396);
  nand ginst14479 (P2_R1233_U398, P2_R1233_U145, P2_R1233_U356);
  nand ginst14480 (P2_R1233_U399, P2_R1233_U230, P2_R1233_U397);
  and ginst14481 (P2_R1233_U4, P2_R1233_U178, P2_R1233_U179);
  nand ginst14482 (P2_R1233_U40, P2_R1233_U205, P2_R1233_U61);
  nand ginst14483 (P2_R1233_U400, P2_R1233_U27, P2_U3070);
  nand ginst14484 (P2_R1233_U401, P2_R1233_U28, P2_U3435);
  nand ginst14485 (P2_R1233_U402, P2_R1233_U147, P2_U3057);
  nand ginst14486 (P2_R1233_U403, P2_R1233_U146, P2_U3960);
  nand ginst14487 (P2_R1233_U404, P2_R1233_U147, P2_U3057);
  nand ginst14488 (P2_R1233_U405, P2_R1233_U146, P2_U3960);
  nand ginst14489 (P2_R1233_U406, P2_R1233_U404, P2_R1233_U405);
  nand ginst14490 (P2_R1233_U407, P2_R1233_U148, P2_R1233_U149);
  nand ginst14491 (P2_R1233_U408, P2_R1233_U305, P2_R1233_U406);
  nand ginst14492 (P2_R1233_U409, P2_R1233_U88, P2_U3056);
  nand ginst14493 (P2_R1233_U41, P2_R1233_U117, P2_R1233_U193);
  nand ginst14494 (P2_R1233_U410, P2_R1233_U87, P2_U3949);
  nand ginst14495 (P2_R1233_U411, P2_R1233_U88, P2_U3056);
  nand ginst14496 (P2_R1233_U412, P2_R1233_U87, P2_U3949);
  nand ginst14497 (P2_R1233_U413, P2_R1233_U411, P2_R1233_U412);
  nand ginst14498 (P2_R1233_U414, P2_R1233_U150, P2_R1233_U151);
  nand ginst14499 (P2_R1233_U415, P2_R1233_U303, P2_R1233_U413);
  nand ginst14500 (P2_R1233_U416, P2_R1233_U46, P2_U3055);
  nand ginst14501 (P2_R1233_U417, P2_R1233_U47, P2_U3950);
  nand ginst14502 (P2_R1233_U418, P2_R1233_U46, P2_U3055);
  nand ginst14503 (P2_R1233_U419, P2_R1233_U47, P2_U3950);
  nand ginst14504 (P2_R1233_U42, P2_R1233_U182, P2_R1233_U183);
  nand ginst14505 (P2_R1233_U420, P2_R1233_U418, P2_R1233_U419);
  nand ginst14506 (P2_R1233_U421, P2_R1233_U152, P2_R1233_U153);
  nand ginst14507 (P2_R1233_U422, P2_R1233_U300, P2_R1233_U420);
  nand ginst14508 (P2_R1233_U423, P2_R1233_U49, P2_U3059);
  nand ginst14509 (P2_R1233_U424, P2_R1233_U48, P2_U3951);
  nand ginst14510 (P2_R1233_U425, P2_R1233_U50, P2_U3060);
  nand ginst14511 (P2_R1233_U426, P2_R1233_U51, P2_U3952);
  nand ginst14512 (P2_R1233_U427, P2_R1233_U425, P2_R1233_U426);
  nand ginst14513 (P2_R1233_U428, P2_R1233_U357, P2_R1233_U89);
  nand ginst14514 (P2_R1233_U429, P2_R1233_U307, P2_R1233_U427);
  nand ginst14515 (P2_R1233_U43, P2_U3080, P2_U3432);
  nand ginst14516 (P2_R1233_U430, P2_R1233_U52, P2_U3067);
  nand ginst14517 (P2_R1233_U431, P2_R1233_U53, P2_U3953);
  nand ginst14518 (P2_R1233_U432, P2_R1233_U430, P2_R1233_U431);
  nand ginst14519 (P2_R1233_U433, P2_R1233_U155, P2_R1233_U358);
  nand ginst14520 (P2_R1233_U434, P2_R1233_U294, P2_R1233_U432);
  nand ginst14521 (P2_R1233_U435, P2_R1233_U84, P2_U3068);
  nand ginst14522 (P2_R1233_U436, P2_R1233_U85, P2_U3954);
  nand ginst14523 (P2_R1233_U437, P2_R1233_U84, P2_U3068);
  nand ginst14524 (P2_R1233_U438, P2_R1233_U85, P2_U3954);
  nand ginst14525 (P2_R1233_U439, P2_R1233_U437, P2_R1233_U438);
  nand ginst14526 (P2_R1233_U44, P2_R1233_U122, P2_R1233_U219);
  nand ginst14527 (P2_R1233_U440, P2_R1233_U156, P2_R1233_U157);
  nand ginst14528 (P2_R1233_U441, P2_R1233_U290, P2_R1233_U439);
  nand ginst14529 (P2_R1233_U442, P2_R1233_U82, P2_U3063);
  nand ginst14530 (P2_R1233_U443, P2_R1233_U83, P2_U3955);
  nand ginst14531 (P2_R1233_U444, P2_R1233_U82, P2_U3063);
  nand ginst14532 (P2_R1233_U445, P2_R1233_U83, P2_U3955);
  nand ginst14533 (P2_R1233_U446, P2_R1233_U444, P2_R1233_U445);
  nand ginst14534 (P2_R1233_U447, P2_R1233_U158, P2_R1233_U159);
  nand ginst14535 (P2_R1233_U448, P2_R1233_U286, P2_R1233_U446);
  nand ginst14536 (P2_R1233_U449, P2_R1233_U54, P2_U3077);
  nand ginst14537 (P2_R1233_U45, P2_R1233_U215, P2_R1233_U216);
  nand ginst14538 (P2_R1233_U450, P2_R1233_U55, P2_U3956);
  nand ginst14539 (P2_R1233_U451, P2_R1233_U54, P2_U3077);
  nand ginst14540 (P2_R1233_U452, P2_R1233_U55, P2_U3956);
  nand ginst14541 (P2_R1233_U453, P2_R1233_U451, P2_R1233_U452);
  nand ginst14542 (P2_R1233_U454, P2_R1233_U81, P2_U3078);
  nand ginst14543 (P2_R1233_U455, P2_R1233_U90, P2_U3957);
  nand ginst14544 (P2_R1233_U456, P2_R1233_U161, P2_R1233_U182);
  nand ginst14545 (P2_R1233_U457, P2_R1233_U31, P2_R1233_U328);
  nand ginst14546 (P2_R1233_U458, P2_R1233_U78, P2_U3083);
  nand ginst14547 (P2_R1233_U459, P2_R1233_U79, P2_U3485);
  not ginst14548 (P2_R1233_U46, P2_U3950);
  nand ginst14549 (P2_R1233_U460, P2_R1233_U458, P2_R1233_U459);
  nand ginst14550 (P2_R1233_U461, P2_R1233_U359, P2_R1233_U91);
  nand ginst14551 (P2_R1233_U462, P2_R1233_U316, P2_R1233_U460);
  nand ginst14552 (P2_R1233_U463, P2_R1233_U75, P2_U3084);
  nand ginst14553 (P2_R1233_U464, P2_R1233_U76, P2_U3483);
  nand ginst14554 (P2_R1233_U465, P2_R1233_U463, P2_R1233_U464);
  nand ginst14555 (P2_R1233_U466, P2_R1233_U162, P2_R1233_U360);
  nand ginst14556 (P2_R1233_U467, P2_R1233_U270, P2_R1233_U465);
  nand ginst14557 (P2_R1233_U468, P2_R1233_U60, P2_U3071);
  nand ginst14558 (P2_R1233_U469, P2_R1233_U58, P2_U3480);
  not ginst14559 (P2_R1233_U47, P2_U3055);
  nand ginst14560 (P2_R1233_U470, P2_R1233_U56, P2_U3075);
  nand ginst14561 (P2_R1233_U471, P2_R1233_U57, P2_U3477);
  nand ginst14562 (P2_R1233_U472, P2_R1233_U470, P2_R1233_U471);
  nand ginst14563 (P2_R1233_U473, P2_R1233_U361, P2_R1233_U92);
  nand ginst14564 (P2_R1233_U474, P2_R1233_U262, P2_R1233_U472);
  nand ginst14565 (P2_R1233_U475, P2_R1233_U73, P2_U3076);
  nand ginst14566 (P2_R1233_U476, P2_R1233_U74, P2_U3474);
  nand ginst14567 (P2_R1233_U477, P2_R1233_U73, P2_U3076);
  nand ginst14568 (P2_R1233_U478, P2_R1233_U74, P2_U3474);
  nand ginst14569 (P2_R1233_U479, P2_R1233_U477, P2_R1233_U478);
  not ginst14570 (P2_R1233_U48, P2_U3059);
  nand ginst14571 (P2_R1233_U480, P2_R1233_U163, P2_R1233_U164);
  nand ginst14572 (P2_R1233_U481, P2_R1233_U258, P2_R1233_U479);
  nand ginst14573 (P2_R1233_U482, P2_R1233_U71, P2_U3081);
  nand ginst14574 (P2_R1233_U483, P2_R1233_U72, P2_U3471);
  nand ginst14575 (P2_R1233_U484, P2_R1233_U71, P2_U3081);
  nand ginst14576 (P2_R1233_U485, P2_R1233_U72, P2_U3471);
  nand ginst14577 (P2_R1233_U486, P2_R1233_U484, P2_R1233_U485);
  nand ginst14578 (P2_R1233_U487, P2_R1233_U165, P2_R1233_U166);
  nand ginst14579 (P2_R1233_U488, P2_R1233_U254, P2_R1233_U486);
  nand ginst14580 (P2_R1233_U489, P2_R1233_U69, P2_U3082);
  not ginst14581 (P2_R1233_U49, P2_U3951);
  nand ginst14582 (P2_R1233_U490, P2_R1233_U70, P2_U3468);
  nand ginst14583 (P2_R1233_U491, P2_R1233_U64, P2_U3074);
  nand ginst14584 (P2_R1233_U492, P2_R1233_U65, P2_U3465);
  nand ginst14585 (P2_R1233_U493, P2_R1233_U491, P2_R1233_U492);
  nand ginst14586 (P2_R1233_U494, P2_R1233_U362, P2_R1233_U93);
  nand ginst14587 (P2_R1233_U495, P2_R1233_U338, P2_R1233_U493);
  nand ginst14588 (P2_R1233_U496, P2_R1233_U66, P2_U3065);
  nand ginst14589 (P2_R1233_U497, P2_R1233_U67, P2_U3462);
  nand ginst14590 (P2_R1233_U498, P2_R1233_U496, P2_R1233_U497);
  nand ginst14591 (P2_R1233_U499, P2_R1233_U167, P2_R1233_U363);
  and ginst14592 (P2_R1233_U5, P2_R1233_U196, P2_R1233_U197);
  not ginst14593 (P2_R1233_U50, P2_U3952);
  nand ginst14594 (P2_R1233_U500, P2_R1233_U244, P2_R1233_U498);
  nand ginst14595 (P2_R1233_U501, P2_R1233_U62, P2_U3064);
  nand ginst14596 (P2_R1233_U502, P2_R1233_U63, P2_U3459);
  nand ginst14597 (P2_R1233_U503, P2_R1233_U29, P2_U3079);
  nand ginst14598 (P2_R1233_U504, P2_R1233_U30, P2_U3427);
  not ginst14599 (P2_R1233_U51, P2_U3060);
  not ginst14600 (P2_R1233_U52, P2_U3953);
  not ginst14601 (P2_R1233_U53, P2_U3067);
  not ginst14602 (P2_R1233_U54, P2_U3956);
  not ginst14603 (P2_R1233_U55, P2_U3077);
  not ginst14604 (P2_R1233_U56, P2_U3477);
  not ginst14605 (P2_R1233_U57, P2_U3075);
  not ginst14606 (P2_R1233_U58, P2_U3071);
  nand ginst14607 (P2_R1233_U59, P2_U3075, P2_U3477);
  and ginst14608 (P2_R1233_U6, P2_R1233_U236, P2_R1233_U237);
  not ginst14609 (P2_R1233_U60, P2_U3480);
  nand ginst14610 (P2_R1233_U61, P2_U3086, P2_U3453);
  not ginst14611 (P2_R1233_U62, P2_U3459);
  not ginst14612 (P2_R1233_U63, P2_U3064);
  not ginst14613 (P2_R1233_U64, P2_U3465);
  not ginst14614 (P2_R1233_U65, P2_U3074);
  not ginst14615 (P2_R1233_U66, P2_U3462);
  not ginst14616 (P2_R1233_U67, P2_U3065);
  nand ginst14617 (P2_R1233_U68, P2_U3065, P2_U3462);
  not ginst14618 (P2_R1233_U69, P2_U3468);
  and ginst14619 (P2_R1233_U7, P2_R1233_U245, P2_R1233_U246);
  not ginst14620 (P2_R1233_U70, P2_U3082);
  not ginst14621 (P2_R1233_U71, P2_U3471);
  not ginst14622 (P2_R1233_U72, P2_U3081);
  not ginst14623 (P2_R1233_U73, P2_U3474);
  not ginst14624 (P2_R1233_U74, P2_U3076);
  not ginst14625 (P2_R1233_U75, P2_U3483);
  not ginst14626 (P2_R1233_U76, P2_U3084);
  nand ginst14627 (P2_R1233_U77, P2_U3084, P2_U3483);
  not ginst14628 (P2_R1233_U78, P2_U3485);
  not ginst14629 (P2_R1233_U79, P2_U3083);
  and ginst14630 (P2_R1233_U8, P2_R1233_U263, P2_R1233_U264);
  nand ginst14631 (P2_R1233_U80, P2_U3083, P2_U3485);
  not ginst14632 (P2_R1233_U81, P2_U3957);
  not ginst14633 (P2_R1233_U82, P2_U3955);
  not ginst14634 (P2_R1233_U83, P2_U3063);
  not ginst14635 (P2_R1233_U84, P2_U3954);
  not ginst14636 (P2_R1233_U85, P2_U3068);
  nand ginst14637 (P2_R1233_U86, P2_U3059, P2_U3951);
  not ginst14638 (P2_R1233_U87, P2_U3056);
  not ginst14639 (P2_R1233_U88, P2_U3949);
  nand ginst14640 (P2_R1233_U89, P2_R1233_U176, P2_R1233_U306);
  and ginst14641 (P2_R1233_U9, P2_R1233_U271, P2_R1233_U272);
  not ginst14642 (P2_R1233_U90, P2_U3078);
  nand ginst14643 (P2_R1233_U91, P2_R1233_U315, P2_R1233_U77);
  nand ginst14644 (P2_R1233_U92, P2_R1233_U260, P2_R1233_U261);
  nand ginst14645 (P2_R1233_U93, P2_R1233_U337, P2_R1233_U68);
  nand ginst14646 (P2_R1233_U94, P2_R1233_U456, P2_R1233_U457);
  nand ginst14647 (P2_R1233_U95, P2_R1233_U503, P2_R1233_U504);
  nand ginst14648 (P2_R1233_U96, P2_R1233_U374, P2_R1233_U375);
  nand ginst14649 (P2_R1233_U97, P2_R1233_U379, P2_R1233_U380);
  nand ginst14650 (P2_R1233_U98, P2_R1233_U386, P2_R1233_U387);
  nand ginst14651 (P2_R1233_U99, P2_R1233_U393, P2_R1233_U394);
  and ginst14652 (P2_R1275_U10, P2_R1275_U129, P2_R1275_U39);
  not ginst14653 (P2_R1275_U100, P2_R1275_U36);
  not ginst14654 (P2_R1275_U101, P2_R1275_U37);
  not ginst14655 (P2_R1275_U102, P2_R1275_U38);
  not ginst14656 (P2_R1275_U103, P2_R1275_U39);
  not ginst14657 (P2_R1275_U104, P2_R1275_U40);
  not ginst14658 (P2_R1275_U105, P2_R1275_U41);
  not ginst14659 (P2_R1275_U106, P2_R1275_U42);
  not ginst14660 (P2_R1275_U107, P2_R1275_U43);
  not ginst14661 (P2_R1275_U108, P2_R1275_U44);
  not ginst14662 (P2_R1275_U109, P2_R1275_U45);
  and ginst14663 (P2_R1275_U11, P2_R1275_U128, P2_R1275_U40);
  not ginst14664 (P2_R1275_U110, P2_R1275_U46);
  not ginst14665 (P2_R1275_U111, P2_R1275_U67);
  nand ginst14666 (P2_R1275_U112, P2_R1275_U110, P2_R1275_U69);
  nand ginst14667 (P2_R1275_U113, P2_R1275_U112, P2_U3959);
  or ginst14668 (P2_R1275_U114, P2_U3427, P2_U3432);
  nand ginst14669 (P2_R1275_U115, P2_R1275_U114, P2_U3435);
  nand ginst14670 (P2_R1275_U116, P2_R1275_U109, P2_R1275_U71);
  nand ginst14671 (P2_R1275_U117, P2_R1275_U116, P2_U3949);
  nand ginst14672 (P2_R1275_U118, P2_R1275_U108, P2_R1275_U73);
  nand ginst14673 (P2_R1275_U119, P2_R1275_U118, P2_U3951);
  and ginst14674 (P2_R1275_U12, P2_R1275_U127, P2_R1275_U41);
  nand ginst14675 (P2_R1275_U120, P2_R1275_U107, P2_R1275_U75);
  nand ginst14676 (P2_R1275_U121, P2_R1275_U120, P2_U3953);
  nand ginst14677 (P2_R1275_U122, P2_R1275_U106, P2_R1275_U77);
  nand ginst14678 (P2_R1275_U123, P2_R1275_U122, P2_U3955);
  nand ginst14679 (P2_R1275_U124, P2_R1275_U105, P2_R1275_U81);
  nand ginst14680 (P2_R1275_U125, P2_R1275_U124, P2_U3957);
  nand ginst14681 (P2_R1275_U126, P2_R1275_U104, P2_R1275_U83);
  nand ginst14682 (P2_R1275_U127, P2_R1275_U126, P2_U3483);
  nand ginst14683 (P2_R1275_U128, P2_R1275_U39, P2_U3477);
  nand ginst14684 (P2_R1275_U129, P2_R1275_U38, P2_U3474);
  and ginst14685 (P2_R1275_U13, P2_R1275_U125, P2_R1275_U42);
  nand ginst14686 (P2_R1275_U130, P2_R1275_U101, P2_R1275_U85);
  nand ginst14687 (P2_R1275_U131, P2_R1275_U130, P2_U3471);
  nand ginst14688 (P2_R1275_U132, P2_R1275_U36, P2_U3465);
  nand ginst14689 (P2_R1275_U133, P2_R1275_U35, P2_U3462);
  nand ginst14690 (P2_R1275_U134, P2_R1275_U62, P2_R1275_U92);
  nand ginst14691 (P2_R1275_U135, P2_R1275_U134, P2_U3459);
  nand ginst14692 (P2_R1275_U136, P2_R1275_U30, P2_U3456);
  nand ginst14693 (P2_R1275_U137, P2_R1275_U62, P2_R1275_U92);
  nand ginst14694 (P2_R1275_U138, P2_R1275_U27, P2_U3444);
  nand ginst14695 (P2_R1275_U139, P2_R1275_U64, P2_R1275_U89);
  and ginst14696 (P2_R1275_U14, P2_R1275_U123, P2_R1275_U43);
  nand ginst14697 (P2_R1275_U140, P2_R1275_U67, P2_U3958);
  nand ginst14698 (P2_R1275_U141, P2_R1275_U111, P2_R1275_U66);
  nand ginst14699 (P2_R1275_U142, P2_R1275_U46, P2_U3960);
  nand ginst14700 (P2_R1275_U143, P2_R1275_U110, P2_R1275_U69);
  nand ginst14701 (P2_R1275_U144, P2_R1275_U45, P2_U3950);
  nand ginst14702 (P2_R1275_U145, P2_R1275_U109, P2_R1275_U71);
  nand ginst14703 (P2_R1275_U146, P2_R1275_U44, P2_U3952);
  nand ginst14704 (P2_R1275_U147, P2_R1275_U108, P2_R1275_U73);
  nand ginst14705 (P2_R1275_U148, P2_R1275_U43, P2_U3954);
  nand ginst14706 (P2_R1275_U149, P2_R1275_U107, P2_R1275_U75);
  and ginst14707 (P2_R1275_U15, P2_R1275_U121, P2_R1275_U44);
  nand ginst14708 (P2_R1275_U150, P2_R1275_U42, P2_U3956);
  nand ginst14709 (P2_R1275_U151, P2_R1275_U106, P2_R1275_U77);
  nand ginst14710 (P2_R1275_U152, P2_R1275_U80, P2_U3432);
  nand ginst14711 (P2_R1275_U153, P2_R1275_U79, P2_U3427);
  nand ginst14712 (P2_R1275_U154, P2_R1275_U41, P2_U3485);
  nand ginst14713 (P2_R1275_U155, P2_R1275_U105, P2_R1275_U81);
  nand ginst14714 (P2_R1275_U156, P2_R1275_U40, P2_U3480);
  nand ginst14715 (P2_R1275_U157, P2_R1275_U104, P2_R1275_U83);
  nand ginst14716 (P2_R1275_U158, P2_R1275_U37, P2_U3468);
  nand ginst14717 (P2_R1275_U159, P2_R1275_U101, P2_R1275_U85);
  and ginst14718 (P2_R1275_U16, P2_R1275_U119, P2_R1275_U45);
  and ginst14719 (P2_R1275_U17, P2_R1275_U117, P2_R1275_U46);
  and ginst14720 (P2_R1275_U18, P2_R1275_U115, P2_R1275_U25);
  and ginst14721 (P2_R1275_U19, P2_R1275_U113, P2_R1275_U67);
  and ginst14722 (P2_R1275_U20, P2_R1275_U26, P2_R1275_U98);
  and ginst14723 (P2_R1275_U21, P2_R1275_U27, P2_R1275_U97);
  and ginst14724 (P2_R1275_U22, P2_R1275_U28, P2_R1275_U96);
  and ginst14725 (P2_R1275_U23, P2_R1275_U29, P2_R1275_U94);
  and ginst14726 (P2_R1275_U24, P2_R1275_U30, P2_R1275_U93);
  or ginst14727 (P2_R1275_U25, P2_U3427, P2_U3432, P2_U3435);
  nand ginst14728 (P2_R1275_U26, P2_R1275_U34, P2_R1275_U87);
  nand ginst14729 (P2_R1275_U27, P2_R1275_U33, P2_R1275_U88);
  nand ginst14730 (P2_R1275_U28, P2_R1275_U56, P2_R1275_U89);
  nand ginst14731 (P2_R1275_U29, P2_R1275_U32, P2_R1275_U90);
  nand ginst14732 (P2_R1275_U30, P2_R1275_U31, P2_R1275_U91);
  not ginst14733 (P2_R1275_U31, P2_U3453);
  not ginst14734 (P2_R1275_U32, P2_U3450);
  not ginst14735 (P2_R1275_U33, P2_U3441);
  not ginst14736 (P2_R1275_U34, P2_U3438);
  nand ginst14737 (P2_R1275_U35, P2_R1275_U57, P2_R1275_U92);
  nand ginst14738 (P2_R1275_U36, P2_R1275_U54, P2_R1275_U99);
  nand ginst14739 (P2_R1275_U37, P2_R1275_U100, P2_R1275_U53);
  nand ginst14740 (P2_R1275_U38, P2_R1275_U101, P2_R1275_U58);
  nand ginst14741 (P2_R1275_U39, P2_R1275_U102, P2_R1275_U52);
  nand ginst14742 (P2_R1275_U40, P2_R1275_U103, P2_R1275_U51);
  nand ginst14743 (P2_R1275_U41, P2_R1275_U104, P2_R1275_U59);
  nand ginst14744 (P2_R1275_U42, P2_R1275_U105, P2_R1275_U60);
  nand ginst14745 (P2_R1275_U43, P2_R1275_U106, P2_R1275_U61);
  nand ginst14746 (P2_R1275_U44, P2_R1275_U107, P2_R1275_U50, P2_R1275_U75);
  nand ginst14747 (P2_R1275_U45, P2_R1275_U108, P2_R1275_U49, P2_R1275_U73);
  nand ginst14748 (P2_R1275_U46, P2_R1275_U109, P2_R1275_U48, P2_R1275_U71);
  not ginst14749 (P2_R1275_U47, P2_U3959);
  not ginst14750 (P2_R1275_U48, P2_U3949);
  not ginst14751 (P2_R1275_U49, P2_U3951);
  not ginst14752 (P2_R1275_U50, P2_U3953);
  not ginst14753 (P2_R1275_U51, P2_U3477);
  not ginst14754 (P2_R1275_U52, P2_U3474);
  not ginst14755 (P2_R1275_U53, P2_U3465);
  not ginst14756 (P2_R1275_U54, P2_U3462);
  nand ginst14757 (P2_R1275_U55, P2_R1275_U152, P2_R1275_U153);
  nor ginst14758 (P2_R1275_U56, P2_U3444, P2_U3447);
  nor ginst14759 (P2_R1275_U57, P2_U3456, P2_U3459);
  nor ginst14760 (P2_R1275_U58, P2_U3468, P2_U3471);
  nor ginst14761 (P2_R1275_U59, P2_U3480, P2_U3483);
  and ginst14762 (P2_R1275_U6, P2_R1275_U135, P2_R1275_U35);
  nor ginst14763 (P2_R1275_U60, P2_U3485, P2_U3957);
  nor ginst14764 (P2_R1275_U61, P2_U3955, P2_U3956);
  not ginst14765 (P2_R1275_U62, P2_U3456);
  and ginst14766 (P2_R1275_U63, P2_R1275_U136, P2_R1275_U137);
  not ginst14767 (P2_R1275_U64, P2_U3444);
  and ginst14768 (P2_R1275_U65, P2_R1275_U138, P2_R1275_U139);
  not ginst14769 (P2_R1275_U66, P2_U3958);
  nand ginst14770 (P2_R1275_U67, P2_R1275_U110, P2_R1275_U47, P2_R1275_U69);
  and ginst14771 (P2_R1275_U68, P2_R1275_U140, P2_R1275_U141);
  not ginst14772 (P2_R1275_U69, P2_U3960);
  and ginst14773 (P2_R1275_U7, P2_R1275_U133, P2_R1275_U36);
  and ginst14774 (P2_R1275_U70, P2_R1275_U142, P2_R1275_U143);
  not ginst14775 (P2_R1275_U71, P2_U3950);
  and ginst14776 (P2_R1275_U72, P2_R1275_U144, P2_R1275_U145);
  not ginst14777 (P2_R1275_U73, P2_U3952);
  and ginst14778 (P2_R1275_U74, P2_R1275_U146, P2_R1275_U147);
  not ginst14779 (P2_R1275_U75, P2_U3954);
  and ginst14780 (P2_R1275_U76, P2_R1275_U148, P2_R1275_U149);
  not ginst14781 (P2_R1275_U77, P2_U3956);
  and ginst14782 (P2_R1275_U78, P2_R1275_U150, P2_R1275_U151);
  not ginst14783 (P2_R1275_U79, P2_U3432);
  and ginst14784 (P2_R1275_U8, P2_R1275_U132, P2_R1275_U37);
  not ginst14785 (P2_R1275_U80, P2_U3427);
  not ginst14786 (P2_R1275_U81, P2_U3485);
  and ginst14787 (P2_R1275_U82, P2_R1275_U154, P2_R1275_U155);
  not ginst14788 (P2_R1275_U83, P2_U3480);
  and ginst14789 (P2_R1275_U84, P2_R1275_U156, P2_R1275_U157);
  not ginst14790 (P2_R1275_U85, P2_U3468);
  and ginst14791 (P2_R1275_U86, P2_R1275_U158, P2_R1275_U159);
  not ginst14792 (P2_R1275_U87, P2_R1275_U25);
  not ginst14793 (P2_R1275_U88, P2_R1275_U26);
  not ginst14794 (P2_R1275_U89, P2_R1275_U27);
  and ginst14795 (P2_R1275_U9, P2_R1275_U131, P2_R1275_U38);
  not ginst14796 (P2_R1275_U90, P2_R1275_U28);
  not ginst14797 (P2_R1275_U91, P2_R1275_U29);
  not ginst14798 (P2_R1275_U92, P2_R1275_U30);
  nand ginst14799 (P2_R1275_U93, P2_R1275_U29, P2_U3453);
  nand ginst14800 (P2_R1275_U94, P2_R1275_U28, P2_U3450);
  nand ginst14801 (P2_R1275_U95, P2_R1275_U64, P2_R1275_U89);
  nand ginst14802 (P2_R1275_U96, P2_R1275_U95, P2_U3447);
  nand ginst14803 (P2_R1275_U97, P2_R1275_U26, P2_U3441);
  nand ginst14804 (P2_R1275_U98, P2_R1275_U25, P2_U3438);
  not ginst14805 (P2_R1275_U99, P2_R1275_U35);
  and ginst14806 (P2_R1299_U6, P2_R1299_U7, P2_U3061);
  not ginst14807 (P2_R1299_U7, P2_U3058);
  and ginst14808 (P2_R1312_U10, P2_R1312_U212, P2_R1312_U213);
  and ginst14809 (P2_R1312_U100, P2_R1312_U13, P2_U3141);
  and ginst14810 (P2_R1312_U101, P2_R1312_U167, P2_R1312_U168, P2_R1312_U177, P2_R1312_U33);
  and ginst14811 (P2_R1312_U102, P2_R1312_U103, P2_R1312_U13);
  and ginst14812 (P2_R1312_U103, P2_R1312_U178, P2_U3143);
  and ginst14813 (P2_R1312_U104, P2_R1312_U166, P2_R1312_U167, P2_R1312_U168, P2_R1312_U49);
  and ginst14814 (P2_R1312_U105, P2_R1312_U164, P2_R1312_U166, P2_R1312_U167, P2_R1312_U168, P2_R1312_U47);
  and ginst14815 (P2_R1312_U106, P2_R1312_U167, P2_R1312_U168, P2_R1312_U169, P2_R1312_U45);
  and ginst14816 (P2_R1312_U107, P2_R1312_U16, P2_U3131);
  and ginst14817 (P2_R1312_U108, P2_R1312_U167, P2_R1312_U168, P2_R1312_U171, P2_R1312_U41);
  and ginst14818 (P2_R1312_U109, P2_R1312_U16, P2_U3134);
  and ginst14819 (P2_R1312_U11, P2_R1312_U14, P2_R1312_U169, P2_R1312_U82);
  and ginst14820 (P2_R1312_U110, P2_R1312_U167, P2_R1312_U168, P2_R1312_U170, P2_R1312_U43);
  and ginst14821 (P2_R1312_U111, P2_R1312_U11, P2_R1312_U112, P2_R1312_U166, P2_R1312_U17, P2_R1312_U171);
  and ginst14822 (P2_R1312_U112, P2_R1312_U16, P2_U3135);
  and ginst14823 (P2_R1312_U113, P2_R1312_U166, P2_R1312_U167, P2_R1312_U27);
  and ginst14824 (P2_R1312_U114, P2_R1312_U168, P2_U3137);
  and ginst14825 (P2_R1312_U115, P2_R1312_U157, P2_R1312_U166, P2_R1312_U167, P2_R1312_U37);
  and ginst14826 (P2_R1312_U116, P2_R1312_U156, P2_R1312_U157, P2_R1312_U166, P2_R1312_U167, P2_R1312_U35);
  and ginst14827 (P2_R1312_U117, P2_R1312_U166, P2_R1312_U167, P2_R1312_U168, P2_R1312_U42);
  and ginst14828 (P2_R1312_U118, P2_R1312_U16, P2_U3133);
  and ginst14829 (P2_R1312_U119, P2_R1312_U166, P2_R1312_U167, P2_R1312_U168, P2_R1312_U30);
  and ginst14830 (P2_R1312_U12, P2_R1312_U154, P2_R1312_U155, P2_R1312_U156, P2_R1312_U157);
  and ginst14831 (P2_R1312_U120, P2_R1312_U173, P2_R1312_U174, P2_U3139);
  and ginst14832 (P2_R1312_U121, P2_R1312_U166, P2_R1312_U167, P2_R1312_U168, P2_R1312_U38);
  and ginst14833 (P2_R1312_U122, P2_R1312_U161, P2_R1312_U164, P2_R1312_U166, P2_R1312_U167, P2_R1312_U48);
  and ginst14834 (P2_R1312_U123, P2_R1312_U168, P2_R1312_U169);
  and ginst14835 (P2_R1312_U124, P2_R1312_U160, P2_R1312_U166, P2_R1312_U167, P2_R1312_U168, P2_R1312_U44);
  and ginst14836 (P2_R1312_U125, P2_R1312_U16, P2_U3132);
  and ginst14837 (P2_R1312_U126, P2_R1312_U167, P2_R1312_U39);
  and ginst14838 (P2_R1312_U127, P2_R1312_U126, P2_R1312_U168, P2_R1312_U17);
  and ginst14839 (P2_R1312_U128, P2_R1312_U6, P2_U3136);
  and ginst14840 (P2_R1312_U129, P2_R1312_U166, P2_R1312_U167, P2_R1312_U168, P2_R1312_U28);
  and ginst14841 (P2_R1312_U13, P2_R1312_U173, P2_R1312_U174, P2_R1312_U175, P2_R1312_U176);
  and ginst14842 (P2_R1312_U130, P2_R1312_U173, P2_U3138);
  and ginst14843 (P2_R1312_U131, P2_R1312_U166, P2_R1312_U167, P2_R1312_U168, P2_R1312_U32);
  and ginst14844 (P2_R1312_U132, P2_R1312_U13, P2_R1312_U133);
  and ginst14845 (P2_R1312_U133, P2_R1312_U177, P2_U3142);
  and ginst14846 (P2_R1312_U134, P2_R1312_U167, P2_R1312_U168, P2_R1312_U177, P2_R1312_U34);
  and ginst14847 (P2_R1312_U135, P2_R1312_U13, P2_R1312_U136);
  and ginst14848 (P2_R1312_U136, P2_R1312_U178, P2_R1312_U179, P2_U3144);
  and ginst14849 (P2_R1312_U137, P2_R1312_U154, P2_R1312_U156, P2_R1312_U157, P2_R1312_U166, P2_R1312_U36);
  and ginst14850 (P2_R1312_U138, P2_R1312_U167, P2_R1312_U168, P2_R1312_U8, P2_U3148);
  and ginst14851 (P2_R1312_U139, P2_R1312_U167, P2_R1312_U168, P2_R1312_U221, P2_R1312_U52);
  and ginst14852 (P2_R1312_U14, P2_R1312_U161, P2_R1312_U162, P2_R1312_U164);
  and ginst14853 (P2_R1312_U140, P2_R1312_U12, P2_U3150);
  and ginst14854 (P2_R1312_U141, P2_R1312_U153, P2_R1312_U181);
  and ginst14855 (P2_R1312_U142, P2_R1312_U188, P2_R1312_U192);
  and ginst14856 (P2_R1312_U143, P2_R1312_U197, P2_R1312_U198, P2_R1312_U199);
  and ginst14857 (P2_R1312_U144, P2_R1312_U141, P2_R1312_U142, P2_R1312_U143);
  and ginst14858 (P2_R1312_U145, P2_R1312_U202, P2_R1312_U203);
  and ginst14859 (P2_R1312_U146, P2_R1312_U204, P2_R1312_U205);
  and ginst14860 (P2_R1312_U147, P2_R1312_U145, P2_R1312_U146, P2_R1312_U200, P2_R1312_U201, P2_R1312_U206);
  and ginst14861 (P2_R1312_U148, P2_R1312_U209, P2_R1312_U210);
  and ginst14862 (P2_R1312_U149, P2_R1312_U214, P2_R1312_U215);
  and ginst14863 (P2_R1312_U15, P2_R1312_U11, P2_R1312_U165, P2_R1312_U17, P2_R1312_U6, P2_R1312_U83);
  and ginst14864 (P2_R1312_U150, P2_R1312_U148, P2_R1312_U149, P2_R1312_U207, P2_R1312_U208, P2_R1312_U211);
  and ginst14865 (P2_R1312_U151, P2_R1312_U216, P2_R1312_U217, P2_R1312_U218, P2_R1312_U219);
  and ginst14866 (P2_R1312_U152, P2_R1312_U10, P2_R1312_U220, P2_R1312_U222);
  nand ginst14867 (P2_R1312_U153, P2_R1312_U191, P2_R1312_U81);
  nand ginst14868 (P2_R1312_U154, P2_R1312_U68, P2_U3115);
  nand ginst14869 (P2_R1312_U155, P2_R1312_U78, P2_U3116);
  nand ginst14870 (P2_R1312_U156, P2_R1312_U67, P2_U3114);
  nand ginst14871 (P2_R1312_U157, P2_R1312_U71, P2_U3113);
  nand ginst14872 (P2_R1312_U158, P2_R1312_U74, P2_U3104);
  nand ginst14873 (P2_R1312_U159, P2_R1312_U73, P2_U3100);
  and ginst14874 (P2_R1312_U16, P2_R1312_U163, P2_R1312_U165);
  nand ginst14875 (P2_R1312_U160, P2_R1312_U63, P2_U3099);
  nand ginst14876 (P2_R1312_U161, P2_R1312_U62, P2_U3097);
  nand ginst14877 (P2_R1312_U162, P2_R1312_U72, P2_U3098);
  nand ginst14878 (P2_R1312_U163, P2_R1312_U23, P2_U3094);
  nand ginst14879 (P2_R1312_U164, P2_R1312_U61, P2_U3096);
  nand ginst14880 (P2_R1312_U165, P2_R1312_U56, P2_U3093);
  nand ginst14881 (P2_R1312_U166, P2_R1312_U80, P2_U3090);
  nand ginst14882 (P2_R1312_U167, P2_R1312_U24, P2_U3091);
  nand ginst14883 (P2_R1312_U168, P2_R1312_U57, P2_U3092);
  nand ginst14884 (P2_R1312_U169, P2_R1312_U55, P2_U3095);
  and ginst14885 (P2_R1312_U17, P2_R1312_U224, P2_R1312_U225);
  nand ginst14886 (P2_R1312_U170, P2_R1312_U64, P2_U3102);
  nand ginst14887 (P2_R1312_U171, P2_R1312_U69, P2_U3101);
  nand ginst14888 (P2_R1312_U172, P2_R1312_U65, P2_U3103);
  nand ginst14889 (P2_R1312_U173, P2_R1312_U66, P2_U3105);
  nand ginst14890 (P2_R1312_U174, P2_R1312_U75, P2_U3106);
  nand ginst14891 (P2_R1312_U175, P2_R1312_U58, P2_U3108);
  nand ginst14892 (P2_R1312_U176, P2_R1312_U70, P2_U3107);
  nand ginst14893 (P2_R1312_U177, P2_R1312_U59, P2_U3109);
  nand ginst14894 (P2_R1312_U178, P2_R1312_U76, P2_U3110);
  nand ginst14895 (P2_R1312_U179, P2_R1312_U60, P2_U3111);
  nand ginst14896 (P2_R1312_U18, P2_R1312_U144, P2_R1312_U147, P2_R1312_U150, P2_R1312_U151, P2_R1312_U152);
  nand ginst14897 (P2_R1312_U180, P2_R1312_U77, P2_U3112);
  nand ginst14898 (P2_R1312_U181, P2_R1312_U15, P2_R1312_U8, P2_R1312_U86, P2_R1312_U87);
  nand ginst14899 (P2_R1312_U182, P2_R1312_U50, P2_U3117);
  nand ginst14900 (P2_R1312_U183, P2_R1312_U79, P2_U3118);
  nand ginst14901 (P2_R1312_U184, P2_U3152, P2_U3153);
  nand ginst14902 (P2_R1312_U185, P2_R1312_U184, P2_U3120);
  nand ginst14903 (P2_R1312_U186, P2_R1312_U54, P2_U3119);
  or ginst14904 (P2_R1312_U187, P2_U3152, P2_U3153);
  nand ginst14905 (P2_R1312_U188, P2_R1312_U15, P2_R1312_U89, P2_R1312_U90);
  nand ginst14906 (P2_R1312_U189, P2_R1312_U165, P2_R1312_U167, P2_R1312_U168, P2_R1312_U40, P2_U3126);
  not ginst14907 (P2_R1312_U19, P2_U3090);
  nand ginst14908 (P2_R1312_U190, P2_R1312_U21, P2_U3123);
  nand ginst14909 (P2_R1312_U191, P2_R1312_U189, P2_R1312_U190);
  nand ginst14910 (P2_R1312_U192, P2_R1312_U15, P2_R1312_U168, P2_R1312_U8, P2_R1312_U92, P2_R1312_U93);
  nand ginst14911 (P2_R1312_U193, P2_R1312_U16, P2_R1312_U94);
  nand ginst14912 (P2_R1312_U194, P2_R1312_U20, P2_U3125);
  nand ginst14913 (P2_R1312_U195, P2_R1312_U22, P2_U3124);
  nand ginst14914 (P2_R1312_U196, P2_R1312_U193, P2_R1312_U95);
  nand ginst14915 (P2_R1312_U197, P2_R1312_U17, P2_R1312_U196, P2_R1312_U96);
  nand ginst14916 (P2_R1312_U198, P2_R1312_U15, P2_R1312_U166, P2_R1312_U97, P2_R1312_U98);
  nand ginst14917 (P2_R1312_U199, P2_R1312_U100, P2_R1312_U15, P2_R1312_U99);
  not ginst14918 (P2_R1312_U20, P2_U3093);
  nand ginst14919 (P2_R1312_U200, P2_R1312_U101, P2_R1312_U102, P2_R1312_U15, P2_R1312_U166);
  nand ginst14920 (P2_R1312_U201, P2_R1312_U104, P2_R1312_U16, P2_R1312_U169, P2_R1312_U17, P2_U3128);
  nand ginst14921 (P2_R1312_U202, P2_R1312_U105, P2_R1312_U16, P2_R1312_U169, P2_R1312_U17, P2_U3129);
  nand ginst14922 (P2_R1312_U203, P2_R1312_U106, P2_R1312_U107, P2_R1312_U14, P2_R1312_U166, P2_R1312_U17);
  nand ginst14923 (P2_R1312_U204, P2_R1312_U108, P2_R1312_U109, P2_R1312_U11, P2_R1312_U166, P2_R1312_U17);
  nand ginst14924 (P2_R1312_U205, P2_R1312_U110, P2_R1312_U111);
  nand ginst14925 (P2_R1312_U206, P2_R1312_U113, P2_R1312_U114, P2_R1312_U15);
  nand ginst14926 (P2_R1312_U207, P2_R1312_U115, P2_R1312_U15, P2_R1312_U168, P2_R1312_U8, P2_U3146);
  nand ginst14927 (P2_R1312_U208, P2_R1312_U116, P2_R1312_U15, P2_R1312_U168, P2_R1312_U8, P2_U3147);
  nand ginst14928 (P2_R1312_U209, P2_R1312_U11, P2_R1312_U117, P2_R1312_U118, P2_R1312_U17);
  not ginst14929 (P2_R1312_U21, P2_U3091);
  nand ginst14930 (P2_R1312_U210, P2_R1312_U119, P2_R1312_U120, P2_R1312_U15);
  nand ginst14931 (P2_R1312_U211, P2_R1312_U121, P2_R1312_U15, P2_R1312_U8, P2_U3145);
  nand ginst14932 (P2_R1312_U212, P2_R1312_U223, P2_R1312_U226, P2_R1312_U227);
  nand ginst14933 (P2_R1312_U213, P2_R1312_U17, P2_R1312_U19, P2_U3122);
  nand ginst14934 (P2_R1312_U214, P2_R1312_U122, P2_R1312_U123, P2_R1312_U16, P2_R1312_U17, P2_U3130);
  nand ginst14935 (P2_R1312_U215, P2_R1312_U124, P2_R1312_U125, P2_R1312_U14, P2_R1312_U169, P2_R1312_U17);
  nand ginst14936 (P2_R1312_U216, P2_R1312_U11, P2_R1312_U127, P2_R1312_U128, P2_R1312_U16, P2_R1312_U166);
  nand ginst14937 (P2_R1312_U217, P2_R1312_U129, P2_R1312_U130, P2_R1312_U15);
  nand ginst14938 (P2_R1312_U218, P2_R1312_U131, P2_R1312_U132, P2_R1312_U15);
  nand ginst14939 (P2_R1312_U219, P2_R1312_U134, P2_R1312_U135, P2_R1312_U15, P2_R1312_U166);
  not ginst14940 (P2_R1312_U22, P2_U3092);
  nand ginst14941 (P2_R1312_U220, P2_R1312_U137, P2_R1312_U138, P2_R1312_U15);
  nand ginst14942 (P2_R1312_U221, P2_R1312_U50, P2_U3117);
  nand ginst14943 (P2_R1312_U222, P2_R1312_U139, P2_R1312_U140, P2_R1312_U15, P2_R1312_U166, P2_R1312_U8);
  nand ginst14944 (P2_R1312_U223, P2_U3089, P2_U3121);
  nand ginst14945 (P2_R1312_U224, P2_R1312_U26, P2_U3089);
  nand ginst14946 (P2_R1312_U225, P2_R1312_U25, P2_U3121);
  or ginst14947 (P2_R1312_U226, P2_U3121, P2_U3154);
  nand ginst14948 (P2_R1312_U227, P2_R1312_U25, P2_U3154);
  not ginst14949 (P2_R1312_U23, P2_U3126);
  not ginst14950 (P2_R1312_U24, P2_U3123);
  not ginst14951 (P2_R1312_U25, P2_U3089);
  not ginst14952 (P2_R1312_U26, P2_U3121);
  not ginst14953 (P2_R1312_U27, P2_U3105);
  not ginst14954 (P2_R1312_U28, P2_U3106);
  not ginst14955 (P2_R1312_U29, P2_U3108);
  not ginst14956 (P2_R1312_U30, P2_U3107);
  not ginst14957 (P2_R1312_U31, P2_U3109);
  not ginst14958 (P2_R1312_U32, P2_U3110);
  not ginst14959 (P2_R1312_U33, P2_U3111);
  not ginst14960 (P2_R1312_U34, P2_U3112);
  not ginst14961 (P2_R1312_U35, P2_U3115);
  not ginst14962 (P2_R1312_U36, P2_U3116);
  not ginst14963 (P2_R1312_U37, P2_U3114);
  not ginst14964 (P2_R1312_U38, P2_U3113);
  not ginst14965 (P2_R1312_U39, P2_U3104);
  not ginst14966 (P2_R1312_U40, P2_U3094);
  not ginst14967 (P2_R1312_U41, P2_U3102);
  not ginst14968 (P2_R1312_U42, P2_U3101);
  not ginst14969 (P2_R1312_U43, P2_U3103);
  not ginst14970 (P2_R1312_U44, P2_U3100);
  not ginst14971 (P2_R1312_U45, P2_U3099);
  not ginst14972 (P2_R1312_U46, P2_U3095);
  not ginst14973 (P2_R1312_U47, P2_U3097);
  not ginst14974 (P2_R1312_U48, P2_U3098);
  not ginst14975 (P2_R1312_U49, P2_U3096);
  not ginst14976 (P2_R1312_U50, P2_U3149);
  not ginst14977 (P2_R1312_U51, P2_U3117);
  not ginst14978 (P2_R1312_U52, P2_U3118);
  not ginst14979 (P2_R1312_U53, P2_U3119);
  not ginst14980 (P2_R1312_U54, P2_U3151);
  not ginst14981 (P2_R1312_U55, P2_U3127);
  not ginst14982 (P2_R1312_U56, P2_U3125);
  not ginst14983 (P2_R1312_U57, P2_U3124);
  not ginst14984 (P2_R1312_U58, P2_U3140);
  not ginst14985 (P2_R1312_U59, P2_U3141);
  and ginst14986 (P2_R1312_U6, P2_R1312_U170, P2_R1312_U171, P2_R1312_U172);
  not ginst14987 (P2_R1312_U60, P2_U3143);
  not ginst14988 (P2_R1312_U61, P2_U3128);
  not ginst14989 (P2_R1312_U62, P2_U3129);
  not ginst14990 (P2_R1312_U63, P2_U3131);
  not ginst14991 (P2_R1312_U64, P2_U3134);
  not ginst14992 (P2_R1312_U65, P2_U3135);
  not ginst14993 (P2_R1312_U66, P2_U3137);
  not ginst14994 (P2_R1312_U67, P2_U3146);
  not ginst14995 (P2_R1312_U68, P2_U3147);
  not ginst14996 (P2_R1312_U69, P2_U3133);
  and ginst14997 (P2_R1312_U7, P2_R1312_U84, P2_R1312_U85);
  not ginst14998 (P2_R1312_U70, P2_U3139);
  not ginst14999 (P2_R1312_U71, P2_U3145);
  not ginst15000 (P2_R1312_U72, P2_U3130);
  not ginst15001 (P2_R1312_U73, P2_U3132);
  not ginst15002 (P2_R1312_U74, P2_U3136);
  not ginst15003 (P2_R1312_U75, P2_U3138);
  not ginst15004 (P2_R1312_U76, P2_U3142);
  not ginst15005 (P2_R1312_U77, P2_U3144);
  not ginst15006 (P2_R1312_U78, P2_U3148);
  not ginst15007 (P2_R1312_U79, P2_U3150);
  and ginst15008 (P2_R1312_U8, P2_R1312_U173, P2_R1312_U7);
  not ginst15009 (P2_R1312_U80, P2_U3122);
  and ginst15010 (P2_R1312_U81, P2_R1312_U166, P2_R1312_U17);
  and ginst15011 (P2_R1312_U82, P2_R1312_U159, P2_R1312_U160);
  and ginst15012 (P2_R1312_U83, P2_R1312_U158, P2_R1312_U163);
  and ginst15013 (P2_R1312_U84, P2_R1312_U174, P2_R1312_U175, P2_R1312_U176, P2_R1312_U177);
  and ginst15014 (P2_R1312_U85, P2_R1312_U178, P2_R1312_U179, P2_R1312_U180);
  and ginst15015 (P2_R1312_U86, P2_R1312_U166, P2_R1312_U167, P2_R1312_U168, P2_R1312_U51);
  and ginst15016 (P2_R1312_U87, P2_R1312_U12, P2_U3149);
  and ginst15017 (P2_R1312_U88, P2_R1312_U173, P2_R1312_U186);
  and ginst15018 (P2_R1312_U89, P2_R1312_U166, P2_R1312_U167, P2_R1312_U168, P2_R1312_U185, P2_R1312_U88);
  and ginst15019 (P2_R1312_U9, P2_R1312_U182, P2_R1312_U183);
  and ginst15020 (P2_R1312_U90, P2_R1312_U187, P2_R1312_U7, P2_R1312_U91);
  and ginst15021 (P2_R1312_U91, P2_R1312_U12, P2_R1312_U9);
  and ginst15022 (P2_R1312_U92, P2_R1312_U166, P2_R1312_U167, P2_R1312_U53);
  and ginst15023 (P2_R1312_U93, P2_R1312_U12, P2_R1312_U9, P2_U3151);
  and ginst15024 (P2_R1312_U94, P2_R1312_U46, P2_U3127);
  and ginst15025 (P2_R1312_U95, P2_R1312_U194, P2_R1312_U195);
  and ginst15026 (P2_R1312_U96, P2_R1312_U166, P2_R1312_U167, P2_R1312_U168);
  and ginst15027 (P2_R1312_U97, P2_R1312_U167, P2_R1312_U168, P2_R1312_U173, P2_R1312_U29);
  and ginst15028 (P2_R1312_U98, P2_R1312_U174, P2_R1312_U176, P2_U3140);
  and ginst15029 (P2_R1312_U99, P2_R1312_U166, P2_R1312_U167, P2_R1312_U168, P2_R1312_U31);
  nand ginst15030 (P2_R1335_U10, P2_R1335_U7, P2_U3061);
  not ginst15031 (P2_R1335_U6, P2_U3061);
  not ginst15032 (P2_R1335_U7, P2_U3058);
  and ginst15033 (P2_R1335_U8, P2_R1335_U10, P2_R1335_U9);
  nand ginst15034 (P2_R1335_U9, P2_R1335_U6, P2_U3058);
  and ginst15035 (P2_SUB_1108_U10, P2_SUB_1108_U143, P2_SUB_1108_U166);
  not ginst15036 (P2_SUB_1108_U100, P2_IR_REG_5__SCAN_IN);
  and ginst15037 (P2_SUB_1108_U101, P2_SUB_1108_U177, P2_SUB_1108_U178);
  not ginst15038 (P2_SUB_1108_U102, P2_IR_REG_31__SCAN_IN);
  not ginst15039 (P2_SUB_1108_U103, P2_IR_REG_30__SCAN_IN);
  and ginst15040 (P2_SUB_1108_U104, P2_SUB_1108_U181, P2_SUB_1108_U182);
  not ginst15041 (P2_SUB_1108_U105, P2_IR_REG_28__SCAN_IN);
  nand ginst15042 (P2_SUB_1108_U106, P2_SUB_1108_U72, P2_SUB_1108_U77);
  and ginst15043 (P2_SUB_1108_U107, P2_SUB_1108_U183, P2_SUB_1108_U184);
  not ginst15044 (P2_SUB_1108_U108, P2_IR_REG_27__SCAN_IN);
  nand ginst15045 (P2_SUB_1108_U109, P2_SUB_1108_U82, P2_SUB_1108_U87);
  and ginst15046 (P2_SUB_1108_U11, P2_SUB_1108_U165, P2_SUB_1108_U30);
  and ginst15047 (P2_SUB_1108_U110, P2_SUB_1108_U185, P2_SUB_1108_U186);
  not ginst15048 (P2_SUB_1108_U111, P2_IR_REG_25__SCAN_IN);
  and ginst15049 (P2_SUB_1108_U112, P2_SUB_1108_U187, P2_SUB_1108_U188);
  not ginst15050 (P2_SUB_1108_U113, P2_IR_REG_22__SCAN_IN);
  and ginst15051 (P2_SUB_1108_U114, P2_SUB_1108_U189, P2_SUB_1108_U190);
  not ginst15052 (P2_SUB_1108_U115, P2_IR_REG_21__SCAN_IN);
  and ginst15053 (P2_SUB_1108_U116, P2_SUB_1108_U191, P2_SUB_1108_U192);
  not ginst15054 (P2_SUB_1108_U117, P2_IR_REG_20__SCAN_IN);
  nand ginst15055 (P2_SUB_1108_U118, P2_SUB_1108_U122, P2_SUB_1108_U145);
  and ginst15056 (P2_SUB_1108_U119, P2_SUB_1108_U193, P2_SUB_1108_U194);
  and ginst15057 (P2_SUB_1108_U12, P2_SUB_1108_U164, P2_SUB_1108_U36);
  not ginst15058 (P2_SUB_1108_U120, P2_IR_REG_1__SCAN_IN);
  not ginst15059 (P2_SUB_1108_U121, P2_IR_REG_0__SCAN_IN);
  not ginst15060 (P2_SUB_1108_U122, P2_IR_REG_19__SCAN_IN);
  and ginst15061 (P2_SUB_1108_U123, P2_SUB_1108_U197, P2_SUB_1108_U198);
  not ginst15062 (P2_SUB_1108_U124, P2_IR_REG_17__SCAN_IN);
  and ginst15063 (P2_SUB_1108_U125, P2_SUB_1108_U199, P2_SUB_1108_U200);
  not ginst15064 (P2_SUB_1108_U126, P2_IR_REG_13__SCAN_IN);
  and ginst15065 (P2_SUB_1108_U127, P2_SUB_1108_U201, P2_SUB_1108_U202);
  nand ginst15066 (P2_SUB_1108_U128, P2_SUB_1108_U174, P2_SUB_1108_U28);
  not ginst15067 (P2_SUB_1108_U129, P2_SUB_1108_U25);
  and ginst15068 (P2_SUB_1108_U13, P2_SUB_1108_U162, P2_SUB_1108_U32);
  not ginst15069 (P2_SUB_1108_U130, P2_SUB_1108_U26);
  nand ginst15070 (P2_SUB_1108_U131, P2_SUB_1108_U130, P2_SUB_1108_U27);
  not ginst15071 (P2_SUB_1108_U132, P2_SUB_1108_U24);
  nand ginst15072 (P2_SUB_1108_U133, P2_IR_REG_8__SCAN_IN, P2_SUB_1108_U131);
  nand ginst15073 (P2_SUB_1108_U134, P2_IR_REG_7__SCAN_IN, P2_SUB_1108_U26);
  nand ginst15074 (P2_SUB_1108_U135, P2_SUB_1108_U100, P2_SUB_1108_U129);
  nand ginst15075 (P2_SUB_1108_U136, P2_IR_REG_6__SCAN_IN, P2_SUB_1108_U135);
  nand ginst15076 (P2_SUB_1108_U137, P2_IR_REG_4__SCAN_IN, P2_SUB_1108_U128);
  nand ginst15077 (P2_SUB_1108_U138, P2_IR_REG_3__SCAN_IN, P2_SUB_1108_U23);
  not ginst15078 (P2_SUB_1108_U139, P2_SUB_1108_U40);
  and ginst15079 (P2_SUB_1108_U14, P2_SUB_1108_U160, P2_SUB_1108_U33);
  nand ginst15080 (P2_SUB_1108_U140, P2_SUB_1108_U139, P2_SUB_1108_U41);
  not ginst15081 (P2_SUB_1108_U141, P2_SUB_1108_U37);
  not ginst15082 (P2_SUB_1108_U142, P2_SUB_1108_U38);
  nand ginst15083 (P2_SUB_1108_U143, P2_SUB_1108_U142, P2_SUB_1108_U39);
  not ginst15084 (P2_SUB_1108_U144, P2_SUB_1108_U30);
  not ginst15085 (P2_SUB_1108_U145, P2_SUB_1108_U36);
  not ginst15086 (P2_SUB_1108_U146, P2_SUB_1108_U118);
  not ginst15087 (P2_SUB_1108_U147, P2_SUB_1108_U31);
  not ginst15088 (P2_SUB_1108_U148, P2_SUB_1108_U35);
  not ginst15089 (P2_SUB_1108_U149, P2_SUB_1108_U32);
  and ginst15090 (P2_SUB_1108_U15, P2_SUB_1108_U109, P2_SUB_1108_U159);
  not ginst15091 (P2_SUB_1108_U150, P2_SUB_1108_U33);
  not ginst15092 (P2_SUB_1108_U151, P2_SUB_1108_U109);
  not ginst15093 (P2_SUB_1108_U152, P2_SUB_1108_U106);
  not ginst15094 (P2_SUB_1108_U153, P2_SUB_1108_U29);
  or ginst15095 (P2_SUB_1108_U154, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN);
  nand ginst15096 (P2_SUB_1108_U155, P2_IR_REG_2__SCAN_IN, P2_SUB_1108_U154);
  nand ginst15097 (P2_SUB_1108_U156, P2_SUB_1108_U62, P2_SUB_1108_U67);
  nand ginst15098 (P2_SUB_1108_U157, P2_IR_REG_29__SCAN_IN, P2_SUB_1108_U156);
  nand ginst15099 (P2_SUB_1108_U158, P2_SUB_1108_U111, P2_SUB_1108_U150);
  nand ginst15100 (P2_SUB_1108_U159, P2_IR_REG_26__SCAN_IN, P2_SUB_1108_U158);
  and ginst15101 (P2_SUB_1108_U16, P2_SUB_1108_U157, P2_SUB_1108_U29);
  nand ginst15102 (P2_SUB_1108_U160, P2_IR_REG_24__SCAN_IN, P2_SUB_1108_U32);
  nand ginst15103 (P2_SUB_1108_U161, P2_SUB_1108_U113, P2_SUB_1108_U148);
  nand ginst15104 (P2_SUB_1108_U162, P2_IR_REG_23__SCAN_IN, P2_SUB_1108_U161);
  nand ginst15105 (P2_SUB_1108_U163, P2_SUB_1108_U124, P2_SUB_1108_U144);
  nand ginst15106 (P2_SUB_1108_U164, P2_IR_REG_18__SCAN_IN, P2_SUB_1108_U163);
  nand ginst15107 (P2_SUB_1108_U165, P2_IR_REG_16__SCAN_IN, P2_SUB_1108_U143);
  nand ginst15108 (P2_SUB_1108_U166, P2_IR_REG_15__SCAN_IN, P2_SUB_1108_U38);
  nand ginst15109 (P2_SUB_1108_U167, P2_SUB_1108_U126, P2_SUB_1108_U141);
  nand ginst15110 (P2_SUB_1108_U168, P2_IR_REG_14__SCAN_IN, P2_SUB_1108_U167);
  nand ginst15111 (P2_SUB_1108_U169, P2_IR_REG_12__SCAN_IN, P2_SUB_1108_U140);
  and ginst15112 (P2_SUB_1108_U17, P2_SUB_1108_U155, P2_SUB_1108_U23);
  nand ginst15113 (P2_SUB_1108_U170, P2_IR_REG_11__SCAN_IN, P2_SUB_1108_U40);
  nand ginst15114 (P2_SUB_1108_U171, P2_SUB_1108_U132, P2_SUB_1108_U98);
  nand ginst15115 (P2_SUB_1108_U172, P2_IR_REG_10__SCAN_IN, P2_SUB_1108_U171);
  nand ginst15116 (P2_SUB_1108_U173, P2_SUB_1108_U103, P2_SUB_1108_U153);
  not ginst15117 (P2_SUB_1108_U174, P2_SUB_1108_U23);
  nand ginst15118 (P2_SUB_1108_U175, P2_IR_REG_9__SCAN_IN, P2_SUB_1108_U24);
  nand ginst15119 (P2_SUB_1108_U176, P2_SUB_1108_U132, P2_SUB_1108_U98);
  nand ginst15120 (P2_SUB_1108_U177, P2_IR_REG_5__SCAN_IN, P2_SUB_1108_U25);
  nand ginst15121 (P2_SUB_1108_U178, P2_SUB_1108_U100, P2_SUB_1108_U129);
  nand ginst15122 (P2_SUB_1108_U179, P2_SUB_1108_U102, P2_SUB_1108_U173);
  and ginst15123 (P2_SUB_1108_U18, P2_SUB_1108_U128, P2_SUB_1108_U138);
  nand ginst15124 (P2_SUB_1108_U180, P2_IR_REG_31__SCAN_IN, P2_SUB_1108_U103, P2_SUB_1108_U153);
  nand ginst15125 (P2_SUB_1108_U181, P2_IR_REG_30__SCAN_IN, P2_SUB_1108_U29);
  nand ginst15126 (P2_SUB_1108_U182, P2_SUB_1108_U103, P2_SUB_1108_U153);
  nand ginst15127 (P2_SUB_1108_U183, P2_IR_REG_28__SCAN_IN, P2_SUB_1108_U106);
  nand ginst15128 (P2_SUB_1108_U184, P2_SUB_1108_U105, P2_SUB_1108_U152);
  nand ginst15129 (P2_SUB_1108_U185, P2_IR_REG_27__SCAN_IN, P2_SUB_1108_U109);
  nand ginst15130 (P2_SUB_1108_U186, P2_SUB_1108_U108, P2_SUB_1108_U151);
  nand ginst15131 (P2_SUB_1108_U187, P2_IR_REG_25__SCAN_IN, P2_SUB_1108_U33);
  nand ginst15132 (P2_SUB_1108_U188, P2_SUB_1108_U111, P2_SUB_1108_U150);
  nand ginst15133 (P2_SUB_1108_U189, P2_IR_REG_22__SCAN_IN, P2_SUB_1108_U35);
  and ginst15134 (P2_SUB_1108_U19, P2_SUB_1108_U137, P2_SUB_1108_U25);
  nand ginst15135 (P2_SUB_1108_U190, P2_SUB_1108_U113, P2_SUB_1108_U148);
  nand ginst15136 (P2_SUB_1108_U191, P2_IR_REG_21__SCAN_IN, P2_SUB_1108_U31);
  nand ginst15137 (P2_SUB_1108_U192, P2_SUB_1108_U115, P2_SUB_1108_U147);
  nand ginst15138 (P2_SUB_1108_U193, P2_IR_REG_20__SCAN_IN, P2_SUB_1108_U118);
  nand ginst15139 (P2_SUB_1108_U194, P2_SUB_1108_U117, P2_SUB_1108_U146);
  nand ginst15140 (P2_SUB_1108_U195, P2_IR_REG_1__SCAN_IN, P2_SUB_1108_U121);
  nand ginst15141 (P2_SUB_1108_U196, P2_IR_REG_0__SCAN_IN, P2_SUB_1108_U120);
  nand ginst15142 (P2_SUB_1108_U197, P2_IR_REG_19__SCAN_IN, P2_SUB_1108_U36);
  nand ginst15143 (P2_SUB_1108_U198, P2_SUB_1108_U122, P2_SUB_1108_U145);
  nand ginst15144 (P2_SUB_1108_U199, P2_IR_REG_17__SCAN_IN, P2_SUB_1108_U30);
  and ginst15145 (P2_SUB_1108_U20, P2_SUB_1108_U136, P2_SUB_1108_U26);
  nand ginst15146 (P2_SUB_1108_U200, P2_SUB_1108_U124, P2_SUB_1108_U144);
  nand ginst15147 (P2_SUB_1108_U201, P2_IR_REG_13__SCAN_IN, P2_SUB_1108_U37);
  nand ginst15148 (P2_SUB_1108_U202, P2_SUB_1108_U126, P2_SUB_1108_U141);
  and ginst15149 (P2_SUB_1108_U21, P2_SUB_1108_U131, P2_SUB_1108_U134);
  and ginst15150 (P2_SUB_1108_U22, P2_SUB_1108_U133, P2_SUB_1108_U24);
  or ginst15151 (P2_SUB_1108_U23, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN, P2_IR_REG_2__SCAN_IN);
  nand ginst15152 (P2_SUB_1108_U24, P2_SUB_1108_U174, P2_SUB_1108_U44, P2_SUB_1108_U45);
  nand ginst15153 (P2_SUB_1108_U25, P2_SUB_1108_U174, P2_SUB_1108_U46);
  nand ginst15154 (P2_SUB_1108_U26, P2_SUB_1108_U129, P2_SUB_1108_U47);
  not ginst15155 (P2_SUB_1108_U27, P2_IR_REG_7__SCAN_IN);
  not ginst15156 (P2_SUB_1108_U28, P2_IR_REG_3__SCAN_IN);
  nand ginst15157 (P2_SUB_1108_U29, P2_SUB_1108_U52, P2_SUB_1108_U57);
  nand ginst15158 (P2_SUB_1108_U30, P2_SUB_1108_U88, P2_SUB_1108_U89, P2_SUB_1108_U90, P2_SUB_1108_U91);
  nand ginst15159 (P2_SUB_1108_U31, P2_SUB_1108_U144, P2_SUB_1108_U92);
  nand ginst15160 (P2_SUB_1108_U32, P2_SUB_1108_U147, P2_SUB_1108_U93);
  nand ginst15161 (P2_SUB_1108_U33, P2_SUB_1108_U149, P2_SUB_1108_U34);
  not ginst15162 (P2_SUB_1108_U34, P2_IR_REG_24__SCAN_IN);
  nand ginst15163 (P2_SUB_1108_U35, P2_SUB_1108_U115, P2_SUB_1108_U147);
  nand ginst15164 (P2_SUB_1108_U36, P2_SUB_1108_U144, P2_SUB_1108_U94);
  nand ginst15165 (P2_SUB_1108_U37, P2_SUB_1108_U132, P2_SUB_1108_U95);
  nand ginst15166 (P2_SUB_1108_U38, P2_SUB_1108_U141, P2_SUB_1108_U96);
  not ginst15167 (P2_SUB_1108_U39, P2_IR_REG_15__SCAN_IN);
  nand ginst15168 (P2_SUB_1108_U40, P2_SUB_1108_U132, P2_SUB_1108_U97);
  not ginst15169 (P2_SUB_1108_U41, P2_IR_REG_11__SCAN_IN);
  nand ginst15170 (P2_SUB_1108_U42, P2_SUB_1108_U195, P2_SUB_1108_U196);
  nand ginst15171 (P2_SUB_1108_U43, P2_SUB_1108_U179, P2_SUB_1108_U180);
  nor ginst15172 (P2_SUB_1108_U44, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN, P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN);
  nor ginst15173 (P2_SUB_1108_U45, P2_IR_REG_7__SCAN_IN, P2_IR_REG_8__SCAN_IN);
  nor ginst15174 (P2_SUB_1108_U46, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN);
  nor ginst15175 (P2_SUB_1108_U47, P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN);
  nor ginst15176 (P2_SUB_1108_U48, P2_IR_REG_10__SCAN_IN, P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN);
  nor ginst15177 (P2_SUB_1108_U49, P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN, P2_IR_REG_17__SCAN_IN);
  nor ginst15178 (P2_SUB_1108_U50, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN);
  nor ginst15179 (P2_SUB_1108_U51, P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN);
  and ginst15180 (P2_SUB_1108_U52, P2_SUB_1108_U48, P2_SUB_1108_U49, P2_SUB_1108_U50, P2_SUB_1108_U51);
  nor ginst15181 (P2_SUB_1108_U53, P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN, P2_IR_REG_26__SCAN_IN);
  nor ginst15182 (P2_SUB_1108_U54, P2_IR_REG_2__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN, P2_IR_REG_29__SCAN_IN);
  nor ginst15183 (P2_SUB_1108_U55, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN, P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN);
  nor ginst15184 (P2_SUB_1108_U56, P2_IR_REG_7__SCAN_IN, P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN);
  and ginst15185 (P2_SUB_1108_U57, P2_SUB_1108_U53, P2_SUB_1108_U54, P2_SUB_1108_U55, P2_SUB_1108_U56);
  nor ginst15186 (P2_SUB_1108_U58, P2_IR_REG_10__SCAN_IN, P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN);
  nor ginst15187 (P2_SUB_1108_U59, P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN, P2_IR_REG_17__SCAN_IN);
  and ginst15188 (P2_SUB_1108_U6, P2_SUB_1108_U172, P2_SUB_1108_U40);
  nor ginst15189 (P2_SUB_1108_U60, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN);
  nor ginst15190 (P2_SUB_1108_U61, P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN);
  and ginst15191 (P2_SUB_1108_U62, P2_SUB_1108_U58, P2_SUB_1108_U59, P2_SUB_1108_U60, P2_SUB_1108_U61);
  nor ginst15192 (P2_SUB_1108_U63, P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN, P2_IR_REG_26__SCAN_IN);
  nor ginst15193 (P2_SUB_1108_U64, P2_IR_REG_2__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN);
  nor ginst15194 (P2_SUB_1108_U65, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN, P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN);
  nor ginst15195 (P2_SUB_1108_U66, P2_IR_REG_7__SCAN_IN, P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN);
  and ginst15196 (P2_SUB_1108_U67, P2_SUB_1108_U63, P2_SUB_1108_U64, P2_SUB_1108_U65, P2_SUB_1108_U66);
  nor ginst15197 (P2_SUB_1108_U68, P2_IR_REG_10__SCAN_IN, P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN);
  nor ginst15198 (P2_SUB_1108_U69, P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN);
  and ginst15199 (P2_SUB_1108_U7, P2_SUB_1108_U140, P2_SUB_1108_U170);
  nor ginst15200 (P2_SUB_1108_U70, P2_IR_REG_1__SCAN_IN, P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN);
  nor ginst15201 (P2_SUB_1108_U71, P2_IR_REG_0__SCAN_IN, P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN);
  and ginst15202 (P2_SUB_1108_U72, P2_SUB_1108_U68, P2_SUB_1108_U69, P2_SUB_1108_U70, P2_SUB_1108_U71);
  nor ginst15203 (P2_SUB_1108_U73, P2_IR_REG_22__SCAN_IN, P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN);
  nor ginst15204 (P2_SUB_1108_U74, P2_IR_REG_2__SCAN_IN, P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN);
  nor ginst15205 (P2_SUB_1108_U75, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN, P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN);
  nor ginst15206 (P2_SUB_1108_U76, P2_IR_REG_7__SCAN_IN, P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN);
  and ginst15207 (P2_SUB_1108_U77, P2_SUB_1108_U73, P2_SUB_1108_U74, P2_SUB_1108_U75, P2_SUB_1108_U76);
  nor ginst15208 (P2_SUB_1108_U78, P2_IR_REG_10__SCAN_IN, P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN);
  nor ginst15209 (P2_SUB_1108_U79, P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN);
  and ginst15210 (P2_SUB_1108_U8, P2_SUB_1108_U169, P2_SUB_1108_U37);
  nor ginst15211 (P2_SUB_1108_U80, P2_IR_REG_1__SCAN_IN, P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN);
  nor ginst15212 (P2_SUB_1108_U81, P2_IR_REG_0__SCAN_IN, P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN);
  and ginst15213 (P2_SUB_1108_U82, P2_SUB_1108_U78, P2_SUB_1108_U79, P2_SUB_1108_U80, P2_SUB_1108_U81);
  nor ginst15214 (P2_SUB_1108_U83, P2_IR_REG_22__SCAN_IN, P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN);
  nor ginst15215 (P2_SUB_1108_U84, P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_26__SCAN_IN);
  nor ginst15216 (P2_SUB_1108_U85, P2_IR_REG_4__SCAN_IN, P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN);
  nor ginst15217 (P2_SUB_1108_U86, P2_IR_REG_7__SCAN_IN, P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN);
  and ginst15218 (P2_SUB_1108_U87, P2_SUB_1108_U83, P2_SUB_1108_U84, P2_SUB_1108_U85, P2_SUB_1108_U86);
  nor ginst15219 (P2_SUB_1108_U88, P2_IR_REG_10__SCAN_IN, P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN, P2_IR_REG_14__SCAN_IN);
  nor ginst15220 (P2_SUB_1108_U89, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN);
  and ginst15221 (P2_SUB_1108_U9, P2_SUB_1108_U168, P2_SUB_1108_U38);
  nor ginst15222 (P2_SUB_1108_U90, P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN, P2_IR_REG_5__SCAN_IN);
  nor ginst15223 (P2_SUB_1108_U91, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN, P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN);
  nor ginst15224 (P2_SUB_1108_U92, P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN, P2_IR_REG_20__SCAN_IN);
  nor ginst15225 (P2_SUB_1108_U93, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN, P2_IR_REG_23__SCAN_IN);
  nor ginst15226 (P2_SUB_1108_U94, P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN);
  nor ginst15227 (P2_SUB_1108_U95, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN, P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN);
  nor ginst15228 (P2_SUB_1108_U96, P2_IR_REG_13__SCAN_IN, P2_IR_REG_14__SCAN_IN);
  nor ginst15229 (P2_SUB_1108_U97, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN);
  not ginst15230 (P2_SUB_1108_U98, P2_IR_REG_9__SCAN_IN);
  and ginst15231 (P2_SUB_1108_U99, P2_SUB_1108_U175, P2_SUB_1108_U176);
  and ginst15232 (P2_U3014, P2_U3924, P2_U5671);
  and ginst15233 (P2_U3015, P2_U3419, P2_U3937);
  and ginst15234 (P2_U3016, P2_U3570, P2_U3575);
  and ginst15235 (P2_U3017, P2_U3423, P2_U5688);
  and ginst15236 (P2_U3018, P2_U3423, P2_U3426);
  and ginst15237 (P2_U3019, P2_U3421, P2_U3422);
  and ginst15238 (P2_U3020, P2_U3421, P2_U5680);
  and ginst15239 (P2_U3021, P2_U3422, P2_U5677);
  and ginst15240 (P2_U3022, P2_U5677, P2_U5680);
  and ginst15241 (P2_U3023, P2_STATE_REG_SCAN_IN, P2_U3048);
  and ginst15242 (P2_U3024, P2_U3401, P2_U3757);
  and ginst15243 (P2_U3025, P2_U3976, P2_U5671);
  and ginst15244 (P2_U3026, P2_U3963, P2_U5683);
  and ginst15245 (P2_U3027, P2_U3944, P2_U5671);
  and ginst15246 (P2_U3028, P2_U3803, P2_U3946);
  and ginst15247 (P2_U3029, P2_R1299_U6, P2_U3411);
  and ginst15248 (P2_U3030, P2_STATE_REG_SCAN_IN, P2_U3329);
  and ginst15249 (P2_U3031, P2_U3932, P2_U3964);
  and ginst15250 (P2_U3032, P2_U3398, P2_U3964);
  and ginst15251 (P2_U3033, P2_U3933, P2_U3964);
  and ginst15252 (P2_U3034, P2_U3938, P2_U3964);
  and ginst15253 (P2_U3035, P2_U3423, P2_U3963);
  and ginst15254 (P2_U3036, P2_U3946, P2_U5683);
  and ginst15255 (P2_U3037, P2_U3026, P2_U3964);
  and ginst15256 (P2_U3038, P2_U3423, P2_U3946);
  and ginst15257 (P2_U3039, P2_U4854, P2_U5688);
  and ginst15258 (P2_U3040, P2_U3024, P2_U5688);
  and ginst15259 (P2_U3041, P2_U4854, P2_U5683);
  and ginst15260 (P2_U3042, P2_U3024, P2_U5683);
  and ginst15261 (P2_U3043, P2_U3018, P2_U4854);
  and ginst15262 (P2_U3044, P2_U3018, P2_U3024);
  and ginst15263 (P2_U3045, P2_U3023, P2_U3401);
  and ginst15264 (P2_U3046, P2_STATE_REG_SCAN_IN, P2_U5184);
  and ginst15265 (P2_U3047, P2_U3023, P2_U5186);
  and ginst15266 (P2_U3048, P2_U3396, P2_U5658);
  and ginst15267 (P2_U3049, P2_U3418, P2_U5668);
  and ginst15268 (P2_U3050, P2_U3016, P2_U3576);
  and ginst15269 (P2_U3051, P2_U3337, P2_U3338, P2_U3341, P2_U3392, P2_U3402);
  and ginst15270 (P2_U3052, P2_STATE_REG_SCAN_IN, P2_U3399);
  and ginst15271 (P2_U3053, P2_U3819, P2_U3820, P2_U5439);
  and ginst15272 (P2_U3054, P2_U5460, P2_U5461);
  nand ginst15273 (P2_U3055, P2_U4610, P2_U4611, P2_U4612, P2_U4613);
  nand ginst15274 (P2_U3056, P2_U4629, P2_U4630, P2_U4631, P2_U4632);
  nand ginst15275 (P2_U3057, P2_U4648, P2_U4649, P2_U4650, P2_U4651);
  nand ginst15276 (P2_U3058, P2_U4687, P2_U4688, P2_U4689);
  nand ginst15277 (P2_U3059, P2_U4591, P2_U4592, P2_U4593, P2_U4594);
  nand ginst15278 (P2_U3060, P2_U4572, P2_U4573, P2_U4574, P2_U4575);
  nand ginst15279 (P2_U3061, P2_U4667, P2_U4668, P2_U4669);
  nand ginst15280 (P2_U3062, P2_U4173, P2_U4174, P2_U4175, P2_U4176);
  nand ginst15281 (P2_U3063, P2_U4515, P2_U4516, P2_U4517, P2_U4518);
  nand ginst15282 (P2_U3064, P2_U4287, P2_U4288, P2_U4289, P2_U4290);
  nand ginst15283 (P2_U3065, P2_U4306, P2_U4307, P2_U4308, P2_U4309);
  nand ginst15284 (P2_U3066, P2_U4154, P2_U4155, P2_U4156, P2_U4157);
  nand ginst15285 (P2_U3067, P2_U4553, P2_U4554, P2_U4555, P2_U4556);
  nand ginst15286 (P2_U3068, P2_U4534, P2_U4535, P2_U4536, P2_U4537);
  nand ginst15287 (P2_U3069, P2_U4192, P2_U4193, P2_U4194, P2_U4195);
  nand ginst15288 (P2_U3070, P2_U4130, P2_U4131, P2_U4132, P2_U4133);
  nand ginst15289 (P2_U3071, P2_U4420, P2_U4421, P2_U4422, P2_U4423);
  nand ginst15290 (P2_U3072, P2_U4230, P2_U4231, P2_U4232, P2_U4233);
  nand ginst15291 (P2_U3073, P2_U4211, P2_U4212, P2_U4213, P2_U4214);
  nand ginst15292 (P2_U3074, P2_U4325, P2_U4326, P2_U4327, P2_U4328);
  nand ginst15293 (P2_U3075, P2_U4401, P2_U4402, P2_U4403, P2_U4404);
  nand ginst15294 (P2_U3076, P2_U4382, P2_U4383, P2_U4384, P2_U4385);
  nand ginst15295 (P2_U3077, P2_U4496, P2_U4497, P2_U4498, P2_U4499);
  nand ginst15296 (P2_U3078, P2_U4477, P2_U4478, P2_U4479, P2_U4480);
  nand ginst15297 (P2_U3079, P2_U4135, P2_U4136, P2_U4137, P2_U4138);
  nand ginst15298 (P2_U3080, P2_U4111, P2_U4112, P2_U4113, P2_U4114);
  nand ginst15299 (P2_U3081, P2_U4363, P2_U4364, P2_U4365, P2_U4366);
  nand ginst15300 (P2_U3082, P2_U4344, P2_U4345, P2_U4346, P2_U4347);
  nand ginst15301 (P2_U3083, P2_U4458, P2_U4459, P2_U4460, P2_U4461);
  nand ginst15302 (P2_U3084, P2_U4439, P2_U4440, P2_U4441, P2_U4442);
  nand ginst15303 (P2_U3085, P2_U4268, P2_U4269, P2_U4270, P2_U4271);
  nand ginst15304 (P2_U3086, P2_U4249, P2_U4250, P2_U4251, P2_U4252);
  nand ginst15305 (P2_U3087, P2_U3815, P2_U5434);
  not ginst15306 (P2_U3088, P2_STATE_REG_SCAN_IN);
  nand ginst15307 (P2_U3089, P2_U5556, P2_U5557);
  nand ginst15308 (P2_U3090, P2_U5558, P2_U5559);
  nand ginst15309 (P2_U3091, P2_U3859, P2_U5563);
  nand ginst15310 (P2_U3092, P2_U3860, P2_U5566);
  nand ginst15311 (P2_U3093, P2_U3861, P2_U5569);
  nand ginst15312 (P2_U3094, P2_U3862, P2_U5572);
  nand ginst15313 (P2_U3095, P2_U3863, P2_U5575);
  nand ginst15314 (P2_U3096, P2_U3864, P2_U5578);
  nand ginst15315 (P2_U3097, P2_U3865, P2_U5581);
  nand ginst15316 (P2_U3098, P2_U3866, P2_U5584);
  nand ginst15317 (P2_U3099, P2_U3867, P2_U5587);
  nand ginst15318 (P2_U3100, P2_U3868, P2_U5590);
  nand ginst15319 (P2_U3101, P2_U3869, P2_U5596);
  nand ginst15320 (P2_U3102, P2_U3870, P2_U5599);
  nand ginst15321 (P2_U3103, P2_U3871, P2_U5602);
  nand ginst15322 (P2_U3104, P2_U3872, P2_U5605);
  nand ginst15323 (P2_U3105, P2_U3873, P2_U5608);
  nand ginst15324 (P2_U3106, P2_U3874, P2_U5611);
  nand ginst15325 (P2_U3107, P2_U3875, P2_U5614);
  nand ginst15326 (P2_U3108, P2_U3876, P2_U5617);
  nand ginst15327 (P2_U3109, P2_U3877, P2_U5620);
  nand ginst15328 (P2_U3110, P2_U3878, P2_U5623);
  nand ginst15329 (P2_U3111, P2_U3857, P2_U5538);
  nand ginst15330 (P2_U3112, P2_U3858, P2_U5541);
  nand ginst15331 (P2_U3113, P2_U5544, P2_U5545, P2_U5546);
  nand ginst15332 (P2_U3114, P2_U5547, P2_U5548, P2_U5549);
  nand ginst15333 (P2_U3115, P2_U5550, P2_U5551, P2_U5552);
  nand ginst15334 (P2_U3116, P2_U5553, P2_U5554, P2_U5555);
  nand ginst15335 (P2_U3117, P2_U5560, P2_U5561, P2_U5562);
  nand ginst15336 (P2_U3118, P2_U5593, P2_U5594, P2_U5595);
  nand ginst15337 (P2_U3119, P2_U5626, P2_U5627, P2_U5628);
  nand ginst15338 (P2_U3120, P2_U5629, P2_U5630);
  and ginst15339 (P2_U3121, P2_U5632, P2_U5637, P2_U5638);
  nand ginst15340 (P2_U3122, P2_U5462, P2_U5463, P2_U5464);
  nand ginst15341 (P2_U3123, P2_U3831, P2_U5469, P2_U5470);
  nand ginst15342 (P2_U3124, P2_U3832, P2_U5472, P2_U5473);
  nand ginst15343 (P2_U3125, P2_U3833, P2_U5475, P2_U5476);
  nand ginst15344 (P2_U3126, P2_U3834, P2_U5478, P2_U5479);
  nand ginst15345 (P2_U3127, P2_U3835, P2_U5481, P2_U5482);
  nand ginst15346 (P2_U3128, P2_U3836, P2_U5484, P2_U5485);
  nand ginst15347 (P2_U3129, P2_U3837, P2_U5487, P2_U5488);
  nand ginst15348 (P2_U3130, P2_U3838, P2_U5490, P2_U5491);
  nand ginst15349 (P2_U3131, P2_U3839, P2_U5493, P2_U5494);
  nand ginst15350 (P2_U3132, P2_U3840, P2_U5496, P2_U5497);
  nand ginst15351 (P2_U3133, P2_U3843, P2_U5502, P2_U5503);
  nand ginst15352 (P2_U3134, P2_U3844, P2_U5505, P2_U5506);
  nand ginst15353 (P2_U3135, P2_U3845, P2_U5508, P2_U5509);
  nand ginst15354 (P2_U3136, P2_U3846, P2_U5511, P2_U5512);
  nand ginst15355 (P2_U3137, P2_U3847, P2_U5514, P2_U5515);
  nand ginst15356 (P2_U3138, P2_U3848, P2_U5517, P2_U5518);
  nand ginst15357 (P2_U3139, P2_U3849, P2_U5520, P2_U5521);
  nand ginst15358 (P2_U3140, P2_U3850, P2_U5523, P2_U5524);
  nand ginst15359 (P2_U3141, P2_U3851, P2_U5525, P2_U5526);
  nand ginst15360 (P2_U3142, P2_U3852, P2_U5528, P2_U5529);
  nand ginst15361 (P2_U3143, P2_U3821, P2_U5442, P2_U5443);
  nand ginst15362 (P2_U3144, P2_U3822, P2_U5445, P2_U5446);
  nand ginst15363 (P2_U3145, P2_U3823, P2_U5448, P2_U5449);
  nand ginst15364 (P2_U3146, P2_U3824, P2_U5451, P2_U5452);
  nand ginst15365 (P2_U3147, P2_U3825, P2_U5454, P2_U5455);
  nand ginst15366 (P2_U3148, P2_U3826, P2_U5458);
  nand ginst15367 (P2_U3149, P2_U3829, P2_U5466);
  nand ginst15368 (P2_U3150, P2_U3841, P2_U5499);
  nand ginst15369 (P2_U3151, P2_U3853, P2_U5532);
  nand ginst15370 (P2_U3152, P2_U3855, P2_U5535);
  nand ginst15371 (P2_U3153, P2_U3345, P2_U3415, P2_U3817);
  nand ginst15372 (P2_U3154, P2_U3015, P2_U5658);
  and ginst15373 (P2_U3155, P2_U3056, P2_U5437);
  and ginst15374 (P2_U3156, P2_U3055, P2_U5437);
  and ginst15375 (P2_U3157, P2_U3059, P2_U5437);
  and ginst15376 (P2_U3158, P2_U3060, P2_U5437);
  and ginst15377 (P2_U3159, P2_U3067, P2_U5437);
  and ginst15378 (P2_U3160, P2_U3068, P2_U5437);
  and ginst15379 (P2_U3161, P2_U3063, P2_U5437);
  and ginst15380 (P2_U3162, P2_U3077, P2_U5437);
  and ginst15381 (P2_U3163, P2_U3078, P2_U5437);
  and ginst15382 (P2_U3164, P2_U3083, P2_U5437);
  and ginst15383 (P2_U3165, P2_U3084, P2_U5437);
  and ginst15384 (P2_U3166, P2_U3071, P2_U5437);
  and ginst15385 (P2_U3167, P2_U3075, P2_U5437);
  and ginst15386 (P2_U3168, P2_U3076, P2_U5437);
  and ginst15387 (P2_U3169, P2_U3081, P2_U5437);
  and ginst15388 (P2_U3170, P2_U3082, P2_U5437);
  and ginst15389 (P2_U3171, P2_U3074, P2_U5437);
  and ginst15390 (P2_U3172, P2_U3065, P2_U5437);
  and ginst15391 (P2_U3173, P2_U3064, P2_U5437);
  and ginst15392 (P2_U3174, P2_U3085, P2_U5437);
  and ginst15393 (P2_U3175, P2_U3086, P2_U5437);
  and ginst15394 (P2_U3176, P2_U3072, P2_U5437);
  and ginst15395 (P2_U3177, P2_U3073, P2_U5437);
  and ginst15396 (P2_U3178, P2_U3069, P2_U5437);
  and ginst15397 (P2_U3179, P2_U3062, P2_U5437);
  and ginst15398 (P2_U3180, P2_U3066, P2_U5437);
  and ginst15399 (P2_U3181, P2_U3070, P2_U5437);
  and ginst15400 (P2_U3182, P2_U3080, P2_U5437);
  and ginst15401 (P2_U3183, P2_U3079, P2_U5437);
  nand ginst15402 (P2_U3184, P2_U3343, P2_U3404, P2_U5436);
  nand ginst15403 (P2_U3185, P2_U3814, P2_U5430, P2_U5432, P2_U5433);
  nand ginst15404 (P2_U3186, P2_U5420, P2_U5421, P2_U5422, P2_U5423, P2_U5424);
  nand ginst15405 (P2_U3187, P2_U5411, P2_U5412, P2_U5413, P2_U5414, P2_U5415);
  nand ginst15406 (P2_U3188, P2_U5402, P2_U5403, P2_U5404, P2_U5405, P2_U5406);
  nand ginst15407 (P2_U3189, P2_U5393, P2_U5394, P2_U5395, P2_U5396, P2_U5397);
  nand ginst15408 (P2_U3190, P2_U3813, P2_U5385, P2_U5387, P2_U5388);
  nand ginst15409 (P2_U3191, P2_U5375, P2_U5376, P2_U5377, P2_U5378, P2_U5379);
  nand ginst15410 (P2_U3192, P2_U5366, P2_U5367, P2_U5368, P2_U5369, P2_U5370);
  nand ginst15411 (P2_U3193, P2_U3812, P2_U5358, P2_U5360, P2_U5361);
  nand ginst15412 (P2_U3194, P2_U3811, P2_U5349, P2_U5351, P2_U5352);
  nand ginst15413 (P2_U3195, P2_U5339, P2_U5340, P2_U5341, P2_U5342, P2_U5343);
  nand ginst15414 (P2_U3196, P2_U5330, P2_U5331, P2_U5332, P2_U5333, P2_U5334);
  nand ginst15415 (P2_U3197, P2_U5321, P2_U5322, P2_U5323, P2_U5324, P2_U5325);
  nand ginst15416 (P2_U3198, P2_U5312, P2_U5313, P2_U5314, P2_U5315, P2_U5316);
  nand ginst15417 (P2_U3199, P2_U3810, P2_U5304, P2_U5306, P2_U5307);
  nand ginst15418 (P2_U3200, P2_U5294, P2_U5295, P2_U5296, P2_U5297, P2_U5298);
  nand ginst15419 (P2_U3201, P2_U5285, P2_U5286, P2_U5287, P2_U5288, P2_U5289);
  nand ginst15420 (P2_U3202, P2_U3809, P2_U5277, P2_U5279, P2_U5280);
  nand ginst15421 (P2_U3203, P2_U5267, P2_U5268, P2_U5269, P2_U5270, P2_U5271);
  nand ginst15422 (P2_U3204, P2_U3807, P2_U3808, P2_U5260);
  nand ginst15423 (P2_U3205, P2_U5250, P2_U5251, P2_U5252, P2_U5253, P2_U5254);
  nand ginst15424 (P2_U3206, P2_U5241, P2_U5242, P2_U5243, P2_U5244, P2_U5245);
  nand ginst15425 (P2_U3207, P2_U5232, P2_U5233, P2_U5234, P2_U5235, P2_U5236);
  nand ginst15426 (P2_U3208, P2_U5223, P2_U5224, P2_U5225, P2_U5226, P2_U5227);
  nand ginst15427 (P2_U3209, P2_U3805, P2_U5215, P2_U5217, P2_U5218);
  nand ginst15428 (P2_U3210, P2_U5205, P2_U5206, P2_U5207, P2_U5208, P2_U5209);
  nand ginst15429 (P2_U3211, P2_U3804, P2_U5197, P2_U5199, P2_U5200);
  nand ginst15430 (P2_U3212, P2_U5187, P2_U5188, P2_U5189, P2_U5190, P2_U5191);
  nand ginst15431 (P2_U3213, P2_U5174, P2_U5175, P2_U5176, P2_U5177, P2_U5178);
  nand ginst15432 (P2_U3214, P2_U3785, P2_U3786, P2_U5149, P2_U5150);
  nand ginst15433 (P2_U3215, P2_U3783, P2_U3784, P2_U5134, P2_U5135);
  nand ginst15434 (P2_U3216, P2_U3781, P2_U3782, P2_U5119, P2_U5120);
  nand ginst15435 (P2_U3217, P2_U3779, P2_U3780, P2_U5104, P2_U5105);
  nand ginst15436 (P2_U3218, P2_U3777, P2_U3778, P2_U5089, P2_U5090);
  nand ginst15437 (P2_U3219, P2_U3775, P2_U3776, P2_U5074, P2_U5075);
  nand ginst15438 (P2_U3220, P2_U3773, P2_U3774, P2_U5059, P2_U5060);
  nand ginst15439 (P2_U3221, P2_U3771, P2_U3772, P2_U5044, P2_U5045);
  nand ginst15440 (P2_U3222, P2_U3769, P2_U3770, P2_U5029, P2_U5030);
  nand ginst15441 (P2_U3223, P2_U3768, P2_U5014, P2_U5015);
  nand ginst15442 (P2_U3224, P2_U3767, P2_U4999, P2_U5000);
  nand ginst15443 (P2_U3225, P2_U3766, P2_U4984, P2_U4985);
  nand ginst15444 (P2_U3226, P2_U3765, P2_U4969, P2_U4970);
  nand ginst15445 (P2_U3227, P2_U3764, P2_U4954, P2_U4955);
  nand ginst15446 (P2_U3228, P2_U3763, P2_U4939, P2_U4940);
  nand ginst15447 (P2_U3229, P2_U3762, P2_U4924, P2_U4925);
  nand ginst15448 (P2_U3230, P2_U3761, P2_U4909, P2_U4910);
  nand ginst15449 (P2_U3231, P2_U3760, P2_U4894, P2_U4895);
  nand ginst15450 (P2_U3232, P2_U3759, P2_U4879, P2_U4880);
  nand ginst15451 (P2_U3233, P2_U3758, P2_U4864, P2_U4865);
  nand ginst15452 (P2_U3234, P2_U3915, P2_U4852, P2_U4853);
  nand ginst15453 (P2_U3235, P2_U3914, P2_U4850, P2_U4851);
  nand ginst15454 (P2_U3236, P2_U3912, P2_U4846, P2_U4847, P2_U4848, P2_U4849);
  nand ginst15455 (P2_U3237, P2_U3753, P2_U3754, P2_U3911, P2_U4842);
  nand ginst15456 (P2_U3238, P2_U3751, P2_U3752, P2_U3910, P2_U4837);
  nand ginst15457 (P2_U3239, P2_U3749, P2_U3750, P2_U3909, P2_U4832);
  nand ginst15458 (P2_U3240, P2_U3747, P2_U3748, P2_U3908, P2_U4827);
  nand ginst15459 (P2_U3241, P2_U3745, P2_U3746, P2_U3907, P2_U4822);
  nand ginst15460 (P2_U3242, P2_U3743, P2_U3744, P2_U3906, P2_U4817);
  nand ginst15461 (P2_U3243, P2_U3741, P2_U3742, P2_U3905, P2_U4812);
  nand ginst15462 (P2_U3244, P2_U3739, P2_U3740, P2_U3904, P2_U4807);
  nand ginst15463 (P2_U3245, P2_U3737, P2_U3738, P2_U3903, P2_U4802);
  nand ginst15464 (P2_U3246, P2_U3735, P2_U3736, P2_U3902, P2_U4797);
  nand ginst15465 (P2_U3247, P2_U3733, P2_U3734, P2_U3901, P2_U4792);
  nand ginst15466 (P2_U3248, P2_U3731, P2_U3732, P2_U3900, P2_U4787);
  nand ginst15467 (P2_U3249, P2_U3729, P2_U3730, P2_U3899, P2_U4782);
  nand ginst15468 (P2_U3250, P2_U3727, P2_U3728, P2_U3898);
  nand ginst15469 (P2_U3251, P2_U3725, P2_U3726, P2_U3897);
  nand ginst15470 (P2_U3252, P2_U3723, P2_U3724, P2_U3896);
  nand ginst15471 (P2_U3253, P2_U3721, P2_U3722, P2_U3895);
  nand ginst15472 (P2_U3254, P2_U3719, P2_U3720, P2_U3894);
  nand ginst15473 (P2_U3255, P2_U3717, P2_U3718, P2_U3893);
  nand ginst15474 (P2_U3256, P2_U3715, P2_U3716);
  nand ginst15475 (P2_U3257, P2_U3713, P2_U3714);
  nand ginst15476 (P2_U3258, P2_U3711, P2_U3712);
  nand ginst15477 (P2_U3259, P2_U3709, P2_U3710);
  nand ginst15478 (P2_U3260, P2_U3707, P2_U3708);
  nand ginst15479 (P2_U3261, P2_U3705, P2_U3706);
  nand ginst15480 (P2_U3262, P2_U3703, P2_U3704);
  nand ginst15481 (P2_U3263, P2_U3701, P2_U3702);
  nand ginst15482 (P2_U3264, P2_U3699, P2_U3700);
  nand ginst15483 (P2_U3265, P2_U3697, P2_U3698);
  and ginst15484 (P2_U3266, P2_D_REG_31__SCAN_IN, P2_U3880);
  and ginst15485 (P2_U3267, P2_D_REG_30__SCAN_IN, P2_U3880);
  and ginst15486 (P2_U3268, P2_D_REG_29__SCAN_IN, P2_U3880);
  and ginst15487 (P2_U3269, P2_D_REG_28__SCAN_IN, P2_U3880);
  and ginst15488 (P2_U3270, P2_D_REG_27__SCAN_IN, P2_U3880);
  and ginst15489 (P2_U3271, P2_D_REG_26__SCAN_IN, P2_U3880);
  and ginst15490 (P2_U3272, P2_D_REG_25__SCAN_IN, P2_U3880);
  and ginst15491 (P2_U3273, P2_D_REG_24__SCAN_IN, P2_U3880);
  and ginst15492 (P2_U3274, P2_D_REG_23__SCAN_IN, P2_U3880);
  and ginst15493 (P2_U3275, P2_D_REG_22__SCAN_IN, P2_U3880);
  and ginst15494 (P2_U3276, P2_D_REG_21__SCAN_IN, P2_U3880);
  and ginst15495 (P2_U3277, P2_D_REG_20__SCAN_IN, P2_U3880);
  and ginst15496 (P2_U3278, P2_D_REG_19__SCAN_IN, P2_U3880);
  and ginst15497 (P2_U3279, P2_D_REG_18__SCAN_IN, P2_U3880);
  and ginst15498 (P2_U3280, P2_D_REG_17__SCAN_IN, P2_U3880);
  and ginst15499 (P2_U3281, P2_D_REG_16__SCAN_IN, P2_U3880);
  and ginst15500 (P2_U3282, P2_D_REG_15__SCAN_IN, P2_U3880);
  and ginst15501 (P2_U3283, P2_D_REG_14__SCAN_IN, P2_U3880);
  and ginst15502 (P2_U3284, P2_D_REG_13__SCAN_IN, P2_U3880);
  and ginst15503 (P2_U3285, P2_D_REG_12__SCAN_IN, P2_U3880);
  and ginst15504 (P2_U3286, P2_D_REG_11__SCAN_IN, P2_U3880);
  and ginst15505 (P2_U3287, P2_D_REG_10__SCAN_IN, P2_U3880);
  and ginst15506 (P2_U3288, P2_D_REG_9__SCAN_IN, P2_U3880);
  and ginst15507 (P2_U3289, P2_D_REG_8__SCAN_IN, P2_U3880);
  and ginst15508 (P2_U3290, P2_D_REG_7__SCAN_IN, P2_U3880);
  and ginst15509 (P2_U3291, P2_D_REG_6__SCAN_IN, P2_U3880);
  and ginst15510 (P2_U3292, P2_D_REG_5__SCAN_IN, P2_U3880);
  and ginst15511 (P2_U3293, P2_D_REG_4__SCAN_IN, P2_U3880);
  and ginst15512 (P2_U3294, P2_D_REG_3__SCAN_IN, P2_U3880);
  and ginst15513 (P2_U3295, P2_D_REG_2__SCAN_IN, P2_U3880);
  nand ginst15514 (P2_U3296, P2_U4072, P2_U4073, P2_U4074);
  nand ginst15515 (P2_U3297, P2_U4069, P2_U4070, P2_U4071);
  nand ginst15516 (P2_U3298, P2_U4066, P2_U4067, P2_U4068);
  nand ginst15517 (P2_U3299, P2_U4063, P2_U4064, P2_U4065);
  nand ginst15518 (P2_U3300, P2_U4060, P2_U4061, P2_U4062);
  nand ginst15519 (P2_U3301, P2_U4057, P2_U4058, P2_U4059);
  nand ginst15520 (P2_U3302, P2_U4054, P2_U4055, P2_U4056);
  nand ginst15521 (P2_U3303, P2_U4051, P2_U4052, P2_U4053);
  nand ginst15522 (P2_U3304, P2_U4048, P2_U4049, P2_U4050);
  nand ginst15523 (P2_U3305, P2_U4045, P2_U4046, P2_U4047);
  nand ginst15524 (P2_U3306, P2_U4042, P2_U4043, P2_U4044);
  nand ginst15525 (P2_U3307, P2_U4039, P2_U4040, P2_U4041);
  nand ginst15526 (P2_U3308, P2_U4036, P2_U4037, P2_U4038);
  nand ginst15527 (P2_U3309, P2_U4033, P2_U4034, P2_U4035);
  nand ginst15528 (P2_U3310, P2_U4030, P2_U4031, P2_U4032);
  nand ginst15529 (P2_U3311, P2_U4027, P2_U4028, P2_U4029);
  nand ginst15530 (P2_U3312, P2_U4024, P2_U4025, P2_U4026);
  nand ginst15531 (P2_U3313, P2_U4021, P2_U4022, P2_U4023);
  nand ginst15532 (P2_U3314, P2_U4018, P2_U4019, P2_U4020);
  nand ginst15533 (P2_U3315, P2_U4015, P2_U4016, P2_U4017);
  nand ginst15534 (P2_U3316, P2_U4012, P2_U4013, P2_U4014);
  nand ginst15535 (P2_U3317, P2_U4009, P2_U4010, P2_U4011);
  nand ginst15536 (P2_U3318, P2_U4006, P2_U4007, P2_U4008);
  nand ginst15537 (P2_U3319, P2_U4003, P2_U4004, P2_U4005);
  nand ginst15538 (P2_U3320, P2_U4000, P2_U4001, P2_U4002);
  nand ginst15539 (P2_U3321, P2_U3997, P2_U3998, P2_U3999);
  nand ginst15540 (P2_U3322, P2_U3994, P2_U3995, P2_U3996);
  nand ginst15541 (P2_U3323, P2_U3991, P2_U3992, P2_U3993);
  nand ginst15542 (P2_U3324, P2_U3988, P2_U3989, P2_U3990);
  nand ginst15543 (P2_U3325, P2_U3985, P2_U3986, P2_U3987);
  nand ginst15544 (P2_U3326, P2_U3982, P2_U3983, P2_U3984);
  nand ginst15545 (P2_U3327, P2_U3979, P2_U3980, P2_U3981);
  and ginst15546 (P2_U3328, P2_U3797, P2_U5641);
  nand ginst15547 (P2_U3329, P2_STATE_REG_SCAN_IN, P2_U3879);
  not ginst15548 (P2_U3330, U69);
  not ginst15549 (P2_U3331, P2_B_REG_SCAN_IN);
  nand ginst15550 (P2_U3332, P2_U3414, P2_U5649);
  nand ginst15551 (P2_U3333, P2_U3414, P2_U4075);
  nand ginst15552 (P2_U3334, P2_U3420, P2_U3424, P2_U5671);
  nand ginst15553 (P2_U3335, P2_U3418, P2_U3420, P2_U3424);
  nand ginst15554 (P2_U3336, P2_U3049, P2_U3420);
  nand ginst15555 (P2_U3337, P2_U3418, P2_U3419, P2_U3424);
  nand ginst15556 (P2_U3338, P2_U3049, P2_U3419);
  nand ginst15557 (P2_U3339, P2_U3420, P2_U5668, P2_U5674);
  nand ginst15558 (P2_U3340, P2_U5668, P2_U5671);
  nand ginst15559 (P2_U3341, P2_U3419, P2_U3974);
  nand ginst15560 (P2_U3342, P2_U3939, P2_U5665);
  nand ginst15561 (P2_U3343, P2_U5665, P2_U5674);
  nand ginst15562 (P2_U3344, P2_U3419, P2_U3420);
  nand ginst15563 (P2_U3345, P2_U3424, P2_U5665);
  nand ginst15564 (P2_U3346, P2_U3049, P2_U5665);
  nand ginst15565 (P2_U3347, P2_U5683, P2_U5688);
  nand ginst15566 (P2_U3348, P2_U3563, P2_U3564, P2_U4123);
  nand ginst15567 (P2_U3349, P2_U3578, P2_U3580, P2_U4140, P2_U4141);
  nand ginst15568 (P2_U3350, P2_U3582, P2_U3584, P2_U4159, P2_U4160);
  nand ginst15569 (P2_U3351, P2_U3586, P2_U3588, P2_U4178, P2_U4179);
  nand ginst15570 (P2_U3352, P2_U3590, P2_U3592, P2_U4197, P2_U4198);
  nand ginst15571 (P2_U3353, P2_U3594, P2_U3596, P2_U4216, P2_U4217);
  nand ginst15572 (P2_U3354, P2_U3598, P2_U3600, P2_U4235, P2_U4236);
  nand ginst15573 (P2_U3355, P2_U3602, P2_U3604, P2_U4254, P2_U4255);
  nand ginst15574 (P2_U3356, P2_U3606, P2_U3608, P2_U4273, P2_U4274);
  nand ginst15575 (P2_U3357, P2_U3610, P2_U3612, P2_U4292, P2_U4293);
  nand ginst15576 (P2_U3358, P2_U3614, P2_U3616, P2_U4311, P2_U4312);
  nand ginst15577 (P2_U3359, P2_U3618, P2_U3620, P2_U4330, P2_U4331);
  nand ginst15578 (P2_U3360, P2_U3622, P2_U3624, P2_U4349, P2_U4350);
  nand ginst15579 (P2_U3361, P2_U3626, P2_U3628, P2_U4368, P2_U4369);
  nand ginst15580 (P2_U3362, P2_U3630, P2_U3632, P2_U4387, P2_U4388);
  nand ginst15581 (P2_U3363, P2_U3634, P2_U3636, P2_U4406, P2_U4407);
  nand ginst15582 (P2_U3364, P2_U3638, P2_U3640, P2_U4425, P2_U4426);
  nand ginst15583 (P2_U3365, P2_U3642, P2_U3644, P2_U4444, P2_U4445);
  nand ginst15584 (P2_U3366, P2_U3646, P2_U3648, P2_U4463, P2_U4464);
  nand ginst15585 (P2_U3367, P2_U3650, P2_U3652, P2_U4482, P2_U4483);
  nand ginst15586 (P2_U3368, P2_U3347, U81);
  nand ginst15587 (P2_U3369, P2_U3654, P2_U3656, P2_U4501, P2_U4502);
  nand ginst15588 (P2_U3370, P2_U3347, U80);
  nand ginst15589 (P2_U3371, P2_U3658, P2_U3660, P2_U4520, P2_U4521);
  nand ginst15590 (P2_U3372, P2_U3347, U79);
  nand ginst15591 (P2_U3373, P2_U3662, P2_U3664, P2_U4539, P2_U4540);
  nand ginst15592 (P2_U3374, P2_U3347, U78);
  nand ginst15593 (P2_U3375, P2_U3666, P2_U3668, P2_U4558, P2_U4559);
  nand ginst15594 (P2_U3376, P2_U3347, U77);
  nand ginst15595 (P2_U3377, P2_U3670, P2_U3672, P2_U4577, P2_U4578);
  nand ginst15596 (P2_U3378, P2_U3347, U76);
  nand ginst15597 (P2_U3379, P2_U3674, P2_U3676, P2_U4596, P2_U4597);
  nand ginst15598 (P2_U3380, P2_U3347, U75);
  nand ginst15599 (P2_U3381, P2_U3678, P2_U3680, P2_U4615, P2_U4616);
  nand ginst15600 (P2_U3382, P2_U3347, U74);
  nand ginst15601 (P2_U3383, P2_U3682, P2_U3684, P2_U4634, P2_U4635);
  nand ginst15602 (P2_U3384, P2_U3347, U73);
  nand ginst15603 (P2_U3385, P2_U3687, P2_U4653, P2_U4654, P2_U4655, P2_U4656);
  nand ginst15604 (P2_U3386, P2_U3347, U72);
  nand ginst15605 (P2_U3387, P2_U3690, P2_U3692, P2_U4673, P2_U4674, P2_U4675);
  nand ginst15606 (P2_U3388, P2_U3347, U70);
  nand ginst15607 (P2_U3389, P2_U3347, U69);
  nand ginst15608 (P2_U3390, P2_U3424, P2_U3944);
  nand ginst15609 (P2_U3391, P2_U3023, P2_U4698);
  nand ginst15610 (P2_U3392, P2_U3419, P2_U3424, P2_U5671);
  nand ginst15611 (P2_U3393, P2_U3921, P2_U5671);
  nand ginst15612 (P2_U3394, P2_U3944, P2_U5668);
  nand ginst15613 (P2_U3395, P2_U3927, P2_U5671);
  nand ginst15614 (P2_U3396, P2_U3412, P2_U3413, P2_U3414);
  nand ginst15615 (P2_U3397, P2_U3344, P2_U3347);
  nand ginst15616 (P2_U3398, P2_U3934, P2_U4699);
  nand ginst15617 (P2_U3399, P2_U3962, P2_U5658);
  nand ginst15618 (P2_U3400, P2_STATE_REG_SCAN_IN, P2_U3977);
  nand ginst15619 (P2_U3401, P2_U3052, P2_U3756);
  nand ginst15620 (P2_U3402, P2_U3420, P2_U3974);
  nand ginst15621 (P2_U3403, P2_U3015, P2_U3018);
  nand ginst15622 (P2_U3404, P2_U3424, P2_U5674);
  nand ginst15623 (P2_U3405, P2_U3023, P2_U3398);
  nand ginst15624 (P2_U3406, P2_U3016, P2_U3798);
  nand ginst15625 (P2_U3407, P2_STATE_REG_SCAN_IN, P2_U3396, P2_U5168);
  nand ginst15626 (P2_U3408, P2_U3802, P2_U5172);
  not ginst15627 (P2_U3409, P2_R1299_U6);
  nand ginst15628 (P2_U3410, P2_U3938, P2_U5665);
  nand ginst15629 (P2_U3411, P2_U3335, P2_U3336, P2_U3346, P2_U3923);
  nand ginst15630 (P2_U3412, P2_U5644, P2_U5645);
  nand ginst15631 (P2_U3413, P2_U5647, P2_U5648);
  nand ginst15632 (P2_U3414, P2_U5650, P2_U5651);
  nand ginst15633 (P2_U3415, P2_U5656, P2_U5657);
  nand ginst15634 (P2_U3416, P2_U5659, P2_U5660);
  nand ginst15635 (P2_U3417, P2_U5661, P2_U5662);
  nand ginst15636 (P2_U3418, P2_U5669, P2_U5670);
  nand ginst15637 (P2_U3419, P2_U5672, P2_U5673);
  nand ginst15638 (P2_U3420, P2_U5663, P2_U5664);
  nand ginst15639 (P2_U3421, P2_U5675, P2_U5676);
  nand ginst15640 (P2_U3422, P2_U5678, P2_U5679);
  nand ginst15641 (P2_U3423, P2_U5681, P2_U5682);
  nand ginst15642 (P2_U3424, P2_U5666, P2_U5667);
  nand ginst15643 (P2_U3425, P2_U5684, P2_U5685);
  nand ginst15644 (P2_U3426, P2_U5686, P2_U5687);
  nand ginst15645 (P2_U3427, P2_U5689, P2_U5690);
  nand ginst15646 (P2_U3428, P2_U5697, P2_U5698);
  nand ginst15647 (P2_U3429, P2_U5694, P2_U5695);
  nand ginst15648 (P2_U3430, P2_U5700, P2_U5701);
  nand ginst15649 (P2_U3431, P2_U5702, P2_U5703);
  nand ginst15650 (P2_U3432, P2_U5704, P2_U5705);
  nand ginst15651 (P2_U3433, P2_U5707, P2_U5708);
  nand ginst15652 (P2_U3434, P2_U5709, P2_U5710);
  nand ginst15653 (P2_U3435, P2_U5711, P2_U5712);
  nand ginst15654 (P2_U3436, P2_U5714, P2_U5715);
  nand ginst15655 (P2_U3437, P2_U5716, P2_U5717);
  nand ginst15656 (P2_U3438, P2_U5718, P2_U5719);
  nand ginst15657 (P2_U3439, P2_U5721, P2_U5722);
  nand ginst15658 (P2_U3440, P2_U5723, P2_U5724);
  nand ginst15659 (P2_U3441, P2_U5725, P2_U5726);
  nand ginst15660 (P2_U3442, P2_U5728, P2_U5729);
  nand ginst15661 (P2_U3443, P2_U5730, P2_U5731);
  nand ginst15662 (P2_U3444, P2_U5732, P2_U5733);
  nand ginst15663 (P2_U3445, P2_U5735, P2_U5736);
  nand ginst15664 (P2_U3446, P2_U5737, P2_U5738);
  nand ginst15665 (P2_U3447, P2_U5739, P2_U5740);
  nand ginst15666 (P2_U3448, P2_U5742, P2_U5743);
  nand ginst15667 (P2_U3449, P2_U5744, P2_U5745);
  nand ginst15668 (P2_U3450, P2_U5746, P2_U5747);
  nand ginst15669 (P2_U3451, P2_U5749, P2_U5750);
  nand ginst15670 (P2_U3452, P2_U5751, P2_U5752);
  nand ginst15671 (P2_U3453, P2_U5753, P2_U5754);
  nand ginst15672 (P2_U3454, P2_U5756, P2_U5757);
  nand ginst15673 (P2_U3455, P2_U5758, P2_U5759);
  nand ginst15674 (P2_U3456, P2_U5760, P2_U5761);
  nand ginst15675 (P2_U3457, P2_U5763, P2_U5764);
  nand ginst15676 (P2_U3458, P2_U5765, P2_U5766);
  nand ginst15677 (P2_U3459, P2_U5767, P2_U5768);
  nand ginst15678 (P2_U3460, P2_U5770, P2_U5771);
  nand ginst15679 (P2_U3461, P2_U5772, P2_U5773);
  nand ginst15680 (P2_U3462, P2_U5774, P2_U5775);
  nand ginst15681 (P2_U3463, P2_U5777, P2_U5778);
  nand ginst15682 (P2_U3464, P2_U5779, P2_U5780);
  nand ginst15683 (P2_U3465, P2_U5781, P2_U5782);
  nand ginst15684 (P2_U3466, P2_U5784, P2_U5785);
  nand ginst15685 (P2_U3467, P2_U5786, P2_U5787);
  nand ginst15686 (P2_U3468, P2_U5788, P2_U5789);
  nand ginst15687 (P2_U3469, P2_U5791, P2_U5792);
  nand ginst15688 (P2_U3470, P2_U5793, P2_U5794);
  nand ginst15689 (P2_U3471, P2_U5795, P2_U5796);
  nand ginst15690 (P2_U3472, P2_U5798, P2_U5799);
  nand ginst15691 (P2_U3473, P2_U5800, P2_U5801);
  nand ginst15692 (P2_U3474, P2_U5802, P2_U5803);
  nand ginst15693 (P2_U3475, P2_U5805, P2_U5806);
  nand ginst15694 (P2_U3476, P2_U5807, P2_U5808);
  nand ginst15695 (P2_U3477, P2_U5809, P2_U5810);
  nand ginst15696 (P2_U3478, P2_U5812, P2_U5813);
  nand ginst15697 (P2_U3479, P2_U5814, P2_U5815);
  nand ginst15698 (P2_U3480, P2_U5816, P2_U5817);
  nand ginst15699 (P2_U3481, P2_U5819, P2_U5820);
  nand ginst15700 (P2_U3482, P2_U5821, P2_U5822);
  nand ginst15701 (P2_U3483, P2_U5823, P2_U5824);
  nand ginst15702 (P2_U3484, P2_U5826, P2_U5827);
  nand ginst15703 (P2_U3485, P2_U5828, P2_U5829);
  nand ginst15704 (P2_U3486, P2_U5831, P2_U5832);
  nand ginst15705 (P2_U3487, P2_U5833, P2_U5834);
  nand ginst15706 (P2_U3488, P2_U5835, P2_U5836);
  nand ginst15707 (P2_U3489, P2_U5837, P2_U5838);
  nand ginst15708 (P2_U3490, P2_U5839, P2_U5840);
  nand ginst15709 (P2_U3491, P2_U5841, P2_U5842);
  nand ginst15710 (P2_U3492, P2_U5843, P2_U5844);
  nand ginst15711 (P2_U3493, P2_U5845, P2_U5846);
  nand ginst15712 (P2_U3494, P2_U5847, P2_U5848);
  nand ginst15713 (P2_U3495, P2_U5849, P2_U5850);
  nand ginst15714 (P2_U3496, P2_U5851, P2_U5852);
  nand ginst15715 (P2_U3497, P2_U5853, P2_U5854);
  nand ginst15716 (P2_U3498, P2_U5855, P2_U5856);
  nand ginst15717 (P2_U3499, P2_U5857, P2_U5858);
  nand ginst15718 (P2_U3500, P2_U5859, P2_U5860);
  nand ginst15719 (P2_U3501, P2_U5861, P2_U5862);
  nand ginst15720 (P2_U3502, P2_U5863, P2_U5864);
  nand ginst15721 (P2_U3503, P2_U5865, P2_U5866);
  nand ginst15722 (P2_U3504, P2_U5867, P2_U5868);
  nand ginst15723 (P2_U3505, P2_U5869, P2_U5870);
  nand ginst15724 (P2_U3506, P2_U5871, P2_U5872);
  nand ginst15725 (P2_U3507, P2_U5873, P2_U5874);
  nand ginst15726 (P2_U3508, P2_U5875, P2_U5876);
  nand ginst15727 (P2_U3509, P2_U5877, P2_U5878);
  nand ginst15728 (P2_U3510, P2_U5879, P2_U5880);
  nand ginst15729 (P2_U3511, P2_U5881, P2_U5882);
  nand ginst15730 (P2_U3512, P2_U5883, P2_U5884);
  nand ginst15731 (P2_U3513, P2_U5885, P2_U5886);
  nand ginst15732 (P2_U3514, P2_U5887, P2_U5888);
  nand ginst15733 (P2_U3515, P2_U5889, P2_U5890);
  nand ginst15734 (P2_U3516, P2_U5891, P2_U5892);
  nand ginst15735 (P2_U3517, P2_U5893, P2_U5894);
  nand ginst15736 (P2_U3518, P2_U5895, P2_U5896);
  nand ginst15737 (P2_U3519, P2_U5897, P2_U5898);
  xor ginst15738 (P2_U3520, P2_U3520_in, flip_signal);
  nand ginst15739 (P2_U3520_in, P2_U5899, P2_U5900);
  nand ginst15740 (P2_U3521, P2_U5901, P2_U5902);
  nand ginst15741 (P2_U3522, P2_U5903, P2_U5904);
  nand ginst15742 (P2_U3523, P2_U5905, P2_U5906);
  nand ginst15743 (P2_U3524, P2_U5907, P2_U5908);
  nand ginst15744 (P2_U3525, P2_U5909, P2_U5910);
  nand ginst15745 (P2_U3526, P2_U5911, P2_U5912);
  nand ginst15746 (P2_U3527, P2_U5913, P2_U5914);
  nand ginst15747 (P2_U3528, P2_U5915, P2_U5916);
  nand ginst15748 (P2_U3529, P2_U5917, P2_U5918);
  nand ginst15749 (P2_U3530, P2_U5919, P2_U5920);
  nand ginst15750 (P2_U3531, P2_U5985, P2_U5986);
  nand ginst15751 (P2_U3532, P2_U5987, P2_U5988);
  nand ginst15752 (P2_U3533, P2_U5989, P2_U5990);
  nand ginst15753 (P2_U3534, P2_U5991, P2_U5992);
  nand ginst15754 (P2_U3535, P2_U5993, P2_U5994);
  nand ginst15755 (P2_U3536, P2_U5995, P2_U5996);
  nand ginst15756 (P2_U3537, P2_U5997, P2_U5998);
  nand ginst15757 (P2_U3538, P2_U5999, P2_U6000);
  nand ginst15758 (P2_U3539, P2_U6001, P2_U6002);
  nand ginst15759 (P2_U3540, P2_U6003, P2_U6004);
  nand ginst15760 (P2_U3541, P2_U6005, P2_U6006);
  nand ginst15761 (P2_U3542, P2_U6007, P2_U6008);
  nand ginst15762 (P2_U3543, P2_U6009, P2_U6010);
  nand ginst15763 (P2_U3544, P2_U6011, P2_U6012);
  nand ginst15764 (P2_U3545, P2_U6013, P2_U6014);
  nand ginst15765 (P2_U3546, P2_U6015, P2_U6016);
  nand ginst15766 (P2_U3547, P2_U6017, P2_U6018);
  nand ginst15767 (P2_U3548, P2_U6019, P2_U6020);
  nand ginst15768 (P2_U3549, P2_U6021, P2_U6022);
  nand ginst15769 (P2_U3550, P2_U6023, P2_U6024);
  nand ginst15770 (P2_U3551, P2_U6025, P2_U6026);
  nand ginst15771 (P2_U3552, P2_U6027, P2_U6028);
  nand ginst15772 (P2_U3553, P2_U6029, P2_U6030);
  nand ginst15773 (P2_U3554, P2_U6031, P2_U6032);
  nand ginst15774 (P2_U3555, P2_U6033, P2_U6034);
  nand ginst15775 (P2_U3556, P2_U6035, P2_U6036);
  nand ginst15776 (P2_U3557, P2_U6037, P2_U6038);
  nand ginst15777 (P2_U3558, P2_U6039, P2_U6040);
  nand ginst15778 (P2_U3559, P2_U6041, P2_U6042);
  nand ginst15779 (P2_U3560, P2_U6043, P2_U6044);
  nand ginst15780 (P2_U3561, P2_U6045, P2_U6046);
  nand ginst15781 (P2_U3562, P2_U6047, P2_U6048);
  and ginst15782 (P2_U3563, P2_U4117, P2_U4118, P2_U4119, P2_U4120);
  and ginst15783 (P2_U3564, P2_U4121, P2_U4122);
  and ginst15784 (P2_U3565, P2_U4125, P2_U4127);
  and ginst15785 (P2_U3566, P2_U4079, P2_U4080, P2_U4081, P2_U4082);
  and ginst15786 (P2_U3567, P2_U4083, P2_U4084, P2_U4085, P2_U4086);
  and ginst15787 (P2_U3568, P2_U4087, P2_U4088, P2_U4089, P2_U4090);
  and ginst15788 (P2_U3569, P2_U4091, P2_U4092, P2_U4093);
  and ginst15789 (P2_U3570, P2_U3566, P2_U3567, P2_U3568, P2_U3569);
  and ginst15790 (P2_U3571, P2_U4094, P2_U4095, P2_U4096, P2_U4097);
  and ginst15791 (P2_U3572, P2_U4098, P2_U4099, P2_U4100, P2_U4101);
  and ginst15792 (P2_U3573, P2_U4102, P2_U4103, P2_U4104, P2_U4105);
  and ginst15793 (P2_U3574, P2_U4106, P2_U4107, P2_U4108);
  and ginst15794 (P2_U3575, P2_U3571, P2_U3572, P2_U3573, P2_U3574);
  and ginst15795 (P2_U3576, P2_U4110, P2_U5696);
  and ginst15796 (P2_U3577, P2_U3023, P2_U5699);
  and ginst15797 (P2_U3578, P2_U4142, P2_U4143);
  and ginst15798 (P2_U3579, P2_U4144, P2_U4145);
  and ginst15799 (P2_U3580, P2_U3579, P2_U4146, P2_U4147);
  and ginst15800 (P2_U3581, P2_U4149, P2_U4150, P2_U4151, P2_U4152);
  and ginst15801 (P2_U3582, P2_U4161, P2_U4162);
  and ginst15802 (P2_U3583, P2_U4163, P2_U4164);
  and ginst15803 (P2_U3584, P2_U3583, P2_U4165, P2_U4166);
  and ginst15804 (P2_U3585, P2_U4168, P2_U4169, P2_U4170, P2_U4171);
  and ginst15805 (P2_U3586, P2_U4180, P2_U4181);
  and ginst15806 (P2_U3587, P2_U4182, P2_U4183);
  and ginst15807 (P2_U3588, P2_U3587, P2_U4184, P2_U4185);
  and ginst15808 (P2_U3589, P2_U4187, P2_U4188, P2_U4189, P2_U4190);
  and ginst15809 (P2_U3590, P2_U4199, P2_U4200);
  and ginst15810 (P2_U3591, P2_U4201, P2_U4202);
  and ginst15811 (P2_U3592, P2_U3591, P2_U4203, P2_U4204);
  and ginst15812 (P2_U3593, P2_U4206, P2_U4207, P2_U4208, P2_U4209);
  and ginst15813 (P2_U3594, P2_U4218, P2_U4219);
  and ginst15814 (P2_U3595, P2_U4220, P2_U4221);
  and ginst15815 (P2_U3596, P2_U3595, P2_U4222, P2_U4223);
  and ginst15816 (P2_U3597, P2_U4225, P2_U4226, P2_U4227, P2_U4228);
  and ginst15817 (P2_U3598, P2_U4237, P2_U4238);
  and ginst15818 (P2_U3599, P2_U4239, P2_U4240);
  and ginst15819 (P2_U3600, P2_U3599, P2_U4241, P2_U4242);
  and ginst15820 (P2_U3601, P2_U4244, P2_U4245, P2_U4246, P2_U4247);
  and ginst15821 (P2_U3602, P2_U4256, P2_U4257);
  and ginst15822 (P2_U3603, P2_U4258, P2_U4259);
  and ginst15823 (P2_U3604, P2_U3603, P2_U4260, P2_U4261);
  and ginst15824 (P2_U3605, P2_U4263, P2_U4264, P2_U4265, P2_U4266);
  and ginst15825 (P2_U3606, P2_U4275, P2_U4276);
  and ginst15826 (P2_U3607, P2_U4277, P2_U4278);
  and ginst15827 (P2_U3608, P2_U3607, P2_U4279, P2_U4280);
  and ginst15828 (P2_U3609, P2_U4282, P2_U4283, P2_U4284, P2_U4285);
  and ginst15829 (P2_U3610, P2_U4294, P2_U4295);
  and ginst15830 (P2_U3611, P2_U4296, P2_U4297);
  and ginst15831 (P2_U3612, P2_U3611, P2_U4298, P2_U4299);
  and ginst15832 (P2_U3613, P2_U4301, P2_U4302, P2_U4303, P2_U4304);
  and ginst15833 (P2_U3614, P2_U4313, P2_U4314);
  and ginst15834 (P2_U3615, P2_U4315, P2_U4316);
  and ginst15835 (P2_U3616, P2_U3615, P2_U4317, P2_U4318);
  and ginst15836 (P2_U3617, P2_U4320, P2_U4321, P2_U4322, P2_U4323);
  and ginst15837 (P2_U3618, P2_U4332, P2_U4333);
  and ginst15838 (P2_U3619, P2_U4334, P2_U4335);
  and ginst15839 (P2_U3620, P2_U3619, P2_U4336, P2_U4337);
  and ginst15840 (P2_U3621, P2_U4339, P2_U4340, P2_U4341, P2_U4342);
  and ginst15841 (P2_U3622, P2_U4351, P2_U4352);
  and ginst15842 (P2_U3623, P2_U4353, P2_U4354);
  and ginst15843 (P2_U3624, P2_U3623, P2_U4355, P2_U4356);
  and ginst15844 (P2_U3625, P2_U4358, P2_U4359, P2_U4360, P2_U4361);
  and ginst15845 (P2_U3626, P2_U4370, P2_U4371);
  and ginst15846 (P2_U3627, P2_U4372, P2_U4373);
  and ginst15847 (P2_U3628, P2_U3627, P2_U4374, P2_U4375);
  and ginst15848 (P2_U3629, P2_U4377, P2_U4378, P2_U4379, P2_U4380);
  and ginst15849 (P2_U3630, P2_U4389, P2_U4390);
  and ginst15850 (P2_U3631, P2_U4391, P2_U4392);
  and ginst15851 (P2_U3632, P2_U3631, P2_U4393, P2_U4394);
  and ginst15852 (P2_U3633, P2_U4396, P2_U4397, P2_U4398, P2_U4399);
  and ginst15853 (P2_U3634, P2_U4408, P2_U4409);
  and ginst15854 (P2_U3635, P2_U4410, P2_U4411);
  and ginst15855 (P2_U3636, P2_U3635, P2_U4412, P2_U4413);
  and ginst15856 (P2_U3637, P2_U4415, P2_U4416, P2_U4417, P2_U4418);
  and ginst15857 (P2_U3638, P2_U4427, P2_U4428);
  and ginst15858 (P2_U3639, P2_U4429, P2_U4430);
  and ginst15859 (P2_U3640, P2_U3639, P2_U4431, P2_U4432);
  and ginst15860 (P2_U3641, P2_U4434, P2_U4435, P2_U4436, P2_U4437);
  and ginst15861 (P2_U3642, P2_U4446, P2_U4447);
  and ginst15862 (P2_U3643, P2_U4448, P2_U4449);
  and ginst15863 (P2_U3644, P2_U3643, P2_U4450, P2_U4451);
  and ginst15864 (P2_U3645, P2_U4453, P2_U4454, P2_U4455, P2_U4456);
  and ginst15865 (P2_U3646, P2_U4465, P2_U4466);
  and ginst15866 (P2_U3647, P2_U4467, P2_U4468);
  and ginst15867 (P2_U3648, P2_U3647, P2_U4469, P2_U4470);
  and ginst15868 (P2_U3649, P2_U4472, P2_U4473, P2_U4474, P2_U4475);
  and ginst15869 (P2_U3650, P2_U4484, P2_U4485);
  and ginst15870 (P2_U3651, P2_U4486, P2_U4487);
  and ginst15871 (P2_U3652, P2_U3651, P2_U4488, P2_U4489);
  and ginst15872 (P2_U3653, P2_U4491, P2_U4492, P2_U4493, P2_U4494);
  and ginst15873 (P2_U3654, P2_U4503, P2_U4504);
  and ginst15874 (P2_U3655, P2_U4505, P2_U4506);
  and ginst15875 (P2_U3656, P2_U3655, P2_U4507, P2_U4508);
  and ginst15876 (P2_U3657, P2_U4510, P2_U4511, P2_U4512, P2_U4513);
  and ginst15877 (P2_U3658, P2_U4522, P2_U4523);
  and ginst15878 (P2_U3659, P2_U4524, P2_U4525);
  and ginst15879 (P2_U3660, P2_U3659, P2_U4526, P2_U4527);
  and ginst15880 (P2_U3661, P2_U4529, P2_U4530, P2_U4531, P2_U4532);
  and ginst15881 (P2_U3662, P2_U4541, P2_U4542);
  and ginst15882 (P2_U3663, P2_U4543, P2_U4544);
  and ginst15883 (P2_U3664, P2_U3663, P2_U4545, P2_U4546);
  and ginst15884 (P2_U3665, P2_U4548, P2_U4549, P2_U4550, P2_U4551);
  and ginst15885 (P2_U3666, P2_U4560, P2_U4561);
  and ginst15886 (P2_U3667, P2_U4562, P2_U4563);
  and ginst15887 (P2_U3668, P2_U3667, P2_U4564, P2_U4565);
  and ginst15888 (P2_U3669, P2_U4567, P2_U4568, P2_U4569, P2_U4570);
  and ginst15889 (P2_U3670, P2_U4579, P2_U4580);
  and ginst15890 (P2_U3671, P2_U4581, P2_U4582);
  and ginst15891 (P2_U3672, P2_U3671, P2_U4583, P2_U4584);
  and ginst15892 (P2_U3673, P2_U4586, P2_U4587, P2_U4588, P2_U4589);
  and ginst15893 (P2_U3674, P2_U4598, P2_U4599);
  and ginst15894 (P2_U3675, P2_U4600, P2_U4601);
  and ginst15895 (P2_U3676, P2_U3675, P2_U4602, P2_U4603);
  and ginst15896 (P2_U3677, P2_U4605, P2_U4606, P2_U4607, P2_U4608);
  and ginst15897 (P2_U3678, P2_U4617, P2_U4618);
  and ginst15898 (P2_U3679, P2_U4619, P2_U4620);
  and ginst15899 (P2_U3680, P2_U3679, P2_U4621, P2_U4622);
  and ginst15900 (P2_U3681, P2_U4624, P2_U4625, P2_U4626, P2_U4627);
  and ginst15901 (P2_U3682, P2_U4636, P2_U4637);
  and ginst15902 (P2_U3683, P2_U4638, P2_U4639);
  and ginst15903 (P2_U3684, P2_U3683, P2_U4640, P2_U4641);
  and ginst15904 (P2_U3685, P2_U4643, P2_U4644, P2_U4645, P2_U4646);
  and ginst15905 (P2_U3686, P2_U4657, P2_U4658);
  and ginst15906 (P2_U3687, P2_U3686, P2_U4659, P2_U4660);
  and ginst15907 (P2_U3688, P2_U4662, P2_U4663, P2_U4664, P2_U4665);
  and ginst15908 (P2_U3689, P2_U3963, P2_U4672);
  and ginst15909 (P2_U3690, P2_U4676, P2_U4677);
  and ginst15910 (P2_U3691, P2_U4678, P2_U4679);
  and ginst15911 (P2_U3692, P2_U3691, P2_U4680, P2_U4681);
  and ginst15912 (P2_U3693, P2_U4683, P2_U4684, P2_U4685);
  and ginst15913 (P2_U3694, P2_U3963, P2_U4672);
  and ginst15914 (P2_U3695, P2_U3023, P2_U3428);
  and ginst15915 (P2_U3696, P2_U3429, P2_U3935, P2_U5699);
  and ginst15916 (P2_U3697, P2_U4701, P2_U4702, P2_U4703);
  and ginst15917 (P2_U3698, P2_U3883, P2_U4704, P2_U4705);
  and ginst15918 (P2_U3699, P2_U4706, P2_U4707, P2_U4708);
  and ginst15919 (P2_U3700, P2_U3884, P2_U4709, P2_U4710);
  and ginst15920 (P2_U3701, P2_U4711, P2_U4712, P2_U4713);
  and ginst15921 (P2_U3702, P2_U3885, P2_U4714, P2_U4715);
  and ginst15922 (P2_U3703, P2_U4716, P2_U4717, P2_U4718);
  and ginst15923 (P2_U3704, P2_U3886, P2_U4719, P2_U4720);
  and ginst15924 (P2_U3705, P2_U4721, P2_U4722, P2_U4723);
  and ginst15925 (P2_U3706, P2_U3887, P2_U4724, P2_U4725);
  and ginst15926 (P2_U3707, P2_U4726, P2_U4727, P2_U4728);
  and ginst15927 (P2_U3708, P2_U3888, P2_U4729, P2_U4730);
  and ginst15928 (P2_U3709, P2_U4731, P2_U4732, P2_U4733);
  and ginst15929 (P2_U3710, P2_U3889, P2_U4734, P2_U4735);
  and ginst15930 (P2_U3711, P2_U4736, P2_U4737, P2_U4738);
  and ginst15931 (P2_U3712, P2_U3890, P2_U4739, P2_U4740);
  and ginst15932 (P2_U3713, P2_U4741, P2_U4742, P2_U4743);
  and ginst15933 (P2_U3714, P2_U3891, P2_U4744, P2_U4745);
  and ginst15934 (P2_U3715, P2_U4746, P2_U4747, P2_U4748);
  and ginst15935 (P2_U3716, P2_U3892, P2_U4749, P2_U4750);
  and ginst15936 (P2_U3717, P2_U4751, P2_U4752, P2_U4753);
  and ginst15937 (P2_U3718, P2_U4754, P2_U4755);
  and ginst15938 (P2_U3719, P2_U4756, P2_U4757, P2_U4758);
  and ginst15939 (P2_U3720, P2_U4759, P2_U4760);
  and ginst15940 (P2_U3721, P2_U4761, P2_U4762, P2_U4763);
  and ginst15941 (P2_U3722, P2_U4764, P2_U4765);
  and ginst15942 (P2_U3723, P2_U4766, P2_U4767, P2_U4768);
  and ginst15943 (P2_U3724, P2_U4769, P2_U4770);
  and ginst15944 (P2_U3725, P2_U4771, P2_U4772, P2_U4773);
  and ginst15945 (P2_U3726, P2_U4774, P2_U4775);
  and ginst15946 (P2_U3727, P2_U4776, P2_U4777, P2_U4778);
  and ginst15947 (P2_U3728, P2_U4779, P2_U4780);
  and ginst15948 (P2_U3729, P2_U4781, P2_U4783);
  and ginst15949 (P2_U3730, P2_U4784, P2_U4785);
  and ginst15950 (P2_U3731, P2_U4786, P2_U4788);
  and ginst15951 (P2_U3732, P2_U4789, P2_U4790);
  and ginst15952 (P2_U3733, P2_U4791, P2_U4793);
  and ginst15953 (P2_U3734, P2_U4794, P2_U4795);
  and ginst15954 (P2_U3735, P2_U4796, P2_U4798);
  and ginst15955 (P2_U3736, P2_U4799, P2_U4800);
  and ginst15956 (P2_U3737, P2_U4801, P2_U4803);
  and ginst15957 (P2_U3738, P2_U4804, P2_U4805);
  and ginst15958 (P2_U3739, P2_U4806, P2_U4808);
  and ginst15959 (P2_U3740, P2_U4809, P2_U4810);
  and ginst15960 (P2_U3741, P2_U4811, P2_U4813);
  and ginst15961 (P2_U3742, P2_U4814, P2_U4815);
  and ginst15962 (P2_U3743, P2_U4816, P2_U4818);
  and ginst15963 (P2_U3744, P2_U4819, P2_U4820);
  and ginst15964 (P2_U3745, P2_U4821, P2_U4823);
  and ginst15965 (P2_U3746, P2_U4824, P2_U4825);
  and ginst15966 (P2_U3747, P2_U4826, P2_U4828);
  and ginst15967 (P2_U3748, P2_U4829, P2_U4830);
  and ginst15968 (P2_U3749, P2_U4831, P2_U4833);
  and ginst15969 (P2_U3750, P2_U4834, P2_U4835);
  and ginst15970 (P2_U3751, P2_U4836, P2_U4838);
  and ginst15971 (P2_U3752, P2_U4839, P2_U4840);
  and ginst15972 (P2_U3753, P2_U4841, P2_U4843);
  and ginst15973 (P2_U3754, P2_U4844, P2_U4845);
  and ginst15974 (P2_U3755, P2_U3334, P2_U3335, P2_U3336);
  and ginst15975 (P2_U3756, P2_U3397, P2_U5643);
  and ginst15976 (P2_U3757, P2_STATE_REG_SCAN_IN, P2_U3415);
  and ginst15977 (P2_U3758, P2_U4866, P2_U4867, P2_U4868, P2_U4869, P2_U4870);
  and ginst15978 (P2_U3759, P2_U4881, P2_U4882, P2_U4883, P2_U4884, P2_U4885);
  and ginst15979 (P2_U3760, P2_U4896, P2_U4897, P2_U4898, P2_U4899, P2_U4900);
  and ginst15980 (P2_U3761, P2_U4911, P2_U4912, P2_U4913, P2_U4914, P2_U4915);
  and ginst15981 (P2_U3762, P2_U4926, P2_U4927, P2_U4928, P2_U4929, P2_U4930);
  and ginst15982 (P2_U3763, P2_U4941, P2_U4942, P2_U4943, P2_U4944, P2_U4945);
  and ginst15983 (P2_U3764, P2_U4956, P2_U4957, P2_U4958, P2_U4959, P2_U4960);
  and ginst15984 (P2_U3765, P2_U4971, P2_U4972, P2_U4973, P2_U4974, P2_U4975);
  and ginst15985 (P2_U3766, P2_U4986, P2_U4987, P2_U4988, P2_U4989, P2_U4990);
  and ginst15986 (P2_U3767, P2_U5001, P2_U5002, P2_U5003, P2_U5004, P2_U5005);
  and ginst15987 (P2_U3768, P2_U5016, P2_U5017, P2_U5018, P2_U5019, P2_U5020);
  and ginst15988 (P2_U3769, P2_U5031, P2_U5032);
  and ginst15989 (P2_U3770, P2_U5033, P2_U5034, P2_U5035);
  and ginst15990 (P2_U3771, P2_U5046, P2_U5047);
  and ginst15991 (P2_U3772, P2_U5048, P2_U5049, P2_U5050);
  and ginst15992 (P2_U3773, P2_U5061, P2_U5062);
  and ginst15993 (P2_U3774, P2_U5063, P2_U5064, P2_U5065);
  and ginst15994 (P2_U3775, P2_U5076, P2_U5077);
  and ginst15995 (P2_U3776, P2_U5078, P2_U5079, P2_U5080);
  and ginst15996 (P2_U3777, P2_U5091, P2_U5092);
  and ginst15997 (P2_U3778, P2_U5093, P2_U5094, P2_U5095);
  and ginst15998 (P2_U3779, P2_U5106, P2_U5107);
  and ginst15999 (P2_U3780, P2_U5108, P2_U5109, P2_U5110);
  and ginst16000 (P2_U3781, P2_U5121, P2_U5122);
  and ginst16001 (P2_U3782, P2_U5123, P2_U5124, P2_U5125);
  and ginst16002 (P2_U3783, P2_U5136, P2_U5137);
  and ginst16003 (P2_U3784, P2_U5138, P2_U5139, P2_U5140);
  and ginst16004 (P2_U3785, P2_U5151, P2_U5152);
  and ginst16005 (P2_U3786, P2_U5153, P2_U5154, P2_U5155);
  and ginst16006 (P2_U3787, P2_U5639, P2_U5658);
  and ginst16007 (P2_U3788, P2_U6100, P2_U6103, P2_U6106);
  and ginst16008 (P2_U3789, P2_U6088, P2_U6091, P2_U6094, P2_U6097);
  and ginst16009 (P2_U3790, P2_U6112, P2_U6115, P2_U6118, P2_U6121);
  and ginst16010 (P2_U3791, P2_U6124, P2_U6127, P2_U6130, P2_U6133);
  and ginst16011 (P2_U3792, P2_U3788, P2_U3789, P2_U3790, P2_U3791, P2_U6109);
  and ginst16012 (P2_U3793, P2_U3795, P2_U3796, P2_U6055, P2_U6058, P2_U6061);
  and ginst16013 (P2_U3794, P2_U6136, P2_U6139, P2_U6142, P2_U6145, P2_U6148);
  and ginst16014 (P2_U3795, P2_U6064, P2_U6067, P2_U6070, P2_U6073);
  and ginst16015 (P2_U3796, P2_U6076, P2_U6079);
  and ginst16016 (P2_U3797, P2_U5631, P2_U5640);
  and ginst16017 (P2_U3798, P2_U3428, P2_U3429);
  and ginst16018 (P2_U3799, P2_U3339, P2_U3928);
  and ginst16019 (P2_U3800, P2_U3342, P2_U3799);
  and ginst16020 (P2_U3801, P2_U3395, P2_U3410);
  and ginst16021 (P2_U3802, P2_U3399, P2_U3935, P2_U5658);
  and ginst16022 (P2_U3803, P2_U3023, P2_U5171);
  and ginst16023 (P2_U3804, P2_U5196, P2_U5198);
  and ginst16024 (P2_U3805, P2_U5214, P2_U5216);
  and ginst16025 (P2_U3806, P2_U3080, P2_U3969);
  and ginst16026 (P2_U3807, P2_U5258, P2_U5259);
  and ginst16027 (P2_U3808, P2_U5261, P2_U5262);
  and ginst16028 (P2_U3809, P2_U5276, P2_U5278);
  and ginst16029 (P2_U3810, P2_U5303, P2_U5305);
  and ginst16030 (P2_U3811, P2_U5348, P2_U5350);
  and ginst16031 (P2_U3812, P2_U5357, P2_U5359);
  and ginst16032 (P2_U3813, P2_U5384, P2_U5386);
  and ginst16033 (P2_U3814, P2_U5429, P2_U5431);
  and ginst16034 (P2_U3815, P2_STATE_REG_SCAN_IN, P2_U5435);
  and ginst16035 (P2_U3816, P2_U3919, P2_U3920, P2_U3936);
  and ginst16036 (P2_U3817, P2_U3419, P2_U5671);
  and ginst16037 (P2_U3818, P2_U3339, P2_U3394);
  and ginst16038 (P2_U3819, P2_U3342, P2_U3390, P2_U3818);
  and ginst16039 (P2_U3820, P2_U3334, P2_U3928);
  and ginst16040 (P2_U3821, P2_U3415, P2_U5444);
  and ginst16041 (P2_U3822, P2_U3415, P2_U5447);
  and ginst16042 (P2_U3823, P2_U3415, P2_U5450);
  and ginst16043 (P2_U3824, P2_U3415, P2_U5453);
  and ginst16044 (P2_U3825, P2_U3415, P2_U5456);
  and ginst16045 (P2_U3826, P2_U3827, P2_U5457);
  and ginst16046 (P2_U3827, P2_U3415, P2_U5459);
  and ginst16047 (P2_U3828, P2_U3410, P2_U5460);
  and ginst16048 (P2_U3829, P2_U3830, P2_U5465);
  and ginst16049 (P2_U3830, P2_U3415, P2_U5467);
  and ginst16050 (P2_U3831, P2_U3415, P2_U5468);
  and ginst16051 (P2_U3832, P2_U3415, P2_U5471);
  and ginst16052 (P2_U3833, P2_U3415, P2_U5474);
  and ginst16053 (P2_U3834, P2_U3415, P2_U5477);
  and ginst16054 (P2_U3835, P2_U3415, P2_U5480);
  and ginst16055 (P2_U3836, P2_U3415, P2_U5483);
  and ginst16056 (P2_U3837, P2_U3415, P2_U5486);
  and ginst16057 (P2_U3838, P2_U3415, P2_U5489);
  and ginst16058 (P2_U3839, P2_U3415, P2_U5492);
  and ginst16059 (P2_U3840, P2_U3415, P2_U5495);
  and ginst16060 (P2_U3841, P2_U3842, P2_U5498);
  and ginst16061 (P2_U3842, P2_U3415, P2_U5500);
  and ginst16062 (P2_U3843, P2_U3415, P2_U5501);
  and ginst16063 (P2_U3844, P2_U3415, P2_U5504);
  and ginst16064 (P2_U3845, P2_U3415, P2_U5507);
  and ginst16065 (P2_U3846, P2_U3415, P2_U5510);
  and ginst16066 (P2_U3847, P2_U3415, P2_U5513);
  and ginst16067 (P2_U3848, P2_U3415, P2_U5516);
  and ginst16068 (P2_U3849, P2_U3415, P2_U5519);
  and ginst16069 (P2_U3850, P2_U3415, P2_U5522);
  and ginst16070 (P2_U3851, P2_U3415, P2_U5527);
  and ginst16071 (P2_U3852, P2_U3415, P2_U5530);
  and ginst16072 (P2_U3853, P2_U3854, P2_U5531);
  and ginst16073 (P2_U3854, P2_U3415, P2_U5533);
  and ginst16074 (P2_U3855, P2_U3856, P2_U5534);
  and ginst16075 (P2_U3856, P2_U3415, P2_U5536);
  and ginst16076 (P2_U3857, P2_U5539, P2_U5540);
  and ginst16077 (P2_U3858, P2_U5542, P2_U5543);
  and ginst16078 (P2_U3859, P2_U5564, P2_U5565);
  and ginst16079 (P2_U3860, P2_U5567, P2_U5568);
  and ginst16080 (P2_U3861, P2_U5570, P2_U5571);
  and ginst16081 (P2_U3862, P2_U5573, P2_U5574);
  and ginst16082 (P2_U3863, P2_U5576, P2_U5577);
  and ginst16083 (P2_U3864, P2_U5579, P2_U5580);
  and ginst16084 (P2_U3865, P2_U5582, P2_U5583);
  and ginst16085 (P2_U3866, P2_U5585, P2_U5586);
  and ginst16086 (P2_U3867, P2_U5588, P2_U5589);
  and ginst16087 (P2_U3868, P2_U5591, P2_U5592);
  and ginst16088 (P2_U3869, P2_U5597, P2_U5598);
  and ginst16089 (P2_U3870, P2_U5600, P2_U5601);
  and ginst16090 (P2_U3871, P2_U5603, P2_U5604);
  and ginst16091 (P2_U3872, P2_U5606, P2_U5607);
  and ginst16092 (P2_U3873, P2_U5609, P2_U5610);
  and ginst16093 (P2_U3874, P2_U5612, P2_U5613);
  and ginst16094 (P2_U3875, P2_U5615, P2_U5616);
  and ginst16095 (P2_U3876, P2_U5618, P2_U5619);
  and ginst16096 (P2_U3877, P2_U5621, P2_U5622);
  and ginst16097 (P2_U3878, P2_U5624, P2_U5625);
  not ginst16098 (P2_U3879, P2_IR_REG_31__SCAN_IN);
  nand ginst16099 (P2_U3880, P2_U3023, P2_U3333);
  nand ginst16100 (P2_U3881, P2_U3050, P2_U3577);
  nand ginst16101 (P2_U3882, P2_U3050, P2_U3695);
  and ginst16102 (P2_U3883, P2_U5921, P2_U5922);
  and ginst16103 (P2_U3884, P2_U5923, P2_U5924);
  and ginst16104 (P2_U3885, P2_U5925, P2_U5926);
  and ginst16105 (P2_U3886, P2_U5927, P2_U5928);
  and ginst16106 (P2_U3887, P2_U5929, P2_U5930);
  and ginst16107 (P2_U3888, P2_U5931, P2_U5932);
  and ginst16108 (P2_U3889, P2_U5933, P2_U5934);
  and ginst16109 (P2_U3890, P2_U5935, P2_U5936);
  and ginst16110 (P2_U3891, P2_U5937, P2_U5938);
  and ginst16111 (P2_U3892, P2_U5939, P2_U5940);
  and ginst16112 (P2_U3893, P2_U5941, P2_U5942);
  and ginst16113 (P2_U3894, P2_U5943, P2_U5944);
  and ginst16114 (P2_U3895, P2_U5945, P2_U5946);
  and ginst16115 (P2_U3896, P2_U5947, P2_U5948);
  and ginst16116 (P2_U3897, P2_U5949, P2_U5950);
  and ginst16117 (P2_U3898, P2_U5951, P2_U5952);
  and ginst16118 (P2_U3899, P2_U5953, P2_U5954);
  and ginst16119 (P2_U3900, P2_U5955, P2_U5956);
  and ginst16120 (P2_U3901, P2_U5957, P2_U5958);
  and ginst16121 (P2_U3902, P2_U5959, P2_U5960);
  and ginst16122 (P2_U3903, P2_U5961, P2_U5962);
  and ginst16123 (P2_U3904, P2_U5963, P2_U5964);
  and ginst16124 (P2_U3905, P2_U5965, P2_U5966);
  and ginst16125 (P2_U3906, P2_U5967, P2_U5968);
  and ginst16126 (P2_U3907, P2_U5969, P2_U5970);
  and ginst16127 (P2_U3908, P2_U5971, P2_U5972);
  and ginst16128 (P2_U3909, P2_U5973, P2_U5974);
  and ginst16129 (P2_U3910, P2_U5975, P2_U5976);
  and ginst16130 (P2_U3911, P2_U5977, P2_U5978);
  and ginst16131 (P2_U3912, P2_U5979, P2_U5980);
  nand ginst16132 (P2_U3913, P2_U3058, P2_U3694);
  and ginst16133 (P2_U3914, P2_U5981, P2_U5982);
  and ginst16134 (P2_U3915, P2_U5983, P2_U5984);
  not ginst16135 (P2_U3916, P2_R1312_U18);
  and ginst16136 (P2_U3917, P2_U6049, P2_U6050);
  nand ginst16137 (P2_U3918, P2_U3792, P2_U3793, P2_U3794, P2_U6082, P2_U6085);
  nand ginst16138 (P2_U3919, P2_U3049, P2_U5674);
  nand ginst16139 (P2_U3920, P2_U3418, P2_U3973);
  not ginst16140 (P2_U3921, P2_U3390);
  not ginst16141 (P2_U3922, P2_U3342);
  nand ginst16142 (P2_U3923, P2_U3418, P2_U3976);
  not ginst16143 (P2_U3924, P2_U3339);
  not ginst16144 (P2_U3925, P2_U3346);
  not ginst16145 (P2_U3926, P2_U3336);
  not ginst16146 (P2_U3927, P2_U3394);
  nand ginst16147 (P2_U3928, P2_U3420, P2_U3973);
  not ginst16148 (P2_U3929, P2_U3410);
  not ginst16149 (P2_U3930, P2_U3335);
  not ginst16150 (P2_U3931, P2_U3334);
  not ginst16151 (P2_U3932, P2_U3395);
  not ginst16152 (P2_U3933, P2_U3393);
  nand ginst16153 (P2_U3934, P2_U3925, P2_U5674);
  nand ginst16154 (P2_U3935, P2_U3340, P2_U3963);
  nand ginst16155 (P2_U3936, P2_U3973, P2_U5671);
  not ginst16156 (P2_U3937, P2_U3402);
  not ginst16157 (P2_U3938, P2_U3392);
  not ginst16158 (P2_U3939, P2_U3341);
  not ginst16159 (P2_U3940, P2_U3919);
  not ginst16160 (P2_U3941, P2_U3337);
  not ginst16161 (P2_U3942, P2_U3920);
  not ginst16162 (P2_U3943, P2_U3338);
  not ginst16163 (P2_U3944, P2_U3343);
  not ginst16164 (P2_U3945, P2_U3347);
  not ginst16165 (P2_U3946, P2_U3406);
  not ginst16166 (P2_U3947, P2_U3400);
  not ginst16167 (P2_U3948, P2_U3397);
  not ginst16168 (P2_U3949, P2_U3384);
  not ginst16169 (P2_U3950, P2_U3382);
  not ginst16170 (P2_U3951, P2_U3380);
  not ginst16171 (P2_U3952, P2_U3378);
  not ginst16172 (P2_U3953, P2_U3376);
  not ginst16173 (P2_U3954, P2_U3374);
  not ginst16174 (P2_U3955, P2_U3372);
  not ginst16175 (P2_U3956, P2_U3370);
  not ginst16176 (P2_U3957, P2_U3368);
  not ginst16177 (P2_U3958, P2_U3389);
  not ginst16178 (P2_U3959, P2_U3388);
  not ginst16179 (P2_U3960, P2_U3386);
  not ginst16180 (P2_U3961, P2_U3403);
  not ginst16181 (P2_U3962, P2_U3396);
  not ginst16182 (P2_U3963, P2_U3344);
  not ginst16183 (P2_U3964, P2_U3391);
  not ginst16184 (P2_U3965, P2_U3882);
  not ginst16185 (P2_U3966, P2_U3881);
  not ginst16186 (P2_U3967, P2_U3880);
  not ginst16187 (P2_U3968, P2_U3913);
  not ginst16188 (P2_U3969, P2_U3407);
  nand ginst16189 (P2_U3970, P2_STATE_REG_SCAN_IN, P2_U3408);
  nand ginst16190 (P2_U3971, P2_U3023, P2_U3933);
  not ginst16191 (P2_U3972, P2_U3405);
  not ginst16192 (P2_U3973, P2_U3404);
  not ginst16193 (P2_U3974, P2_U3340);
  not ginst16194 (P2_U3975, P2_U3332);
  not ginst16195 (P2_U3976, P2_U3345);
  not ginst16196 (P2_U3977, P2_U3399);
  not ginst16197 (P2_U3978, P2_U3329);
  nand ginst16198 (P2_U3979, P2_U3088, U93);
  nand ginst16199 (P2_U3980, P2_IR_REG_0__SCAN_IN, P2_U3030);
  nand ginst16200 (P2_U3981, P2_IR_REG_0__SCAN_IN, P2_U3978);
  nand ginst16201 (P2_U3982, P2_U3088, U82);
  nand ginst16202 (P2_U3983, P2_SUB_1108_U42, P2_U3030);
  nand ginst16203 (P2_U3984, P2_IR_REG_1__SCAN_IN, P2_U3978);
  nand ginst16204 (P2_U3985, P2_U3088, U71);
  nand ginst16205 (P2_U3986, P2_SUB_1108_U17, P2_U3030);
  nand ginst16206 (P2_U3987, P2_IR_REG_2__SCAN_IN, P2_U3978);
  nand ginst16207 (P2_U3988, P2_U3088, U68);
  nand ginst16208 (P2_U3989, P2_SUB_1108_U18, P2_U3030);
  nand ginst16209 (P2_U3990, P2_IR_REG_3__SCAN_IN, P2_U3978);
  nand ginst16210 (P2_U3991, P2_U3088, U67);
  nand ginst16211 (P2_U3992, P2_SUB_1108_U19, P2_U3030);
  nand ginst16212 (P2_U3993, P2_IR_REG_4__SCAN_IN, P2_U3978);
  nand ginst16213 (P2_U3994, P2_U3088, U66);
  nand ginst16214 (P2_U3995, P2_SUB_1108_U101, P2_U3030);
  nand ginst16215 (P2_U3996, P2_IR_REG_5__SCAN_IN, P2_U3978);
  nand ginst16216 (P2_U3997, P2_U3088, U65);
  nand ginst16217 (P2_U3998, P2_SUB_1108_U20, P2_U3030);
  nand ginst16218 (P2_U3999, P2_IR_REG_6__SCAN_IN, P2_U3978);
  nand ginst16219 (P2_U4000, P2_U3088, U64);
  nand ginst16220 (P2_U4001, P2_SUB_1108_U21, P2_U3030);
  nand ginst16221 (P2_U4002, P2_IR_REG_7__SCAN_IN, P2_U3978);
  nand ginst16222 (P2_U4003, P2_U3088, U63);
  nand ginst16223 (P2_U4004, P2_SUB_1108_U22, P2_U3030);
  nand ginst16224 (P2_U4005, P2_IR_REG_8__SCAN_IN, P2_U3978);
  nand ginst16225 (P2_U4006, P2_U3088, U62);
  nand ginst16226 (P2_U4007, P2_SUB_1108_U99, P2_U3030);
  nand ginst16227 (P2_U4008, P2_IR_REG_9__SCAN_IN, P2_U3978);
  nand ginst16228 (P2_U4009, P2_U3088, U92);
  nand ginst16229 (P2_U4010, P2_SUB_1108_U6, P2_U3030);
  nand ginst16230 (P2_U4011, P2_IR_REG_10__SCAN_IN, P2_U3978);
  nand ginst16231 (P2_U4012, P2_U3088, U91);
  nand ginst16232 (P2_U4013, P2_SUB_1108_U7, P2_U3030);
  nand ginst16233 (P2_U4014, P2_IR_REG_11__SCAN_IN, P2_U3978);
  nand ginst16234 (P2_U4015, P2_U3088, U90);
  nand ginst16235 (P2_U4016, P2_SUB_1108_U8, P2_U3030);
  nand ginst16236 (P2_U4017, P2_IR_REG_12__SCAN_IN, P2_U3978);
  nand ginst16237 (P2_U4018, P2_U3088, U89);
  nand ginst16238 (P2_U4019, P2_SUB_1108_U127, P2_U3030);
  nand ginst16239 (P2_U4020, P2_IR_REG_13__SCAN_IN, P2_U3978);
  nand ginst16240 (P2_U4021, P2_U3088, U88);
  nand ginst16241 (P2_U4022, P2_SUB_1108_U9, P2_U3030);
  nand ginst16242 (P2_U4023, P2_IR_REG_14__SCAN_IN, P2_U3978);
  nand ginst16243 (P2_U4024, P2_U3088, U87);
  nand ginst16244 (P2_U4025, P2_SUB_1108_U10, P2_U3030);
  nand ginst16245 (P2_U4026, P2_IR_REG_15__SCAN_IN, P2_U3978);
  nand ginst16246 (P2_U4027, P2_U3088, U86);
  nand ginst16247 (P2_U4028, P2_SUB_1108_U11, P2_U3030);
  nand ginst16248 (P2_U4029, P2_IR_REG_16__SCAN_IN, P2_U3978);
  nand ginst16249 (P2_U4030, P2_U3088, U85);
  nand ginst16250 (P2_U4031, P2_SUB_1108_U125, P2_U3030);
  nand ginst16251 (P2_U4032, P2_IR_REG_17__SCAN_IN, P2_U3978);
  nand ginst16252 (P2_U4033, P2_U3088, U84);
  nand ginst16253 (P2_U4034, P2_SUB_1108_U12, P2_U3030);
  nand ginst16254 (P2_U4035, P2_IR_REG_18__SCAN_IN, P2_U3978);
  nand ginst16255 (P2_U4036, P2_U3088, U83);
  nand ginst16256 (P2_U4037, P2_SUB_1108_U123, P2_U3030);
  nand ginst16257 (P2_U4038, P2_IR_REG_19__SCAN_IN, P2_U3978);
  nand ginst16258 (P2_U4039, P2_U3088, U81);
  nand ginst16259 (P2_U4040, P2_SUB_1108_U119, P2_U3030);
  nand ginst16260 (P2_U4041, P2_IR_REG_20__SCAN_IN, P2_U3978);
  nand ginst16261 (P2_U4042, P2_U3088, U80);
  nand ginst16262 (P2_U4043, P2_SUB_1108_U116, P2_U3030);
  nand ginst16263 (P2_U4044, P2_IR_REG_21__SCAN_IN, P2_U3978);
  nand ginst16264 (P2_U4045, P2_U3088, U79);
  nand ginst16265 (P2_U4046, P2_SUB_1108_U114, P2_U3030);
  nand ginst16266 (P2_U4047, P2_IR_REG_22__SCAN_IN, P2_U3978);
  nand ginst16267 (P2_U4048, P2_U3088, U78);
  nand ginst16268 (P2_U4049, P2_SUB_1108_U13, P2_U3030);
  nand ginst16269 (P2_U4050, P2_IR_REG_23__SCAN_IN, P2_U3978);
  nand ginst16270 (P2_U4051, P2_U3088, U77);
  nand ginst16271 (P2_U4052, P2_SUB_1108_U14, P2_U3030);
  nand ginst16272 (P2_U4053, P2_IR_REG_24__SCAN_IN, P2_U3978);
  nand ginst16273 (P2_U4054, P2_U3088, U76);
  nand ginst16274 (P2_U4055, P2_SUB_1108_U112, P2_U3030);
  nand ginst16275 (P2_U4056, P2_IR_REG_25__SCAN_IN, P2_U3978);
  nand ginst16276 (P2_U4057, P2_U3088, U75);
  nand ginst16277 (P2_U4058, P2_SUB_1108_U15, P2_U3030);
  nand ginst16278 (P2_U4059, P2_IR_REG_26__SCAN_IN, P2_U3978);
  nand ginst16279 (P2_U4060, P2_U3088, U74);
  nand ginst16280 (P2_U4061, P2_SUB_1108_U110, P2_U3030);
  nand ginst16281 (P2_U4062, P2_IR_REG_27__SCAN_IN, P2_U3978);
  nand ginst16282 (P2_U4063, P2_U3088, U73);
  nand ginst16283 (P2_U4064, P2_SUB_1108_U107, P2_U3030);
  nand ginst16284 (P2_U4065, P2_IR_REG_28__SCAN_IN, P2_U3978);
  nand ginst16285 (P2_U4066, P2_U3088, U72);
  nand ginst16286 (P2_U4067, P2_SUB_1108_U16, P2_U3030);
  nand ginst16287 (P2_U4068, P2_IR_REG_29__SCAN_IN, P2_U3978);
  nand ginst16288 (P2_U4069, P2_U3088, U70);
  nand ginst16289 (P2_U4070, P2_SUB_1108_U104, P2_U3030);
  nand ginst16290 (P2_U4071, P2_IR_REG_30__SCAN_IN, P2_U3978);
  nand ginst16291 (P2_U4072, P2_U3088, U69);
  nand ginst16292 (P2_U4073, P2_SUB_1108_U43, P2_U3030);
  nand ginst16293 (P2_U4074, P2_IR_REG_31__SCAN_IN, P2_U3978);
  nand ginst16294 (P2_U4075, P2_U3975, P2_U5655);
  not ginst16295 (P2_U4076, P2_U3333);
  nand ginst16296 (P2_U4077, P2_U3332, P2_U5646);
  nand ginst16297 (P2_U4078, P2_U3332, P2_U5649);
  nand ginst16298 (P2_U4079, P2_D_REG_10__SCAN_IN, P2_U4076);
  nand ginst16299 (P2_U4080, P2_D_REG_11__SCAN_IN, P2_U4076);
  nand ginst16300 (P2_U4081, P2_D_REG_12__SCAN_IN, P2_U4076);
  nand ginst16301 (P2_U4082, P2_D_REG_13__SCAN_IN, P2_U4076);
  nand ginst16302 (P2_U4083, P2_D_REG_14__SCAN_IN, P2_U4076);
  nand ginst16303 (P2_U4084, P2_D_REG_15__SCAN_IN, P2_U4076);
  nand ginst16304 (P2_U4085, P2_D_REG_16__SCAN_IN, P2_U4076);
  nand ginst16305 (P2_U4086, P2_D_REG_17__SCAN_IN, P2_U4076);
  nand ginst16306 (P2_U4087, P2_D_REG_18__SCAN_IN, P2_U4076);
  nand ginst16307 (P2_U4088, P2_D_REG_19__SCAN_IN, P2_U4076);
  nand ginst16308 (P2_U4089, P2_D_REG_20__SCAN_IN, P2_U4076);
  nand ginst16309 (P2_U4090, P2_D_REG_21__SCAN_IN, P2_U4076);
  nand ginst16310 (P2_U4091, P2_D_REG_22__SCAN_IN, P2_U4076);
  nand ginst16311 (P2_U4092, P2_D_REG_23__SCAN_IN, P2_U4076);
  nand ginst16312 (P2_U4093, P2_D_REG_24__SCAN_IN, P2_U4076);
  nand ginst16313 (P2_U4094, P2_D_REG_25__SCAN_IN, P2_U4076);
  nand ginst16314 (P2_U4095, P2_D_REG_26__SCAN_IN, P2_U4076);
  nand ginst16315 (P2_U4096, P2_D_REG_27__SCAN_IN, P2_U4076);
  nand ginst16316 (P2_U4097, P2_D_REG_28__SCAN_IN, P2_U4076);
  nand ginst16317 (P2_U4098, P2_D_REG_29__SCAN_IN, P2_U4076);
  nand ginst16318 (P2_U4099, P2_D_REG_2__SCAN_IN, P2_U4076);
  nand ginst16319 (P2_U4100, P2_D_REG_30__SCAN_IN, P2_U4076);
  nand ginst16320 (P2_U4101, P2_D_REG_31__SCAN_IN, P2_U4076);
  nand ginst16321 (P2_U4102, P2_D_REG_3__SCAN_IN, P2_U4076);
  nand ginst16322 (P2_U4103, P2_D_REG_4__SCAN_IN, P2_U4076);
  nand ginst16323 (P2_U4104, P2_D_REG_5__SCAN_IN, P2_U4076);
  nand ginst16324 (P2_U4105, P2_D_REG_6__SCAN_IN, P2_U4076);
  nand ginst16325 (P2_U4106, P2_D_REG_7__SCAN_IN, P2_U4076);
  nand ginst16326 (P2_U4107, P2_D_REG_8__SCAN_IN, P2_U4076);
  nand ginst16327 (P2_U4108, P2_D_REG_9__SCAN_IN, P2_U4076);
  nand ginst16328 (P2_U4109, P2_U5671, P2_U5674);
  nand ginst16329 (P2_U4110, P2_U3340, P2_U5692, P2_U5693);
  nand ginst16330 (P2_U4111, P2_REG2_REG_1__SCAN_IN, P2_U3020);
  nand ginst16331 (P2_U4112, P2_REG1_REG_1__SCAN_IN, P2_U3021);
  nand ginst16332 (P2_U4113, P2_REG0_REG_1__SCAN_IN, P2_U3022);
  nand ginst16333 (P2_U4114, P2_REG3_REG_1__SCAN_IN, P2_U3019);
  not ginst16334 (P2_U4115, P2_U3080);
  nand ginst16335 (P2_U4116, P2_U3390, P2_U3934);
  nand ginst16336 (P2_U4117, P2_R1146_U20, P2_U3931);
  nand ginst16337 (P2_U4118, P2_R1113_U20, P2_U3930);
  nand ginst16338 (P2_U4119, P2_R1131_U95, P2_U3926);
  nand ginst16339 (P2_U4120, P2_R1179_U20, P2_U3941);
  nand ginst16340 (P2_U4121, P2_R1203_U20, P2_U3943);
  nand ginst16341 (P2_U4122, P2_R1164_U95, P2_U3014);
  nand ginst16342 (P2_U4123, P2_R1233_U95, P2_U3922);
  not ginst16343 (P2_U4124, P2_U3348);
  nand ginst16344 (P2_U4125, P2_U3027, P2_U3427);
  nand ginst16345 (P2_U4126, P2_U3026, P2_U3080);
  nand ginst16346 (P2_U4127, P2_R1215_U96, P2_U3025);
  nand ginst16347 (P2_U4128, P2_U3427, P2_U4116);
  nand ginst16348 (P2_U4129, P2_U3565, P2_U4124, P2_U4126, P2_U4128);
  nand ginst16349 (P2_U4130, P2_REG2_REG_2__SCAN_IN, P2_U3020);
  nand ginst16350 (P2_U4131, P2_REG1_REG_2__SCAN_IN, P2_U3021);
  nand ginst16351 (P2_U4132, P2_REG0_REG_2__SCAN_IN, P2_U3022);
  nand ginst16352 (P2_U4133, P2_REG3_REG_2__SCAN_IN, P2_U3019);
  not ginst16353 (P2_U4134, P2_U3070);
  nand ginst16354 (P2_U4135, P2_REG2_REG_0__SCAN_IN, P2_U3020);
  nand ginst16355 (P2_U4136, P2_REG1_REG_0__SCAN_IN, P2_U3021);
  nand ginst16356 (P2_U4137, P2_REG0_REG_0__SCAN_IN, P2_U3022);
  nand ginst16357 (P2_U4138, P2_REG3_REG_0__SCAN_IN, P2_U3019);
  not ginst16358 (P2_U4139, P2_U3079);
  nand ginst16359 (P2_U4140, P2_U3035, P2_U3079);
  nand ginst16360 (P2_U4141, P2_R1146_U97, P2_U3931);
  nand ginst16361 (P2_U4142, P2_R1113_U97, P2_U3930);
  nand ginst16362 (P2_U4143, P2_R1131_U94, P2_U3926);
  nand ginst16363 (P2_U4144, P2_R1179_U97, P2_U3941);
  nand ginst16364 (P2_U4145, P2_R1203_U97, P2_U3943);
  nand ginst16365 (P2_U4146, P2_R1164_U94, P2_U3014);
  nand ginst16366 (P2_U4147, P2_R1233_U94, P2_U3922);
  not ginst16367 (P2_U4148, P2_U3349);
  nand ginst16368 (P2_U4149, P2_R1275_U55, P2_U3027);
  nand ginst16369 (P2_U4150, P2_U3026, P2_U3070);
  nand ginst16370 (P2_U4151, P2_R1215_U95, P2_U3025);
  nand ginst16371 (P2_U4152, P2_U3432, P2_U4116);
  nand ginst16372 (P2_U4153, P2_U3581, P2_U4148);
  nand ginst16373 (P2_U4154, P2_REG2_REG_3__SCAN_IN, P2_U3020);
  nand ginst16374 (P2_U4155, P2_REG1_REG_3__SCAN_IN, P2_U3021);
  nand ginst16375 (P2_U4156, P2_REG0_REG_3__SCAN_IN, P2_U3022);
  nand ginst16376 (P2_U4157, P2_ADD_1119_U4, P2_U3019);
  not ginst16377 (P2_U4158, P2_U3066);
  nand ginst16378 (P2_U4159, P2_U3035, P2_U3080);
  nand ginst16379 (P2_U4160, P2_R1146_U107, P2_U3931);
  nand ginst16380 (P2_U4161, P2_R1113_U107, P2_U3930);
  nand ginst16381 (P2_U4162, P2_R1131_U16, P2_U3926);
  nand ginst16382 (P2_U4163, P2_R1179_U107, P2_U3941);
  nand ginst16383 (P2_U4164, P2_R1203_U107, P2_U3943);
  nand ginst16384 (P2_U4165, P2_R1164_U16, P2_U3014);
  nand ginst16385 (P2_U4166, P2_R1233_U16, P2_U3922);
  not ginst16386 (P2_U4167, P2_U3350);
  nand ginst16387 (P2_U4168, P2_R1275_U18, P2_U3027);
  nand ginst16388 (P2_U4169, P2_U3026, P2_U3066);
  nand ginst16389 (P2_U4170, P2_R1215_U17, P2_U3025);
  nand ginst16390 (P2_U4171, P2_U3435, P2_U4116);
  nand ginst16391 (P2_U4172, P2_U3585, P2_U4167);
  nand ginst16392 (P2_U4173, P2_REG2_REG_4__SCAN_IN, P2_U3020);
  nand ginst16393 (P2_U4174, P2_REG1_REG_4__SCAN_IN, P2_U3021);
  nand ginst16394 (P2_U4175, P2_REG0_REG_4__SCAN_IN, P2_U3022);
  nand ginst16395 (P2_U4176, P2_ADD_1119_U55, P2_U3019);
  not ginst16396 (P2_U4177, P2_U3062);
  nand ginst16397 (P2_U4178, P2_U3035, P2_U3070);
  nand ginst16398 (P2_U4179, P2_R1146_U17, P2_U3931);
  nand ginst16399 (P2_U4180, P2_R1113_U17, P2_U3930);
  nand ginst16400 (P2_U4181, P2_R1131_U100, P2_U3926);
  nand ginst16401 (P2_U4182, P2_R1179_U17, P2_U3941);
  nand ginst16402 (P2_U4183, P2_R1203_U17, P2_U3943);
  nand ginst16403 (P2_U4184, P2_R1164_U100, P2_U3014);
  nand ginst16404 (P2_U4185, P2_R1233_U100, P2_U3922);
  not ginst16405 (P2_U4186, P2_U3351);
  nand ginst16406 (P2_U4187, P2_R1275_U20, P2_U3027);
  nand ginst16407 (P2_U4188, P2_U3026, P2_U3062);
  nand ginst16408 (P2_U4189, P2_R1215_U101, P2_U3025);
  nand ginst16409 (P2_U4190, P2_U3438, P2_U4116);
  nand ginst16410 (P2_U4191, P2_U3589, P2_U4186);
  nand ginst16411 (P2_U4192, P2_REG2_REG_5__SCAN_IN, P2_U3020);
  nand ginst16412 (P2_U4193, P2_REG1_REG_5__SCAN_IN, P2_U3021);
  nand ginst16413 (P2_U4194, P2_REG0_REG_5__SCAN_IN, P2_U3022);
  nand ginst16414 (P2_U4195, P2_ADD_1119_U54, P2_U3019);
  not ginst16415 (P2_U4196, P2_U3069);
  nand ginst16416 (P2_U4197, P2_U3035, P2_U3066);
  nand ginst16417 (P2_U4198, P2_R1146_U106, P2_U3931);
  nand ginst16418 (P2_U4199, P2_R1113_U106, P2_U3930);
  nand ginst16419 (P2_U4200, P2_R1131_U99, P2_U3926);
  nand ginst16420 (P2_U4201, P2_R1179_U106, P2_U3941);
  nand ginst16421 (P2_U4202, P2_R1203_U106, P2_U3943);
  nand ginst16422 (P2_U4203, P2_R1164_U99, P2_U3014);
  nand ginst16423 (P2_U4204, P2_R1233_U99, P2_U3922);
  not ginst16424 (P2_U4205, P2_U3352);
  nand ginst16425 (P2_U4206, P2_R1275_U21, P2_U3027);
  nand ginst16426 (P2_U4207, P2_U3026, P2_U3069);
  nand ginst16427 (P2_U4208, P2_R1215_U100, P2_U3025);
  nand ginst16428 (P2_U4209, P2_U3441, P2_U4116);
  nand ginst16429 (P2_U4210, P2_U3593, P2_U4205);
  nand ginst16430 (P2_U4211, P2_REG2_REG_6__SCAN_IN, P2_U3020);
  nand ginst16431 (P2_U4212, P2_REG1_REG_6__SCAN_IN, P2_U3021);
  nand ginst16432 (P2_U4213, P2_REG0_REG_6__SCAN_IN, P2_U3022);
  nand ginst16433 (P2_U4214, P2_ADD_1119_U53, P2_U3019);
  not ginst16434 (P2_U4215, P2_U3073);
  nand ginst16435 (P2_U4216, P2_U3035, P2_U3062);
  nand ginst16436 (P2_U4217, P2_R1146_U105, P2_U3931);
  nand ginst16437 (P2_U4218, P2_R1113_U105, P2_U3930);
  nand ginst16438 (P2_U4219, P2_R1131_U17, P2_U3926);
  nand ginst16439 (P2_U4220, P2_R1179_U105, P2_U3941);
  nand ginst16440 (P2_U4221, P2_R1203_U105, P2_U3943);
  nand ginst16441 (P2_U4222, P2_R1164_U17, P2_U3014);
  nand ginst16442 (P2_U4223, P2_R1233_U17, P2_U3922);
  not ginst16443 (P2_U4224, P2_U3353);
  nand ginst16444 (P2_U4225, P2_R1275_U65, P2_U3027);
  nand ginst16445 (P2_U4226, P2_U3026, P2_U3073);
  nand ginst16446 (P2_U4227, P2_R1215_U18, P2_U3025);
  nand ginst16447 (P2_U4228, P2_U3444, P2_U4116);
  nand ginst16448 (P2_U4229, P2_U3597, P2_U4224);
  nand ginst16449 (P2_U4230, P2_REG2_REG_7__SCAN_IN, P2_U3020);
  nand ginst16450 (P2_U4231, P2_REG1_REG_7__SCAN_IN, P2_U3021);
  nand ginst16451 (P2_U4232, P2_REG0_REG_7__SCAN_IN, P2_U3022);
  nand ginst16452 (P2_U4233, P2_ADD_1119_U52, P2_U3019);
  not ginst16453 (P2_U4234, P2_U3072);
  nand ginst16454 (P2_U4235, P2_U3035, P2_U3069);
  nand ginst16455 (P2_U4236, P2_R1146_U18, P2_U3931);
  nand ginst16456 (P2_U4237, P2_R1113_U18, P2_U3930);
  nand ginst16457 (P2_U4238, P2_R1131_U98, P2_U3926);
  nand ginst16458 (P2_U4239, P2_R1179_U18, P2_U3941);
  nand ginst16459 (P2_U4240, P2_R1203_U18, P2_U3943);
  nand ginst16460 (P2_U4241, P2_R1164_U98, P2_U3014);
  nand ginst16461 (P2_U4242, P2_R1233_U98, P2_U3922);
  not ginst16462 (P2_U4243, P2_U3354);
  nand ginst16463 (P2_U4244, P2_R1275_U22, P2_U3027);
  nand ginst16464 (P2_U4245, P2_U3026, P2_U3072);
  nand ginst16465 (P2_U4246, P2_R1215_U99, P2_U3025);
  nand ginst16466 (P2_U4247, P2_U3447, P2_U4116);
  nand ginst16467 (P2_U4248, P2_U3601, P2_U4243);
  nand ginst16468 (P2_U4249, P2_REG2_REG_8__SCAN_IN, P2_U3020);
  nand ginst16469 (P2_U4250, P2_REG1_REG_8__SCAN_IN, P2_U3021);
  nand ginst16470 (P2_U4251, P2_REG0_REG_8__SCAN_IN, P2_U3022);
  nand ginst16471 (P2_U4252, P2_ADD_1119_U51, P2_U3019);
  not ginst16472 (P2_U4253, P2_U3086);
  nand ginst16473 (P2_U4254, P2_U3035, P2_U3073);
  nand ginst16474 (P2_U4255, P2_R1146_U104, P2_U3931);
  nand ginst16475 (P2_U4256, P2_R1113_U104, P2_U3930);
  nand ginst16476 (P2_U4257, P2_R1131_U18, P2_U3926);
  nand ginst16477 (P2_U4258, P2_R1179_U104, P2_U3941);
  nand ginst16478 (P2_U4259, P2_R1203_U104, P2_U3943);
  nand ginst16479 (P2_U4260, P2_R1164_U18, P2_U3014);
  nand ginst16480 (P2_U4261, P2_R1233_U18, P2_U3922);
  not ginst16481 (P2_U4262, P2_U3355);
  nand ginst16482 (P2_U4263, P2_R1275_U23, P2_U3027);
  nand ginst16483 (P2_U4264, P2_U3026, P2_U3086);
  nand ginst16484 (P2_U4265, P2_R1215_U19, P2_U3025);
  nand ginst16485 (P2_U4266, P2_U3450, P2_U4116);
  nand ginst16486 (P2_U4267, P2_U3605, P2_U4262);
  nand ginst16487 (P2_U4268, P2_REG2_REG_9__SCAN_IN, P2_U3020);
  nand ginst16488 (P2_U4269, P2_REG1_REG_9__SCAN_IN, P2_U3021);
  nand ginst16489 (P2_U4270, P2_REG0_REG_9__SCAN_IN, P2_U3022);
  nand ginst16490 (P2_U4271, P2_ADD_1119_U50, P2_U3019);
  not ginst16491 (P2_U4272, P2_U3085);
  nand ginst16492 (P2_U4273, P2_U3035, P2_U3072);
  nand ginst16493 (P2_U4274, P2_R1146_U19, P2_U3931);
  nand ginst16494 (P2_U4275, P2_R1113_U19, P2_U3930);
  nand ginst16495 (P2_U4276, P2_R1131_U97, P2_U3926);
  nand ginst16496 (P2_U4277, P2_R1179_U19, P2_U3941);
  nand ginst16497 (P2_U4278, P2_R1203_U19, P2_U3943);
  nand ginst16498 (P2_U4279, P2_R1164_U97, P2_U3014);
  nand ginst16499 (P2_U4280, P2_R1233_U97, P2_U3922);
  not ginst16500 (P2_U4281, P2_U3356);
  nand ginst16501 (P2_U4282, P2_R1275_U24, P2_U3027);
  nand ginst16502 (P2_U4283, P2_U3026, P2_U3085);
  nand ginst16503 (P2_U4284, P2_R1215_U98, P2_U3025);
  nand ginst16504 (P2_U4285, P2_U3453, P2_U4116);
  nand ginst16505 (P2_U4286, P2_U3609, P2_U4281);
  nand ginst16506 (P2_U4287, P2_REG2_REG_10__SCAN_IN, P2_U3020);
  nand ginst16507 (P2_U4288, P2_REG1_REG_10__SCAN_IN, P2_U3021);
  nand ginst16508 (P2_U4289, P2_REG0_REG_10__SCAN_IN, P2_U3022);
  nand ginst16509 (P2_U4290, P2_ADD_1119_U74, P2_U3019);
  not ginst16510 (P2_U4291, P2_U3064);
  nand ginst16511 (P2_U4292, P2_U3035, P2_U3086);
  nand ginst16512 (P2_U4293, P2_R1146_U103, P2_U3931);
  nand ginst16513 (P2_U4294, P2_R1113_U103, P2_U3930);
  nand ginst16514 (P2_U4295, P2_R1131_U96, P2_U3926);
  nand ginst16515 (P2_U4296, P2_R1179_U103, P2_U3941);
  nand ginst16516 (P2_U4297, P2_R1203_U103, P2_U3943);
  nand ginst16517 (P2_U4298, P2_R1164_U96, P2_U3014);
  nand ginst16518 (P2_U4299, P2_R1233_U96, P2_U3922);
  not ginst16519 (P2_U4300, P2_U3357);
  nand ginst16520 (P2_U4301, P2_R1275_U63, P2_U3027);
  nand ginst16521 (P2_U4302, P2_U3026, P2_U3064);
  nand ginst16522 (P2_U4303, P2_R1215_U97, P2_U3025);
  nand ginst16523 (P2_U4304, P2_U3456, P2_U4116);
  nand ginst16524 (P2_U4305, P2_U3613, P2_U4300);
  nand ginst16525 (P2_U4306, P2_REG2_REG_11__SCAN_IN, P2_U3020);
  nand ginst16526 (P2_U4307, P2_REG1_REG_11__SCAN_IN, P2_U3021);
  nand ginst16527 (P2_U4308, P2_REG0_REG_11__SCAN_IN, P2_U3022);
  nand ginst16528 (P2_U4309, P2_ADD_1119_U73, P2_U3019);
  not ginst16529 (P2_U4310, P2_U3065);
  nand ginst16530 (P2_U4311, P2_U3035, P2_U3085);
  nand ginst16531 (P2_U4312, P2_R1146_U113, P2_U3931);
  nand ginst16532 (P2_U4313, P2_R1113_U113, P2_U3930);
  nand ginst16533 (P2_U4314, P2_R1131_U10, P2_U3926);
  nand ginst16534 (P2_U4315, P2_R1179_U113, P2_U3941);
  nand ginst16535 (P2_U4316, P2_R1203_U113, P2_U3943);
  nand ginst16536 (P2_U4317, P2_R1164_U10, P2_U3014);
  nand ginst16537 (P2_U4318, P2_R1233_U10, P2_U3922);
  not ginst16538 (P2_U4319, P2_U3358);
  nand ginst16539 (P2_U4320, P2_R1275_U6, P2_U3027);
  nand ginst16540 (P2_U4321, P2_U3026, P2_U3065);
  nand ginst16541 (P2_U4322, P2_R1215_U11, P2_U3025);
  nand ginst16542 (P2_U4323, P2_U3459, P2_U4116);
  nand ginst16543 (P2_U4324, P2_U3617, P2_U4319);
  nand ginst16544 (P2_U4325, P2_REG2_REG_12__SCAN_IN, P2_U3020);
  nand ginst16545 (P2_U4326, P2_REG1_REG_12__SCAN_IN, P2_U3021);
  nand ginst16546 (P2_U4327, P2_REG0_REG_12__SCAN_IN, P2_U3022);
  nand ginst16547 (P2_U4328, P2_ADD_1119_U72, P2_U3019);
  not ginst16548 (P2_U4329, P2_U3074);
  nand ginst16549 (P2_U4330, P2_U3035, P2_U3064);
  nand ginst16550 (P2_U4331, P2_R1146_U12, P2_U3931);
  nand ginst16551 (P2_U4332, P2_R1113_U12, P2_U3930);
  nand ginst16552 (P2_U4333, P2_R1131_U114, P2_U3926);
  nand ginst16553 (P2_U4334, P2_R1179_U12, P2_U3941);
  nand ginst16554 (P2_U4335, P2_R1203_U12, P2_U3943);
  nand ginst16555 (P2_U4336, P2_R1164_U114, P2_U3014);
  nand ginst16556 (P2_U4337, P2_R1233_U114, P2_U3922);
  not ginst16557 (P2_U4338, P2_U3359);
  nand ginst16558 (P2_U4339, P2_R1275_U7, P2_U3027);
  nand ginst16559 (P2_U4340, P2_U3026, P2_U3074);
  nand ginst16560 (P2_U4341, P2_R1215_U115, P2_U3025);
  nand ginst16561 (P2_U4342, P2_U3462, P2_U4116);
  nand ginst16562 (P2_U4343, P2_U3621, P2_U4338);
  nand ginst16563 (P2_U4344, P2_REG2_REG_13__SCAN_IN, P2_U3020);
  nand ginst16564 (P2_U4345, P2_REG1_REG_13__SCAN_IN, P2_U3021);
  nand ginst16565 (P2_U4346, P2_REG0_REG_13__SCAN_IN, P2_U3022);
  nand ginst16566 (P2_U4347, P2_ADD_1119_U71, P2_U3019);
  not ginst16567 (P2_U4348, P2_U3082);
  nand ginst16568 (P2_U4349, P2_U3035, P2_U3065);
  nand ginst16569 (P2_U4350, P2_R1146_U102, P2_U3931);
  nand ginst16570 (P2_U4351, P2_R1113_U102, P2_U3930);
  nand ginst16571 (P2_U4352, P2_R1131_U113, P2_U3926);
  nand ginst16572 (P2_U4353, P2_R1179_U102, P2_U3941);
  nand ginst16573 (P2_U4354, P2_R1203_U102, P2_U3943);
  nand ginst16574 (P2_U4355, P2_R1164_U113, P2_U3014);
  nand ginst16575 (P2_U4356, P2_R1233_U113, P2_U3922);
  not ginst16576 (P2_U4357, P2_U3360);
  nand ginst16577 (P2_U4358, P2_R1275_U8, P2_U3027);
  nand ginst16578 (P2_U4359, P2_U3026, P2_U3082);
  nand ginst16579 (P2_U4360, P2_R1215_U114, P2_U3025);
  nand ginst16580 (P2_U4361, P2_U3465, P2_U4116);
  nand ginst16581 (P2_U4362, P2_U3625, P2_U4357);
  nand ginst16582 (P2_U4363, P2_REG2_REG_14__SCAN_IN, P2_U3020);
  nand ginst16583 (P2_U4364, P2_REG1_REG_14__SCAN_IN, P2_U3021);
  nand ginst16584 (P2_U4365, P2_REG0_REG_14__SCAN_IN, P2_U3022);
  nand ginst16585 (P2_U4366, P2_ADD_1119_U70, P2_U3019);
  not ginst16586 (P2_U4367, P2_U3081);
  nand ginst16587 (P2_U4368, P2_U3035, P2_U3074);
  nand ginst16588 (P2_U4369, P2_R1146_U101, P2_U3931);
  nand ginst16589 (P2_U4370, P2_R1113_U101, P2_U3930);
  nand ginst16590 (P2_U4371, P2_R1131_U11, P2_U3926);
  nand ginst16591 (P2_U4372, P2_R1179_U101, P2_U3941);
  nand ginst16592 (P2_U4373, P2_R1203_U101, P2_U3943);
  nand ginst16593 (P2_U4374, P2_R1164_U11, P2_U3014);
  nand ginst16594 (P2_U4375, P2_R1233_U11, P2_U3922);
  not ginst16595 (P2_U4376, P2_U3361);
  nand ginst16596 (P2_U4377, P2_R1275_U86, P2_U3027);
  nand ginst16597 (P2_U4378, P2_U3026, P2_U3081);
  nand ginst16598 (P2_U4379, P2_R1215_U12, P2_U3025);
  nand ginst16599 (P2_U4380, P2_U3468, P2_U4116);
  nand ginst16600 (P2_U4381, P2_U3629, P2_U4376);
  nand ginst16601 (P2_U4382, P2_REG2_REG_15__SCAN_IN, P2_U3020);
  nand ginst16602 (P2_U4383, P2_REG1_REG_15__SCAN_IN, P2_U3021);
  nand ginst16603 (P2_U4384, P2_REG0_REG_15__SCAN_IN, P2_U3022);
  nand ginst16604 (P2_U4385, P2_ADD_1119_U69, P2_U3019);
  not ginst16605 (P2_U4386, P2_U3076);
  nand ginst16606 (P2_U4387, P2_U3035, P2_U3082);
  nand ginst16607 (P2_U4388, P2_R1146_U112, P2_U3931);
  nand ginst16608 (P2_U4389, P2_R1113_U112, P2_U3930);
  nand ginst16609 (P2_U4390, P2_R1131_U112, P2_U3926);
  nand ginst16610 (P2_U4391, P2_R1179_U112, P2_U3941);
  nand ginst16611 (P2_U4392, P2_R1203_U112, P2_U3943);
  nand ginst16612 (P2_U4393, P2_R1164_U112, P2_U3014);
  nand ginst16613 (P2_U4394, P2_R1233_U112, P2_U3922);
  not ginst16614 (P2_U4395, P2_U3362);
  nand ginst16615 (P2_U4396, P2_R1275_U9, P2_U3027);
  nand ginst16616 (P2_U4397, P2_U3026, P2_U3076);
  nand ginst16617 (P2_U4398, P2_R1215_U113, P2_U3025);
  nand ginst16618 (P2_U4399, P2_U3471, P2_U4116);
  nand ginst16619 (P2_U4400, P2_U3633, P2_U4395);
  nand ginst16620 (P2_U4401, P2_REG2_REG_16__SCAN_IN, P2_U3020);
  nand ginst16621 (P2_U4402, P2_REG1_REG_16__SCAN_IN, P2_U3021);
  nand ginst16622 (P2_U4403, P2_REG0_REG_16__SCAN_IN, P2_U3022);
  nand ginst16623 (P2_U4404, P2_ADD_1119_U68, P2_U3019);
  not ginst16624 (P2_U4405, P2_U3075);
  nand ginst16625 (P2_U4406, P2_U3035, P2_U3081);
  nand ginst16626 (P2_U4407, P2_R1146_U111, P2_U3931);
  nand ginst16627 (P2_U4408, P2_R1113_U111, P2_U3930);
  nand ginst16628 (P2_U4409, P2_R1131_U111, P2_U3926);
  nand ginst16629 (P2_U4410, P2_R1179_U111, P2_U3941);
  nand ginst16630 (P2_U4411, P2_R1203_U111, P2_U3943);
  nand ginst16631 (P2_U4412, P2_R1164_U111, P2_U3014);
  nand ginst16632 (P2_U4413, P2_R1233_U111, P2_U3922);
  not ginst16633 (P2_U4414, P2_U3363);
  nand ginst16634 (P2_U4415, P2_R1275_U10, P2_U3027);
  nand ginst16635 (P2_U4416, P2_U3026, P2_U3075);
  nand ginst16636 (P2_U4417, P2_R1215_U112, P2_U3025);
  nand ginst16637 (P2_U4418, P2_U3474, P2_U4116);
  nand ginst16638 (P2_U4419, P2_U3637, P2_U4414);
  nand ginst16639 (P2_U4420, P2_REG2_REG_17__SCAN_IN, P2_U3020);
  nand ginst16640 (P2_U4421, P2_REG1_REG_17__SCAN_IN, P2_U3021);
  nand ginst16641 (P2_U4422, P2_REG0_REG_17__SCAN_IN, P2_U3022);
  nand ginst16642 (P2_U4423, P2_ADD_1119_U67, P2_U3019);
  not ginst16643 (P2_U4424, P2_U3071);
  nand ginst16644 (P2_U4425, P2_U3035, P2_U3076);
  nand ginst16645 (P2_U4426, P2_R1146_U13, P2_U3931);
  nand ginst16646 (P2_U4427, P2_R1113_U13, P2_U3930);
  nand ginst16647 (P2_U4428, P2_R1131_U110, P2_U3926);
  nand ginst16648 (P2_U4429, P2_R1179_U13, P2_U3941);
  nand ginst16649 (P2_U4430, P2_R1203_U13, P2_U3943);
  nand ginst16650 (P2_U4431, P2_R1164_U110, P2_U3014);
  nand ginst16651 (P2_U4432, P2_R1233_U110, P2_U3922);
  not ginst16652 (P2_U4433, P2_U3364);
  nand ginst16653 (P2_U4434, P2_R1275_U11, P2_U3027);
  nand ginst16654 (P2_U4435, P2_U3026, P2_U3071);
  nand ginst16655 (P2_U4436, P2_R1215_U111, P2_U3025);
  nand ginst16656 (P2_U4437, P2_U3477, P2_U4116);
  nand ginst16657 (P2_U4438, P2_U3641, P2_U4433);
  nand ginst16658 (P2_U4439, P2_REG2_REG_18__SCAN_IN, P2_U3020);
  nand ginst16659 (P2_U4440, P2_REG1_REG_18__SCAN_IN, P2_U3021);
  nand ginst16660 (P2_U4441, P2_REG0_REG_18__SCAN_IN, P2_U3022);
  nand ginst16661 (P2_U4442, P2_ADD_1119_U66, P2_U3019);
  not ginst16662 (P2_U4443, P2_U3084);
  nand ginst16663 (P2_U4444, P2_U3035, P2_U3075);
  nand ginst16664 (P2_U4445, P2_R1146_U100, P2_U3931);
  nand ginst16665 (P2_U4446, P2_R1113_U100, P2_U3930);
  nand ginst16666 (P2_U4447, P2_R1131_U12, P2_U3926);
  nand ginst16667 (P2_U4448, P2_R1179_U100, P2_U3941);
  nand ginst16668 (P2_U4449, P2_R1203_U100, P2_U3943);
  nand ginst16669 (P2_U4450, P2_R1164_U12, P2_U3014);
  nand ginst16670 (P2_U4451, P2_R1233_U12, P2_U3922);
  not ginst16671 (P2_U4452, P2_U3365);
  nand ginst16672 (P2_U4453, P2_R1275_U84, P2_U3027);
  nand ginst16673 (P2_U4454, P2_U3026, P2_U3084);
  nand ginst16674 (P2_U4455, P2_R1215_U13, P2_U3025);
  nand ginst16675 (P2_U4456, P2_U3480, P2_U4116);
  nand ginst16676 (P2_U4457, P2_U3645, P2_U4452);
  nand ginst16677 (P2_U4458, P2_REG2_REG_19__SCAN_IN, P2_U3020);
  nand ginst16678 (P2_U4459, P2_REG1_REG_19__SCAN_IN, P2_U3021);
  nand ginst16679 (P2_U4460, P2_REG0_REG_19__SCAN_IN, P2_U3022);
  nand ginst16680 (P2_U4461, P2_ADD_1119_U65, P2_U3019);
  not ginst16681 (P2_U4462, P2_U3083);
  nand ginst16682 (P2_U4463, P2_U3035, P2_U3071);
  nand ginst16683 (P2_U4464, P2_R1146_U99, P2_U3931);
  nand ginst16684 (P2_U4465, P2_R1113_U99, P2_U3930);
  nand ginst16685 (P2_U4466, P2_R1131_U109, P2_U3926);
  nand ginst16686 (P2_U4467, P2_R1179_U99, P2_U3941);
  nand ginst16687 (P2_U4468, P2_R1203_U99, P2_U3943);
  nand ginst16688 (P2_U4469, P2_R1164_U109, P2_U3014);
  nand ginst16689 (P2_U4470, P2_R1233_U109, P2_U3922);
  not ginst16690 (P2_U4471, P2_U3366);
  nand ginst16691 (P2_U4472, P2_R1275_U12, P2_U3027);
  nand ginst16692 (P2_U4473, P2_U3026, P2_U3083);
  nand ginst16693 (P2_U4474, P2_R1215_U110, P2_U3025);
  nand ginst16694 (P2_U4475, P2_U3483, P2_U4116);
  nand ginst16695 (P2_U4476, P2_U3649, P2_U4471);
  nand ginst16696 (P2_U4477, P2_REG2_REG_20__SCAN_IN, P2_U3020);
  nand ginst16697 (P2_U4478, P2_REG1_REG_20__SCAN_IN, P2_U3021);
  nand ginst16698 (P2_U4479, P2_REG0_REG_20__SCAN_IN, P2_U3022);
  nand ginst16699 (P2_U4480, P2_ADD_1119_U64, P2_U3019);
  not ginst16700 (P2_U4481, P2_U3078);
  nand ginst16701 (P2_U4482, P2_U3035, P2_U3084);
  nand ginst16702 (P2_U4483, P2_R1146_U98, P2_U3931);
  nand ginst16703 (P2_U4484, P2_R1113_U98, P2_U3930);
  nand ginst16704 (P2_U4485, P2_R1131_U108, P2_U3926);
  nand ginst16705 (P2_U4486, P2_R1179_U98, P2_U3941);
  nand ginst16706 (P2_U4487, P2_R1203_U98, P2_U3943);
  nand ginst16707 (P2_U4488, P2_R1164_U108, P2_U3014);
  nand ginst16708 (P2_U4489, P2_R1233_U108, P2_U3922);
  not ginst16709 (P2_U4490, P2_U3367);
  nand ginst16710 (P2_U4491, P2_R1275_U82, P2_U3027);
  nand ginst16711 (P2_U4492, P2_U3026, P2_U3078);
  nand ginst16712 (P2_U4493, P2_R1215_U109, P2_U3025);
  nand ginst16713 (P2_U4494, P2_U3485, P2_U4116);
  nand ginst16714 (P2_U4495, P2_U3653, P2_U4490);
  nand ginst16715 (P2_U4496, P2_REG2_REG_21__SCAN_IN, P2_U3020);
  nand ginst16716 (P2_U4497, P2_REG1_REG_21__SCAN_IN, P2_U3021);
  nand ginst16717 (P2_U4498, P2_REG0_REG_21__SCAN_IN, P2_U3022);
  nand ginst16718 (P2_U4499, P2_ADD_1119_U63, P2_U3019);
  not ginst16719 (P2_U4500, P2_U3077);
  nand ginst16720 (P2_U4501, P2_U3035, P2_U3083);
  nand ginst16721 (P2_U4502, P2_R1146_U96, P2_U3931);
  nand ginst16722 (P2_U4503, P2_R1113_U96, P2_U3930);
  nand ginst16723 (P2_U4504, P2_R1131_U13, P2_U3926);
  nand ginst16724 (P2_U4505, P2_R1179_U96, P2_U3941);
  nand ginst16725 (P2_U4506, P2_R1203_U96, P2_U3943);
  nand ginst16726 (P2_U4507, P2_R1164_U13, P2_U3014);
  nand ginst16727 (P2_U4508, P2_R1233_U13, P2_U3922);
  not ginst16728 (P2_U4509, P2_U3369);
  nand ginst16729 (P2_U4510, P2_R1275_U13, P2_U3027);
  nand ginst16730 (P2_U4511, P2_U3026, P2_U3077);
  nand ginst16731 (P2_U4512, P2_R1215_U14, P2_U3025);
  nand ginst16732 (P2_U4513, P2_U3957, P2_U4116);
  nand ginst16733 (P2_U4514, P2_U3657, P2_U4509);
  nand ginst16734 (P2_U4515, P2_REG2_REG_22__SCAN_IN, P2_U3020);
  nand ginst16735 (P2_U4516, P2_REG1_REG_22__SCAN_IN, P2_U3021);
  nand ginst16736 (P2_U4517, P2_REG0_REG_22__SCAN_IN, P2_U3022);
  nand ginst16737 (P2_U4518, P2_ADD_1119_U62, P2_U3019);
  not ginst16738 (P2_U4519, P2_U3063);
  nand ginst16739 (P2_U4520, P2_U3035, P2_U3078);
  nand ginst16740 (P2_U4521, P2_R1146_U110, P2_U3931);
  nand ginst16741 (P2_U4522, P2_R1113_U110, P2_U3930);
  nand ginst16742 (P2_U4523, P2_R1131_U14, P2_U3926);
  nand ginst16743 (P2_U4524, P2_R1179_U110, P2_U3941);
  nand ginst16744 (P2_U4525, P2_R1203_U110, P2_U3943);
  nand ginst16745 (P2_U4526, P2_R1164_U14, P2_U3014);
  nand ginst16746 (P2_U4527, P2_R1233_U14, P2_U3922);
  not ginst16747 (P2_U4528, P2_U3371);
  nand ginst16748 (P2_U4529, P2_R1275_U78, P2_U3027);
  nand ginst16749 (P2_U4530, P2_U3026, P2_U3063);
  nand ginst16750 (P2_U4531, P2_R1215_U15, P2_U3025);
  nand ginst16751 (P2_U4532, P2_U3956, P2_U4116);
  nand ginst16752 (P2_U4533, P2_U3661, P2_U4528);
  nand ginst16753 (P2_U4534, P2_REG2_REG_23__SCAN_IN, P2_U3020);
  nand ginst16754 (P2_U4535, P2_REG1_REG_23__SCAN_IN, P2_U3021);
  nand ginst16755 (P2_U4536, P2_REG0_REG_23__SCAN_IN, P2_U3022);
  nand ginst16756 (P2_U4537, P2_ADD_1119_U61, P2_U3019);
  not ginst16757 (P2_U4538, P2_U3068);
  nand ginst16758 (P2_U4539, P2_U3035, P2_U3077);
  nand ginst16759 (P2_U4540, P2_R1146_U109, P2_U3931);
  nand ginst16760 (P2_U4541, P2_R1113_U109, P2_U3930);
  nand ginst16761 (P2_U4542, P2_R1131_U107, P2_U3926);
  nand ginst16762 (P2_U4543, P2_R1179_U109, P2_U3941);
  nand ginst16763 (P2_U4544, P2_R1203_U109, P2_U3943);
  nand ginst16764 (P2_U4545, P2_R1164_U107, P2_U3014);
  nand ginst16765 (P2_U4546, P2_R1233_U107, P2_U3922);
  not ginst16766 (P2_U4547, P2_U3373);
  nand ginst16767 (P2_U4548, P2_R1275_U14, P2_U3027);
  nand ginst16768 (P2_U4549, P2_U3026, P2_U3068);
  nand ginst16769 (P2_U4550, P2_R1215_U108, P2_U3025);
  nand ginst16770 (P2_U4551, P2_U3955, P2_U4116);
  nand ginst16771 (P2_U4552, P2_U3665, P2_U4547);
  nand ginst16772 (P2_U4553, P2_REG2_REG_24__SCAN_IN, P2_U3020);
  nand ginst16773 (P2_U4554, P2_REG1_REG_24__SCAN_IN, P2_U3021);
  nand ginst16774 (P2_U4555, P2_REG0_REG_24__SCAN_IN, P2_U3022);
  nand ginst16775 (P2_U4556, P2_ADD_1119_U60, P2_U3019);
  not ginst16776 (P2_U4557, P2_U3067);
  nand ginst16777 (P2_U4558, P2_U3035, P2_U3063);
  nand ginst16778 (P2_U4559, P2_R1146_U14, P2_U3931);
  nand ginst16779 (P2_U4560, P2_R1113_U14, P2_U3930);
  nand ginst16780 (P2_U4561, P2_R1131_U106, P2_U3926);
  nand ginst16781 (P2_U4562, P2_R1179_U14, P2_U3941);
  nand ginst16782 (P2_U4563, P2_R1203_U14, P2_U3943);
  nand ginst16783 (P2_U4564, P2_R1164_U106, P2_U3014);
  nand ginst16784 (P2_U4565, P2_R1233_U106, P2_U3922);
  not ginst16785 (P2_U4566, P2_U3375);
  nand ginst16786 (P2_U4567, P2_R1275_U76, P2_U3027);
  nand ginst16787 (P2_U4568, P2_U3026, P2_U3067);
  nand ginst16788 (P2_U4569, P2_R1215_U107, P2_U3025);
  nand ginst16789 (P2_U4570, P2_U3954, P2_U4116);
  nand ginst16790 (P2_U4571, P2_U3669, P2_U4566);
  nand ginst16791 (P2_U4572, P2_REG2_REG_25__SCAN_IN, P2_U3020);
  nand ginst16792 (P2_U4573, P2_REG1_REG_25__SCAN_IN, P2_U3021);
  nand ginst16793 (P2_U4574, P2_REG0_REG_25__SCAN_IN, P2_U3022);
  nand ginst16794 (P2_U4575, P2_ADD_1119_U59, P2_U3019);
  not ginst16795 (P2_U4576, P2_U3060);
  nand ginst16796 (P2_U4577, P2_U3035, P2_U3068);
  nand ginst16797 (P2_U4578, P2_R1146_U95, P2_U3931);
  nand ginst16798 (P2_U4579, P2_R1113_U95, P2_U3930);
  nand ginst16799 (P2_U4580, P2_R1131_U105, P2_U3926);
  nand ginst16800 (P2_U4581, P2_R1179_U95, P2_U3941);
  nand ginst16801 (P2_U4582, P2_R1203_U95, P2_U3943);
  nand ginst16802 (P2_U4583, P2_R1164_U105, P2_U3014);
  nand ginst16803 (P2_U4584, P2_R1233_U105, P2_U3922);
  not ginst16804 (P2_U4585, P2_U3377);
  nand ginst16805 (P2_U4586, P2_R1275_U15, P2_U3027);
  nand ginst16806 (P2_U4587, P2_U3026, P2_U3060);
  nand ginst16807 (P2_U4588, P2_R1215_U106, P2_U3025);
  nand ginst16808 (P2_U4589, P2_U3953, P2_U4116);
  nand ginst16809 (P2_U4590, P2_U3673, P2_U4585);
  nand ginst16810 (P2_U4591, P2_REG2_REG_26__SCAN_IN, P2_U3020);
  nand ginst16811 (P2_U4592, P2_REG1_REG_26__SCAN_IN, P2_U3021);
  nand ginst16812 (P2_U4593, P2_REG0_REG_26__SCAN_IN, P2_U3022);
  nand ginst16813 (P2_U4594, P2_ADD_1119_U58, P2_U3019);
  not ginst16814 (P2_U4595, P2_U3059);
  nand ginst16815 (P2_U4596, P2_U3035, P2_U3067);
  nand ginst16816 (P2_U4597, P2_R1146_U94, P2_U3931);
  nand ginst16817 (P2_U4598, P2_R1113_U94, P2_U3930);
  nand ginst16818 (P2_U4599, P2_R1131_U104, P2_U3926);
  nand ginst16819 (P2_U4600, P2_R1179_U94, P2_U3941);
  nand ginst16820 (P2_U4601, P2_R1203_U94, P2_U3943);
  nand ginst16821 (P2_U4602, P2_R1164_U104, P2_U3014);
  nand ginst16822 (P2_U4603, P2_R1233_U104, P2_U3922);
  not ginst16823 (P2_U4604, P2_U3379);
  nand ginst16824 (P2_U4605, P2_R1275_U74, P2_U3027);
  nand ginst16825 (P2_U4606, P2_U3026, P2_U3059);
  nand ginst16826 (P2_U4607, P2_R1215_U105, P2_U3025);
  nand ginst16827 (P2_U4608, P2_U3952, P2_U4116);
  nand ginst16828 (P2_U4609, P2_U3677, P2_U4604);
  nand ginst16829 (P2_U4610, P2_REG2_REG_27__SCAN_IN, P2_U3020);
  nand ginst16830 (P2_U4611, P2_REG1_REG_27__SCAN_IN, P2_U3021);
  nand ginst16831 (P2_U4612, P2_REG0_REG_27__SCAN_IN, P2_U3022);
  nand ginst16832 (P2_U4613, P2_ADD_1119_U57, P2_U3019);
  not ginst16833 (P2_U4614, P2_U3055);
  nand ginst16834 (P2_U4615, P2_U3035, P2_U3060);
  nand ginst16835 (P2_U4616, P2_R1146_U108, P2_U3931);
  nand ginst16836 (P2_U4617, P2_R1113_U108, P2_U3930);
  nand ginst16837 (P2_U4618, P2_R1131_U15, P2_U3926);
  nand ginst16838 (P2_U4619, P2_R1179_U108, P2_U3941);
  nand ginst16839 (P2_U4620, P2_R1203_U108, P2_U3943);
  nand ginst16840 (P2_U4621, P2_R1164_U15, P2_U3014);
  nand ginst16841 (P2_U4622, P2_R1233_U15, P2_U3922);
  not ginst16842 (P2_U4623, P2_U3381);
  nand ginst16843 (P2_U4624, P2_R1275_U16, P2_U3027);
  nand ginst16844 (P2_U4625, P2_U3026, P2_U3055);
  nand ginst16845 (P2_U4626, P2_R1215_U16, P2_U3025);
  nand ginst16846 (P2_U4627, P2_U3951, P2_U4116);
  nand ginst16847 (P2_U4628, P2_U3681, P2_U4623);
  nand ginst16848 (P2_U4629, P2_REG2_REG_28__SCAN_IN, P2_U3020);
  nand ginst16849 (P2_U4630, P2_REG1_REG_28__SCAN_IN, P2_U3021);
  nand ginst16850 (P2_U4631, P2_REG0_REG_28__SCAN_IN, P2_U3022);
  nand ginst16851 (P2_U4632, P2_ADD_1119_U56, P2_U3019);
  not ginst16852 (P2_U4633, P2_U3056);
  nand ginst16853 (P2_U4634, P2_U3035, P2_U3059);
  nand ginst16854 (P2_U4635, P2_R1146_U15, P2_U3931);
  nand ginst16855 (P2_U4636, P2_R1113_U15, P2_U3930);
  nand ginst16856 (P2_U4637, P2_R1131_U103, P2_U3926);
  nand ginst16857 (P2_U4638, P2_R1179_U15, P2_U3941);
  nand ginst16858 (P2_U4639, P2_R1203_U15, P2_U3943);
  nand ginst16859 (P2_U4640, P2_R1164_U103, P2_U3014);
  nand ginst16860 (P2_U4641, P2_R1233_U103, P2_U3922);
  not ginst16861 (P2_U4642, P2_U3383);
  nand ginst16862 (P2_U4643, P2_R1275_U72, P2_U3027);
  nand ginst16863 (P2_U4644, P2_U3026, P2_U3056);
  nand ginst16864 (P2_U4645, P2_R1215_U104, P2_U3025);
  nand ginst16865 (P2_U4646, P2_U3950, P2_U4116);
  nand ginst16866 (P2_U4647, P2_U3685, P2_U4642);
  nand ginst16867 (P2_U4648, P2_ADD_1119_U5, P2_U3019);
  nand ginst16868 (P2_U4649, P2_REG2_REG_29__SCAN_IN, P2_U3020);
  nand ginst16869 (P2_U4650, P2_REG1_REG_29__SCAN_IN, P2_U3021);
  nand ginst16870 (P2_U4651, P2_REG0_REG_29__SCAN_IN, P2_U3022);
  not ginst16871 (P2_U4652, P2_U3057);
  nand ginst16872 (P2_U4653, P2_U3035, P2_U3055);
  nand ginst16873 (P2_U4654, P2_R1146_U93, P2_U3931);
  nand ginst16874 (P2_U4655, P2_R1113_U93, P2_U3930);
  nand ginst16875 (P2_U4656, P2_R1131_U102, P2_U3926);
  nand ginst16876 (P2_U4657, P2_R1179_U93, P2_U3941);
  nand ginst16877 (P2_U4658, P2_R1203_U93, P2_U3943);
  nand ginst16878 (P2_U4659, P2_R1164_U102, P2_U3014);
  nand ginst16879 (P2_U4660, P2_R1233_U102, P2_U3922);
  not ginst16880 (P2_U4661, P2_U3385);
  nand ginst16881 (P2_U4662, P2_R1275_U17, P2_U3027);
  nand ginst16882 (P2_U4663, P2_U3026, P2_U3057);
  nand ginst16883 (P2_U4664, P2_R1215_U103, P2_U3025);
  nand ginst16884 (P2_U4665, P2_U3949, P2_U4116);
  nand ginst16885 (P2_U4666, P2_U3688, P2_U4661);
  nand ginst16886 (P2_U4667, P2_REG2_REG_30__SCAN_IN, P2_U3020);
  nand ginst16887 (P2_U4668, P2_REG1_REG_30__SCAN_IN, P2_U3021);
  nand ginst16888 (P2_U4669, P2_REG0_REG_30__SCAN_IN, P2_U3022);
  not ginst16889 (P2_U4670, P2_U3061);
  nand ginst16890 (P2_U4671, P2_U3331, P2_U5683);
  nand ginst16891 (P2_U4672, P2_U3347, P2_U4671);
  nand ginst16892 (P2_U4673, P2_U3061, P2_U3689);
  nand ginst16893 (P2_U4674, P2_U3035, P2_U3056);
  nand ginst16894 (P2_U4675, P2_R1146_U16, P2_U3931);
  nand ginst16895 (P2_U4676, P2_R1113_U16, P2_U3930);
  nand ginst16896 (P2_U4677, P2_R1131_U101, P2_U3926);
  nand ginst16897 (P2_U4678, P2_R1179_U16, P2_U3941);
  nand ginst16898 (P2_U4679, P2_R1203_U16, P2_U3943);
  nand ginst16899 (P2_U4680, P2_R1164_U101, P2_U3014);
  nand ginst16900 (P2_U4681, P2_R1233_U101, P2_U3922);
  not ginst16901 (P2_U4682, P2_U3387);
  nand ginst16902 (P2_U4683, P2_R1275_U70, P2_U3027);
  nand ginst16903 (P2_U4684, P2_R1215_U102, P2_U3025);
  nand ginst16904 (P2_U4685, P2_U3960, P2_U4116);
  nand ginst16905 (P2_U4686, P2_U3693, P2_U4682);
  nand ginst16906 (P2_U4687, P2_REG2_REG_31__SCAN_IN, P2_U3020);
  nand ginst16907 (P2_U4688, P2_REG1_REG_31__SCAN_IN, P2_U3021);
  nand ginst16908 (P2_U4689, P2_REG0_REG_31__SCAN_IN, P2_U3022);
  not ginst16909 (P2_U4690, P2_U3058);
  nand ginst16910 (P2_U4691, P2_R1275_U19, P2_U3027);
  nand ginst16911 (P2_U4692, P2_U3959, P2_U4116);
  nand ginst16912 (P2_U4693, P2_U3913, P2_U4691, P2_U4692);
  nand ginst16913 (P2_U4694, P2_R1275_U68, P2_U3027);
  nand ginst16914 (P2_U4695, P2_U3958, P2_U4116);
  nand ginst16915 (P2_U4696, P2_U3913, P2_U4694, P2_U4695);
  nand ginst16916 (P2_U4697, P2_U3016, P2_U3696);
  nand ginst16917 (P2_U4698, P2_U3393, P2_U4697);
  nand ginst16918 (P2_U4699, P2_U3418, P2_U3921);
  not ginst16919 (P2_U4700, P2_U3398);
  nand ginst16920 (P2_U4701, P2_U3037, P2_U3080);
  nand ginst16921 (P2_U4702, P2_R1215_U96, P2_U3034);
  nand ginst16922 (P2_U4703, P2_REG3_REG_0__SCAN_IN, P2_U3033);
  nand ginst16923 (P2_U4704, P2_U3032, P2_U3427);
  nand ginst16924 (P2_U4705, P2_U3031, P2_U3427);
  nand ginst16925 (P2_U4706, P2_U3037, P2_U3070);
  nand ginst16926 (P2_U4707, P2_R1215_U95, P2_U3034);
  nand ginst16927 (P2_U4708, P2_REG3_REG_1__SCAN_IN, P2_U3033);
  nand ginst16928 (P2_U4709, P2_U3032, P2_U3432);
  nand ginst16929 (P2_U4710, P2_R1275_U55, P2_U3031);
  nand ginst16930 (P2_U4711, P2_U3037, P2_U3066);
  nand ginst16931 (P2_U4712, P2_R1215_U17, P2_U3034);
  nand ginst16932 (P2_U4713, P2_REG3_REG_2__SCAN_IN, P2_U3033);
  nand ginst16933 (P2_U4714, P2_U3032, P2_U3435);
  nand ginst16934 (P2_U4715, P2_R1275_U18, P2_U3031);
  nand ginst16935 (P2_U4716, P2_U3037, P2_U3062);
  nand ginst16936 (P2_U4717, P2_R1215_U101, P2_U3034);
  nand ginst16937 (P2_U4718, P2_ADD_1119_U4, P2_U3033);
  nand ginst16938 (P2_U4719, P2_U3032, P2_U3438);
  nand ginst16939 (P2_U4720, P2_R1275_U20, P2_U3031);
  nand ginst16940 (P2_U4721, P2_U3037, P2_U3069);
  nand ginst16941 (P2_U4722, P2_R1215_U100, P2_U3034);
  nand ginst16942 (P2_U4723, P2_ADD_1119_U55, P2_U3033);
  nand ginst16943 (P2_U4724, P2_U3032, P2_U3441);
  nand ginst16944 (P2_U4725, P2_R1275_U21, P2_U3031);
  nand ginst16945 (P2_U4726, P2_U3037, P2_U3073);
  nand ginst16946 (P2_U4727, P2_R1215_U18, P2_U3034);
  nand ginst16947 (P2_U4728, P2_ADD_1119_U54, P2_U3033);
  nand ginst16948 (P2_U4729, P2_U3032, P2_U3444);
  nand ginst16949 (P2_U4730, P2_R1275_U65, P2_U3031);
  nand ginst16950 (P2_U4731, P2_U3037, P2_U3072);
  nand ginst16951 (P2_U4732, P2_R1215_U99, P2_U3034);
  nand ginst16952 (P2_U4733, P2_ADD_1119_U53, P2_U3033);
  nand ginst16953 (P2_U4734, P2_U3032, P2_U3447);
  nand ginst16954 (P2_U4735, P2_R1275_U22, P2_U3031);
  nand ginst16955 (P2_U4736, P2_U3037, P2_U3086);
  nand ginst16956 (P2_U4737, P2_R1215_U19, P2_U3034);
  nand ginst16957 (P2_U4738, P2_ADD_1119_U52, P2_U3033);
  nand ginst16958 (P2_U4739, P2_U3032, P2_U3450);
  nand ginst16959 (P2_U4740, P2_R1275_U23, P2_U3031);
  nand ginst16960 (P2_U4741, P2_U3037, P2_U3085);
  nand ginst16961 (P2_U4742, P2_R1215_U98, P2_U3034);
  nand ginst16962 (P2_U4743, P2_ADD_1119_U51, P2_U3033);
  nand ginst16963 (P2_U4744, P2_U3032, P2_U3453);
  nand ginst16964 (P2_U4745, P2_R1275_U24, P2_U3031);
  nand ginst16965 (P2_U4746, P2_U3037, P2_U3064);
  nand ginst16966 (P2_U4747, P2_R1215_U97, P2_U3034);
  nand ginst16967 (P2_U4748, P2_ADD_1119_U50, P2_U3033);
  nand ginst16968 (P2_U4749, P2_U3032, P2_U3456);
  nand ginst16969 (P2_U4750, P2_R1275_U63, P2_U3031);
  nand ginst16970 (P2_U4751, P2_U3037, P2_U3065);
  nand ginst16971 (P2_U4752, P2_R1215_U11, P2_U3034);
  nand ginst16972 (P2_U4753, P2_ADD_1119_U74, P2_U3033);
  nand ginst16973 (P2_U4754, P2_U3032, P2_U3459);
  nand ginst16974 (P2_U4755, P2_R1275_U6, P2_U3031);
  nand ginst16975 (P2_U4756, P2_U3037, P2_U3074);
  nand ginst16976 (P2_U4757, P2_R1215_U115, P2_U3034);
  nand ginst16977 (P2_U4758, P2_ADD_1119_U73, P2_U3033);
  nand ginst16978 (P2_U4759, P2_U3032, P2_U3462);
  nand ginst16979 (P2_U4760, P2_R1275_U7, P2_U3031);
  nand ginst16980 (P2_U4761, P2_U3037, P2_U3082);
  nand ginst16981 (P2_U4762, P2_R1215_U114, P2_U3034);
  nand ginst16982 (P2_U4763, P2_ADD_1119_U72, P2_U3033);
  nand ginst16983 (P2_U4764, P2_U3032, P2_U3465);
  nand ginst16984 (P2_U4765, P2_R1275_U8, P2_U3031);
  nand ginst16985 (P2_U4766, P2_U3037, P2_U3081);
  nand ginst16986 (P2_U4767, P2_R1215_U12, P2_U3034);
  nand ginst16987 (P2_U4768, P2_ADD_1119_U71, P2_U3033);
  nand ginst16988 (P2_U4769, P2_U3032, P2_U3468);
  nand ginst16989 (P2_U4770, P2_R1275_U86, P2_U3031);
  nand ginst16990 (P2_U4771, P2_U3037, P2_U3076);
  nand ginst16991 (P2_U4772, P2_R1215_U113, P2_U3034);
  nand ginst16992 (P2_U4773, P2_ADD_1119_U70, P2_U3033);
  nand ginst16993 (P2_U4774, P2_U3032, P2_U3471);
  nand ginst16994 (P2_U4775, P2_R1275_U9, P2_U3031);
  nand ginst16995 (P2_U4776, P2_U3037, P2_U3075);
  nand ginst16996 (P2_U4777, P2_R1215_U112, P2_U3034);
  nand ginst16997 (P2_U4778, P2_ADD_1119_U69, P2_U3033);
  nand ginst16998 (P2_U4779, P2_U3032, P2_U3474);
  nand ginst16999 (P2_U4780, P2_R1275_U10, P2_U3031);
  nand ginst17000 (P2_U4781, P2_U3037, P2_U3071);
  nand ginst17001 (P2_U4782, P2_R1215_U111, P2_U3034);
  nand ginst17002 (P2_U4783, P2_ADD_1119_U68, P2_U3033);
  nand ginst17003 (P2_U4784, P2_U3032, P2_U3477);
  nand ginst17004 (P2_U4785, P2_R1275_U11, P2_U3031);
  nand ginst17005 (P2_U4786, P2_U3037, P2_U3084);
  nand ginst17006 (P2_U4787, P2_R1215_U13, P2_U3034);
  nand ginst17007 (P2_U4788, P2_ADD_1119_U67, P2_U3033);
  nand ginst17008 (P2_U4789, P2_U3032, P2_U3480);
  nand ginst17009 (P2_U4790, P2_R1275_U84, P2_U3031);
  nand ginst17010 (P2_U4791, P2_U3037, P2_U3083);
  nand ginst17011 (P2_U4792, P2_R1215_U110, P2_U3034);
  nand ginst17012 (P2_U4793, P2_ADD_1119_U66, P2_U3033);
  nand ginst17013 (P2_U4794, P2_U3032, P2_U3483);
  nand ginst17014 (P2_U4795, P2_R1275_U12, P2_U3031);
  nand ginst17015 (P2_U4796, P2_U3037, P2_U3078);
  nand ginst17016 (P2_U4797, P2_R1215_U109, P2_U3034);
  nand ginst17017 (P2_U4798, P2_ADD_1119_U65, P2_U3033);
  nand ginst17018 (P2_U4799, P2_U3032, P2_U3485);
  nand ginst17019 (P2_U4800, P2_R1275_U82, P2_U3031);
  nand ginst17020 (P2_U4801, P2_U3037, P2_U3077);
  nand ginst17021 (P2_U4802, P2_R1215_U14, P2_U3034);
  nand ginst17022 (P2_U4803, P2_ADD_1119_U64, P2_U3033);
  nand ginst17023 (P2_U4804, P2_U3032, P2_U3957);
  nand ginst17024 (P2_U4805, P2_R1275_U13, P2_U3031);
  nand ginst17025 (P2_U4806, P2_U3037, P2_U3063);
  nand ginst17026 (P2_U4807, P2_R1215_U15, P2_U3034);
  nand ginst17027 (P2_U4808, P2_ADD_1119_U63, P2_U3033);
  nand ginst17028 (P2_U4809, P2_U3032, P2_U3956);
  nand ginst17029 (P2_U4810, P2_R1275_U78, P2_U3031);
  nand ginst17030 (P2_U4811, P2_U3037, P2_U3068);
  nand ginst17031 (P2_U4812, P2_R1215_U108, P2_U3034);
  nand ginst17032 (P2_U4813, P2_ADD_1119_U62, P2_U3033);
  nand ginst17033 (P2_U4814, P2_U3032, P2_U3955);
  nand ginst17034 (P2_U4815, P2_R1275_U14, P2_U3031);
  nand ginst17035 (P2_U4816, P2_U3037, P2_U3067);
  nand ginst17036 (P2_U4817, P2_R1215_U107, P2_U3034);
  nand ginst17037 (P2_U4818, P2_ADD_1119_U61, P2_U3033);
  nand ginst17038 (P2_U4819, P2_U3032, P2_U3954);
  nand ginst17039 (P2_U4820, P2_R1275_U76, P2_U3031);
  nand ginst17040 (P2_U4821, P2_U3037, P2_U3060);
  nand ginst17041 (P2_U4822, P2_R1215_U106, P2_U3034);
  nand ginst17042 (P2_U4823, P2_ADD_1119_U60, P2_U3033);
  nand ginst17043 (P2_U4824, P2_U3032, P2_U3953);
  nand ginst17044 (P2_U4825, P2_R1275_U15, P2_U3031);
  nand ginst17045 (P2_U4826, P2_U3037, P2_U3059);
  nand ginst17046 (P2_U4827, P2_R1215_U105, P2_U3034);
  nand ginst17047 (P2_U4828, P2_ADD_1119_U59, P2_U3033);
  nand ginst17048 (P2_U4829, P2_U3032, P2_U3952);
  nand ginst17049 (P2_U4830, P2_R1275_U74, P2_U3031);
  nand ginst17050 (P2_U4831, P2_U3037, P2_U3055);
  nand ginst17051 (P2_U4832, P2_R1215_U16, P2_U3034);
  nand ginst17052 (P2_U4833, P2_ADD_1119_U58, P2_U3033);
  nand ginst17053 (P2_U4834, P2_U3032, P2_U3951);
  nand ginst17054 (P2_U4835, P2_R1275_U16, P2_U3031);
  nand ginst17055 (P2_U4836, P2_U3037, P2_U3056);
  nand ginst17056 (P2_U4837, P2_R1215_U104, P2_U3034);
  nand ginst17057 (P2_U4838, P2_ADD_1119_U57, P2_U3033);
  nand ginst17058 (P2_U4839, P2_U3032, P2_U3950);
  nand ginst17059 (P2_U4840, P2_R1275_U72, P2_U3031);
  nand ginst17060 (P2_U4841, P2_U3037, P2_U3057);
  nand ginst17061 (P2_U4842, P2_R1215_U103, P2_U3034);
  nand ginst17062 (P2_U4843, P2_ADD_1119_U56, P2_U3033);
  nand ginst17063 (P2_U4844, P2_U3032, P2_U3949);
  nand ginst17064 (P2_U4845, P2_R1275_U17, P2_U3031);
  nand ginst17065 (P2_U4846, P2_R1215_U102, P2_U3034);
  nand ginst17066 (P2_U4847, P2_ADD_1119_U5, P2_U3033);
  nand ginst17067 (P2_U4848, P2_U3032, P2_U3960);
  nand ginst17068 (P2_U4849, P2_R1275_U70, P2_U3031);
  nand ginst17069 (P2_U4850, P2_U3032, P2_U3959);
  nand ginst17070 (P2_U4851, P2_R1275_U19, P2_U3031);
  nand ginst17071 (P2_U4852, P2_U3032, P2_U3958);
  nand ginst17072 (P2_U4853, P2_R1275_U68, P2_U3031);
  nand ginst17073 (P2_U4854, P2_U3051, P2_U3393, P2_U3395, P2_U3755, P2_U4700);
  nand ginst17074 (P2_U4855, P2_R1170_U13, P2_U3043);
  nand ginst17075 (P2_U4856, P2_U3041, P2_U3424);
  nand ginst17076 (P2_U4857, P2_R1209_U13, P2_U3039);
  nand ginst17077 (P2_U4858, P2_U4855, P2_U4856, P2_U4857);
  nand ginst17078 (P2_U4859, P2_R1170_U13, P2_U3018);
  nand ginst17079 (P2_U4860, P2_R1209_U13, P2_U3017);
  nand ginst17080 (P2_U4861, P2_U3424, P2_U5683);
  nand ginst17081 (P2_U4862, P2_U4859, P2_U4860, P2_U4861);
  not ginst17082 (P2_U4863, P2_U3401);
  nand ginst17083 (P2_U4864, P2_U3045, P2_U4858);
  nand ginst17084 (P2_U4865, P2_U3947, P2_U4862);
  nand ginst17085 (P2_U4866, P2_R1170_U13, P2_U3044);
  nand ginst17086 (P2_U4867, P2_REG3_REG_19__SCAN_IN, P2_U3088);
  nand ginst17087 (P2_U4868, P2_U3042, P2_U3424);
  nand ginst17088 (P2_U4869, P2_R1209_U13, P2_U3040);
  nand ginst17089 (P2_U4870, P2_ADDR_REG_19__SCAN_IN, P2_U4863);
  nand ginst17090 (P2_U4871, P2_R1170_U75, P2_U3043);
  nand ginst17091 (P2_U4872, P2_U3041, P2_U3482);
  nand ginst17092 (P2_U4873, P2_R1209_U75, P2_U3039);
  nand ginst17093 (P2_U4874, P2_U4871, P2_U4872, P2_U4873);
  nand ginst17094 (P2_U4875, P2_R1170_U75, P2_U3018);
  nand ginst17095 (P2_U4876, P2_R1209_U75, P2_U3017);
  nand ginst17096 (P2_U4877, P2_U3482, P2_U5683);
  nand ginst17097 (P2_U4878, P2_U4875, P2_U4876, P2_U4877);
  nand ginst17098 (P2_U4879, P2_U3045, P2_U4874);
  nand ginst17099 (P2_U4880, P2_U3947, P2_U4878);
  nand ginst17100 (P2_U4881, P2_R1170_U75, P2_U3044);
  nand ginst17101 (P2_U4882, P2_REG3_REG_18__SCAN_IN, P2_U3088);
  nand ginst17102 (P2_U4883, P2_U3042, P2_U3482);
  nand ginst17103 (P2_U4884, P2_R1209_U75, P2_U3040);
  nand ginst17104 (P2_U4885, P2_ADDR_REG_18__SCAN_IN, P2_U4863);
  nand ginst17105 (P2_U4886, P2_R1170_U12, P2_U3043);
  nand ginst17106 (P2_U4887, P2_U3041, P2_U3479);
  nand ginst17107 (P2_U4888, P2_R1209_U12, P2_U3039);
  nand ginst17108 (P2_U4889, P2_U4886, P2_U4887, P2_U4888);
  nand ginst17109 (P2_U4890, P2_R1170_U12, P2_U3018);
  nand ginst17110 (P2_U4891, P2_R1209_U12, P2_U3017);
  nand ginst17111 (P2_U4892, P2_U3479, P2_U5683);
  nand ginst17112 (P2_U4893, P2_U4890, P2_U4891, P2_U4892);
  nand ginst17113 (P2_U4894, P2_U3045, P2_U4889);
  nand ginst17114 (P2_U4895, P2_U3947, P2_U4893);
  nand ginst17115 (P2_U4896, P2_R1170_U12, P2_U3044);
  nand ginst17116 (P2_U4897, P2_REG3_REG_17__SCAN_IN, P2_U3088);
  nand ginst17117 (P2_U4898, P2_U3042, P2_U3479);
  nand ginst17118 (P2_U4899, P2_R1209_U12, P2_U3040);
  nand ginst17119 (P2_U4900, P2_ADDR_REG_17__SCAN_IN, P2_U4863);
  nand ginst17120 (P2_U4901, P2_R1170_U76, P2_U3043);
  nand ginst17121 (P2_U4902, P2_U3041, P2_U3476);
  nand ginst17122 (P2_U4903, P2_R1209_U76, P2_U3039);
  nand ginst17123 (P2_U4904, P2_U4901, P2_U4902, P2_U4903);
  nand ginst17124 (P2_U4905, P2_R1170_U76, P2_U3018);
  nand ginst17125 (P2_U4906, P2_R1209_U76, P2_U3017);
  nand ginst17126 (P2_U4907, P2_U3476, P2_U5683);
  nand ginst17127 (P2_U4908, P2_U4905, P2_U4906, P2_U4907);
  nand ginst17128 (P2_U4909, P2_U3045, P2_U4904);
  nand ginst17129 (P2_U4910, P2_U3947, P2_U4908);
  nand ginst17130 (P2_U4911, P2_R1170_U76, P2_U3044);
  nand ginst17131 (P2_U4912, P2_REG3_REG_16__SCAN_IN, P2_U3088);
  nand ginst17132 (P2_U4913, P2_U3042, P2_U3476);
  nand ginst17133 (P2_U4914, P2_R1209_U76, P2_U3040);
  nand ginst17134 (P2_U4915, P2_ADDR_REG_16__SCAN_IN, P2_U4863);
  nand ginst17135 (P2_U4916, P2_R1170_U77, P2_U3043);
  nand ginst17136 (P2_U4917, P2_U3041, P2_U3473);
  nand ginst17137 (P2_U4918, P2_R1209_U77, P2_U3039);
  nand ginst17138 (P2_U4919, P2_U4916, P2_U4917, P2_U4918);
  nand ginst17139 (P2_U4920, P2_R1170_U77, P2_U3018);
  nand ginst17140 (P2_U4921, P2_R1209_U77, P2_U3017);
  nand ginst17141 (P2_U4922, P2_U3473, P2_U5683);
  nand ginst17142 (P2_U4923, P2_U4920, P2_U4921, P2_U4922);
  nand ginst17143 (P2_U4924, P2_U3045, P2_U4919);
  nand ginst17144 (P2_U4925, P2_U3947, P2_U4923);
  nand ginst17145 (P2_U4926, P2_R1170_U77, P2_U3044);
  nand ginst17146 (P2_U4927, P2_REG3_REG_15__SCAN_IN, P2_U3088);
  nand ginst17147 (P2_U4928, P2_U3042, P2_U3473);
  nand ginst17148 (P2_U4929, P2_R1209_U77, P2_U3040);
  nand ginst17149 (P2_U4930, P2_ADDR_REG_15__SCAN_IN, P2_U4863);
  nand ginst17150 (P2_U4931, P2_R1170_U78, P2_U3043);
  nand ginst17151 (P2_U4932, P2_U3041, P2_U3470);
  nand ginst17152 (P2_U4933, P2_R1209_U78, P2_U3039);
  nand ginst17153 (P2_U4934, P2_U4931, P2_U4932, P2_U4933);
  nand ginst17154 (P2_U4935, P2_R1170_U78, P2_U3018);
  nand ginst17155 (P2_U4936, P2_R1209_U78, P2_U3017);
  nand ginst17156 (P2_U4937, P2_U3470, P2_U5683);
  nand ginst17157 (P2_U4938, P2_U4935, P2_U4936, P2_U4937);
  nand ginst17158 (P2_U4939, P2_U3045, P2_U4934);
  nand ginst17159 (P2_U4940, P2_U3947, P2_U4938);
  nand ginst17160 (P2_U4941, P2_R1170_U78, P2_U3044);
  nand ginst17161 (P2_U4942, P2_REG3_REG_14__SCAN_IN, P2_U3088);
  nand ginst17162 (P2_U4943, P2_U3042, P2_U3470);
  nand ginst17163 (P2_U4944, P2_R1209_U78, P2_U3040);
  nand ginst17164 (P2_U4945, P2_ADDR_REG_14__SCAN_IN, P2_U4863);
  nand ginst17165 (P2_U4946, P2_R1170_U11, P2_U3043);
  nand ginst17166 (P2_U4947, P2_U3041, P2_U3467);
  nand ginst17167 (P2_U4948, P2_R1209_U11, P2_U3039);
  nand ginst17168 (P2_U4949, P2_U4946, P2_U4947, P2_U4948);
  nand ginst17169 (P2_U4950, P2_R1170_U11, P2_U3018);
  nand ginst17170 (P2_U4951, P2_R1209_U11, P2_U3017);
  nand ginst17171 (P2_U4952, P2_U3467, P2_U5683);
  nand ginst17172 (P2_U4953, P2_U4950, P2_U4951, P2_U4952);
  nand ginst17173 (P2_U4954, P2_U3045, P2_U4949);
  nand ginst17174 (P2_U4955, P2_U3947, P2_U4953);
  nand ginst17175 (P2_U4956, P2_R1170_U11, P2_U3044);
  nand ginst17176 (P2_U4957, P2_REG3_REG_13__SCAN_IN, P2_U3088);
  nand ginst17177 (P2_U4958, P2_U3042, P2_U3467);
  nand ginst17178 (P2_U4959, P2_R1209_U11, P2_U3040);
  nand ginst17179 (P2_U4960, P2_ADDR_REG_13__SCAN_IN, P2_U4863);
  nand ginst17180 (P2_U4961, P2_R1170_U79, P2_U3043);
  nand ginst17181 (P2_U4962, P2_U3041, P2_U3464);
  nand ginst17182 (P2_U4963, P2_R1209_U79, P2_U3039);
  nand ginst17183 (P2_U4964, P2_U4961, P2_U4962, P2_U4963);
  nand ginst17184 (P2_U4965, P2_R1170_U79, P2_U3018);
  nand ginst17185 (P2_U4966, P2_R1209_U79, P2_U3017);
  nand ginst17186 (P2_U4967, P2_U3464, P2_U5683);
  nand ginst17187 (P2_U4968, P2_U4965, P2_U4966, P2_U4967);
  nand ginst17188 (P2_U4969, P2_U3045, P2_U4964);
  nand ginst17189 (P2_U4970, P2_U3947, P2_U4968);
  nand ginst17190 (P2_U4971, P2_R1170_U79, P2_U3044);
  nand ginst17191 (P2_U4972, P2_REG3_REG_12__SCAN_IN, P2_U3088);
  nand ginst17192 (P2_U4973, P2_U3042, P2_U3464);
  nand ginst17193 (P2_U4974, P2_R1209_U79, P2_U3040);
  nand ginst17194 (P2_U4975, P2_ADDR_REG_12__SCAN_IN, P2_U4863);
  nand ginst17195 (P2_U4976, P2_R1170_U80, P2_U3043);
  nand ginst17196 (P2_U4977, P2_U3041, P2_U3461);
  nand ginst17197 (P2_U4978, P2_R1209_U80, P2_U3039);
  nand ginst17198 (P2_U4979, P2_U4976, P2_U4977, P2_U4978);
  nand ginst17199 (P2_U4980, P2_R1170_U80, P2_U3018);
  nand ginst17200 (P2_U4981, P2_R1209_U80, P2_U3017);
  nand ginst17201 (P2_U4982, P2_U3461, P2_U5683);
  nand ginst17202 (P2_U4983, P2_U4980, P2_U4981, P2_U4982);
  nand ginst17203 (P2_U4984, P2_U3045, P2_U4979);
  nand ginst17204 (P2_U4985, P2_U3947, P2_U4983);
  nand ginst17205 (P2_U4986, P2_R1170_U80, P2_U3044);
  nand ginst17206 (P2_U4987, P2_REG3_REG_11__SCAN_IN, P2_U3088);
  nand ginst17207 (P2_U4988, P2_U3042, P2_U3461);
  nand ginst17208 (P2_U4989, P2_R1209_U80, P2_U3040);
  nand ginst17209 (P2_U4990, P2_ADDR_REG_11__SCAN_IN, P2_U4863);
  nand ginst17210 (P2_U4991, P2_R1170_U10, P2_U3043);
  nand ginst17211 (P2_U4992, P2_U3041, P2_U3458);
  nand ginst17212 (P2_U4993, P2_R1209_U10, P2_U3039);
  nand ginst17213 (P2_U4994, P2_U4991, P2_U4992, P2_U4993);
  nand ginst17214 (P2_U4995, P2_R1170_U10, P2_U3018);
  nand ginst17215 (P2_U4996, P2_R1209_U10, P2_U3017);
  nand ginst17216 (P2_U4997, P2_U3458, P2_U5683);
  nand ginst17217 (P2_U4998, P2_U4995, P2_U4996, P2_U4997);
  nand ginst17218 (P2_U4999, P2_U3045, P2_U4994);
  nand ginst17219 (P2_U5000, P2_U3947, P2_U4998);
  nand ginst17220 (P2_U5001, P2_R1170_U10, P2_U3044);
  nand ginst17221 (P2_U5002, P2_REG3_REG_10__SCAN_IN, P2_U3088);
  nand ginst17222 (P2_U5003, P2_U3042, P2_U3458);
  nand ginst17223 (P2_U5004, P2_R1209_U10, P2_U3040);
  nand ginst17224 (P2_U5005, P2_ADDR_REG_10__SCAN_IN, P2_U4863);
  nand ginst17225 (P2_U5006, P2_R1170_U70, P2_U3043);
  nand ginst17226 (P2_U5007, P2_U3041, P2_U3455);
  nand ginst17227 (P2_U5008, P2_R1209_U70, P2_U3039);
  nand ginst17228 (P2_U5009, P2_U5006, P2_U5007, P2_U5008);
  nand ginst17229 (P2_U5010, P2_R1170_U70, P2_U3018);
  nand ginst17230 (P2_U5011, P2_R1209_U70, P2_U3017);
  nand ginst17231 (P2_U5012, P2_U3455, P2_U5683);
  nand ginst17232 (P2_U5013, P2_U5010, P2_U5011, P2_U5012);
  nand ginst17233 (P2_U5014, P2_U3045, P2_U5009);
  nand ginst17234 (P2_U5015, P2_U3947, P2_U5013);
  nand ginst17235 (P2_U5016, P2_R1170_U70, P2_U3044);
  nand ginst17236 (P2_U5017, P2_REG3_REG_9__SCAN_IN, P2_U3088);
  nand ginst17237 (P2_U5018, P2_U3042, P2_U3455);
  nand ginst17238 (P2_U5019, P2_R1209_U70, P2_U3040);
  nand ginst17239 (P2_U5020, P2_ADDR_REG_9__SCAN_IN, P2_U4863);
  nand ginst17240 (P2_U5021, P2_R1170_U71, P2_U3043);
  nand ginst17241 (P2_U5022, P2_U3041, P2_U3452);
  nand ginst17242 (P2_U5023, P2_R1209_U71, P2_U3039);
  nand ginst17243 (P2_U5024, P2_U5021, P2_U5022, P2_U5023);
  nand ginst17244 (P2_U5025, P2_R1170_U71, P2_U3018);
  nand ginst17245 (P2_U5026, P2_R1209_U71, P2_U3017);
  nand ginst17246 (P2_U5027, P2_U3452, P2_U5683);
  nand ginst17247 (P2_U5028, P2_U5025, P2_U5026, P2_U5027);
  nand ginst17248 (P2_U5029, P2_U3045, P2_U5024);
  nand ginst17249 (P2_U5030, P2_U3947, P2_U5028);
  nand ginst17250 (P2_U5031, P2_R1170_U71, P2_U3044);
  nand ginst17251 (P2_U5032, P2_REG3_REG_8__SCAN_IN, P2_U3088);
  nand ginst17252 (P2_U5033, P2_U3042, P2_U3452);
  nand ginst17253 (P2_U5034, P2_R1209_U71, P2_U3040);
  nand ginst17254 (P2_U5035, P2_ADDR_REG_8__SCAN_IN, P2_U4863);
  nand ginst17255 (P2_U5036, P2_R1170_U16, P2_U3043);
  nand ginst17256 (P2_U5037, P2_U3041, P2_U3449);
  nand ginst17257 (P2_U5038, P2_R1209_U16, P2_U3039);
  nand ginst17258 (P2_U5039, P2_U5036, P2_U5037, P2_U5038);
  nand ginst17259 (P2_U5040, P2_R1170_U16, P2_U3018);
  nand ginst17260 (P2_U5041, P2_R1209_U16, P2_U3017);
  nand ginst17261 (P2_U5042, P2_U3449, P2_U5683);
  nand ginst17262 (P2_U5043, P2_U5040, P2_U5041, P2_U5042);
  nand ginst17263 (P2_U5044, P2_U3045, P2_U5039);
  nand ginst17264 (P2_U5045, P2_U3947, P2_U5043);
  nand ginst17265 (P2_U5046, P2_R1170_U16, P2_U3044);
  nand ginst17266 (P2_U5047, P2_REG3_REG_7__SCAN_IN, P2_U3088);
  nand ginst17267 (P2_U5048, P2_U3042, P2_U3449);
  nand ginst17268 (P2_U5049, P2_R1209_U16, P2_U3040);
  nand ginst17269 (P2_U5050, P2_ADDR_REG_7__SCAN_IN, P2_U4863);
  nand ginst17270 (P2_U5051, P2_R1170_U72, P2_U3043);
  nand ginst17271 (P2_U5052, P2_U3041, P2_U3446);
  nand ginst17272 (P2_U5053, P2_R1209_U72, P2_U3039);
  nand ginst17273 (P2_U5054, P2_U5051, P2_U5052, P2_U5053);
  nand ginst17274 (P2_U5055, P2_R1170_U72, P2_U3018);
  nand ginst17275 (P2_U5056, P2_R1209_U72, P2_U3017);
  nand ginst17276 (P2_U5057, P2_U3446, P2_U5683);
  nand ginst17277 (P2_U5058, P2_U5055, P2_U5056, P2_U5057);
  nand ginst17278 (P2_U5059, P2_U3045, P2_U5054);
  nand ginst17279 (P2_U5060, P2_U3947, P2_U5058);
  nand ginst17280 (P2_U5061, P2_R1170_U72, P2_U3044);
  nand ginst17281 (P2_U5062, P2_REG3_REG_6__SCAN_IN, P2_U3088);
  nand ginst17282 (P2_U5063, P2_U3042, P2_U3446);
  nand ginst17283 (P2_U5064, P2_R1209_U72, P2_U3040);
  nand ginst17284 (P2_U5065, P2_ADDR_REG_6__SCAN_IN, P2_U4863);
  nand ginst17285 (P2_U5066, P2_R1170_U15, P2_U3043);
  nand ginst17286 (P2_U5067, P2_U3041, P2_U3443);
  nand ginst17287 (P2_U5068, P2_R1209_U15, P2_U3039);
  nand ginst17288 (P2_U5069, P2_U5066, P2_U5067, P2_U5068);
  nand ginst17289 (P2_U5070, P2_R1170_U15, P2_U3018);
  nand ginst17290 (P2_U5071, P2_R1209_U15, P2_U3017);
  nand ginst17291 (P2_U5072, P2_U3443, P2_U5683);
  nand ginst17292 (P2_U5073, P2_U5070, P2_U5071, P2_U5072);
  nand ginst17293 (P2_U5074, P2_U3045, P2_U5069);
  nand ginst17294 (P2_U5075, P2_U3947, P2_U5073);
  nand ginst17295 (P2_U5076, P2_R1170_U15, P2_U3044);
  nand ginst17296 (P2_U5077, P2_REG3_REG_5__SCAN_IN, P2_U3088);
  nand ginst17297 (P2_U5078, P2_U3042, P2_U3443);
  nand ginst17298 (P2_U5079, P2_R1209_U15, P2_U3040);
  nand ginst17299 (P2_U5080, P2_ADDR_REG_5__SCAN_IN, P2_U4863);
  nand ginst17300 (P2_U5081, P2_R1170_U73, P2_U3043);
  nand ginst17301 (P2_U5082, P2_U3041, P2_U3440);
  nand ginst17302 (P2_U5083, P2_R1209_U73, P2_U3039);
  nand ginst17303 (P2_U5084, P2_U5081, P2_U5082, P2_U5083);
  nand ginst17304 (P2_U5085, P2_R1170_U73, P2_U3018);
  nand ginst17305 (P2_U5086, P2_R1209_U73, P2_U3017);
  nand ginst17306 (P2_U5087, P2_U3440, P2_U5683);
  nand ginst17307 (P2_U5088, P2_U5085, P2_U5086, P2_U5087);
  nand ginst17308 (P2_U5089, P2_U3045, P2_U5084);
  nand ginst17309 (P2_U5090, P2_U3947, P2_U5088);
  nand ginst17310 (P2_U5091, P2_R1170_U73, P2_U3044);
  nand ginst17311 (P2_U5092, P2_REG3_REG_4__SCAN_IN, P2_U3088);
  nand ginst17312 (P2_U5093, P2_U3042, P2_U3440);
  nand ginst17313 (P2_U5094, P2_R1209_U73, P2_U3040);
  nand ginst17314 (P2_U5095, P2_ADDR_REG_4__SCAN_IN, P2_U4863);
  nand ginst17315 (P2_U5096, P2_R1170_U74, P2_U3043);
  nand ginst17316 (P2_U5097, P2_U3041, P2_U3437);
  nand ginst17317 (P2_U5098, P2_R1209_U74, P2_U3039);
  nand ginst17318 (P2_U5099, P2_U5096, P2_U5097, P2_U5098);
  nand ginst17319 (P2_U5100, P2_R1170_U74, P2_U3018);
  nand ginst17320 (P2_U5101, P2_R1209_U74, P2_U3017);
  nand ginst17321 (P2_U5102, P2_U3437, P2_U5683);
  nand ginst17322 (P2_U5103, P2_U5100, P2_U5101, P2_U5102);
  nand ginst17323 (P2_U5104, P2_U3045, P2_U5099);
  nand ginst17324 (P2_U5105, P2_U3947, P2_U5103);
  nand ginst17325 (P2_U5106, P2_R1170_U74, P2_U3044);
  nand ginst17326 (P2_U5107, P2_REG3_REG_3__SCAN_IN, P2_U3088);
  nand ginst17327 (P2_U5108, P2_U3042, P2_U3437);
  nand ginst17328 (P2_U5109, P2_R1209_U74, P2_U3040);
  nand ginst17329 (P2_U5110, P2_ADDR_REG_3__SCAN_IN, P2_U4863);
  nand ginst17330 (P2_U5111, P2_R1170_U14, P2_U3043);
  nand ginst17331 (P2_U5112, P2_U3041, P2_U3434);
  nand ginst17332 (P2_U5113, P2_R1209_U14, P2_U3039);
  nand ginst17333 (P2_U5114, P2_U5111, P2_U5112, P2_U5113);
  nand ginst17334 (P2_U5115, P2_R1170_U14, P2_U3018);
  nand ginst17335 (P2_U5116, P2_R1209_U14, P2_U3017);
  nand ginst17336 (P2_U5117, P2_U3434, P2_U5683);
  nand ginst17337 (P2_U5118, P2_U5115, P2_U5116, P2_U5117);
  nand ginst17338 (P2_U5119, P2_U3045, P2_U5114);
  nand ginst17339 (P2_U5120, P2_U3947, P2_U5118);
  nand ginst17340 (P2_U5121, P2_R1170_U14, P2_U3044);
  nand ginst17341 (P2_U5122, P2_REG3_REG_2__SCAN_IN, P2_U3088);
  nand ginst17342 (P2_U5123, P2_U3042, P2_U3434);
  nand ginst17343 (P2_U5124, P2_R1209_U14, P2_U3040);
  nand ginst17344 (P2_U5125, P2_ADDR_REG_2__SCAN_IN, P2_U4863);
  nand ginst17345 (P2_U5126, P2_R1170_U68, P2_U3043);
  nand ginst17346 (P2_U5127, P2_U3041, P2_U3431);
  nand ginst17347 (P2_U5128, P2_R1209_U68, P2_U3039);
  nand ginst17348 (P2_U5129, P2_U5126, P2_U5127, P2_U5128);
  nand ginst17349 (P2_U5130, P2_R1170_U68, P2_U3018);
  nand ginst17350 (P2_U5131, P2_R1209_U68, P2_U3017);
  nand ginst17351 (P2_U5132, P2_U3431, P2_U5683);
  nand ginst17352 (P2_U5133, P2_U5130, P2_U5131, P2_U5132);
  nand ginst17353 (P2_U5134, P2_U3045, P2_U5129);
  nand ginst17354 (P2_U5135, P2_U3947, P2_U5133);
  nand ginst17355 (P2_U5136, P2_R1170_U68, P2_U3044);
  nand ginst17356 (P2_U5137, P2_REG3_REG_1__SCAN_IN, P2_U3088);
  nand ginst17357 (P2_U5138, P2_U3042, P2_U3431);
  nand ginst17358 (P2_U5139, P2_R1209_U68, P2_U3040);
  nand ginst17359 (P2_U5140, P2_ADDR_REG_1__SCAN_IN, P2_U4863);
  nand ginst17360 (P2_U5141, P2_R1170_U69, P2_U3043);
  nand ginst17361 (P2_U5142, P2_U3041, P2_U3425);
  nand ginst17362 (P2_U5143, P2_R1209_U69, P2_U3039);
  nand ginst17363 (P2_U5144, P2_U5141, P2_U5142, P2_U5143);
  nand ginst17364 (P2_U5145, P2_R1170_U69, P2_U3018);
  nand ginst17365 (P2_U5146, P2_R1209_U69, P2_U3017);
  nand ginst17366 (P2_U5147, P2_U3425, P2_U5683);
  nand ginst17367 (P2_U5148, P2_U5145, P2_U5146, P2_U5147);
  nand ginst17368 (P2_U5149, P2_U3045, P2_U5144);
  nand ginst17369 (P2_U5150, P2_U3947, P2_U5148);
  nand ginst17370 (P2_U5151, P2_R1170_U69, P2_U3044);
  nand ginst17371 (P2_U5152, P2_REG3_REG_0__SCAN_IN, P2_U3088);
  nand ginst17372 (P2_U5153, P2_U3042, P2_U3425);
  nand ginst17373 (P2_U5154, P2_R1209_U69, P2_U3040);
  nand ginst17374 (P2_U5155, P2_ADDR_REG_0__SCAN_IN, P2_U4863);
  not ginst17375 (P2_U5156, P2_U3918);
  nand ginst17376 (P2_U5157, P2_U3334, P2_U3337, P2_U3936);
  nand ginst17377 (P2_U5158, P2_U5665, P2_U5671);
  nand ginst17378 (P2_U5159, P2_U3424, P2_U5158);
  nand ginst17379 (P2_U5160, P2_U3419, P2_U5159);
  nand ginst17380 (P2_U5161, P2_U3340, P2_U5160);
  nand ginst17381 (P2_U5162, P2_U3052, P2_U6051, P2_U6052);
  nand ginst17382 (P2_U5163, P2_B_REG_SCAN_IN, P2_U5162);
  nand ginst17383 (P2_U5164, P2_U3038, P2_U3081);
  nand ginst17384 (P2_U5165, P2_U3036, P2_U3075);
  nand ginst17385 (P2_U5166, P2_ADD_1119_U69, P2_U3406);
  nand ginst17386 (P2_U5167, P2_U5164, P2_U5165, P2_U5166);
  not ginst17387 (P2_U5168, P2_U3154);
  nand ginst17388 (P2_U5169, P2_U3346, P2_U3923);
  nand ginst17389 (P2_U5170, P2_U3419, P2_U5169);
  nand ginst17390 (P2_U5171, P2_U3800, P2_U3801, P2_U5170);
  nand ginst17391 (P2_U5172, P2_U3406, P2_U5171);
  not ginst17392 (P2_U5173, P2_U3408);
  nand ginst17393 (P2_U5174, P2_U3474, P2_U5636);
  nand ginst17394 (P2_U5175, P2_ADD_1119_U69, P2_U5635);
  nand ginst17395 (P2_U5176, P2_R1176_U111, P2_U3028);
  nand ginst17396 (P2_U5177, P2_U3969, P2_U5167);
  nand ginst17397 (P2_U5178, P2_REG3_REG_15__SCAN_IN, P2_U3088);
  nand ginst17398 (P2_U5179, P2_U3038, P2_U3060);
  nand ginst17399 (P2_U5180, P2_U3036, P2_U3055);
  nand ginst17400 (P2_U5181, P2_ADD_1119_U58, P2_U3406);
  nand ginst17401 (P2_U5182, P2_U5179, P2_U5180, P2_U5181);
  nand ginst17402 (P2_U5183, P2_U3398, P2_U3406);
  nand ginst17403 (P2_U5184, P2_U5173, P2_U5183);
  nand ginst17404 (P2_U5185, P2_U3398, P2_U3946);
  nand ginst17405 (P2_U5186, P2_U3393, P2_U5185);
  nand ginst17406 (P2_U5187, P2_U3047, P2_U3951);
  nand ginst17407 (P2_U5188, P2_ADD_1119_U58, P2_U3046);
  nand ginst17408 (P2_U5189, P2_R1176_U16, P2_U3028);
  nand ginst17409 (P2_U5190, P2_U3969, P2_U5182);
  nand ginst17410 (P2_U5191, P2_REG3_REG_26__SCAN_IN, P2_U3088);
  nand ginst17411 (P2_U5192, P2_U3038, P2_U3069);
  nand ginst17412 (P2_U5193, P2_U3036, P2_U3072);
  nand ginst17413 (P2_U5194, P2_ADD_1119_U53, P2_U3406);
  nand ginst17414 (P2_U5195, P2_U5192, P2_U5193, P2_U5194);
  nand ginst17415 (P2_U5196, P2_U3447, P2_U5636);
  nand ginst17416 (P2_U5197, P2_ADD_1119_U53, P2_U5635);
  nand ginst17417 (P2_U5198, P2_R1176_U96, P2_U3028);
  nand ginst17418 (P2_U5199, P2_U3969, P2_U5195);
  nand ginst17419 (P2_U5200, P2_REG3_REG_6__SCAN_IN, P2_U3088);
  nand ginst17420 (P2_U5201, P2_U3038, P2_U3071);
  nand ginst17421 (P2_U5202, P2_U3036, P2_U3083);
  nand ginst17422 (P2_U5203, P2_ADD_1119_U66, P2_U3406);
  nand ginst17423 (P2_U5204, P2_U5201, P2_U5202, P2_U5203);
  nand ginst17424 (P2_U5205, P2_U3483, P2_U5636);
  nand ginst17425 (P2_U5206, P2_ADD_1119_U66, P2_U5635);
  nand ginst17426 (P2_U5207, P2_R1176_U109, P2_U3028);
  nand ginst17427 (P2_U5208, P2_U3969, P2_U5204);
  nand ginst17428 (P2_U5209, P2_REG3_REG_18__SCAN_IN, P2_U3088);
  nand ginst17429 (P2_U5210, P2_U3038, P2_U3080);
  nand ginst17430 (P2_U5211, P2_U3036, P2_U3066);
  nand ginst17431 (P2_U5212, P2_REG3_REG_2__SCAN_IN, P2_U3406);
  nand ginst17432 (P2_U5213, P2_U5210, P2_U5211, P2_U5212);
  nand ginst17433 (P2_U5214, P2_U3435, P2_U5636);
  nand ginst17434 (P2_U5215, P2_REG3_REG_2__SCAN_IN, P2_U5635);
  nand ginst17435 (P2_U5216, P2_R1176_U99, P2_U3028);
  nand ginst17436 (P2_U5217, P2_U3969, P2_U5213);
  nand ginst17437 (P2_U5218, P2_REG3_REG_2__SCAN_IN, P2_U3088);
  nand ginst17438 (P2_U5219, P2_U3038, P2_U3064);
  nand ginst17439 (P2_U5220, P2_U3036, P2_U3074);
  nand ginst17440 (P2_U5221, P2_ADD_1119_U73, P2_U3406);
  nand ginst17441 (P2_U5222, P2_U5219, P2_U5220, P2_U5221);
  nand ginst17442 (P2_U5223, P2_U3462, P2_U5636);
  nand ginst17443 (P2_U5224, P2_ADD_1119_U73, P2_U5635);
  nand ginst17444 (P2_U5225, P2_R1176_U114, P2_U3028);
  nand ginst17445 (P2_U5226, P2_U3969, P2_U5222);
  nand ginst17446 (P2_U5227, P2_REG3_REG_11__SCAN_IN, P2_U3088);
  nand ginst17447 (P2_U5228, P2_U3038, P2_U3077);
  nand ginst17448 (P2_U5229, P2_U3036, P2_U3068);
  nand ginst17449 (P2_U5230, P2_ADD_1119_U62, P2_U3406);
  nand ginst17450 (P2_U5231, P2_U5228, P2_U5229, P2_U5230);
  nand ginst17451 (P2_U5232, P2_U3047, P2_U3955);
  nand ginst17452 (P2_U5233, P2_ADD_1119_U62, P2_U3046);
  nand ginst17453 (P2_U5234, P2_R1176_U105, P2_U3028);
  nand ginst17454 (P2_U5235, P2_U3969, P2_U5231);
  nand ginst17455 (P2_U5236, P2_REG3_REG_22__SCAN_IN, P2_U3088);
  nand ginst17456 (P2_U5237, P2_U3038, P2_U3074);
  nand ginst17457 (P2_U5238, P2_U3036, P2_U3081);
  nand ginst17458 (P2_U5239, P2_ADD_1119_U71, P2_U3406);
  nand ginst17459 (P2_U5240, P2_U5237, P2_U5238, P2_U5239);
  nand ginst17460 (P2_U5241, P2_U3468, P2_U5636);
  nand ginst17461 (P2_U5242, P2_ADD_1119_U71, P2_U5635);
  nand ginst17462 (P2_U5243, P2_R1176_U13, P2_U3028);
  nand ginst17463 (P2_U5244, P2_U3969, P2_U5240);
  nand ginst17464 (P2_U5245, P2_REG3_REG_13__SCAN_IN, P2_U3088);
  nand ginst17465 (P2_U5246, P2_U3038, P2_U3083);
  nand ginst17466 (P2_U5247, P2_U3036, P2_U3077);
  nand ginst17467 (P2_U5248, P2_ADD_1119_U64, P2_U3406);
  nand ginst17468 (P2_U5249, P2_U5246, P2_U5247, P2_U5248);
  nand ginst17469 (P2_U5250, P2_U3047, P2_U3957);
  nand ginst17470 (P2_U5251, P2_ADD_1119_U64, P2_U3046);
  nand ginst17471 (P2_U5252, P2_R1176_U106, P2_U3028);
  nand ginst17472 (P2_U5253, P2_U3969, P2_U5249);
  nand ginst17473 (P2_U5254, P2_REG3_REG_20__SCAN_IN, P2_U3088);
  nand ginst17474 (P2_U5255, P2_U3405, P2_U3407);
  nand ginst17475 (P2_U5256, P2_U3406, P2_U5255);
  nand ginst17476 (P2_U5257, P2_U3970, P2_U5256);
  nand ginst17477 (P2_U5258, P2_U3036, P2_U3806);
  nand ginst17478 (P2_U5259, P2_U3427, P2_U5636);
  nand ginst17479 (P2_U5260, P2_REG3_REG_0__SCAN_IN, P2_U5257);
  nand ginst17480 (P2_U5261, P2_R1176_U93, P2_U3028);
  nand ginst17481 (P2_U5262, P2_REG3_REG_0__SCAN_IN, P2_U3088);
  nand ginst17482 (P2_U5263, P2_U3038, P2_U3086);
  nand ginst17483 (P2_U5264, P2_U3036, P2_U3064);
  nand ginst17484 (P2_U5265, P2_ADD_1119_U50, P2_U3406);
  nand ginst17485 (P2_U5266, P2_U5263, P2_U5264, P2_U5265);
  nand ginst17486 (P2_U5267, P2_U3456, P2_U5636);
  nand ginst17487 (P2_U5268, P2_ADD_1119_U50, P2_U5635);
  nand ginst17488 (P2_U5269, P2_R1176_U94, P2_U3028);
  nand ginst17489 (P2_U5270, P2_U3969, P2_U5266);
  nand ginst17490 (P2_U5271, P2_REG3_REG_9__SCAN_IN, P2_U3088);
  nand ginst17491 (P2_U5272, P2_U3038, P2_U3066);
  nand ginst17492 (P2_U5273, P2_U3036, P2_U3069);
  nand ginst17493 (P2_U5274, P2_ADD_1119_U55, P2_U3406);
  nand ginst17494 (P2_U5275, P2_U5272, P2_U5273, P2_U5274);
  nand ginst17495 (P2_U5276, P2_U3441, P2_U5636);
  nand ginst17496 (P2_U5277, P2_ADD_1119_U55, P2_U5635);
  nand ginst17497 (P2_U5278, P2_R1176_U98, P2_U3028);
  nand ginst17498 (P2_U5279, P2_U3969, P2_U5275);
  nand ginst17499 (P2_U5280, P2_REG3_REG_4__SCAN_IN, P2_U3088);
  nand ginst17500 (P2_U5281, P2_U3038, P2_U3068);
  nand ginst17501 (P2_U5282, P2_U3036, P2_U3060);
  nand ginst17502 (P2_U5283, P2_ADD_1119_U60, P2_U3406);
  nand ginst17503 (P2_U5284, P2_U5281, P2_U5282, P2_U5283);
  nand ginst17504 (P2_U5285, P2_U3047, P2_U3953);
  nand ginst17505 (P2_U5286, P2_ADD_1119_U60, P2_U3046);
  nand ginst17506 (P2_U5287, P2_R1176_U103, P2_U3028);
  nand ginst17507 (P2_U5288, P2_U3969, P2_U5284);
  nand ginst17508 (P2_U5289, P2_REG3_REG_24__SCAN_IN, P2_U3088);
  nand ginst17509 (P2_U5290, P2_U3038, P2_U3075);
  nand ginst17510 (P2_U5291, P2_U3036, P2_U3084);
  nand ginst17511 (P2_U5292, P2_ADD_1119_U67, P2_U3406);
  nand ginst17512 (P2_U5293, P2_U5290, P2_U5291, P2_U5292);
  nand ginst17513 (P2_U5294, P2_U3480, P2_U5636);
  nand ginst17514 (P2_U5295, P2_ADD_1119_U67, P2_U5635);
  nand ginst17515 (P2_U5296, P2_R1176_U14, P2_U3028);
  nand ginst17516 (P2_U5297, P2_U3969, P2_U5293);
  nand ginst17517 (P2_U5298, P2_REG3_REG_17__SCAN_IN, P2_U3088);
  nand ginst17518 (P2_U5299, P2_U3038, P2_U3062);
  nand ginst17519 (P2_U5300, P2_U3036, P2_U3073);
  nand ginst17520 (P2_U5301, P2_ADD_1119_U54, P2_U3406);
  nand ginst17521 (P2_U5302, P2_U5299, P2_U5300, P2_U5301);
  nand ginst17522 (P2_U5303, P2_U3444, P2_U5636);
  nand ginst17523 (P2_U5304, P2_ADD_1119_U54, P2_U5635);
  nand ginst17524 (P2_U5305, P2_R1176_U97, P2_U3028);
  nand ginst17525 (P2_U5306, P2_U3969, P2_U5302);
  nand ginst17526 (P2_U5307, P2_REG3_REG_5__SCAN_IN, P2_U3088);
  nand ginst17527 (P2_U5308, P2_U3038, P2_U3076);
  nand ginst17528 (P2_U5309, P2_U3036, P2_U3071);
  nand ginst17529 (P2_U5310, P2_ADD_1119_U68, P2_U3406);
  nand ginst17530 (P2_U5311, P2_U5308, P2_U5309, P2_U5310);
  nand ginst17531 (P2_U5312, P2_U3477, P2_U5636);
  nand ginst17532 (P2_U5313, P2_ADD_1119_U68, P2_U5635);
  nand ginst17533 (P2_U5314, P2_R1176_U110, P2_U3028);
  nand ginst17534 (P2_U5315, P2_U3969, P2_U5311);
  nand ginst17535 (P2_U5316, P2_REG3_REG_16__SCAN_IN, P2_U3088);
  nand ginst17536 (P2_U5317, P2_U3038, P2_U3067);
  nand ginst17537 (P2_U5318, P2_U3036, P2_U3059);
  nand ginst17538 (P2_U5319, P2_ADD_1119_U59, P2_U3406);
  nand ginst17539 (P2_U5320, P2_U5317, P2_U5318, P2_U5319);
  nand ginst17540 (P2_U5321, P2_U3047, P2_U3952);
  nand ginst17541 (P2_U5322, P2_ADD_1119_U59, P2_U3046);
  nand ginst17542 (P2_U5323, P2_R1176_U102, P2_U3028);
  nand ginst17543 (P2_U5324, P2_U3969, P2_U5320);
  nand ginst17544 (P2_U5325, P2_REG3_REG_25__SCAN_IN, P2_U3088);
  nand ginst17545 (P2_U5326, P2_U3038, P2_U3065);
  nand ginst17546 (P2_U5327, P2_U3036, P2_U3082);
  nand ginst17547 (P2_U5328, P2_ADD_1119_U72, P2_U3406);
  nand ginst17548 (P2_U5329, P2_U5326, P2_U5327, P2_U5328);
  nand ginst17549 (P2_U5330, P2_U3465, P2_U5636);
  nand ginst17550 (P2_U5331, P2_ADD_1119_U72, P2_U5635);
  nand ginst17551 (P2_U5332, P2_R1176_U113, P2_U3028);
  nand ginst17552 (P2_U5333, P2_U3969, P2_U5329);
  nand ginst17553 (P2_U5334, P2_REG3_REG_12__SCAN_IN, P2_U3088);
  nand ginst17554 (P2_U5335, P2_U3038, P2_U3078);
  nand ginst17555 (P2_U5336, P2_U3036, P2_U3063);
  nand ginst17556 (P2_U5337, P2_ADD_1119_U63, P2_U3406);
  nand ginst17557 (P2_U5338, P2_U5335, P2_U5336, P2_U5337);
  nand ginst17558 (P2_U5339, P2_U3047, P2_U3956);
  nand ginst17559 (P2_U5340, P2_ADD_1119_U63, P2_U3046);
  nand ginst17560 (P2_U5341, P2_R1176_U15, P2_U3028);
  nand ginst17561 (P2_U5342, P2_U3969, P2_U5338);
  nand ginst17562 (P2_U5343, P2_REG3_REG_21__SCAN_IN, P2_U3088);
  nand ginst17563 (P2_U5344, P2_U3038, P2_U3079);
  nand ginst17564 (P2_U5345, P2_U3036, P2_U3070);
  nand ginst17565 (P2_U5346, P2_REG3_REG_1__SCAN_IN, P2_U3406);
  nand ginst17566 (P2_U5347, P2_U5344, P2_U5345, P2_U5346);
  nand ginst17567 (P2_U5348, P2_U3432, P2_U5636);
  nand ginst17568 (P2_U5349, P2_REG3_REG_1__SCAN_IN, P2_U5635);
  nand ginst17569 (P2_U5350, P2_R1176_U107, P2_U3028);
  nand ginst17570 (P2_U5351, P2_U3969, P2_U5347);
  nand ginst17571 (P2_U5352, P2_REG3_REG_1__SCAN_IN, P2_U3088);
  nand ginst17572 (P2_U5353, P2_U3038, P2_U3072);
  nand ginst17573 (P2_U5354, P2_U3036, P2_U3085);
  nand ginst17574 (P2_U5355, P2_ADD_1119_U51, P2_U3406);
  nand ginst17575 (P2_U5356, P2_U5353, P2_U5354, P2_U5355);
  nand ginst17576 (P2_U5357, P2_U3453, P2_U5636);
  nand ginst17577 (P2_U5358, P2_ADD_1119_U51, P2_U5635);
  nand ginst17578 (P2_U5359, P2_R1176_U95, P2_U3028);
  nand ginst17579 (P2_U5360, P2_U3969, P2_U5356);
  nand ginst17580 (P2_U5361, P2_REG3_REG_8__SCAN_IN, P2_U3088);
  nand ginst17581 (P2_U5362, P2_U3038, P2_U3055);
  nand ginst17582 (P2_U5363, P2_U3036, P2_U3057);
  nand ginst17583 (P2_U5364, P2_ADD_1119_U56, P2_U3406);
  nand ginst17584 (P2_U5365, P2_U5362, P2_U5363, P2_U5364);
  nand ginst17585 (P2_U5366, P2_U3047, P2_U3949);
  nand ginst17586 (P2_U5367, P2_ADD_1119_U56, P2_U3046);
  nand ginst17587 (P2_U5368, P2_R1176_U100, P2_U3028);
  nand ginst17588 (P2_U5369, P2_U3969, P2_U5365);
  nand ginst17589 (P2_U5370, P2_REG3_REG_28__SCAN_IN, P2_U3088);
  nand ginst17590 (P2_U5371, P2_U3038, P2_U3084);
  nand ginst17591 (P2_U5372, P2_U3036, P2_U3078);
  nand ginst17592 (P2_U5373, P2_ADD_1119_U65, P2_U3406);
  nand ginst17593 (P2_U5374, P2_U5371, P2_U5372, P2_U5373);
  nand ginst17594 (P2_U5375, P2_U3485, P2_U5636);
  nand ginst17595 (P2_U5376, P2_ADD_1119_U65, P2_U5635);
  nand ginst17596 (P2_U5377, P2_R1176_U108, P2_U3028);
  nand ginst17597 (P2_U5378, P2_U3969, P2_U5374);
  nand ginst17598 (P2_U5379, P2_REG3_REG_19__SCAN_IN, P2_U3088);
  nand ginst17599 (P2_U5380, P2_U3038, P2_U3070);
  nand ginst17600 (P2_U5381, P2_U3036, P2_U3062);
  nand ginst17601 (P2_U5382, P2_ADD_1119_U4, P2_U3406);
  nand ginst17602 (P2_U5383, P2_U5380, P2_U5381, P2_U5382);
  nand ginst17603 (P2_U5384, P2_U3438, P2_U5636);
  nand ginst17604 (P2_U5385, P2_ADD_1119_U4, P2_U5635);
  nand ginst17605 (P2_U5386, P2_R1176_U17, P2_U3028);
  nand ginst17606 (P2_U5387, P2_U3969, P2_U5383);
  nand ginst17607 (P2_U5388, P2_REG3_REG_3__SCAN_IN, P2_U3088);
  nand ginst17608 (P2_U5389, P2_U3038, P2_U3085);
  nand ginst17609 (P2_U5390, P2_U3036, P2_U3065);
  nand ginst17610 (P2_U5391, P2_ADD_1119_U74, P2_U3406);
  nand ginst17611 (P2_U5392, P2_U5389, P2_U5390, P2_U5391);
  nand ginst17612 (P2_U5393, P2_U3459, P2_U5636);
  nand ginst17613 (P2_U5394, P2_ADD_1119_U74, P2_U5635);
  nand ginst17614 (P2_U5395, P2_R1176_U115, P2_U3028);
  nand ginst17615 (P2_U5396, P2_U3969, P2_U5392);
  nand ginst17616 (P2_U5397, P2_REG3_REG_10__SCAN_IN, P2_U3088);
  nand ginst17617 (P2_U5398, P2_U3038, P2_U3063);
  nand ginst17618 (P2_U5399, P2_U3036, P2_U3067);
  nand ginst17619 (P2_U5400, P2_ADD_1119_U61, P2_U3406);
  nand ginst17620 (P2_U5401, P2_U5398, P2_U5399, P2_U5400);
  nand ginst17621 (P2_U5402, P2_U3047, P2_U3954);
  nand ginst17622 (P2_U5403, P2_ADD_1119_U61, P2_U3046);
  nand ginst17623 (P2_U5404, P2_R1176_U104, P2_U3028);
  nand ginst17624 (P2_U5405, P2_U3969, P2_U5401);
  nand ginst17625 (P2_U5406, P2_REG3_REG_23__SCAN_IN, P2_U3088);
  nand ginst17626 (P2_U5407, P2_U3038, P2_U3082);
  nand ginst17627 (P2_U5408, P2_U3036, P2_U3076);
  nand ginst17628 (P2_U5409, P2_ADD_1119_U70, P2_U3406);
  nand ginst17629 (P2_U5410, P2_U5407, P2_U5408, P2_U5409);
  nand ginst17630 (P2_U5411, P2_U3471, P2_U5636);
  nand ginst17631 (P2_U5412, P2_ADD_1119_U70, P2_U5635);
  nand ginst17632 (P2_U5413, P2_R1176_U112, P2_U3028);
  nand ginst17633 (P2_U5414, P2_U3969, P2_U5410);
  nand ginst17634 (P2_U5415, P2_REG3_REG_14__SCAN_IN, P2_U3088);
  nand ginst17635 (P2_U5416, P2_U3038, P2_U3059);
  nand ginst17636 (P2_U5417, P2_U3036, P2_U3056);
  nand ginst17637 (P2_U5418, P2_ADD_1119_U57, P2_U3406);
  nand ginst17638 (P2_U5419, P2_U5416, P2_U5417, P2_U5418);
  nand ginst17639 (P2_U5420, P2_U3047, P2_U3950);
  nand ginst17640 (P2_U5421, P2_ADD_1119_U57, P2_U3046);
  nand ginst17641 (P2_U5422, P2_R1176_U101, P2_U3028);
  nand ginst17642 (P2_U5423, P2_U3969, P2_U5419);
  nand ginst17643 (P2_U5424, P2_REG3_REG_27__SCAN_IN, P2_U3088);
  nand ginst17644 (P2_U5425, P2_U3038, P2_U3073);
  nand ginst17645 (P2_U5426, P2_U3036, P2_U3086);
  nand ginst17646 (P2_U5427, P2_ADD_1119_U52, P2_U3406);
  nand ginst17647 (P2_U5428, P2_U5425, P2_U5426, P2_U5427);
  nand ginst17648 (P2_U5429, P2_U3450, P2_U5636);
  nand ginst17649 (P2_U5430, P2_ADD_1119_U52, P2_U5635);
  nand ginst17650 (P2_U5431, P2_R1176_U18, P2_U3028);
  nand ginst17651 (P2_U5432, P2_U3969, P2_U5428);
  nand ginst17652 (P2_U5433, P2_REG3_REG_7__SCAN_IN, P2_U3088);
  nand ginst17653 (P2_U5434, P2_U3048, P2_U3948);
  nand ginst17654 (P2_U5435, P2_U3347, P2_U3415);
  nand ginst17655 (P2_U5436, P2_U3418, P2_U3419);
  nand ginst17656 (P2_U5437, P2_U3051, P2_U3816);
  not ginst17657 (P2_U5438, P2_U3411);
  nand ginst17658 (P2_U5439, P2_U3015, P2_U3415);
  nand ginst17659 (P2_U5440, P2_U3409, P2_U3411);
  nand ginst17660 (P2_U5441, P2_U3053, P2_U5440);
  nand ginst17661 (P2_U5442, P2_U3029, P2_U3085);
  nand ginst17662 (P2_U5443, P2_U3085, P2_U5441);
  nand ginst17663 (P2_U5444, P2_U3456, P2_U3929);
  nand ginst17664 (P2_U5445, P2_U3029, P2_U3086);
  nand ginst17665 (P2_U5446, P2_U3086, P2_U5441);
  nand ginst17666 (P2_U5447, P2_U3453, P2_U3929);
  nand ginst17667 (P2_U5448, P2_U3029, P2_U3072);
  nand ginst17668 (P2_U5449, P2_U3072, P2_U5441);
  nand ginst17669 (P2_U5450, P2_U3450, P2_U3929);
  nand ginst17670 (P2_U5451, P2_U3029, P2_U3073);
  nand ginst17671 (P2_U5452, P2_U3073, P2_U5441);
  nand ginst17672 (P2_U5453, P2_U3447, P2_U3929);
  nand ginst17673 (P2_U5454, P2_U3029, P2_U3069);
  nand ginst17674 (P2_U5455, P2_U3069, P2_U5441);
  nand ginst17675 (P2_U5456, P2_U3444, P2_U3929);
  nand ginst17676 (P2_U5457, P2_U3029, P2_U3062);
  nand ginst17677 (P2_U5458, P2_U3062, P2_U5441);
  nand ginst17678 (P2_U5459, P2_U3441, P2_U3929);
  nand ginst17679 (P2_U5460, P2_R1335_U8, P2_U3029);
  nand ginst17680 (P2_U5461, P2_U3058, P2_U5441);
  nand ginst17681 (P2_U5462, P2_R1335_U6, P2_U3029);
  nand ginst17682 (P2_U5463, P2_U3061, P2_U5441);
  nand ginst17683 (P2_U5464, P2_U3347, P2_U3929, U70);
  nand ginst17684 (P2_U5465, P2_U3029, P2_U3066);
  nand ginst17685 (P2_U5466, P2_U3066, P2_U5441);
  nand ginst17686 (P2_U5467, P2_U3438, P2_U3929);
  nand ginst17687 (P2_U5468, P2_U3029, P2_U3057);
  nand ginst17688 (P2_U5469, P2_U3057, P2_U5441);
  nand ginst17689 (P2_U5470, P2_U3929, P2_U3960);
  nand ginst17690 (P2_U5471, P2_U3029, P2_U3056);
  nand ginst17691 (P2_U5472, P2_U3056, P2_U5441);
  nand ginst17692 (P2_U5473, P2_U3929, P2_U3949);
  nand ginst17693 (P2_U5474, P2_U3029, P2_U3055);
  nand ginst17694 (P2_U5475, P2_U3055, P2_U5441);
  nand ginst17695 (P2_U5476, P2_U3929, P2_U3950);
  nand ginst17696 (P2_U5477, P2_U3029, P2_U3059);
  nand ginst17697 (P2_U5478, P2_U3059, P2_U5441);
  nand ginst17698 (P2_U5479, P2_U3929, P2_U3951);
  nand ginst17699 (P2_U5480, P2_U3029, P2_U3060);
  nand ginst17700 (P2_U5481, P2_U3060, P2_U5441);
  nand ginst17701 (P2_U5482, P2_U3929, P2_U3952);
  nand ginst17702 (P2_U5483, P2_U3029, P2_U3067);
  nand ginst17703 (P2_U5484, P2_U3067, P2_U5441);
  nand ginst17704 (P2_U5485, P2_U3929, P2_U3953);
  nand ginst17705 (P2_U5486, P2_U3029, P2_U3068);
  nand ginst17706 (P2_U5487, P2_U3068, P2_U5441);
  nand ginst17707 (P2_U5488, P2_U3929, P2_U3954);
  nand ginst17708 (P2_U5489, P2_U3029, P2_U3063);
  nand ginst17709 (P2_U5490, P2_U3063, P2_U5441);
  nand ginst17710 (P2_U5491, P2_U3929, P2_U3955);
  nand ginst17711 (P2_U5492, P2_U3029, P2_U3077);
  nand ginst17712 (P2_U5493, P2_U3077, P2_U5441);
  nand ginst17713 (P2_U5494, P2_U3929, P2_U3956);
  nand ginst17714 (P2_U5495, P2_U3029, P2_U3078);
  nand ginst17715 (P2_U5496, P2_U3078, P2_U5441);
  nand ginst17716 (P2_U5497, P2_U3929, P2_U3957);
  nand ginst17717 (P2_U5498, P2_U3029, P2_U3070);
  nand ginst17718 (P2_U5499, P2_U3070, P2_U5441);
  nand ginst17719 (P2_U5500, P2_U3435, P2_U3929);
  nand ginst17720 (P2_U5501, P2_U3029, P2_U3083);
  nand ginst17721 (P2_U5502, P2_U3083, P2_U5441);
  nand ginst17722 (P2_U5503, P2_U3485, P2_U3929);
  nand ginst17723 (P2_U5504, P2_U3029, P2_U3084);
  nand ginst17724 (P2_U5505, P2_U3084, P2_U5441);
  nand ginst17725 (P2_U5506, P2_U3483, P2_U3929);
  nand ginst17726 (P2_U5507, P2_U3029, P2_U3071);
  nand ginst17727 (P2_U5508, P2_U3071, P2_U5441);
  nand ginst17728 (P2_U5509, P2_U3480, P2_U3929);
  nand ginst17729 (P2_U5510, P2_U3029, P2_U3075);
  nand ginst17730 (P2_U5511, P2_U3075, P2_U5441);
  nand ginst17731 (P2_U5512, P2_U3477, P2_U3929);
  nand ginst17732 (P2_U5513, P2_U3029, P2_U3076);
  nand ginst17733 (P2_U5514, P2_U3076, P2_U5441);
  nand ginst17734 (P2_U5515, P2_U3474, P2_U3929);
  nand ginst17735 (P2_U5516, P2_U3029, P2_U3081);
  nand ginst17736 (P2_U5517, P2_U3081, P2_U5441);
  nand ginst17737 (P2_U5518, P2_U3471, P2_U3929);
  nand ginst17738 (P2_U5519, P2_U3029, P2_U3082);
  nand ginst17739 (P2_U5520, P2_U3082, P2_U5441);
  nand ginst17740 (P2_U5521, P2_U3468, P2_U3929);
  nand ginst17741 (P2_U5522, P2_U3029, P2_U3074);
  nand ginst17742 (P2_U5523, P2_U3074, P2_U5441);
  nand ginst17743 (P2_U5524, P2_U3465, P2_U3929);
  nand ginst17744 (P2_U5525, P2_U3029, P2_U3065);
  nand ginst17745 (P2_U5526, P2_U3065, P2_U5441);
  nand ginst17746 (P2_U5527, P2_U3462, P2_U3929);
  nand ginst17747 (P2_U5528, P2_U3029, P2_U3064);
  nand ginst17748 (P2_U5529, P2_U3064, P2_U5441);
  nand ginst17749 (P2_U5530, P2_U3459, P2_U3929);
  nand ginst17750 (P2_U5531, P2_U3029, P2_U3080);
  nand ginst17751 (P2_U5532, P2_U3080, P2_U5441);
  nand ginst17752 (P2_U5533, P2_U3432, P2_U3929);
  nand ginst17753 (P2_U5534, P2_U3029, P2_U3079);
  nand ginst17754 (P2_U5535, P2_U3079, P2_U5441);
  nand ginst17755 (P2_U5536, P2_U3427, P2_U3929);
  nand ginst17756 (P2_U5537, P2_U3053, P2_U5438);
  nand ginst17757 (P2_U5538, P2_U3456, P2_U5537);
  nand ginst17758 (P2_U5539, P2_U3085, P2_U3929);
  nand ginst17759 (P2_U5540, P2_U3086, P2_U5658);
  nand ginst17760 (P2_U5541, P2_U3453, P2_U5537);
  nand ginst17761 (P2_U5542, P2_U3086, P2_U3929);
  nand ginst17762 (P2_U5543, P2_U3072, P2_U5658);
  nand ginst17763 (P2_U5544, P2_U3450, P2_U5537);
  nand ginst17764 (P2_U5545, P2_U3072, P2_U3929);
  nand ginst17765 (P2_U5546, P2_U3073, P2_U5658);
  nand ginst17766 (P2_U5547, P2_U3447, P2_U5537);
  nand ginst17767 (P2_U5548, P2_U3073, P2_U3929);
  nand ginst17768 (P2_U5549, P2_U3069, P2_U5658);
  nand ginst17769 (P2_U5550, P2_U3444, P2_U5537);
  nand ginst17770 (P2_U5551, P2_U3069, P2_U3929);
  nand ginst17771 (P2_U5552, P2_U3062, P2_U5658);
  nand ginst17772 (P2_U5553, P2_U3441, P2_U5537);
  nand ginst17773 (P2_U5554, P2_U3062, P2_U3929);
  nand ginst17774 (P2_U5555, P2_U3066, P2_U5658);
  nand ginst17775 (P2_U5556, P2_U3347, P2_U5537, U69);
  nand ginst17776 (P2_U5557, P2_U3058, P2_U3929);
  nand ginst17777 (P2_U5558, P2_U3959, P2_U5537);
  nand ginst17778 (P2_U5559, P2_U3061, P2_U3929);
  nand ginst17779 (P2_U5560, P2_U3438, P2_U5537);
  nand ginst17780 (P2_U5561, P2_U3066, P2_U3929);
  nand ginst17781 (P2_U5562, P2_U3070, P2_U5658);
  nand ginst17782 (P2_U5563, P2_U3960, P2_U5537);
  nand ginst17783 (P2_U5564, P2_U3057, P2_U3929);
  nand ginst17784 (P2_U5565, P2_U3056, P2_U5658);
  nand ginst17785 (P2_U5566, P2_U3949, P2_U5537);
  nand ginst17786 (P2_U5567, P2_U3056, P2_U3929);
  nand ginst17787 (P2_U5568, P2_U3055, P2_U5658);
  nand ginst17788 (P2_U5569, P2_U3950, P2_U5537);
  nand ginst17789 (P2_U5570, P2_U3055, P2_U3929);
  nand ginst17790 (P2_U5571, P2_U3059, P2_U5658);
  nand ginst17791 (P2_U5572, P2_U3951, P2_U5537);
  nand ginst17792 (P2_U5573, P2_U3059, P2_U3929);
  nand ginst17793 (P2_U5574, P2_U3060, P2_U5658);
  nand ginst17794 (P2_U5575, P2_U3952, P2_U5537);
  nand ginst17795 (P2_U5576, P2_U3060, P2_U3929);
  nand ginst17796 (P2_U5577, P2_U3067, P2_U5658);
  nand ginst17797 (P2_U5578, P2_U3953, P2_U5537);
  nand ginst17798 (P2_U5579, P2_U3067, P2_U3929);
  nand ginst17799 (P2_U5580, P2_U3068, P2_U5658);
  nand ginst17800 (P2_U5581, P2_U3954, P2_U5537);
  nand ginst17801 (P2_U5582, P2_U3068, P2_U3929);
  nand ginst17802 (P2_U5583, P2_U3063, P2_U5658);
  nand ginst17803 (P2_U5584, P2_U3955, P2_U5537);
  nand ginst17804 (P2_U5585, P2_U3063, P2_U3929);
  nand ginst17805 (P2_U5586, P2_U3077, P2_U5658);
  nand ginst17806 (P2_U5587, P2_U3956, P2_U5537);
  nand ginst17807 (P2_U5588, P2_U3077, P2_U3929);
  nand ginst17808 (P2_U5589, P2_U3078, P2_U5658);
  nand ginst17809 (P2_U5590, P2_U3957, P2_U5537);
  nand ginst17810 (P2_U5591, P2_U3078, P2_U3929);
  nand ginst17811 (P2_U5592, P2_U3083, P2_U5658);
  nand ginst17812 (P2_U5593, P2_U3435, P2_U5537);
  nand ginst17813 (P2_U5594, P2_U3070, P2_U3929);
  nand ginst17814 (P2_U5595, P2_U3080, P2_U5658);
  nand ginst17815 (P2_U5596, P2_U3485, P2_U5537);
  nand ginst17816 (P2_U5597, P2_U3083, P2_U3929);
  nand ginst17817 (P2_U5598, P2_U3084, P2_U5658);
  nand ginst17818 (P2_U5599, P2_U3483, P2_U5537);
  nand ginst17819 (P2_U5600, P2_U3084, P2_U3929);
  nand ginst17820 (P2_U5601, P2_U3071, P2_U5658);
  nand ginst17821 (P2_U5602, P2_U3480, P2_U5537);
  nand ginst17822 (P2_U5603, P2_U3071, P2_U3929);
  nand ginst17823 (P2_U5604, P2_U3075, P2_U5658);
  nand ginst17824 (P2_U5605, P2_U3477, P2_U5537);
  nand ginst17825 (P2_U5606, P2_U3075, P2_U3929);
  nand ginst17826 (P2_U5607, P2_U3076, P2_U5658);
  nand ginst17827 (P2_U5608, P2_U3474, P2_U5537);
  nand ginst17828 (P2_U5609, P2_U3076, P2_U3929);
  nand ginst17829 (P2_U5610, P2_U3081, P2_U5658);
  nand ginst17830 (P2_U5611, P2_U3471, P2_U5537);
  nand ginst17831 (P2_U5612, P2_U3081, P2_U3929);
  nand ginst17832 (P2_U5613, P2_U3082, P2_U5658);
  nand ginst17833 (P2_U5614, P2_U3468, P2_U5537);
  nand ginst17834 (P2_U5615, P2_U3082, P2_U3929);
  nand ginst17835 (P2_U5616, P2_U3074, P2_U5658);
  nand ginst17836 (P2_U5617, P2_U3465, P2_U5537);
  nand ginst17837 (P2_U5618, P2_U3074, P2_U3929);
  nand ginst17838 (P2_U5619, P2_U3065, P2_U5658);
  nand ginst17839 (P2_U5620, P2_U3462, P2_U5537);
  nand ginst17840 (P2_U5621, P2_U3065, P2_U3929);
  nand ginst17841 (P2_U5622, P2_U3064, P2_U5658);
  nand ginst17842 (P2_U5623, P2_U3459, P2_U5537);
  nand ginst17843 (P2_U5624, P2_U3064, P2_U3929);
  nand ginst17844 (P2_U5625, P2_U3085, P2_U5658);
  nand ginst17845 (P2_U5626, P2_U3432, P2_U5537);
  nand ginst17846 (P2_U5627, P2_U3080, P2_U3929);
  nand ginst17847 (P2_U5628, P2_U3079, P2_U5658);
  nand ginst17848 (P2_U5629, P2_U3427, P2_U5537);
  nand ginst17849 (P2_U5630, P2_U3079, P2_U3929);
  nand ginst17850 (P2_U5631, P2_U3088, P2_U5163);
  nand ginst17851 (P2_U5632, P2_U3828, P2_U5461);
  nand ginst17852 (P2_U5633, P2_U3406, P2_U3972);
  nand ginst17853 (P2_U5634, P2_U3946, P2_U3972);
  nand ginst17854 (P2_U5635, P2_U3970, P2_U5633);
  nand ginst17855 (P2_U5636, P2_U3971, P2_U5634);
  nand ginst17856 (P2_U5637, P2_U3054, P2_U3945);
  nand ginst17857 (P2_U5638, P2_U3054, P2_U3330);
  nand ginst17858 (P2_U5639, P2_U3023, P2_U3961);
  nand ginst17859 (P2_U5640, P2_U3787, P2_U5163);
  nand ginst17860 (P2_U5641, P2_U3917, P2_U5163, P2_U6149, P2_U6150);
  nand ginst17861 (P2_U5642, P2_U5646, P2_U5652);
  nand ginst17862 (P2_U5643, P2_U3347, P2_U3415);
  nand ginst17863 (P2_U5644, P2_IR_REG_24__SCAN_IN, P2_U3879);
  nand ginst17864 (P2_U5645, P2_IR_REG_31__SCAN_IN, P2_SUB_1108_U14);
  not ginst17865 (P2_U5646, P2_U3412);
  nand ginst17866 (P2_U5647, P2_IR_REG_25__SCAN_IN, P2_U3879);
  nand ginst17867 (P2_U5648, P2_IR_REG_31__SCAN_IN, P2_SUB_1108_U112);
  not ginst17868 (P2_U5649, P2_U3413);
  nand ginst17869 (P2_U5650, P2_IR_REG_26__SCAN_IN, P2_U3879);
  nand ginst17870 (P2_U5651, P2_IR_REG_31__SCAN_IN, P2_SUB_1108_U15);
  not ginst17871 (P2_U5652, P2_U3414);
  nand ginst17872 (P2_U5653, P2_B_REG_SCAN_IN, P2_U5646);
  nand ginst17873 (P2_U5654, P2_U3331, P2_U3412);
  nand ginst17874 (P2_U5655, P2_U5653, P2_U5654);
  nand ginst17875 (P2_U5656, P2_IR_REG_23__SCAN_IN, P2_U3879);
  nand ginst17876 (P2_U5657, P2_IR_REG_31__SCAN_IN, P2_SUB_1108_U13);
  not ginst17877 (P2_U5658, P2_U3415);
  nand ginst17878 (P2_U5659, P2_D_REG_0__SCAN_IN, P2_U3880);
  nand ginst17879 (P2_U5660, P2_U3967, P2_U4077);
  nand ginst17880 (P2_U5661, P2_D_REG_1__SCAN_IN, P2_U3880);
  nand ginst17881 (P2_U5662, P2_U3967, P2_U4078);
  nand ginst17882 (P2_U5663, P2_IR_REG_22__SCAN_IN, P2_U3879);
  nand ginst17883 (P2_U5664, P2_IR_REG_31__SCAN_IN, P2_SUB_1108_U114);
  not ginst17884 (P2_U5665, P2_U3420);
  nand ginst17885 (P2_U5666, P2_IR_REG_19__SCAN_IN, P2_U3879);
  nand ginst17886 (P2_U5667, P2_IR_REG_31__SCAN_IN, P2_SUB_1108_U123);
  not ginst17887 (P2_U5668, P2_U3424);
  nand ginst17888 (P2_U5669, P2_IR_REG_20__SCAN_IN, P2_U3879);
  nand ginst17889 (P2_U5670, P2_IR_REG_31__SCAN_IN, P2_SUB_1108_U119);
  not ginst17890 (P2_U5671, P2_U3418);
  nand ginst17891 (P2_U5672, P2_IR_REG_21__SCAN_IN, P2_U3879);
  nand ginst17892 (P2_U5673, P2_IR_REG_31__SCAN_IN, P2_SUB_1108_U116);
  not ginst17893 (P2_U5674, P2_U3419);
  nand ginst17894 (P2_U5675, P2_IR_REG_30__SCAN_IN, P2_U3879);
  nand ginst17895 (P2_U5676, P2_IR_REG_31__SCAN_IN, P2_SUB_1108_U104);
  not ginst17896 (P2_U5677, P2_U3421);
  nand ginst17897 (P2_U5678, P2_IR_REG_29__SCAN_IN, P2_U3879);
  nand ginst17898 (P2_U5679, P2_IR_REG_31__SCAN_IN, P2_SUB_1108_U16);
  not ginst17899 (P2_U5680, P2_U3422);
  nand ginst17900 (P2_U5681, P2_IR_REG_28__SCAN_IN, P2_U3879);
  nand ginst17901 (P2_U5682, P2_IR_REG_31__SCAN_IN, P2_SUB_1108_U107);
  not ginst17902 (P2_U5683, P2_U3423);
  nand ginst17903 (P2_U5684, P2_IR_REG_0__SCAN_IN, P2_U3879);
  nand ginst17904 (P2_U5685, P2_IR_REG_0__SCAN_IN, P2_IR_REG_31__SCAN_IN);
  nand ginst17905 (P2_U5686, P2_IR_REG_27__SCAN_IN, P2_U3879);
  nand ginst17906 (P2_U5687, P2_IR_REG_31__SCAN_IN, P2_SUB_1108_U110);
  not ginst17907 (P2_U5688, P2_U3426);
  nand ginst17908 (P2_U5689, P2_U3347, U93);
  nand ginst17909 (P2_U5690, P2_U3425, P2_U3945);
  not ginst17910 (P2_U5691, P2_U3427);
  nand ginst17911 (P2_U5692, P2_U3420, P2_U5674);
  nand ginst17912 (P2_U5693, P2_U4109, P2_U5665);
  nand ginst17913 (P2_U5694, P2_D_REG_1__SCAN_IN, P2_U4076);
  nand ginst17914 (P2_U5695, P2_U3333, P2_U4078);
  not ginst17915 (P2_U5696, P2_U3429);
  nand ginst17916 (P2_U5697, P2_U3333, P2_U5642);
  nand ginst17917 (P2_U5698, P2_D_REG_0__SCAN_IN, P2_U4076);
  not ginst17918 (P2_U5699, P2_U3428);
  nand ginst17919 (P2_U5700, P2_REG0_REG_0__SCAN_IN, P2_U3881);
  nand ginst17920 (P2_U5701, P2_U3966, P2_U4129);
  nand ginst17921 (P2_U5702, P2_IR_REG_1__SCAN_IN, P2_U3879);
  nand ginst17922 (P2_U5703, P2_IR_REG_31__SCAN_IN, P2_SUB_1108_U42);
  nand ginst17923 (P2_U5704, P2_U3347, U82);
  nand ginst17924 (P2_U5705, P2_U3431, P2_U3945);
  not ginst17925 (P2_U5706, P2_U3432);
  nand ginst17926 (P2_U5707, P2_REG0_REG_1__SCAN_IN, P2_U3881);
  nand ginst17927 (P2_U5708, P2_U3966, P2_U4153);
  nand ginst17928 (P2_U5709, P2_IR_REG_2__SCAN_IN, P2_U3879);
  nand ginst17929 (P2_U5710, P2_IR_REG_31__SCAN_IN, P2_SUB_1108_U17);
  nand ginst17930 (P2_U5711, P2_U3347, U71);
  nand ginst17931 (P2_U5712, P2_U3434, P2_U3945);
  not ginst17932 (P2_U5713, P2_U3435);
  nand ginst17933 (P2_U5714, P2_REG0_REG_2__SCAN_IN, P2_U3881);
  nand ginst17934 (P2_U5715, P2_U3966, P2_U4172);
  nand ginst17935 (P2_U5716, P2_IR_REG_3__SCAN_IN, P2_U3879);
  nand ginst17936 (P2_U5717, P2_IR_REG_31__SCAN_IN, P2_SUB_1108_U18);
  nand ginst17937 (P2_U5718, P2_U3347, U68);
  nand ginst17938 (P2_U5719, P2_U3437, P2_U3945);
  not ginst17939 (P2_U5720, P2_U3438);
  nand ginst17940 (P2_U5721, P2_REG0_REG_3__SCAN_IN, P2_U3881);
  nand ginst17941 (P2_U5722, P2_U3966, P2_U4191);
  nand ginst17942 (P2_U5723, P2_IR_REG_4__SCAN_IN, P2_U3879);
  nand ginst17943 (P2_U5724, P2_IR_REG_31__SCAN_IN, P2_SUB_1108_U19);
  nand ginst17944 (P2_U5725, P2_U3347, U67);
  nand ginst17945 (P2_U5726, P2_U3440, P2_U3945);
  not ginst17946 (P2_U5727, P2_U3441);
  nand ginst17947 (P2_U5728, P2_REG0_REG_4__SCAN_IN, P2_U3881);
  nand ginst17948 (P2_U5729, P2_U3966, P2_U4210);
  nand ginst17949 (P2_U5730, P2_IR_REG_5__SCAN_IN, P2_U3879);
  nand ginst17950 (P2_U5731, P2_IR_REG_31__SCAN_IN, P2_SUB_1108_U101);
  nand ginst17951 (P2_U5732, P2_U3347, U66);
  nand ginst17952 (P2_U5733, P2_U3443, P2_U3945);
  not ginst17953 (P2_U5734, P2_U3444);
  nand ginst17954 (P2_U5735, P2_REG0_REG_5__SCAN_IN, P2_U3881);
  nand ginst17955 (P2_U5736, P2_U3966, P2_U4229);
  nand ginst17956 (P2_U5737, P2_IR_REG_6__SCAN_IN, P2_U3879);
  nand ginst17957 (P2_U5738, P2_IR_REG_31__SCAN_IN, P2_SUB_1108_U20);
  nand ginst17958 (P2_U5739, P2_U3347, U65);
  nand ginst17959 (P2_U5740, P2_U3446, P2_U3945);
  not ginst17960 (P2_U5741, P2_U3447);
  nand ginst17961 (P2_U5742, P2_REG0_REG_6__SCAN_IN, P2_U3881);
  nand ginst17962 (P2_U5743, P2_U3966, P2_U4248);
  nand ginst17963 (P2_U5744, P2_IR_REG_7__SCAN_IN, P2_U3879);
  nand ginst17964 (P2_U5745, P2_IR_REG_31__SCAN_IN, P2_SUB_1108_U21);
  nand ginst17965 (P2_U5746, P2_U3347, U64);
  nand ginst17966 (P2_U5747, P2_U3449, P2_U3945);
  not ginst17967 (P2_U5748, P2_U3450);
  nand ginst17968 (P2_U5749, P2_REG0_REG_7__SCAN_IN, P2_U3881);
  nand ginst17969 (P2_U5750, P2_U3966, P2_U4267);
  nand ginst17970 (P2_U5751, P2_IR_REG_8__SCAN_IN, P2_U3879);
  nand ginst17971 (P2_U5752, P2_IR_REG_31__SCAN_IN, P2_SUB_1108_U22);
  nand ginst17972 (P2_U5753, P2_U3347, U63);
  nand ginst17973 (P2_U5754, P2_U3452, P2_U3945);
  not ginst17974 (P2_U5755, P2_U3453);
  nand ginst17975 (P2_U5756, P2_REG0_REG_8__SCAN_IN, P2_U3881);
  nand ginst17976 (P2_U5757, P2_U3966, P2_U4286);
  nand ginst17977 (P2_U5758, P2_IR_REG_9__SCAN_IN, P2_U3879);
  nand ginst17978 (P2_U5759, P2_IR_REG_31__SCAN_IN, P2_SUB_1108_U99);
  nand ginst17979 (P2_U5760, P2_U3347, U62);
  nand ginst17980 (P2_U5761, P2_U3455, P2_U3945);
  not ginst17981 (P2_U5762, P2_U3456);
  nand ginst17982 (P2_U5763, P2_REG0_REG_9__SCAN_IN, P2_U3881);
  nand ginst17983 (P2_U5764, P2_U3966, P2_U4305);
  nand ginst17984 (P2_U5765, P2_IR_REG_10__SCAN_IN, P2_U3879);
  nand ginst17985 (P2_U5766, P2_IR_REG_31__SCAN_IN, P2_SUB_1108_U6);
  nand ginst17986 (P2_U5767, P2_U3347, U92);
  nand ginst17987 (P2_U5768, P2_U3458, P2_U3945);
  not ginst17988 (P2_U5769, P2_U3459);
  nand ginst17989 (P2_U5770, P2_REG0_REG_10__SCAN_IN, P2_U3881);
  nand ginst17990 (P2_U5771, P2_U3966, P2_U4324);
  nand ginst17991 (P2_U5772, P2_IR_REG_11__SCAN_IN, P2_U3879);
  nand ginst17992 (P2_U5773, P2_IR_REG_31__SCAN_IN, P2_SUB_1108_U7);
  nand ginst17993 (P2_U5774, P2_U3347, U91);
  nand ginst17994 (P2_U5775, P2_U3461, P2_U3945);
  not ginst17995 (P2_U5776, P2_U3462);
  nand ginst17996 (P2_U5777, P2_REG0_REG_11__SCAN_IN, P2_U3881);
  nand ginst17997 (P2_U5778, P2_U3966, P2_U4343);
  nand ginst17998 (P2_U5779, P2_IR_REG_12__SCAN_IN, P2_U3879);
  nand ginst17999 (P2_U5780, P2_IR_REG_31__SCAN_IN, P2_SUB_1108_U8);
  nand ginst18000 (P2_U5781, P2_U3347, U90);
  nand ginst18001 (P2_U5782, P2_U3464, P2_U3945);
  not ginst18002 (P2_U5783, P2_U3465);
  nand ginst18003 (P2_U5784, P2_REG0_REG_12__SCAN_IN, P2_U3881);
  nand ginst18004 (P2_U5785, P2_U3966, P2_U4362);
  nand ginst18005 (P2_U5786, P2_IR_REG_13__SCAN_IN, P2_U3879);
  nand ginst18006 (P2_U5787, P2_IR_REG_31__SCAN_IN, P2_SUB_1108_U127);
  nand ginst18007 (P2_U5788, P2_U3347, U89);
  nand ginst18008 (P2_U5789, P2_U3467, P2_U3945);
  not ginst18009 (P2_U5790, P2_U3468);
  nand ginst18010 (P2_U5791, P2_REG0_REG_13__SCAN_IN, P2_U3881);
  nand ginst18011 (P2_U5792, P2_U3966, P2_U4381);
  nand ginst18012 (P2_U5793, P2_IR_REG_14__SCAN_IN, P2_U3879);
  nand ginst18013 (P2_U5794, P2_IR_REG_31__SCAN_IN, P2_SUB_1108_U9);
  nand ginst18014 (P2_U5795, P2_U3347, U88);
  nand ginst18015 (P2_U5796, P2_U3470, P2_U3945);
  not ginst18016 (P2_U5797, P2_U3471);
  nand ginst18017 (P2_U5798, P2_REG0_REG_14__SCAN_IN, P2_U3881);
  nand ginst18018 (P2_U5799, P2_U3966, P2_U4400);
  nand ginst18019 (P2_U5800, P2_IR_REG_15__SCAN_IN, P2_U3879);
  nand ginst18020 (P2_U5801, P2_IR_REG_31__SCAN_IN, P2_SUB_1108_U10);
  nand ginst18021 (P2_U5802, P2_U3347, U87);
  nand ginst18022 (P2_U5803, P2_U3473, P2_U3945);
  not ginst18023 (P2_U5804, P2_U3474);
  nand ginst18024 (P2_U5805, P2_REG0_REG_15__SCAN_IN, P2_U3881);
  nand ginst18025 (P2_U5806, P2_U3966, P2_U4419);
  nand ginst18026 (P2_U5807, P2_IR_REG_16__SCAN_IN, P2_U3879);
  nand ginst18027 (P2_U5808, P2_IR_REG_31__SCAN_IN, P2_SUB_1108_U11);
  nand ginst18028 (P2_U5809, P2_U3347, U86);
  nand ginst18029 (P2_U5810, P2_U3476, P2_U3945);
  not ginst18030 (P2_U5811, P2_U3477);
  nand ginst18031 (P2_U5812, P2_REG0_REG_16__SCAN_IN, P2_U3881);
  nand ginst18032 (P2_U5813, P2_U3966, P2_U4438);
  nand ginst18033 (P2_U5814, P2_IR_REG_17__SCAN_IN, P2_U3879);
  nand ginst18034 (P2_U5815, P2_IR_REG_31__SCAN_IN, P2_SUB_1108_U125);
  nand ginst18035 (P2_U5816, P2_U3347, U85);
  nand ginst18036 (P2_U5817, P2_U3479, P2_U3945);
  not ginst18037 (P2_U5818, P2_U3480);
  nand ginst18038 (P2_U5819, P2_REG0_REG_17__SCAN_IN, P2_U3881);
  nand ginst18039 (P2_U5820, P2_U3966, P2_U4457);
  nand ginst18040 (P2_U5821, P2_IR_REG_18__SCAN_IN, P2_U3879);
  nand ginst18041 (P2_U5822, P2_IR_REG_31__SCAN_IN, P2_SUB_1108_U12);
  nand ginst18042 (P2_U5823, P2_U3347, U84);
  nand ginst18043 (P2_U5824, P2_U3482, P2_U3945);
  not ginst18044 (P2_U5825, P2_U3483);
  nand ginst18045 (P2_U5826, P2_REG0_REG_18__SCAN_IN, P2_U3881);
  nand ginst18046 (P2_U5827, P2_U3966, P2_U4476);
  nand ginst18047 (P2_U5828, P2_U3347, U83);
  nand ginst18048 (P2_U5829, P2_U3424, P2_U3945);
  not ginst18049 (P2_U5830, P2_U3485);
  nand ginst18050 (P2_U5831, P2_REG0_REG_19__SCAN_IN, P2_U3881);
  nand ginst18051 (P2_U5832, P2_U3966, P2_U4495);
  nand ginst18052 (P2_U5833, P2_REG0_REG_20__SCAN_IN, P2_U3881);
  nand ginst18053 (P2_U5834, P2_U3966, P2_U4514);
  nand ginst18054 (P2_U5835, P2_REG0_REG_21__SCAN_IN, P2_U3881);
  nand ginst18055 (P2_U5836, P2_U3966, P2_U4533);
  nand ginst18056 (P2_U5837, P2_REG0_REG_22__SCAN_IN, P2_U3881);
  nand ginst18057 (P2_U5838, P2_U3966, P2_U4552);
  nand ginst18058 (P2_U5839, P2_REG0_REG_23__SCAN_IN, P2_U3881);
  nand ginst18059 (P2_U5840, P2_U3966, P2_U4571);
  nand ginst18060 (P2_U5841, P2_REG0_REG_24__SCAN_IN, P2_U3881);
  nand ginst18061 (P2_U5842, P2_U3966, P2_U4590);
  nand ginst18062 (P2_U5843, P2_REG0_REG_25__SCAN_IN, P2_U3881);
  nand ginst18063 (P2_U5844, P2_U3966, P2_U4609);
  nand ginst18064 (P2_U5845, P2_REG0_REG_26__SCAN_IN, P2_U3881);
  nand ginst18065 (P2_U5846, P2_U3966, P2_U4628);
  nand ginst18066 (P2_U5847, P2_REG0_REG_27__SCAN_IN, P2_U3881);
  nand ginst18067 (P2_U5848, P2_U3966, P2_U4647);
  nand ginst18068 (P2_U5849, P2_REG0_REG_28__SCAN_IN, P2_U3881);
  nand ginst18069 (P2_U5850, P2_U3966, P2_U4666);
  nand ginst18070 (P2_U5851, P2_REG0_REG_29__SCAN_IN, P2_U3881);
  nand ginst18071 (P2_U5852, P2_U3966, P2_U4686);
  nand ginst18072 (P2_U5853, P2_REG0_REG_30__SCAN_IN, P2_U3881);
  nand ginst18073 (P2_U5854, P2_U3966, P2_U4693);
  nand ginst18074 (P2_U5855, P2_REG0_REG_31__SCAN_IN, P2_U3881);
  nand ginst18075 (P2_U5856, P2_U3966, P2_U4696);
  nand ginst18076 (P2_U5857, P2_REG1_REG_0__SCAN_IN, P2_U3882);
  nand ginst18077 (P2_U5858, P2_U3965, P2_U4129);
  nand ginst18078 (P2_U5859, P2_REG1_REG_1__SCAN_IN, P2_U3882);
  nand ginst18079 (P2_U5860, P2_U3965, P2_U4153);
  nand ginst18080 (P2_U5861, P2_REG1_REG_2__SCAN_IN, P2_U3882);
  nand ginst18081 (P2_U5862, P2_U3965, P2_U4172);
  nand ginst18082 (P2_U5863, P2_REG1_REG_3__SCAN_IN, P2_U3882);
  nand ginst18083 (P2_U5864, P2_U3965, P2_U4191);
  nand ginst18084 (P2_U5865, P2_REG1_REG_4__SCAN_IN, P2_U3882);
  nand ginst18085 (P2_U5866, P2_U3965, P2_U4210);
  nand ginst18086 (P2_U5867, P2_REG1_REG_5__SCAN_IN, P2_U3882);
  nand ginst18087 (P2_U5868, P2_U3965, P2_U4229);
  nand ginst18088 (P2_U5869, P2_REG1_REG_6__SCAN_IN, P2_U3882);
  nand ginst18089 (P2_U5870, P2_U3965, P2_U4248);
  nand ginst18090 (P2_U5871, P2_REG1_REG_7__SCAN_IN, P2_U3882);
  nand ginst18091 (P2_U5872, P2_U3965, P2_U4267);
  nand ginst18092 (P2_U5873, P2_REG1_REG_8__SCAN_IN, P2_U3882);
  nand ginst18093 (P2_U5874, P2_U3965, P2_U4286);
  nand ginst18094 (P2_U5875, P2_REG1_REG_9__SCAN_IN, P2_U3882);
  nand ginst18095 (P2_U5876, P2_U3965, P2_U4305);
  nand ginst18096 (P2_U5877, P2_REG1_REG_10__SCAN_IN, P2_U3882);
  nand ginst18097 (P2_U5878, P2_U3965, P2_U4324);
  nand ginst18098 (P2_U5879, P2_REG1_REG_11__SCAN_IN, P2_U3882);
  nand ginst18099 (P2_U5880, P2_U3965, P2_U4343);
  nand ginst18100 (P2_U5881, P2_REG1_REG_12__SCAN_IN, P2_U3882);
  nand ginst18101 (P2_U5882, P2_U3965, P2_U4362);
  nand ginst18102 (P2_U5883, P2_REG1_REG_13__SCAN_IN, P2_U3882);
  nand ginst18103 (P2_U5884, P2_U3965, P2_U4381);
  nand ginst18104 (P2_U5885, P2_REG1_REG_14__SCAN_IN, P2_U3882);
  nand ginst18105 (P2_U5886, P2_U3965, P2_U4400);
  nand ginst18106 (P2_U5887, P2_REG1_REG_15__SCAN_IN, P2_U3882);
  nand ginst18107 (P2_U5888, P2_U3965, P2_U4419);
  nand ginst18108 (P2_U5889, P2_REG1_REG_16__SCAN_IN, P2_U3882);
  nand ginst18109 (P2_U5890, P2_U3965, P2_U4438);
  nand ginst18110 (P2_U5891, P2_REG1_REG_17__SCAN_IN, P2_U3882);
  nand ginst18111 (P2_U5892, P2_U3965, P2_U4457);
  nand ginst18112 (P2_U5893, P2_REG1_REG_18__SCAN_IN, P2_U3882);
  nand ginst18113 (P2_U5894, P2_U3965, P2_U4476);
  nand ginst18114 (P2_U5895, P2_REG1_REG_19__SCAN_IN, P2_U3882);
  nand ginst18115 (P2_U5896, P2_U3965, P2_U4495);
  nand ginst18116 (P2_U5897, P2_REG1_REG_20__SCAN_IN, P2_U3882);
  nand ginst18117 (P2_U5898, P2_U3965, P2_U4514);
  nand ginst18118 (P2_U5899, P2_REG1_REG_21__SCAN_IN, P2_U3882);
  nand ginst18119 (P2_U5900, P2_U3965, P2_U4533);
  nand ginst18120 (P2_U5901, P2_REG1_REG_22__SCAN_IN, P2_U3882);
  nand ginst18121 (P2_U5902, P2_U3965, P2_U4552);
  nand ginst18122 (P2_U5903, P2_REG1_REG_23__SCAN_IN, P2_U3882);
  nand ginst18123 (P2_U5904, P2_U3965, P2_U4571);
  nand ginst18124 (P2_U5905, P2_REG1_REG_24__SCAN_IN, P2_U3882);
  nand ginst18125 (P2_U5906, P2_U3965, P2_U4590);
  nand ginst18126 (P2_U5907, P2_REG1_REG_25__SCAN_IN, P2_U3882);
  nand ginst18127 (P2_U5908, P2_U3965, P2_U4609);
  nand ginst18128 (P2_U5909, P2_REG1_REG_26__SCAN_IN, P2_U3882);
  nand ginst18129 (P2_U5910, P2_U3965, P2_U4628);
  nand ginst18130 (P2_U5911, P2_REG1_REG_27__SCAN_IN, P2_U3882);
  nand ginst18131 (P2_U5912, P2_U3965, P2_U4647);
  nand ginst18132 (P2_U5913, P2_REG1_REG_28__SCAN_IN, P2_U3882);
  nand ginst18133 (P2_U5914, P2_U3965, P2_U4666);
  nand ginst18134 (P2_U5915, P2_REG1_REG_29__SCAN_IN, P2_U3882);
  nand ginst18135 (P2_U5916, P2_U3965, P2_U4686);
  nand ginst18136 (P2_U5917, P2_REG1_REG_30__SCAN_IN, P2_U3882);
  nand ginst18137 (P2_U5918, P2_U3965, P2_U4693);
  nand ginst18138 (P2_U5919, P2_REG1_REG_31__SCAN_IN, P2_U3882);
  nand ginst18139 (P2_U5920, P2_U3965, P2_U4696);
  nand ginst18140 (P2_U5921, P2_REG2_REG_0__SCAN_IN, P2_U3391);
  nand ginst18141 (P2_U5922, P2_U3348, P2_U3964);
  nand ginst18142 (P2_U5923, P2_REG2_REG_1__SCAN_IN, P2_U3391);
  nand ginst18143 (P2_U5924, P2_U3349, P2_U3964);
  nand ginst18144 (P2_U5925, P2_REG2_REG_2__SCAN_IN, P2_U3391);
  nand ginst18145 (P2_U5926, P2_U3350, P2_U3964);
  nand ginst18146 (P2_U5927, P2_REG2_REG_3__SCAN_IN, P2_U3391);
  nand ginst18147 (P2_U5928, P2_U3351, P2_U3964);
  nand ginst18148 (P2_U5929, P2_REG2_REG_4__SCAN_IN, P2_U3391);
  nand ginst18149 (P2_U5930, P2_U3352, P2_U3964);
  nand ginst18150 (P2_U5931, P2_REG2_REG_5__SCAN_IN, P2_U3391);
  nand ginst18151 (P2_U5932, P2_U3353, P2_U3964);
  nand ginst18152 (P2_U5933, P2_REG2_REG_6__SCAN_IN, P2_U3391);
  nand ginst18153 (P2_U5934, P2_U3354, P2_U3964);
  nand ginst18154 (P2_U5935, P2_REG2_REG_7__SCAN_IN, P2_U3391);
  nand ginst18155 (P2_U5936, P2_U3355, P2_U3964);
  nand ginst18156 (P2_U5937, P2_REG2_REG_8__SCAN_IN, P2_U3391);
  nand ginst18157 (P2_U5938, P2_U3356, P2_U3964);
  nand ginst18158 (P2_U5939, P2_REG2_REG_9__SCAN_IN, P2_U3391);
  nand ginst18159 (P2_U5940, P2_U3357, P2_U3964);
  nand ginst18160 (P2_U5941, P2_REG2_REG_10__SCAN_IN, P2_U3391);
  nand ginst18161 (P2_U5942, P2_U3358, P2_U3964);
  nand ginst18162 (P2_U5943, P2_REG2_REG_11__SCAN_IN, P2_U3391);
  nand ginst18163 (P2_U5944, P2_U3359, P2_U3964);
  nand ginst18164 (P2_U5945, P2_REG2_REG_12__SCAN_IN, P2_U3391);
  nand ginst18165 (P2_U5946, P2_U3360, P2_U3964);
  nand ginst18166 (P2_U5947, P2_REG2_REG_13__SCAN_IN, P2_U3391);
  nand ginst18167 (P2_U5948, P2_U3361, P2_U3964);
  nand ginst18168 (P2_U5949, P2_REG2_REG_14__SCAN_IN, P2_U3391);
  nand ginst18169 (P2_U5950, P2_U3362, P2_U3964);
  nand ginst18170 (P2_U5951, P2_REG2_REG_15__SCAN_IN, P2_U3391);
  nand ginst18171 (P2_U5952, P2_U3363, P2_U3964);
  nand ginst18172 (P2_U5953, P2_REG2_REG_16__SCAN_IN, P2_U3391);
  nand ginst18173 (P2_U5954, P2_U3364, P2_U3964);
  nand ginst18174 (P2_U5955, P2_REG2_REG_17__SCAN_IN, P2_U3391);
  nand ginst18175 (P2_U5956, P2_U3365, P2_U3964);
  nand ginst18176 (P2_U5957, P2_REG2_REG_18__SCAN_IN, P2_U3391);
  nand ginst18177 (P2_U5958, P2_U3366, P2_U3964);
  nand ginst18178 (P2_U5959, P2_REG2_REG_19__SCAN_IN, P2_U3391);
  nand ginst18179 (P2_U5960, P2_U3367, P2_U3964);
  nand ginst18180 (P2_U5961, P2_REG2_REG_20__SCAN_IN, P2_U3391);
  nand ginst18181 (P2_U5962, P2_U3369, P2_U3964);
  nand ginst18182 (P2_U5963, P2_REG2_REG_21__SCAN_IN, P2_U3391);
  nand ginst18183 (P2_U5964, P2_U3371, P2_U3964);
  nand ginst18184 (P2_U5965, P2_REG2_REG_22__SCAN_IN, P2_U3391);
  nand ginst18185 (P2_U5966, P2_U3373, P2_U3964);
  nand ginst18186 (P2_U5967, P2_REG2_REG_23__SCAN_IN, P2_U3391);
  nand ginst18187 (P2_U5968, P2_U3375, P2_U3964);
  nand ginst18188 (P2_U5969, P2_REG2_REG_24__SCAN_IN, P2_U3391);
  nand ginst18189 (P2_U5970, P2_U3377, P2_U3964);
  nand ginst18190 (P2_U5971, P2_REG2_REG_25__SCAN_IN, P2_U3391);
  nand ginst18191 (P2_U5972, P2_U3379, P2_U3964);
  nand ginst18192 (P2_U5973, P2_REG2_REG_26__SCAN_IN, P2_U3391);
  nand ginst18193 (P2_U5974, P2_U3381, P2_U3964);
  nand ginst18194 (P2_U5975, P2_REG2_REG_27__SCAN_IN, P2_U3391);
  nand ginst18195 (P2_U5976, P2_U3383, P2_U3964);
  nand ginst18196 (P2_U5977, P2_REG2_REG_28__SCAN_IN, P2_U3391);
  nand ginst18197 (P2_U5978, P2_U3385, P2_U3964);
  nand ginst18198 (P2_U5979, P2_REG2_REG_29__SCAN_IN, P2_U3391);
  nand ginst18199 (P2_U5980, P2_U3387, P2_U3964);
  nand ginst18200 (P2_U5981, P2_REG2_REG_30__SCAN_IN, P2_U3391);
  nand ginst18201 (P2_U5982, P2_U3964, P2_U3968);
  nand ginst18202 (P2_U5983, P2_REG2_REG_31__SCAN_IN, P2_U3391);
  nand ginst18203 (P2_U5984, P2_U3964, P2_U3968);
  nand ginst18204 (P2_U5985, P2_DATAO_REG_0__SCAN_IN, P2_U3400);
  nand ginst18205 (P2_U5986, P2_U3079, P2_U3947);
  nand ginst18206 (P2_U5987, P2_DATAO_REG_1__SCAN_IN, P2_U3400);
  nand ginst18207 (P2_U5988, P2_U3080, P2_U3947);
  nand ginst18208 (P2_U5989, P2_DATAO_REG_2__SCAN_IN, P2_U3400);
  nand ginst18209 (P2_U5990, P2_U3070, P2_U3947);
  nand ginst18210 (P2_U5991, P2_DATAO_REG_3__SCAN_IN, P2_U3400);
  nand ginst18211 (P2_U5992, P2_U3066, P2_U3947);
  nand ginst18212 (P2_U5993, P2_DATAO_REG_4__SCAN_IN, P2_U3400);
  nand ginst18213 (P2_U5994, P2_U3062, P2_U3947);
  nand ginst18214 (P2_U5995, P2_DATAO_REG_5__SCAN_IN, P2_U3400);
  nand ginst18215 (P2_U5996, P2_U3069, P2_U3947);
  nand ginst18216 (P2_U5997, P2_DATAO_REG_6__SCAN_IN, P2_U3400);
  nand ginst18217 (P2_U5998, P2_U3073, P2_U3947);
  nand ginst18218 (P2_U5999, P2_DATAO_REG_7__SCAN_IN, P2_U3400);
  nand ginst18219 (P2_U6000, P2_U3072, P2_U3947);
  nand ginst18220 (P2_U6001, P2_DATAO_REG_8__SCAN_IN, P2_U3400);
  nand ginst18221 (P2_U6002, P2_U3086, P2_U3947);
  nand ginst18222 (P2_U6003, P2_DATAO_REG_9__SCAN_IN, P2_U3400);
  nand ginst18223 (P2_U6004, P2_U3085, P2_U3947);
  nand ginst18224 (P2_U6005, P2_DATAO_REG_10__SCAN_IN, P2_U3400);
  nand ginst18225 (P2_U6006, P2_U3064, P2_U3947);
  nand ginst18226 (P2_U6007, P2_DATAO_REG_11__SCAN_IN, P2_U3400);
  nand ginst18227 (P2_U6008, P2_U3065, P2_U3947);
  nand ginst18228 (P2_U6009, P2_DATAO_REG_12__SCAN_IN, P2_U3400);
  nand ginst18229 (P2_U6010, P2_U3074, P2_U3947);
  nand ginst18230 (P2_U6011, P2_DATAO_REG_13__SCAN_IN, P2_U3400);
  nand ginst18231 (P2_U6012, P2_U3082, P2_U3947);
  nand ginst18232 (P2_U6013, P2_DATAO_REG_14__SCAN_IN, P2_U3400);
  nand ginst18233 (P2_U6014, P2_U3081, P2_U3947);
  nand ginst18234 (P2_U6015, P2_DATAO_REG_15__SCAN_IN, P2_U3400);
  nand ginst18235 (P2_U6016, P2_U3076, P2_U3947);
  nand ginst18236 (P2_U6017, P2_DATAO_REG_16__SCAN_IN, P2_U3400);
  nand ginst18237 (P2_U6018, P2_U3075, P2_U3947);
  nand ginst18238 (P2_U6019, P2_DATAO_REG_17__SCAN_IN, P2_U3400);
  nand ginst18239 (P2_U6020, P2_U3071, P2_U3947);
  nand ginst18240 (P2_U6021, P2_DATAO_REG_18__SCAN_IN, P2_U3400);
  nand ginst18241 (P2_U6022, P2_U3084, P2_U3947);
  nand ginst18242 (P2_U6023, P2_DATAO_REG_19__SCAN_IN, P2_U3400);
  nand ginst18243 (P2_U6024, P2_U3083, P2_U3947);
  nand ginst18244 (P2_U6025, P2_DATAO_REG_20__SCAN_IN, P2_U3400);
  nand ginst18245 (P2_U6026, P2_U3078, P2_U3947);
  nand ginst18246 (P2_U6027, P2_DATAO_REG_21__SCAN_IN, P2_U3400);
  nand ginst18247 (P2_U6028, P2_U3077, P2_U3947);
  nand ginst18248 (P2_U6029, P2_DATAO_REG_22__SCAN_IN, P2_U3400);
  nand ginst18249 (P2_U6030, P2_U3063, P2_U3947);
  nand ginst18250 (P2_U6031, P2_DATAO_REG_23__SCAN_IN, P2_U3400);
  nand ginst18251 (P2_U6032, P2_U3068, P2_U3947);
  nand ginst18252 (P2_U6033, P2_DATAO_REG_24__SCAN_IN, P2_U3400);
  nand ginst18253 (P2_U6034, P2_U3067, P2_U3947);
  nand ginst18254 (P2_U6035, P2_DATAO_REG_25__SCAN_IN, P2_U3400);
  nand ginst18255 (P2_U6036, P2_U3060, P2_U3947);
  nand ginst18256 (P2_U6037, P2_DATAO_REG_26__SCAN_IN, P2_U3400);
  nand ginst18257 (P2_U6038, P2_U3059, P2_U3947);
  nand ginst18258 (P2_U6039, P2_DATAO_REG_27__SCAN_IN, P2_U3400);
  nand ginst18259 (P2_U6040, P2_U3055, P2_U3947);
  nand ginst18260 (P2_U6041, P2_DATAO_REG_28__SCAN_IN, P2_U3400);
  nand ginst18261 (P2_U6042, P2_U3056, P2_U3947);
  nand ginst18262 (P2_U6043, P2_DATAO_REG_29__SCAN_IN, P2_U3400);
  nand ginst18263 (P2_U6044, P2_U3057, P2_U3947);
  nand ginst18264 (P2_U6045, P2_DATAO_REG_30__SCAN_IN, P2_U3400);
  nand ginst18265 (P2_U6046, P2_U3061, P2_U3947);
  nand ginst18266 (P2_U6047, P2_DATAO_REG_31__SCAN_IN, P2_U3400);
  nand ginst18267 (P2_U6048, P2_U3058, P2_U3947);
  nand ginst18268 (P2_U6049, P2_R1312_U18, P2_U5157);
  nand ginst18269 (P2_U6050, P2_U3916, P2_U5161);
  nand ginst18270 (P2_U6051, P2_U3403, P2_U5658);
  nand ginst18271 (P2_U6052, P2_U3415, P2_U3420);
  nand ginst18272 (P2_U6053, P2_U3057, P2_U3960);
  nand ginst18273 (P2_U6054, P2_U3386, P2_U4652);
  nand ginst18274 (P2_U6055, P2_U6053, P2_U6054);
  nand ginst18275 (P2_U6056, P2_U3056, P2_U3949);
  nand ginst18276 (P2_U6057, P2_U3384, P2_U4633);
  nand ginst18277 (P2_U6058, P2_U6056, P2_U6057);
  nand ginst18278 (P2_U6059, P2_U3055, P2_U3950);
  nand ginst18279 (P2_U6060, P2_U3382, P2_U4614);
  nand ginst18280 (P2_U6061, P2_U6059, P2_U6060);
  nand ginst18281 (P2_U6062, P2_U3067, P2_U3953);
  nand ginst18282 (P2_U6063, P2_U3376, P2_U4557);
  nand ginst18283 (P2_U6064, P2_U6062, P2_U6063);
  nand ginst18284 (P2_U6065, P2_U3068, P2_U3954);
  nand ginst18285 (P2_U6066, P2_U3374, P2_U4538);
  nand ginst18286 (P2_U6067, P2_U6065, P2_U6066);
  nand ginst18287 (P2_U6068, P2_U3077, P2_U3956);
  nand ginst18288 (P2_U6069, P2_U3370, P2_U4500);
  nand ginst18289 (P2_U6070, P2_U6068, P2_U6069);
  nand ginst18290 (P2_U6071, P2_U3063, P2_U3955);
  nand ginst18291 (P2_U6072, P2_U3372, P2_U4519);
  nand ginst18292 (P2_U6073, P2_U6071, P2_U6072);
  nand ginst18293 (P2_U6074, P2_U3060, P2_U3952);
  nand ginst18294 (P2_U6075, P2_U3378, P2_U4576);
  nand ginst18295 (P2_U6076, P2_U6074, P2_U6075);
  nand ginst18296 (P2_U6077, P2_U3059, P2_U3951);
  nand ginst18297 (P2_U6078, P2_U3380, P2_U4595);
  nand ginst18298 (P2_U6079, P2_U6077, P2_U6078);
  nand ginst18299 (P2_U6080, P2_U3061, P2_U3959);
  nand ginst18300 (P2_U6081, P2_U3388, P2_U4670);
  nand ginst18301 (P2_U6082, P2_U6080, P2_U6081);
  nand ginst18302 (P2_U6083, P2_U3058, P2_U3958);
  nand ginst18303 (P2_U6084, P2_U3389, P2_U4690);
  nand ginst18304 (P2_U6085, P2_U6083, P2_U6084);
  nand ginst18305 (P2_U6086, P2_U4367, P2_U5797);
  nand ginst18306 (P2_U6087, P2_U3081, P2_U3471);
  nand ginst18307 (P2_U6088, P2_U6086, P2_U6087);
  nand ginst18308 (P2_U6089, P2_U4115, P2_U5706);
  nand ginst18309 (P2_U6090, P2_U3080, P2_U3432);
  nand ginst18310 (P2_U6091, P2_U6089, P2_U6090);
  nand ginst18311 (P2_U6092, P2_U4139, P2_U5691);
  nand ginst18312 (P2_U6093, P2_U3079, P2_U3427);
  nand ginst18313 (P2_U6094, P2_U6092, P2_U6093);
  nand ginst18314 (P2_U6095, P2_U4386, P2_U5804);
  nand ginst18315 (P2_U6096, P2_U3076, P2_U3474);
  nand ginst18316 (P2_U6097, P2_U6095, P2_U6096);
  nand ginst18317 (P2_U6098, P2_U4253, P2_U5755);
  nand ginst18318 (P2_U6099, P2_U3086, P2_U3453);
  nand ginst18319 (P2_U6100, P2_U6098, P2_U6099);
  nand ginst18320 (P2_U6101, P2_U4272, P2_U5762);
  nand ginst18321 (P2_U6102, P2_U3085, P2_U3456);
  nand ginst18322 (P2_U6103, P2_U6101, P2_U6102);
  nand ginst18323 (P2_U6104, P2_U4348, P2_U5790);
  nand ginst18324 (P2_U6105, P2_U3082, P2_U3468);
  nand ginst18325 (P2_U6106, P2_U6104, P2_U6105);
  nand ginst18326 (P2_U6107, P2_U4443, P2_U5825);
  nand ginst18327 (P2_U6108, P2_U3084, P2_U3483);
  nand ginst18328 (P2_U6109, P2_U6107, P2_U6108);
  nand ginst18329 (P2_U6110, P2_U4405, P2_U5811);
  nand ginst18330 (P2_U6111, P2_U3075, P2_U3477);
  nand ginst18331 (P2_U6112, P2_U6110, P2_U6111);
  nand ginst18332 (P2_U6113, P2_U4329, P2_U5783);
  nand ginst18333 (P2_U6114, P2_U3074, P2_U3465);
  nand ginst18334 (P2_U6115, P2_U6113, P2_U6114);
  nand ginst18335 (P2_U6116, P2_U4215, P2_U5741);
  nand ginst18336 (P2_U6117, P2_U3073, P2_U3447);
  nand ginst18337 (P2_U6118, P2_U6116, P2_U6117);
  nand ginst18338 (P2_U6119, P2_U4234, P2_U5748);
  nand ginst18339 (P2_U6120, P2_U3072, P2_U3450);
  nand ginst18340 (P2_U6121, P2_U6119, P2_U6120);
  nand ginst18341 (P2_U6122, P2_U4196, P2_U5734);
  nand ginst18342 (P2_U6123, P2_U3069, P2_U3444);
  nand ginst18343 (P2_U6124, P2_U6122, P2_U6123);
  nand ginst18344 (P2_U6125, P2_U4158, P2_U5720);
  nand ginst18345 (P2_U6126, P2_U3066, P2_U3438);
  nand ginst18346 (P2_U6127, P2_U6125, P2_U6126);
  nand ginst18347 (P2_U6128, P2_U4134, P2_U5713);
  nand ginst18348 (P2_U6129, P2_U3070, P2_U3435);
  nand ginst18349 (P2_U6130, P2_U6128, P2_U6129);
  nand ginst18350 (P2_U6131, P2_U4424, P2_U5818);
  nand ginst18351 (P2_U6132, P2_U3071, P2_U3480);
  nand ginst18352 (P2_U6133, P2_U6131, P2_U6132);
  nand ginst18353 (P2_U6134, P2_U4462, P2_U5830);
  nand ginst18354 (P2_U6135, P2_U3083, P2_U3485);
  nand ginst18355 (P2_U6136, P2_U6134, P2_U6135);
  nand ginst18356 (P2_U6137, P2_U4177, P2_U5727);
  nand ginst18357 (P2_U6138, P2_U3062, P2_U3441);
  nand ginst18358 (P2_U6139, P2_U6137, P2_U6138);
  nand ginst18359 (P2_U6140, P2_U4310, P2_U5776);
  nand ginst18360 (P2_U6141, P2_U3065, P2_U3462);
  nand ginst18361 (P2_U6142, P2_U6140, P2_U6141);
  nand ginst18362 (P2_U6143, P2_U4291, P2_U5769);
  nand ginst18363 (P2_U6144, P2_U3064, P2_U3459);
  nand ginst18364 (P2_U6145, P2_U6143, P2_U6144);
  nand ginst18365 (P2_U6146, P2_U3078, P2_U3957);
  nand ginst18366 (P2_U6147, P2_U3368, P2_U4481);
  nand ginst18367 (P2_U6148, P2_U6146, P2_U6147);
  nand ginst18368 (P2_U6149, P2_U3940, P2_U5156);
  nand ginst18369 (P2_U6150, P2_U3918, P2_U3942);
  and ginst18370 (P3_R1054_U10, P3_R1054_U100, P3_R1054_U174);
  nand ginst18371 (P3_R1054_U100, P3_R1054_U56, P3_U3433);
  nand ginst18372 (P3_R1054_U101, P3_R1054_U24, P3_U3394);
  nand ginst18373 (P3_R1054_U102, P3_R1054_U31, P3_U3403);
  nand ginst18374 (P3_R1054_U103, P3_R1054_U35, P3_U3409);
  not ginst18375 (P3_R1054_U104, P3_R1054_U58);
  not ginst18376 (P3_R1054_U105, P3_R1054_U33);
  not ginst18377 (P3_R1054_U106, P3_R1054_U47);
  not ginst18378 (P3_R1054_U107, P3_R1054_U21);
  nand ginst18379 (P3_R1054_U108, P3_R1054_U107, P3_R1054_U22);
  nand ginst18380 (P3_R1054_U109, P3_R1054_U108, P3_R1054_U88);
  and ginst18381 (P3_R1054_U11, P3_R1054_U175, P3_R1054_U176);
  nand ginst18382 (P3_R1054_U110, P3_R1054_U21, P3_U3573);
  not ginst18383 (P3_R1054_U111, P3_R1054_U42);
  nand ginst18384 (P3_R1054_U112, P3_R1054_U26, P3_U3397);
  nand ginst18385 (P3_R1054_U113, P3_R1054_U101, P3_R1054_U112, P3_R1054_U42);
  nand ginst18386 (P3_R1054_U114, P3_R1054_U25, P3_R1054_U26);
  nand ginst18387 (P3_R1054_U115, P3_R1054_U114, P3_R1054_U23);
  nand ginst18388 (P3_R1054_U116, P3_R1054_U97, P3_U3561);
  not ginst18389 (P3_R1054_U117, P3_R1054_U87);
  nand ginst18390 (P3_R1054_U118, P3_R1054_U30, P3_U3406);
  nand ginst18391 (P3_R1054_U119, P3_R1054_U27, P3_U3558);
  nand ginst18392 (P3_R1054_U12, P3_R1054_U207, P3_R1054_U210);
  nand ginst18393 (P3_R1054_U120, P3_R1054_U28, P3_U3559);
  nand ginst18394 (P3_R1054_U121, P3_R1054_U105, P3_R1054_U6);
  nand ginst18395 (P3_R1054_U122, P3_R1054_U121, P3_R1054_U7);
  nand ginst18396 (P3_R1054_U123, P3_R1054_U32, P3_U3400);
  nand ginst18397 (P3_R1054_U124, P3_R1054_U30, P3_U3406);
  nand ginst18398 (P3_R1054_U125, P3_R1054_U123, P3_R1054_U6, P3_R1054_U87);
  nand ginst18399 (P3_R1054_U126, P3_R1054_U122, P3_R1054_U124);
  not ginst18400 (P3_R1054_U127, P3_R1054_U40);
  nand ginst18401 (P3_R1054_U128, P3_R1054_U37, P3_U3412);
  nand ginst18402 (P3_R1054_U129, P3_R1054_U103, P3_R1054_U128, P3_R1054_U40);
  nand ginst18403 (P3_R1054_U13, P3_R1054_U196, P3_R1054_U199);
  nand ginst18404 (P3_R1054_U130, P3_R1054_U36, P3_R1054_U37);
  nand ginst18405 (P3_R1054_U131, P3_R1054_U130, P3_R1054_U34);
  nand ginst18406 (P3_R1054_U132, P3_R1054_U98, P3_U3556);
  not ginst18407 (P3_R1054_U133, P3_R1054_U86);
  nand ginst18408 (P3_R1054_U134, P3_R1054_U39, P3_U3415);
  nand ginst18409 (P3_R1054_U135, P3_R1054_U134, P3_R1054_U47);
  nand ginst18410 (P3_R1054_U136, P3_R1054_U127, P3_R1054_U36);
  nand ginst18411 (P3_R1054_U137, P3_R1054_U103, P3_R1054_U136, P3_R1054_U222);
  nand ginst18412 (P3_R1054_U138, P3_R1054_U103, P3_R1054_U40);
  nand ginst18413 (P3_R1054_U139, P3_R1054_U138, P3_R1054_U218, P3_R1054_U219, P3_R1054_U36);
  nand ginst18414 (P3_R1054_U14, P3_R1054_U153, P3_R1054_U155);
  nand ginst18415 (P3_R1054_U140, P3_R1054_U103, P3_R1054_U36);
  nand ginst18416 (P3_R1054_U141, P3_R1054_U123, P3_R1054_U87);
  not ginst18417 (P3_R1054_U142, P3_R1054_U41);
  nand ginst18418 (P3_R1054_U143, P3_R1054_U28, P3_U3559);
  nand ginst18419 (P3_R1054_U144, P3_R1054_U142, P3_R1054_U143);
  nand ginst18420 (P3_R1054_U145, P3_R1054_U102, P3_R1054_U144, P3_R1054_U229);
  nand ginst18421 (P3_R1054_U146, P3_R1054_U102, P3_R1054_U41);
  nand ginst18422 (P3_R1054_U147, P3_R1054_U30, P3_U3406);
  nand ginst18423 (P3_R1054_U148, P3_R1054_U146, P3_R1054_U147, P3_R1054_U7);
  nand ginst18424 (P3_R1054_U149, P3_R1054_U28, P3_U3559);
  nand ginst18425 (P3_R1054_U15, P3_R1054_U145, P3_R1054_U148);
  nand ginst18426 (P3_R1054_U150, P3_R1054_U102, P3_R1054_U149);
  nand ginst18427 (P3_R1054_U151, P3_R1054_U123, P3_R1054_U33);
  nand ginst18428 (P3_R1054_U152, P3_R1054_U111, P3_R1054_U25);
  nand ginst18429 (P3_R1054_U153, P3_R1054_U101, P3_R1054_U152, P3_R1054_U242);
  nand ginst18430 (P3_R1054_U154, P3_R1054_U101, P3_R1054_U42);
  nand ginst18431 (P3_R1054_U155, P3_R1054_U154, P3_R1054_U238, P3_R1054_U239, P3_R1054_U25);
  nand ginst18432 (P3_R1054_U156, P3_R1054_U101, P3_R1054_U25);
  nand ginst18433 (P3_R1054_U157, P3_R1054_U45, P3_U3421);
  nand ginst18434 (P3_R1054_U158, P3_R1054_U43, P3_U3571);
  nand ginst18435 (P3_R1054_U159, P3_R1054_U44, P3_U3572);
  nand ginst18436 (P3_R1054_U16, P3_R1054_U137, P3_R1054_U139);
  nand ginst18437 (P3_R1054_U160, P3_R1054_U106, P3_R1054_U8);
  nand ginst18438 (P3_R1054_U161, P3_R1054_U160, P3_R1054_U9);
  nand ginst18439 (P3_R1054_U162, P3_R1054_U45, P3_U3421);
  nand ginst18440 (P3_R1054_U163, P3_R1054_U134, P3_R1054_U8, P3_R1054_U86);
  nand ginst18441 (P3_R1054_U164, P3_R1054_U161, P3_R1054_U162);
  not ginst18442 (P3_R1054_U165, P3_R1054_U96);
  nand ginst18443 (P3_R1054_U166, P3_R1054_U49, P3_U3424);
  nand ginst18444 (P3_R1054_U167, P3_R1054_U166, P3_R1054_U96);
  nand ginst18445 (P3_R1054_U168, P3_R1054_U48, P3_U3570);
  not ginst18446 (P3_R1054_U169, P3_R1054_U95);
  nand ginst18447 (P3_R1054_U17, P3_R1054_U21, P3_R1054_U213);
  nand ginst18448 (P3_R1054_U170, P3_R1054_U51, P3_U3427);
  nand ginst18449 (P3_R1054_U171, P3_R1054_U170, P3_R1054_U95);
  nand ginst18450 (P3_R1054_U172, P3_R1054_U50, P3_U3569);
  not ginst18451 (P3_R1054_U173, P3_R1054_U94);
  nand ginst18452 (P3_R1054_U174, P3_R1054_U55, P3_U3436);
  nand ginst18453 (P3_R1054_U175, P3_R1054_U52, P3_U3566);
  nand ginst18454 (P3_R1054_U176, P3_R1054_U53, P3_U3567);
  nand ginst18455 (P3_R1054_U177, P3_R1054_U10, P3_R1054_U104);
  nand ginst18456 (P3_R1054_U178, P3_R1054_U11, P3_R1054_U177);
  nand ginst18457 (P3_R1054_U179, P3_R1054_U57, P3_U3430);
  not ginst18458 (P3_R1054_U18, P3_U3409);
  nand ginst18459 (P3_R1054_U180, P3_R1054_U55, P3_U3436);
  nand ginst18460 (P3_R1054_U181, P3_R1054_U10, P3_R1054_U179, P3_R1054_U94);
  nand ginst18461 (P3_R1054_U182, P3_R1054_U178, P3_R1054_U180);
  not ginst18462 (P3_R1054_U183, P3_R1054_U93);
  nand ginst18463 (P3_R1054_U184, P3_R1054_U60, P3_U3439);
  nand ginst18464 (P3_R1054_U185, P3_R1054_U184, P3_R1054_U93);
  nand ginst18465 (P3_R1054_U186, P3_R1054_U59, P3_U3565);
  not ginst18466 (P3_R1054_U187, P3_R1054_U61);
  nand ginst18467 (P3_R1054_U188, P3_R1054_U187, P3_R1054_U62);
  nand ginst18468 (P3_R1054_U189, P3_R1054_U188, P3_R1054_U92);
  not ginst18469 (P3_R1054_U19, P3_U3394);
  nand ginst18470 (P3_R1054_U190, P3_R1054_U61, P3_U3564);
  not ginst18471 (P3_R1054_U191, P3_R1054_U91);
  nand ginst18472 (P3_R1054_U192, P3_R1054_U179, P3_R1054_U94);
  not ginst18473 (P3_R1054_U193, P3_R1054_U63);
  nand ginst18474 (P3_R1054_U194, P3_R1054_U53, P3_U3567);
  nand ginst18475 (P3_R1054_U195, P3_R1054_U193, P3_R1054_U194);
  nand ginst18476 (P3_R1054_U196, P3_R1054_U100, P3_R1054_U195, P3_R1054_U269);
  nand ginst18477 (P3_R1054_U197, P3_R1054_U100, P3_R1054_U63);
  nand ginst18478 (P3_R1054_U198, P3_R1054_U55, P3_U3436);
  nand ginst18479 (P3_R1054_U199, P3_R1054_U11, P3_R1054_U197, P3_R1054_U198);
  not ginst18480 (P3_R1054_U20, P3_U3386);
  nand ginst18481 (P3_R1054_U200, P3_R1054_U53, P3_U3567);
  nand ginst18482 (P3_R1054_U201, P3_R1054_U100, P3_R1054_U200);
  nand ginst18483 (P3_R1054_U202, P3_R1054_U179, P3_R1054_U58);
  nand ginst18484 (P3_R1054_U203, P3_R1054_U134, P3_R1054_U86);
  not ginst18485 (P3_R1054_U204, P3_R1054_U64);
  nand ginst18486 (P3_R1054_U205, P3_R1054_U44, P3_U3572);
  nand ginst18487 (P3_R1054_U206, P3_R1054_U204, P3_R1054_U205);
  nand ginst18488 (P3_R1054_U207, P3_R1054_U206, P3_R1054_U290, P3_R1054_U99);
  nand ginst18489 (P3_R1054_U208, P3_R1054_U64, P3_R1054_U99);
  nand ginst18490 (P3_R1054_U209, P3_R1054_U45, P3_U3421);
  nand ginst18491 (P3_R1054_U21, P3_R1054_U65, P3_U3386);
  nand ginst18492 (P3_R1054_U210, P3_R1054_U208, P3_R1054_U209, P3_R1054_U9);
  nand ginst18493 (P3_R1054_U211, P3_R1054_U44, P3_U3572);
  nand ginst18494 (P3_R1054_U212, P3_R1054_U211, P3_R1054_U99);
  nand ginst18495 (P3_R1054_U213, P3_R1054_U20, P3_U3574);
  nand ginst18496 (P3_R1054_U214, P3_R1054_U39, P3_U3415);
  nand ginst18497 (P3_R1054_U215, P3_R1054_U38, P3_U3555);
  nand ginst18498 (P3_R1054_U216, P3_R1054_U135, P3_R1054_U86);
  nand ginst18499 (P3_R1054_U217, P3_R1054_U133, P3_R1054_U214, P3_R1054_U215);
  nand ginst18500 (P3_R1054_U218, P3_R1054_U37, P3_U3412);
  nand ginst18501 (P3_R1054_U219, P3_R1054_U34, P3_U3556);
  not ginst18502 (P3_R1054_U22, P3_U3573);
  nand ginst18503 (P3_R1054_U220, P3_R1054_U37, P3_U3412);
  nand ginst18504 (P3_R1054_U221, P3_R1054_U34, P3_U3556);
  nand ginst18505 (P3_R1054_U222, P3_R1054_U220, P3_R1054_U221);
  nand ginst18506 (P3_R1054_U223, P3_R1054_U35, P3_U3409);
  nand ginst18507 (P3_R1054_U224, P3_R1054_U18, P3_U3557);
  nand ginst18508 (P3_R1054_U225, P3_R1054_U140, P3_R1054_U40);
  nand ginst18509 (P3_R1054_U226, P3_R1054_U127, P3_R1054_U223, P3_R1054_U224);
  nand ginst18510 (P3_R1054_U227, P3_R1054_U30, P3_U3406);
  nand ginst18511 (P3_R1054_U228, P3_R1054_U27, P3_U3558);
  nand ginst18512 (P3_R1054_U229, P3_R1054_U227, P3_R1054_U228);
  not ginst18513 (P3_R1054_U23, P3_U3397);
  nand ginst18514 (P3_R1054_U230, P3_R1054_U31, P3_U3403);
  nand ginst18515 (P3_R1054_U231, P3_R1054_U28, P3_U3559);
  nand ginst18516 (P3_R1054_U232, P3_R1054_U150, P3_R1054_U41);
  nand ginst18517 (P3_R1054_U233, P3_R1054_U142, P3_R1054_U230, P3_R1054_U231);
  nand ginst18518 (P3_R1054_U234, P3_R1054_U32, P3_U3400);
  nand ginst18519 (P3_R1054_U235, P3_R1054_U29, P3_U3560);
  nand ginst18520 (P3_R1054_U236, P3_R1054_U151, P3_R1054_U87);
  nand ginst18521 (P3_R1054_U237, P3_R1054_U117, P3_R1054_U234, P3_R1054_U235);
  nand ginst18522 (P3_R1054_U238, P3_R1054_U26, P3_U3397);
  nand ginst18523 (P3_R1054_U239, P3_R1054_U23, P3_U3561);
  not ginst18524 (P3_R1054_U24, P3_U3562);
  nand ginst18525 (P3_R1054_U240, P3_R1054_U26, P3_U3397);
  nand ginst18526 (P3_R1054_U241, P3_R1054_U23, P3_U3561);
  nand ginst18527 (P3_R1054_U242, P3_R1054_U240, P3_R1054_U241);
  nand ginst18528 (P3_R1054_U243, P3_R1054_U24, P3_U3394);
  nand ginst18529 (P3_R1054_U244, P3_R1054_U19, P3_U3562);
  nand ginst18530 (P3_R1054_U245, P3_R1054_U156, P3_R1054_U42);
  nand ginst18531 (P3_R1054_U246, P3_R1054_U111, P3_R1054_U243, P3_R1054_U244);
  nand ginst18532 (P3_R1054_U247, P3_R1054_U22, P3_U3391);
  nand ginst18533 (P3_R1054_U248, P3_R1054_U88, P3_U3573);
  not ginst18534 (P3_R1054_U249, P3_R1054_U80);
  nand ginst18535 (P3_R1054_U25, P3_R1054_U19, P3_U3562);
  nand ginst18536 (P3_R1054_U250, P3_R1054_U107, P3_R1054_U249);
  nand ginst18537 (P3_R1054_U251, P3_R1054_U21, P3_R1054_U80);
  nand ginst18538 (P3_R1054_U252, P3_R1054_U90, P3_U3379);
  nand ginst18539 (P3_R1054_U253, P3_R1054_U89, P3_U3563);
  not ginst18540 (P3_R1054_U254, P3_R1054_U81);
  nand ginst18541 (P3_R1054_U255, P3_R1054_U191, P3_R1054_U254);
  nand ginst18542 (P3_R1054_U256, P3_R1054_U81, P3_R1054_U91);
  nand ginst18543 (P3_R1054_U257, P3_R1054_U62, P3_U3442);
  nand ginst18544 (P3_R1054_U258, P3_R1054_U92, P3_U3564);
  not ginst18545 (P3_R1054_U259, P3_R1054_U82);
  not ginst18546 (P3_R1054_U26, P3_U3561);
  nand ginst18547 (P3_R1054_U260, P3_R1054_U187, P3_R1054_U259);
  nand ginst18548 (P3_R1054_U261, P3_R1054_U61, P3_R1054_U82);
  nand ginst18549 (P3_R1054_U262, P3_R1054_U60, P3_U3439);
  nand ginst18550 (P3_R1054_U263, P3_R1054_U59, P3_U3565);
  not ginst18551 (P3_R1054_U264, P3_R1054_U83);
  nand ginst18552 (P3_R1054_U265, P3_R1054_U183, P3_R1054_U264);
  nand ginst18553 (P3_R1054_U266, P3_R1054_U83, P3_R1054_U93);
  nand ginst18554 (P3_R1054_U267, P3_R1054_U55, P3_U3436);
  nand ginst18555 (P3_R1054_U268, P3_R1054_U52, P3_U3566);
  nand ginst18556 (P3_R1054_U269, P3_R1054_U267, P3_R1054_U268);
  not ginst18557 (P3_R1054_U27, P3_U3406);
  nand ginst18558 (P3_R1054_U270, P3_R1054_U56, P3_U3433);
  nand ginst18559 (P3_R1054_U271, P3_R1054_U53, P3_U3567);
  nand ginst18560 (P3_R1054_U272, P3_R1054_U201, P3_R1054_U63);
  nand ginst18561 (P3_R1054_U273, P3_R1054_U193, P3_R1054_U270, P3_R1054_U271);
  nand ginst18562 (P3_R1054_U274, P3_R1054_U57, P3_U3430);
  nand ginst18563 (P3_R1054_U275, P3_R1054_U54, P3_U3568);
  nand ginst18564 (P3_R1054_U276, P3_R1054_U202, P3_R1054_U94);
  nand ginst18565 (P3_R1054_U277, P3_R1054_U173, P3_R1054_U274, P3_R1054_U275);
  nand ginst18566 (P3_R1054_U278, P3_R1054_U51, P3_U3427);
  nand ginst18567 (P3_R1054_U279, P3_R1054_U50, P3_U3569);
  not ginst18568 (P3_R1054_U28, P3_U3403);
  not ginst18569 (P3_R1054_U280, P3_R1054_U84);
  nand ginst18570 (P3_R1054_U281, P3_R1054_U169, P3_R1054_U280);
  nand ginst18571 (P3_R1054_U282, P3_R1054_U84, P3_R1054_U95);
  nand ginst18572 (P3_R1054_U283, P3_R1054_U49, P3_U3424);
  nand ginst18573 (P3_R1054_U284, P3_R1054_U48, P3_U3570);
  not ginst18574 (P3_R1054_U285, P3_R1054_U85);
  nand ginst18575 (P3_R1054_U286, P3_R1054_U165, P3_R1054_U285);
  nand ginst18576 (P3_R1054_U287, P3_R1054_U85, P3_R1054_U96);
  nand ginst18577 (P3_R1054_U288, P3_R1054_U45, P3_U3421);
  nand ginst18578 (P3_R1054_U289, P3_R1054_U43, P3_U3571);
  not ginst18579 (P3_R1054_U29, P3_U3400);
  nand ginst18580 (P3_R1054_U290, P3_R1054_U288, P3_R1054_U289);
  nand ginst18581 (P3_R1054_U291, P3_R1054_U46, P3_U3418);
  nand ginst18582 (P3_R1054_U292, P3_R1054_U44, P3_U3572);
  nand ginst18583 (P3_R1054_U293, P3_R1054_U212, P3_R1054_U64);
  nand ginst18584 (P3_R1054_U294, P3_R1054_U204, P3_R1054_U291, P3_R1054_U292);
  not ginst18585 (P3_R1054_U30, P3_U3558);
  not ginst18586 (P3_R1054_U31, P3_U3559);
  not ginst18587 (P3_R1054_U32, P3_U3560);
  nand ginst18588 (P3_R1054_U33, P3_R1054_U29, P3_U3560);
  not ginst18589 (P3_R1054_U34, P3_U3412);
  not ginst18590 (P3_R1054_U35, P3_U3557);
  nand ginst18591 (P3_R1054_U36, P3_R1054_U18, P3_U3557);
  not ginst18592 (P3_R1054_U37, P3_U3556);
  not ginst18593 (P3_R1054_U38, P3_U3415);
  not ginst18594 (P3_R1054_U39, P3_U3555);
  nand ginst18595 (P3_R1054_U40, P3_R1054_U125, P3_R1054_U126);
  nand ginst18596 (P3_R1054_U41, P3_R1054_U141, P3_R1054_U33);
  nand ginst18597 (P3_R1054_U42, P3_R1054_U109, P3_R1054_U110);
  not ginst18598 (P3_R1054_U43, P3_U3421);
  not ginst18599 (P3_R1054_U44, P3_U3418);
  not ginst18600 (P3_R1054_U45, P3_U3571);
  not ginst18601 (P3_R1054_U46, P3_U3572);
  nand ginst18602 (P3_R1054_U47, P3_R1054_U38, P3_U3555);
  not ginst18603 (P3_R1054_U48, P3_U3424);
  not ginst18604 (P3_R1054_U49, P3_U3570);
  not ginst18605 (P3_R1054_U50, P3_U3427);
  not ginst18606 (P3_R1054_U51, P3_U3569);
  not ginst18607 (P3_R1054_U52, P3_U3436);
  not ginst18608 (P3_R1054_U53, P3_U3433);
  not ginst18609 (P3_R1054_U54, P3_U3430);
  not ginst18610 (P3_R1054_U55, P3_U3566);
  not ginst18611 (P3_R1054_U56, P3_U3567);
  not ginst18612 (P3_R1054_U57, P3_U3568);
  nand ginst18613 (P3_R1054_U58, P3_R1054_U54, P3_U3568);
  not ginst18614 (P3_R1054_U59, P3_U3439);
  and ginst18615 (P3_R1054_U6, P3_R1054_U102, P3_R1054_U118);
  not ginst18616 (P3_R1054_U60, P3_U3565);
  nand ginst18617 (P3_R1054_U61, P3_R1054_U185, P3_R1054_U186);
  not ginst18618 (P3_R1054_U62, P3_U3564);
  nand ginst18619 (P3_R1054_U63, P3_R1054_U192, P3_R1054_U58);
  nand ginst18620 (P3_R1054_U64, P3_R1054_U203, P3_R1054_U47);
  not ginst18621 (P3_R1054_U65, P3_U3574);
  nand ginst18622 (P3_R1054_U66, P3_R1054_U250, P3_R1054_U251);
  nand ginst18623 (P3_R1054_U67, P3_R1054_U255, P3_R1054_U256);
  nand ginst18624 (P3_R1054_U68, P3_R1054_U260, P3_R1054_U261);
  nand ginst18625 (P3_R1054_U69, P3_R1054_U265, P3_R1054_U266);
  and ginst18626 (P3_R1054_U7, P3_R1054_U119, P3_R1054_U120);
  nand ginst18627 (P3_R1054_U70, P3_R1054_U281, P3_R1054_U282);
  nand ginst18628 (P3_R1054_U71, P3_R1054_U286, P3_R1054_U287);
  nand ginst18629 (P3_R1054_U72, P3_R1054_U216, P3_R1054_U217);
  nand ginst18630 (P3_R1054_U73, P3_R1054_U225, P3_R1054_U226);
  nand ginst18631 (P3_R1054_U74, P3_R1054_U232, P3_R1054_U233);
  nand ginst18632 (P3_R1054_U75, P3_R1054_U236, P3_R1054_U237);
  nand ginst18633 (P3_R1054_U76, P3_R1054_U245, P3_R1054_U246);
  nand ginst18634 (P3_R1054_U77, P3_R1054_U272, P3_R1054_U273);
  nand ginst18635 (P3_R1054_U78, P3_R1054_U276, P3_R1054_U277);
  nand ginst18636 (P3_R1054_U79, P3_R1054_U293, P3_R1054_U294);
  and ginst18637 (P3_R1054_U8, P3_R1054_U157, P3_R1054_U99);
  nand ginst18638 (P3_R1054_U80, P3_R1054_U247, P3_R1054_U248);
  nand ginst18639 (P3_R1054_U81, P3_R1054_U252, P3_R1054_U253);
  nand ginst18640 (P3_R1054_U82, P3_R1054_U257, P3_R1054_U258);
  nand ginst18641 (P3_R1054_U83, P3_R1054_U262, P3_R1054_U263);
  nand ginst18642 (P3_R1054_U84, P3_R1054_U278, P3_R1054_U279);
  nand ginst18643 (P3_R1054_U85, P3_R1054_U283, P3_R1054_U284);
  nand ginst18644 (P3_R1054_U86, P3_R1054_U129, P3_R1054_U131, P3_R1054_U132);
  nand ginst18645 (P3_R1054_U87, P3_R1054_U113, P3_R1054_U115, P3_R1054_U116);
  not ginst18646 (P3_R1054_U88, P3_U3391);
  not ginst18647 (P3_R1054_U89, P3_U3379);
  and ginst18648 (P3_R1054_U9, P3_R1054_U158, P3_R1054_U159);
  not ginst18649 (P3_R1054_U90, P3_U3563);
  nand ginst18650 (P3_R1054_U91, P3_R1054_U189, P3_R1054_U190);
  not ginst18651 (P3_R1054_U92, P3_U3442);
  nand ginst18652 (P3_R1054_U93, P3_R1054_U181, P3_R1054_U182);
  nand ginst18653 (P3_R1054_U94, P3_R1054_U171, P3_R1054_U172);
  nand ginst18654 (P3_R1054_U95, P3_R1054_U167, P3_R1054_U168);
  nand ginst18655 (P3_R1054_U96, P3_R1054_U163, P3_R1054_U164);
  not ginst18656 (P3_R1054_U97, P3_R1054_U25);
  not ginst18657 (P3_R1054_U98, P3_R1054_U36);
  nand ginst18658 (P3_R1054_U99, P3_R1054_U46, P3_U3418);
  and ginst18659 (P3_R1077_U10, P3_R1077_U348, P3_R1077_U351);
  nand ginst18660 (P3_R1077_U100, P3_R1077_U398, P3_R1077_U399);
  nand ginst18661 (P3_R1077_U101, P3_R1077_U407, P3_R1077_U408);
  nand ginst18662 (P3_R1077_U102, P3_R1077_U414, P3_R1077_U415);
  nand ginst18663 (P3_R1077_U103, P3_R1077_U421, P3_R1077_U422);
  nand ginst18664 (P3_R1077_U104, P3_R1077_U428, P3_R1077_U429);
  nand ginst18665 (P3_R1077_U105, P3_R1077_U433, P3_R1077_U434);
  nand ginst18666 (P3_R1077_U106, P3_R1077_U440, P3_R1077_U441);
  nand ginst18667 (P3_R1077_U107, P3_R1077_U447, P3_R1077_U448);
  nand ginst18668 (P3_R1077_U108, P3_R1077_U461, P3_R1077_U462);
  nand ginst18669 (P3_R1077_U109, P3_R1077_U466, P3_R1077_U467);
  and ginst18670 (P3_R1077_U11, P3_R1077_U341, P3_R1077_U344);
  nand ginst18671 (P3_R1077_U110, P3_R1077_U473, P3_R1077_U474);
  nand ginst18672 (P3_R1077_U111, P3_R1077_U480, P3_R1077_U481);
  nand ginst18673 (P3_R1077_U112, P3_R1077_U487, P3_R1077_U488);
  nand ginst18674 (P3_R1077_U113, P3_R1077_U494, P3_R1077_U495);
  nand ginst18675 (P3_R1077_U114, P3_R1077_U499, P3_R1077_U500);
  and ginst18676 (P3_R1077_U115, P3_R1077_U187, P3_R1077_U189);
  and ginst18677 (P3_R1077_U116, P3_R1077_U180, P3_R1077_U4);
  and ginst18678 (P3_R1077_U117, P3_R1077_U192, P3_R1077_U194);
  and ginst18679 (P3_R1077_U118, P3_R1077_U200, P3_R1077_U201);
  and ginst18680 (P3_R1077_U119, P3_R1077_U22, P3_R1077_U381, P3_R1077_U382);
  and ginst18681 (P3_R1077_U12, P3_R1077_U332, P3_R1077_U335);
  and ginst18682 (P3_R1077_U120, P3_R1077_U212, P3_R1077_U5);
  and ginst18683 (P3_R1077_U121, P3_R1077_U180, P3_R1077_U181);
  and ginst18684 (P3_R1077_U122, P3_R1077_U218, P3_R1077_U220);
  and ginst18685 (P3_R1077_U123, P3_R1077_U34, P3_R1077_U388, P3_R1077_U389);
  and ginst18686 (P3_R1077_U124, P3_R1077_U226, P3_R1077_U4);
  and ginst18687 (P3_R1077_U125, P3_R1077_U181, P3_R1077_U234);
  and ginst18688 (P3_R1077_U126, P3_R1077_U204, P3_R1077_U6);
  and ginst18689 (P3_R1077_U127, P3_R1077_U171, P3_R1077_U239);
  and ginst18690 (P3_R1077_U128, P3_R1077_U250, P3_R1077_U7);
  and ginst18691 (P3_R1077_U129, P3_R1077_U172, P3_R1077_U248);
  and ginst18692 (P3_R1077_U13, P3_R1077_U323, P3_R1077_U326);
  and ginst18693 (P3_R1077_U130, P3_R1077_U267, P3_R1077_U268);
  and ginst18694 (P3_R1077_U131, P3_R1077_U273, P3_R1077_U282, P3_R1077_U9);
  and ginst18695 (P3_R1077_U132, P3_R1077_U280, P3_R1077_U285);
  and ginst18696 (P3_R1077_U133, P3_R1077_U298, P3_R1077_U301);
  and ginst18697 (P3_R1077_U134, P3_R1077_U302, P3_R1077_U368);
  and ginst18698 (P3_R1077_U135, P3_R1077_U160, P3_R1077_U278);
  and ginst18699 (P3_R1077_U136, P3_R1077_U454, P3_R1077_U455, P3_R1077_U80);
  and ginst18700 (P3_R1077_U137, P3_R1077_U325, P3_R1077_U9);
  and ginst18701 (P3_R1077_U138, P3_R1077_U468, P3_R1077_U469, P3_R1077_U59);
  and ginst18702 (P3_R1077_U139, P3_R1077_U334, P3_R1077_U8);
  and ginst18703 (P3_R1077_U14, P3_R1077_U318, P3_R1077_U320);
  and ginst18704 (P3_R1077_U140, P3_R1077_U172, P3_R1077_U489, P3_R1077_U490);
  and ginst18705 (P3_R1077_U141, P3_R1077_U343, P3_R1077_U7);
  and ginst18706 (P3_R1077_U142, P3_R1077_U171, P3_R1077_U501, P3_R1077_U502);
  and ginst18707 (P3_R1077_U143, P3_R1077_U350, P3_R1077_U6);
  nand ginst18708 (P3_R1077_U144, P3_R1077_U118, P3_R1077_U202);
  nand ginst18709 (P3_R1077_U145, P3_R1077_U217, P3_R1077_U229);
  not ginst18710 (P3_R1077_U146, P3_U3054);
  not ginst18711 (P3_R1077_U147, P3_U3908);
  and ginst18712 (P3_R1077_U148, P3_R1077_U402, P3_R1077_U403);
  nand ginst18713 (P3_R1077_U149, P3_R1077_U169, P3_R1077_U304, P3_R1077_U364);
  and ginst18714 (P3_R1077_U15, P3_R1077_U310, P3_R1077_U313);
  and ginst18715 (P3_R1077_U150, P3_R1077_U409, P3_R1077_U410);
  nand ginst18716 (P3_R1077_U151, P3_R1077_U134, P3_R1077_U369, P3_R1077_U370);
  and ginst18717 (P3_R1077_U152, P3_R1077_U416, P3_R1077_U417);
  nand ginst18718 (P3_R1077_U153, P3_R1077_U299, P3_R1077_U365, P3_R1077_U86);
  and ginst18719 (P3_R1077_U154, P3_R1077_U423, P3_R1077_U424);
  nand ginst18720 (P3_R1077_U155, P3_R1077_U292, P3_R1077_U293);
  and ginst18721 (P3_R1077_U156, P3_R1077_U435, P3_R1077_U436);
  nand ginst18722 (P3_R1077_U157, P3_R1077_U288, P3_R1077_U289);
  and ginst18723 (P3_R1077_U158, P3_R1077_U442, P3_R1077_U443);
  nand ginst18724 (P3_R1077_U159, P3_R1077_U132, P3_R1077_U284);
  and ginst18725 (P3_R1077_U16, P3_R1077_U232, P3_R1077_U235);
  and ginst18726 (P3_R1077_U160, P3_R1077_U449, P3_R1077_U450);
  nand ginst18727 (P3_R1077_U161, P3_R1077_U327, P3_R1077_U43);
  nand ginst18728 (P3_R1077_U162, P3_R1077_U130, P3_R1077_U269);
  and ginst18729 (P3_R1077_U163, P3_R1077_U475, P3_R1077_U476);
  nand ginst18730 (P3_R1077_U164, P3_R1077_U256, P3_R1077_U257);
  and ginst18731 (P3_R1077_U165, P3_R1077_U482, P3_R1077_U483);
  nand ginst18732 (P3_R1077_U166, P3_R1077_U252, P3_R1077_U253);
  nand ginst18733 (P3_R1077_U167, P3_R1077_U242, P3_R1077_U243);
  nand ginst18734 (P3_R1077_U168, P3_R1077_U366, P3_R1077_U367);
  nand ginst18735 (P3_R1077_U169, P3_R1077_U151, P3_U3053);
  and ginst18736 (P3_R1077_U17, P3_R1077_U224, P3_R1077_U227);
  not ginst18737 (P3_R1077_U170, P3_R1077_U34);
  nand ginst18738 (P3_R1077_U171, P3_U3082, P3_U3416);
  nand ginst18739 (P3_R1077_U172, P3_U3071, P3_U3425);
  nand ginst18740 (P3_R1077_U173, P3_U3057, P3_U3902);
  not ginst18741 (P3_R1077_U174, P3_R1077_U68);
  not ginst18742 (P3_R1077_U175, P3_R1077_U77);
  nand ginst18743 (P3_R1077_U176, P3_U3064, P3_U3903);
  not ginst18744 (P3_R1077_U177, P3_R1077_U61);
  or ginst18745 (P3_R1077_U178, P3_U3066, P3_U3404);
  or ginst18746 (P3_R1077_U179, P3_U3059, P3_U3401);
  and ginst18747 (P3_R1077_U18, P3_R1077_U210, P3_R1077_U213);
  or ginst18748 (P3_R1077_U180, P3_U3063, P3_U3398);
  or ginst18749 (P3_R1077_U181, P3_U3067, P3_U3395);
  not ginst18750 (P3_R1077_U182, P3_R1077_U31);
  or ginst18751 (P3_R1077_U183, P3_U3077, P3_U3392);
  not ginst18752 (P3_R1077_U184, P3_R1077_U42);
  not ginst18753 (P3_R1077_U185, P3_R1077_U43);
  nand ginst18754 (P3_R1077_U186, P3_R1077_U42, P3_R1077_U43);
  nand ginst18755 (P3_R1077_U187, P3_U3067, P3_U3395);
  nand ginst18756 (P3_R1077_U188, P3_R1077_U181, P3_R1077_U186);
  nand ginst18757 (P3_R1077_U189, P3_U3063, P3_U3398);
  not ginst18758 (P3_R1077_U19, P3_U3407);
  nand ginst18759 (P3_R1077_U190, P3_R1077_U115, P3_R1077_U188);
  nand ginst18760 (P3_R1077_U191, P3_R1077_U34, P3_R1077_U35);
  nand ginst18761 (P3_R1077_U192, P3_R1077_U191, P3_U3066);
  nand ginst18762 (P3_R1077_U193, P3_R1077_U116, P3_R1077_U190);
  nand ginst18763 (P3_R1077_U194, P3_R1077_U170, P3_U3404);
  not ginst18764 (P3_R1077_U195, P3_R1077_U41);
  or ginst18765 (P3_R1077_U196, P3_U3069, P3_U3410);
  or ginst18766 (P3_R1077_U197, P3_U3070, P3_U3407);
  not ginst18767 (P3_R1077_U198, P3_R1077_U22);
  nand ginst18768 (P3_R1077_U199, P3_R1077_U22, P3_R1077_U23);
  not ginst18769 (P3_R1077_U20, P3_U3070);
  nand ginst18770 (P3_R1077_U200, P3_R1077_U199, P3_U3069);
  nand ginst18771 (P3_R1077_U201, P3_R1077_U198, P3_U3410);
  nand ginst18772 (P3_R1077_U202, P3_R1077_U41, P3_R1077_U5);
  not ginst18773 (P3_R1077_U203, P3_R1077_U144);
  or ginst18774 (P3_R1077_U204, P3_U3083, P3_U3413);
  nand ginst18775 (P3_R1077_U205, P3_R1077_U144, P3_R1077_U204);
  not ginst18776 (P3_R1077_U206, P3_R1077_U40);
  or ginst18777 (P3_R1077_U207, P3_U3082, P3_U3416);
  or ginst18778 (P3_R1077_U208, P3_U3070, P3_U3407);
  nand ginst18779 (P3_R1077_U209, P3_R1077_U208, P3_R1077_U41);
  not ginst18780 (P3_R1077_U21, P3_U3069);
  nand ginst18781 (P3_R1077_U210, P3_R1077_U119, P3_R1077_U209);
  nand ginst18782 (P3_R1077_U211, P3_R1077_U195, P3_R1077_U22);
  nand ginst18783 (P3_R1077_U212, P3_U3069, P3_U3410);
  nand ginst18784 (P3_R1077_U213, P3_R1077_U120, P3_R1077_U211);
  or ginst18785 (P3_R1077_U214, P3_U3070, P3_U3407);
  nand ginst18786 (P3_R1077_U215, P3_R1077_U181, P3_R1077_U185);
  nand ginst18787 (P3_R1077_U216, P3_U3067, P3_U3395);
  not ginst18788 (P3_R1077_U217, P3_R1077_U45);
  nand ginst18789 (P3_R1077_U218, P3_R1077_U121, P3_R1077_U184);
  nand ginst18790 (P3_R1077_U219, P3_R1077_U180, P3_R1077_U45);
  nand ginst18791 (P3_R1077_U22, P3_U3070, P3_U3407);
  nand ginst18792 (P3_R1077_U220, P3_U3063, P3_U3398);
  not ginst18793 (P3_R1077_U221, P3_R1077_U44);
  or ginst18794 (P3_R1077_U222, P3_U3059, P3_U3401);
  nand ginst18795 (P3_R1077_U223, P3_R1077_U222, P3_R1077_U44);
  nand ginst18796 (P3_R1077_U224, P3_R1077_U123, P3_R1077_U223);
  nand ginst18797 (P3_R1077_U225, P3_R1077_U221, P3_R1077_U34);
  nand ginst18798 (P3_R1077_U226, P3_U3066, P3_U3404);
  nand ginst18799 (P3_R1077_U227, P3_R1077_U124, P3_R1077_U225);
  or ginst18800 (P3_R1077_U228, P3_U3059, P3_U3401);
  nand ginst18801 (P3_R1077_U229, P3_R1077_U181, P3_R1077_U184);
  not ginst18802 (P3_R1077_U23, P3_U3410);
  not ginst18803 (P3_R1077_U230, P3_R1077_U145);
  nand ginst18804 (P3_R1077_U231, P3_U3063, P3_U3398);
  nand ginst18805 (P3_R1077_U232, P3_R1077_U400, P3_R1077_U401, P3_R1077_U42, P3_R1077_U43);
  nand ginst18806 (P3_R1077_U233, P3_R1077_U42, P3_R1077_U43);
  nand ginst18807 (P3_R1077_U234, P3_U3067, P3_U3395);
  nand ginst18808 (P3_R1077_U235, P3_R1077_U125, P3_R1077_U233);
  or ginst18809 (P3_R1077_U236, P3_U3082, P3_U3416);
  or ginst18810 (P3_R1077_U237, P3_U3061, P3_U3419);
  nand ginst18811 (P3_R1077_U238, P3_R1077_U177, P3_R1077_U6);
  nand ginst18812 (P3_R1077_U239, P3_U3061, P3_U3419);
  not ginst18813 (P3_R1077_U24, P3_U3401);
  nand ginst18814 (P3_R1077_U240, P3_R1077_U127, P3_R1077_U238);
  or ginst18815 (P3_R1077_U241, P3_U3061, P3_U3419);
  nand ginst18816 (P3_R1077_U242, P3_R1077_U126, P3_R1077_U144);
  nand ginst18817 (P3_R1077_U243, P3_R1077_U240, P3_R1077_U241);
  not ginst18818 (P3_R1077_U244, P3_R1077_U167);
  or ginst18819 (P3_R1077_U245, P3_U3079, P3_U3428);
  or ginst18820 (P3_R1077_U246, P3_U3071, P3_U3425);
  nand ginst18821 (P3_R1077_U247, P3_R1077_U174, P3_R1077_U7);
  nand ginst18822 (P3_R1077_U248, P3_U3079, P3_U3428);
  nand ginst18823 (P3_R1077_U249, P3_R1077_U129, P3_R1077_U247);
  not ginst18824 (P3_R1077_U25, P3_U3059);
  or ginst18825 (P3_R1077_U250, P3_U3062, P3_U3422);
  or ginst18826 (P3_R1077_U251, P3_U3079, P3_U3428);
  nand ginst18827 (P3_R1077_U252, P3_R1077_U128, P3_R1077_U167);
  nand ginst18828 (P3_R1077_U253, P3_R1077_U249, P3_R1077_U251);
  not ginst18829 (P3_R1077_U254, P3_R1077_U166);
  or ginst18830 (P3_R1077_U255, P3_U3078, P3_U3431);
  nand ginst18831 (P3_R1077_U256, P3_R1077_U166, P3_R1077_U255);
  nand ginst18832 (P3_R1077_U257, P3_U3078, P3_U3431);
  not ginst18833 (P3_R1077_U258, P3_R1077_U164);
  or ginst18834 (P3_R1077_U259, P3_U3073, P3_U3434);
  not ginst18835 (P3_R1077_U26, P3_U3066);
  nand ginst18836 (P3_R1077_U260, P3_R1077_U164, P3_R1077_U259);
  nand ginst18837 (P3_R1077_U261, P3_U3073, P3_U3434);
  not ginst18838 (P3_R1077_U262, P3_R1077_U92);
  or ginst18839 (P3_R1077_U263, P3_U3068, P3_U3440);
  or ginst18840 (P3_R1077_U264, P3_U3072, P3_U3437);
  not ginst18841 (P3_R1077_U265, P3_R1077_U59);
  nand ginst18842 (P3_R1077_U266, P3_R1077_U59, P3_R1077_U60);
  nand ginst18843 (P3_R1077_U267, P3_R1077_U266, P3_U3068);
  nand ginst18844 (P3_R1077_U268, P3_R1077_U265, P3_U3440);
  nand ginst18845 (P3_R1077_U269, P3_R1077_U8, P3_R1077_U92);
  not ginst18846 (P3_R1077_U27, P3_U3395);
  not ginst18847 (P3_R1077_U270, P3_R1077_U162);
  or ginst18848 (P3_R1077_U271, P3_U3075, P3_U3907);
  or ginst18849 (P3_R1077_U272, P3_U3080, P3_U3445);
  or ginst18850 (P3_R1077_U273, P3_U3074, P3_U3906);
  not ginst18851 (P3_R1077_U274, P3_R1077_U80);
  nand ginst18852 (P3_R1077_U275, P3_R1077_U274, P3_U3907);
  nand ginst18853 (P3_R1077_U276, P3_R1077_U275, P3_R1077_U90);
  nand ginst18854 (P3_R1077_U277, P3_R1077_U80, P3_R1077_U81);
  nand ginst18855 (P3_R1077_U278, P3_R1077_U276, P3_R1077_U277);
  nand ginst18856 (P3_R1077_U279, P3_R1077_U175, P3_R1077_U9);
  not ginst18857 (P3_R1077_U28, P3_U3067);
  nand ginst18858 (P3_R1077_U280, P3_U3074, P3_U3906);
  nand ginst18859 (P3_R1077_U281, P3_R1077_U278, P3_R1077_U279);
  or ginst18860 (P3_R1077_U282, P3_U3081, P3_U3443);
  or ginst18861 (P3_R1077_U283, P3_U3074, P3_U3906);
  nand ginst18862 (P3_R1077_U284, P3_R1077_U131, P3_R1077_U162);
  nand ginst18863 (P3_R1077_U285, P3_R1077_U281, P3_R1077_U283);
  not ginst18864 (P3_R1077_U286, P3_R1077_U159);
  or ginst18865 (P3_R1077_U287, P3_U3060, P3_U3905);
  nand ginst18866 (P3_R1077_U288, P3_R1077_U159, P3_R1077_U287);
  nand ginst18867 (P3_R1077_U289, P3_U3060, P3_U3905);
  not ginst18868 (P3_R1077_U29, P3_U3387);
  not ginst18869 (P3_R1077_U290, P3_R1077_U157);
  or ginst18870 (P3_R1077_U291, P3_U3065, P3_U3904);
  nand ginst18871 (P3_R1077_U292, P3_R1077_U157, P3_R1077_U291);
  nand ginst18872 (P3_R1077_U293, P3_U3065, P3_U3904);
  not ginst18873 (P3_R1077_U294, P3_R1077_U155);
  or ginst18874 (P3_R1077_U295, P3_U3057, P3_U3902);
  nand ginst18875 (P3_R1077_U296, P3_R1077_U173, P3_R1077_U176);
  not ginst18876 (P3_R1077_U297, P3_R1077_U86);
  or ginst18877 (P3_R1077_U298, P3_U3064, P3_U3903);
  nand ginst18878 (P3_R1077_U299, P3_R1077_U155, P3_R1077_U168, P3_R1077_U298);
  not ginst18879 (P3_R1077_U30, P3_U3076);
  not ginst18880 (P3_R1077_U300, P3_R1077_U153);
  or ginst18881 (P3_R1077_U301, P3_U3052, P3_U3900);
  nand ginst18882 (P3_R1077_U302, P3_U3052, P3_U3900);
  not ginst18883 (P3_R1077_U303, P3_R1077_U151);
  nand ginst18884 (P3_R1077_U304, P3_R1077_U151, P3_U3899);
  not ginst18885 (P3_R1077_U305, P3_R1077_U149);
  nand ginst18886 (P3_R1077_U306, P3_R1077_U155, P3_R1077_U298);
  not ginst18887 (P3_R1077_U307, P3_R1077_U89);
  or ginst18888 (P3_R1077_U308, P3_U3057, P3_U3902);
  nand ginst18889 (P3_R1077_U309, P3_R1077_U308, P3_R1077_U89);
  nand ginst18890 (P3_R1077_U31, P3_U3076, P3_U3387);
  nand ginst18891 (P3_R1077_U310, P3_R1077_U154, P3_R1077_U173, P3_R1077_U309);
  nand ginst18892 (P3_R1077_U311, P3_R1077_U173, P3_R1077_U307);
  nand ginst18893 (P3_R1077_U312, P3_U3056, P3_U3901);
  nand ginst18894 (P3_R1077_U313, P3_R1077_U168, P3_R1077_U311, P3_R1077_U312);
  or ginst18895 (P3_R1077_U314, P3_U3057, P3_U3902);
  nand ginst18896 (P3_R1077_U315, P3_R1077_U162, P3_R1077_U282);
  not ginst18897 (P3_R1077_U316, P3_R1077_U91);
  nand ginst18898 (P3_R1077_U317, P3_R1077_U9, P3_R1077_U91);
  nand ginst18899 (P3_R1077_U318, P3_R1077_U135, P3_R1077_U317);
  nand ginst18900 (P3_R1077_U319, P3_R1077_U278, P3_R1077_U317);
  not ginst18901 (P3_R1077_U32, P3_U3398);
  nand ginst18902 (P3_R1077_U320, P3_R1077_U319, P3_R1077_U453);
  or ginst18903 (P3_R1077_U321, P3_U3080, P3_U3445);
  nand ginst18904 (P3_R1077_U322, P3_R1077_U321, P3_R1077_U91);
  nand ginst18905 (P3_R1077_U323, P3_R1077_U136, P3_R1077_U322);
  nand ginst18906 (P3_R1077_U324, P3_R1077_U316, P3_R1077_U80);
  nand ginst18907 (P3_R1077_U325, P3_U3075, P3_U3907);
  nand ginst18908 (P3_R1077_U326, P3_R1077_U137, P3_R1077_U324);
  or ginst18909 (P3_R1077_U327, P3_U3077, P3_U3392);
  not ginst18910 (P3_R1077_U328, P3_R1077_U161);
  or ginst18911 (P3_R1077_U329, P3_U3080, P3_U3445);
  not ginst18912 (P3_R1077_U33, P3_U3063);
  or ginst18913 (P3_R1077_U330, P3_U3072, P3_U3437);
  nand ginst18914 (P3_R1077_U331, P3_R1077_U330, P3_R1077_U92);
  nand ginst18915 (P3_R1077_U332, P3_R1077_U138, P3_R1077_U331);
  nand ginst18916 (P3_R1077_U333, P3_R1077_U262, P3_R1077_U59);
  nand ginst18917 (P3_R1077_U334, P3_U3068, P3_U3440);
  nand ginst18918 (P3_R1077_U335, P3_R1077_U139, P3_R1077_U333);
  or ginst18919 (P3_R1077_U336, P3_U3072, P3_U3437);
  nand ginst18920 (P3_R1077_U337, P3_R1077_U167, P3_R1077_U250);
  not ginst18921 (P3_R1077_U338, P3_R1077_U93);
  or ginst18922 (P3_R1077_U339, P3_U3071, P3_U3425);
  nand ginst18923 (P3_R1077_U34, P3_U3059, P3_U3401);
  nand ginst18924 (P3_R1077_U340, P3_R1077_U339, P3_R1077_U93);
  nand ginst18925 (P3_R1077_U341, P3_R1077_U140, P3_R1077_U340);
  nand ginst18926 (P3_R1077_U342, P3_R1077_U172, P3_R1077_U338);
  nand ginst18927 (P3_R1077_U343, P3_U3079, P3_U3428);
  nand ginst18928 (P3_R1077_U344, P3_R1077_U141, P3_R1077_U342);
  or ginst18929 (P3_R1077_U345, P3_U3071, P3_U3425);
  or ginst18930 (P3_R1077_U346, P3_U3082, P3_U3416);
  nand ginst18931 (P3_R1077_U347, P3_R1077_U346, P3_R1077_U40);
  nand ginst18932 (P3_R1077_U348, P3_R1077_U142, P3_R1077_U347);
  nand ginst18933 (P3_R1077_U349, P3_R1077_U171, P3_R1077_U206);
  not ginst18934 (P3_R1077_U35, P3_U3404);
  nand ginst18935 (P3_R1077_U350, P3_U3061, P3_U3419);
  nand ginst18936 (P3_R1077_U351, P3_R1077_U143, P3_R1077_U349);
  nand ginst18937 (P3_R1077_U352, P3_R1077_U171, P3_R1077_U207);
  nand ginst18938 (P3_R1077_U353, P3_R1077_U204, P3_R1077_U61);
  nand ginst18939 (P3_R1077_U354, P3_R1077_U214, P3_R1077_U22);
  nand ginst18940 (P3_R1077_U355, P3_R1077_U228, P3_R1077_U34);
  nand ginst18941 (P3_R1077_U356, P3_R1077_U180, P3_R1077_U231);
  nand ginst18942 (P3_R1077_U357, P3_R1077_U173, P3_R1077_U314);
  nand ginst18943 (P3_R1077_U358, P3_R1077_U176, P3_R1077_U298);
  nand ginst18944 (P3_R1077_U359, P3_R1077_U329, P3_R1077_U80);
  not ginst18945 (P3_R1077_U36, P3_U3413);
  nand ginst18946 (P3_R1077_U360, P3_R1077_U282, P3_R1077_U77);
  nand ginst18947 (P3_R1077_U361, P3_R1077_U336, P3_R1077_U59);
  nand ginst18948 (P3_R1077_U362, P3_R1077_U172, P3_R1077_U345);
  nand ginst18949 (P3_R1077_U363, P3_R1077_U250, P3_R1077_U68);
  nand ginst18950 (P3_R1077_U364, P3_U3053, P3_U3899);
  nand ginst18951 (P3_R1077_U365, P3_R1077_U168, P3_R1077_U296);
  nand ginst18952 (P3_R1077_U366, P3_R1077_U295, P3_U3056);
  nand ginst18953 (P3_R1077_U367, P3_R1077_U295, P3_U3901);
  nand ginst18954 (P3_R1077_U368, P3_R1077_U168, P3_R1077_U296, P3_R1077_U301);
  nand ginst18955 (P3_R1077_U369, P3_R1077_U133, P3_R1077_U155, P3_R1077_U168);
  not ginst18956 (P3_R1077_U37, P3_U3083);
  nand ginst18957 (P3_R1077_U370, P3_R1077_U297, P3_R1077_U301);
  nand ginst18958 (P3_R1077_U371, P3_R1077_U39, P3_U3082);
  nand ginst18959 (P3_R1077_U372, P3_R1077_U38, P3_U3416);
  nand ginst18960 (P3_R1077_U373, P3_R1077_U371, P3_R1077_U372);
  nand ginst18961 (P3_R1077_U374, P3_R1077_U352, P3_R1077_U40);
  nand ginst18962 (P3_R1077_U375, P3_R1077_U206, P3_R1077_U373);
  nand ginst18963 (P3_R1077_U376, P3_R1077_U36, P3_U3083);
  nand ginst18964 (P3_R1077_U377, P3_R1077_U37, P3_U3413);
  nand ginst18965 (P3_R1077_U378, P3_R1077_U376, P3_R1077_U377);
  nand ginst18966 (P3_R1077_U379, P3_R1077_U144, P3_R1077_U353);
  not ginst18967 (P3_R1077_U38, P3_U3082);
  nand ginst18968 (P3_R1077_U380, P3_R1077_U203, P3_R1077_U378);
  nand ginst18969 (P3_R1077_U381, P3_R1077_U23, P3_U3069);
  nand ginst18970 (P3_R1077_U382, P3_R1077_U21, P3_U3410);
  nand ginst18971 (P3_R1077_U383, P3_R1077_U19, P3_U3070);
  nand ginst18972 (P3_R1077_U384, P3_R1077_U20, P3_U3407);
  nand ginst18973 (P3_R1077_U385, P3_R1077_U383, P3_R1077_U384);
  nand ginst18974 (P3_R1077_U386, P3_R1077_U354, P3_R1077_U41);
  nand ginst18975 (P3_R1077_U387, P3_R1077_U195, P3_R1077_U385);
  nand ginst18976 (P3_R1077_U388, P3_R1077_U35, P3_U3066);
  nand ginst18977 (P3_R1077_U389, P3_R1077_U26, P3_U3404);
  not ginst18978 (P3_R1077_U39, P3_U3416);
  nand ginst18979 (P3_R1077_U390, P3_R1077_U24, P3_U3059);
  nand ginst18980 (P3_R1077_U391, P3_R1077_U25, P3_U3401);
  nand ginst18981 (P3_R1077_U392, P3_R1077_U390, P3_R1077_U391);
  nand ginst18982 (P3_R1077_U393, P3_R1077_U355, P3_R1077_U44);
  nand ginst18983 (P3_R1077_U394, P3_R1077_U221, P3_R1077_U392);
  nand ginst18984 (P3_R1077_U395, P3_R1077_U32, P3_U3063);
  nand ginst18985 (P3_R1077_U396, P3_R1077_U33, P3_U3398);
  nand ginst18986 (P3_R1077_U397, P3_R1077_U395, P3_R1077_U396);
  nand ginst18987 (P3_R1077_U398, P3_R1077_U145, P3_R1077_U356);
  nand ginst18988 (P3_R1077_U399, P3_R1077_U230, P3_R1077_U397);
  and ginst18989 (P3_R1077_U4, P3_R1077_U178, P3_R1077_U179);
  nand ginst18990 (P3_R1077_U40, P3_R1077_U205, P3_R1077_U61);
  nand ginst18991 (P3_R1077_U400, P3_R1077_U27, P3_U3067);
  nand ginst18992 (P3_R1077_U401, P3_R1077_U28, P3_U3395);
  nand ginst18993 (P3_R1077_U402, P3_R1077_U147, P3_U3054);
  nand ginst18994 (P3_R1077_U403, P3_R1077_U146, P3_U3908);
  nand ginst18995 (P3_R1077_U404, P3_R1077_U147, P3_U3054);
  nand ginst18996 (P3_R1077_U405, P3_R1077_U146, P3_U3908);
  nand ginst18997 (P3_R1077_U406, P3_R1077_U404, P3_R1077_U405);
  nand ginst18998 (P3_R1077_U407, P3_R1077_U148, P3_R1077_U149);
  nand ginst18999 (P3_R1077_U408, P3_R1077_U305, P3_R1077_U406);
  nand ginst19000 (P3_R1077_U409, P3_R1077_U88, P3_U3053);
  nand ginst19001 (P3_R1077_U41, P3_R1077_U117, P3_R1077_U193);
  nand ginst19002 (P3_R1077_U410, P3_R1077_U87, P3_U3899);
  nand ginst19003 (P3_R1077_U411, P3_R1077_U88, P3_U3053);
  nand ginst19004 (P3_R1077_U412, P3_R1077_U87, P3_U3899);
  nand ginst19005 (P3_R1077_U413, P3_R1077_U411, P3_R1077_U412);
  nand ginst19006 (P3_R1077_U414, P3_R1077_U150, P3_R1077_U151);
  nand ginst19007 (P3_R1077_U415, P3_R1077_U303, P3_R1077_U413);
  nand ginst19008 (P3_R1077_U416, P3_R1077_U46, P3_U3052);
  nand ginst19009 (P3_R1077_U417, P3_R1077_U47, P3_U3900);
  nand ginst19010 (P3_R1077_U418, P3_R1077_U46, P3_U3052);
  nand ginst19011 (P3_R1077_U419, P3_R1077_U47, P3_U3900);
  nand ginst19012 (P3_R1077_U42, P3_R1077_U182, P3_R1077_U183);
  nand ginst19013 (P3_R1077_U420, P3_R1077_U418, P3_R1077_U419);
  nand ginst19014 (P3_R1077_U421, P3_R1077_U152, P3_R1077_U153);
  nand ginst19015 (P3_R1077_U422, P3_R1077_U300, P3_R1077_U420);
  nand ginst19016 (P3_R1077_U423, P3_R1077_U49, P3_U3056);
  nand ginst19017 (P3_R1077_U424, P3_R1077_U48, P3_U3901);
  nand ginst19018 (P3_R1077_U425, P3_R1077_U50, P3_U3057);
  nand ginst19019 (P3_R1077_U426, P3_R1077_U51, P3_U3902);
  nand ginst19020 (P3_R1077_U427, P3_R1077_U425, P3_R1077_U426);
  nand ginst19021 (P3_R1077_U428, P3_R1077_U357, P3_R1077_U89);
  nand ginst19022 (P3_R1077_U429, P3_R1077_U307, P3_R1077_U427);
  nand ginst19023 (P3_R1077_U43, P3_U3077, P3_U3392);
  nand ginst19024 (P3_R1077_U430, P3_R1077_U52, P3_U3064);
  nand ginst19025 (P3_R1077_U431, P3_R1077_U53, P3_U3903);
  nand ginst19026 (P3_R1077_U432, P3_R1077_U430, P3_R1077_U431);
  nand ginst19027 (P3_R1077_U433, P3_R1077_U155, P3_R1077_U358);
  nand ginst19028 (P3_R1077_U434, P3_R1077_U294, P3_R1077_U432);
  nand ginst19029 (P3_R1077_U435, P3_R1077_U84, P3_U3065);
  nand ginst19030 (P3_R1077_U436, P3_R1077_U85, P3_U3904);
  nand ginst19031 (P3_R1077_U437, P3_R1077_U84, P3_U3065);
  nand ginst19032 (P3_R1077_U438, P3_R1077_U85, P3_U3904);
  nand ginst19033 (P3_R1077_U439, P3_R1077_U437, P3_R1077_U438);
  nand ginst19034 (P3_R1077_U44, P3_R1077_U122, P3_R1077_U219);
  nand ginst19035 (P3_R1077_U440, P3_R1077_U156, P3_R1077_U157);
  nand ginst19036 (P3_R1077_U441, P3_R1077_U290, P3_R1077_U439);
  nand ginst19037 (P3_R1077_U442, P3_R1077_U82, P3_U3060);
  nand ginst19038 (P3_R1077_U443, P3_R1077_U83, P3_U3905);
  nand ginst19039 (P3_R1077_U444, P3_R1077_U82, P3_U3060);
  nand ginst19040 (P3_R1077_U445, P3_R1077_U83, P3_U3905);
  nand ginst19041 (P3_R1077_U446, P3_R1077_U444, P3_R1077_U445);
  nand ginst19042 (P3_R1077_U447, P3_R1077_U158, P3_R1077_U159);
  nand ginst19043 (P3_R1077_U448, P3_R1077_U286, P3_R1077_U446);
  nand ginst19044 (P3_R1077_U449, P3_R1077_U54, P3_U3074);
  nand ginst19045 (P3_R1077_U45, P3_R1077_U215, P3_R1077_U216);
  nand ginst19046 (P3_R1077_U450, P3_R1077_U55, P3_U3906);
  nand ginst19047 (P3_R1077_U451, P3_R1077_U54, P3_U3074);
  nand ginst19048 (P3_R1077_U452, P3_R1077_U55, P3_U3906);
  nand ginst19049 (P3_R1077_U453, P3_R1077_U451, P3_R1077_U452);
  nand ginst19050 (P3_R1077_U454, P3_R1077_U81, P3_U3075);
  nand ginst19051 (P3_R1077_U455, P3_R1077_U90, P3_U3907);
  nand ginst19052 (P3_R1077_U456, P3_R1077_U161, P3_R1077_U182);
  nand ginst19053 (P3_R1077_U457, P3_R1077_U31, P3_R1077_U328);
  nand ginst19054 (P3_R1077_U458, P3_R1077_U78, P3_U3080);
  nand ginst19055 (P3_R1077_U459, P3_R1077_U79, P3_U3445);
  not ginst19056 (P3_R1077_U46, P3_U3900);
  nand ginst19057 (P3_R1077_U460, P3_R1077_U458, P3_R1077_U459);
  nand ginst19058 (P3_R1077_U461, P3_R1077_U359, P3_R1077_U91);
  nand ginst19059 (P3_R1077_U462, P3_R1077_U316, P3_R1077_U460);
  nand ginst19060 (P3_R1077_U463, P3_R1077_U75, P3_U3081);
  nand ginst19061 (P3_R1077_U464, P3_R1077_U76, P3_U3443);
  nand ginst19062 (P3_R1077_U465, P3_R1077_U463, P3_R1077_U464);
  nand ginst19063 (P3_R1077_U466, P3_R1077_U162, P3_R1077_U360);
  nand ginst19064 (P3_R1077_U467, P3_R1077_U270, P3_R1077_U465);
  nand ginst19065 (P3_R1077_U468, P3_R1077_U60, P3_U3068);
  nand ginst19066 (P3_R1077_U469, P3_R1077_U58, P3_U3440);
  not ginst19067 (P3_R1077_U47, P3_U3052);
  nand ginst19068 (P3_R1077_U470, P3_R1077_U56, P3_U3072);
  nand ginst19069 (P3_R1077_U471, P3_R1077_U57, P3_U3437);
  nand ginst19070 (P3_R1077_U472, P3_R1077_U470, P3_R1077_U471);
  nand ginst19071 (P3_R1077_U473, P3_R1077_U361, P3_R1077_U92);
  nand ginst19072 (P3_R1077_U474, P3_R1077_U262, P3_R1077_U472);
  nand ginst19073 (P3_R1077_U475, P3_R1077_U73, P3_U3073);
  nand ginst19074 (P3_R1077_U476, P3_R1077_U74, P3_U3434);
  nand ginst19075 (P3_R1077_U477, P3_R1077_U73, P3_U3073);
  nand ginst19076 (P3_R1077_U478, P3_R1077_U74, P3_U3434);
  nand ginst19077 (P3_R1077_U479, P3_R1077_U477, P3_R1077_U478);
  not ginst19078 (P3_R1077_U48, P3_U3056);
  nand ginst19079 (P3_R1077_U480, P3_R1077_U163, P3_R1077_U164);
  nand ginst19080 (P3_R1077_U481, P3_R1077_U258, P3_R1077_U479);
  nand ginst19081 (P3_R1077_U482, P3_R1077_U71, P3_U3078);
  nand ginst19082 (P3_R1077_U483, P3_R1077_U72, P3_U3431);
  nand ginst19083 (P3_R1077_U484, P3_R1077_U71, P3_U3078);
  nand ginst19084 (P3_R1077_U485, P3_R1077_U72, P3_U3431);
  nand ginst19085 (P3_R1077_U486, P3_R1077_U484, P3_R1077_U485);
  nand ginst19086 (P3_R1077_U487, P3_R1077_U165, P3_R1077_U166);
  nand ginst19087 (P3_R1077_U488, P3_R1077_U254, P3_R1077_U486);
  nand ginst19088 (P3_R1077_U489, P3_R1077_U69, P3_U3079);
  not ginst19089 (P3_R1077_U49, P3_U3901);
  nand ginst19090 (P3_R1077_U490, P3_R1077_U70, P3_U3428);
  nand ginst19091 (P3_R1077_U491, P3_R1077_U64, P3_U3071);
  nand ginst19092 (P3_R1077_U492, P3_R1077_U65, P3_U3425);
  nand ginst19093 (P3_R1077_U493, P3_R1077_U491, P3_R1077_U492);
  nand ginst19094 (P3_R1077_U494, P3_R1077_U362, P3_R1077_U93);
  nand ginst19095 (P3_R1077_U495, P3_R1077_U338, P3_R1077_U493);
  nand ginst19096 (P3_R1077_U496, P3_R1077_U66, P3_U3062);
  nand ginst19097 (P3_R1077_U497, P3_R1077_U67, P3_U3422);
  nand ginst19098 (P3_R1077_U498, P3_R1077_U496, P3_R1077_U497);
  nand ginst19099 (P3_R1077_U499, P3_R1077_U167, P3_R1077_U363);
  and ginst19100 (P3_R1077_U5, P3_R1077_U196, P3_R1077_U197);
  not ginst19101 (P3_R1077_U50, P3_U3902);
  nand ginst19102 (P3_R1077_U500, P3_R1077_U244, P3_R1077_U498);
  nand ginst19103 (P3_R1077_U501, P3_R1077_U62, P3_U3061);
  nand ginst19104 (P3_R1077_U502, P3_R1077_U63, P3_U3419);
  nand ginst19105 (P3_R1077_U503, P3_R1077_U29, P3_U3076);
  nand ginst19106 (P3_R1077_U504, P3_R1077_U30, P3_U3387);
  not ginst19107 (P3_R1077_U51, P3_U3057);
  not ginst19108 (P3_R1077_U52, P3_U3903);
  not ginst19109 (P3_R1077_U53, P3_U3064);
  not ginst19110 (P3_R1077_U54, P3_U3906);
  not ginst19111 (P3_R1077_U55, P3_U3074);
  not ginst19112 (P3_R1077_U56, P3_U3437);
  not ginst19113 (P3_R1077_U57, P3_U3072);
  not ginst19114 (P3_R1077_U58, P3_U3068);
  nand ginst19115 (P3_R1077_U59, P3_U3072, P3_U3437);
  and ginst19116 (P3_R1077_U6, P3_R1077_U236, P3_R1077_U237);
  not ginst19117 (P3_R1077_U60, P3_U3440);
  nand ginst19118 (P3_R1077_U61, P3_U3083, P3_U3413);
  not ginst19119 (P3_R1077_U62, P3_U3419);
  not ginst19120 (P3_R1077_U63, P3_U3061);
  not ginst19121 (P3_R1077_U64, P3_U3425);
  not ginst19122 (P3_R1077_U65, P3_U3071);
  not ginst19123 (P3_R1077_U66, P3_U3422);
  not ginst19124 (P3_R1077_U67, P3_U3062);
  nand ginst19125 (P3_R1077_U68, P3_U3062, P3_U3422);
  not ginst19126 (P3_R1077_U69, P3_U3428);
  and ginst19127 (P3_R1077_U7, P3_R1077_U245, P3_R1077_U246);
  not ginst19128 (P3_R1077_U70, P3_U3079);
  not ginst19129 (P3_R1077_U71, P3_U3431);
  not ginst19130 (P3_R1077_U72, P3_U3078);
  not ginst19131 (P3_R1077_U73, P3_U3434);
  not ginst19132 (P3_R1077_U74, P3_U3073);
  not ginst19133 (P3_R1077_U75, P3_U3443);
  not ginst19134 (P3_R1077_U76, P3_U3081);
  nand ginst19135 (P3_R1077_U77, P3_U3081, P3_U3443);
  not ginst19136 (P3_R1077_U78, P3_U3445);
  not ginst19137 (P3_R1077_U79, P3_U3080);
  and ginst19138 (P3_R1077_U8, P3_R1077_U263, P3_R1077_U264);
  nand ginst19139 (P3_R1077_U80, P3_U3080, P3_U3445);
  not ginst19140 (P3_R1077_U81, P3_U3907);
  not ginst19141 (P3_R1077_U82, P3_U3905);
  not ginst19142 (P3_R1077_U83, P3_U3060);
  not ginst19143 (P3_R1077_U84, P3_U3904);
  not ginst19144 (P3_R1077_U85, P3_U3065);
  nand ginst19145 (P3_R1077_U86, P3_U3056, P3_U3901);
  not ginst19146 (P3_R1077_U87, P3_U3053);
  not ginst19147 (P3_R1077_U88, P3_U3899);
  nand ginst19148 (P3_R1077_U89, P3_R1077_U176, P3_R1077_U306);
  and ginst19149 (P3_R1077_U9, P3_R1077_U271, P3_R1077_U272);
  not ginst19150 (P3_R1077_U90, P3_U3075);
  nand ginst19151 (P3_R1077_U91, P3_R1077_U315, P3_R1077_U77);
  nand ginst19152 (P3_R1077_U92, P3_R1077_U260, P3_R1077_U261);
  nand ginst19153 (P3_R1077_U93, P3_R1077_U337, P3_R1077_U68);
  nand ginst19154 (P3_R1077_U94, P3_R1077_U456, P3_R1077_U457);
  nand ginst19155 (P3_R1077_U95, P3_R1077_U503, P3_R1077_U504);
  nand ginst19156 (P3_R1077_U96, P3_R1077_U374, P3_R1077_U375);
  nand ginst19157 (P3_R1077_U97, P3_R1077_U379, P3_R1077_U380);
  nand ginst19158 (P3_R1077_U98, P3_R1077_U386, P3_R1077_U387);
  nand ginst19159 (P3_R1077_U99, P3_R1077_U393, P3_R1077_U394);
  and ginst19160 (P3_R1095_U10, P3_R1095_U263, P3_R1095_U264);
  nand ginst19161 (P3_R1095_U100, P3_R1095_U441, P3_R1095_U442);
  nand ginst19162 (P3_R1095_U101, P3_R1095_U446, P3_R1095_U447);
  nand ginst19163 (P3_R1095_U102, P3_R1095_U451, P3_R1095_U452);
  nand ginst19164 (P3_R1095_U103, P3_R1095_U456, P3_R1095_U457);
  nand ginst19165 (P3_R1095_U104, P3_R1095_U472, P3_R1095_U473);
  nand ginst19166 (P3_R1095_U105, P3_R1095_U477, P3_R1095_U478);
  nand ginst19167 (P3_R1095_U106, P3_R1095_U360, P3_R1095_U361);
  nand ginst19168 (P3_R1095_U107, P3_R1095_U369, P3_R1095_U370);
  nand ginst19169 (P3_R1095_U108, P3_R1095_U376, P3_R1095_U377);
  nand ginst19170 (P3_R1095_U109, P3_R1095_U380, P3_R1095_U381);
  and ginst19171 (P3_R1095_U11, P3_R1095_U191, P3_R1095_U286);
  nand ginst19172 (P3_R1095_U110, P3_R1095_U389, P3_R1095_U390);
  nand ginst19173 (P3_R1095_U111, P3_R1095_U410, P3_R1095_U411);
  nand ginst19174 (P3_R1095_U112, P3_R1095_U427, P3_R1095_U428);
  nand ginst19175 (P3_R1095_U113, P3_R1095_U431, P3_R1095_U432);
  nand ginst19176 (P3_R1095_U114, P3_R1095_U463, P3_R1095_U464);
  nand ginst19177 (P3_R1095_U115, P3_R1095_U467, P3_R1095_U468);
  nand ginst19178 (P3_R1095_U116, P3_R1095_U484, P3_R1095_U485);
  and ginst19179 (P3_R1095_U117, P3_R1095_U193, P3_R1095_U352);
  and ginst19180 (P3_R1095_U118, P3_R1095_U205, P3_R1095_U206);
  and ginst19181 (P3_R1095_U119, P3_R1095_U13, P3_R1095_U14);
  and ginst19182 (P3_R1095_U12, P3_R1095_U287, P3_R1095_U288);
  and ginst19183 (P3_R1095_U120, P3_R1095_U354, P3_R1095_U357);
  and ginst19184 (P3_R1095_U121, P3_R1095_U26, P3_R1095_U362, P3_R1095_U363);
  and ginst19185 (P3_R1095_U122, P3_R1095_U195, P3_R1095_U366);
  and ginst19186 (P3_R1095_U123, P3_R1095_U235, P3_R1095_U6);
  and ginst19187 (P3_R1095_U124, P3_R1095_U194, P3_R1095_U373);
  and ginst19188 (P3_R1095_U125, P3_R1095_U34, P3_R1095_U382, P3_R1095_U383);
  and ginst19189 (P3_R1095_U126, P3_R1095_U193, P3_R1095_U386);
  and ginst19190 (P3_R1095_U127, P3_R1095_U222, P3_R1095_U7);
  and ginst19191 (P3_R1095_U128, P3_R1095_U267, P3_R1095_U9);
  and ginst19192 (P3_R1095_U129, P3_R1095_U11, P3_R1095_U291);
  and ginst19193 (P3_R1095_U13, P3_R1095_U194, P3_R1095_U208, P3_R1095_U213);
  and ginst19194 (P3_R1095_U130, P3_R1095_U192, P3_R1095_U355);
  and ginst19195 (P3_R1095_U131, P3_R1095_U306, P3_R1095_U307);
  and ginst19196 (P3_R1095_U132, P3_R1095_U309, P3_R1095_U395);
  and ginst19197 (P3_R1095_U133, P3_R1095_U306, P3_R1095_U307);
  and ginst19198 (P3_R1095_U134, P3_R1095_U15, P3_R1095_U310);
  nand ginst19199 (P3_R1095_U135, P3_R1095_U398, P3_R1095_U399);
  and ginst19200 (P3_R1095_U136, P3_R1095_U403, P3_R1095_U404, P3_R1095_U87);
  and ginst19201 (P3_R1095_U137, P3_R1095_U192, P3_R1095_U407);
  nand ginst19202 (P3_R1095_U138, P3_R1095_U412, P3_R1095_U413);
  nand ginst19203 (P3_R1095_U139, P3_R1095_U417, P3_R1095_U418);
  and ginst19204 (P3_R1095_U14, P3_R1095_U195, P3_R1095_U218);
  and ginst19205 (P3_R1095_U140, P3_R1095_U12, P3_R1095_U322);
  and ginst19206 (P3_R1095_U141, P3_R1095_U191, P3_R1095_U424);
  nand ginst19207 (P3_R1095_U142, P3_R1095_U433, P3_R1095_U434);
  nand ginst19208 (P3_R1095_U143, P3_R1095_U438, P3_R1095_U439);
  nand ginst19209 (P3_R1095_U144, P3_R1095_U443, P3_R1095_U444);
  nand ginst19210 (P3_R1095_U145, P3_R1095_U448, P3_R1095_U449);
  nand ginst19211 (P3_R1095_U146, P3_R1095_U453, P3_R1095_U454);
  and ginst19212 (P3_R1095_U147, P3_R1095_U10, P3_R1095_U333);
  and ginst19213 (P3_R1095_U148, P3_R1095_U190, P3_R1095_U460);
  nand ginst19214 (P3_R1095_U149, P3_R1095_U469, P3_R1095_U470);
  and ginst19215 (P3_R1095_U15, P3_R1095_U391, P3_R1095_U392);
  nand ginst19216 (P3_R1095_U150, P3_R1095_U474, P3_R1095_U475);
  and ginst19217 (P3_R1095_U151, P3_R1095_U344, P3_R1095_U8);
  and ginst19218 (P3_R1095_U152, P3_R1095_U189, P3_R1095_U481);
  and ginst19219 (P3_R1095_U153, P3_R1095_U358, P3_R1095_U359);
  nand ginst19220 (P3_R1095_U154, P3_R1095_U120, P3_R1095_U356);
  and ginst19221 (P3_R1095_U155, P3_R1095_U367, P3_R1095_U368);
  and ginst19222 (P3_R1095_U156, P3_R1095_U374, P3_R1095_U375);
  and ginst19223 (P3_R1095_U157, P3_R1095_U378, P3_R1095_U379);
  nand ginst19224 (P3_R1095_U158, P3_R1095_U118, P3_R1095_U203);
  and ginst19225 (P3_R1095_U159, P3_R1095_U387, P3_R1095_U388);
  nand ginst19226 (P3_R1095_U16, P3_R1095_U342, P3_R1095_U345);
  not ginst19227 (P3_R1095_U160, P3_U3908);
  not ginst19228 (P3_R1095_U161, P3_U3054);
  and ginst19229 (P3_R1095_U162, P3_R1095_U396, P3_R1095_U397);
  nand ginst19230 (P3_R1095_U163, P3_R1095_U131, P3_R1095_U304);
  and ginst19231 (P3_R1095_U164, P3_R1095_U408, P3_R1095_U409);
  nand ginst19232 (P3_R1095_U165, P3_R1095_U297, P3_R1095_U298);
  nand ginst19233 (P3_R1095_U166, P3_R1095_U293, P3_R1095_U294);
  and ginst19234 (P3_R1095_U167, P3_R1095_U425, P3_R1095_U426);
  and ginst19235 (P3_R1095_U168, P3_R1095_U429, P3_R1095_U430);
  nand ginst19236 (P3_R1095_U169, P3_R1095_U283, P3_R1095_U284);
  nand ginst19237 (P3_R1095_U17, P3_R1095_U331, P3_R1095_U334);
  nand ginst19238 (P3_R1095_U170, P3_R1095_U279, P3_R1095_U280);
  not ginst19239 (P3_R1095_U171, P3_U3392);
  nand ginst19240 (P3_R1095_U172, P3_R1095_U95, P3_U3387);
  nand ginst19241 (P3_R1095_U173, P3_R1095_U184, P3_R1095_U276, P3_R1095_U350);
  not ginst19242 (P3_R1095_U174, P3_U3443);
  nand ginst19243 (P3_R1095_U175, P3_R1095_U273, P3_R1095_U274);
  nand ginst19244 (P3_R1095_U176, P3_R1095_U269, P3_R1095_U270);
  and ginst19245 (P3_R1095_U177, P3_R1095_U461, P3_R1095_U462);
  and ginst19246 (P3_R1095_U178, P3_R1095_U465, P3_R1095_U466);
  nand ginst19247 (P3_R1095_U179, P3_R1095_U259, P3_R1095_U260);
  nand ginst19248 (P3_R1095_U18, P3_R1095_U320, P3_R1095_U323);
  nand ginst19249 (P3_R1095_U180, P3_R1095_U255, P3_R1095_U256);
  nand ginst19250 (P3_R1095_U181, P3_R1095_U251, P3_R1095_U252);
  and ginst19251 (P3_R1095_U182, P3_R1095_U482, P3_R1095_U483);
  nand ginst19252 (P3_R1095_U183, P3_R1095_U132, P3_R1095_U163);
  nand ginst19253 (P3_R1095_U184, P3_R1095_U174, P3_R1095_U175);
  nand ginst19254 (P3_R1095_U185, P3_R1095_U171, P3_R1095_U172);
  not ginst19255 (P3_R1095_U186, P3_R1095_U87);
  not ginst19256 (P3_R1095_U187, P3_R1095_U34);
  not ginst19257 (P3_R1095_U188, P3_R1095_U26);
  nand ginst19258 (P3_R1095_U189, P3_R1095_U54, P3_U3419);
  nand ginst19259 (P3_R1095_U19, P3_R1095_U312, P3_R1095_U314);
  nand ginst19260 (P3_R1095_U190, P3_R1095_U64, P3_U3434);
  nand ginst19261 (P3_R1095_U191, P3_R1095_U78, P3_U3905);
  nand ginst19262 (P3_R1095_U192, P3_R1095_U86, P3_U3901);
  nand ginst19263 (P3_R1095_U193, P3_R1095_U33, P3_U3395);
  nand ginst19264 (P3_R1095_U194, P3_R1095_U41, P3_U3404);
  nand ginst19265 (P3_R1095_U195, P3_R1095_U25, P3_U3410);
  not ginst19266 (P3_R1095_U196, P3_R1095_U66);
  not ginst19267 (P3_R1095_U197, P3_R1095_U80);
  not ginst19268 (P3_R1095_U198, P3_R1095_U43);
  not ginst19269 (P3_R1095_U199, P3_R1095_U55);
  nand ginst19270 (P3_R1095_U20, P3_R1095_U162, P3_R1095_U183, P3_R1095_U351);
  not ginst19271 (P3_R1095_U200, P3_R1095_U172);
  nand ginst19272 (P3_R1095_U201, P3_R1095_U172, P3_U3077);
  not ginst19273 (P3_R1095_U202, P3_R1095_U49);
  nand ginst19274 (P3_R1095_U203, P3_R1095_U117, P3_R1095_U49);
  nand ginst19275 (P3_R1095_U204, P3_R1095_U34, P3_R1095_U35);
  nand ginst19276 (P3_R1095_U205, P3_R1095_U204, P3_R1095_U32);
  nand ginst19277 (P3_R1095_U206, P3_R1095_U187, P3_U3063);
  not ginst19278 (P3_R1095_U207, P3_R1095_U158);
  nand ginst19279 (P3_R1095_U208, P3_R1095_U40, P3_U3407);
  nand ginst19280 (P3_R1095_U209, P3_R1095_U37, P3_U3070);
  nand ginst19281 (P3_R1095_U21, P3_R1095_U241, P3_R1095_U243);
  nand ginst19282 (P3_R1095_U210, P3_R1095_U36, P3_U3066);
  nand ginst19283 (P3_R1095_U211, P3_R1095_U194, P3_R1095_U198);
  nand ginst19284 (P3_R1095_U212, P3_R1095_U211, P3_R1095_U6);
  nand ginst19285 (P3_R1095_U213, P3_R1095_U42, P3_U3401);
  nand ginst19286 (P3_R1095_U214, P3_R1095_U40, P3_U3407);
  nand ginst19287 (P3_R1095_U215, P3_R1095_U13, P3_R1095_U158);
  not ginst19288 (P3_R1095_U216, P3_R1095_U44);
  not ginst19289 (P3_R1095_U217, P3_R1095_U47);
  nand ginst19290 (P3_R1095_U218, P3_R1095_U27, P3_U3413);
  nand ginst19291 (P3_R1095_U219, P3_R1095_U26, P3_R1095_U27);
  nand ginst19292 (P3_R1095_U22, P3_R1095_U233, P3_R1095_U236);
  nand ginst19293 (P3_R1095_U220, P3_R1095_U188, P3_U3083);
  not ginst19294 (P3_R1095_U221, P3_R1095_U154);
  nand ginst19295 (P3_R1095_U222, P3_R1095_U46, P3_U3416);
  nand ginst19296 (P3_R1095_U223, P3_R1095_U222, P3_R1095_U55);
  nand ginst19297 (P3_R1095_U224, P3_R1095_U217, P3_R1095_U26);
  nand ginst19298 (P3_R1095_U225, P3_R1095_U122, P3_R1095_U224);
  nand ginst19299 (P3_R1095_U226, P3_R1095_U195, P3_R1095_U47);
  nand ginst19300 (P3_R1095_U227, P3_R1095_U121, P3_R1095_U226);
  nand ginst19301 (P3_R1095_U228, P3_R1095_U195, P3_R1095_U26);
  nand ginst19302 (P3_R1095_U229, P3_R1095_U158, P3_R1095_U213);
  nand ginst19303 (P3_R1095_U23, P3_R1095_U225, P3_R1095_U227);
  not ginst19304 (P3_R1095_U230, P3_R1095_U48);
  nand ginst19305 (P3_R1095_U231, P3_R1095_U36, P3_U3066);
  nand ginst19306 (P3_R1095_U232, P3_R1095_U230, P3_R1095_U231);
  nand ginst19307 (P3_R1095_U233, P3_R1095_U124, P3_R1095_U232);
  nand ginst19308 (P3_R1095_U234, P3_R1095_U194, P3_R1095_U48);
  nand ginst19309 (P3_R1095_U235, P3_R1095_U40, P3_U3407);
  nand ginst19310 (P3_R1095_U236, P3_R1095_U123, P3_R1095_U234);
  nand ginst19311 (P3_R1095_U237, P3_R1095_U36, P3_U3066);
  nand ginst19312 (P3_R1095_U238, P3_R1095_U194, P3_R1095_U237);
  nand ginst19313 (P3_R1095_U239, P3_R1095_U213, P3_R1095_U43);
  nand ginst19314 (P3_R1095_U24, P3_R1095_U172, P3_R1095_U348);
  nand ginst19315 (P3_R1095_U240, P3_R1095_U202, P3_R1095_U34);
  nand ginst19316 (P3_R1095_U241, P3_R1095_U126, P3_R1095_U240);
  nand ginst19317 (P3_R1095_U242, P3_R1095_U193, P3_R1095_U49);
  nand ginst19318 (P3_R1095_U243, P3_R1095_U125, P3_R1095_U242);
  nand ginst19319 (P3_R1095_U244, P3_R1095_U193, P3_R1095_U34);
  nand ginst19320 (P3_R1095_U245, P3_R1095_U53, P3_U3422);
  nand ginst19321 (P3_R1095_U246, P3_R1095_U51, P3_U3062);
  nand ginst19322 (P3_R1095_U247, P3_R1095_U52, P3_U3061);
  nand ginst19323 (P3_R1095_U248, P3_R1095_U199, P3_R1095_U7);
  nand ginst19324 (P3_R1095_U249, P3_R1095_U248, P3_R1095_U8);
  not ginst19325 (P3_R1095_U25, P3_U3069);
  nand ginst19326 (P3_R1095_U250, P3_R1095_U53, P3_U3422);
  nand ginst19327 (P3_R1095_U251, P3_R1095_U127, P3_R1095_U154);
  nand ginst19328 (P3_R1095_U252, P3_R1095_U249, P3_R1095_U250);
  not ginst19329 (P3_R1095_U253, P3_R1095_U181);
  nand ginst19330 (P3_R1095_U254, P3_R1095_U57, P3_U3425);
  nand ginst19331 (P3_R1095_U255, P3_R1095_U181, P3_R1095_U254);
  nand ginst19332 (P3_R1095_U256, P3_R1095_U56, P3_U3071);
  not ginst19333 (P3_R1095_U257, P3_R1095_U180);
  nand ginst19334 (P3_R1095_U258, P3_R1095_U59, P3_U3428);
  nand ginst19335 (P3_R1095_U259, P3_R1095_U180, P3_R1095_U258);
  nand ginst19336 (P3_R1095_U26, P3_R1095_U39, P3_U3069);
  nand ginst19337 (P3_R1095_U260, P3_R1095_U58, P3_U3079);
  not ginst19338 (P3_R1095_U261, P3_R1095_U179);
  nand ginst19339 (P3_R1095_U262, P3_R1095_U63, P3_U3437);
  nand ginst19340 (P3_R1095_U263, P3_R1095_U60, P3_U3072);
  nand ginst19341 (P3_R1095_U264, P3_R1095_U61, P3_U3073);
  nand ginst19342 (P3_R1095_U265, P3_R1095_U196, P3_R1095_U9);
  nand ginst19343 (P3_R1095_U266, P3_R1095_U10, P3_R1095_U265);
  nand ginst19344 (P3_R1095_U267, P3_R1095_U65, P3_U3431);
  nand ginst19345 (P3_R1095_U268, P3_R1095_U63, P3_U3437);
  nand ginst19346 (P3_R1095_U269, P3_R1095_U128, P3_R1095_U179);
  not ginst19347 (P3_R1095_U27, P3_U3083);
  nand ginst19348 (P3_R1095_U270, P3_R1095_U266, P3_R1095_U268);
  not ginst19349 (P3_R1095_U271, P3_R1095_U176);
  nand ginst19350 (P3_R1095_U272, P3_R1095_U68, P3_U3440);
  nand ginst19351 (P3_R1095_U273, P3_R1095_U176, P3_R1095_U272);
  nand ginst19352 (P3_R1095_U274, P3_R1095_U67, P3_U3068);
  not ginst19353 (P3_R1095_U275, P3_R1095_U175);
  nand ginst19354 (P3_R1095_U276, P3_R1095_U175, P3_U3081);
  not ginst19355 (P3_R1095_U277, P3_R1095_U173);
  nand ginst19356 (P3_R1095_U278, P3_R1095_U71, P3_U3445);
  nand ginst19357 (P3_R1095_U279, P3_R1095_U173, P3_R1095_U278);
  not ginst19358 (P3_R1095_U28, P3_U3413);
  nand ginst19359 (P3_R1095_U280, P3_R1095_U70, P3_U3080);
  not ginst19360 (P3_R1095_U281, P3_R1095_U170);
  nand ginst19361 (P3_R1095_U282, P3_R1095_U73, P3_U3907);
  nand ginst19362 (P3_R1095_U283, P3_R1095_U170, P3_R1095_U282);
  nand ginst19363 (P3_R1095_U284, P3_R1095_U72, P3_U3075);
  not ginst19364 (P3_R1095_U285, P3_R1095_U169);
  nand ginst19365 (P3_R1095_U286, P3_R1095_U77, P3_U3904);
  nand ginst19366 (P3_R1095_U287, P3_R1095_U74, P3_U3065);
  nand ginst19367 (P3_R1095_U288, P3_R1095_U75, P3_U3060);
  nand ginst19368 (P3_R1095_U289, P3_R1095_U11, P3_R1095_U197);
  not ginst19369 (P3_R1095_U29, P3_U3395);
  nand ginst19370 (P3_R1095_U290, P3_R1095_U12, P3_R1095_U289);
  nand ginst19371 (P3_R1095_U291, P3_R1095_U79, P3_U3906);
  nand ginst19372 (P3_R1095_U292, P3_R1095_U77, P3_U3904);
  nand ginst19373 (P3_R1095_U293, P3_R1095_U129, P3_R1095_U169);
  nand ginst19374 (P3_R1095_U294, P3_R1095_U290, P3_R1095_U292);
  not ginst19375 (P3_R1095_U295, P3_R1095_U166);
  nand ginst19376 (P3_R1095_U296, P3_R1095_U82, P3_U3903);
  nand ginst19377 (P3_R1095_U297, P3_R1095_U166, P3_R1095_U296);
  nand ginst19378 (P3_R1095_U298, P3_R1095_U81, P3_U3064);
  not ginst19379 (P3_R1095_U299, P3_R1095_U165);
  not ginst19380 (P3_R1095_U30, P3_U3387);
  nand ginst19381 (P3_R1095_U300, P3_R1095_U84, P3_U3902);
  nand ginst19382 (P3_R1095_U301, P3_R1095_U165, P3_R1095_U300);
  nand ginst19383 (P3_R1095_U302, P3_R1095_U83, P3_U3057);
  not ginst19384 (P3_R1095_U303, P3_R1095_U91);
  nand ginst19385 (P3_R1095_U304, P3_R1095_U130, P3_R1095_U91);
  nand ginst19386 (P3_R1095_U305, P3_R1095_U87, P3_R1095_U88);
  nand ginst19387 (P3_R1095_U306, P3_R1095_U305, P3_R1095_U85);
  nand ginst19388 (P3_R1095_U307, P3_R1095_U186, P3_U3052);
  not ginst19389 (P3_R1095_U308, P3_R1095_U163);
  nand ginst19390 (P3_R1095_U309, P3_R1095_U90, P3_U3899);
  not ginst19391 (P3_R1095_U31, P3_U3077);
  nand ginst19392 (P3_R1095_U310, P3_R1095_U89, P3_U3053);
  nand ginst19393 (P3_R1095_U311, P3_R1095_U303, P3_R1095_U87);
  nand ginst19394 (P3_R1095_U312, P3_R1095_U137, P3_R1095_U311);
  nand ginst19395 (P3_R1095_U313, P3_R1095_U192, P3_R1095_U91);
  nand ginst19396 (P3_R1095_U314, P3_R1095_U136, P3_R1095_U313);
  nand ginst19397 (P3_R1095_U315, P3_R1095_U192, P3_R1095_U87);
  nand ginst19398 (P3_R1095_U316, P3_R1095_U169, P3_R1095_U291);
  not ginst19399 (P3_R1095_U317, P3_R1095_U92);
  nand ginst19400 (P3_R1095_U318, P3_R1095_U75, P3_U3060);
  nand ginst19401 (P3_R1095_U319, P3_R1095_U317, P3_R1095_U318);
  not ginst19402 (P3_R1095_U32, P3_U3398);
  nand ginst19403 (P3_R1095_U320, P3_R1095_U141, P3_R1095_U319);
  nand ginst19404 (P3_R1095_U321, P3_R1095_U191, P3_R1095_U92);
  nand ginst19405 (P3_R1095_U322, P3_R1095_U77, P3_U3904);
  nand ginst19406 (P3_R1095_U323, P3_R1095_U140, P3_R1095_U321);
  nand ginst19407 (P3_R1095_U324, P3_R1095_U75, P3_U3060);
  nand ginst19408 (P3_R1095_U325, P3_R1095_U191, P3_R1095_U324);
  nand ginst19409 (P3_R1095_U326, P3_R1095_U291, P3_R1095_U80);
  nand ginst19410 (P3_R1095_U327, P3_R1095_U179, P3_R1095_U267);
  not ginst19411 (P3_R1095_U328, P3_R1095_U93);
  nand ginst19412 (P3_R1095_U329, P3_R1095_U61, P3_U3073);
  not ginst19413 (P3_R1095_U33, P3_U3067);
  nand ginst19414 (P3_R1095_U330, P3_R1095_U328, P3_R1095_U329);
  nand ginst19415 (P3_R1095_U331, P3_R1095_U148, P3_R1095_U330);
  nand ginst19416 (P3_R1095_U332, P3_R1095_U190, P3_R1095_U93);
  nand ginst19417 (P3_R1095_U333, P3_R1095_U63, P3_U3437);
  nand ginst19418 (P3_R1095_U334, P3_R1095_U147, P3_R1095_U332);
  nand ginst19419 (P3_R1095_U335, P3_R1095_U61, P3_U3073);
  nand ginst19420 (P3_R1095_U336, P3_R1095_U190, P3_R1095_U335);
  nand ginst19421 (P3_R1095_U337, P3_R1095_U267, P3_R1095_U66);
  nand ginst19422 (P3_R1095_U338, P3_R1095_U154, P3_R1095_U222);
  not ginst19423 (P3_R1095_U339, P3_R1095_U94);
  nand ginst19424 (P3_R1095_U34, P3_R1095_U29, P3_U3067);
  nand ginst19425 (P3_R1095_U340, P3_R1095_U52, P3_U3061);
  nand ginst19426 (P3_R1095_U341, P3_R1095_U339, P3_R1095_U340);
  nand ginst19427 (P3_R1095_U342, P3_R1095_U152, P3_R1095_U341);
  nand ginst19428 (P3_R1095_U343, P3_R1095_U189, P3_R1095_U94);
  nand ginst19429 (P3_R1095_U344, P3_R1095_U53, P3_U3422);
  nand ginst19430 (P3_R1095_U345, P3_R1095_U151, P3_R1095_U343);
  nand ginst19431 (P3_R1095_U346, P3_R1095_U52, P3_U3061);
  nand ginst19432 (P3_R1095_U347, P3_R1095_U189, P3_R1095_U346);
  nand ginst19433 (P3_R1095_U348, P3_R1095_U30, P3_U3076);
  nand ginst19434 (P3_R1095_U349, P3_R1095_U171, P3_U3077);
  not ginst19435 (P3_R1095_U35, P3_U3063);
  nand ginst19436 (P3_R1095_U350, P3_R1095_U174, P3_U3081);
  nand ginst19437 (P3_R1095_U351, P3_R1095_U133, P3_R1095_U134, P3_R1095_U304);
  nand ginst19438 (P3_R1095_U352, P3_R1095_U35, P3_U3398);
  nand ginst19439 (P3_R1095_U353, P3_R1095_U220, P3_U3413);
  nand ginst19440 (P3_R1095_U354, P3_R1095_U219, P3_R1095_U353);
  nand ginst19441 (P3_R1095_U355, P3_R1095_U88, P3_U3900);
  nand ginst19442 (P3_R1095_U356, P3_R1095_U119, P3_R1095_U158);
  nand ginst19443 (P3_R1095_U357, P3_R1095_U14, P3_R1095_U216);
  nand ginst19444 (P3_R1095_U358, P3_R1095_U46, P3_U3416);
  nand ginst19445 (P3_R1095_U359, P3_R1095_U45, P3_U3082);
  not ginst19446 (P3_R1095_U36, P3_U3404);
  nand ginst19447 (P3_R1095_U360, P3_R1095_U154, P3_R1095_U223);
  nand ginst19448 (P3_R1095_U361, P3_R1095_U153, P3_R1095_U221);
  nand ginst19449 (P3_R1095_U362, P3_R1095_U27, P3_U3413);
  nand ginst19450 (P3_R1095_U363, P3_R1095_U28, P3_U3083);
  nand ginst19451 (P3_R1095_U364, P3_R1095_U27, P3_U3413);
  nand ginst19452 (P3_R1095_U365, P3_R1095_U28, P3_U3083);
  nand ginst19453 (P3_R1095_U366, P3_R1095_U364, P3_R1095_U365);
  nand ginst19454 (P3_R1095_U367, P3_R1095_U25, P3_U3410);
  nand ginst19455 (P3_R1095_U368, P3_R1095_U39, P3_U3069);
  nand ginst19456 (P3_R1095_U369, P3_R1095_U228, P3_R1095_U47);
  not ginst19457 (P3_R1095_U37, P3_U3407);
  nand ginst19458 (P3_R1095_U370, P3_R1095_U155, P3_R1095_U217);
  nand ginst19459 (P3_R1095_U371, P3_R1095_U40, P3_U3407);
  nand ginst19460 (P3_R1095_U372, P3_R1095_U37, P3_U3070);
  nand ginst19461 (P3_R1095_U373, P3_R1095_U371, P3_R1095_U372);
  nand ginst19462 (P3_R1095_U374, P3_R1095_U41, P3_U3404);
  nand ginst19463 (P3_R1095_U375, P3_R1095_U36, P3_U3066);
  nand ginst19464 (P3_R1095_U376, P3_R1095_U238, P3_R1095_U48);
  nand ginst19465 (P3_R1095_U377, P3_R1095_U156, P3_R1095_U230);
  nand ginst19466 (P3_R1095_U378, P3_R1095_U42, P3_U3401);
  nand ginst19467 (P3_R1095_U379, P3_R1095_U38, P3_U3059);
  not ginst19468 (P3_R1095_U38, P3_U3401);
  nand ginst19469 (P3_R1095_U380, P3_R1095_U158, P3_R1095_U239);
  nand ginst19470 (P3_R1095_U381, P3_R1095_U157, P3_R1095_U207);
  nand ginst19471 (P3_R1095_U382, P3_R1095_U35, P3_U3398);
  nand ginst19472 (P3_R1095_U383, P3_R1095_U32, P3_U3063);
  nand ginst19473 (P3_R1095_U384, P3_R1095_U35, P3_U3398);
  nand ginst19474 (P3_R1095_U385, P3_R1095_U32, P3_U3063);
  nand ginst19475 (P3_R1095_U386, P3_R1095_U384, P3_R1095_U385);
  nand ginst19476 (P3_R1095_U387, P3_R1095_U33, P3_U3395);
  nand ginst19477 (P3_R1095_U388, P3_R1095_U29, P3_U3067);
  nand ginst19478 (P3_R1095_U389, P3_R1095_U244, P3_R1095_U49);
  not ginst19479 (P3_R1095_U39, P3_U3410);
  nand ginst19480 (P3_R1095_U390, P3_R1095_U159, P3_R1095_U202);
  nand ginst19481 (P3_R1095_U391, P3_R1095_U161, P3_U3908);
  nand ginst19482 (P3_R1095_U392, P3_R1095_U160, P3_U3054);
  nand ginst19483 (P3_R1095_U393, P3_R1095_U161, P3_U3908);
  nand ginst19484 (P3_R1095_U394, P3_R1095_U160, P3_U3054);
  nand ginst19485 (P3_R1095_U395, P3_R1095_U393, P3_R1095_U394);
  nand ginst19486 (P3_R1095_U396, P3_R1095_U395, P3_R1095_U89, P3_U3053);
  nand ginst19487 (P3_R1095_U397, P3_R1095_U15, P3_R1095_U90, P3_U3899);
  nand ginst19488 (P3_R1095_U398, P3_R1095_U90, P3_U3899);
  nand ginst19489 (P3_R1095_U399, P3_R1095_U89, P3_U3053);
  not ginst19490 (P3_R1095_U40, P3_U3070);
  not ginst19491 (P3_R1095_U400, P3_R1095_U135);
  nand ginst19492 (P3_R1095_U401, P3_R1095_U308, P3_R1095_U400);
  nand ginst19493 (P3_R1095_U402, P3_R1095_U135, P3_R1095_U163);
  nand ginst19494 (P3_R1095_U403, P3_R1095_U88, P3_U3900);
  nand ginst19495 (P3_R1095_U404, P3_R1095_U85, P3_U3052);
  nand ginst19496 (P3_R1095_U405, P3_R1095_U88, P3_U3900);
  nand ginst19497 (P3_R1095_U406, P3_R1095_U85, P3_U3052);
  nand ginst19498 (P3_R1095_U407, P3_R1095_U405, P3_R1095_U406);
  nand ginst19499 (P3_R1095_U408, P3_R1095_U86, P3_U3901);
  nand ginst19500 (P3_R1095_U409, P3_R1095_U50, P3_U3056);
  not ginst19501 (P3_R1095_U41, P3_U3066);
  nand ginst19502 (P3_R1095_U410, P3_R1095_U315, P3_R1095_U91);
  nand ginst19503 (P3_R1095_U411, P3_R1095_U164, P3_R1095_U303);
  nand ginst19504 (P3_R1095_U412, P3_R1095_U84, P3_U3902);
  nand ginst19505 (P3_R1095_U413, P3_R1095_U83, P3_U3057);
  not ginst19506 (P3_R1095_U414, P3_R1095_U138);
  nand ginst19507 (P3_R1095_U415, P3_R1095_U299, P3_R1095_U414);
  nand ginst19508 (P3_R1095_U416, P3_R1095_U138, P3_R1095_U165);
  nand ginst19509 (P3_R1095_U417, P3_R1095_U82, P3_U3903);
  nand ginst19510 (P3_R1095_U418, P3_R1095_U81, P3_U3064);
  not ginst19511 (P3_R1095_U419, P3_R1095_U139);
  not ginst19512 (P3_R1095_U42, P3_U3059);
  nand ginst19513 (P3_R1095_U420, P3_R1095_U295, P3_R1095_U419);
  nand ginst19514 (P3_R1095_U421, P3_R1095_U139, P3_R1095_U166);
  nand ginst19515 (P3_R1095_U422, P3_R1095_U77, P3_U3904);
  nand ginst19516 (P3_R1095_U423, P3_R1095_U74, P3_U3065);
  nand ginst19517 (P3_R1095_U424, P3_R1095_U422, P3_R1095_U423);
  nand ginst19518 (P3_R1095_U425, P3_R1095_U78, P3_U3905);
  nand ginst19519 (P3_R1095_U426, P3_R1095_U75, P3_U3060);
  nand ginst19520 (P3_R1095_U427, P3_R1095_U325, P3_R1095_U92);
  nand ginst19521 (P3_R1095_U428, P3_R1095_U167, P3_R1095_U317);
  nand ginst19522 (P3_R1095_U429, P3_R1095_U79, P3_U3906);
  nand ginst19523 (P3_R1095_U43, P3_R1095_U38, P3_U3059);
  nand ginst19524 (P3_R1095_U430, P3_R1095_U76, P3_U3074);
  nand ginst19525 (P3_R1095_U431, P3_R1095_U169, P3_R1095_U326);
  nand ginst19526 (P3_R1095_U432, P3_R1095_U168, P3_R1095_U285);
  nand ginst19527 (P3_R1095_U433, P3_R1095_U73, P3_U3907);
  nand ginst19528 (P3_R1095_U434, P3_R1095_U72, P3_U3075);
  not ginst19529 (P3_R1095_U435, P3_R1095_U142);
  nand ginst19530 (P3_R1095_U436, P3_R1095_U281, P3_R1095_U435);
  nand ginst19531 (P3_R1095_U437, P3_R1095_U142, P3_R1095_U170);
  nand ginst19532 (P3_R1095_U438, P3_R1095_U31, P3_U3392);
  nand ginst19533 (P3_R1095_U439, P3_R1095_U171, P3_U3077);
  nand ginst19534 (P3_R1095_U44, P3_R1095_U212, P3_R1095_U214);
  not ginst19535 (P3_R1095_U440, P3_R1095_U143);
  nand ginst19536 (P3_R1095_U441, P3_R1095_U200, P3_R1095_U440);
  nand ginst19537 (P3_R1095_U442, P3_R1095_U143, P3_R1095_U172);
  nand ginst19538 (P3_R1095_U443, P3_R1095_U71, P3_U3445);
  nand ginst19539 (P3_R1095_U444, P3_R1095_U70, P3_U3080);
  not ginst19540 (P3_R1095_U445, P3_R1095_U144);
  nand ginst19541 (P3_R1095_U446, P3_R1095_U277, P3_R1095_U445);
  nand ginst19542 (P3_R1095_U447, P3_R1095_U144, P3_R1095_U173);
  nand ginst19543 (P3_R1095_U448, P3_R1095_U69, P3_U3443);
  nand ginst19544 (P3_R1095_U449, P3_R1095_U174, P3_U3081);
  not ginst19545 (P3_R1095_U45, P3_U3416);
  not ginst19546 (P3_R1095_U450, P3_R1095_U145);
  nand ginst19547 (P3_R1095_U451, P3_R1095_U275, P3_R1095_U450);
  nand ginst19548 (P3_R1095_U452, P3_R1095_U145, P3_R1095_U175);
  nand ginst19549 (P3_R1095_U453, P3_R1095_U68, P3_U3440);
  nand ginst19550 (P3_R1095_U454, P3_R1095_U67, P3_U3068);
  not ginst19551 (P3_R1095_U455, P3_R1095_U146);
  nand ginst19552 (P3_R1095_U456, P3_R1095_U271, P3_R1095_U455);
  nand ginst19553 (P3_R1095_U457, P3_R1095_U146, P3_R1095_U176);
  nand ginst19554 (P3_R1095_U458, P3_R1095_U63, P3_U3437);
  nand ginst19555 (P3_R1095_U459, P3_R1095_U60, P3_U3072);
  not ginst19556 (P3_R1095_U46, P3_U3082);
  nand ginst19557 (P3_R1095_U460, P3_R1095_U458, P3_R1095_U459);
  nand ginst19558 (P3_R1095_U461, P3_R1095_U64, P3_U3434);
  nand ginst19559 (P3_R1095_U462, P3_R1095_U61, P3_U3073);
  nand ginst19560 (P3_R1095_U463, P3_R1095_U336, P3_R1095_U93);
  nand ginst19561 (P3_R1095_U464, P3_R1095_U177, P3_R1095_U328);
  nand ginst19562 (P3_R1095_U465, P3_R1095_U65, P3_U3431);
  nand ginst19563 (P3_R1095_U466, P3_R1095_U62, P3_U3078);
  nand ginst19564 (P3_R1095_U467, P3_R1095_U179, P3_R1095_U337);
  nand ginst19565 (P3_R1095_U468, P3_R1095_U178, P3_R1095_U261);
  nand ginst19566 (P3_R1095_U469, P3_R1095_U59, P3_U3428);
  nand ginst19567 (P3_R1095_U47, P3_R1095_U215, P3_R1095_U44);
  nand ginst19568 (P3_R1095_U470, P3_R1095_U58, P3_U3079);
  not ginst19569 (P3_R1095_U471, P3_R1095_U149);
  nand ginst19570 (P3_R1095_U472, P3_R1095_U257, P3_R1095_U471);
  nand ginst19571 (P3_R1095_U473, P3_R1095_U149, P3_R1095_U180);
  nand ginst19572 (P3_R1095_U474, P3_R1095_U57, P3_U3425);
  nand ginst19573 (P3_R1095_U475, P3_R1095_U56, P3_U3071);
  not ginst19574 (P3_R1095_U476, P3_R1095_U150);
  nand ginst19575 (P3_R1095_U477, P3_R1095_U253, P3_R1095_U476);
  nand ginst19576 (P3_R1095_U478, P3_R1095_U150, P3_R1095_U181);
  nand ginst19577 (P3_R1095_U479, P3_R1095_U53, P3_U3422);
  nand ginst19578 (P3_R1095_U48, P3_R1095_U229, P3_R1095_U43);
  nand ginst19579 (P3_R1095_U480, P3_R1095_U51, P3_U3062);
  nand ginst19580 (P3_R1095_U481, P3_R1095_U479, P3_R1095_U480);
  nand ginst19581 (P3_R1095_U482, P3_R1095_U54, P3_U3419);
  nand ginst19582 (P3_R1095_U483, P3_R1095_U52, P3_U3061);
  nand ginst19583 (P3_R1095_U484, P3_R1095_U347, P3_R1095_U94);
  nand ginst19584 (P3_R1095_U485, P3_R1095_U182, P3_R1095_U339);
  nand ginst19585 (P3_R1095_U49, P3_R1095_U185, P3_R1095_U201, P3_R1095_U349);
  not ginst19586 (P3_R1095_U50, P3_U3901);
  not ginst19587 (P3_R1095_U51, P3_U3422);
  not ginst19588 (P3_R1095_U52, P3_U3419);
  not ginst19589 (P3_R1095_U53, P3_U3062);
  not ginst19590 (P3_R1095_U54, P3_U3061);
  nand ginst19591 (P3_R1095_U55, P3_R1095_U45, P3_U3082);
  not ginst19592 (P3_R1095_U56, P3_U3425);
  not ginst19593 (P3_R1095_U57, P3_U3071);
  not ginst19594 (P3_R1095_U58, P3_U3428);
  not ginst19595 (P3_R1095_U59, P3_U3079);
  and ginst19596 (P3_R1095_U6, P3_R1095_U209, P3_R1095_U210);
  not ginst19597 (P3_R1095_U60, P3_U3437);
  not ginst19598 (P3_R1095_U61, P3_U3434);
  not ginst19599 (P3_R1095_U62, P3_U3431);
  not ginst19600 (P3_R1095_U63, P3_U3072);
  not ginst19601 (P3_R1095_U64, P3_U3073);
  not ginst19602 (P3_R1095_U65, P3_U3078);
  nand ginst19603 (P3_R1095_U66, P3_R1095_U62, P3_U3078);
  not ginst19604 (P3_R1095_U67, P3_U3440);
  not ginst19605 (P3_R1095_U68, P3_U3068);
  not ginst19606 (P3_R1095_U69, P3_U3081);
  and ginst19607 (P3_R1095_U7, P3_R1095_U189, P3_R1095_U245);
  not ginst19608 (P3_R1095_U70, P3_U3445);
  not ginst19609 (P3_R1095_U71, P3_U3080);
  not ginst19610 (P3_R1095_U72, P3_U3907);
  not ginst19611 (P3_R1095_U73, P3_U3075);
  not ginst19612 (P3_R1095_U74, P3_U3904);
  not ginst19613 (P3_R1095_U75, P3_U3905);
  not ginst19614 (P3_R1095_U76, P3_U3906);
  not ginst19615 (P3_R1095_U77, P3_U3065);
  not ginst19616 (P3_R1095_U78, P3_U3060);
  not ginst19617 (P3_R1095_U79, P3_U3074);
  and ginst19618 (P3_R1095_U8, P3_R1095_U246, P3_R1095_U247);
  nand ginst19619 (P3_R1095_U80, P3_R1095_U76, P3_U3074);
  not ginst19620 (P3_R1095_U81, P3_U3903);
  not ginst19621 (P3_R1095_U82, P3_U3064);
  not ginst19622 (P3_R1095_U83, P3_U3902);
  not ginst19623 (P3_R1095_U84, P3_U3057);
  not ginst19624 (P3_R1095_U85, P3_U3900);
  not ginst19625 (P3_R1095_U86, P3_U3056);
  nand ginst19626 (P3_R1095_U87, P3_R1095_U50, P3_U3056);
  not ginst19627 (P3_R1095_U88, P3_U3052);
  not ginst19628 (P3_R1095_U89, P3_U3899);
  and ginst19629 (P3_R1095_U9, P3_R1095_U190, P3_R1095_U262);
  not ginst19630 (P3_R1095_U90, P3_U3053);
  nand ginst19631 (P3_R1095_U91, P3_R1095_U301, P3_R1095_U302);
  nand ginst19632 (P3_R1095_U92, P3_R1095_U316, P3_R1095_U80);
  nand ginst19633 (P3_R1095_U93, P3_R1095_U327, P3_R1095_U66);
  nand ginst19634 (P3_R1095_U94, P3_R1095_U338, P3_R1095_U55);
  not ginst19635 (P3_R1095_U95, P3_U3076);
  nand ginst19636 (P3_R1095_U96, P3_R1095_U401, P3_R1095_U402);
  nand ginst19637 (P3_R1095_U97, P3_R1095_U415, P3_R1095_U416);
  nand ginst19638 (P3_R1095_U98, P3_R1095_U420, P3_R1095_U421);
  nand ginst19639 (P3_R1095_U99, P3_R1095_U436, P3_R1095_U437);
  and ginst19640 (P3_R1110_U10, P3_R1110_U348, P3_R1110_U351);
  nand ginst19641 (P3_R1110_U100, P3_R1110_U398, P3_R1110_U399);
  nand ginst19642 (P3_R1110_U101, P3_R1110_U407, P3_R1110_U408);
  nand ginst19643 (P3_R1110_U102, P3_R1110_U414, P3_R1110_U415);
  nand ginst19644 (P3_R1110_U103, P3_R1110_U421, P3_R1110_U422);
  nand ginst19645 (P3_R1110_U104, P3_R1110_U428, P3_R1110_U429);
  nand ginst19646 (P3_R1110_U105, P3_R1110_U433, P3_R1110_U434);
  nand ginst19647 (P3_R1110_U106, P3_R1110_U440, P3_R1110_U441);
  nand ginst19648 (P3_R1110_U107, P3_R1110_U447, P3_R1110_U448);
  nand ginst19649 (P3_R1110_U108, P3_R1110_U461, P3_R1110_U462);
  nand ginst19650 (P3_R1110_U109, P3_R1110_U466, P3_R1110_U467);
  and ginst19651 (P3_R1110_U11, P3_R1110_U341, P3_R1110_U344);
  nand ginst19652 (P3_R1110_U110, P3_R1110_U473, P3_R1110_U474);
  nand ginst19653 (P3_R1110_U111, P3_R1110_U480, P3_R1110_U481);
  nand ginst19654 (P3_R1110_U112, P3_R1110_U487, P3_R1110_U488);
  nand ginst19655 (P3_R1110_U113, P3_R1110_U494, P3_R1110_U495);
  nand ginst19656 (P3_R1110_U114, P3_R1110_U499, P3_R1110_U500);
  and ginst19657 (P3_R1110_U115, P3_R1110_U187, P3_R1110_U189);
  and ginst19658 (P3_R1110_U116, P3_R1110_U180, P3_R1110_U4);
  and ginst19659 (P3_R1110_U117, P3_R1110_U192, P3_R1110_U194);
  and ginst19660 (P3_R1110_U118, P3_R1110_U200, P3_R1110_U201);
  and ginst19661 (P3_R1110_U119, P3_R1110_U22, P3_R1110_U381, P3_R1110_U382);
  and ginst19662 (P3_R1110_U12, P3_R1110_U332, P3_R1110_U335);
  and ginst19663 (P3_R1110_U120, P3_R1110_U212, P3_R1110_U5);
  and ginst19664 (P3_R1110_U121, P3_R1110_U180, P3_R1110_U181);
  and ginst19665 (P3_R1110_U122, P3_R1110_U218, P3_R1110_U220);
  and ginst19666 (P3_R1110_U123, P3_R1110_U34, P3_R1110_U388, P3_R1110_U389);
  and ginst19667 (P3_R1110_U124, P3_R1110_U226, P3_R1110_U4);
  and ginst19668 (P3_R1110_U125, P3_R1110_U181, P3_R1110_U234);
  and ginst19669 (P3_R1110_U126, P3_R1110_U204, P3_R1110_U6);
  and ginst19670 (P3_R1110_U127, P3_R1110_U171, P3_R1110_U239);
  and ginst19671 (P3_R1110_U128, P3_R1110_U250, P3_R1110_U7);
  and ginst19672 (P3_R1110_U129, P3_R1110_U172, P3_R1110_U248);
  and ginst19673 (P3_R1110_U13, P3_R1110_U323, P3_R1110_U326);
  and ginst19674 (P3_R1110_U130, P3_R1110_U267, P3_R1110_U268);
  and ginst19675 (P3_R1110_U131, P3_R1110_U273, P3_R1110_U282, P3_R1110_U9);
  and ginst19676 (P3_R1110_U132, P3_R1110_U280, P3_R1110_U285);
  and ginst19677 (P3_R1110_U133, P3_R1110_U298, P3_R1110_U301);
  and ginst19678 (P3_R1110_U134, P3_R1110_U302, P3_R1110_U368);
  and ginst19679 (P3_R1110_U135, P3_R1110_U160, P3_R1110_U278);
  and ginst19680 (P3_R1110_U136, P3_R1110_U454, P3_R1110_U455, P3_R1110_U80);
  and ginst19681 (P3_R1110_U137, P3_R1110_U325, P3_R1110_U9);
  and ginst19682 (P3_R1110_U138, P3_R1110_U468, P3_R1110_U469, P3_R1110_U59);
  and ginst19683 (P3_R1110_U139, P3_R1110_U334, P3_R1110_U8);
  and ginst19684 (P3_R1110_U14, P3_R1110_U318, P3_R1110_U320);
  and ginst19685 (P3_R1110_U140, P3_R1110_U172, P3_R1110_U489, P3_R1110_U490);
  and ginst19686 (P3_R1110_U141, P3_R1110_U343, P3_R1110_U7);
  and ginst19687 (P3_R1110_U142, P3_R1110_U171, P3_R1110_U501, P3_R1110_U502);
  and ginst19688 (P3_R1110_U143, P3_R1110_U350, P3_R1110_U6);
  nand ginst19689 (P3_R1110_U144, P3_R1110_U118, P3_R1110_U202);
  nand ginst19690 (P3_R1110_U145, P3_R1110_U217, P3_R1110_U229);
  not ginst19691 (P3_R1110_U146, P3_U3054);
  not ginst19692 (P3_R1110_U147, P3_U3908);
  and ginst19693 (P3_R1110_U148, P3_R1110_U402, P3_R1110_U403);
  nand ginst19694 (P3_R1110_U149, P3_R1110_U169, P3_R1110_U304, P3_R1110_U364);
  and ginst19695 (P3_R1110_U15, P3_R1110_U310, P3_R1110_U313);
  and ginst19696 (P3_R1110_U150, P3_R1110_U409, P3_R1110_U410);
  nand ginst19697 (P3_R1110_U151, P3_R1110_U134, P3_R1110_U369, P3_R1110_U370);
  and ginst19698 (P3_R1110_U152, P3_R1110_U416, P3_R1110_U417);
  nand ginst19699 (P3_R1110_U153, P3_R1110_U299, P3_R1110_U365, P3_R1110_U86);
  and ginst19700 (P3_R1110_U154, P3_R1110_U423, P3_R1110_U424);
  nand ginst19701 (P3_R1110_U155, P3_R1110_U292, P3_R1110_U293);
  and ginst19702 (P3_R1110_U156, P3_R1110_U435, P3_R1110_U436);
  nand ginst19703 (P3_R1110_U157, P3_R1110_U288, P3_R1110_U289);
  and ginst19704 (P3_R1110_U158, P3_R1110_U442, P3_R1110_U443);
  nand ginst19705 (P3_R1110_U159, P3_R1110_U132, P3_R1110_U284);
  and ginst19706 (P3_R1110_U16, P3_R1110_U232, P3_R1110_U235);
  and ginst19707 (P3_R1110_U160, P3_R1110_U449, P3_R1110_U450);
  nand ginst19708 (P3_R1110_U161, P3_R1110_U327, P3_R1110_U43);
  nand ginst19709 (P3_R1110_U162, P3_R1110_U130, P3_R1110_U269);
  and ginst19710 (P3_R1110_U163, P3_R1110_U475, P3_R1110_U476);
  nand ginst19711 (P3_R1110_U164, P3_R1110_U256, P3_R1110_U257);
  and ginst19712 (P3_R1110_U165, P3_R1110_U482, P3_R1110_U483);
  nand ginst19713 (P3_R1110_U166, P3_R1110_U252, P3_R1110_U253);
  nand ginst19714 (P3_R1110_U167, P3_R1110_U242, P3_R1110_U243);
  nand ginst19715 (P3_R1110_U168, P3_R1110_U366, P3_R1110_U367);
  nand ginst19716 (P3_R1110_U169, P3_R1110_U151, P3_U3053);
  and ginst19717 (P3_R1110_U17, P3_R1110_U224, P3_R1110_U227);
  not ginst19718 (P3_R1110_U170, P3_R1110_U34);
  nand ginst19719 (P3_R1110_U171, P3_U3082, P3_U3416);
  nand ginst19720 (P3_R1110_U172, P3_U3071, P3_U3425);
  nand ginst19721 (P3_R1110_U173, P3_U3057, P3_U3902);
  not ginst19722 (P3_R1110_U174, P3_R1110_U68);
  not ginst19723 (P3_R1110_U175, P3_R1110_U77);
  nand ginst19724 (P3_R1110_U176, P3_U3064, P3_U3903);
  not ginst19725 (P3_R1110_U177, P3_R1110_U61);
  or ginst19726 (P3_R1110_U178, P3_U3066, P3_U3404);
  or ginst19727 (P3_R1110_U179, P3_U3059, P3_U3401);
  and ginst19728 (P3_R1110_U18, P3_R1110_U210, P3_R1110_U213);
  or ginst19729 (P3_R1110_U180, P3_U3063, P3_U3398);
  or ginst19730 (P3_R1110_U181, P3_U3067, P3_U3395);
  not ginst19731 (P3_R1110_U182, P3_R1110_U31);
  or ginst19732 (P3_R1110_U183, P3_U3077, P3_U3392);
  not ginst19733 (P3_R1110_U184, P3_R1110_U42);
  not ginst19734 (P3_R1110_U185, P3_R1110_U43);
  nand ginst19735 (P3_R1110_U186, P3_R1110_U42, P3_R1110_U43);
  nand ginst19736 (P3_R1110_U187, P3_U3067, P3_U3395);
  nand ginst19737 (P3_R1110_U188, P3_R1110_U181, P3_R1110_U186);
  nand ginst19738 (P3_R1110_U189, P3_U3063, P3_U3398);
  not ginst19739 (P3_R1110_U19, P3_U3407);
  nand ginst19740 (P3_R1110_U190, P3_R1110_U115, P3_R1110_U188);
  nand ginst19741 (P3_R1110_U191, P3_R1110_U34, P3_R1110_U35);
  nand ginst19742 (P3_R1110_U192, P3_R1110_U191, P3_U3066);
  nand ginst19743 (P3_R1110_U193, P3_R1110_U116, P3_R1110_U190);
  nand ginst19744 (P3_R1110_U194, P3_R1110_U170, P3_U3404);
  not ginst19745 (P3_R1110_U195, P3_R1110_U41);
  or ginst19746 (P3_R1110_U196, P3_U3069, P3_U3410);
  or ginst19747 (P3_R1110_U197, P3_U3070, P3_U3407);
  not ginst19748 (P3_R1110_U198, P3_R1110_U22);
  nand ginst19749 (P3_R1110_U199, P3_R1110_U22, P3_R1110_U23);
  not ginst19750 (P3_R1110_U20, P3_U3070);
  nand ginst19751 (P3_R1110_U200, P3_R1110_U199, P3_U3069);
  nand ginst19752 (P3_R1110_U201, P3_R1110_U198, P3_U3410);
  nand ginst19753 (P3_R1110_U202, P3_R1110_U41, P3_R1110_U5);
  not ginst19754 (P3_R1110_U203, P3_R1110_U144);
  or ginst19755 (P3_R1110_U204, P3_U3083, P3_U3413);
  nand ginst19756 (P3_R1110_U205, P3_R1110_U144, P3_R1110_U204);
  not ginst19757 (P3_R1110_U206, P3_R1110_U40);
  or ginst19758 (P3_R1110_U207, P3_U3082, P3_U3416);
  or ginst19759 (P3_R1110_U208, P3_U3070, P3_U3407);
  nand ginst19760 (P3_R1110_U209, P3_R1110_U208, P3_R1110_U41);
  not ginst19761 (P3_R1110_U21, P3_U3069);
  nand ginst19762 (P3_R1110_U210, P3_R1110_U119, P3_R1110_U209);
  nand ginst19763 (P3_R1110_U211, P3_R1110_U195, P3_R1110_U22);
  nand ginst19764 (P3_R1110_U212, P3_U3069, P3_U3410);
  nand ginst19765 (P3_R1110_U213, P3_R1110_U120, P3_R1110_U211);
  or ginst19766 (P3_R1110_U214, P3_U3070, P3_U3407);
  nand ginst19767 (P3_R1110_U215, P3_R1110_U181, P3_R1110_U185);
  nand ginst19768 (P3_R1110_U216, P3_U3067, P3_U3395);
  not ginst19769 (P3_R1110_U217, P3_R1110_U45);
  nand ginst19770 (P3_R1110_U218, P3_R1110_U121, P3_R1110_U184);
  nand ginst19771 (P3_R1110_U219, P3_R1110_U180, P3_R1110_U45);
  nand ginst19772 (P3_R1110_U22, P3_U3070, P3_U3407);
  nand ginst19773 (P3_R1110_U220, P3_U3063, P3_U3398);
  not ginst19774 (P3_R1110_U221, P3_R1110_U44);
  or ginst19775 (P3_R1110_U222, P3_U3059, P3_U3401);
  nand ginst19776 (P3_R1110_U223, P3_R1110_U222, P3_R1110_U44);
  nand ginst19777 (P3_R1110_U224, P3_R1110_U123, P3_R1110_U223);
  nand ginst19778 (P3_R1110_U225, P3_R1110_U221, P3_R1110_U34);
  nand ginst19779 (P3_R1110_U226, P3_U3066, P3_U3404);
  nand ginst19780 (P3_R1110_U227, P3_R1110_U124, P3_R1110_U225);
  or ginst19781 (P3_R1110_U228, P3_U3059, P3_U3401);
  nand ginst19782 (P3_R1110_U229, P3_R1110_U181, P3_R1110_U184);
  not ginst19783 (P3_R1110_U23, P3_U3410);
  not ginst19784 (P3_R1110_U230, P3_R1110_U145);
  nand ginst19785 (P3_R1110_U231, P3_U3063, P3_U3398);
  nand ginst19786 (P3_R1110_U232, P3_R1110_U400, P3_R1110_U401, P3_R1110_U42, P3_R1110_U43);
  nand ginst19787 (P3_R1110_U233, P3_R1110_U42, P3_R1110_U43);
  nand ginst19788 (P3_R1110_U234, P3_U3067, P3_U3395);
  nand ginst19789 (P3_R1110_U235, P3_R1110_U125, P3_R1110_U233);
  or ginst19790 (P3_R1110_U236, P3_U3082, P3_U3416);
  or ginst19791 (P3_R1110_U237, P3_U3061, P3_U3419);
  nand ginst19792 (P3_R1110_U238, P3_R1110_U177, P3_R1110_U6);
  nand ginst19793 (P3_R1110_U239, P3_U3061, P3_U3419);
  not ginst19794 (P3_R1110_U24, P3_U3401);
  nand ginst19795 (P3_R1110_U240, P3_R1110_U127, P3_R1110_U238);
  or ginst19796 (P3_R1110_U241, P3_U3061, P3_U3419);
  nand ginst19797 (P3_R1110_U242, P3_R1110_U126, P3_R1110_U144);
  nand ginst19798 (P3_R1110_U243, P3_R1110_U240, P3_R1110_U241);
  not ginst19799 (P3_R1110_U244, P3_R1110_U167);
  or ginst19800 (P3_R1110_U245, P3_U3079, P3_U3428);
  or ginst19801 (P3_R1110_U246, P3_U3071, P3_U3425);
  nand ginst19802 (P3_R1110_U247, P3_R1110_U174, P3_R1110_U7);
  nand ginst19803 (P3_R1110_U248, P3_U3079, P3_U3428);
  nand ginst19804 (P3_R1110_U249, P3_R1110_U129, P3_R1110_U247);
  not ginst19805 (P3_R1110_U25, P3_U3059);
  or ginst19806 (P3_R1110_U250, P3_U3062, P3_U3422);
  or ginst19807 (P3_R1110_U251, P3_U3079, P3_U3428);
  nand ginst19808 (P3_R1110_U252, P3_R1110_U128, P3_R1110_U167);
  nand ginst19809 (P3_R1110_U253, P3_R1110_U249, P3_R1110_U251);
  not ginst19810 (P3_R1110_U254, P3_R1110_U166);
  or ginst19811 (P3_R1110_U255, P3_U3078, P3_U3431);
  nand ginst19812 (P3_R1110_U256, P3_R1110_U166, P3_R1110_U255);
  nand ginst19813 (P3_R1110_U257, P3_U3078, P3_U3431);
  not ginst19814 (P3_R1110_U258, P3_R1110_U164);
  or ginst19815 (P3_R1110_U259, P3_U3073, P3_U3434);
  not ginst19816 (P3_R1110_U26, P3_U3066);
  nand ginst19817 (P3_R1110_U260, P3_R1110_U164, P3_R1110_U259);
  nand ginst19818 (P3_R1110_U261, P3_U3073, P3_U3434);
  not ginst19819 (P3_R1110_U262, P3_R1110_U92);
  or ginst19820 (P3_R1110_U263, P3_U3068, P3_U3440);
  or ginst19821 (P3_R1110_U264, P3_U3072, P3_U3437);
  not ginst19822 (P3_R1110_U265, P3_R1110_U59);
  nand ginst19823 (P3_R1110_U266, P3_R1110_U59, P3_R1110_U60);
  nand ginst19824 (P3_R1110_U267, P3_R1110_U266, P3_U3068);
  nand ginst19825 (P3_R1110_U268, P3_R1110_U265, P3_U3440);
  nand ginst19826 (P3_R1110_U269, P3_R1110_U8, P3_R1110_U92);
  not ginst19827 (P3_R1110_U27, P3_U3395);
  not ginst19828 (P3_R1110_U270, P3_R1110_U162);
  or ginst19829 (P3_R1110_U271, P3_U3075, P3_U3907);
  or ginst19830 (P3_R1110_U272, P3_U3080, P3_U3445);
  or ginst19831 (P3_R1110_U273, P3_U3074, P3_U3906);
  not ginst19832 (P3_R1110_U274, P3_R1110_U80);
  nand ginst19833 (P3_R1110_U275, P3_R1110_U274, P3_U3907);
  nand ginst19834 (P3_R1110_U276, P3_R1110_U275, P3_R1110_U90);
  nand ginst19835 (P3_R1110_U277, P3_R1110_U80, P3_R1110_U81);
  nand ginst19836 (P3_R1110_U278, P3_R1110_U276, P3_R1110_U277);
  nand ginst19837 (P3_R1110_U279, P3_R1110_U175, P3_R1110_U9);
  not ginst19838 (P3_R1110_U28, P3_U3067);
  nand ginst19839 (P3_R1110_U280, P3_U3074, P3_U3906);
  nand ginst19840 (P3_R1110_U281, P3_R1110_U278, P3_R1110_U279);
  or ginst19841 (P3_R1110_U282, P3_U3081, P3_U3443);
  or ginst19842 (P3_R1110_U283, P3_U3074, P3_U3906);
  nand ginst19843 (P3_R1110_U284, P3_R1110_U131, P3_R1110_U162);
  nand ginst19844 (P3_R1110_U285, P3_R1110_U281, P3_R1110_U283);
  not ginst19845 (P3_R1110_U286, P3_R1110_U159);
  or ginst19846 (P3_R1110_U287, P3_U3060, P3_U3905);
  nand ginst19847 (P3_R1110_U288, P3_R1110_U159, P3_R1110_U287);
  nand ginst19848 (P3_R1110_U289, P3_U3060, P3_U3905);
  not ginst19849 (P3_R1110_U29, P3_U3387);
  not ginst19850 (P3_R1110_U290, P3_R1110_U157);
  or ginst19851 (P3_R1110_U291, P3_U3065, P3_U3904);
  nand ginst19852 (P3_R1110_U292, P3_R1110_U157, P3_R1110_U291);
  nand ginst19853 (P3_R1110_U293, P3_U3065, P3_U3904);
  not ginst19854 (P3_R1110_U294, P3_R1110_U155);
  or ginst19855 (P3_R1110_U295, P3_U3057, P3_U3902);
  nand ginst19856 (P3_R1110_U296, P3_R1110_U173, P3_R1110_U176);
  not ginst19857 (P3_R1110_U297, P3_R1110_U86);
  or ginst19858 (P3_R1110_U298, P3_U3064, P3_U3903);
  nand ginst19859 (P3_R1110_U299, P3_R1110_U155, P3_R1110_U168, P3_R1110_U298);
  not ginst19860 (P3_R1110_U30, P3_U3076);
  not ginst19861 (P3_R1110_U300, P3_R1110_U153);
  or ginst19862 (P3_R1110_U301, P3_U3052, P3_U3900);
  nand ginst19863 (P3_R1110_U302, P3_U3052, P3_U3900);
  not ginst19864 (P3_R1110_U303, P3_R1110_U151);
  nand ginst19865 (P3_R1110_U304, P3_R1110_U151, P3_U3899);
  not ginst19866 (P3_R1110_U305, P3_R1110_U149);
  nand ginst19867 (P3_R1110_U306, P3_R1110_U155, P3_R1110_U298);
  not ginst19868 (P3_R1110_U307, P3_R1110_U89);
  or ginst19869 (P3_R1110_U308, P3_U3057, P3_U3902);
  nand ginst19870 (P3_R1110_U309, P3_R1110_U308, P3_R1110_U89);
  nand ginst19871 (P3_R1110_U31, P3_U3076, P3_U3387);
  nand ginst19872 (P3_R1110_U310, P3_R1110_U154, P3_R1110_U173, P3_R1110_U309);
  nand ginst19873 (P3_R1110_U311, P3_R1110_U173, P3_R1110_U307);
  nand ginst19874 (P3_R1110_U312, P3_U3056, P3_U3901);
  nand ginst19875 (P3_R1110_U313, P3_R1110_U168, P3_R1110_U311, P3_R1110_U312);
  or ginst19876 (P3_R1110_U314, P3_U3057, P3_U3902);
  nand ginst19877 (P3_R1110_U315, P3_R1110_U162, P3_R1110_U282);
  not ginst19878 (P3_R1110_U316, P3_R1110_U91);
  nand ginst19879 (P3_R1110_U317, P3_R1110_U9, P3_R1110_U91);
  nand ginst19880 (P3_R1110_U318, P3_R1110_U135, P3_R1110_U317);
  nand ginst19881 (P3_R1110_U319, P3_R1110_U278, P3_R1110_U317);
  not ginst19882 (P3_R1110_U32, P3_U3398);
  nand ginst19883 (P3_R1110_U320, P3_R1110_U319, P3_R1110_U453);
  or ginst19884 (P3_R1110_U321, P3_U3080, P3_U3445);
  nand ginst19885 (P3_R1110_U322, P3_R1110_U321, P3_R1110_U91);
  nand ginst19886 (P3_R1110_U323, P3_R1110_U136, P3_R1110_U322);
  nand ginst19887 (P3_R1110_U324, P3_R1110_U316, P3_R1110_U80);
  nand ginst19888 (P3_R1110_U325, P3_U3075, P3_U3907);
  nand ginst19889 (P3_R1110_U326, P3_R1110_U137, P3_R1110_U324);
  or ginst19890 (P3_R1110_U327, P3_U3077, P3_U3392);
  not ginst19891 (P3_R1110_U328, P3_R1110_U161);
  or ginst19892 (P3_R1110_U329, P3_U3080, P3_U3445);
  not ginst19893 (P3_R1110_U33, P3_U3063);
  or ginst19894 (P3_R1110_U330, P3_U3072, P3_U3437);
  nand ginst19895 (P3_R1110_U331, P3_R1110_U330, P3_R1110_U92);
  nand ginst19896 (P3_R1110_U332, P3_R1110_U138, P3_R1110_U331);
  nand ginst19897 (P3_R1110_U333, P3_R1110_U262, P3_R1110_U59);
  nand ginst19898 (P3_R1110_U334, P3_U3068, P3_U3440);
  nand ginst19899 (P3_R1110_U335, P3_R1110_U139, P3_R1110_U333);
  or ginst19900 (P3_R1110_U336, P3_U3072, P3_U3437);
  nand ginst19901 (P3_R1110_U337, P3_R1110_U167, P3_R1110_U250);
  not ginst19902 (P3_R1110_U338, P3_R1110_U93);
  or ginst19903 (P3_R1110_U339, P3_U3071, P3_U3425);
  nand ginst19904 (P3_R1110_U34, P3_U3059, P3_U3401);
  nand ginst19905 (P3_R1110_U340, P3_R1110_U339, P3_R1110_U93);
  nand ginst19906 (P3_R1110_U341, P3_R1110_U140, P3_R1110_U340);
  nand ginst19907 (P3_R1110_U342, P3_R1110_U172, P3_R1110_U338);
  nand ginst19908 (P3_R1110_U343, P3_U3079, P3_U3428);
  nand ginst19909 (P3_R1110_U344, P3_R1110_U141, P3_R1110_U342);
  or ginst19910 (P3_R1110_U345, P3_U3071, P3_U3425);
  or ginst19911 (P3_R1110_U346, P3_U3082, P3_U3416);
  nand ginst19912 (P3_R1110_U347, P3_R1110_U346, P3_R1110_U40);
  nand ginst19913 (P3_R1110_U348, P3_R1110_U142, P3_R1110_U347);
  nand ginst19914 (P3_R1110_U349, P3_R1110_U171, P3_R1110_U206);
  not ginst19915 (P3_R1110_U35, P3_U3404);
  nand ginst19916 (P3_R1110_U350, P3_U3061, P3_U3419);
  nand ginst19917 (P3_R1110_U351, P3_R1110_U143, P3_R1110_U349);
  nand ginst19918 (P3_R1110_U352, P3_R1110_U171, P3_R1110_U207);
  nand ginst19919 (P3_R1110_U353, P3_R1110_U204, P3_R1110_U61);
  nand ginst19920 (P3_R1110_U354, P3_R1110_U214, P3_R1110_U22);
  nand ginst19921 (P3_R1110_U355, P3_R1110_U228, P3_R1110_U34);
  nand ginst19922 (P3_R1110_U356, P3_R1110_U180, P3_R1110_U231);
  nand ginst19923 (P3_R1110_U357, P3_R1110_U173, P3_R1110_U314);
  nand ginst19924 (P3_R1110_U358, P3_R1110_U176, P3_R1110_U298);
  nand ginst19925 (P3_R1110_U359, P3_R1110_U329, P3_R1110_U80);
  not ginst19926 (P3_R1110_U36, P3_U3413);
  nand ginst19927 (P3_R1110_U360, P3_R1110_U282, P3_R1110_U77);
  nand ginst19928 (P3_R1110_U361, P3_R1110_U336, P3_R1110_U59);
  nand ginst19929 (P3_R1110_U362, P3_R1110_U172, P3_R1110_U345);
  nand ginst19930 (P3_R1110_U363, P3_R1110_U250, P3_R1110_U68);
  nand ginst19931 (P3_R1110_U364, P3_U3053, P3_U3899);
  nand ginst19932 (P3_R1110_U365, P3_R1110_U168, P3_R1110_U296);
  nand ginst19933 (P3_R1110_U366, P3_R1110_U295, P3_U3056);
  nand ginst19934 (P3_R1110_U367, P3_R1110_U295, P3_U3901);
  nand ginst19935 (P3_R1110_U368, P3_R1110_U168, P3_R1110_U296, P3_R1110_U301);
  nand ginst19936 (P3_R1110_U369, P3_R1110_U133, P3_R1110_U155, P3_R1110_U168);
  not ginst19937 (P3_R1110_U37, P3_U3083);
  nand ginst19938 (P3_R1110_U370, P3_R1110_U297, P3_R1110_U301);
  nand ginst19939 (P3_R1110_U371, P3_R1110_U39, P3_U3082);
  nand ginst19940 (P3_R1110_U372, P3_R1110_U38, P3_U3416);
  nand ginst19941 (P3_R1110_U373, P3_R1110_U371, P3_R1110_U372);
  nand ginst19942 (P3_R1110_U374, P3_R1110_U352, P3_R1110_U40);
  nand ginst19943 (P3_R1110_U375, P3_R1110_U206, P3_R1110_U373);
  nand ginst19944 (P3_R1110_U376, P3_R1110_U36, P3_U3083);
  nand ginst19945 (P3_R1110_U377, P3_R1110_U37, P3_U3413);
  nand ginst19946 (P3_R1110_U378, P3_R1110_U376, P3_R1110_U377);
  nand ginst19947 (P3_R1110_U379, P3_R1110_U144, P3_R1110_U353);
  not ginst19948 (P3_R1110_U38, P3_U3082);
  nand ginst19949 (P3_R1110_U380, P3_R1110_U203, P3_R1110_U378);
  nand ginst19950 (P3_R1110_U381, P3_R1110_U23, P3_U3069);
  nand ginst19951 (P3_R1110_U382, P3_R1110_U21, P3_U3410);
  nand ginst19952 (P3_R1110_U383, P3_R1110_U19, P3_U3070);
  nand ginst19953 (P3_R1110_U384, P3_R1110_U20, P3_U3407);
  nand ginst19954 (P3_R1110_U385, P3_R1110_U383, P3_R1110_U384);
  nand ginst19955 (P3_R1110_U386, P3_R1110_U354, P3_R1110_U41);
  nand ginst19956 (P3_R1110_U387, P3_R1110_U195, P3_R1110_U385);
  nand ginst19957 (P3_R1110_U388, P3_R1110_U35, P3_U3066);
  nand ginst19958 (P3_R1110_U389, P3_R1110_U26, P3_U3404);
  not ginst19959 (P3_R1110_U39, P3_U3416);
  nand ginst19960 (P3_R1110_U390, P3_R1110_U24, P3_U3059);
  nand ginst19961 (P3_R1110_U391, P3_R1110_U25, P3_U3401);
  nand ginst19962 (P3_R1110_U392, P3_R1110_U390, P3_R1110_U391);
  nand ginst19963 (P3_R1110_U393, P3_R1110_U355, P3_R1110_U44);
  nand ginst19964 (P3_R1110_U394, P3_R1110_U221, P3_R1110_U392);
  nand ginst19965 (P3_R1110_U395, P3_R1110_U32, P3_U3063);
  nand ginst19966 (P3_R1110_U396, P3_R1110_U33, P3_U3398);
  nand ginst19967 (P3_R1110_U397, P3_R1110_U395, P3_R1110_U396);
  nand ginst19968 (P3_R1110_U398, P3_R1110_U145, P3_R1110_U356);
  nand ginst19969 (P3_R1110_U399, P3_R1110_U230, P3_R1110_U397);
  and ginst19970 (P3_R1110_U4, P3_R1110_U178, P3_R1110_U179);
  nand ginst19971 (P3_R1110_U40, P3_R1110_U205, P3_R1110_U61);
  nand ginst19972 (P3_R1110_U400, P3_R1110_U27, P3_U3067);
  nand ginst19973 (P3_R1110_U401, P3_R1110_U28, P3_U3395);
  nand ginst19974 (P3_R1110_U402, P3_R1110_U147, P3_U3054);
  nand ginst19975 (P3_R1110_U403, P3_R1110_U146, P3_U3908);
  nand ginst19976 (P3_R1110_U404, P3_R1110_U147, P3_U3054);
  nand ginst19977 (P3_R1110_U405, P3_R1110_U146, P3_U3908);
  nand ginst19978 (P3_R1110_U406, P3_R1110_U404, P3_R1110_U405);
  nand ginst19979 (P3_R1110_U407, P3_R1110_U148, P3_R1110_U149);
  nand ginst19980 (P3_R1110_U408, P3_R1110_U305, P3_R1110_U406);
  nand ginst19981 (P3_R1110_U409, P3_R1110_U88, P3_U3053);
  nand ginst19982 (P3_R1110_U41, P3_R1110_U117, P3_R1110_U193);
  nand ginst19983 (P3_R1110_U410, P3_R1110_U87, P3_U3899);
  nand ginst19984 (P3_R1110_U411, P3_R1110_U88, P3_U3053);
  nand ginst19985 (P3_R1110_U412, P3_R1110_U87, P3_U3899);
  nand ginst19986 (P3_R1110_U413, P3_R1110_U411, P3_R1110_U412);
  nand ginst19987 (P3_R1110_U414, P3_R1110_U150, P3_R1110_U151);
  nand ginst19988 (P3_R1110_U415, P3_R1110_U303, P3_R1110_U413);
  nand ginst19989 (P3_R1110_U416, P3_R1110_U46, P3_U3052);
  nand ginst19990 (P3_R1110_U417, P3_R1110_U47, P3_U3900);
  nand ginst19991 (P3_R1110_U418, P3_R1110_U46, P3_U3052);
  nand ginst19992 (P3_R1110_U419, P3_R1110_U47, P3_U3900);
  nand ginst19993 (P3_R1110_U42, P3_R1110_U182, P3_R1110_U183);
  nand ginst19994 (P3_R1110_U420, P3_R1110_U418, P3_R1110_U419);
  nand ginst19995 (P3_R1110_U421, P3_R1110_U152, P3_R1110_U153);
  nand ginst19996 (P3_R1110_U422, P3_R1110_U300, P3_R1110_U420);
  nand ginst19997 (P3_R1110_U423, P3_R1110_U49, P3_U3056);
  nand ginst19998 (P3_R1110_U424, P3_R1110_U48, P3_U3901);
  nand ginst19999 (P3_R1110_U425, P3_R1110_U50, P3_U3057);
  nand ginst20000 (P3_R1110_U426, P3_R1110_U51, P3_U3902);
  nand ginst20001 (P3_R1110_U427, P3_R1110_U425, P3_R1110_U426);
  nand ginst20002 (P3_R1110_U428, P3_R1110_U357, P3_R1110_U89);
  nand ginst20003 (P3_R1110_U429, P3_R1110_U307, P3_R1110_U427);
  nand ginst20004 (P3_R1110_U43, P3_U3077, P3_U3392);
  nand ginst20005 (P3_R1110_U430, P3_R1110_U52, P3_U3064);
  nand ginst20006 (P3_R1110_U431, P3_R1110_U53, P3_U3903);
  nand ginst20007 (P3_R1110_U432, P3_R1110_U430, P3_R1110_U431);
  nand ginst20008 (P3_R1110_U433, P3_R1110_U155, P3_R1110_U358);
  nand ginst20009 (P3_R1110_U434, P3_R1110_U294, P3_R1110_U432);
  nand ginst20010 (P3_R1110_U435, P3_R1110_U84, P3_U3065);
  nand ginst20011 (P3_R1110_U436, P3_R1110_U85, P3_U3904);
  nand ginst20012 (P3_R1110_U437, P3_R1110_U84, P3_U3065);
  nand ginst20013 (P3_R1110_U438, P3_R1110_U85, P3_U3904);
  nand ginst20014 (P3_R1110_U439, P3_R1110_U437, P3_R1110_U438);
  nand ginst20015 (P3_R1110_U44, P3_R1110_U122, P3_R1110_U219);
  nand ginst20016 (P3_R1110_U440, P3_R1110_U156, P3_R1110_U157);
  nand ginst20017 (P3_R1110_U441, P3_R1110_U290, P3_R1110_U439);
  nand ginst20018 (P3_R1110_U442, P3_R1110_U82, P3_U3060);
  nand ginst20019 (P3_R1110_U443, P3_R1110_U83, P3_U3905);
  nand ginst20020 (P3_R1110_U444, P3_R1110_U82, P3_U3060);
  nand ginst20021 (P3_R1110_U445, P3_R1110_U83, P3_U3905);
  nand ginst20022 (P3_R1110_U446, P3_R1110_U444, P3_R1110_U445);
  nand ginst20023 (P3_R1110_U447, P3_R1110_U158, P3_R1110_U159);
  nand ginst20024 (P3_R1110_U448, P3_R1110_U286, P3_R1110_U446);
  nand ginst20025 (P3_R1110_U449, P3_R1110_U54, P3_U3074);
  nand ginst20026 (P3_R1110_U45, P3_R1110_U215, P3_R1110_U216);
  nand ginst20027 (P3_R1110_U450, P3_R1110_U55, P3_U3906);
  nand ginst20028 (P3_R1110_U451, P3_R1110_U54, P3_U3074);
  nand ginst20029 (P3_R1110_U452, P3_R1110_U55, P3_U3906);
  nand ginst20030 (P3_R1110_U453, P3_R1110_U451, P3_R1110_U452);
  nand ginst20031 (P3_R1110_U454, P3_R1110_U81, P3_U3075);
  nand ginst20032 (P3_R1110_U455, P3_R1110_U90, P3_U3907);
  nand ginst20033 (P3_R1110_U456, P3_R1110_U161, P3_R1110_U182);
  nand ginst20034 (P3_R1110_U457, P3_R1110_U31, P3_R1110_U328);
  nand ginst20035 (P3_R1110_U458, P3_R1110_U78, P3_U3080);
  nand ginst20036 (P3_R1110_U459, P3_R1110_U79, P3_U3445);
  not ginst20037 (P3_R1110_U46, P3_U3900);
  nand ginst20038 (P3_R1110_U460, P3_R1110_U458, P3_R1110_U459);
  nand ginst20039 (P3_R1110_U461, P3_R1110_U359, P3_R1110_U91);
  nand ginst20040 (P3_R1110_U462, P3_R1110_U316, P3_R1110_U460);
  nand ginst20041 (P3_R1110_U463, P3_R1110_U75, P3_U3081);
  nand ginst20042 (P3_R1110_U464, P3_R1110_U76, P3_U3443);
  nand ginst20043 (P3_R1110_U465, P3_R1110_U463, P3_R1110_U464);
  nand ginst20044 (P3_R1110_U466, P3_R1110_U162, P3_R1110_U360);
  nand ginst20045 (P3_R1110_U467, P3_R1110_U270, P3_R1110_U465);
  nand ginst20046 (P3_R1110_U468, P3_R1110_U60, P3_U3068);
  nand ginst20047 (P3_R1110_U469, P3_R1110_U58, P3_U3440);
  not ginst20048 (P3_R1110_U47, P3_U3052);
  nand ginst20049 (P3_R1110_U470, P3_R1110_U56, P3_U3072);
  nand ginst20050 (P3_R1110_U471, P3_R1110_U57, P3_U3437);
  nand ginst20051 (P3_R1110_U472, P3_R1110_U470, P3_R1110_U471);
  nand ginst20052 (P3_R1110_U473, P3_R1110_U361, P3_R1110_U92);
  nand ginst20053 (P3_R1110_U474, P3_R1110_U262, P3_R1110_U472);
  nand ginst20054 (P3_R1110_U475, P3_R1110_U73, P3_U3073);
  nand ginst20055 (P3_R1110_U476, P3_R1110_U74, P3_U3434);
  nand ginst20056 (P3_R1110_U477, P3_R1110_U73, P3_U3073);
  nand ginst20057 (P3_R1110_U478, P3_R1110_U74, P3_U3434);
  nand ginst20058 (P3_R1110_U479, P3_R1110_U477, P3_R1110_U478);
  not ginst20059 (P3_R1110_U48, P3_U3056);
  nand ginst20060 (P3_R1110_U480, P3_R1110_U163, P3_R1110_U164);
  nand ginst20061 (P3_R1110_U481, P3_R1110_U258, P3_R1110_U479);
  nand ginst20062 (P3_R1110_U482, P3_R1110_U71, P3_U3078);
  nand ginst20063 (P3_R1110_U483, P3_R1110_U72, P3_U3431);
  nand ginst20064 (P3_R1110_U484, P3_R1110_U71, P3_U3078);
  nand ginst20065 (P3_R1110_U485, P3_R1110_U72, P3_U3431);
  nand ginst20066 (P3_R1110_U486, P3_R1110_U484, P3_R1110_U485);
  nand ginst20067 (P3_R1110_U487, P3_R1110_U165, P3_R1110_U166);
  nand ginst20068 (P3_R1110_U488, P3_R1110_U254, P3_R1110_U486);
  nand ginst20069 (P3_R1110_U489, P3_R1110_U69, P3_U3079);
  not ginst20070 (P3_R1110_U49, P3_U3901);
  nand ginst20071 (P3_R1110_U490, P3_R1110_U70, P3_U3428);
  nand ginst20072 (P3_R1110_U491, P3_R1110_U64, P3_U3071);
  nand ginst20073 (P3_R1110_U492, P3_R1110_U65, P3_U3425);
  nand ginst20074 (P3_R1110_U493, P3_R1110_U491, P3_R1110_U492);
  nand ginst20075 (P3_R1110_U494, P3_R1110_U362, P3_R1110_U93);
  nand ginst20076 (P3_R1110_U495, P3_R1110_U338, P3_R1110_U493);
  nand ginst20077 (P3_R1110_U496, P3_R1110_U66, P3_U3062);
  nand ginst20078 (P3_R1110_U497, P3_R1110_U67, P3_U3422);
  nand ginst20079 (P3_R1110_U498, P3_R1110_U496, P3_R1110_U497);
  nand ginst20080 (P3_R1110_U499, P3_R1110_U167, P3_R1110_U363);
  and ginst20081 (P3_R1110_U5, P3_R1110_U196, P3_R1110_U197);
  not ginst20082 (P3_R1110_U50, P3_U3902);
  nand ginst20083 (P3_R1110_U500, P3_R1110_U244, P3_R1110_U498);
  nand ginst20084 (P3_R1110_U501, P3_R1110_U62, P3_U3061);
  nand ginst20085 (P3_R1110_U502, P3_R1110_U63, P3_U3419);
  nand ginst20086 (P3_R1110_U503, P3_R1110_U29, P3_U3076);
  nand ginst20087 (P3_R1110_U504, P3_R1110_U30, P3_U3387);
  not ginst20088 (P3_R1110_U51, P3_U3057);
  not ginst20089 (P3_R1110_U52, P3_U3903);
  not ginst20090 (P3_R1110_U53, P3_U3064);
  not ginst20091 (P3_R1110_U54, P3_U3906);
  not ginst20092 (P3_R1110_U55, P3_U3074);
  not ginst20093 (P3_R1110_U56, P3_U3437);
  not ginst20094 (P3_R1110_U57, P3_U3072);
  not ginst20095 (P3_R1110_U58, P3_U3068);
  nand ginst20096 (P3_R1110_U59, P3_U3072, P3_U3437);
  and ginst20097 (P3_R1110_U6, P3_R1110_U236, P3_R1110_U237);
  not ginst20098 (P3_R1110_U60, P3_U3440);
  nand ginst20099 (P3_R1110_U61, P3_U3083, P3_U3413);
  not ginst20100 (P3_R1110_U62, P3_U3419);
  not ginst20101 (P3_R1110_U63, P3_U3061);
  not ginst20102 (P3_R1110_U64, P3_U3425);
  not ginst20103 (P3_R1110_U65, P3_U3071);
  not ginst20104 (P3_R1110_U66, P3_U3422);
  not ginst20105 (P3_R1110_U67, P3_U3062);
  nand ginst20106 (P3_R1110_U68, P3_U3062, P3_U3422);
  not ginst20107 (P3_R1110_U69, P3_U3428);
  and ginst20108 (P3_R1110_U7, P3_R1110_U245, P3_R1110_U246);
  not ginst20109 (P3_R1110_U70, P3_U3079);
  not ginst20110 (P3_R1110_U71, P3_U3431);
  not ginst20111 (P3_R1110_U72, P3_U3078);
  not ginst20112 (P3_R1110_U73, P3_U3434);
  not ginst20113 (P3_R1110_U74, P3_U3073);
  not ginst20114 (P3_R1110_U75, P3_U3443);
  not ginst20115 (P3_R1110_U76, P3_U3081);
  nand ginst20116 (P3_R1110_U77, P3_U3081, P3_U3443);
  not ginst20117 (P3_R1110_U78, P3_U3445);
  not ginst20118 (P3_R1110_U79, P3_U3080);
  and ginst20119 (P3_R1110_U8, P3_R1110_U263, P3_R1110_U264);
  nand ginst20120 (P3_R1110_U80, P3_U3080, P3_U3445);
  not ginst20121 (P3_R1110_U81, P3_U3907);
  not ginst20122 (P3_R1110_U82, P3_U3905);
  not ginst20123 (P3_R1110_U83, P3_U3060);
  not ginst20124 (P3_R1110_U84, P3_U3904);
  not ginst20125 (P3_R1110_U85, P3_U3065);
  nand ginst20126 (P3_R1110_U86, P3_U3056, P3_U3901);
  not ginst20127 (P3_R1110_U87, P3_U3053);
  not ginst20128 (P3_R1110_U88, P3_U3899);
  nand ginst20129 (P3_R1110_U89, P3_R1110_U176, P3_R1110_U306);
  and ginst20130 (P3_R1110_U9, P3_R1110_U271, P3_R1110_U272);
  not ginst20131 (P3_R1110_U90, P3_U3075);
  nand ginst20132 (P3_R1110_U91, P3_R1110_U315, P3_R1110_U77);
  nand ginst20133 (P3_R1110_U92, P3_R1110_U260, P3_R1110_U261);
  nand ginst20134 (P3_R1110_U93, P3_R1110_U337, P3_R1110_U68);
  nand ginst20135 (P3_R1110_U94, P3_R1110_U456, P3_R1110_U457);
  nand ginst20136 (P3_R1110_U95, P3_R1110_U503, P3_R1110_U504);
  nand ginst20137 (P3_R1110_U96, P3_R1110_U374, P3_R1110_U375);
  nand ginst20138 (P3_R1110_U97, P3_R1110_U379, P3_R1110_U380);
  nand ginst20139 (P3_R1110_U98, P3_R1110_U386, P3_R1110_U387);
  nand ginst20140 (P3_R1110_U99, P3_R1110_U393, P3_R1110_U394);
  and ginst20141 (P3_R1131_U10, P3_R1131_U263, P3_R1131_U264);
  nand ginst20142 (P3_R1131_U100, P3_R1131_U441, P3_R1131_U442);
  nand ginst20143 (P3_R1131_U101, P3_R1131_U446, P3_R1131_U447);
  nand ginst20144 (P3_R1131_U102, P3_R1131_U451, P3_R1131_U452);
  nand ginst20145 (P3_R1131_U103, P3_R1131_U456, P3_R1131_U457);
  nand ginst20146 (P3_R1131_U104, P3_R1131_U472, P3_R1131_U473);
  nand ginst20147 (P3_R1131_U105, P3_R1131_U477, P3_R1131_U478);
  nand ginst20148 (P3_R1131_U106, P3_R1131_U360, P3_R1131_U361);
  nand ginst20149 (P3_R1131_U107, P3_R1131_U369, P3_R1131_U370);
  nand ginst20150 (P3_R1131_U108, P3_R1131_U376, P3_R1131_U377);
  nand ginst20151 (P3_R1131_U109, P3_R1131_U380, P3_R1131_U381);
  and ginst20152 (P3_R1131_U11, P3_R1131_U191, P3_R1131_U286);
  nand ginst20153 (P3_R1131_U110, P3_R1131_U389, P3_R1131_U390);
  nand ginst20154 (P3_R1131_U111, P3_R1131_U410, P3_R1131_U411);
  nand ginst20155 (P3_R1131_U112, P3_R1131_U427, P3_R1131_U428);
  nand ginst20156 (P3_R1131_U113, P3_R1131_U431, P3_R1131_U432);
  nand ginst20157 (P3_R1131_U114, P3_R1131_U463, P3_R1131_U464);
  nand ginst20158 (P3_R1131_U115, P3_R1131_U467, P3_R1131_U468);
  nand ginst20159 (P3_R1131_U116, P3_R1131_U484, P3_R1131_U485);
  and ginst20160 (P3_R1131_U117, P3_R1131_U193, P3_R1131_U352);
  and ginst20161 (P3_R1131_U118, P3_R1131_U205, P3_R1131_U206);
  and ginst20162 (P3_R1131_U119, P3_R1131_U13, P3_R1131_U14);
  and ginst20163 (P3_R1131_U12, P3_R1131_U287, P3_R1131_U288);
  and ginst20164 (P3_R1131_U120, P3_R1131_U354, P3_R1131_U357);
  and ginst20165 (P3_R1131_U121, P3_R1131_U26, P3_R1131_U362, P3_R1131_U363);
  and ginst20166 (P3_R1131_U122, P3_R1131_U195, P3_R1131_U366);
  and ginst20167 (P3_R1131_U123, P3_R1131_U235, P3_R1131_U6);
  and ginst20168 (P3_R1131_U124, P3_R1131_U194, P3_R1131_U373);
  and ginst20169 (P3_R1131_U125, P3_R1131_U34, P3_R1131_U382, P3_R1131_U383);
  and ginst20170 (P3_R1131_U126, P3_R1131_U193, P3_R1131_U386);
  and ginst20171 (P3_R1131_U127, P3_R1131_U222, P3_R1131_U7);
  and ginst20172 (P3_R1131_U128, P3_R1131_U267, P3_R1131_U9);
  and ginst20173 (P3_R1131_U129, P3_R1131_U11, P3_R1131_U291);
  and ginst20174 (P3_R1131_U13, P3_R1131_U194, P3_R1131_U208, P3_R1131_U213);
  and ginst20175 (P3_R1131_U130, P3_R1131_U192, P3_R1131_U355);
  and ginst20176 (P3_R1131_U131, P3_R1131_U306, P3_R1131_U307);
  and ginst20177 (P3_R1131_U132, P3_R1131_U309, P3_R1131_U395);
  and ginst20178 (P3_R1131_U133, P3_R1131_U306, P3_R1131_U307);
  and ginst20179 (P3_R1131_U134, P3_R1131_U15, P3_R1131_U310);
  nand ginst20180 (P3_R1131_U135, P3_R1131_U398, P3_R1131_U399);
  and ginst20181 (P3_R1131_U136, P3_R1131_U403, P3_R1131_U404, P3_R1131_U87);
  and ginst20182 (P3_R1131_U137, P3_R1131_U192, P3_R1131_U407);
  nand ginst20183 (P3_R1131_U138, P3_R1131_U412, P3_R1131_U413);
  nand ginst20184 (P3_R1131_U139, P3_R1131_U417, P3_R1131_U418);
  and ginst20185 (P3_R1131_U14, P3_R1131_U195, P3_R1131_U218);
  and ginst20186 (P3_R1131_U140, P3_R1131_U12, P3_R1131_U322);
  and ginst20187 (P3_R1131_U141, P3_R1131_U191, P3_R1131_U424);
  nand ginst20188 (P3_R1131_U142, P3_R1131_U433, P3_R1131_U434);
  nand ginst20189 (P3_R1131_U143, P3_R1131_U438, P3_R1131_U439);
  nand ginst20190 (P3_R1131_U144, P3_R1131_U443, P3_R1131_U444);
  nand ginst20191 (P3_R1131_U145, P3_R1131_U448, P3_R1131_U449);
  nand ginst20192 (P3_R1131_U146, P3_R1131_U453, P3_R1131_U454);
  and ginst20193 (P3_R1131_U147, P3_R1131_U10, P3_R1131_U333);
  and ginst20194 (P3_R1131_U148, P3_R1131_U190, P3_R1131_U460);
  nand ginst20195 (P3_R1131_U149, P3_R1131_U469, P3_R1131_U470);
  and ginst20196 (P3_R1131_U15, P3_R1131_U391, P3_R1131_U392);
  nand ginst20197 (P3_R1131_U150, P3_R1131_U474, P3_R1131_U475);
  and ginst20198 (P3_R1131_U151, P3_R1131_U344, P3_R1131_U8);
  and ginst20199 (P3_R1131_U152, P3_R1131_U189, P3_R1131_U481);
  and ginst20200 (P3_R1131_U153, P3_R1131_U358, P3_R1131_U359);
  nand ginst20201 (P3_R1131_U154, P3_R1131_U120, P3_R1131_U356);
  and ginst20202 (P3_R1131_U155, P3_R1131_U367, P3_R1131_U368);
  and ginst20203 (P3_R1131_U156, P3_R1131_U374, P3_R1131_U375);
  and ginst20204 (P3_R1131_U157, P3_R1131_U378, P3_R1131_U379);
  nand ginst20205 (P3_R1131_U158, P3_R1131_U118, P3_R1131_U203);
  and ginst20206 (P3_R1131_U159, P3_R1131_U387, P3_R1131_U388);
  nand ginst20207 (P3_R1131_U16, P3_R1131_U342, P3_R1131_U345);
  not ginst20208 (P3_R1131_U160, P3_U3908);
  not ginst20209 (P3_R1131_U161, P3_U3054);
  and ginst20210 (P3_R1131_U162, P3_R1131_U396, P3_R1131_U397);
  nand ginst20211 (P3_R1131_U163, P3_R1131_U131, P3_R1131_U304);
  and ginst20212 (P3_R1131_U164, P3_R1131_U408, P3_R1131_U409);
  nand ginst20213 (P3_R1131_U165, P3_R1131_U297, P3_R1131_U298);
  nand ginst20214 (P3_R1131_U166, P3_R1131_U293, P3_R1131_U294);
  and ginst20215 (P3_R1131_U167, P3_R1131_U425, P3_R1131_U426);
  and ginst20216 (P3_R1131_U168, P3_R1131_U429, P3_R1131_U430);
  nand ginst20217 (P3_R1131_U169, P3_R1131_U283, P3_R1131_U284);
  nand ginst20218 (P3_R1131_U17, P3_R1131_U331, P3_R1131_U334);
  nand ginst20219 (P3_R1131_U170, P3_R1131_U279, P3_R1131_U280);
  not ginst20220 (P3_R1131_U171, P3_U3392);
  nand ginst20221 (P3_R1131_U172, P3_R1131_U95, P3_U3387);
  nand ginst20222 (P3_R1131_U173, P3_R1131_U184, P3_R1131_U276, P3_R1131_U350);
  not ginst20223 (P3_R1131_U174, P3_U3443);
  nand ginst20224 (P3_R1131_U175, P3_R1131_U273, P3_R1131_U274);
  nand ginst20225 (P3_R1131_U176, P3_R1131_U269, P3_R1131_U270);
  and ginst20226 (P3_R1131_U177, P3_R1131_U461, P3_R1131_U462);
  and ginst20227 (P3_R1131_U178, P3_R1131_U465, P3_R1131_U466);
  nand ginst20228 (P3_R1131_U179, P3_R1131_U259, P3_R1131_U260);
  nand ginst20229 (P3_R1131_U18, P3_R1131_U320, P3_R1131_U323);
  nand ginst20230 (P3_R1131_U180, P3_R1131_U255, P3_R1131_U256);
  nand ginst20231 (P3_R1131_U181, P3_R1131_U251, P3_R1131_U252);
  and ginst20232 (P3_R1131_U182, P3_R1131_U482, P3_R1131_U483);
  nand ginst20233 (P3_R1131_U183, P3_R1131_U132, P3_R1131_U163);
  nand ginst20234 (P3_R1131_U184, P3_R1131_U174, P3_R1131_U175);
  nand ginst20235 (P3_R1131_U185, P3_R1131_U171, P3_R1131_U172);
  not ginst20236 (P3_R1131_U186, P3_R1131_U87);
  not ginst20237 (P3_R1131_U187, P3_R1131_U34);
  not ginst20238 (P3_R1131_U188, P3_R1131_U26);
  nand ginst20239 (P3_R1131_U189, P3_R1131_U54, P3_U3419);
  nand ginst20240 (P3_R1131_U19, P3_R1131_U312, P3_R1131_U314);
  nand ginst20241 (P3_R1131_U190, P3_R1131_U64, P3_U3434);
  nand ginst20242 (P3_R1131_U191, P3_R1131_U78, P3_U3905);
  nand ginst20243 (P3_R1131_U192, P3_R1131_U86, P3_U3901);
  nand ginst20244 (P3_R1131_U193, P3_R1131_U33, P3_U3395);
  nand ginst20245 (P3_R1131_U194, P3_R1131_U41, P3_U3404);
  nand ginst20246 (P3_R1131_U195, P3_R1131_U25, P3_U3410);
  not ginst20247 (P3_R1131_U196, P3_R1131_U66);
  not ginst20248 (P3_R1131_U197, P3_R1131_U80);
  not ginst20249 (P3_R1131_U198, P3_R1131_U43);
  not ginst20250 (P3_R1131_U199, P3_R1131_U55);
  nand ginst20251 (P3_R1131_U20, P3_R1131_U162, P3_R1131_U183, P3_R1131_U351);
  not ginst20252 (P3_R1131_U200, P3_R1131_U172);
  nand ginst20253 (P3_R1131_U201, P3_R1131_U172, P3_U3077);
  not ginst20254 (P3_R1131_U202, P3_R1131_U49);
  nand ginst20255 (P3_R1131_U203, P3_R1131_U117, P3_R1131_U49);
  nand ginst20256 (P3_R1131_U204, P3_R1131_U34, P3_R1131_U35);
  nand ginst20257 (P3_R1131_U205, P3_R1131_U204, P3_R1131_U32);
  nand ginst20258 (P3_R1131_U206, P3_R1131_U187, P3_U3063);
  not ginst20259 (P3_R1131_U207, P3_R1131_U158);
  nand ginst20260 (P3_R1131_U208, P3_R1131_U40, P3_U3407);
  nand ginst20261 (P3_R1131_U209, P3_R1131_U37, P3_U3070);
  nand ginst20262 (P3_R1131_U21, P3_R1131_U241, P3_R1131_U243);
  nand ginst20263 (P3_R1131_U210, P3_R1131_U36, P3_U3066);
  nand ginst20264 (P3_R1131_U211, P3_R1131_U194, P3_R1131_U198);
  nand ginst20265 (P3_R1131_U212, P3_R1131_U211, P3_R1131_U6);
  nand ginst20266 (P3_R1131_U213, P3_R1131_U42, P3_U3401);
  nand ginst20267 (P3_R1131_U214, P3_R1131_U40, P3_U3407);
  nand ginst20268 (P3_R1131_U215, P3_R1131_U13, P3_R1131_U158);
  not ginst20269 (P3_R1131_U216, P3_R1131_U44);
  not ginst20270 (P3_R1131_U217, P3_R1131_U47);
  nand ginst20271 (P3_R1131_U218, P3_R1131_U27, P3_U3413);
  nand ginst20272 (P3_R1131_U219, P3_R1131_U26, P3_R1131_U27);
  nand ginst20273 (P3_R1131_U22, P3_R1131_U233, P3_R1131_U236);
  nand ginst20274 (P3_R1131_U220, P3_R1131_U188, P3_U3083);
  not ginst20275 (P3_R1131_U221, P3_R1131_U154);
  nand ginst20276 (P3_R1131_U222, P3_R1131_U46, P3_U3416);
  nand ginst20277 (P3_R1131_U223, P3_R1131_U222, P3_R1131_U55);
  nand ginst20278 (P3_R1131_U224, P3_R1131_U217, P3_R1131_U26);
  nand ginst20279 (P3_R1131_U225, P3_R1131_U122, P3_R1131_U224);
  nand ginst20280 (P3_R1131_U226, P3_R1131_U195, P3_R1131_U47);
  nand ginst20281 (P3_R1131_U227, P3_R1131_U121, P3_R1131_U226);
  nand ginst20282 (P3_R1131_U228, P3_R1131_U195, P3_R1131_U26);
  nand ginst20283 (P3_R1131_U229, P3_R1131_U158, P3_R1131_U213);
  nand ginst20284 (P3_R1131_U23, P3_R1131_U225, P3_R1131_U227);
  not ginst20285 (P3_R1131_U230, P3_R1131_U48);
  nand ginst20286 (P3_R1131_U231, P3_R1131_U36, P3_U3066);
  nand ginst20287 (P3_R1131_U232, P3_R1131_U230, P3_R1131_U231);
  nand ginst20288 (P3_R1131_U233, P3_R1131_U124, P3_R1131_U232);
  nand ginst20289 (P3_R1131_U234, P3_R1131_U194, P3_R1131_U48);
  nand ginst20290 (P3_R1131_U235, P3_R1131_U40, P3_U3407);
  nand ginst20291 (P3_R1131_U236, P3_R1131_U123, P3_R1131_U234);
  nand ginst20292 (P3_R1131_U237, P3_R1131_U36, P3_U3066);
  nand ginst20293 (P3_R1131_U238, P3_R1131_U194, P3_R1131_U237);
  nand ginst20294 (P3_R1131_U239, P3_R1131_U213, P3_R1131_U43);
  nand ginst20295 (P3_R1131_U24, P3_R1131_U172, P3_R1131_U348);
  nand ginst20296 (P3_R1131_U240, P3_R1131_U202, P3_R1131_U34);
  nand ginst20297 (P3_R1131_U241, P3_R1131_U126, P3_R1131_U240);
  nand ginst20298 (P3_R1131_U242, P3_R1131_U193, P3_R1131_U49);
  nand ginst20299 (P3_R1131_U243, P3_R1131_U125, P3_R1131_U242);
  nand ginst20300 (P3_R1131_U244, P3_R1131_U193, P3_R1131_U34);
  nand ginst20301 (P3_R1131_U245, P3_R1131_U53, P3_U3422);
  nand ginst20302 (P3_R1131_U246, P3_R1131_U51, P3_U3062);
  nand ginst20303 (P3_R1131_U247, P3_R1131_U52, P3_U3061);
  nand ginst20304 (P3_R1131_U248, P3_R1131_U199, P3_R1131_U7);
  nand ginst20305 (P3_R1131_U249, P3_R1131_U248, P3_R1131_U8);
  not ginst20306 (P3_R1131_U25, P3_U3069);
  nand ginst20307 (P3_R1131_U250, P3_R1131_U53, P3_U3422);
  nand ginst20308 (P3_R1131_U251, P3_R1131_U127, P3_R1131_U154);
  nand ginst20309 (P3_R1131_U252, P3_R1131_U249, P3_R1131_U250);
  not ginst20310 (P3_R1131_U253, P3_R1131_U181);
  nand ginst20311 (P3_R1131_U254, P3_R1131_U57, P3_U3425);
  nand ginst20312 (P3_R1131_U255, P3_R1131_U181, P3_R1131_U254);
  nand ginst20313 (P3_R1131_U256, P3_R1131_U56, P3_U3071);
  not ginst20314 (P3_R1131_U257, P3_R1131_U180);
  nand ginst20315 (P3_R1131_U258, P3_R1131_U59, P3_U3428);
  nand ginst20316 (P3_R1131_U259, P3_R1131_U180, P3_R1131_U258);
  nand ginst20317 (P3_R1131_U26, P3_R1131_U39, P3_U3069);
  nand ginst20318 (P3_R1131_U260, P3_R1131_U58, P3_U3079);
  not ginst20319 (P3_R1131_U261, P3_R1131_U179);
  nand ginst20320 (P3_R1131_U262, P3_R1131_U63, P3_U3437);
  nand ginst20321 (P3_R1131_U263, P3_R1131_U60, P3_U3072);
  nand ginst20322 (P3_R1131_U264, P3_R1131_U61, P3_U3073);
  nand ginst20323 (P3_R1131_U265, P3_R1131_U196, P3_R1131_U9);
  nand ginst20324 (P3_R1131_U266, P3_R1131_U10, P3_R1131_U265);
  nand ginst20325 (P3_R1131_U267, P3_R1131_U65, P3_U3431);
  nand ginst20326 (P3_R1131_U268, P3_R1131_U63, P3_U3437);
  nand ginst20327 (P3_R1131_U269, P3_R1131_U128, P3_R1131_U179);
  not ginst20328 (P3_R1131_U27, P3_U3083);
  nand ginst20329 (P3_R1131_U270, P3_R1131_U266, P3_R1131_U268);
  not ginst20330 (P3_R1131_U271, P3_R1131_U176);
  nand ginst20331 (P3_R1131_U272, P3_R1131_U68, P3_U3440);
  nand ginst20332 (P3_R1131_U273, P3_R1131_U176, P3_R1131_U272);
  nand ginst20333 (P3_R1131_U274, P3_R1131_U67, P3_U3068);
  not ginst20334 (P3_R1131_U275, P3_R1131_U175);
  nand ginst20335 (P3_R1131_U276, P3_R1131_U175, P3_U3081);
  not ginst20336 (P3_R1131_U277, P3_R1131_U173);
  nand ginst20337 (P3_R1131_U278, P3_R1131_U71, P3_U3445);
  nand ginst20338 (P3_R1131_U279, P3_R1131_U173, P3_R1131_U278);
  not ginst20339 (P3_R1131_U28, P3_U3413);
  nand ginst20340 (P3_R1131_U280, P3_R1131_U70, P3_U3080);
  not ginst20341 (P3_R1131_U281, P3_R1131_U170);
  nand ginst20342 (P3_R1131_U282, P3_R1131_U73, P3_U3907);
  nand ginst20343 (P3_R1131_U283, P3_R1131_U170, P3_R1131_U282);
  nand ginst20344 (P3_R1131_U284, P3_R1131_U72, P3_U3075);
  not ginst20345 (P3_R1131_U285, P3_R1131_U169);
  nand ginst20346 (P3_R1131_U286, P3_R1131_U77, P3_U3904);
  nand ginst20347 (P3_R1131_U287, P3_R1131_U74, P3_U3065);
  nand ginst20348 (P3_R1131_U288, P3_R1131_U75, P3_U3060);
  nand ginst20349 (P3_R1131_U289, P3_R1131_U11, P3_R1131_U197);
  not ginst20350 (P3_R1131_U29, P3_U3395);
  nand ginst20351 (P3_R1131_U290, P3_R1131_U12, P3_R1131_U289);
  nand ginst20352 (P3_R1131_U291, P3_R1131_U79, P3_U3906);
  nand ginst20353 (P3_R1131_U292, P3_R1131_U77, P3_U3904);
  nand ginst20354 (P3_R1131_U293, P3_R1131_U129, P3_R1131_U169);
  nand ginst20355 (P3_R1131_U294, P3_R1131_U290, P3_R1131_U292);
  not ginst20356 (P3_R1131_U295, P3_R1131_U166);
  nand ginst20357 (P3_R1131_U296, P3_R1131_U82, P3_U3903);
  nand ginst20358 (P3_R1131_U297, P3_R1131_U166, P3_R1131_U296);
  nand ginst20359 (P3_R1131_U298, P3_R1131_U81, P3_U3064);
  not ginst20360 (P3_R1131_U299, P3_R1131_U165);
  not ginst20361 (P3_R1131_U30, P3_U3387);
  nand ginst20362 (P3_R1131_U300, P3_R1131_U84, P3_U3902);
  nand ginst20363 (P3_R1131_U301, P3_R1131_U165, P3_R1131_U300);
  nand ginst20364 (P3_R1131_U302, P3_R1131_U83, P3_U3057);
  not ginst20365 (P3_R1131_U303, P3_R1131_U91);
  nand ginst20366 (P3_R1131_U304, P3_R1131_U130, P3_R1131_U91);
  nand ginst20367 (P3_R1131_U305, P3_R1131_U87, P3_R1131_U88);
  nand ginst20368 (P3_R1131_U306, P3_R1131_U305, P3_R1131_U85);
  nand ginst20369 (P3_R1131_U307, P3_R1131_U186, P3_U3052);
  not ginst20370 (P3_R1131_U308, P3_R1131_U163);
  nand ginst20371 (P3_R1131_U309, P3_R1131_U90, P3_U3899);
  not ginst20372 (P3_R1131_U31, P3_U3077);
  nand ginst20373 (P3_R1131_U310, P3_R1131_U89, P3_U3053);
  nand ginst20374 (P3_R1131_U311, P3_R1131_U303, P3_R1131_U87);
  nand ginst20375 (P3_R1131_U312, P3_R1131_U137, P3_R1131_U311);
  nand ginst20376 (P3_R1131_U313, P3_R1131_U192, P3_R1131_U91);
  nand ginst20377 (P3_R1131_U314, P3_R1131_U136, P3_R1131_U313);
  nand ginst20378 (P3_R1131_U315, P3_R1131_U192, P3_R1131_U87);
  nand ginst20379 (P3_R1131_U316, P3_R1131_U169, P3_R1131_U291);
  not ginst20380 (P3_R1131_U317, P3_R1131_U92);
  nand ginst20381 (P3_R1131_U318, P3_R1131_U75, P3_U3060);
  nand ginst20382 (P3_R1131_U319, P3_R1131_U317, P3_R1131_U318);
  not ginst20383 (P3_R1131_U32, P3_U3398);
  nand ginst20384 (P3_R1131_U320, P3_R1131_U141, P3_R1131_U319);
  nand ginst20385 (P3_R1131_U321, P3_R1131_U191, P3_R1131_U92);
  nand ginst20386 (P3_R1131_U322, P3_R1131_U77, P3_U3904);
  nand ginst20387 (P3_R1131_U323, P3_R1131_U140, P3_R1131_U321);
  nand ginst20388 (P3_R1131_U324, P3_R1131_U75, P3_U3060);
  nand ginst20389 (P3_R1131_U325, P3_R1131_U191, P3_R1131_U324);
  nand ginst20390 (P3_R1131_U326, P3_R1131_U291, P3_R1131_U80);
  nand ginst20391 (P3_R1131_U327, P3_R1131_U179, P3_R1131_U267);
  not ginst20392 (P3_R1131_U328, P3_R1131_U93);
  nand ginst20393 (P3_R1131_U329, P3_R1131_U61, P3_U3073);
  not ginst20394 (P3_R1131_U33, P3_U3067);
  nand ginst20395 (P3_R1131_U330, P3_R1131_U328, P3_R1131_U329);
  nand ginst20396 (P3_R1131_U331, P3_R1131_U148, P3_R1131_U330);
  nand ginst20397 (P3_R1131_U332, P3_R1131_U190, P3_R1131_U93);
  nand ginst20398 (P3_R1131_U333, P3_R1131_U63, P3_U3437);
  nand ginst20399 (P3_R1131_U334, P3_R1131_U147, P3_R1131_U332);
  nand ginst20400 (P3_R1131_U335, P3_R1131_U61, P3_U3073);
  nand ginst20401 (P3_R1131_U336, P3_R1131_U190, P3_R1131_U335);
  nand ginst20402 (P3_R1131_U337, P3_R1131_U267, P3_R1131_U66);
  nand ginst20403 (P3_R1131_U338, P3_R1131_U154, P3_R1131_U222);
  not ginst20404 (P3_R1131_U339, P3_R1131_U94);
  nand ginst20405 (P3_R1131_U34, P3_R1131_U29, P3_U3067);
  nand ginst20406 (P3_R1131_U340, P3_R1131_U52, P3_U3061);
  nand ginst20407 (P3_R1131_U341, P3_R1131_U339, P3_R1131_U340);
  nand ginst20408 (P3_R1131_U342, P3_R1131_U152, P3_R1131_U341);
  nand ginst20409 (P3_R1131_U343, P3_R1131_U189, P3_R1131_U94);
  nand ginst20410 (P3_R1131_U344, P3_R1131_U53, P3_U3422);
  nand ginst20411 (P3_R1131_U345, P3_R1131_U151, P3_R1131_U343);
  nand ginst20412 (P3_R1131_U346, P3_R1131_U52, P3_U3061);
  nand ginst20413 (P3_R1131_U347, P3_R1131_U189, P3_R1131_U346);
  nand ginst20414 (P3_R1131_U348, P3_R1131_U30, P3_U3076);
  nand ginst20415 (P3_R1131_U349, P3_R1131_U171, P3_U3077);
  not ginst20416 (P3_R1131_U35, P3_U3063);
  nand ginst20417 (P3_R1131_U350, P3_R1131_U174, P3_U3081);
  nand ginst20418 (P3_R1131_U351, P3_R1131_U133, P3_R1131_U134, P3_R1131_U304);
  nand ginst20419 (P3_R1131_U352, P3_R1131_U35, P3_U3398);
  nand ginst20420 (P3_R1131_U353, P3_R1131_U220, P3_U3413);
  nand ginst20421 (P3_R1131_U354, P3_R1131_U219, P3_R1131_U353);
  nand ginst20422 (P3_R1131_U355, P3_R1131_U88, P3_U3900);
  nand ginst20423 (P3_R1131_U356, P3_R1131_U119, P3_R1131_U158);
  nand ginst20424 (P3_R1131_U357, P3_R1131_U14, P3_R1131_U216);
  nand ginst20425 (P3_R1131_U358, P3_R1131_U46, P3_U3416);
  nand ginst20426 (P3_R1131_U359, P3_R1131_U45, P3_U3082);
  not ginst20427 (P3_R1131_U36, P3_U3404);
  nand ginst20428 (P3_R1131_U360, P3_R1131_U154, P3_R1131_U223);
  nand ginst20429 (P3_R1131_U361, P3_R1131_U153, P3_R1131_U221);
  nand ginst20430 (P3_R1131_U362, P3_R1131_U27, P3_U3413);
  nand ginst20431 (P3_R1131_U363, P3_R1131_U28, P3_U3083);
  nand ginst20432 (P3_R1131_U364, P3_R1131_U27, P3_U3413);
  nand ginst20433 (P3_R1131_U365, P3_R1131_U28, P3_U3083);
  nand ginst20434 (P3_R1131_U366, P3_R1131_U364, P3_R1131_U365);
  nand ginst20435 (P3_R1131_U367, P3_R1131_U25, P3_U3410);
  nand ginst20436 (P3_R1131_U368, P3_R1131_U39, P3_U3069);
  nand ginst20437 (P3_R1131_U369, P3_R1131_U228, P3_R1131_U47);
  not ginst20438 (P3_R1131_U37, P3_U3407);
  nand ginst20439 (P3_R1131_U370, P3_R1131_U155, P3_R1131_U217);
  nand ginst20440 (P3_R1131_U371, P3_R1131_U40, P3_U3407);
  nand ginst20441 (P3_R1131_U372, P3_R1131_U37, P3_U3070);
  nand ginst20442 (P3_R1131_U373, P3_R1131_U371, P3_R1131_U372);
  nand ginst20443 (P3_R1131_U374, P3_R1131_U41, P3_U3404);
  nand ginst20444 (P3_R1131_U375, P3_R1131_U36, P3_U3066);
  nand ginst20445 (P3_R1131_U376, P3_R1131_U238, P3_R1131_U48);
  nand ginst20446 (P3_R1131_U377, P3_R1131_U156, P3_R1131_U230);
  nand ginst20447 (P3_R1131_U378, P3_R1131_U42, P3_U3401);
  nand ginst20448 (P3_R1131_U379, P3_R1131_U38, P3_U3059);
  not ginst20449 (P3_R1131_U38, P3_U3401);
  nand ginst20450 (P3_R1131_U380, P3_R1131_U158, P3_R1131_U239);
  nand ginst20451 (P3_R1131_U381, P3_R1131_U157, P3_R1131_U207);
  nand ginst20452 (P3_R1131_U382, P3_R1131_U35, P3_U3398);
  nand ginst20453 (P3_R1131_U383, P3_R1131_U32, P3_U3063);
  nand ginst20454 (P3_R1131_U384, P3_R1131_U35, P3_U3398);
  nand ginst20455 (P3_R1131_U385, P3_R1131_U32, P3_U3063);
  nand ginst20456 (P3_R1131_U386, P3_R1131_U384, P3_R1131_U385);
  nand ginst20457 (P3_R1131_U387, P3_R1131_U33, P3_U3395);
  nand ginst20458 (P3_R1131_U388, P3_R1131_U29, P3_U3067);
  nand ginst20459 (P3_R1131_U389, P3_R1131_U244, P3_R1131_U49);
  not ginst20460 (P3_R1131_U39, P3_U3410);
  nand ginst20461 (P3_R1131_U390, P3_R1131_U159, P3_R1131_U202);
  nand ginst20462 (P3_R1131_U391, P3_R1131_U161, P3_U3908);
  nand ginst20463 (P3_R1131_U392, P3_R1131_U160, P3_U3054);
  nand ginst20464 (P3_R1131_U393, P3_R1131_U161, P3_U3908);
  nand ginst20465 (P3_R1131_U394, P3_R1131_U160, P3_U3054);
  nand ginst20466 (P3_R1131_U395, P3_R1131_U393, P3_R1131_U394);
  nand ginst20467 (P3_R1131_U396, P3_R1131_U395, P3_R1131_U89, P3_U3053);
  nand ginst20468 (P3_R1131_U397, P3_R1131_U15, P3_R1131_U90, P3_U3899);
  nand ginst20469 (P3_R1131_U398, P3_R1131_U90, P3_U3899);
  nand ginst20470 (P3_R1131_U399, P3_R1131_U89, P3_U3053);
  not ginst20471 (P3_R1131_U40, P3_U3070);
  not ginst20472 (P3_R1131_U400, P3_R1131_U135);
  nand ginst20473 (P3_R1131_U401, P3_R1131_U308, P3_R1131_U400);
  nand ginst20474 (P3_R1131_U402, P3_R1131_U135, P3_R1131_U163);
  nand ginst20475 (P3_R1131_U403, P3_R1131_U88, P3_U3900);
  nand ginst20476 (P3_R1131_U404, P3_R1131_U85, P3_U3052);
  nand ginst20477 (P3_R1131_U405, P3_R1131_U88, P3_U3900);
  nand ginst20478 (P3_R1131_U406, P3_R1131_U85, P3_U3052);
  nand ginst20479 (P3_R1131_U407, P3_R1131_U405, P3_R1131_U406);
  nand ginst20480 (P3_R1131_U408, P3_R1131_U86, P3_U3901);
  nand ginst20481 (P3_R1131_U409, P3_R1131_U50, P3_U3056);
  not ginst20482 (P3_R1131_U41, P3_U3066);
  nand ginst20483 (P3_R1131_U410, P3_R1131_U315, P3_R1131_U91);
  nand ginst20484 (P3_R1131_U411, P3_R1131_U164, P3_R1131_U303);
  nand ginst20485 (P3_R1131_U412, P3_R1131_U84, P3_U3902);
  nand ginst20486 (P3_R1131_U413, P3_R1131_U83, P3_U3057);
  not ginst20487 (P3_R1131_U414, P3_R1131_U138);
  nand ginst20488 (P3_R1131_U415, P3_R1131_U299, P3_R1131_U414);
  nand ginst20489 (P3_R1131_U416, P3_R1131_U138, P3_R1131_U165);
  nand ginst20490 (P3_R1131_U417, P3_R1131_U82, P3_U3903);
  nand ginst20491 (P3_R1131_U418, P3_R1131_U81, P3_U3064);
  not ginst20492 (P3_R1131_U419, P3_R1131_U139);
  not ginst20493 (P3_R1131_U42, P3_U3059);
  nand ginst20494 (P3_R1131_U420, P3_R1131_U295, P3_R1131_U419);
  nand ginst20495 (P3_R1131_U421, P3_R1131_U139, P3_R1131_U166);
  nand ginst20496 (P3_R1131_U422, P3_R1131_U77, P3_U3904);
  nand ginst20497 (P3_R1131_U423, P3_R1131_U74, P3_U3065);
  nand ginst20498 (P3_R1131_U424, P3_R1131_U422, P3_R1131_U423);
  nand ginst20499 (P3_R1131_U425, P3_R1131_U78, P3_U3905);
  nand ginst20500 (P3_R1131_U426, P3_R1131_U75, P3_U3060);
  nand ginst20501 (P3_R1131_U427, P3_R1131_U325, P3_R1131_U92);
  nand ginst20502 (P3_R1131_U428, P3_R1131_U167, P3_R1131_U317);
  nand ginst20503 (P3_R1131_U429, P3_R1131_U79, P3_U3906);
  nand ginst20504 (P3_R1131_U43, P3_R1131_U38, P3_U3059);
  nand ginst20505 (P3_R1131_U430, P3_R1131_U76, P3_U3074);
  nand ginst20506 (P3_R1131_U431, P3_R1131_U169, P3_R1131_U326);
  nand ginst20507 (P3_R1131_U432, P3_R1131_U168, P3_R1131_U285);
  nand ginst20508 (P3_R1131_U433, P3_R1131_U73, P3_U3907);
  nand ginst20509 (P3_R1131_U434, P3_R1131_U72, P3_U3075);
  not ginst20510 (P3_R1131_U435, P3_R1131_U142);
  nand ginst20511 (P3_R1131_U436, P3_R1131_U281, P3_R1131_U435);
  nand ginst20512 (P3_R1131_U437, P3_R1131_U142, P3_R1131_U170);
  nand ginst20513 (P3_R1131_U438, P3_R1131_U31, P3_U3392);
  nand ginst20514 (P3_R1131_U439, P3_R1131_U171, P3_U3077);
  nand ginst20515 (P3_R1131_U44, P3_R1131_U212, P3_R1131_U214);
  not ginst20516 (P3_R1131_U440, P3_R1131_U143);
  nand ginst20517 (P3_R1131_U441, P3_R1131_U200, P3_R1131_U440);
  nand ginst20518 (P3_R1131_U442, P3_R1131_U143, P3_R1131_U172);
  nand ginst20519 (P3_R1131_U443, P3_R1131_U71, P3_U3445);
  nand ginst20520 (P3_R1131_U444, P3_R1131_U70, P3_U3080);
  not ginst20521 (P3_R1131_U445, P3_R1131_U144);
  nand ginst20522 (P3_R1131_U446, P3_R1131_U277, P3_R1131_U445);
  nand ginst20523 (P3_R1131_U447, P3_R1131_U144, P3_R1131_U173);
  nand ginst20524 (P3_R1131_U448, P3_R1131_U69, P3_U3443);
  nand ginst20525 (P3_R1131_U449, P3_R1131_U174, P3_U3081);
  not ginst20526 (P3_R1131_U45, P3_U3416);
  not ginst20527 (P3_R1131_U450, P3_R1131_U145);
  nand ginst20528 (P3_R1131_U451, P3_R1131_U275, P3_R1131_U450);
  nand ginst20529 (P3_R1131_U452, P3_R1131_U145, P3_R1131_U175);
  nand ginst20530 (P3_R1131_U453, P3_R1131_U68, P3_U3440);
  nand ginst20531 (P3_R1131_U454, P3_R1131_U67, P3_U3068);
  not ginst20532 (P3_R1131_U455, P3_R1131_U146);
  nand ginst20533 (P3_R1131_U456, P3_R1131_U271, P3_R1131_U455);
  nand ginst20534 (P3_R1131_U457, P3_R1131_U146, P3_R1131_U176);
  nand ginst20535 (P3_R1131_U458, P3_R1131_U63, P3_U3437);
  nand ginst20536 (P3_R1131_U459, P3_R1131_U60, P3_U3072);
  not ginst20537 (P3_R1131_U46, P3_U3082);
  nand ginst20538 (P3_R1131_U460, P3_R1131_U458, P3_R1131_U459);
  nand ginst20539 (P3_R1131_U461, P3_R1131_U64, P3_U3434);
  nand ginst20540 (P3_R1131_U462, P3_R1131_U61, P3_U3073);
  nand ginst20541 (P3_R1131_U463, P3_R1131_U336, P3_R1131_U93);
  nand ginst20542 (P3_R1131_U464, P3_R1131_U177, P3_R1131_U328);
  nand ginst20543 (P3_R1131_U465, P3_R1131_U65, P3_U3431);
  nand ginst20544 (P3_R1131_U466, P3_R1131_U62, P3_U3078);
  nand ginst20545 (P3_R1131_U467, P3_R1131_U179, P3_R1131_U337);
  nand ginst20546 (P3_R1131_U468, P3_R1131_U178, P3_R1131_U261);
  nand ginst20547 (P3_R1131_U469, P3_R1131_U59, P3_U3428);
  nand ginst20548 (P3_R1131_U47, P3_R1131_U215, P3_R1131_U44);
  nand ginst20549 (P3_R1131_U470, P3_R1131_U58, P3_U3079);
  not ginst20550 (P3_R1131_U471, P3_R1131_U149);
  nand ginst20551 (P3_R1131_U472, P3_R1131_U257, P3_R1131_U471);
  nand ginst20552 (P3_R1131_U473, P3_R1131_U149, P3_R1131_U180);
  nand ginst20553 (P3_R1131_U474, P3_R1131_U57, P3_U3425);
  nand ginst20554 (P3_R1131_U475, P3_R1131_U56, P3_U3071);
  not ginst20555 (P3_R1131_U476, P3_R1131_U150);
  nand ginst20556 (P3_R1131_U477, P3_R1131_U253, P3_R1131_U476);
  nand ginst20557 (P3_R1131_U478, P3_R1131_U150, P3_R1131_U181);
  nand ginst20558 (P3_R1131_U479, P3_R1131_U53, P3_U3422);
  nand ginst20559 (P3_R1131_U48, P3_R1131_U229, P3_R1131_U43);
  nand ginst20560 (P3_R1131_U480, P3_R1131_U51, P3_U3062);
  nand ginst20561 (P3_R1131_U481, P3_R1131_U479, P3_R1131_U480);
  nand ginst20562 (P3_R1131_U482, P3_R1131_U54, P3_U3419);
  nand ginst20563 (P3_R1131_U483, P3_R1131_U52, P3_U3061);
  nand ginst20564 (P3_R1131_U484, P3_R1131_U347, P3_R1131_U94);
  nand ginst20565 (P3_R1131_U485, P3_R1131_U182, P3_R1131_U339);
  nand ginst20566 (P3_R1131_U49, P3_R1131_U185, P3_R1131_U201, P3_R1131_U349);
  not ginst20567 (P3_R1131_U50, P3_U3901);
  not ginst20568 (P3_R1131_U51, P3_U3422);
  not ginst20569 (P3_R1131_U52, P3_U3419);
  not ginst20570 (P3_R1131_U53, P3_U3062);
  not ginst20571 (P3_R1131_U54, P3_U3061);
  nand ginst20572 (P3_R1131_U55, P3_R1131_U45, P3_U3082);
  not ginst20573 (P3_R1131_U56, P3_U3425);
  not ginst20574 (P3_R1131_U57, P3_U3071);
  not ginst20575 (P3_R1131_U58, P3_U3428);
  not ginst20576 (P3_R1131_U59, P3_U3079);
  and ginst20577 (P3_R1131_U6, P3_R1131_U209, P3_R1131_U210);
  not ginst20578 (P3_R1131_U60, P3_U3437);
  not ginst20579 (P3_R1131_U61, P3_U3434);
  not ginst20580 (P3_R1131_U62, P3_U3431);
  not ginst20581 (P3_R1131_U63, P3_U3072);
  not ginst20582 (P3_R1131_U64, P3_U3073);
  not ginst20583 (P3_R1131_U65, P3_U3078);
  nand ginst20584 (P3_R1131_U66, P3_R1131_U62, P3_U3078);
  not ginst20585 (P3_R1131_U67, P3_U3440);
  not ginst20586 (P3_R1131_U68, P3_U3068);
  not ginst20587 (P3_R1131_U69, P3_U3081);
  and ginst20588 (P3_R1131_U7, P3_R1131_U189, P3_R1131_U245);
  not ginst20589 (P3_R1131_U70, P3_U3445);
  not ginst20590 (P3_R1131_U71, P3_U3080);
  not ginst20591 (P3_R1131_U72, P3_U3907);
  not ginst20592 (P3_R1131_U73, P3_U3075);
  not ginst20593 (P3_R1131_U74, P3_U3904);
  not ginst20594 (P3_R1131_U75, P3_U3905);
  not ginst20595 (P3_R1131_U76, P3_U3906);
  not ginst20596 (P3_R1131_U77, P3_U3065);
  not ginst20597 (P3_R1131_U78, P3_U3060);
  not ginst20598 (P3_R1131_U79, P3_U3074);
  and ginst20599 (P3_R1131_U8, P3_R1131_U246, P3_R1131_U247);
  nand ginst20600 (P3_R1131_U80, P3_R1131_U76, P3_U3074);
  not ginst20601 (P3_R1131_U81, P3_U3903);
  not ginst20602 (P3_R1131_U82, P3_U3064);
  not ginst20603 (P3_R1131_U83, P3_U3902);
  not ginst20604 (P3_R1131_U84, P3_U3057);
  not ginst20605 (P3_R1131_U85, P3_U3900);
  not ginst20606 (P3_R1131_U86, P3_U3056);
  nand ginst20607 (P3_R1131_U87, P3_R1131_U50, P3_U3056);
  not ginst20608 (P3_R1131_U88, P3_U3052);
  not ginst20609 (P3_R1131_U89, P3_U3899);
  and ginst20610 (P3_R1131_U9, P3_R1131_U190, P3_R1131_U262);
  not ginst20611 (P3_R1131_U90, P3_U3053);
  nand ginst20612 (P3_R1131_U91, P3_R1131_U301, P3_R1131_U302);
  nand ginst20613 (P3_R1131_U92, P3_R1131_U316, P3_R1131_U80);
  nand ginst20614 (P3_R1131_U93, P3_R1131_U327, P3_R1131_U66);
  nand ginst20615 (P3_R1131_U94, P3_R1131_U338, P3_R1131_U55);
  not ginst20616 (P3_R1131_U95, P3_U3076);
  nand ginst20617 (P3_R1131_U96, P3_R1131_U401, P3_R1131_U402);
  nand ginst20618 (P3_R1131_U97, P3_R1131_U415, P3_R1131_U416);
  nand ginst20619 (P3_R1131_U98, P3_R1131_U420, P3_R1131_U421);
  nand ginst20620 (P3_R1131_U99, P3_R1131_U436, P3_R1131_U437);
  and ginst20621 (P3_R1143_U10, P3_R1143_U348, P3_R1143_U351);
  nand ginst20622 (P3_R1143_U100, P3_R1143_U398, P3_R1143_U399);
  nand ginst20623 (P3_R1143_U101, P3_R1143_U407, P3_R1143_U408);
  nand ginst20624 (P3_R1143_U102, P3_R1143_U414, P3_R1143_U415);
  nand ginst20625 (P3_R1143_U103, P3_R1143_U421, P3_R1143_U422);
  nand ginst20626 (P3_R1143_U104, P3_R1143_U428, P3_R1143_U429);
  nand ginst20627 (P3_R1143_U105, P3_R1143_U433, P3_R1143_U434);
  nand ginst20628 (P3_R1143_U106, P3_R1143_U440, P3_R1143_U441);
  nand ginst20629 (P3_R1143_U107, P3_R1143_U447, P3_R1143_U448);
  nand ginst20630 (P3_R1143_U108, P3_R1143_U461, P3_R1143_U462);
  nand ginst20631 (P3_R1143_U109, P3_R1143_U466, P3_R1143_U467);
  and ginst20632 (P3_R1143_U11, P3_R1143_U341, P3_R1143_U344);
  nand ginst20633 (P3_R1143_U110, P3_R1143_U473, P3_R1143_U474);
  nand ginst20634 (P3_R1143_U111, P3_R1143_U480, P3_R1143_U481);
  nand ginst20635 (P3_R1143_U112, P3_R1143_U487, P3_R1143_U488);
  nand ginst20636 (P3_R1143_U113, P3_R1143_U494, P3_R1143_U495);
  nand ginst20637 (P3_R1143_U114, P3_R1143_U499, P3_R1143_U500);
  and ginst20638 (P3_R1143_U115, P3_R1143_U187, P3_R1143_U189);
  and ginst20639 (P3_R1143_U116, P3_R1143_U180, P3_R1143_U4);
  and ginst20640 (P3_R1143_U117, P3_R1143_U192, P3_R1143_U194);
  and ginst20641 (P3_R1143_U118, P3_R1143_U200, P3_R1143_U201);
  and ginst20642 (P3_R1143_U119, P3_R1143_U22, P3_R1143_U381, P3_R1143_U382);
  and ginst20643 (P3_R1143_U12, P3_R1143_U332, P3_R1143_U335);
  and ginst20644 (P3_R1143_U120, P3_R1143_U212, P3_R1143_U5);
  and ginst20645 (P3_R1143_U121, P3_R1143_U180, P3_R1143_U181);
  and ginst20646 (P3_R1143_U122, P3_R1143_U218, P3_R1143_U220);
  and ginst20647 (P3_R1143_U123, P3_R1143_U34, P3_R1143_U388, P3_R1143_U389);
  and ginst20648 (P3_R1143_U124, P3_R1143_U226, P3_R1143_U4);
  and ginst20649 (P3_R1143_U125, P3_R1143_U181, P3_R1143_U234);
  and ginst20650 (P3_R1143_U126, P3_R1143_U204, P3_R1143_U6);
  and ginst20651 (P3_R1143_U127, P3_R1143_U239, P3_R1143_U243);
  and ginst20652 (P3_R1143_U128, P3_R1143_U250, P3_R1143_U7);
  and ginst20653 (P3_R1143_U129, P3_R1143_U172, P3_R1143_U248);
  and ginst20654 (P3_R1143_U13, P3_R1143_U323, P3_R1143_U326);
  and ginst20655 (P3_R1143_U130, P3_R1143_U267, P3_R1143_U268);
  and ginst20656 (P3_R1143_U131, P3_R1143_U273, P3_R1143_U282, P3_R1143_U9);
  and ginst20657 (P3_R1143_U132, P3_R1143_U280, P3_R1143_U285);
  and ginst20658 (P3_R1143_U133, P3_R1143_U298, P3_R1143_U301);
  and ginst20659 (P3_R1143_U134, P3_R1143_U302, P3_R1143_U368);
  and ginst20660 (P3_R1143_U135, P3_R1143_U160, P3_R1143_U278);
  and ginst20661 (P3_R1143_U136, P3_R1143_U454, P3_R1143_U455, P3_R1143_U80);
  and ginst20662 (P3_R1143_U137, P3_R1143_U325, P3_R1143_U9);
  and ginst20663 (P3_R1143_U138, P3_R1143_U468, P3_R1143_U469, P3_R1143_U59);
  and ginst20664 (P3_R1143_U139, P3_R1143_U334, P3_R1143_U8);
  and ginst20665 (P3_R1143_U14, P3_R1143_U318, P3_R1143_U320);
  and ginst20666 (P3_R1143_U140, P3_R1143_U172, P3_R1143_U489, P3_R1143_U490);
  and ginst20667 (P3_R1143_U141, P3_R1143_U343, P3_R1143_U7);
  and ginst20668 (P3_R1143_U142, P3_R1143_U171, P3_R1143_U501, P3_R1143_U502);
  and ginst20669 (P3_R1143_U143, P3_R1143_U350, P3_R1143_U6);
  nand ginst20670 (P3_R1143_U144, P3_R1143_U118, P3_R1143_U202);
  nand ginst20671 (P3_R1143_U145, P3_R1143_U217, P3_R1143_U229);
  not ginst20672 (P3_R1143_U146, P3_U3054);
  not ginst20673 (P3_R1143_U147, P3_U3908);
  and ginst20674 (P3_R1143_U148, P3_R1143_U402, P3_R1143_U403);
  nand ginst20675 (P3_R1143_U149, P3_R1143_U169, P3_R1143_U304, P3_R1143_U364);
  and ginst20676 (P3_R1143_U15, P3_R1143_U310, P3_R1143_U313);
  and ginst20677 (P3_R1143_U150, P3_R1143_U409, P3_R1143_U410);
  nand ginst20678 (P3_R1143_U151, P3_R1143_U134, P3_R1143_U369, P3_R1143_U370);
  and ginst20679 (P3_R1143_U152, P3_R1143_U416, P3_R1143_U417);
  nand ginst20680 (P3_R1143_U153, P3_R1143_U299, P3_R1143_U365, P3_R1143_U86);
  and ginst20681 (P3_R1143_U154, P3_R1143_U423, P3_R1143_U424);
  nand ginst20682 (P3_R1143_U155, P3_R1143_U292, P3_R1143_U293);
  and ginst20683 (P3_R1143_U156, P3_R1143_U435, P3_R1143_U436);
  nand ginst20684 (P3_R1143_U157, P3_R1143_U288, P3_R1143_U289);
  and ginst20685 (P3_R1143_U158, P3_R1143_U442, P3_R1143_U443);
  nand ginst20686 (P3_R1143_U159, P3_R1143_U132, P3_R1143_U284);
  and ginst20687 (P3_R1143_U16, P3_R1143_U232, P3_R1143_U235);
  and ginst20688 (P3_R1143_U160, P3_R1143_U449, P3_R1143_U450);
  nand ginst20689 (P3_R1143_U161, P3_R1143_U327, P3_R1143_U43);
  nand ginst20690 (P3_R1143_U162, P3_R1143_U130, P3_R1143_U269);
  and ginst20691 (P3_R1143_U163, P3_R1143_U475, P3_R1143_U476);
  nand ginst20692 (P3_R1143_U164, P3_R1143_U256, P3_R1143_U257);
  and ginst20693 (P3_R1143_U165, P3_R1143_U482, P3_R1143_U483);
  nand ginst20694 (P3_R1143_U166, P3_R1143_U252, P3_R1143_U253);
  nand ginst20695 (P3_R1143_U167, P3_R1143_U127, P3_R1143_U242);
  nand ginst20696 (P3_R1143_U168, P3_R1143_U366, P3_R1143_U367);
  nand ginst20697 (P3_R1143_U169, P3_R1143_U151, P3_U3053);
  and ginst20698 (P3_R1143_U17, P3_R1143_U224, P3_R1143_U227);
  not ginst20699 (P3_R1143_U170, P3_R1143_U34);
  nand ginst20700 (P3_R1143_U171, P3_U3082, P3_U3416);
  nand ginst20701 (P3_R1143_U172, P3_U3071, P3_U3425);
  nand ginst20702 (P3_R1143_U173, P3_U3057, P3_U3902);
  not ginst20703 (P3_R1143_U174, P3_R1143_U68);
  not ginst20704 (P3_R1143_U175, P3_R1143_U77);
  nand ginst20705 (P3_R1143_U176, P3_U3064, P3_U3903);
  not ginst20706 (P3_R1143_U177, P3_R1143_U63);
  or ginst20707 (P3_R1143_U178, P3_U3066, P3_U3404);
  or ginst20708 (P3_R1143_U179, P3_U3059, P3_U3401);
  and ginst20709 (P3_R1143_U18, P3_R1143_U210, P3_R1143_U213);
  or ginst20710 (P3_R1143_U180, P3_U3063, P3_U3398);
  or ginst20711 (P3_R1143_U181, P3_U3067, P3_U3395);
  not ginst20712 (P3_R1143_U182, P3_R1143_U31);
  or ginst20713 (P3_R1143_U183, P3_U3077, P3_U3392);
  not ginst20714 (P3_R1143_U184, P3_R1143_U42);
  not ginst20715 (P3_R1143_U185, P3_R1143_U43);
  nand ginst20716 (P3_R1143_U186, P3_R1143_U42, P3_R1143_U43);
  nand ginst20717 (P3_R1143_U187, P3_U3067, P3_U3395);
  nand ginst20718 (P3_R1143_U188, P3_R1143_U181, P3_R1143_U186);
  nand ginst20719 (P3_R1143_U189, P3_U3063, P3_U3398);
  not ginst20720 (P3_R1143_U19, P3_U3407);
  nand ginst20721 (P3_R1143_U190, P3_R1143_U115, P3_R1143_U188);
  nand ginst20722 (P3_R1143_U191, P3_R1143_U34, P3_R1143_U35);
  nand ginst20723 (P3_R1143_U192, P3_R1143_U191, P3_U3066);
  nand ginst20724 (P3_R1143_U193, P3_R1143_U116, P3_R1143_U190);
  nand ginst20725 (P3_R1143_U194, P3_R1143_U170, P3_U3404);
  not ginst20726 (P3_R1143_U195, P3_R1143_U41);
  or ginst20727 (P3_R1143_U196, P3_U3069, P3_U3410);
  or ginst20728 (P3_R1143_U197, P3_U3070, P3_U3407);
  not ginst20729 (P3_R1143_U198, P3_R1143_U22);
  nand ginst20730 (P3_R1143_U199, P3_R1143_U22, P3_R1143_U23);
  not ginst20731 (P3_R1143_U20, P3_U3070);
  nand ginst20732 (P3_R1143_U200, P3_R1143_U199, P3_U3069);
  nand ginst20733 (P3_R1143_U201, P3_R1143_U198, P3_U3410);
  nand ginst20734 (P3_R1143_U202, P3_R1143_U41, P3_R1143_U5);
  not ginst20735 (P3_R1143_U203, P3_R1143_U144);
  or ginst20736 (P3_R1143_U204, P3_U3083, P3_U3413);
  nand ginst20737 (P3_R1143_U205, P3_R1143_U144, P3_R1143_U204);
  not ginst20738 (P3_R1143_U206, P3_R1143_U40);
  or ginst20739 (P3_R1143_U207, P3_U3082, P3_U3416);
  or ginst20740 (P3_R1143_U208, P3_U3070, P3_U3407);
  nand ginst20741 (P3_R1143_U209, P3_R1143_U208, P3_R1143_U41);
  not ginst20742 (P3_R1143_U21, P3_U3069);
  nand ginst20743 (P3_R1143_U210, P3_R1143_U119, P3_R1143_U209);
  nand ginst20744 (P3_R1143_U211, P3_R1143_U195, P3_R1143_U22);
  nand ginst20745 (P3_R1143_U212, P3_U3069, P3_U3410);
  nand ginst20746 (P3_R1143_U213, P3_R1143_U120, P3_R1143_U211);
  or ginst20747 (P3_R1143_U214, P3_U3070, P3_U3407);
  nand ginst20748 (P3_R1143_U215, P3_R1143_U181, P3_R1143_U185);
  nand ginst20749 (P3_R1143_U216, P3_U3067, P3_U3395);
  not ginst20750 (P3_R1143_U217, P3_R1143_U45);
  nand ginst20751 (P3_R1143_U218, P3_R1143_U121, P3_R1143_U184);
  nand ginst20752 (P3_R1143_U219, P3_R1143_U180, P3_R1143_U45);
  nand ginst20753 (P3_R1143_U22, P3_U3070, P3_U3407);
  nand ginst20754 (P3_R1143_U220, P3_U3063, P3_U3398);
  not ginst20755 (P3_R1143_U221, P3_R1143_U44);
  or ginst20756 (P3_R1143_U222, P3_U3059, P3_U3401);
  nand ginst20757 (P3_R1143_U223, P3_R1143_U222, P3_R1143_U44);
  nand ginst20758 (P3_R1143_U224, P3_R1143_U123, P3_R1143_U223);
  nand ginst20759 (P3_R1143_U225, P3_R1143_U221, P3_R1143_U34);
  nand ginst20760 (P3_R1143_U226, P3_U3066, P3_U3404);
  nand ginst20761 (P3_R1143_U227, P3_R1143_U124, P3_R1143_U225);
  or ginst20762 (P3_R1143_U228, P3_U3059, P3_U3401);
  nand ginst20763 (P3_R1143_U229, P3_R1143_U181, P3_R1143_U184);
  not ginst20764 (P3_R1143_U23, P3_U3410);
  not ginst20765 (P3_R1143_U230, P3_R1143_U145);
  nand ginst20766 (P3_R1143_U231, P3_U3063, P3_U3398);
  nand ginst20767 (P3_R1143_U232, P3_R1143_U400, P3_R1143_U401, P3_R1143_U42, P3_R1143_U43);
  nand ginst20768 (P3_R1143_U233, P3_R1143_U42, P3_R1143_U43);
  nand ginst20769 (P3_R1143_U234, P3_U3067, P3_U3395);
  nand ginst20770 (P3_R1143_U235, P3_R1143_U125, P3_R1143_U233);
  or ginst20771 (P3_R1143_U236, P3_U3082, P3_U3416);
  or ginst20772 (P3_R1143_U237, P3_U3061, P3_U3419);
  nand ginst20773 (P3_R1143_U238, P3_R1143_U177, P3_R1143_U6);
  nand ginst20774 (P3_R1143_U239, P3_U3061, P3_U3419);
  not ginst20775 (P3_R1143_U24, P3_U3401);
  nand ginst20776 (P3_R1143_U240, P3_R1143_U171, P3_R1143_U238);
  or ginst20777 (P3_R1143_U241, P3_U3061, P3_U3419);
  nand ginst20778 (P3_R1143_U242, P3_R1143_U126, P3_R1143_U144);
  nand ginst20779 (P3_R1143_U243, P3_R1143_U240, P3_R1143_U241);
  not ginst20780 (P3_R1143_U244, P3_R1143_U167);
  or ginst20781 (P3_R1143_U245, P3_U3079, P3_U3428);
  or ginst20782 (P3_R1143_U246, P3_U3071, P3_U3425);
  nand ginst20783 (P3_R1143_U247, P3_R1143_U174, P3_R1143_U7);
  nand ginst20784 (P3_R1143_U248, P3_U3079, P3_U3428);
  nand ginst20785 (P3_R1143_U249, P3_R1143_U129, P3_R1143_U247);
  not ginst20786 (P3_R1143_U25, P3_U3059);
  or ginst20787 (P3_R1143_U250, P3_U3062, P3_U3422);
  or ginst20788 (P3_R1143_U251, P3_U3079, P3_U3428);
  nand ginst20789 (P3_R1143_U252, P3_R1143_U128, P3_R1143_U167);
  nand ginst20790 (P3_R1143_U253, P3_R1143_U249, P3_R1143_U251);
  not ginst20791 (P3_R1143_U254, P3_R1143_U166);
  or ginst20792 (P3_R1143_U255, P3_U3078, P3_U3431);
  nand ginst20793 (P3_R1143_U256, P3_R1143_U166, P3_R1143_U255);
  nand ginst20794 (P3_R1143_U257, P3_U3078, P3_U3431);
  not ginst20795 (P3_R1143_U258, P3_R1143_U164);
  or ginst20796 (P3_R1143_U259, P3_U3073, P3_U3434);
  not ginst20797 (P3_R1143_U26, P3_U3066);
  nand ginst20798 (P3_R1143_U260, P3_R1143_U164, P3_R1143_U259);
  nand ginst20799 (P3_R1143_U261, P3_U3073, P3_U3434);
  not ginst20800 (P3_R1143_U262, P3_R1143_U92);
  or ginst20801 (P3_R1143_U263, P3_U3068, P3_U3440);
  or ginst20802 (P3_R1143_U264, P3_U3072, P3_U3437);
  not ginst20803 (P3_R1143_U265, P3_R1143_U59);
  nand ginst20804 (P3_R1143_U266, P3_R1143_U59, P3_R1143_U60);
  nand ginst20805 (P3_R1143_U267, P3_R1143_U266, P3_U3068);
  nand ginst20806 (P3_R1143_U268, P3_R1143_U265, P3_U3440);
  nand ginst20807 (P3_R1143_U269, P3_R1143_U8, P3_R1143_U92);
  not ginst20808 (P3_R1143_U27, P3_U3395);
  not ginst20809 (P3_R1143_U270, P3_R1143_U162);
  or ginst20810 (P3_R1143_U271, P3_U3075, P3_U3907);
  or ginst20811 (P3_R1143_U272, P3_U3080, P3_U3445);
  or ginst20812 (P3_R1143_U273, P3_U3074, P3_U3906);
  not ginst20813 (P3_R1143_U274, P3_R1143_U80);
  nand ginst20814 (P3_R1143_U275, P3_R1143_U274, P3_U3907);
  nand ginst20815 (P3_R1143_U276, P3_R1143_U275, P3_R1143_U90);
  nand ginst20816 (P3_R1143_U277, P3_R1143_U80, P3_R1143_U81);
  nand ginst20817 (P3_R1143_U278, P3_R1143_U276, P3_R1143_U277);
  nand ginst20818 (P3_R1143_U279, P3_R1143_U175, P3_R1143_U9);
  not ginst20819 (P3_R1143_U28, P3_U3067);
  nand ginst20820 (P3_R1143_U280, P3_U3074, P3_U3906);
  nand ginst20821 (P3_R1143_U281, P3_R1143_U278, P3_R1143_U279);
  or ginst20822 (P3_R1143_U282, P3_U3081, P3_U3443);
  or ginst20823 (P3_R1143_U283, P3_U3074, P3_U3906);
  nand ginst20824 (P3_R1143_U284, P3_R1143_U131, P3_R1143_U162);
  nand ginst20825 (P3_R1143_U285, P3_R1143_U281, P3_R1143_U283);
  not ginst20826 (P3_R1143_U286, P3_R1143_U159);
  or ginst20827 (P3_R1143_U287, P3_U3060, P3_U3905);
  nand ginst20828 (P3_R1143_U288, P3_R1143_U159, P3_R1143_U287);
  nand ginst20829 (P3_R1143_U289, P3_U3060, P3_U3905);
  not ginst20830 (P3_R1143_U29, P3_U3387);
  not ginst20831 (P3_R1143_U290, P3_R1143_U157);
  or ginst20832 (P3_R1143_U291, P3_U3065, P3_U3904);
  nand ginst20833 (P3_R1143_U292, P3_R1143_U157, P3_R1143_U291);
  nand ginst20834 (P3_R1143_U293, P3_U3065, P3_U3904);
  not ginst20835 (P3_R1143_U294, P3_R1143_U155);
  or ginst20836 (P3_R1143_U295, P3_U3057, P3_U3902);
  nand ginst20837 (P3_R1143_U296, P3_R1143_U173, P3_R1143_U176);
  not ginst20838 (P3_R1143_U297, P3_R1143_U86);
  or ginst20839 (P3_R1143_U298, P3_U3064, P3_U3903);
  nand ginst20840 (P3_R1143_U299, P3_R1143_U155, P3_R1143_U168, P3_R1143_U298);
  not ginst20841 (P3_R1143_U30, P3_U3076);
  not ginst20842 (P3_R1143_U300, P3_R1143_U153);
  or ginst20843 (P3_R1143_U301, P3_U3052, P3_U3900);
  nand ginst20844 (P3_R1143_U302, P3_U3052, P3_U3900);
  not ginst20845 (P3_R1143_U303, P3_R1143_U151);
  nand ginst20846 (P3_R1143_U304, P3_R1143_U151, P3_U3899);
  not ginst20847 (P3_R1143_U305, P3_R1143_U149);
  nand ginst20848 (P3_R1143_U306, P3_R1143_U155, P3_R1143_U298);
  not ginst20849 (P3_R1143_U307, P3_R1143_U89);
  or ginst20850 (P3_R1143_U308, P3_U3057, P3_U3902);
  nand ginst20851 (P3_R1143_U309, P3_R1143_U308, P3_R1143_U89);
  nand ginst20852 (P3_R1143_U31, P3_U3076, P3_U3387);
  nand ginst20853 (P3_R1143_U310, P3_R1143_U154, P3_R1143_U173, P3_R1143_U309);
  nand ginst20854 (P3_R1143_U311, P3_R1143_U173, P3_R1143_U307);
  nand ginst20855 (P3_R1143_U312, P3_U3056, P3_U3901);
  nand ginst20856 (P3_R1143_U313, P3_R1143_U168, P3_R1143_U311, P3_R1143_U312);
  or ginst20857 (P3_R1143_U314, P3_U3057, P3_U3902);
  nand ginst20858 (P3_R1143_U315, P3_R1143_U162, P3_R1143_U282);
  not ginst20859 (P3_R1143_U316, P3_R1143_U91);
  nand ginst20860 (P3_R1143_U317, P3_R1143_U9, P3_R1143_U91);
  nand ginst20861 (P3_R1143_U318, P3_R1143_U135, P3_R1143_U317);
  nand ginst20862 (P3_R1143_U319, P3_R1143_U278, P3_R1143_U317);
  not ginst20863 (P3_R1143_U32, P3_U3398);
  nand ginst20864 (P3_R1143_U320, P3_R1143_U319, P3_R1143_U453);
  or ginst20865 (P3_R1143_U321, P3_U3080, P3_U3445);
  nand ginst20866 (P3_R1143_U322, P3_R1143_U321, P3_R1143_U91);
  nand ginst20867 (P3_R1143_U323, P3_R1143_U136, P3_R1143_U322);
  nand ginst20868 (P3_R1143_U324, P3_R1143_U316, P3_R1143_U80);
  nand ginst20869 (P3_R1143_U325, P3_U3075, P3_U3907);
  nand ginst20870 (P3_R1143_U326, P3_R1143_U137, P3_R1143_U324);
  or ginst20871 (P3_R1143_U327, P3_U3077, P3_U3392);
  not ginst20872 (P3_R1143_U328, P3_R1143_U161);
  or ginst20873 (P3_R1143_U329, P3_U3080, P3_U3445);
  not ginst20874 (P3_R1143_U33, P3_U3063);
  or ginst20875 (P3_R1143_U330, P3_U3072, P3_U3437);
  nand ginst20876 (P3_R1143_U331, P3_R1143_U330, P3_R1143_U92);
  nand ginst20877 (P3_R1143_U332, P3_R1143_U138, P3_R1143_U331);
  nand ginst20878 (P3_R1143_U333, P3_R1143_U262, P3_R1143_U59);
  nand ginst20879 (P3_R1143_U334, P3_U3068, P3_U3440);
  nand ginst20880 (P3_R1143_U335, P3_R1143_U139, P3_R1143_U333);
  or ginst20881 (P3_R1143_U336, P3_U3072, P3_U3437);
  nand ginst20882 (P3_R1143_U337, P3_R1143_U167, P3_R1143_U250);
  not ginst20883 (P3_R1143_U338, P3_R1143_U93);
  or ginst20884 (P3_R1143_U339, P3_U3071, P3_U3425);
  nand ginst20885 (P3_R1143_U34, P3_U3059, P3_U3401);
  nand ginst20886 (P3_R1143_U340, P3_R1143_U339, P3_R1143_U93);
  nand ginst20887 (P3_R1143_U341, P3_R1143_U140, P3_R1143_U340);
  nand ginst20888 (P3_R1143_U342, P3_R1143_U172, P3_R1143_U338);
  nand ginst20889 (P3_R1143_U343, P3_U3079, P3_U3428);
  nand ginst20890 (P3_R1143_U344, P3_R1143_U141, P3_R1143_U342);
  or ginst20891 (P3_R1143_U345, P3_U3071, P3_U3425);
  or ginst20892 (P3_R1143_U346, P3_U3082, P3_U3416);
  nand ginst20893 (P3_R1143_U347, P3_R1143_U346, P3_R1143_U40);
  nand ginst20894 (P3_R1143_U348, P3_R1143_U142, P3_R1143_U347);
  nand ginst20895 (P3_R1143_U349, P3_R1143_U171, P3_R1143_U206);
  not ginst20896 (P3_R1143_U35, P3_U3404);
  nand ginst20897 (P3_R1143_U350, P3_U3061, P3_U3419);
  nand ginst20898 (P3_R1143_U351, P3_R1143_U143, P3_R1143_U349);
  nand ginst20899 (P3_R1143_U352, P3_R1143_U171, P3_R1143_U207);
  nand ginst20900 (P3_R1143_U353, P3_R1143_U204, P3_R1143_U63);
  nand ginst20901 (P3_R1143_U354, P3_R1143_U214, P3_R1143_U22);
  nand ginst20902 (P3_R1143_U355, P3_R1143_U228, P3_R1143_U34);
  nand ginst20903 (P3_R1143_U356, P3_R1143_U180, P3_R1143_U231);
  nand ginst20904 (P3_R1143_U357, P3_R1143_U173, P3_R1143_U314);
  nand ginst20905 (P3_R1143_U358, P3_R1143_U176, P3_R1143_U298);
  nand ginst20906 (P3_R1143_U359, P3_R1143_U329, P3_R1143_U80);
  not ginst20907 (P3_R1143_U36, P3_U3413);
  nand ginst20908 (P3_R1143_U360, P3_R1143_U282, P3_R1143_U77);
  nand ginst20909 (P3_R1143_U361, P3_R1143_U336, P3_R1143_U59);
  nand ginst20910 (P3_R1143_U362, P3_R1143_U172, P3_R1143_U345);
  nand ginst20911 (P3_R1143_U363, P3_R1143_U250, P3_R1143_U68);
  nand ginst20912 (P3_R1143_U364, P3_U3053, P3_U3899);
  nand ginst20913 (P3_R1143_U365, P3_R1143_U168, P3_R1143_U296);
  nand ginst20914 (P3_R1143_U366, P3_R1143_U295, P3_U3056);
  nand ginst20915 (P3_R1143_U367, P3_R1143_U295, P3_U3901);
  nand ginst20916 (P3_R1143_U368, P3_R1143_U168, P3_R1143_U296, P3_R1143_U301);
  nand ginst20917 (P3_R1143_U369, P3_R1143_U133, P3_R1143_U155, P3_R1143_U168);
  not ginst20918 (P3_R1143_U37, P3_U3083);
  nand ginst20919 (P3_R1143_U370, P3_R1143_U297, P3_R1143_U301);
  nand ginst20920 (P3_R1143_U371, P3_R1143_U39, P3_U3082);
  nand ginst20921 (P3_R1143_U372, P3_R1143_U38, P3_U3416);
  nand ginst20922 (P3_R1143_U373, P3_R1143_U371, P3_R1143_U372);
  nand ginst20923 (P3_R1143_U374, P3_R1143_U352, P3_R1143_U40);
  nand ginst20924 (P3_R1143_U375, P3_R1143_U206, P3_R1143_U373);
  nand ginst20925 (P3_R1143_U376, P3_R1143_U36, P3_U3083);
  nand ginst20926 (P3_R1143_U377, P3_R1143_U37, P3_U3413);
  nand ginst20927 (P3_R1143_U378, P3_R1143_U376, P3_R1143_U377);
  nand ginst20928 (P3_R1143_U379, P3_R1143_U144, P3_R1143_U353);
  not ginst20929 (P3_R1143_U38, P3_U3082);
  nand ginst20930 (P3_R1143_U380, P3_R1143_U203, P3_R1143_U378);
  nand ginst20931 (P3_R1143_U381, P3_R1143_U23, P3_U3069);
  nand ginst20932 (P3_R1143_U382, P3_R1143_U21, P3_U3410);
  nand ginst20933 (P3_R1143_U383, P3_R1143_U19, P3_U3070);
  nand ginst20934 (P3_R1143_U384, P3_R1143_U20, P3_U3407);
  nand ginst20935 (P3_R1143_U385, P3_R1143_U383, P3_R1143_U384);
  nand ginst20936 (P3_R1143_U386, P3_R1143_U354, P3_R1143_U41);
  nand ginst20937 (P3_R1143_U387, P3_R1143_U195, P3_R1143_U385);
  nand ginst20938 (P3_R1143_U388, P3_R1143_U35, P3_U3066);
  nand ginst20939 (P3_R1143_U389, P3_R1143_U26, P3_U3404);
  not ginst20940 (P3_R1143_U39, P3_U3416);
  nand ginst20941 (P3_R1143_U390, P3_R1143_U24, P3_U3059);
  nand ginst20942 (P3_R1143_U391, P3_R1143_U25, P3_U3401);
  nand ginst20943 (P3_R1143_U392, P3_R1143_U390, P3_R1143_U391);
  nand ginst20944 (P3_R1143_U393, P3_R1143_U355, P3_R1143_U44);
  nand ginst20945 (P3_R1143_U394, P3_R1143_U221, P3_R1143_U392);
  nand ginst20946 (P3_R1143_U395, P3_R1143_U32, P3_U3063);
  nand ginst20947 (P3_R1143_U396, P3_R1143_U33, P3_U3398);
  nand ginst20948 (P3_R1143_U397, P3_R1143_U395, P3_R1143_U396);
  nand ginst20949 (P3_R1143_U398, P3_R1143_U145, P3_R1143_U356);
  nand ginst20950 (P3_R1143_U399, P3_R1143_U230, P3_R1143_U397);
  and ginst20951 (P3_R1143_U4, P3_R1143_U178, P3_R1143_U179);
  nand ginst20952 (P3_R1143_U40, P3_R1143_U205, P3_R1143_U63);
  nand ginst20953 (P3_R1143_U400, P3_R1143_U27, P3_U3067);
  nand ginst20954 (P3_R1143_U401, P3_R1143_U28, P3_U3395);
  nand ginst20955 (P3_R1143_U402, P3_R1143_U147, P3_U3054);
  nand ginst20956 (P3_R1143_U403, P3_R1143_U146, P3_U3908);
  nand ginst20957 (P3_R1143_U404, P3_R1143_U147, P3_U3054);
  nand ginst20958 (P3_R1143_U405, P3_R1143_U146, P3_U3908);
  nand ginst20959 (P3_R1143_U406, P3_R1143_U404, P3_R1143_U405);
  nand ginst20960 (P3_R1143_U407, P3_R1143_U148, P3_R1143_U149);
  nand ginst20961 (P3_R1143_U408, P3_R1143_U305, P3_R1143_U406);
  nand ginst20962 (P3_R1143_U409, P3_R1143_U88, P3_U3053);
  nand ginst20963 (P3_R1143_U41, P3_R1143_U117, P3_R1143_U193);
  nand ginst20964 (P3_R1143_U410, P3_R1143_U87, P3_U3899);
  nand ginst20965 (P3_R1143_U411, P3_R1143_U88, P3_U3053);
  nand ginst20966 (P3_R1143_U412, P3_R1143_U87, P3_U3899);
  nand ginst20967 (P3_R1143_U413, P3_R1143_U411, P3_R1143_U412);
  nand ginst20968 (P3_R1143_U414, P3_R1143_U150, P3_R1143_U151);
  nand ginst20969 (P3_R1143_U415, P3_R1143_U303, P3_R1143_U413);
  nand ginst20970 (P3_R1143_U416, P3_R1143_U46, P3_U3052);
  nand ginst20971 (P3_R1143_U417, P3_R1143_U47, P3_U3900);
  nand ginst20972 (P3_R1143_U418, P3_R1143_U46, P3_U3052);
  nand ginst20973 (P3_R1143_U419, P3_R1143_U47, P3_U3900);
  nand ginst20974 (P3_R1143_U42, P3_R1143_U182, P3_R1143_U183);
  nand ginst20975 (P3_R1143_U420, P3_R1143_U418, P3_R1143_U419);
  nand ginst20976 (P3_R1143_U421, P3_R1143_U152, P3_R1143_U153);
  nand ginst20977 (P3_R1143_U422, P3_R1143_U300, P3_R1143_U420);
  nand ginst20978 (P3_R1143_U423, P3_R1143_U49, P3_U3056);
  nand ginst20979 (P3_R1143_U424, P3_R1143_U48, P3_U3901);
  nand ginst20980 (P3_R1143_U425, P3_R1143_U50, P3_U3057);
  nand ginst20981 (P3_R1143_U426, P3_R1143_U51, P3_U3902);
  nand ginst20982 (P3_R1143_U427, P3_R1143_U425, P3_R1143_U426);
  nand ginst20983 (P3_R1143_U428, P3_R1143_U357, P3_R1143_U89);
  nand ginst20984 (P3_R1143_U429, P3_R1143_U307, P3_R1143_U427);
  nand ginst20985 (P3_R1143_U43, P3_U3077, P3_U3392);
  nand ginst20986 (P3_R1143_U430, P3_R1143_U52, P3_U3064);
  nand ginst20987 (P3_R1143_U431, P3_R1143_U53, P3_U3903);
  nand ginst20988 (P3_R1143_U432, P3_R1143_U430, P3_R1143_U431);
  nand ginst20989 (P3_R1143_U433, P3_R1143_U155, P3_R1143_U358);
  nand ginst20990 (P3_R1143_U434, P3_R1143_U294, P3_R1143_U432);
  nand ginst20991 (P3_R1143_U435, P3_R1143_U84, P3_U3065);
  nand ginst20992 (P3_R1143_U436, P3_R1143_U85, P3_U3904);
  nand ginst20993 (P3_R1143_U437, P3_R1143_U84, P3_U3065);
  nand ginst20994 (P3_R1143_U438, P3_R1143_U85, P3_U3904);
  nand ginst20995 (P3_R1143_U439, P3_R1143_U437, P3_R1143_U438);
  nand ginst20996 (P3_R1143_U44, P3_R1143_U122, P3_R1143_U219);
  nand ginst20997 (P3_R1143_U440, P3_R1143_U156, P3_R1143_U157);
  nand ginst20998 (P3_R1143_U441, P3_R1143_U290, P3_R1143_U439);
  nand ginst20999 (P3_R1143_U442, P3_R1143_U82, P3_U3060);
  nand ginst21000 (P3_R1143_U443, P3_R1143_U83, P3_U3905);
  nand ginst21001 (P3_R1143_U444, P3_R1143_U82, P3_U3060);
  nand ginst21002 (P3_R1143_U445, P3_R1143_U83, P3_U3905);
  nand ginst21003 (P3_R1143_U446, P3_R1143_U444, P3_R1143_U445);
  nand ginst21004 (P3_R1143_U447, P3_R1143_U158, P3_R1143_U159);
  nand ginst21005 (P3_R1143_U448, P3_R1143_U286, P3_R1143_U446);
  nand ginst21006 (P3_R1143_U449, P3_R1143_U54, P3_U3074);
  nand ginst21007 (P3_R1143_U45, P3_R1143_U215, P3_R1143_U216);
  nand ginst21008 (P3_R1143_U450, P3_R1143_U55, P3_U3906);
  nand ginst21009 (P3_R1143_U451, P3_R1143_U54, P3_U3074);
  nand ginst21010 (P3_R1143_U452, P3_R1143_U55, P3_U3906);
  nand ginst21011 (P3_R1143_U453, P3_R1143_U451, P3_R1143_U452);
  nand ginst21012 (P3_R1143_U454, P3_R1143_U81, P3_U3075);
  nand ginst21013 (P3_R1143_U455, P3_R1143_U90, P3_U3907);
  nand ginst21014 (P3_R1143_U456, P3_R1143_U161, P3_R1143_U182);
  nand ginst21015 (P3_R1143_U457, P3_R1143_U31, P3_R1143_U328);
  nand ginst21016 (P3_R1143_U458, P3_R1143_U78, P3_U3080);
  nand ginst21017 (P3_R1143_U459, P3_R1143_U79, P3_U3445);
  not ginst21018 (P3_R1143_U46, P3_U3900);
  nand ginst21019 (P3_R1143_U460, P3_R1143_U458, P3_R1143_U459);
  nand ginst21020 (P3_R1143_U461, P3_R1143_U359, P3_R1143_U91);
  nand ginst21021 (P3_R1143_U462, P3_R1143_U316, P3_R1143_U460);
  nand ginst21022 (P3_R1143_U463, P3_R1143_U75, P3_U3081);
  nand ginst21023 (P3_R1143_U464, P3_R1143_U76, P3_U3443);
  nand ginst21024 (P3_R1143_U465, P3_R1143_U463, P3_R1143_U464);
  nand ginst21025 (P3_R1143_U466, P3_R1143_U162, P3_R1143_U360);
  nand ginst21026 (P3_R1143_U467, P3_R1143_U270, P3_R1143_U465);
  nand ginst21027 (P3_R1143_U468, P3_R1143_U60, P3_U3068);
  nand ginst21028 (P3_R1143_U469, P3_R1143_U58, P3_U3440);
  not ginst21029 (P3_R1143_U47, P3_U3052);
  nand ginst21030 (P3_R1143_U470, P3_R1143_U56, P3_U3072);
  nand ginst21031 (P3_R1143_U471, P3_R1143_U57, P3_U3437);
  nand ginst21032 (P3_R1143_U472, P3_R1143_U470, P3_R1143_U471);
  nand ginst21033 (P3_R1143_U473, P3_R1143_U361, P3_R1143_U92);
  nand ginst21034 (P3_R1143_U474, P3_R1143_U262, P3_R1143_U472);
  nand ginst21035 (P3_R1143_U475, P3_R1143_U73, P3_U3073);
  nand ginst21036 (P3_R1143_U476, P3_R1143_U74, P3_U3434);
  nand ginst21037 (P3_R1143_U477, P3_R1143_U73, P3_U3073);
  nand ginst21038 (P3_R1143_U478, P3_R1143_U74, P3_U3434);
  nand ginst21039 (P3_R1143_U479, P3_R1143_U477, P3_R1143_U478);
  not ginst21040 (P3_R1143_U48, P3_U3056);
  nand ginst21041 (P3_R1143_U480, P3_R1143_U163, P3_R1143_U164);
  nand ginst21042 (P3_R1143_U481, P3_R1143_U258, P3_R1143_U479);
  nand ginst21043 (P3_R1143_U482, P3_R1143_U71, P3_U3078);
  nand ginst21044 (P3_R1143_U483, P3_R1143_U72, P3_U3431);
  nand ginst21045 (P3_R1143_U484, P3_R1143_U71, P3_U3078);
  nand ginst21046 (P3_R1143_U485, P3_R1143_U72, P3_U3431);
  nand ginst21047 (P3_R1143_U486, P3_R1143_U484, P3_R1143_U485);
  nand ginst21048 (P3_R1143_U487, P3_R1143_U165, P3_R1143_U166);
  nand ginst21049 (P3_R1143_U488, P3_R1143_U254, P3_R1143_U486);
  nand ginst21050 (P3_R1143_U489, P3_R1143_U69, P3_U3079);
  not ginst21051 (P3_R1143_U49, P3_U3901);
  nand ginst21052 (P3_R1143_U490, P3_R1143_U70, P3_U3428);
  nand ginst21053 (P3_R1143_U491, P3_R1143_U64, P3_U3071);
  nand ginst21054 (P3_R1143_U492, P3_R1143_U65, P3_U3425);
  nand ginst21055 (P3_R1143_U493, P3_R1143_U491, P3_R1143_U492);
  nand ginst21056 (P3_R1143_U494, P3_R1143_U362, P3_R1143_U93);
  nand ginst21057 (P3_R1143_U495, P3_R1143_U338, P3_R1143_U493);
  nand ginst21058 (P3_R1143_U496, P3_R1143_U66, P3_U3062);
  nand ginst21059 (P3_R1143_U497, P3_R1143_U67, P3_U3422);
  nand ginst21060 (P3_R1143_U498, P3_R1143_U496, P3_R1143_U497);
  nand ginst21061 (P3_R1143_U499, P3_R1143_U167, P3_R1143_U363);
  and ginst21062 (P3_R1143_U5, P3_R1143_U196, P3_R1143_U197);
  not ginst21063 (P3_R1143_U50, P3_U3902);
  nand ginst21064 (P3_R1143_U500, P3_R1143_U244, P3_R1143_U498);
  nand ginst21065 (P3_R1143_U501, P3_R1143_U61, P3_U3061);
  nand ginst21066 (P3_R1143_U502, P3_R1143_U62, P3_U3419);
  nand ginst21067 (P3_R1143_U503, P3_R1143_U29, P3_U3076);
  nand ginst21068 (P3_R1143_U504, P3_R1143_U30, P3_U3387);
  not ginst21069 (P3_R1143_U51, P3_U3057);
  not ginst21070 (P3_R1143_U52, P3_U3903);
  not ginst21071 (P3_R1143_U53, P3_U3064);
  not ginst21072 (P3_R1143_U54, P3_U3906);
  not ginst21073 (P3_R1143_U55, P3_U3074);
  not ginst21074 (P3_R1143_U56, P3_U3437);
  not ginst21075 (P3_R1143_U57, P3_U3072);
  not ginst21076 (P3_R1143_U58, P3_U3068);
  nand ginst21077 (P3_R1143_U59, P3_U3072, P3_U3437);
  and ginst21078 (P3_R1143_U6, P3_R1143_U236, P3_R1143_U237);
  not ginst21079 (P3_R1143_U60, P3_U3440);
  not ginst21080 (P3_R1143_U61, P3_U3419);
  not ginst21081 (P3_R1143_U62, P3_U3061);
  nand ginst21082 (P3_R1143_U63, P3_U3083, P3_U3413);
  not ginst21083 (P3_R1143_U64, P3_U3425);
  not ginst21084 (P3_R1143_U65, P3_U3071);
  not ginst21085 (P3_R1143_U66, P3_U3422);
  not ginst21086 (P3_R1143_U67, P3_U3062);
  nand ginst21087 (P3_R1143_U68, P3_U3062, P3_U3422);
  not ginst21088 (P3_R1143_U69, P3_U3428);
  and ginst21089 (P3_R1143_U7, P3_R1143_U245, P3_R1143_U246);
  not ginst21090 (P3_R1143_U70, P3_U3079);
  not ginst21091 (P3_R1143_U71, P3_U3431);
  not ginst21092 (P3_R1143_U72, P3_U3078);
  not ginst21093 (P3_R1143_U73, P3_U3434);
  not ginst21094 (P3_R1143_U74, P3_U3073);
  not ginst21095 (P3_R1143_U75, P3_U3443);
  not ginst21096 (P3_R1143_U76, P3_U3081);
  nand ginst21097 (P3_R1143_U77, P3_U3081, P3_U3443);
  not ginst21098 (P3_R1143_U78, P3_U3445);
  not ginst21099 (P3_R1143_U79, P3_U3080);
  and ginst21100 (P3_R1143_U8, P3_R1143_U263, P3_R1143_U264);
  nand ginst21101 (P3_R1143_U80, P3_U3080, P3_U3445);
  not ginst21102 (P3_R1143_U81, P3_U3907);
  not ginst21103 (P3_R1143_U82, P3_U3905);
  not ginst21104 (P3_R1143_U83, P3_U3060);
  not ginst21105 (P3_R1143_U84, P3_U3904);
  not ginst21106 (P3_R1143_U85, P3_U3065);
  nand ginst21107 (P3_R1143_U86, P3_U3056, P3_U3901);
  not ginst21108 (P3_R1143_U87, P3_U3053);
  not ginst21109 (P3_R1143_U88, P3_U3899);
  nand ginst21110 (P3_R1143_U89, P3_R1143_U176, P3_R1143_U306);
  and ginst21111 (P3_R1143_U9, P3_R1143_U271, P3_R1143_U272);
  not ginst21112 (P3_R1143_U90, P3_U3075);
  nand ginst21113 (P3_R1143_U91, P3_R1143_U315, P3_R1143_U77);
  nand ginst21114 (P3_R1143_U92, P3_R1143_U260, P3_R1143_U261);
  nand ginst21115 (P3_R1143_U93, P3_R1143_U337, P3_R1143_U68);
  nand ginst21116 (P3_R1143_U94, P3_R1143_U456, P3_R1143_U457);
  nand ginst21117 (P3_R1143_U95, P3_R1143_U503, P3_R1143_U504);
  nand ginst21118 (P3_R1143_U96, P3_R1143_U374, P3_R1143_U375);
  nand ginst21119 (P3_R1143_U97, P3_R1143_U379, P3_R1143_U380);
  nand ginst21120 (P3_R1143_U98, P3_R1143_U386, P3_R1143_U387);
  nand ginst21121 (P3_R1143_U99, P3_R1143_U393, P3_R1143_U394);
  and ginst21122 (P3_R1158_U10, P3_R1158_U235, P3_R1158_U5);
  nand ginst21123 (P3_R1158_U100, P3_R1158_U463, P3_R1158_U464);
  nand ginst21124 (P3_R1158_U101, P3_R1158_U525, P3_R1158_U526);
  nand ginst21125 (P3_R1158_U102, P3_R1158_U532, P3_R1158_U533);
  and ginst21126 (P3_R1158_U103, P3_R1158_U209, P3_R1158_U320);
  and ginst21127 (P3_R1158_U104, P3_R1158_U12, P3_R1158_U141);
  nand ginst21128 (P3_R1158_U105, P3_R1158_U541, P3_R1158_U542);
  nand ginst21129 (P3_R1158_U106, P3_R1158_U546, P3_R1158_U547);
  nand ginst21130 (P3_R1158_U107, P3_R1158_U553, P3_R1158_U554);
  nand ginst21131 (P3_R1158_U108, P3_R1158_U560, P3_R1158_U561);
  nand ginst21132 (P3_R1158_U109, P3_R1158_U567, P3_R1158_U568);
  and ginst21133 (P3_R1158_U11, P3_R1158_U260, P3_R1158_U9);
  nand ginst21134 (P3_R1158_U110, P3_R1158_U574, P3_R1158_U575);
  nand ginst21135 (P3_R1158_U111, P3_R1158_U579, P3_R1158_U580);
  nand ginst21136 (P3_R1158_U112, P3_R1158_U586, P3_R1158_U587);
  nand ginst21137 (P3_R1158_U113, P3_R1158_U593, P3_R1158_U594);
  nand ginst21138 (P3_R1158_U114, P3_R1158_U600, P3_R1158_U601);
  nand ginst21139 (P3_R1158_U115, P3_R1158_U607, P3_R1158_U608);
  nand ginst21140 (P3_R1158_U116, P3_R1158_U614, P3_R1158_U615);
  nand ginst21141 (P3_R1158_U117, P3_R1158_U619, P3_R1158_U620);
  nand ginst21142 (P3_R1158_U118, P3_R1158_U626, P3_R1158_U627);
  and ginst21143 (P3_R1158_U119, P3_R1158_U73, P3_U3152);
  and ginst21144 (P3_R1158_U12, P3_R1158_U534, P3_R1158_U535);
  and ginst21145 (P3_R1158_U120, P3_R1158_U229, P3_R1158_U230);
  and ginst21146 (P3_R1158_U121, P3_R1158_U10, P3_R1158_U242);
  and ginst21147 (P3_R1158_U122, P3_R1158_U243, P3_R1158_U364);
  and ginst21148 (P3_R1158_U123, P3_R1158_U23, P3_R1158_U437, P3_R1158_U438);
  and ginst21149 (P3_R1158_U124, P3_R1158_U248, P3_R1158_U5);
  and ginst21150 (P3_R1158_U125, P3_R1158_U28, P3_R1158_U458, P3_R1158_U459);
  and ginst21151 (P3_R1158_U126, P3_R1158_U255, P3_R1158_U4);
  and ginst21152 (P3_R1158_U127, P3_R1158_U213, P3_R1158_U265);
  and ginst21153 (P3_R1158_U128, P3_R1158_U11, P3_R1158_U270);
  and ginst21154 (P3_R1158_U129, P3_R1158_U271, P3_R1158_U373);
  and ginst21155 (P3_R1158_U13, P3_R1158_U342, P3_R1158_U345);
  and ginst21156 (P3_R1158_U130, P3_R1158_U280, P3_R1158_U281);
  and ginst21157 (P3_R1158_U131, P3_R1158_U293, P3_R1158_U8);
  and ginst21158 (P3_R1158_U132, P3_R1158_U214, P3_R1158_U291);
  and ginst21159 (P3_R1158_U133, P3_R1158_U314, P3_R1158_U376);
  and ginst21160 (P3_R1158_U134, P3_R1158_U307, P3_R1158_U316);
  and ginst21161 (P3_R1158_U135, P3_R1158_U316, P3_R1158_U369);
  and ginst21162 (P3_R1158_U136, P3_R1158_U315, P3_R1158_U374);
  nand ginst21163 (P3_R1158_U137, P3_R1158_U519, P3_R1158_U520);
  and ginst21164 (P3_R1158_U138, P3_R1158_U38, P3_R1158_U515);
  and ginst21165 (P3_R1158_U139, P3_R1158_U215, P3_R1158_U320);
  and ginst21166 (P3_R1158_U14, P3_R1158_U333, P3_R1158_U336);
  and ginst21167 (P3_R1158_U140, P3_R1158_U218, P3_R1158_U320);
  and ginst21168 (P3_R1158_U141, P3_R1158_U59, P3_R1158_U60);
  and ginst21169 (P3_R1158_U142, P3_R1158_U319, P3_R1158_U391, P3_R1158_U392);
  and ginst21170 (P3_R1158_U143, P3_R1158_U214, P3_R1158_U562, P3_R1158_U563);
  and ginst21171 (P3_R1158_U144, P3_R1158_U328, P3_R1158_U8);
  and ginst21172 (P3_R1158_U145, P3_R1158_U42, P3_R1158_U588, P3_R1158_U589);
  and ginst21173 (P3_R1158_U146, P3_R1158_U335, P3_R1158_U7);
  and ginst21174 (P3_R1158_U147, P3_R1158_U213, P3_R1158_U609, P3_R1158_U610);
  and ginst21175 (P3_R1158_U148, P3_R1158_U344, P3_R1158_U6);
  nand ginst21176 (P3_R1158_U149, P3_R1158_U628, P3_R1158_U629);
  and ginst21177 (P3_R1158_U15, P3_R1158_U326, P3_R1158_U329);
  not ginst21178 (P3_R1158_U150, P3_U3416);
  and ginst21179 (P3_R1158_U151, P3_R1158_U396, P3_R1158_U397);
  not ginst21180 (P3_R1158_U152, P3_U3401);
  not ginst21181 (P3_R1158_U153, P3_U3392);
  not ginst21182 (P3_R1158_U154, P3_U3387);
  not ginst21183 (P3_R1158_U155, P3_U3398);
  not ginst21184 (P3_R1158_U156, P3_U3395);
  not ginst21185 (P3_R1158_U157, P3_U3404);
  not ginst21186 (P3_R1158_U158, P3_U3410);
  not ginst21187 (P3_R1158_U159, P3_U3407);
  and ginst21188 (P3_R1158_U16, P3_R1158_U142, P3_R1158_U536, P3_R1158_U537);
  not ginst21189 (P3_R1158_U160, P3_U3413);
  nand ginst21190 (P3_R1158_U161, P3_R1158_U122, P3_R1158_U383);
  and ginst21191 (P3_R1158_U162, P3_R1158_U430, P3_R1158_U431);
  nand ginst21192 (P3_R1158_U163, P3_R1158_U363, P3_R1158_U381);
  and ginst21193 (P3_R1158_U164, P3_R1158_U444, P3_R1158_U445);
  nand ginst21194 (P3_R1158_U165, P3_R1158_U211, P3_R1158_U233, P3_R1158_U356);
  and ginst21195 (P3_R1158_U166, P3_R1158_U451, P3_R1158_U452);
  nand ginst21196 (P3_R1158_U167, P3_R1158_U120, P3_R1158_U231);
  not ginst21197 (P3_R1158_U168, P3_U3900);
  not ginst21198 (P3_R1158_U169, P3_U3419);
  and ginst21199 (P3_R1158_U17, P3_R1158_U253, P3_R1158_U256);
  not ginst21200 (P3_R1158_U170, P3_U3422);
  not ginst21201 (P3_R1158_U171, P3_U3428);
  not ginst21202 (P3_R1158_U172, P3_U3425);
  not ginst21203 (P3_R1158_U173, P3_U3431);
  not ginst21204 (P3_R1158_U174, P3_U3434);
  not ginst21205 (P3_R1158_U175, P3_U3440);
  not ginst21206 (P3_R1158_U176, P3_U3437);
  not ginst21207 (P3_R1158_U177, P3_U3443);
  not ginst21208 (P3_R1158_U178, P3_U3906);
  not ginst21209 (P3_R1158_U179, P3_U3907);
  and ginst21210 (P3_R1158_U18, P3_R1158_U246, P3_R1158_U249);
  not ginst21211 (P3_R1158_U180, P3_U3445);
  not ginst21212 (P3_R1158_U181, P3_U3905);
  not ginst21213 (P3_R1158_U182, P3_U3904);
  not ginst21214 (P3_R1158_U183, P3_U3901);
  not ginst21215 (P3_R1158_U184, P3_U3902);
  not ginst21216 (P3_R1158_U185, P3_U3903);
  not ginst21217 (P3_R1158_U186, P3_U3053);
  not ginst21218 (P3_R1158_U187, P3_U3899);
  and ginst21219 (P3_R1158_U188, P3_R1158_U527, P3_R1158_U528);
  nand ginst21220 (P3_R1158_U189, P3_R1158_U310, P3_R1158_U311);
  nand ginst21221 (P3_R1158_U19, P3_R1158_U306, P3_U3056);
  nand ginst21222 (P3_R1158_U190, P3_R1158_U192, P3_R1158_U309);
  nand ginst21223 (P3_R1158_U191, P3_R1158_U190, P3_R1158_U60);
  nand ginst21224 (P3_R1158_U192, P3_R1158_U303, P3_R1158_U304);
  and ginst21225 (P3_R1158_U193, P3_R1158_U548, P3_R1158_U549);
  nand ginst21226 (P3_R1158_U194, P3_R1158_U299, P3_R1158_U300);
  and ginst21227 (P3_R1158_U195, P3_R1158_U555, P3_R1158_U556);
  nand ginst21228 (P3_R1158_U196, P3_R1158_U295, P3_R1158_U296);
  and ginst21229 (P3_R1158_U197, P3_R1158_U569, P3_R1158_U570);
  nand ginst21230 (P3_R1158_U198, P3_R1158_U220, P3_R1158_U221);
  nand ginst21231 (P3_R1158_U199, P3_R1158_U285, P3_R1158_U286);
  not ginst21232 (P3_R1158_U20, P3_U3152);
  and ginst21233 (P3_R1158_U200, P3_R1158_U581, P3_R1158_U582);
  nand ginst21234 (P3_R1158_U201, P3_R1158_U130, P3_R1158_U282);
  and ginst21235 (P3_R1158_U202, P3_R1158_U595, P3_R1158_U596);
  nand ginst21236 (P3_R1158_U203, P3_R1158_U129, P3_R1158_U389);
  and ginst21237 (P3_R1158_U204, P3_R1158_U602, P3_R1158_U603);
  nand ginst21238 (P3_R1158_U205, P3_R1158_U372, P3_R1158_U387);
  nand ginst21239 (P3_R1158_U206, P3_R1158_U385, P3_R1158_U50);
  and ginst21240 (P3_R1158_U207, P3_R1158_U621, P3_R1158_U622);
  nand ginst21241 (P3_R1158_U208, P3_R1158_U210, P3_R1158_U258, P3_R1158_U357);
  nand ginst21242 (P3_R1158_U209, P3_R1158_U19, P3_R1158_U367);
  not ginst21243 (P3_R1158_U21, P3_U3083);
  nand ginst21244 (P3_R1158_U210, P3_R1158_U161, P3_R1158_U65);
  nand ginst21245 (P3_R1158_U211, P3_R1158_U167, P3_R1158_U74);
  not ginst21246 (P3_R1158_U212, P3_R1158_U28);
  nand ginst21247 (P3_R1158_U213, P3_R1158_U82, P3_U3071);
  nand ginst21248 (P3_R1158_U214, P3_R1158_U90, P3_U3075);
  not ginst21249 (P3_R1158_U215, P3_R1158_U59);
  not ginst21250 (P3_R1158_U216, P3_R1158_U47);
  not ginst21251 (P3_R1158_U217, P3_R1158_U55);
  not ginst21252 (P3_R1158_U218, P3_R1158_U60);
  nand ginst21253 (P3_R1158_U219, P3_R1158_U20, P3_R1158_U409);
  not ginst21254 (P3_R1158_U22, P3_U3070);
  nand ginst21255 (P3_R1158_U220, P3_R1158_U219, P3_U3076);
  nand ginst21256 (P3_R1158_U221, P3_R1158_U73, P3_U3152);
  not ginst21257 (P3_R1158_U222, P3_R1158_U198);
  nand ginst21258 (P3_R1158_U223, P3_R1158_U30, P3_R1158_U406);
  nand ginst21259 (P3_R1158_U224, P3_R1158_U72, P3_U3077);
  not ginst21260 (P3_R1158_U225, P3_R1158_U36);
  nand ginst21261 (P3_R1158_U226, P3_R1158_U29, P3_R1158_U412);
  nand ginst21262 (P3_R1158_U227, P3_R1158_U27, P3_R1158_U415);
  nand ginst21263 (P3_R1158_U228, P3_R1158_U28, P3_R1158_U29);
  nand ginst21264 (P3_R1158_U229, P3_R1158_U228, P3_R1158_U71);
  nand ginst21265 (P3_R1158_U23, P3_R1158_U67, P3_U3070);
  nand ginst21266 (P3_R1158_U230, P3_R1158_U212, P3_U3063);
  nand ginst21267 (P3_R1158_U231, P3_R1158_U36, P3_R1158_U4);
  not ginst21268 (P3_R1158_U232, P3_R1158_U167);
  nand ginst21269 (P3_R1158_U233, P3_R1158_U167, P3_U3059);
  not ginst21270 (P3_R1158_U234, P3_R1158_U165);
  nand ginst21271 (P3_R1158_U235, P3_R1158_U25, P3_R1158_U418);
  not ginst21272 (P3_R1158_U236, P3_R1158_U26);
  nand ginst21273 (P3_R1158_U237, P3_R1158_U24, P3_R1158_U421);
  nand ginst21274 (P3_R1158_U238, P3_R1158_U22, P3_R1158_U424);
  not ginst21275 (P3_R1158_U239, P3_R1158_U23);
  not ginst21276 (P3_R1158_U24, P3_U3069);
  nand ginst21277 (P3_R1158_U240, P3_R1158_U23, P3_R1158_U24);
  nand ginst21278 (P3_R1158_U241, P3_R1158_U239, P3_U3069);
  nand ginst21279 (P3_R1158_U242, P3_R1158_U21, P3_R1158_U427);
  nand ginst21280 (P3_R1158_U243, P3_R1158_U66, P3_U3083);
  nand ginst21281 (P3_R1158_U244, P3_R1158_U22, P3_R1158_U424);
  nand ginst21282 (P3_R1158_U245, P3_R1158_U244, P3_R1158_U35);
  nand ginst21283 (P3_R1158_U246, P3_R1158_U123, P3_R1158_U245);
  nand ginst21284 (P3_R1158_U247, P3_R1158_U23, P3_R1158_U380);
  nand ginst21285 (P3_R1158_U248, P3_R1158_U68, P3_U3069);
  nand ginst21286 (P3_R1158_U249, P3_R1158_U124, P3_R1158_U247);
  not ginst21287 (P3_R1158_U25, P3_U3066);
  nand ginst21288 (P3_R1158_U250, P3_R1158_U22, P3_R1158_U424);
  nand ginst21289 (P3_R1158_U251, P3_R1158_U27, P3_R1158_U415);
  nand ginst21290 (P3_R1158_U252, P3_R1158_U251, P3_R1158_U36);
  nand ginst21291 (P3_R1158_U253, P3_R1158_U125, P3_R1158_U252);
  nand ginst21292 (P3_R1158_U254, P3_R1158_U225, P3_R1158_U28);
  nand ginst21293 (P3_R1158_U255, P3_R1158_U71, P3_U3063);
  nand ginst21294 (P3_R1158_U256, P3_R1158_U126, P3_R1158_U254);
  nand ginst21295 (P3_R1158_U257, P3_R1158_U27, P3_R1158_U415);
  nand ginst21296 (P3_R1158_U258, P3_R1158_U161, P3_U3082);
  not ginst21297 (P3_R1158_U259, P3_R1158_U208);
  nand ginst21298 (P3_R1158_U26, P3_R1158_U69, P3_U3066);
  nand ginst21299 (P3_R1158_U260, P3_R1158_U470, P3_R1158_U49);
  not ginst21300 (P3_R1158_U261, P3_R1158_U50);
  nand ginst21301 (P3_R1158_U262, P3_R1158_U476, P3_R1158_U48);
  nand ginst21302 (P3_R1158_U263, P3_R1158_U45, P3_R1158_U479);
  nand ginst21303 (P3_R1158_U264, P3_R1158_U216, P3_R1158_U6);
  nand ginst21304 (P3_R1158_U265, P3_R1158_U83, P3_U3079);
  nand ginst21305 (P3_R1158_U266, P3_R1158_U127, P3_R1158_U264);
  nand ginst21306 (P3_R1158_U267, P3_R1158_U46, P3_R1158_U473);
  nand ginst21307 (P3_R1158_U268, P3_R1158_U476, P3_R1158_U48);
  nand ginst21308 (P3_R1158_U269, P3_R1158_U266, P3_R1158_U268);
  not ginst21309 (P3_R1158_U27, P3_U3067);
  nand ginst21310 (P3_R1158_U270, P3_R1158_U44, P3_R1158_U482);
  nand ginst21311 (P3_R1158_U271, P3_R1158_U81, P3_U3078);
  nand ginst21312 (P3_R1158_U272, P3_R1158_U485, P3_R1158_U51);
  nand ginst21313 (P3_R1158_U273, P3_R1158_U203, P3_R1158_U272);
  nand ginst21314 (P3_R1158_U274, P3_R1158_U86, P3_U3073);
  not ginst21315 (P3_R1158_U275, P3_R1158_U62);
  nand ginst21316 (P3_R1158_U276, P3_R1158_U43, P3_R1158_U488);
  nand ginst21317 (P3_R1158_U277, P3_R1158_U41, P3_R1158_U491);
  not ginst21318 (P3_R1158_U278, P3_R1158_U42);
  nand ginst21319 (P3_R1158_U279, P3_R1158_U42, P3_R1158_U43);
  nand ginst21320 (P3_R1158_U28, P3_R1158_U70, P3_U3067);
  nand ginst21321 (P3_R1158_U280, P3_R1158_U279, P3_R1158_U80);
  nand ginst21322 (P3_R1158_U281, P3_R1158_U278, P3_U3068);
  nand ginst21323 (P3_R1158_U282, P3_R1158_U62, P3_R1158_U7);
  not ginst21324 (P3_R1158_U283, P3_R1158_U201);
  nand ginst21325 (P3_R1158_U284, P3_R1158_U494, P3_R1158_U52);
  nand ginst21326 (P3_R1158_U285, P3_R1158_U201, P3_R1158_U284);
  nand ginst21327 (P3_R1158_U286, P3_R1158_U87, P3_U3081);
  not ginst21328 (P3_R1158_U287, P3_R1158_U199);
  nand ginst21329 (P3_R1158_U288, P3_R1158_U497, P3_R1158_U56);
  nand ginst21330 (P3_R1158_U289, P3_R1158_U500, P3_R1158_U53);
  not ginst21331 (P3_R1158_U29, P3_U3063);
  nand ginst21332 (P3_R1158_U290, P3_R1158_U217, P3_R1158_U8);
  nand ginst21333 (P3_R1158_U291, P3_R1158_U89, P3_U3074);
  nand ginst21334 (P3_R1158_U292, P3_R1158_U132, P3_R1158_U290);
  nand ginst21335 (P3_R1158_U293, P3_R1158_U503, P3_R1158_U54);
  nand ginst21336 (P3_R1158_U294, P3_R1158_U497, P3_R1158_U56);
  nand ginst21337 (P3_R1158_U295, P3_R1158_U131, P3_R1158_U199);
  nand ginst21338 (P3_R1158_U296, P3_R1158_U292, P3_R1158_U294);
  not ginst21339 (P3_R1158_U297, P3_R1158_U196);
  nand ginst21340 (P3_R1158_U298, P3_R1158_U506, P3_R1158_U57);
  nand ginst21341 (P3_R1158_U299, P3_R1158_U196, P3_R1158_U298);
  not ginst21342 (P3_R1158_U30, P3_U3077);
  nand ginst21343 (P3_R1158_U300, P3_R1158_U91, P3_U3060);
  not ginst21344 (P3_R1158_U301, P3_R1158_U194);
  nand ginst21345 (P3_R1158_U302, P3_R1158_U509, P3_R1158_U58);
  nand ginst21346 (P3_R1158_U303, P3_R1158_U194, P3_R1158_U302);
  nand ginst21347 (P3_R1158_U304, P3_R1158_U92, P3_U3065);
  not ginst21348 (P3_R1158_U305, P3_R1158_U192);
  nand ginst21349 (P3_R1158_U306, P3_R1158_U38, P3_R1158_U515);
  nand ginst21350 (P3_R1158_U307, P3_R1158_U308, P3_R1158_U59, P3_R1158_U60);
  nand ginst21351 (P3_R1158_U308, P3_R1158_U78, P3_U3056);
  nand ginst21352 (P3_R1158_U309, P3_R1158_U39, P3_R1158_U518);
  not ginst21353 (P3_R1158_U31, P3_U3076);
  nand ginst21354 (P3_R1158_U310, P3_R1158_U192, P3_R1158_U369);
  nand ginst21355 (P3_R1158_U311, P3_R1158_U307, P3_R1158_U366);
  not ginst21356 (P3_R1158_U312, P3_R1158_U189);
  nand ginst21357 (P3_R1158_U313, P3_R1158_U37, P3_R1158_U467);
  nand ginst21358 (P3_R1158_U314, P3_R1158_U75, P3_U3052);
  nand ginst21359 (P3_R1158_U315, P3_R1158_U75, P3_U3052);
  nand ginst21360 (P3_R1158_U316, P3_R1158_U37, P3_R1158_U467);
  not ginst21361 (P3_R1158_U317, P3_R1158_U190);
  not ginst21362 (P3_R1158_U318, P3_R1158_U191);
  nand ginst21363 (P3_R1158_U319, P3_R1158_U12, P3_R1158_U138);
  not ginst21364 (P3_R1158_U32, P3_U3059);
  nand ginst21365 (P3_R1158_U320, P3_R1158_U78, P3_U3056);
  nand ginst21366 (P3_R1158_U321, P3_R1158_U38, P3_R1158_U515);
  nand ginst21367 (P3_R1158_U322, P3_R1158_U199, P3_R1158_U293);
  not ginst21368 (P3_R1158_U323, P3_R1158_U61);
  nand ginst21369 (P3_R1158_U324, P3_R1158_U500, P3_R1158_U53);
  nand ginst21370 (P3_R1158_U325, P3_R1158_U324, P3_R1158_U61);
  nand ginst21371 (P3_R1158_U326, P3_R1158_U143, P3_R1158_U325);
  nand ginst21372 (P3_R1158_U327, P3_R1158_U214, P3_R1158_U323);
  nand ginst21373 (P3_R1158_U328, P3_R1158_U89, P3_U3074);
  nand ginst21374 (P3_R1158_U329, P3_R1158_U144, P3_R1158_U327);
  not ginst21375 (P3_R1158_U33, P3_U3082);
  nand ginst21376 (P3_R1158_U330, P3_R1158_U500, P3_R1158_U53);
  nand ginst21377 (P3_R1158_U331, P3_R1158_U41, P3_R1158_U491);
  nand ginst21378 (P3_R1158_U332, P3_R1158_U331, P3_R1158_U62);
  nand ginst21379 (P3_R1158_U333, P3_R1158_U145, P3_R1158_U332);
  nand ginst21380 (P3_R1158_U334, P3_R1158_U275, P3_R1158_U42);
  nand ginst21381 (P3_R1158_U335, P3_R1158_U80, P3_U3068);
  nand ginst21382 (P3_R1158_U336, P3_R1158_U146, P3_R1158_U334);
  nand ginst21383 (P3_R1158_U337, P3_R1158_U41, P3_R1158_U491);
  nand ginst21384 (P3_R1158_U338, P3_R1158_U206, P3_R1158_U267);
  not ginst21385 (P3_R1158_U339, P3_R1158_U64);
  nand ginst21386 (P3_R1158_U34, P3_R1158_U241, P3_R1158_U359, P3_R1158_U362);
  nand ginst21387 (P3_R1158_U340, P3_R1158_U45, P3_R1158_U479);
  nand ginst21388 (P3_R1158_U341, P3_R1158_U340, P3_R1158_U64);
  nand ginst21389 (P3_R1158_U342, P3_R1158_U147, P3_R1158_U341);
  nand ginst21390 (P3_R1158_U343, P3_R1158_U213, P3_R1158_U339);
  nand ginst21391 (P3_R1158_U344, P3_R1158_U83, P3_U3079);
  nand ginst21392 (P3_R1158_U345, P3_R1158_U148, P3_R1158_U343);
  nand ginst21393 (P3_R1158_U346, P3_R1158_U45, P3_R1158_U479);
  nand ginst21394 (P3_R1158_U347, P3_R1158_U23, P3_R1158_U250);
  nand ginst21395 (P3_R1158_U348, P3_R1158_U257, P3_R1158_U28);
  nand ginst21396 (P3_R1158_U349, P3_R1158_U321, P3_R1158_U59);
  nand ginst21397 (P3_R1158_U35, P3_R1158_U26, P3_R1158_U379);
  nand ginst21398 (P3_R1158_U350, P3_R1158_U309, P3_R1158_U60);
  nand ginst21399 (P3_R1158_U351, P3_R1158_U214, P3_R1158_U330);
  nand ginst21400 (P3_R1158_U352, P3_R1158_U293, P3_R1158_U55);
  nand ginst21401 (P3_R1158_U353, P3_R1158_U337, P3_R1158_U42);
  nand ginst21402 (P3_R1158_U354, P3_R1158_U213, P3_R1158_U346);
  nand ginst21403 (P3_R1158_U355, P3_R1158_U267, P3_R1158_U47);
  nand ginst21404 (P3_R1158_U356, P3_R1158_U74, P3_U3059);
  nand ginst21405 (P3_R1158_U357, P3_R1158_U65, P3_U3082);
  nand ginst21406 (P3_R1158_U358, P3_R1158_U133, P3_R1158_U310);
  nand ginst21407 (P3_R1158_U359, P3_R1158_U240, P3_R1158_U68);
  nand ginst21408 (P3_R1158_U36, P3_R1158_U224, P3_R1158_U360, P3_R1158_U361);
  nand ginst21409 (P3_R1158_U360, P3_R1158_U219, P3_R1158_U223, P3_U3076);
  nand ginst21410 (P3_R1158_U361, P3_R1158_U119, P3_R1158_U223);
  nand ginst21411 (P3_R1158_U362, P3_R1158_U236, P3_R1158_U5);
  not ginst21412 (P3_R1158_U363, P3_R1158_U34);
  nand ginst21413 (P3_R1158_U364, P3_R1158_U242, P3_R1158_U34);
  nand ginst21414 (P3_R1158_U365, P3_R1158_U261, P3_R1158_U9);
  nand ginst21415 (P3_R1158_U366, P3_R1158_U19, P3_R1158_U308, P3_R1158_U367);
  nand ginst21416 (P3_R1158_U367, P3_R1158_U306, P3_R1158_U78);
  not ginst21417 (P3_R1158_U368, P3_R1158_U19);
  nand ginst21418 (P3_R1158_U369, P3_R1158_U370, P3_R1158_U371);
  not ginst21419 (P3_R1158_U37, P3_U3052);
  nand ginst21420 (P3_R1158_U370, P3_R1158_U306, P3_R1158_U309, P3_R1158_U78);
  nand ginst21421 (P3_R1158_U371, P3_R1158_U309, P3_R1158_U368);
  not ginst21422 (P3_R1158_U372, P3_R1158_U63);
  nand ginst21423 (P3_R1158_U373, P3_R1158_U270, P3_R1158_U63);
  nand ginst21424 (P3_R1158_U374, P3_R1158_U134, P3_R1158_U366);
  nand ginst21425 (P3_R1158_U375, P3_R1158_U135, P3_R1158_U192);
  nand ginst21426 (P3_R1158_U376, P3_R1158_U377, P3_R1158_U378);
  nand ginst21427 (P3_R1158_U377, P3_R1158_U308, P3_R1158_U59, P3_R1158_U60);
  nand ginst21428 (P3_R1158_U378, P3_R1158_U19, P3_R1158_U308, P3_R1158_U367);
  nand ginst21429 (P3_R1158_U379, P3_R1158_U165, P3_R1158_U235);
  not ginst21430 (P3_R1158_U38, P3_U3057);
  not ginst21431 (P3_R1158_U380, P3_R1158_U35);
  nand ginst21432 (P3_R1158_U381, P3_R1158_U10, P3_R1158_U165);
  not ginst21433 (P3_R1158_U382, P3_R1158_U163);
  nand ginst21434 (P3_R1158_U383, P3_R1158_U121, P3_R1158_U165);
  not ginst21435 (P3_R1158_U384, P3_R1158_U161);
  nand ginst21436 (P3_R1158_U385, P3_R1158_U208, P3_R1158_U260);
  not ginst21437 (P3_R1158_U386, P3_R1158_U206);
  nand ginst21438 (P3_R1158_U387, P3_R1158_U11, P3_R1158_U208);
  not ginst21439 (P3_R1158_U388, P3_R1158_U205);
  nand ginst21440 (P3_R1158_U389, P3_R1158_U128, P3_R1158_U208);
  not ginst21441 (P3_R1158_U39, P3_U3064);
  not ginst21442 (P3_R1158_U390, P3_R1158_U203);
  nand ginst21443 (P3_R1158_U391, P3_R1158_U139, P3_R1158_U209);
  nand ginst21444 (P3_R1158_U392, P3_R1158_U140, P3_R1158_U209);
  nand ginst21445 (P3_R1158_U393, P3_R1158_U150, P3_U3152);
  nand ginst21446 (P3_R1158_U394, P3_R1158_U20, P3_U3416);
  not ginst21447 (P3_R1158_U395, P3_R1158_U65);
  nand ginst21448 (P3_R1158_U396, P3_R1158_U395, P3_U3082);
  nand ginst21449 (P3_R1158_U397, P3_R1158_U33, P3_R1158_U65);
  nand ginst21450 (P3_R1158_U398, P3_R1158_U395, P3_U3082);
  nand ginst21451 (P3_R1158_U399, P3_R1158_U33, P3_R1158_U65);
  and ginst21452 (P3_R1158_U4, P3_R1158_U226, P3_R1158_U227);
  not ginst21453 (P3_R1158_U40, P3_U3056);
  nand ginst21454 (P3_R1158_U400, P3_R1158_U398, P3_R1158_U399);
  nand ginst21455 (P3_R1158_U401, P3_R1158_U152, P3_U3152);
  nand ginst21456 (P3_R1158_U402, P3_R1158_U20, P3_U3401);
  not ginst21457 (P3_R1158_U403, P3_R1158_U74);
  nand ginst21458 (P3_R1158_U404, P3_R1158_U153, P3_U3152);
  nand ginst21459 (P3_R1158_U405, P3_R1158_U20, P3_U3392);
  not ginst21460 (P3_R1158_U406, P3_R1158_U72);
  nand ginst21461 (P3_R1158_U407, P3_R1158_U154, P3_U3152);
  nand ginst21462 (P3_R1158_U408, P3_R1158_U20, P3_U3387);
  not ginst21463 (P3_R1158_U409, P3_R1158_U73);
  not ginst21464 (P3_R1158_U41, P3_U3072);
  nand ginst21465 (P3_R1158_U410, P3_R1158_U155, P3_U3152);
  nand ginst21466 (P3_R1158_U411, P3_R1158_U20, P3_U3398);
  not ginst21467 (P3_R1158_U412, P3_R1158_U71);
  nand ginst21468 (P3_R1158_U413, P3_R1158_U156, P3_U3152);
  nand ginst21469 (P3_R1158_U414, P3_R1158_U20, P3_U3395);
  not ginst21470 (P3_R1158_U415, P3_R1158_U70);
  nand ginst21471 (P3_R1158_U416, P3_R1158_U157, P3_U3152);
  nand ginst21472 (P3_R1158_U417, P3_R1158_U20, P3_U3404);
  not ginst21473 (P3_R1158_U418, P3_R1158_U69);
  nand ginst21474 (P3_R1158_U419, P3_R1158_U158, P3_U3152);
  nand ginst21475 (P3_R1158_U42, P3_R1158_U79, P3_U3072);
  nand ginst21476 (P3_R1158_U420, P3_R1158_U20, P3_U3410);
  not ginst21477 (P3_R1158_U421, P3_R1158_U68);
  nand ginst21478 (P3_R1158_U422, P3_R1158_U159, P3_U3152);
  nand ginst21479 (P3_R1158_U423, P3_R1158_U20, P3_U3407);
  not ginst21480 (P3_R1158_U424, P3_R1158_U67);
  nand ginst21481 (P3_R1158_U425, P3_R1158_U160, P3_U3152);
  nand ginst21482 (P3_R1158_U426, P3_R1158_U20, P3_U3413);
  not ginst21483 (P3_R1158_U427, P3_R1158_U66);
  nand ginst21484 (P3_R1158_U428, P3_R1158_U151, P3_R1158_U161);
  nand ginst21485 (P3_R1158_U429, P3_R1158_U384, P3_R1158_U400);
  not ginst21486 (P3_R1158_U43, P3_U3068);
  nand ginst21487 (P3_R1158_U430, P3_R1158_U427, P3_U3083);
  nand ginst21488 (P3_R1158_U431, P3_R1158_U21, P3_R1158_U66);
  nand ginst21489 (P3_R1158_U432, P3_R1158_U427, P3_U3083);
  nand ginst21490 (P3_R1158_U433, P3_R1158_U21, P3_R1158_U66);
  nand ginst21491 (P3_R1158_U434, P3_R1158_U432, P3_R1158_U433);
  nand ginst21492 (P3_R1158_U435, P3_R1158_U162, P3_R1158_U163);
  nand ginst21493 (P3_R1158_U436, P3_R1158_U382, P3_R1158_U434);
  nand ginst21494 (P3_R1158_U437, P3_R1158_U421, P3_U3069);
  nand ginst21495 (P3_R1158_U438, P3_R1158_U24, P3_R1158_U68);
  nand ginst21496 (P3_R1158_U439, P3_R1158_U424, P3_U3070);
  not ginst21497 (P3_R1158_U44, P3_U3078);
  nand ginst21498 (P3_R1158_U440, P3_R1158_U22, P3_R1158_U67);
  nand ginst21499 (P3_R1158_U441, P3_R1158_U439, P3_R1158_U440);
  nand ginst21500 (P3_R1158_U442, P3_R1158_U347, P3_R1158_U35);
  nand ginst21501 (P3_R1158_U443, P3_R1158_U380, P3_R1158_U441);
  nand ginst21502 (P3_R1158_U444, P3_R1158_U418, P3_U3066);
  nand ginst21503 (P3_R1158_U445, P3_R1158_U25, P3_R1158_U69);
  nand ginst21504 (P3_R1158_U446, P3_R1158_U418, P3_U3066);
  nand ginst21505 (P3_R1158_U447, P3_R1158_U25, P3_R1158_U69);
  nand ginst21506 (P3_R1158_U448, P3_R1158_U446, P3_R1158_U447);
  nand ginst21507 (P3_R1158_U449, P3_R1158_U164, P3_R1158_U165);
  not ginst21508 (P3_R1158_U45, P3_U3071);
  nand ginst21509 (P3_R1158_U450, P3_R1158_U234, P3_R1158_U448);
  nand ginst21510 (P3_R1158_U451, P3_R1158_U403, P3_U3059);
  nand ginst21511 (P3_R1158_U452, P3_R1158_U32, P3_R1158_U74);
  nand ginst21512 (P3_R1158_U453, P3_R1158_U403, P3_U3059);
  nand ginst21513 (P3_R1158_U454, P3_R1158_U32, P3_R1158_U74);
  nand ginst21514 (P3_R1158_U455, P3_R1158_U453, P3_R1158_U454);
  nand ginst21515 (P3_R1158_U456, P3_R1158_U166, P3_R1158_U167);
  nand ginst21516 (P3_R1158_U457, P3_R1158_U232, P3_R1158_U455);
  nand ginst21517 (P3_R1158_U458, P3_R1158_U412, P3_U3063);
  nand ginst21518 (P3_R1158_U459, P3_R1158_U29, P3_R1158_U71);
  not ginst21519 (P3_R1158_U46, P3_U3062);
  nand ginst21520 (P3_R1158_U460, P3_R1158_U415, P3_U3067);
  nand ginst21521 (P3_R1158_U461, P3_R1158_U27, P3_R1158_U70);
  nand ginst21522 (P3_R1158_U462, P3_R1158_U460, P3_R1158_U461);
  nand ginst21523 (P3_R1158_U463, P3_R1158_U348, P3_R1158_U36);
  nand ginst21524 (P3_R1158_U464, P3_R1158_U225, P3_R1158_U462);
  nand ginst21525 (P3_R1158_U465, P3_R1158_U168, P3_U3152);
  nand ginst21526 (P3_R1158_U466, P3_R1158_U20, P3_U3900);
  not ginst21527 (P3_R1158_U467, P3_R1158_U75);
  nand ginst21528 (P3_R1158_U468, P3_R1158_U169, P3_U3152);
  nand ginst21529 (P3_R1158_U469, P3_R1158_U20, P3_U3419);
  nand ginst21530 (P3_R1158_U47, P3_R1158_U84, P3_U3062);
  not ginst21531 (P3_R1158_U470, P3_R1158_U85);
  nand ginst21532 (P3_R1158_U471, P3_R1158_U170, P3_U3152);
  nand ginst21533 (P3_R1158_U472, P3_R1158_U20, P3_U3422);
  not ginst21534 (P3_R1158_U473, P3_R1158_U84);
  nand ginst21535 (P3_R1158_U474, P3_R1158_U171, P3_U3152);
  nand ginst21536 (P3_R1158_U475, P3_R1158_U20, P3_U3428);
  not ginst21537 (P3_R1158_U476, P3_R1158_U83);
  nand ginst21538 (P3_R1158_U477, P3_R1158_U172, P3_U3152);
  nand ginst21539 (P3_R1158_U478, P3_R1158_U20, P3_U3425);
  not ginst21540 (P3_R1158_U479, P3_R1158_U82);
  not ginst21541 (P3_R1158_U48, P3_U3079);
  nand ginst21542 (P3_R1158_U480, P3_R1158_U173, P3_U3152);
  nand ginst21543 (P3_R1158_U481, P3_R1158_U20, P3_U3431);
  not ginst21544 (P3_R1158_U482, P3_R1158_U81);
  nand ginst21545 (P3_R1158_U483, P3_R1158_U174, P3_U3152);
  nand ginst21546 (P3_R1158_U484, P3_R1158_U20, P3_U3434);
  not ginst21547 (P3_R1158_U485, P3_R1158_U86);
  nand ginst21548 (P3_R1158_U486, P3_R1158_U175, P3_U3152);
  nand ginst21549 (P3_R1158_U487, P3_R1158_U20, P3_U3440);
  not ginst21550 (P3_R1158_U488, P3_R1158_U80);
  nand ginst21551 (P3_R1158_U489, P3_R1158_U176, P3_U3152);
  not ginst21552 (P3_R1158_U49, P3_U3061);
  nand ginst21553 (P3_R1158_U490, P3_R1158_U20, P3_U3437);
  not ginst21554 (P3_R1158_U491, P3_R1158_U79);
  nand ginst21555 (P3_R1158_U492, P3_R1158_U177, P3_U3152);
  nand ginst21556 (P3_R1158_U493, P3_R1158_U20, P3_U3443);
  not ginst21557 (P3_R1158_U494, P3_R1158_U87);
  nand ginst21558 (P3_R1158_U495, P3_R1158_U178, P3_U3152);
  nand ginst21559 (P3_R1158_U496, P3_R1158_U20, P3_U3906);
  not ginst21560 (P3_R1158_U497, P3_R1158_U89);
  nand ginst21561 (P3_R1158_U498, P3_R1158_U179, P3_U3152);
  nand ginst21562 (P3_R1158_U499, P3_R1158_U20, P3_U3907);
  and ginst21563 (P3_R1158_U5, P3_R1158_U237, P3_R1158_U238);
  nand ginst21564 (P3_R1158_U50, P3_R1158_U85, P3_U3061);
  not ginst21565 (P3_R1158_U500, P3_R1158_U90);
  nand ginst21566 (P3_R1158_U501, P3_R1158_U180, P3_U3152);
  nand ginst21567 (P3_R1158_U502, P3_R1158_U20, P3_U3445);
  not ginst21568 (P3_R1158_U503, P3_R1158_U88);
  nand ginst21569 (P3_R1158_U504, P3_R1158_U181, P3_U3152);
  nand ginst21570 (P3_R1158_U505, P3_R1158_U20, P3_U3905);
  not ginst21571 (P3_R1158_U506, P3_R1158_U91);
  nand ginst21572 (P3_R1158_U507, P3_R1158_U182, P3_U3152);
  nand ginst21573 (P3_R1158_U508, P3_R1158_U20, P3_U3904);
  not ginst21574 (P3_R1158_U509, P3_R1158_U92);
  not ginst21575 (P3_R1158_U51, P3_U3073);
  nand ginst21576 (P3_R1158_U510, P3_R1158_U183, P3_U3152);
  nand ginst21577 (P3_R1158_U511, P3_R1158_U20, P3_U3901);
  not ginst21578 (P3_R1158_U512, P3_R1158_U78);
  nand ginst21579 (P3_R1158_U513, P3_R1158_U184, P3_U3152);
  nand ginst21580 (P3_R1158_U514, P3_R1158_U20, P3_U3902);
  not ginst21581 (P3_R1158_U515, P3_R1158_U76);
  nand ginst21582 (P3_R1158_U516, P3_R1158_U185, P3_U3152);
  nand ginst21583 (P3_R1158_U517, P3_R1158_U20, P3_U3903);
  not ginst21584 (P3_R1158_U518, P3_R1158_U77);
  nand ginst21585 (P3_R1158_U519, P3_R1158_U186, P3_U3152);
  not ginst21586 (P3_R1158_U52, P3_U3081);
  nand ginst21587 (P3_R1158_U520, P3_R1158_U20, P3_U3053);
  not ginst21588 (P3_R1158_U521, P3_R1158_U137);
  nand ginst21589 (P3_R1158_U522, P3_R1158_U521, P3_U3899);
  nand ginst21590 (P3_R1158_U523, P3_R1158_U137, P3_R1158_U187);
  not ginst21591 (P3_R1158_U524, P3_R1158_U93);
  nand ginst21592 (P3_R1158_U525, P3_R1158_U313, P3_R1158_U358, P3_R1158_U524);
  nand ginst21593 (P3_R1158_U526, P3_R1158_U136, P3_R1158_U375, P3_R1158_U93);
  nand ginst21594 (P3_R1158_U527, P3_R1158_U467, P3_U3052);
  nand ginst21595 (P3_R1158_U528, P3_R1158_U37, P3_R1158_U75);
  nand ginst21596 (P3_R1158_U529, P3_R1158_U467, P3_U3052);
  not ginst21597 (P3_R1158_U53, P3_U3075);
  nand ginst21598 (P3_R1158_U530, P3_R1158_U37, P3_R1158_U75);
  nand ginst21599 (P3_R1158_U531, P3_R1158_U529, P3_R1158_U530);
  nand ginst21600 (P3_R1158_U532, P3_R1158_U188, P3_R1158_U189);
  nand ginst21601 (P3_R1158_U533, P3_R1158_U312, P3_R1158_U531);
  nand ginst21602 (P3_R1158_U534, P3_R1158_U512, P3_U3056);
  nand ginst21603 (P3_R1158_U535, P3_R1158_U40, P3_R1158_U78);
  nand ginst21604 (P3_R1158_U536, P3_R1158_U104, P3_R1158_U190);
  nand ginst21605 (P3_R1158_U537, P3_R1158_U103, P3_R1158_U317);
  nand ginst21606 (P3_R1158_U538, P3_R1158_U515, P3_U3057);
  nand ginst21607 (P3_R1158_U539, P3_R1158_U38, P3_R1158_U76);
  not ginst21608 (P3_R1158_U54, P3_U3080);
  nand ginst21609 (P3_R1158_U540, P3_R1158_U538, P3_R1158_U539);
  nand ginst21610 (P3_R1158_U541, P3_R1158_U191, P3_R1158_U349);
  nand ginst21611 (P3_R1158_U542, P3_R1158_U318, P3_R1158_U540);
  nand ginst21612 (P3_R1158_U543, P3_R1158_U518, P3_U3064);
  nand ginst21613 (P3_R1158_U544, P3_R1158_U39, P3_R1158_U77);
  nand ginst21614 (P3_R1158_U545, P3_R1158_U543, P3_R1158_U544);
  nand ginst21615 (P3_R1158_U546, P3_R1158_U192, P3_R1158_U350);
  nand ginst21616 (P3_R1158_U547, P3_R1158_U305, P3_R1158_U545);
  nand ginst21617 (P3_R1158_U548, P3_R1158_U509, P3_U3065);
  nand ginst21618 (P3_R1158_U549, P3_R1158_U58, P3_R1158_U92);
  nand ginst21619 (P3_R1158_U55, P3_R1158_U88, P3_U3080);
  nand ginst21620 (P3_R1158_U550, P3_R1158_U509, P3_U3065);
  nand ginst21621 (P3_R1158_U551, P3_R1158_U58, P3_R1158_U92);
  nand ginst21622 (P3_R1158_U552, P3_R1158_U550, P3_R1158_U551);
  nand ginst21623 (P3_R1158_U553, P3_R1158_U193, P3_R1158_U194);
  nand ginst21624 (P3_R1158_U554, P3_R1158_U301, P3_R1158_U552);
  nand ginst21625 (P3_R1158_U555, P3_R1158_U506, P3_U3060);
  nand ginst21626 (P3_R1158_U556, P3_R1158_U57, P3_R1158_U91);
  nand ginst21627 (P3_R1158_U557, P3_R1158_U506, P3_U3060);
  nand ginst21628 (P3_R1158_U558, P3_R1158_U57, P3_R1158_U91);
  nand ginst21629 (P3_R1158_U559, P3_R1158_U557, P3_R1158_U558);
  not ginst21630 (P3_R1158_U56, P3_U3074);
  nand ginst21631 (P3_R1158_U560, P3_R1158_U195, P3_R1158_U196);
  nand ginst21632 (P3_R1158_U561, P3_R1158_U297, P3_R1158_U559);
  nand ginst21633 (P3_R1158_U562, P3_R1158_U497, P3_U3074);
  nand ginst21634 (P3_R1158_U563, P3_R1158_U56, P3_R1158_U89);
  nand ginst21635 (P3_R1158_U564, P3_R1158_U500, P3_U3075);
  nand ginst21636 (P3_R1158_U565, P3_R1158_U53, P3_R1158_U90);
  nand ginst21637 (P3_R1158_U566, P3_R1158_U564, P3_R1158_U565);
  nand ginst21638 (P3_R1158_U567, P3_R1158_U351, P3_R1158_U61);
  nand ginst21639 (P3_R1158_U568, P3_R1158_U323, P3_R1158_U566);
  nand ginst21640 (P3_R1158_U569, P3_R1158_U406, P3_U3077);
  not ginst21641 (P3_R1158_U57, P3_U3060);
  nand ginst21642 (P3_R1158_U570, P3_R1158_U30, P3_R1158_U72);
  nand ginst21643 (P3_R1158_U571, P3_R1158_U406, P3_U3077);
  nand ginst21644 (P3_R1158_U572, P3_R1158_U30, P3_R1158_U72);
  nand ginst21645 (P3_R1158_U573, P3_R1158_U571, P3_R1158_U572);
  nand ginst21646 (P3_R1158_U574, P3_R1158_U197, P3_R1158_U198);
  nand ginst21647 (P3_R1158_U575, P3_R1158_U222, P3_R1158_U573);
  nand ginst21648 (P3_R1158_U576, P3_R1158_U503, P3_U3080);
  nand ginst21649 (P3_R1158_U577, P3_R1158_U54, P3_R1158_U88);
  nand ginst21650 (P3_R1158_U578, P3_R1158_U576, P3_R1158_U577);
  nand ginst21651 (P3_R1158_U579, P3_R1158_U199, P3_R1158_U352);
  not ginst21652 (P3_R1158_U58, P3_U3065);
  nand ginst21653 (P3_R1158_U580, P3_R1158_U287, P3_R1158_U578);
  nand ginst21654 (P3_R1158_U581, P3_R1158_U494, P3_U3081);
  nand ginst21655 (P3_R1158_U582, P3_R1158_U52, P3_R1158_U87);
  nand ginst21656 (P3_R1158_U583, P3_R1158_U494, P3_U3081);
  nand ginst21657 (P3_R1158_U584, P3_R1158_U52, P3_R1158_U87);
  nand ginst21658 (P3_R1158_U585, P3_R1158_U583, P3_R1158_U584);
  nand ginst21659 (P3_R1158_U586, P3_R1158_U200, P3_R1158_U201);
  nand ginst21660 (P3_R1158_U587, P3_R1158_U283, P3_R1158_U585);
  nand ginst21661 (P3_R1158_U588, P3_R1158_U488, P3_U3068);
  nand ginst21662 (P3_R1158_U589, P3_R1158_U43, P3_R1158_U80);
  nand ginst21663 (P3_R1158_U59, P3_R1158_U76, P3_U3057);
  nand ginst21664 (P3_R1158_U590, P3_R1158_U491, P3_U3072);
  nand ginst21665 (P3_R1158_U591, P3_R1158_U41, P3_R1158_U79);
  nand ginst21666 (P3_R1158_U592, P3_R1158_U590, P3_R1158_U591);
  nand ginst21667 (P3_R1158_U593, P3_R1158_U353, P3_R1158_U62);
  nand ginst21668 (P3_R1158_U594, P3_R1158_U275, P3_R1158_U592);
  nand ginst21669 (P3_R1158_U595, P3_R1158_U485, P3_U3073);
  nand ginst21670 (P3_R1158_U596, P3_R1158_U51, P3_R1158_U86);
  nand ginst21671 (P3_R1158_U597, P3_R1158_U485, P3_U3073);
  nand ginst21672 (P3_R1158_U598, P3_R1158_U51, P3_R1158_U86);
  nand ginst21673 (P3_R1158_U599, P3_R1158_U597, P3_R1158_U598);
  and ginst21674 (P3_R1158_U6, P3_R1158_U262, P3_R1158_U263);
  nand ginst21675 (P3_R1158_U60, P3_R1158_U77, P3_U3064);
  nand ginst21676 (P3_R1158_U600, P3_R1158_U202, P3_R1158_U203);
  nand ginst21677 (P3_R1158_U601, P3_R1158_U390, P3_R1158_U599);
  nand ginst21678 (P3_R1158_U602, P3_R1158_U482, P3_U3078);
  nand ginst21679 (P3_R1158_U603, P3_R1158_U44, P3_R1158_U81);
  nand ginst21680 (P3_R1158_U604, P3_R1158_U482, P3_U3078);
  nand ginst21681 (P3_R1158_U605, P3_R1158_U44, P3_R1158_U81);
  nand ginst21682 (P3_R1158_U606, P3_R1158_U604, P3_R1158_U605);
  nand ginst21683 (P3_R1158_U607, P3_R1158_U204, P3_R1158_U205);
  nand ginst21684 (P3_R1158_U608, P3_R1158_U388, P3_R1158_U606);
  nand ginst21685 (P3_R1158_U609, P3_R1158_U476, P3_U3079);
  nand ginst21686 (P3_R1158_U61, P3_R1158_U322, P3_R1158_U55);
  nand ginst21687 (P3_R1158_U610, P3_R1158_U48, P3_R1158_U83);
  nand ginst21688 (P3_R1158_U611, P3_R1158_U479, P3_U3071);
  nand ginst21689 (P3_R1158_U612, P3_R1158_U45, P3_R1158_U82);
  nand ginst21690 (P3_R1158_U613, P3_R1158_U611, P3_R1158_U612);
  nand ginst21691 (P3_R1158_U614, P3_R1158_U354, P3_R1158_U64);
  nand ginst21692 (P3_R1158_U615, P3_R1158_U339, P3_R1158_U613);
  nand ginst21693 (P3_R1158_U616, P3_R1158_U473, P3_U3062);
  nand ginst21694 (P3_R1158_U617, P3_R1158_U46, P3_R1158_U84);
  nand ginst21695 (P3_R1158_U618, P3_R1158_U616, P3_R1158_U617);
  nand ginst21696 (P3_R1158_U619, P3_R1158_U206, P3_R1158_U355);
  nand ginst21697 (P3_R1158_U62, P3_R1158_U273, P3_R1158_U274);
  nand ginst21698 (P3_R1158_U620, P3_R1158_U386, P3_R1158_U618);
  nand ginst21699 (P3_R1158_U621, P3_R1158_U470, P3_U3061);
  nand ginst21700 (P3_R1158_U622, P3_R1158_U49, P3_R1158_U85);
  nand ginst21701 (P3_R1158_U623, P3_R1158_U470, P3_U3061);
  nand ginst21702 (P3_R1158_U624, P3_R1158_U49, P3_R1158_U85);
  nand ginst21703 (P3_R1158_U625, P3_R1158_U623, P3_R1158_U624);
  nand ginst21704 (P3_R1158_U626, P3_R1158_U207, P3_R1158_U208);
  nand ginst21705 (P3_R1158_U627, P3_R1158_U259, P3_R1158_U625);
  nand ginst21706 (P3_R1158_U628, P3_R1158_U20, P3_R1158_U73);
  nand ginst21707 (P3_R1158_U629, P3_R1158_U409, P3_U3152);
  nand ginst21708 (P3_R1158_U63, P3_R1158_U269, P3_R1158_U365);
  not ginst21709 (P3_R1158_U630, P3_R1158_U149);
  nand ginst21710 (P3_R1158_U631, P3_R1158_U630, P3_U3076);
  nand ginst21711 (P3_R1158_U632, P3_R1158_U149, P3_R1158_U31);
  nand ginst21712 (P3_R1158_U64, P3_R1158_U338, P3_R1158_U47);
  nand ginst21713 (P3_R1158_U65, P3_R1158_U393, P3_R1158_U394);
  nand ginst21714 (P3_R1158_U66, P3_R1158_U425, P3_R1158_U426);
  nand ginst21715 (P3_R1158_U67, P3_R1158_U422, P3_R1158_U423);
  nand ginst21716 (P3_R1158_U68, P3_R1158_U419, P3_R1158_U420);
  nand ginst21717 (P3_R1158_U69, P3_R1158_U416, P3_R1158_U417);
  and ginst21718 (P3_R1158_U7, P3_R1158_U276, P3_R1158_U277);
  nand ginst21719 (P3_R1158_U70, P3_R1158_U413, P3_R1158_U414);
  nand ginst21720 (P3_R1158_U71, P3_R1158_U410, P3_R1158_U411);
  nand ginst21721 (P3_R1158_U72, P3_R1158_U404, P3_R1158_U405);
  nand ginst21722 (P3_R1158_U73, P3_R1158_U407, P3_R1158_U408);
  nand ginst21723 (P3_R1158_U74, P3_R1158_U401, P3_R1158_U402);
  nand ginst21724 (P3_R1158_U75, P3_R1158_U465, P3_R1158_U466);
  nand ginst21725 (P3_R1158_U76, P3_R1158_U513, P3_R1158_U514);
  nand ginst21726 (P3_R1158_U77, P3_R1158_U516, P3_R1158_U517);
  nand ginst21727 (P3_R1158_U78, P3_R1158_U510, P3_R1158_U511);
  nand ginst21728 (P3_R1158_U79, P3_R1158_U489, P3_R1158_U490);
  and ginst21729 (P3_R1158_U8, P3_R1158_U288, P3_R1158_U289);
  nand ginst21730 (P3_R1158_U80, P3_R1158_U486, P3_R1158_U487);
  nand ginst21731 (P3_R1158_U81, P3_R1158_U480, P3_R1158_U481);
  nand ginst21732 (P3_R1158_U82, P3_R1158_U477, P3_R1158_U478);
  nand ginst21733 (P3_R1158_U83, P3_R1158_U474, P3_R1158_U475);
  nand ginst21734 (P3_R1158_U84, P3_R1158_U471, P3_R1158_U472);
  nand ginst21735 (P3_R1158_U85, P3_R1158_U468, P3_R1158_U469);
  nand ginst21736 (P3_R1158_U86, P3_R1158_U483, P3_R1158_U484);
  nand ginst21737 (P3_R1158_U87, P3_R1158_U492, P3_R1158_U493);
  nand ginst21738 (P3_R1158_U88, P3_R1158_U501, P3_R1158_U502);
  nand ginst21739 (P3_R1158_U89, P3_R1158_U495, P3_R1158_U496);
  and ginst21740 (P3_R1158_U9, P3_R1158_U267, P3_R1158_U6);
  nand ginst21741 (P3_R1158_U90, P3_R1158_U498, P3_R1158_U499);
  nand ginst21742 (P3_R1158_U91, P3_R1158_U504, P3_R1158_U505);
  nand ginst21743 (P3_R1158_U92, P3_R1158_U507, P3_R1158_U508);
  nand ginst21744 (P3_R1158_U93, P3_R1158_U522, P3_R1158_U523);
  nand ginst21745 (P3_R1158_U94, P3_R1158_U631, P3_R1158_U632);
  nand ginst21746 (P3_R1158_U95, P3_R1158_U428, P3_R1158_U429);
  nand ginst21747 (P3_R1158_U96, P3_R1158_U435, P3_R1158_U436);
  nand ginst21748 (P3_R1158_U97, P3_R1158_U442, P3_R1158_U443);
  nand ginst21749 (P3_R1158_U98, P3_R1158_U449, P3_R1158_U450);
  nand ginst21750 (P3_R1158_U99, P3_R1158_U456, P3_R1158_U457);
  and ginst21751 (P3_R1161_U10, P3_R1161_U348, P3_R1161_U351);
  nand ginst21752 (P3_R1161_U100, P3_R1161_U398, P3_R1161_U399);
  nand ginst21753 (P3_R1161_U101, P3_R1161_U407, P3_R1161_U408);
  nand ginst21754 (P3_R1161_U102, P3_R1161_U414, P3_R1161_U415);
  nand ginst21755 (P3_R1161_U103, P3_R1161_U421, P3_R1161_U422);
  nand ginst21756 (P3_R1161_U104, P3_R1161_U428, P3_R1161_U429);
  nand ginst21757 (P3_R1161_U105, P3_R1161_U433, P3_R1161_U434);
  nand ginst21758 (P3_R1161_U106, P3_R1161_U440, P3_R1161_U441);
  nand ginst21759 (P3_R1161_U107, P3_R1161_U447, P3_R1161_U448);
  nand ginst21760 (P3_R1161_U108, P3_R1161_U461, P3_R1161_U462);
  nand ginst21761 (P3_R1161_U109, P3_R1161_U466, P3_R1161_U467);
  and ginst21762 (P3_R1161_U11, P3_R1161_U341, P3_R1161_U344);
  nand ginst21763 (P3_R1161_U110, P3_R1161_U473, P3_R1161_U474);
  nand ginst21764 (P3_R1161_U111, P3_R1161_U480, P3_R1161_U481);
  nand ginst21765 (P3_R1161_U112, P3_R1161_U487, P3_R1161_U488);
  nand ginst21766 (P3_R1161_U113, P3_R1161_U494, P3_R1161_U495);
  nand ginst21767 (P3_R1161_U114, P3_R1161_U499, P3_R1161_U500);
  and ginst21768 (P3_R1161_U115, P3_R1161_U187, P3_R1161_U189);
  and ginst21769 (P3_R1161_U116, P3_R1161_U180, P3_R1161_U4);
  and ginst21770 (P3_R1161_U117, P3_R1161_U192, P3_R1161_U194);
  and ginst21771 (P3_R1161_U118, P3_R1161_U200, P3_R1161_U201);
  and ginst21772 (P3_R1161_U119, P3_R1161_U22, P3_R1161_U381, P3_R1161_U382);
  and ginst21773 (P3_R1161_U12, P3_R1161_U332, P3_R1161_U335);
  and ginst21774 (P3_R1161_U120, P3_R1161_U212, P3_R1161_U5);
  and ginst21775 (P3_R1161_U121, P3_R1161_U180, P3_R1161_U181);
  and ginst21776 (P3_R1161_U122, P3_R1161_U218, P3_R1161_U220);
  and ginst21777 (P3_R1161_U123, P3_R1161_U34, P3_R1161_U388, P3_R1161_U389);
  and ginst21778 (P3_R1161_U124, P3_R1161_U226, P3_R1161_U4);
  and ginst21779 (P3_R1161_U125, P3_R1161_U181, P3_R1161_U234);
  and ginst21780 (P3_R1161_U126, P3_R1161_U204, P3_R1161_U6);
  and ginst21781 (P3_R1161_U127, P3_R1161_U239, P3_R1161_U243);
  and ginst21782 (P3_R1161_U128, P3_R1161_U250, P3_R1161_U7);
  and ginst21783 (P3_R1161_U129, P3_R1161_U172, P3_R1161_U248);
  and ginst21784 (P3_R1161_U13, P3_R1161_U323, P3_R1161_U326);
  and ginst21785 (P3_R1161_U130, P3_R1161_U267, P3_R1161_U268);
  and ginst21786 (P3_R1161_U131, P3_R1161_U273, P3_R1161_U282, P3_R1161_U9);
  and ginst21787 (P3_R1161_U132, P3_R1161_U280, P3_R1161_U285);
  and ginst21788 (P3_R1161_U133, P3_R1161_U298, P3_R1161_U301);
  and ginst21789 (P3_R1161_U134, P3_R1161_U302, P3_R1161_U368);
  and ginst21790 (P3_R1161_U135, P3_R1161_U160, P3_R1161_U278);
  and ginst21791 (P3_R1161_U136, P3_R1161_U454, P3_R1161_U455, P3_R1161_U80);
  and ginst21792 (P3_R1161_U137, P3_R1161_U325, P3_R1161_U9);
  and ginst21793 (P3_R1161_U138, P3_R1161_U468, P3_R1161_U469, P3_R1161_U59);
  and ginst21794 (P3_R1161_U139, P3_R1161_U334, P3_R1161_U8);
  and ginst21795 (P3_R1161_U14, P3_R1161_U318, P3_R1161_U320);
  and ginst21796 (P3_R1161_U140, P3_R1161_U172, P3_R1161_U489, P3_R1161_U490);
  and ginst21797 (P3_R1161_U141, P3_R1161_U343, P3_R1161_U7);
  and ginst21798 (P3_R1161_U142, P3_R1161_U171, P3_R1161_U501, P3_R1161_U502);
  and ginst21799 (P3_R1161_U143, P3_R1161_U350, P3_R1161_U6);
  nand ginst21800 (P3_R1161_U144, P3_R1161_U118, P3_R1161_U202);
  nand ginst21801 (P3_R1161_U145, P3_R1161_U217, P3_R1161_U229);
  not ginst21802 (P3_R1161_U146, P3_U3054);
  not ginst21803 (P3_R1161_U147, P3_U3908);
  and ginst21804 (P3_R1161_U148, P3_R1161_U402, P3_R1161_U403);
  nand ginst21805 (P3_R1161_U149, P3_R1161_U169, P3_R1161_U304, P3_R1161_U364);
  and ginst21806 (P3_R1161_U15, P3_R1161_U310, P3_R1161_U313);
  and ginst21807 (P3_R1161_U150, P3_R1161_U409, P3_R1161_U410);
  nand ginst21808 (P3_R1161_U151, P3_R1161_U134, P3_R1161_U369, P3_R1161_U370);
  and ginst21809 (P3_R1161_U152, P3_R1161_U416, P3_R1161_U417);
  nand ginst21810 (P3_R1161_U153, P3_R1161_U299, P3_R1161_U365, P3_R1161_U86);
  and ginst21811 (P3_R1161_U154, P3_R1161_U423, P3_R1161_U424);
  nand ginst21812 (P3_R1161_U155, P3_R1161_U292, P3_R1161_U293);
  and ginst21813 (P3_R1161_U156, P3_R1161_U435, P3_R1161_U436);
  nand ginst21814 (P3_R1161_U157, P3_R1161_U288, P3_R1161_U289);
  and ginst21815 (P3_R1161_U158, P3_R1161_U442, P3_R1161_U443);
  nand ginst21816 (P3_R1161_U159, P3_R1161_U132, P3_R1161_U284);
  and ginst21817 (P3_R1161_U16, P3_R1161_U232, P3_R1161_U235);
  and ginst21818 (P3_R1161_U160, P3_R1161_U449, P3_R1161_U450);
  nand ginst21819 (P3_R1161_U161, P3_R1161_U327, P3_R1161_U43);
  nand ginst21820 (P3_R1161_U162, P3_R1161_U130, P3_R1161_U269);
  and ginst21821 (P3_R1161_U163, P3_R1161_U475, P3_R1161_U476);
  nand ginst21822 (P3_R1161_U164, P3_R1161_U256, P3_R1161_U257);
  and ginst21823 (P3_R1161_U165, P3_R1161_U482, P3_R1161_U483);
  nand ginst21824 (P3_R1161_U166, P3_R1161_U252, P3_R1161_U253);
  nand ginst21825 (P3_R1161_U167, P3_R1161_U127, P3_R1161_U242);
  nand ginst21826 (P3_R1161_U168, P3_R1161_U366, P3_R1161_U367);
  nand ginst21827 (P3_R1161_U169, P3_R1161_U151, P3_U3053);
  and ginst21828 (P3_R1161_U17, P3_R1161_U224, P3_R1161_U227);
  not ginst21829 (P3_R1161_U170, P3_R1161_U34);
  nand ginst21830 (P3_R1161_U171, P3_U3082, P3_U3416);
  nand ginst21831 (P3_R1161_U172, P3_U3071, P3_U3425);
  nand ginst21832 (P3_R1161_U173, P3_U3057, P3_U3902);
  not ginst21833 (P3_R1161_U174, P3_R1161_U68);
  not ginst21834 (P3_R1161_U175, P3_R1161_U77);
  nand ginst21835 (P3_R1161_U176, P3_U3064, P3_U3903);
  not ginst21836 (P3_R1161_U177, P3_R1161_U63);
  or ginst21837 (P3_R1161_U178, P3_U3066, P3_U3404);
  or ginst21838 (P3_R1161_U179, P3_U3059, P3_U3401);
  and ginst21839 (P3_R1161_U18, P3_R1161_U210, P3_R1161_U213);
  or ginst21840 (P3_R1161_U180, P3_U3063, P3_U3398);
  or ginst21841 (P3_R1161_U181, P3_U3067, P3_U3395);
  not ginst21842 (P3_R1161_U182, P3_R1161_U31);
  or ginst21843 (P3_R1161_U183, P3_U3077, P3_U3392);
  not ginst21844 (P3_R1161_U184, P3_R1161_U42);
  not ginst21845 (P3_R1161_U185, P3_R1161_U43);
  nand ginst21846 (P3_R1161_U186, P3_R1161_U42, P3_R1161_U43);
  nand ginst21847 (P3_R1161_U187, P3_U3067, P3_U3395);
  nand ginst21848 (P3_R1161_U188, P3_R1161_U181, P3_R1161_U186);
  nand ginst21849 (P3_R1161_U189, P3_U3063, P3_U3398);
  not ginst21850 (P3_R1161_U19, P3_U3407);
  nand ginst21851 (P3_R1161_U190, P3_R1161_U115, P3_R1161_U188);
  nand ginst21852 (P3_R1161_U191, P3_R1161_U34, P3_R1161_U35);
  nand ginst21853 (P3_R1161_U192, P3_R1161_U191, P3_U3066);
  nand ginst21854 (P3_R1161_U193, P3_R1161_U116, P3_R1161_U190);
  nand ginst21855 (P3_R1161_U194, P3_R1161_U170, P3_U3404);
  not ginst21856 (P3_R1161_U195, P3_R1161_U41);
  or ginst21857 (P3_R1161_U196, P3_U3069, P3_U3410);
  or ginst21858 (P3_R1161_U197, P3_U3070, P3_U3407);
  not ginst21859 (P3_R1161_U198, P3_R1161_U22);
  nand ginst21860 (P3_R1161_U199, P3_R1161_U22, P3_R1161_U23);
  not ginst21861 (P3_R1161_U20, P3_U3070);
  nand ginst21862 (P3_R1161_U200, P3_R1161_U199, P3_U3069);
  nand ginst21863 (P3_R1161_U201, P3_R1161_U198, P3_U3410);
  nand ginst21864 (P3_R1161_U202, P3_R1161_U41, P3_R1161_U5);
  not ginst21865 (P3_R1161_U203, P3_R1161_U144);
  or ginst21866 (P3_R1161_U204, P3_U3083, P3_U3413);
  nand ginst21867 (P3_R1161_U205, P3_R1161_U144, P3_R1161_U204);
  not ginst21868 (P3_R1161_U206, P3_R1161_U40);
  or ginst21869 (P3_R1161_U207, P3_U3082, P3_U3416);
  or ginst21870 (P3_R1161_U208, P3_U3070, P3_U3407);
  nand ginst21871 (P3_R1161_U209, P3_R1161_U208, P3_R1161_U41);
  not ginst21872 (P3_R1161_U21, P3_U3069);
  nand ginst21873 (P3_R1161_U210, P3_R1161_U119, P3_R1161_U209);
  nand ginst21874 (P3_R1161_U211, P3_R1161_U195, P3_R1161_U22);
  nand ginst21875 (P3_R1161_U212, P3_U3069, P3_U3410);
  nand ginst21876 (P3_R1161_U213, P3_R1161_U120, P3_R1161_U211);
  or ginst21877 (P3_R1161_U214, P3_U3070, P3_U3407);
  nand ginst21878 (P3_R1161_U215, P3_R1161_U181, P3_R1161_U185);
  nand ginst21879 (P3_R1161_U216, P3_U3067, P3_U3395);
  not ginst21880 (P3_R1161_U217, P3_R1161_U45);
  nand ginst21881 (P3_R1161_U218, P3_R1161_U121, P3_R1161_U184);
  nand ginst21882 (P3_R1161_U219, P3_R1161_U180, P3_R1161_U45);
  nand ginst21883 (P3_R1161_U22, P3_U3070, P3_U3407);
  nand ginst21884 (P3_R1161_U220, P3_U3063, P3_U3398);
  not ginst21885 (P3_R1161_U221, P3_R1161_U44);
  or ginst21886 (P3_R1161_U222, P3_U3059, P3_U3401);
  nand ginst21887 (P3_R1161_U223, P3_R1161_U222, P3_R1161_U44);
  nand ginst21888 (P3_R1161_U224, P3_R1161_U123, P3_R1161_U223);
  nand ginst21889 (P3_R1161_U225, P3_R1161_U221, P3_R1161_U34);
  nand ginst21890 (P3_R1161_U226, P3_U3066, P3_U3404);
  nand ginst21891 (P3_R1161_U227, P3_R1161_U124, P3_R1161_U225);
  or ginst21892 (P3_R1161_U228, P3_U3059, P3_U3401);
  nand ginst21893 (P3_R1161_U229, P3_R1161_U181, P3_R1161_U184);
  not ginst21894 (P3_R1161_U23, P3_U3410);
  not ginst21895 (P3_R1161_U230, P3_R1161_U145);
  nand ginst21896 (P3_R1161_U231, P3_U3063, P3_U3398);
  nand ginst21897 (P3_R1161_U232, P3_R1161_U400, P3_R1161_U401, P3_R1161_U42, P3_R1161_U43);
  nand ginst21898 (P3_R1161_U233, P3_R1161_U42, P3_R1161_U43);
  nand ginst21899 (P3_R1161_U234, P3_U3067, P3_U3395);
  nand ginst21900 (P3_R1161_U235, P3_R1161_U125, P3_R1161_U233);
  or ginst21901 (P3_R1161_U236, P3_U3082, P3_U3416);
  or ginst21902 (P3_R1161_U237, P3_U3061, P3_U3419);
  nand ginst21903 (P3_R1161_U238, P3_R1161_U177, P3_R1161_U6);
  nand ginst21904 (P3_R1161_U239, P3_U3061, P3_U3419);
  not ginst21905 (P3_R1161_U24, P3_U3401);
  nand ginst21906 (P3_R1161_U240, P3_R1161_U171, P3_R1161_U238);
  or ginst21907 (P3_R1161_U241, P3_U3061, P3_U3419);
  nand ginst21908 (P3_R1161_U242, P3_R1161_U126, P3_R1161_U144);
  nand ginst21909 (P3_R1161_U243, P3_R1161_U240, P3_R1161_U241);
  not ginst21910 (P3_R1161_U244, P3_R1161_U167);
  or ginst21911 (P3_R1161_U245, P3_U3079, P3_U3428);
  or ginst21912 (P3_R1161_U246, P3_U3071, P3_U3425);
  nand ginst21913 (P3_R1161_U247, P3_R1161_U174, P3_R1161_U7);
  nand ginst21914 (P3_R1161_U248, P3_U3079, P3_U3428);
  nand ginst21915 (P3_R1161_U249, P3_R1161_U129, P3_R1161_U247);
  not ginst21916 (P3_R1161_U25, P3_U3059);
  or ginst21917 (P3_R1161_U250, P3_U3062, P3_U3422);
  or ginst21918 (P3_R1161_U251, P3_U3079, P3_U3428);
  nand ginst21919 (P3_R1161_U252, P3_R1161_U128, P3_R1161_U167);
  nand ginst21920 (P3_R1161_U253, P3_R1161_U249, P3_R1161_U251);
  not ginst21921 (P3_R1161_U254, P3_R1161_U166);
  or ginst21922 (P3_R1161_U255, P3_U3078, P3_U3431);
  nand ginst21923 (P3_R1161_U256, P3_R1161_U166, P3_R1161_U255);
  nand ginst21924 (P3_R1161_U257, P3_U3078, P3_U3431);
  not ginst21925 (P3_R1161_U258, P3_R1161_U164);
  or ginst21926 (P3_R1161_U259, P3_U3073, P3_U3434);
  not ginst21927 (P3_R1161_U26, P3_U3066);
  nand ginst21928 (P3_R1161_U260, P3_R1161_U164, P3_R1161_U259);
  nand ginst21929 (P3_R1161_U261, P3_U3073, P3_U3434);
  not ginst21930 (P3_R1161_U262, P3_R1161_U92);
  or ginst21931 (P3_R1161_U263, P3_U3068, P3_U3440);
  or ginst21932 (P3_R1161_U264, P3_U3072, P3_U3437);
  not ginst21933 (P3_R1161_U265, P3_R1161_U59);
  nand ginst21934 (P3_R1161_U266, P3_R1161_U59, P3_R1161_U60);
  nand ginst21935 (P3_R1161_U267, P3_R1161_U266, P3_U3068);
  nand ginst21936 (P3_R1161_U268, P3_R1161_U265, P3_U3440);
  nand ginst21937 (P3_R1161_U269, P3_R1161_U8, P3_R1161_U92);
  not ginst21938 (P3_R1161_U27, P3_U3395);
  not ginst21939 (P3_R1161_U270, P3_R1161_U162);
  or ginst21940 (P3_R1161_U271, P3_U3075, P3_U3907);
  or ginst21941 (P3_R1161_U272, P3_U3080, P3_U3445);
  or ginst21942 (P3_R1161_U273, P3_U3074, P3_U3906);
  not ginst21943 (P3_R1161_U274, P3_R1161_U80);
  nand ginst21944 (P3_R1161_U275, P3_R1161_U274, P3_U3907);
  nand ginst21945 (P3_R1161_U276, P3_R1161_U275, P3_R1161_U90);
  nand ginst21946 (P3_R1161_U277, P3_R1161_U80, P3_R1161_U81);
  nand ginst21947 (P3_R1161_U278, P3_R1161_U276, P3_R1161_U277);
  nand ginst21948 (P3_R1161_U279, P3_R1161_U175, P3_R1161_U9);
  not ginst21949 (P3_R1161_U28, P3_U3067);
  nand ginst21950 (P3_R1161_U280, P3_U3074, P3_U3906);
  nand ginst21951 (P3_R1161_U281, P3_R1161_U278, P3_R1161_U279);
  or ginst21952 (P3_R1161_U282, P3_U3081, P3_U3443);
  or ginst21953 (P3_R1161_U283, P3_U3074, P3_U3906);
  nand ginst21954 (P3_R1161_U284, P3_R1161_U131, P3_R1161_U162);
  nand ginst21955 (P3_R1161_U285, P3_R1161_U281, P3_R1161_U283);
  not ginst21956 (P3_R1161_U286, P3_R1161_U159);
  or ginst21957 (P3_R1161_U287, P3_U3060, P3_U3905);
  nand ginst21958 (P3_R1161_U288, P3_R1161_U159, P3_R1161_U287);
  nand ginst21959 (P3_R1161_U289, P3_U3060, P3_U3905);
  not ginst21960 (P3_R1161_U29, P3_U3387);
  not ginst21961 (P3_R1161_U290, P3_R1161_U157);
  or ginst21962 (P3_R1161_U291, P3_U3065, P3_U3904);
  nand ginst21963 (P3_R1161_U292, P3_R1161_U157, P3_R1161_U291);
  nand ginst21964 (P3_R1161_U293, P3_U3065, P3_U3904);
  not ginst21965 (P3_R1161_U294, P3_R1161_U155);
  or ginst21966 (P3_R1161_U295, P3_U3057, P3_U3902);
  nand ginst21967 (P3_R1161_U296, P3_R1161_U173, P3_R1161_U176);
  not ginst21968 (P3_R1161_U297, P3_R1161_U86);
  or ginst21969 (P3_R1161_U298, P3_U3064, P3_U3903);
  nand ginst21970 (P3_R1161_U299, P3_R1161_U155, P3_R1161_U168, P3_R1161_U298);
  not ginst21971 (P3_R1161_U30, P3_U3076);
  not ginst21972 (P3_R1161_U300, P3_R1161_U153);
  or ginst21973 (P3_R1161_U301, P3_U3052, P3_U3900);
  nand ginst21974 (P3_R1161_U302, P3_U3052, P3_U3900);
  not ginst21975 (P3_R1161_U303, P3_R1161_U151);
  nand ginst21976 (P3_R1161_U304, P3_R1161_U151, P3_U3899);
  not ginst21977 (P3_R1161_U305, P3_R1161_U149);
  nand ginst21978 (P3_R1161_U306, P3_R1161_U155, P3_R1161_U298);
  not ginst21979 (P3_R1161_U307, P3_R1161_U89);
  or ginst21980 (P3_R1161_U308, P3_U3057, P3_U3902);
  nand ginst21981 (P3_R1161_U309, P3_R1161_U308, P3_R1161_U89);
  nand ginst21982 (P3_R1161_U31, P3_U3076, P3_U3387);
  nand ginst21983 (P3_R1161_U310, P3_R1161_U154, P3_R1161_U173, P3_R1161_U309);
  nand ginst21984 (P3_R1161_U311, P3_R1161_U173, P3_R1161_U307);
  nand ginst21985 (P3_R1161_U312, P3_U3056, P3_U3901);
  nand ginst21986 (P3_R1161_U313, P3_R1161_U168, P3_R1161_U311, P3_R1161_U312);
  or ginst21987 (P3_R1161_U314, P3_U3057, P3_U3902);
  nand ginst21988 (P3_R1161_U315, P3_R1161_U162, P3_R1161_U282);
  not ginst21989 (P3_R1161_U316, P3_R1161_U91);
  nand ginst21990 (P3_R1161_U317, P3_R1161_U9, P3_R1161_U91);
  nand ginst21991 (P3_R1161_U318, P3_R1161_U135, P3_R1161_U317);
  nand ginst21992 (P3_R1161_U319, P3_R1161_U278, P3_R1161_U317);
  not ginst21993 (P3_R1161_U32, P3_U3398);
  nand ginst21994 (P3_R1161_U320, P3_R1161_U319, P3_R1161_U453);
  or ginst21995 (P3_R1161_U321, P3_U3080, P3_U3445);
  nand ginst21996 (P3_R1161_U322, P3_R1161_U321, P3_R1161_U91);
  nand ginst21997 (P3_R1161_U323, P3_R1161_U136, P3_R1161_U322);
  nand ginst21998 (P3_R1161_U324, P3_R1161_U316, P3_R1161_U80);
  nand ginst21999 (P3_R1161_U325, P3_U3075, P3_U3907);
  nand ginst22000 (P3_R1161_U326, P3_R1161_U137, P3_R1161_U324);
  or ginst22001 (P3_R1161_U327, P3_U3077, P3_U3392);
  not ginst22002 (P3_R1161_U328, P3_R1161_U161);
  or ginst22003 (P3_R1161_U329, P3_U3080, P3_U3445);
  not ginst22004 (P3_R1161_U33, P3_U3063);
  or ginst22005 (P3_R1161_U330, P3_U3072, P3_U3437);
  nand ginst22006 (P3_R1161_U331, P3_R1161_U330, P3_R1161_U92);
  nand ginst22007 (P3_R1161_U332, P3_R1161_U138, P3_R1161_U331);
  nand ginst22008 (P3_R1161_U333, P3_R1161_U262, P3_R1161_U59);
  nand ginst22009 (P3_R1161_U334, P3_U3068, P3_U3440);
  nand ginst22010 (P3_R1161_U335, P3_R1161_U139, P3_R1161_U333);
  or ginst22011 (P3_R1161_U336, P3_U3072, P3_U3437);
  nand ginst22012 (P3_R1161_U337, P3_R1161_U167, P3_R1161_U250);
  not ginst22013 (P3_R1161_U338, P3_R1161_U93);
  or ginst22014 (P3_R1161_U339, P3_U3071, P3_U3425);
  nand ginst22015 (P3_R1161_U34, P3_U3059, P3_U3401);
  nand ginst22016 (P3_R1161_U340, P3_R1161_U339, P3_R1161_U93);
  nand ginst22017 (P3_R1161_U341, P3_R1161_U140, P3_R1161_U340);
  nand ginst22018 (P3_R1161_U342, P3_R1161_U172, P3_R1161_U338);
  nand ginst22019 (P3_R1161_U343, P3_U3079, P3_U3428);
  nand ginst22020 (P3_R1161_U344, P3_R1161_U141, P3_R1161_U342);
  or ginst22021 (P3_R1161_U345, P3_U3071, P3_U3425);
  or ginst22022 (P3_R1161_U346, P3_U3082, P3_U3416);
  nand ginst22023 (P3_R1161_U347, P3_R1161_U346, P3_R1161_U40);
  nand ginst22024 (P3_R1161_U348, P3_R1161_U142, P3_R1161_U347);
  nand ginst22025 (P3_R1161_U349, P3_R1161_U171, P3_R1161_U206);
  not ginst22026 (P3_R1161_U35, P3_U3404);
  nand ginst22027 (P3_R1161_U350, P3_U3061, P3_U3419);
  nand ginst22028 (P3_R1161_U351, P3_R1161_U143, P3_R1161_U349);
  nand ginst22029 (P3_R1161_U352, P3_R1161_U171, P3_R1161_U207);
  nand ginst22030 (P3_R1161_U353, P3_R1161_U204, P3_R1161_U63);
  nand ginst22031 (P3_R1161_U354, P3_R1161_U214, P3_R1161_U22);
  nand ginst22032 (P3_R1161_U355, P3_R1161_U228, P3_R1161_U34);
  nand ginst22033 (P3_R1161_U356, P3_R1161_U180, P3_R1161_U231);
  nand ginst22034 (P3_R1161_U357, P3_R1161_U173, P3_R1161_U314);
  nand ginst22035 (P3_R1161_U358, P3_R1161_U176, P3_R1161_U298);
  nand ginst22036 (P3_R1161_U359, P3_R1161_U329, P3_R1161_U80);
  not ginst22037 (P3_R1161_U36, P3_U3413);
  nand ginst22038 (P3_R1161_U360, P3_R1161_U282, P3_R1161_U77);
  nand ginst22039 (P3_R1161_U361, P3_R1161_U336, P3_R1161_U59);
  nand ginst22040 (P3_R1161_U362, P3_R1161_U172, P3_R1161_U345);
  nand ginst22041 (P3_R1161_U363, P3_R1161_U250, P3_R1161_U68);
  nand ginst22042 (P3_R1161_U364, P3_U3053, P3_U3899);
  nand ginst22043 (P3_R1161_U365, P3_R1161_U168, P3_R1161_U296);
  nand ginst22044 (P3_R1161_U366, P3_R1161_U295, P3_U3056);
  nand ginst22045 (P3_R1161_U367, P3_R1161_U295, P3_U3901);
  nand ginst22046 (P3_R1161_U368, P3_R1161_U168, P3_R1161_U296, P3_R1161_U301);
  nand ginst22047 (P3_R1161_U369, P3_R1161_U133, P3_R1161_U155, P3_R1161_U168);
  not ginst22048 (P3_R1161_U37, P3_U3083);
  nand ginst22049 (P3_R1161_U370, P3_R1161_U297, P3_R1161_U301);
  nand ginst22050 (P3_R1161_U371, P3_R1161_U39, P3_U3082);
  nand ginst22051 (P3_R1161_U372, P3_R1161_U38, P3_U3416);
  nand ginst22052 (P3_R1161_U373, P3_R1161_U371, P3_R1161_U372);
  nand ginst22053 (P3_R1161_U374, P3_R1161_U352, P3_R1161_U40);
  nand ginst22054 (P3_R1161_U375, P3_R1161_U206, P3_R1161_U373);
  nand ginst22055 (P3_R1161_U376, P3_R1161_U36, P3_U3083);
  nand ginst22056 (P3_R1161_U377, P3_R1161_U37, P3_U3413);
  nand ginst22057 (P3_R1161_U378, P3_R1161_U376, P3_R1161_U377);
  nand ginst22058 (P3_R1161_U379, P3_R1161_U144, P3_R1161_U353);
  not ginst22059 (P3_R1161_U38, P3_U3082);
  nand ginst22060 (P3_R1161_U380, P3_R1161_U203, P3_R1161_U378);
  nand ginst22061 (P3_R1161_U381, P3_R1161_U23, P3_U3069);
  nand ginst22062 (P3_R1161_U382, P3_R1161_U21, P3_U3410);
  nand ginst22063 (P3_R1161_U383, P3_R1161_U19, P3_U3070);
  nand ginst22064 (P3_R1161_U384, P3_R1161_U20, P3_U3407);
  nand ginst22065 (P3_R1161_U385, P3_R1161_U383, P3_R1161_U384);
  nand ginst22066 (P3_R1161_U386, P3_R1161_U354, P3_R1161_U41);
  nand ginst22067 (P3_R1161_U387, P3_R1161_U195, P3_R1161_U385);
  nand ginst22068 (P3_R1161_U388, P3_R1161_U35, P3_U3066);
  nand ginst22069 (P3_R1161_U389, P3_R1161_U26, P3_U3404);
  not ginst22070 (P3_R1161_U39, P3_U3416);
  nand ginst22071 (P3_R1161_U390, P3_R1161_U24, P3_U3059);
  nand ginst22072 (P3_R1161_U391, P3_R1161_U25, P3_U3401);
  nand ginst22073 (P3_R1161_U392, P3_R1161_U390, P3_R1161_U391);
  nand ginst22074 (P3_R1161_U393, P3_R1161_U355, P3_R1161_U44);
  nand ginst22075 (P3_R1161_U394, P3_R1161_U221, P3_R1161_U392);
  nand ginst22076 (P3_R1161_U395, P3_R1161_U32, P3_U3063);
  nand ginst22077 (P3_R1161_U396, P3_R1161_U33, P3_U3398);
  nand ginst22078 (P3_R1161_U397, P3_R1161_U395, P3_R1161_U396);
  nand ginst22079 (P3_R1161_U398, P3_R1161_U145, P3_R1161_U356);
  nand ginst22080 (P3_R1161_U399, P3_R1161_U230, P3_R1161_U397);
  and ginst22081 (P3_R1161_U4, P3_R1161_U178, P3_R1161_U179);
  nand ginst22082 (P3_R1161_U40, P3_R1161_U205, P3_R1161_U63);
  nand ginst22083 (P3_R1161_U400, P3_R1161_U27, P3_U3067);
  nand ginst22084 (P3_R1161_U401, P3_R1161_U28, P3_U3395);
  nand ginst22085 (P3_R1161_U402, P3_R1161_U147, P3_U3054);
  nand ginst22086 (P3_R1161_U403, P3_R1161_U146, P3_U3908);
  nand ginst22087 (P3_R1161_U404, P3_R1161_U147, P3_U3054);
  nand ginst22088 (P3_R1161_U405, P3_R1161_U146, P3_U3908);
  nand ginst22089 (P3_R1161_U406, P3_R1161_U404, P3_R1161_U405);
  nand ginst22090 (P3_R1161_U407, P3_R1161_U148, P3_R1161_U149);
  nand ginst22091 (P3_R1161_U408, P3_R1161_U305, P3_R1161_U406);
  nand ginst22092 (P3_R1161_U409, P3_R1161_U88, P3_U3053);
  nand ginst22093 (P3_R1161_U41, P3_R1161_U117, P3_R1161_U193);
  nand ginst22094 (P3_R1161_U410, P3_R1161_U87, P3_U3899);
  nand ginst22095 (P3_R1161_U411, P3_R1161_U88, P3_U3053);
  nand ginst22096 (P3_R1161_U412, P3_R1161_U87, P3_U3899);
  nand ginst22097 (P3_R1161_U413, P3_R1161_U411, P3_R1161_U412);
  nand ginst22098 (P3_R1161_U414, P3_R1161_U150, P3_R1161_U151);
  nand ginst22099 (P3_R1161_U415, P3_R1161_U303, P3_R1161_U413);
  nand ginst22100 (P3_R1161_U416, P3_R1161_U46, P3_U3052);
  nand ginst22101 (P3_R1161_U417, P3_R1161_U47, P3_U3900);
  nand ginst22102 (P3_R1161_U418, P3_R1161_U46, P3_U3052);
  nand ginst22103 (P3_R1161_U419, P3_R1161_U47, P3_U3900);
  nand ginst22104 (P3_R1161_U42, P3_R1161_U182, P3_R1161_U183);
  nand ginst22105 (P3_R1161_U420, P3_R1161_U418, P3_R1161_U419);
  nand ginst22106 (P3_R1161_U421, P3_R1161_U152, P3_R1161_U153);
  nand ginst22107 (P3_R1161_U422, P3_R1161_U300, P3_R1161_U420);
  nand ginst22108 (P3_R1161_U423, P3_R1161_U49, P3_U3056);
  nand ginst22109 (P3_R1161_U424, P3_R1161_U48, P3_U3901);
  nand ginst22110 (P3_R1161_U425, P3_R1161_U50, P3_U3057);
  nand ginst22111 (P3_R1161_U426, P3_R1161_U51, P3_U3902);
  nand ginst22112 (P3_R1161_U427, P3_R1161_U425, P3_R1161_U426);
  nand ginst22113 (P3_R1161_U428, P3_R1161_U357, P3_R1161_U89);
  nand ginst22114 (P3_R1161_U429, P3_R1161_U307, P3_R1161_U427);
  nand ginst22115 (P3_R1161_U43, P3_U3077, P3_U3392);
  nand ginst22116 (P3_R1161_U430, P3_R1161_U52, P3_U3064);
  nand ginst22117 (P3_R1161_U431, P3_R1161_U53, P3_U3903);
  nand ginst22118 (P3_R1161_U432, P3_R1161_U430, P3_R1161_U431);
  nand ginst22119 (P3_R1161_U433, P3_R1161_U155, P3_R1161_U358);
  nand ginst22120 (P3_R1161_U434, P3_R1161_U294, P3_R1161_U432);
  nand ginst22121 (P3_R1161_U435, P3_R1161_U84, P3_U3065);
  nand ginst22122 (P3_R1161_U436, P3_R1161_U85, P3_U3904);
  nand ginst22123 (P3_R1161_U437, P3_R1161_U84, P3_U3065);
  nand ginst22124 (P3_R1161_U438, P3_R1161_U85, P3_U3904);
  nand ginst22125 (P3_R1161_U439, P3_R1161_U437, P3_R1161_U438);
  nand ginst22126 (P3_R1161_U44, P3_R1161_U122, P3_R1161_U219);
  nand ginst22127 (P3_R1161_U440, P3_R1161_U156, P3_R1161_U157);
  nand ginst22128 (P3_R1161_U441, P3_R1161_U290, P3_R1161_U439);
  nand ginst22129 (P3_R1161_U442, P3_R1161_U82, P3_U3060);
  nand ginst22130 (P3_R1161_U443, P3_R1161_U83, P3_U3905);
  nand ginst22131 (P3_R1161_U444, P3_R1161_U82, P3_U3060);
  nand ginst22132 (P3_R1161_U445, P3_R1161_U83, P3_U3905);
  nand ginst22133 (P3_R1161_U446, P3_R1161_U444, P3_R1161_U445);
  nand ginst22134 (P3_R1161_U447, P3_R1161_U158, P3_R1161_U159);
  nand ginst22135 (P3_R1161_U448, P3_R1161_U286, P3_R1161_U446);
  nand ginst22136 (P3_R1161_U449, P3_R1161_U54, P3_U3074);
  nand ginst22137 (P3_R1161_U45, P3_R1161_U215, P3_R1161_U216);
  nand ginst22138 (P3_R1161_U450, P3_R1161_U55, P3_U3906);
  nand ginst22139 (P3_R1161_U451, P3_R1161_U54, P3_U3074);
  nand ginst22140 (P3_R1161_U452, P3_R1161_U55, P3_U3906);
  nand ginst22141 (P3_R1161_U453, P3_R1161_U451, P3_R1161_U452);
  nand ginst22142 (P3_R1161_U454, P3_R1161_U81, P3_U3075);
  nand ginst22143 (P3_R1161_U455, P3_R1161_U90, P3_U3907);
  nand ginst22144 (P3_R1161_U456, P3_R1161_U161, P3_R1161_U182);
  nand ginst22145 (P3_R1161_U457, P3_R1161_U31, P3_R1161_U328);
  nand ginst22146 (P3_R1161_U458, P3_R1161_U78, P3_U3080);
  nand ginst22147 (P3_R1161_U459, P3_R1161_U79, P3_U3445);
  not ginst22148 (P3_R1161_U46, P3_U3900);
  nand ginst22149 (P3_R1161_U460, P3_R1161_U458, P3_R1161_U459);
  nand ginst22150 (P3_R1161_U461, P3_R1161_U359, P3_R1161_U91);
  nand ginst22151 (P3_R1161_U462, P3_R1161_U316, P3_R1161_U460);
  nand ginst22152 (P3_R1161_U463, P3_R1161_U75, P3_U3081);
  nand ginst22153 (P3_R1161_U464, P3_R1161_U76, P3_U3443);
  nand ginst22154 (P3_R1161_U465, P3_R1161_U463, P3_R1161_U464);
  nand ginst22155 (P3_R1161_U466, P3_R1161_U162, P3_R1161_U360);
  nand ginst22156 (P3_R1161_U467, P3_R1161_U270, P3_R1161_U465);
  nand ginst22157 (P3_R1161_U468, P3_R1161_U60, P3_U3068);
  nand ginst22158 (P3_R1161_U469, P3_R1161_U58, P3_U3440);
  not ginst22159 (P3_R1161_U47, P3_U3052);
  nand ginst22160 (P3_R1161_U470, P3_R1161_U56, P3_U3072);
  nand ginst22161 (P3_R1161_U471, P3_R1161_U57, P3_U3437);
  nand ginst22162 (P3_R1161_U472, P3_R1161_U470, P3_R1161_U471);
  nand ginst22163 (P3_R1161_U473, P3_R1161_U361, P3_R1161_U92);
  nand ginst22164 (P3_R1161_U474, P3_R1161_U262, P3_R1161_U472);
  nand ginst22165 (P3_R1161_U475, P3_R1161_U73, P3_U3073);
  nand ginst22166 (P3_R1161_U476, P3_R1161_U74, P3_U3434);
  nand ginst22167 (P3_R1161_U477, P3_R1161_U73, P3_U3073);
  nand ginst22168 (P3_R1161_U478, P3_R1161_U74, P3_U3434);
  nand ginst22169 (P3_R1161_U479, P3_R1161_U477, P3_R1161_U478);
  not ginst22170 (P3_R1161_U48, P3_U3056);
  nand ginst22171 (P3_R1161_U480, P3_R1161_U163, P3_R1161_U164);
  nand ginst22172 (P3_R1161_U481, P3_R1161_U258, P3_R1161_U479);
  nand ginst22173 (P3_R1161_U482, P3_R1161_U71, P3_U3078);
  nand ginst22174 (P3_R1161_U483, P3_R1161_U72, P3_U3431);
  nand ginst22175 (P3_R1161_U484, P3_R1161_U71, P3_U3078);
  nand ginst22176 (P3_R1161_U485, P3_R1161_U72, P3_U3431);
  nand ginst22177 (P3_R1161_U486, P3_R1161_U484, P3_R1161_U485);
  nand ginst22178 (P3_R1161_U487, P3_R1161_U165, P3_R1161_U166);
  nand ginst22179 (P3_R1161_U488, P3_R1161_U254, P3_R1161_U486);
  nand ginst22180 (P3_R1161_U489, P3_R1161_U69, P3_U3079);
  not ginst22181 (P3_R1161_U49, P3_U3901);
  nand ginst22182 (P3_R1161_U490, P3_R1161_U70, P3_U3428);
  nand ginst22183 (P3_R1161_U491, P3_R1161_U64, P3_U3071);
  nand ginst22184 (P3_R1161_U492, P3_R1161_U65, P3_U3425);
  nand ginst22185 (P3_R1161_U493, P3_R1161_U491, P3_R1161_U492);
  nand ginst22186 (P3_R1161_U494, P3_R1161_U362, P3_R1161_U93);
  nand ginst22187 (P3_R1161_U495, P3_R1161_U338, P3_R1161_U493);
  nand ginst22188 (P3_R1161_U496, P3_R1161_U66, P3_U3062);
  nand ginst22189 (P3_R1161_U497, P3_R1161_U67, P3_U3422);
  nand ginst22190 (P3_R1161_U498, P3_R1161_U496, P3_R1161_U497);
  nand ginst22191 (P3_R1161_U499, P3_R1161_U167, P3_R1161_U363);
  and ginst22192 (P3_R1161_U5, P3_R1161_U196, P3_R1161_U197);
  not ginst22193 (P3_R1161_U50, P3_U3902);
  nand ginst22194 (P3_R1161_U500, P3_R1161_U244, P3_R1161_U498);
  nand ginst22195 (P3_R1161_U501, P3_R1161_U61, P3_U3061);
  nand ginst22196 (P3_R1161_U502, P3_R1161_U62, P3_U3419);
  nand ginst22197 (P3_R1161_U503, P3_R1161_U29, P3_U3076);
  nand ginst22198 (P3_R1161_U504, P3_R1161_U30, P3_U3387);
  not ginst22199 (P3_R1161_U51, P3_U3057);
  not ginst22200 (P3_R1161_U52, P3_U3903);
  not ginst22201 (P3_R1161_U53, P3_U3064);
  not ginst22202 (P3_R1161_U54, P3_U3906);
  not ginst22203 (P3_R1161_U55, P3_U3074);
  not ginst22204 (P3_R1161_U56, P3_U3437);
  not ginst22205 (P3_R1161_U57, P3_U3072);
  not ginst22206 (P3_R1161_U58, P3_U3068);
  nand ginst22207 (P3_R1161_U59, P3_U3072, P3_U3437);
  and ginst22208 (P3_R1161_U6, P3_R1161_U236, P3_R1161_U237);
  not ginst22209 (P3_R1161_U60, P3_U3440);
  not ginst22210 (P3_R1161_U61, P3_U3419);
  not ginst22211 (P3_R1161_U62, P3_U3061);
  nand ginst22212 (P3_R1161_U63, P3_U3083, P3_U3413);
  not ginst22213 (P3_R1161_U64, P3_U3425);
  not ginst22214 (P3_R1161_U65, P3_U3071);
  not ginst22215 (P3_R1161_U66, P3_U3422);
  not ginst22216 (P3_R1161_U67, P3_U3062);
  nand ginst22217 (P3_R1161_U68, P3_U3062, P3_U3422);
  not ginst22218 (P3_R1161_U69, P3_U3428);
  and ginst22219 (P3_R1161_U7, P3_R1161_U245, P3_R1161_U246);
  not ginst22220 (P3_R1161_U70, P3_U3079);
  not ginst22221 (P3_R1161_U71, P3_U3431);
  not ginst22222 (P3_R1161_U72, P3_U3078);
  not ginst22223 (P3_R1161_U73, P3_U3434);
  not ginst22224 (P3_R1161_U74, P3_U3073);
  not ginst22225 (P3_R1161_U75, P3_U3443);
  not ginst22226 (P3_R1161_U76, P3_U3081);
  nand ginst22227 (P3_R1161_U77, P3_U3081, P3_U3443);
  not ginst22228 (P3_R1161_U78, P3_U3445);
  not ginst22229 (P3_R1161_U79, P3_U3080);
  and ginst22230 (P3_R1161_U8, P3_R1161_U263, P3_R1161_U264);
  nand ginst22231 (P3_R1161_U80, P3_U3080, P3_U3445);
  not ginst22232 (P3_R1161_U81, P3_U3907);
  not ginst22233 (P3_R1161_U82, P3_U3905);
  not ginst22234 (P3_R1161_U83, P3_U3060);
  not ginst22235 (P3_R1161_U84, P3_U3904);
  not ginst22236 (P3_R1161_U85, P3_U3065);
  nand ginst22237 (P3_R1161_U86, P3_U3056, P3_U3901);
  not ginst22238 (P3_R1161_U87, P3_U3053);
  not ginst22239 (P3_R1161_U88, P3_U3899);
  nand ginst22240 (P3_R1161_U89, P3_R1161_U176, P3_R1161_U306);
  and ginst22241 (P3_R1161_U9, P3_R1161_U271, P3_R1161_U272);
  not ginst22242 (P3_R1161_U90, P3_U3075);
  nand ginst22243 (P3_R1161_U91, P3_R1161_U315, P3_R1161_U77);
  nand ginst22244 (P3_R1161_U92, P3_R1161_U260, P3_R1161_U261);
  nand ginst22245 (P3_R1161_U93, P3_R1161_U337, P3_R1161_U68);
  nand ginst22246 (P3_R1161_U94, P3_R1161_U456, P3_R1161_U457);
  nand ginst22247 (P3_R1161_U95, P3_R1161_U503, P3_R1161_U504);
  nand ginst22248 (P3_R1161_U96, P3_R1161_U374, P3_R1161_U375);
  nand ginst22249 (P3_R1161_U97, P3_R1161_U379, P3_R1161_U380);
  nand ginst22250 (P3_R1161_U98, P3_R1161_U386, P3_R1161_U387);
  nand ginst22251 (P3_R1161_U99, P3_R1161_U393, P3_R1161_U394);
  and ginst22252 (P3_R1179_U10, P3_R1179_U263, P3_R1179_U264);
  nand ginst22253 (P3_R1179_U100, P3_R1179_U441, P3_R1179_U442);
  nand ginst22254 (P3_R1179_U101, P3_R1179_U446, P3_R1179_U447);
  nand ginst22255 (P3_R1179_U102, P3_R1179_U451, P3_R1179_U452);
  nand ginst22256 (P3_R1179_U103, P3_R1179_U456, P3_R1179_U457);
  nand ginst22257 (P3_R1179_U104, P3_R1179_U472, P3_R1179_U473);
  nand ginst22258 (P3_R1179_U105, P3_R1179_U477, P3_R1179_U478);
  nand ginst22259 (P3_R1179_U106, P3_R1179_U360, P3_R1179_U361);
  nand ginst22260 (P3_R1179_U107, P3_R1179_U369, P3_R1179_U370);
  nand ginst22261 (P3_R1179_U108, P3_R1179_U376, P3_R1179_U377);
  nand ginst22262 (P3_R1179_U109, P3_R1179_U380, P3_R1179_U381);
  and ginst22263 (P3_R1179_U11, P3_R1179_U191, P3_R1179_U286);
  nand ginst22264 (P3_R1179_U110, P3_R1179_U389, P3_R1179_U390);
  nand ginst22265 (P3_R1179_U111, P3_R1179_U410, P3_R1179_U411);
  nand ginst22266 (P3_R1179_U112, P3_R1179_U427, P3_R1179_U428);
  nand ginst22267 (P3_R1179_U113, P3_R1179_U431, P3_R1179_U432);
  nand ginst22268 (P3_R1179_U114, P3_R1179_U463, P3_R1179_U464);
  nand ginst22269 (P3_R1179_U115, P3_R1179_U467, P3_R1179_U468);
  nand ginst22270 (P3_R1179_U116, P3_R1179_U484, P3_R1179_U485);
  and ginst22271 (P3_R1179_U117, P3_R1179_U193, P3_R1179_U352);
  and ginst22272 (P3_R1179_U118, P3_R1179_U205, P3_R1179_U206);
  and ginst22273 (P3_R1179_U119, P3_R1179_U13, P3_R1179_U14);
  and ginst22274 (P3_R1179_U12, P3_R1179_U287, P3_R1179_U288);
  and ginst22275 (P3_R1179_U120, P3_R1179_U354, P3_R1179_U357);
  and ginst22276 (P3_R1179_U121, P3_R1179_U26, P3_R1179_U362, P3_R1179_U363);
  and ginst22277 (P3_R1179_U122, P3_R1179_U195, P3_R1179_U366);
  and ginst22278 (P3_R1179_U123, P3_R1179_U235, P3_R1179_U6);
  and ginst22279 (P3_R1179_U124, P3_R1179_U194, P3_R1179_U373);
  and ginst22280 (P3_R1179_U125, P3_R1179_U34, P3_R1179_U382, P3_R1179_U383);
  and ginst22281 (P3_R1179_U126, P3_R1179_U193, P3_R1179_U386);
  and ginst22282 (P3_R1179_U127, P3_R1179_U222, P3_R1179_U7);
  and ginst22283 (P3_R1179_U128, P3_R1179_U267, P3_R1179_U9);
  and ginst22284 (P3_R1179_U129, P3_R1179_U11, P3_R1179_U291);
  and ginst22285 (P3_R1179_U13, P3_R1179_U194, P3_R1179_U208, P3_R1179_U213);
  and ginst22286 (P3_R1179_U130, P3_R1179_U192, P3_R1179_U355);
  and ginst22287 (P3_R1179_U131, P3_R1179_U306, P3_R1179_U307);
  and ginst22288 (P3_R1179_U132, P3_R1179_U309, P3_R1179_U395);
  and ginst22289 (P3_R1179_U133, P3_R1179_U306, P3_R1179_U307);
  and ginst22290 (P3_R1179_U134, P3_R1179_U15, P3_R1179_U310);
  nand ginst22291 (P3_R1179_U135, P3_R1179_U398, P3_R1179_U399);
  and ginst22292 (P3_R1179_U136, P3_R1179_U403, P3_R1179_U404, P3_R1179_U87);
  and ginst22293 (P3_R1179_U137, P3_R1179_U192, P3_R1179_U407);
  nand ginst22294 (P3_R1179_U138, P3_R1179_U412, P3_R1179_U413);
  nand ginst22295 (P3_R1179_U139, P3_R1179_U417, P3_R1179_U418);
  and ginst22296 (P3_R1179_U14, P3_R1179_U195, P3_R1179_U218);
  and ginst22297 (P3_R1179_U140, P3_R1179_U12, P3_R1179_U322);
  and ginst22298 (P3_R1179_U141, P3_R1179_U191, P3_R1179_U424);
  nand ginst22299 (P3_R1179_U142, P3_R1179_U433, P3_R1179_U434);
  nand ginst22300 (P3_R1179_U143, P3_R1179_U438, P3_R1179_U439);
  nand ginst22301 (P3_R1179_U144, P3_R1179_U443, P3_R1179_U444);
  nand ginst22302 (P3_R1179_U145, P3_R1179_U448, P3_R1179_U449);
  nand ginst22303 (P3_R1179_U146, P3_R1179_U453, P3_R1179_U454);
  and ginst22304 (P3_R1179_U147, P3_R1179_U10, P3_R1179_U333);
  and ginst22305 (P3_R1179_U148, P3_R1179_U190, P3_R1179_U460);
  nand ginst22306 (P3_R1179_U149, P3_R1179_U469, P3_R1179_U470);
  and ginst22307 (P3_R1179_U15, P3_R1179_U391, P3_R1179_U392);
  nand ginst22308 (P3_R1179_U150, P3_R1179_U474, P3_R1179_U475);
  and ginst22309 (P3_R1179_U151, P3_R1179_U344, P3_R1179_U8);
  and ginst22310 (P3_R1179_U152, P3_R1179_U189, P3_R1179_U481);
  and ginst22311 (P3_R1179_U153, P3_R1179_U358, P3_R1179_U359);
  nand ginst22312 (P3_R1179_U154, P3_R1179_U120, P3_R1179_U356);
  and ginst22313 (P3_R1179_U155, P3_R1179_U367, P3_R1179_U368);
  and ginst22314 (P3_R1179_U156, P3_R1179_U374, P3_R1179_U375);
  and ginst22315 (P3_R1179_U157, P3_R1179_U378, P3_R1179_U379);
  nand ginst22316 (P3_R1179_U158, P3_R1179_U118, P3_R1179_U203);
  and ginst22317 (P3_R1179_U159, P3_R1179_U387, P3_R1179_U388);
  nand ginst22318 (P3_R1179_U16, P3_R1179_U342, P3_R1179_U345);
  not ginst22319 (P3_R1179_U160, P3_U3908);
  not ginst22320 (P3_R1179_U161, P3_U3054);
  and ginst22321 (P3_R1179_U162, P3_R1179_U396, P3_R1179_U397);
  nand ginst22322 (P3_R1179_U163, P3_R1179_U131, P3_R1179_U304);
  and ginst22323 (P3_R1179_U164, P3_R1179_U408, P3_R1179_U409);
  nand ginst22324 (P3_R1179_U165, P3_R1179_U297, P3_R1179_U298);
  nand ginst22325 (P3_R1179_U166, P3_R1179_U293, P3_R1179_U294);
  and ginst22326 (P3_R1179_U167, P3_R1179_U425, P3_R1179_U426);
  and ginst22327 (P3_R1179_U168, P3_R1179_U429, P3_R1179_U430);
  nand ginst22328 (P3_R1179_U169, P3_R1179_U283, P3_R1179_U284);
  nand ginst22329 (P3_R1179_U17, P3_R1179_U331, P3_R1179_U334);
  nand ginst22330 (P3_R1179_U170, P3_R1179_U279, P3_R1179_U280);
  not ginst22331 (P3_R1179_U171, P3_U3392);
  nand ginst22332 (P3_R1179_U172, P3_R1179_U95, P3_U3387);
  nand ginst22333 (P3_R1179_U173, P3_R1179_U184, P3_R1179_U276, P3_R1179_U350);
  not ginst22334 (P3_R1179_U174, P3_U3443);
  nand ginst22335 (P3_R1179_U175, P3_R1179_U273, P3_R1179_U274);
  nand ginst22336 (P3_R1179_U176, P3_R1179_U269, P3_R1179_U270);
  and ginst22337 (P3_R1179_U177, P3_R1179_U461, P3_R1179_U462);
  and ginst22338 (P3_R1179_U178, P3_R1179_U465, P3_R1179_U466);
  nand ginst22339 (P3_R1179_U179, P3_R1179_U259, P3_R1179_U260);
  nand ginst22340 (P3_R1179_U18, P3_R1179_U320, P3_R1179_U323);
  nand ginst22341 (P3_R1179_U180, P3_R1179_U255, P3_R1179_U256);
  nand ginst22342 (P3_R1179_U181, P3_R1179_U251, P3_R1179_U252);
  and ginst22343 (P3_R1179_U182, P3_R1179_U482, P3_R1179_U483);
  nand ginst22344 (P3_R1179_U183, P3_R1179_U132, P3_R1179_U163);
  nand ginst22345 (P3_R1179_U184, P3_R1179_U174, P3_R1179_U175);
  nand ginst22346 (P3_R1179_U185, P3_R1179_U171, P3_R1179_U172);
  not ginst22347 (P3_R1179_U186, P3_R1179_U87);
  not ginst22348 (P3_R1179_U187, P3_R1179_U34);
  not ginst22349 (P3_R1179_U188, P3_R1179_U26);
  nand ginst22350 (P3_R1179_U189, P3_R1179_U54, P3_U3419);
  nand ginst22351 (P3_R1179_U19, P3_R1179_U312, P3_R1179_U314);
  nand ginst22352 (P3_R1179_U190, P3_R1179_U64, P3_U3434);
  nand ginst22353 (P3_R1179_U191, P3_R1179_U78, P3_U3905);
  nand ginst22354 (P3_R1179_U192, P3_R1179_U86, P3_U3901);
  nand ginst22355 (P3_R1179_U193, P3_R1179_U33, P3_U3395);
  nand ginst22356 (P3_R1179_U194, P3_R1179_U41, P3_U3404);
  nand ginst22357 (P3_R1179_U195, P3_R1179_U25, P3_U3410);
  not ginst22358 (P3_R1179_U196, P3_R1179_U66);
  not ginst22359 (P3_R1179_U197, P3_R1179_U80);
  not ginst22360 (P3_R1179_U198, P3_R1179_U43);
  not ginst22361 (P3_R1179_U199, P3_R1179_U55);
  nand ginst22362 (P3_R1179_U20, P3_R1179_U162, P3_R1179_U183, P3_R1179_U351);
  not ginst22363 (P3_R1179_U200, P3_R1179_U172);
  nand ginst22364 (P3_R1179_U201, P3_R1179_U172, P3_U3077);
  not ginst22365 (P3_R1179_U202, P3_R1179_U49);
  nand ginst22366 (P3_R1179_U203, P3_R1179_U117, P3_R1179_U49);
  nand ginst22367 (P3_R1179_U204, P3_R1179_U34, P3_R1179_U35);
  nand ginst22368 (P3_R1179_U205, P3_R1179_U204, P3_R1179_U32);
  nand ginst22369 (P3_R1179_U206, P3_R1179_U187, P3_U3063);
  not ginst22370 (P3_R1179_U207, P3_R1179_U158);
  nand ginst22371 (P3_R1179_U208, P3_R1179_U40, P3_U3407);
  nand ginst22372 (P3_R1179_U209, P3_R1179_U37, P3_U3070);
  nand ginst22373 (P3_R1179_U21, P3_R1179_U241, P3_R1179_U243);
  nand ginst22374 (P3_R1179_U210, P3_R1179_U36, P3_U3066);
  nand ginst22375 (P3_R1179_U211, P3_R1179_U194, P3_R1179_U198);
  nand ginst22376 (P3_R1179_U212, P3_R1179_U211, P3_R1179_U6);
  nand ginst22377 (P3_R1179_U213, P3_R1179_U42, P3_U3401);
  nand ginst22378 (P3_R1179_U214, P3_R1179_U40, P3_U3407);
  nand ginst22379 (P3_R1179_U215, P3_R1179_U13, P3_R1179_U158);
  not ginst22380 (P3_R1179_U216, P3_R1179_U44);
  not ginst22381 (P3_R1179_U217, P3_R1179_U47);
  nand ginst22382 (P3_R1179_U218, P3_R1179_U27, P3_U3413);
  nand ginst22383 (P3_R1179_U219, P3_R1179_U26, P3_R1179_U27);
  nand ginst22384 (P3_R1179_U22, P3_R1179_U233, P3_R1179_U236);
  nand ginst22385 (P3_R1179_U220, P3_R1179_U188, P3_U3083);
  not ginst22386 (P3_R1179_U221, P3_R1179_U154);
  nand ginst22387 (P3_R1179_U222, P3_R1179_U46, P3_U3416);
  nand ginst22388 (P3_R1179_U223, P3_R1179_U222, P3_R1179_U55);
  nand ginst22389 (P3_R1179_U224, P3_R1179_U217, P3_R1179_U26);
  nand ginst22390 (P3_R1179_U225, P3_R1179_U122, P3_R1179_U224);
  nand ginst22391 (P3_R1179_U226, P3_R1179_U195, P3_R1179_U47);
  nand ginst22392 (P3_R1179_U227, P3_R1179_U121, P3_R1179_U226);
  nand ginst22393 (P3_R1179_U228, P3_R1179_U195, P3_R1179_U26);
  nand ginst22394 (P3_R1179_U229, P3_R1179_U158, P3_R1179_U213);
  nand ginst22395 (P3_R1179_U23, P3_R1179_U225, P3_R1179_U227);
  not ginst22396 (P3_R1179_U230, P3_R1179_U48);
  nand ginst22397 (P3_R1179_U231, P3_R1179_U36, P3_U3066);
  nand ginst22398 (P3_R1179_U232, P3_R1179_U230, P3_R1179_U231);
  nand ginst22399 (P3_R1179_U233, P3_R1179_U124, P3_R1179_U232);
  nand ginst22400 (P3_R1179_U234, P3_R1179_U194, P3_R1179_U48);
  nand ginst22401 (P3_R1179_U235, P3_R1179_U40, P3_U3407);
  nand ginst22402 (P3_R1179_U236, P3_R1179_U123, P3_R1179_U234);
  nand ginst22403 (P3_R1179_U237, P3_R1179_U36, P3_U3066);
  nand ginst22404 (P3_R1179_U238, P3_R1179_U194, P3_R1179_U237);
  nand ginst22405 (P3_R1179_U239, P3_R1179_U213, P3_R1179_U43);
  nand ginst22406 (P3_R1179_U24, P3_R1179_U172, P3_R1179_U348);
  nand ginst22407 (P3_R1179_U240, P3_R1179_U202, P3_R1179_U34);
  nand ginst22408 (P3_R1179_U241, P3_R1179_U126, P3_R1179_U240);
  nand ginst22409 (P3_R1179_U242, P3_R1179_U193, P3_R1179_U49);
  nand ginst22410 (P3_R1179_U243, P3_R1179_U125, P3_R1179_U242);
  nand ginst22411 (P3_R1179_U244, P3_R1179_U193, P3_R1179_U34);
  nand ginst22412 (P3_R1179_U245, P3_R1179_U53, P3_U3422);
  nand ginst22413 (P3_R1179_U246, P3_R1179_U51, P3_U3062);
  nand ginst22414 (P3_R1179_U247, P3_R1179_U52, P3_U3061);
  nand ginst22415 (P3_R1179_U248, P3_R1179_U199, P3_R1179_U7);
  nand ginst22416 (P3_R1179_U249, P3_R1179_U248, P3_R1179_U8);
  not ginst22417 (P3_R1179_U25, P3_U3069);
  nand ginst22418 (P3_R1179_U250, P3_R1179_U53, P3_U3422);
  nand ginst22419 (P3_R1179_U251, P3_R1179_U127, P3_R1179_U154);
  nand ginst22420 (P3_R1179_U252, P3_R1179_U249, P3_R1179_U250);
  not ginst22421 (P3_R1179_U253, P3_R1179_U181);
  nand ginst22422 (P3_R1179_U254, P3_R1179_U57, P3_U3425);
  nand ginst22423 (P3_R1179_U255, P3_R1179_U181, P3_R1179_U254);
  nand ginst22424 (P3_R1179_U256, P3_R1179_U56, P3_U3071);
  not ginst22425 (P3_R1179_U257, P3_R1179_U180);
  nand ginst22426 (P3_R1179_U258, P3_R1179_U59, P3_U3428);
  nand ginst22427 (P3_R1179_U259, P3_R1179_U180, P3_R1179_U258);
  nand ginst22428 (P3_R1179_U26, P3_R1179_U39, P3_U3069);
  nand ginst22429 (P3_R1179_U260, P3_R1179_U58, P3_U3079);
  not ginst22430 (P3_R1179_U261, P3_R1179_U179);
  nand ginst22431 (P3_R1179_U262, P3_R1179_U63, P3_U3437);
  nand ginst22432 (P3_R1179_U263, P3_R1179_U60, P3_U3072);
  nand ginst22433 (P3_R1179_U264, P3_R1179_U61, P3_U3073);
  nand ginst22434 (P3_R1179_U265, P3_R1179_U196, P3_R1179_U9);
  nand ginst22435 (P3_R1179_U266, P3_R1179_U10, P3_R1179_U265);
  nand ginst22436 (P3_R1179_U267, P3_R1179_U65, P3_U3431);
  nand ginst22437 (P3_R1179_U268, P3_R1179_U63, P3_U3437);
  nand ginst22438 (P3_R1179_U269, P3_R1179_U128, P3_R1179_U179);
  not ginst22439 (P3_R1179_U27, P3_U3083);
  nand ginst22440 (P3_R1179_U270, P3_R1179_U266, P3_R1179_U268);
  not ginst22441 (P3_R1179_U271, P3_R1179_U176);
  nand ginst22442 (P3_R1179_U272, P3_R1179_U68, P3_U3440);
  nand ginst22443 (P3_R1179_U273, P3_R1179_U176, P3_R1179_U272);
  nand ginst22444 (P3_R1179_U274, P3_R1179_U67, P3_U3068);
  not ginst22445 (P3_R1179_U275, P3_R1179_U175);
  nand ginst22446 (P3_R1179_U276, P3_R1179_U175, P3_U3081);
  not ginst22447 (P3_R1179_U277, P3_R1179_U173);
  nand ginst22448 (P3_R1179_U278, P3_R1179_U71, P3_U3445);
  nand ginst22449 (P3_R1179_U279, P3_R1179_U173, P3_R1179_U278);
  not ginst22450 (P3_R1179_U28, P3_U3413);
  nand ginst22451 (P3_R1179_U280, P3_R1179_U70, P3_U3080);
  not ginst22452 (P3_R1179_U281, P3_R1179_U170);
  nand ginst22453 (P3_R1179_U282, P3_R1179_U73, P3_U3907);
  nand ginst22454 (P3_R1179_U283, P3_R1179_U170, P3_R1179_U282);
  nand ginst22455 (P3_R1179_U284, P3_R1179_U72, P3_U3075);
  not ginst22456 (P3_R1179_U285, P3_R1179_U169);
  nand ginst22457 (P3_R1179_U286, P3_R1179_U77, P3_U3904);
  nand ginst22458 (P3_R1179_U287, P3_R1179_U74, P3_U3065);
  nand ginst22459 (P3_R1179_U288, P3_R1179_U75, P3_U3060);
  nand ginst22460 (P3_R1179_U289, P3_R1179_U11, P3_R1179_U197);
  not ginst22461 (P3_R1179_U29, P3_U3395);
  nand ginst22462 (P3_R1179_U290, P3_R1179_U12, P3_R1179_U289);
  nand ginst22463 (P3_R1179_U291, P3_R1179_U79, P3_U3906);
  nand ginst22464 (P3_R1179_U292, P3_R1179_U77, P3_U3904);
  nand ginst22465 (P3_R1179_U293, P3_R1179_U129, P3_R1179_U169);
  nand ginst22466 (P3_R1179_U294, P3_R1179_U290, P3_R1179_U292);
  not ginst22467 (P3_R1179_U295, P3_R1179_U166);
  nand ginst22468 (P3_R1179_U296, P3_R1179_U82, P3_U3903);
  nand ginst22469 (P3_R1179_U297, P3_R1179_U166, P3_R1179_U296);
  nand ginst22470 (P3_R1179_U298, P3_R1179_U81, P3_U3064);
  not ginst22471 (P3_R1179_U299, P3_R1179_U165);
  not ginst22472 (P3_R1179_U30, P3_U3387);
  nand ginst22473 (P3_R1179_U300, P3_R1179_U84, P3_U3902);
  nand ginst22474 (P3_R1179_U301, P3_R1179_U165, P3_R1179_U300);
  nand ginst22475 (P3_R1179_U302, P3_R1179_U83, P3_U3057);
  not ginst22476 (P3_R1179_U303, P3_R1179_U91);
  nand ginst22477 (P3_R1179_U304, P3_R1179_U130, P3_R1179_U91);
  nand ginst22478 (P3_R1179_U305, P3_R1179_U87, P3_R1179_U88);
  nand ginst22479 (P3_R1179_U306, P3_R1179_U305, P3_R1179_U85);
  nand ginst22480 (P3_R1179_U307, P3_R1179_U186, P3_U3052);
  not ginst22481 (P3_R1179_U308, P3_R1179_U163);
  nand ginst22482 (P3_R1179_U309, P3_R1179_U90, P3_U3899);
  not ginst22483 (P3_R1179_U31, P3_U3077);
  nand ginst22484 (P3_R1179_U310, P3_R1179_U89, P3_U3053);
  nand ginst22485 (P3_R1179_U311, P3_R1179_U303, P3_R1179_U87);
  nand ginst22486 (P3_R1179_U312, P3_R1179_U137, P3_R1179_U311);
  nand ginst22487 (P3_R1179_U313, P3_R1179_U192, P3_R1179_U91);
  nand ginst22488 (P3_R1179_U314, P3_R1179_U136, P3_R1179_U313);
  nand ginst22489 (P3_R1179_U315, P3_R1179_U192, P3_R1179_U87);
  nand ginst22490 (P3_R1179_U316, P3_R1179_U169, P3_R1179_U291);
  not ginst22491 (P3_R1179_U317, P3_R1179_U92);
  nand ginst22492 (P3_R1179_U318, P3_R1179_U75, P3_U3060);
  nand ginst22493 (P3_R1179_U319, P3_R1179_U317, P3_R1179_U318);
  not ginst22494 (P3_R1179_U32, P3_U3398);
  nand ginst22495 (P3_R1179_U320, P3_R1179_U141, P3_R1179_U319);
  nand ginst22496 (P3_R1179_U321, P3_R1179_U191, P3_R1179_U92);
  nand ginst22497 (P3_R1179_U322, P3_R1179_U77, P3_U3904);
  nand ginst22498 (P3_R1179_U323, P3_R1179_U140, P3_R1179_U321);
  nand ginst22499 (P3_R1179_U324, P3_R1179_U75, P3_U3060);
  nand ginst22500 (P3_R1179_U325, P3_R1179_U191, P3_R1179_U324);
  nand ginst22501 (P3_R1179_U326, P3_R1179_U291, P3_R1179_U80);
  nand ginst22502 (P3_R1179_U327, P3_R1179_U179, P3_R1179_U267);
  not ginst22503 (P3_R1179_U328, P3_R1179_U93);
  nand ginst22504 (P3_R1179_U329, P3_R1179_U61, P3_U3073);
  not ginst22505 (P3_R1179_U33, P3_U3067);
  nand ginst22506 (P3_R1179_U330, P3_R1179_U328, P3_R1179_U329);
  nand ginst22507 (P3_R1179_U331, P3_R1179_U148, P3_R1179_U330);
  nand ginst22508 (P3_R1179_U332, P3_R1179_U190, P3_R1179_U93);
  nand ginst22509 (P3_R1179_U333, P3_R1179_U63, P3_U3437);
  nand ginst22510 (P3_R1179_U334, P3_R1179_U147, P3_R1179_U332);
  nand ginst22511 (P3_R1179_U335, P3_R1179_U61, P3_U3073);
  nand ginst22512 (P3_R1179_U336, P3_R1179_U190, P3_R1179_U335);
  nand ginst22513 (P3_R1179_U337, P3_R1179_U267, P3_R1179_U66);
  nand ginst22514 (P3_R1179_U338, P3_R1179_U154, P3_R1179_U222);
  not ginst22515 (P3_R1179_U339, P3_R1179_U94);
  nand ginst22516 (P3_R1179_U34, P3_R1179_U29, P3_U3067);
  nand ginst22517 (P3_R1179_U340, P3_R1179_U52, P3_U3061);
  nand ginst22518 (P3_R1179_U341, P3_R1179_U339, P3_R1179_U340);
  nand ginst22519 (P3_R1179_U342, P3_R1179_U152, P3_R1179_U341);
  nand ginst22520 (P3_R1179_U343, P3_R1179_U189, P3_R1179_U94);
  nand ginst22521 (P3_R1179_U344, P3_R1179_U53, P3_U3422);
  nand ginst22522 (P3_R1179_U345, P3_R1179_U151, P3_R1179_U343);
  nand ginst22523 (P3_R1179_U346, P3_R1179_U52, P3_U3061);
  nand ginst22524 (P3_R1179_U347, P3_R1179_U189, P3_R1179_U346);
  nand ginst22525 (P3_R1179_U348, P3_R1179_U30, P3_U3076);
  nand ginst22526 (P3_R1179_U349, P3_R1179_U171, P3_U3077);
  not ginst22527 (P3_R1179_U35, P3_U3063);
  nand ginst22528 (P3_R1179_U350, P3_R1179_U174, P3_U3081);
  nand ginst22529 (P3_R1179_U351, P3_R1179_U133, P3_R1179_U134, P3_R1179_U304);
  nand ginst22530 (P3_R1179_U352, P3_R1179_U35, P3_U3398);
  nand ginst22531 (P3_R1179_U353, P3_R1179_U220, P3_U3413);
  nand ginst22532 (P3_R1179_U354, P3_R1179_U219, P3_R1179_U353);
  nand ginst22533 (P3_R1179_U355, P3_R1179_U88, P3_U3900);
  nand ginst22534 (P3_R1179_U356, P3_R1179_U119, P3_R1179_U158);
  nand ginst22535 (P3_R1179_U357, P3_R1179_U14, P3_R1179_U216);
  nand ginst22536 (P3_R1179_U358, P3_R1179_U46, P3_U3416);
  nand ginst22537 (P3_R1179_U359, P3_R1179_U45, P3_U3082);
  not ginst22538 (P3_R1179_U36, P3_U3404);
  nand ginst22539 (P3_R1179_U360, P3_R1179_U154, P3_R1179_U223);
  nand ginst22540 (P3_R1179_U361, P3_R1179_U153, P3_R1179_U221);
  nand ginst22541 (P3_R1179_U362, P3_R1179_U27, P3_U3413);
  nand ginst22542 (P3_R1179_U363, P3_R1179_U28, P3_U3083);
  nand ginst22543 (P3_R1179_U364, P3_R1179_U27, P3_U3413);
  nand ginst22544 (P3_R1179_U365, P3_R1179_U28, P3_U3083);
  nand ginst22545 (P3_R1179_U366, P3_R1179_U364, P3_R1179_U365);
  nand ginst22546 (P3_R1179_U367, P3_R1179_U25, P3_U3410);
  nand ginst22547 (P3_R1179_U368, P3_R1179_U39, P3_U3069);
  nand ginst22548 (P3_R1179_U369, P3_R1179_U228, P3_R1179_U47);
  not ginst22549 (P3_R1179_U37, P3_U3407);
  nand ginst22550 (P3_R1179_U370, P3_R1179_U155, P3_R1179_U217);
  nand ginst22551 (P3_R1179_U371, P3_R1179_U40, P3_U3407);
  nand ginst22552 (P3_R1179_U372, P3_R1179_U37, P3_U3070);
  nand ginst22553 (P3_R1179_U373, P3_R1179_U371, P3_R1179_U372);
  nand ginst22554 (P3_R1179_U374, P3_R1179_U41, P3_U3404);
  nand ginst22555 (P3_R1179_U375, P3_R1179_U36, P3_U3066);
  nand ginst22556 (P3_R1179_U376, P3_R1179_U238, P3_R1179_U48);
  nand ginst22557 (P3_R1179_U377, P3_R1179_U156, P3_R1179_U230);
  nand ginst22558 (P3_R1179_U378, P3_R1179_U42, P3_U3401);
  nand ginst22559 (P3_R1179_U379, P3_R1179_U38, P3_U3059);
  not ginst22560 (P3_R1179_U38, P3_U3401);
  nand ginst22561 (P3_R1179_U380, P3_R1179_U158, P3_R1179_U239);
  nand ginst22562 (P3_R1179_U381, P3_R1179_U157, P3_R1179_U207);
  nand ginst22563 (P3_R1179_U382, P3_R1179_U35, P3_U3398);
  nand ginst22564 (P3_R1179_U383, P3_R1179_U32, P3_U3063);
  nand ginst22565 (P3_R1179_U384, P3_R1179_U35, P3_U3398);
  nand ginst22566 (P3_R1179_U385, P3_R1179_U32, P3_U3063);
  nand ginst22567 (P3_R1179_U386, P3_R1179_U384, P3_R1179_U385);
  nand ginst22568 (P3_R1179_U387, P3_R1179_U33, P3_U3395);
  nand ginst22569 (P3_R1179_U388, P3_R1179_U29, P3_U3067);
  nand ginst22570 (P3_R1179_U389, P3_R1179_U244, P3_R1179_U49);
  not ginst22571 (P3_R1179_U39, P3_U3410);
  nand ginst22572 (P3_R1179_U390, P3_R1179_U159, P3_R1179_U202);
  nand ginst22573 (P3_R1179_U391, P3_R1179_U161, P3_U3908);
  nand ginst22574 (P3_R1179_U392, P3_R1179_U160, P3_U3054);
  nand ginst22575 (P3_R1179_U393, P3_R1179_U161, P3_U3908);
  nand ginst22576 (P3_R1179_U394, P3_R1179_U160, P3_U3054);
  nand ginst22577 (P3_R1179_U395, P3_R1179_U393, P3_R1179_U394);
  nand ginst22578 (P3_R1179_U396, P3_R1179_U395, P3_R1179_U89, P3_U3053);
  nand ginst22579 (P3_R1179_U397, P3_R1179_U15, P3_R1179_U90, P3_U3899);
  nand ginst22580 (P3_R1179_U398, P3_R1179_U90, P3_U3899);
  nand ginst22581 (P3_R1179_U399, P3_R1179_U89, P3_U3053);
  not ginst22582 (P3_R1179_U40, P3_U3070);
  not ginst22583 (P3_R1179_U400, P3_R1179_U135);
  nand ginst22584 (P3_R1179_U401, P3_R1179_U308, P3_R1179_U400);
  nand ginst22585 (P3_R1179_U402, P3_R1179_U135, P3_R1179_U163);
  nand ginst22586 (P3_R1179_U403, P3_R1179_U88, P3_U3900);
  nand ginst22587 (P3_R1179_U404, P3_R1179_U85, P3_U3052);
  nand ginst22588 (P3_R1179_U405, P3_R1179_U88, P3_U3900);
  nand ginst22589 (P3_R1179_U406, P3_R1179_U85, P3_U3052);
  nand ginst22590 (P3_R1179_U407, P3_R1179_U405, P3_R1179_U406);
  nand ginst22591 (P3_R1179_U408, P3_R1179_U86, P3_U3901);
  nand ginst22592 (P3_R1179_U409, P3_R1179_U50, P3_U3056);
  not ginst22593 (P3_R1179_U41, P3_U3066);
  nand ginst22594 (P3_R1179_U410, P3_R1179_U315, P3_R1179_U91);
  nand ginst22595 (P3_R1179_U411, P3_R1179_U164, P3_R1179_U303);
  nand ginst22596 (P3_R1179_U412, P3_R1179_U84, P3_U3902);
  nand ginst22597 (P3_R1179_U413, P3_R1179_U83, P3_U3057);
  not ginst22598 (P3_R1179_U414, P3_R1179_U138);
  nand ginst22599 (P3_R1179_U415, P3_R1179_U299, P3_R1179_U414);
  nand ginst22600 (P3_R1179_U416, P3_R1179_U138, P3_R1179_U165);
  nand ginst22601 (P3_R1179_U417, P3_R1179_U82, P3_U3903);
  nand ginst22602 (P3_R1179_U418, P3_R1179_U81, P3_U3064);
  not ginst22603 (P3_R1179_U419, P3_R1179_U139);
  not ginst22604 (P3_R1179_U42, P3_U3059);
  nand ginst22605 (P3_R1179_U420, P3_R1179_U295, P3_R1179_U419);
  nand ginst22606 (P3_R1179_U421, P3_R1179_U139, P3_R1179_U166);
  nand ginst22607 (P3_R1179_U422, P3_R1179_U77, P3_U3904);
  nand ginst22608 (P3_R1179_U423, P3_R1179_U74, P3_U3065);
  nand ginst22609 (P3_R1179_U424, P3_R1179_U422, P3_R1179_U423);
  nand ginst22610 (P3_R1179_U425, P3_R1179_U78, P3_U3905);
  nand ginst22611 (P3_R1179_U426, P3_R1179_U75, P3_U3060);
  nand ginst22612 (P3_R1179_U427, P3_R1179_U325, P3_R1179_U92);
  nand ginst22613 (P3_R1179_U428, P3_R1179_U167, P3_R1179_U317);
  nand ginst22614 (P3_R1179_U429, P3_R1179_U79, P3_U3906);
  nand ginst22615 (P3_R1179_U43, P3_R1179_U38, P3_U3059);
  nand ginst22616 (P3_R1179_U430, P3_R1179_U76, P3_U3074);
  nand ginst22617 (P3_R1179_U431, P3_R1179_U169, P3_R1179_U326);
  nand ginst22618 (P3_R1179_U432, P3_R1179_U168, P3_R1179_U285);
  nand ginst22619 (P3_R1179_U433, P3_R1179_U73, P3_U3907);
  nand ginst22620 (P3_R1179_U434, P3_R1179_U72, P3_U3075);
  not ginst22621 (P3_R1179_U435, P3_R1179_U142);
  nand ginst22622 (P3_R1179_U436, P3_R1179_U281, P3_R1179_U435);
  nand ginst22623 (P3_R1179_U437, P3_R1179_U142, P3_R1179_U170);
  nand ginst22624 (P3_R1179_U438, P3_R1179_U31, P3_U3392);
  nand ginst22625 (P3_R1179_U439, P3_R1179_U171, P3_U3077);
  nand ginst22626 (P3_R1179_U44, P3_R1179_U212, P3_R1179_U214);
  not ginst22627 (P3_R1179_U440, P3_R1179_U143);
  nand ginst22628 (P3_R1179_U441, P3_R1179_U200, P3_R1179_U440);
  nand ginst22629 (P3_R1179_U442, P3_R1179_U143, P3_R1179_U172);
  nand ginst22630 (P3_R1179_U443, P3_R1179_U71, P3_U3445);
  nand ginst22631 (P3_R1179_U444, P3_R1179_U70, P3_U3080);
  not ginst22632 (P3_R1179_U445, P3_R1179_U144);
  nand ginst22633 (P3_R1179_U446, P3_R1179_U277, P3_R1179_U445);
  nand ginst22634 (P3_R1179_U447, P3_R1179_U144, P3_R1179_U173);
  nand ginst22635 (P3_R1179_U448, P3_R1179_U69, P3_U3443);
  nand ginst22636 (P3_R1179_U449, P3_R1179_U174, P3_U3081);
  not ginst22637 (P3_R1179_U45, P3_U3416);
  not ginst22638 (P3_R1179_U450, P3_R1179_U145);
  nand ginst22639 (P3_R1179_U451, P3_R1179_U275, P3_R1179_U450);
  nand ginst22640 (P3_R1179_U452, P3_R1179_U145, P3_R1179_U175);
  nand ginst22641 (P3_R1179_U453, P3_R1179_U68, P3_U3440);
  nand ginst22642 (P3_R1179_U454, P3_R1179_U67, P3_U3068);
  not ginst22643 (P3_R1179_U455, P3_R1179_U146);
  nand ginst22644 (P3_R1179_U456, P3_R1179_U271, P3_R1179_U455);
  nand ginst22645 (P3_R1179_U457, P3_R1179_U146, P3_R1179_U176);
  nand ginst22646 (P3_R1179_U458, P3_R1179_U63, P3_U3437);
  nand ginst22647 (P3_R1179_U459, P3_R1179_U60, P3_U3072);
  not ginst22648 (P3_R1179_U46, P3_U3082);
  nand ginst22649 (P3_R1179_U460, P3_R1179_U458, P3_R1179_U459);
  nand ginst22650 (P3_R1179_U461, P3_R1179_U64, P3_U3434);
  nand ginst22651 (P3_R1179_U462, P3_R1179_U61, P3_U3073);
  nand ginst22652 (P3_R1179_U463, P3_R1179_U336, P3_R1179_U93);
  nand ginst22653 (P3_R1179_U464, P3_R1179_U177, P3_R1179_U328);
  nand ginst22654 (P3_R1179_U465, P3_R1179_U65, P3_U3431);
  nand ginst22655 (P3_R1179_U466, P3_R1179_U62, P3_U3078);
  nand ginst22656 (P3_R1179_U467, P3_R1179_U179, P3_R1179_U337);
  nand ginst22657 (P3_R1179_U468, P3_R1179_U178, P3_R1179_U261);
  nand ginst22658 (P3_R1179_U469, P3_R1179_U59, P3_U3428);
  nand ginst22659 (P3_R1179_U47, P3_R1179_U215, P3_R1179_U44);
  nand ginst22660 (P3_R1179_U470, P3_R1179_U58, P3_U3079);
  not ginst22661 (P3_R1179_U471, P3_R1179_U149);
  nand ginst22662 (P3_R1179_U472, P3_R1179_U257, P3_R1179_U471);
  nand ginst22663 (P3_R1179_U473, P3_R1179_U149, P3_R1179_U180);
  nand ginst22664 (P3_R1179_U474, P3_R1179_U57, P3_U3425);
  nand ginst22665 (P3_R1179_U475, P3_R1179_U56, P3_U3071);
  not ginst22666 (P3_R1179_U476, P3_R1179_U150);
  nand ginst22667 (P3_R1179_U477, P3_R1179_U253, P3_R1179_U476);
  nand ginst22668 (P3_R1179_U478, P3_R1179_U150, P3_R1179_U181);
  nand ginst22669 (P3_R1179_U479, P3_R1179_U53, P3_U3422);
  nand ginst22670 (P3_R1179_U48, P3_R1179_U229, P3_R1179_U43);
  nand ginst22671 (P3_R1179_U480, P3_R1179_U51, P3_U3062);
  nand ginst22672 (P3_R1179_U481, P3_R1179_U479, P3_R1179_U480);
  nand ginst22673 (P3_R1179_U482, P3_R1179_U54, P3_U3419);
  nand ginst22674 (P3_R1179_U483, P3_R1179_U52, P3_U3061);
  nand ginst22675 (P3_R1179_U484, P3_R1179_U347, P3_R1179_U94);
  nand ginst22676 (P3_R1179_U485, P3_R1179_U182, P3_R1179_U339);
  nand ginst22677 (P3_R1179_U49, P3_R1179_U185, P3_R1179_U201, P3_R1179_U349);
  not ginst22678 (P3_R1179_U50, P3_U3901);
  not ginst22679 (P3_R1179_U51, P3_U3422);
  not ginst22680 (P3_R1179_U52, P3_U3419);
  not ginst22681 (P3_R1179_U53, P3_U3062);
  not ginst22682 (P3_R1179_U54, P3_U3061);
  nand ginst22683 (P3_R1179_U55, P3_R1179_U45, P3_U3082);
  not ginst22684 (P3_R1179_U56, P3_U3425);
  not ginst22685 (P3_R1179_U57, P3_U3071);
  not ginst22686 (P3_R1179_U58, P3_U3428);
  not ginst22687 (P3_R1179_U59, P3_U3079);
  and ginst22688 (P3_R1179_U6, P3_R1179_U209, P3_R1179_U210);
  not ginst22689 (P3_R1179_U60, P3_U3437);
  not ginst22690 (P3_R1179_U61, P3_U3434);
  not ginst22691 (P3_R1179_U62, P3_U3431);
  not ginst22692 (P3_R1179_U63, P3_U3072);
  not ginst22693 (P3_R1179_U64, P3_U3073);
  not ginst22694 (P3_R1179_U65, P3_U3078);
  nand ginst22695 (P3_R1179_U66, P3_R1179_U62, P3_U3078);
  not ginst22696 (P3_R1179_U67, P3_U3440);
  not ginst22697 (P3_R1179_U68, P3_U3068);
  not ginst22698 (P3_R1179_U69, P3_U3081);
  and ginst22699 (P3_R1179_U7, P3_R1179_U189, P3_R1179_U245);
  not ginst22700 (P3_R1179_U70, P3_U3445);
  not ginst22701 (P3_R1179_U71, P3_U3080);
  not ginst22702 (P3_R1179_U72, P3_U3907);
  not ginst22703 (P3_R1179_U73, P3_U3075);
  not ginst22704 (P3_R1179_U74, P3_U3904);
  not ginst22705 (P3_R1179_U75, P3_U3905);
  not ginst22706 (P3_R1179_U76, P3_U3906);
  not ginst22707 (P3_R1179_U77, P3_U3065);
  not ginst22708 (P3_R1179_U78, P3_U3060);
  not ginst22709 (P3_R1179_U79, P3_U3074);
  and ginst22710 (P3_R1179_U8, P3_R1179_U246, P3_R1179_U247);
  nand ginst22711 (P3_R1179_U80, P3_R1179_U76, P3_U3074);
  not ginst22712 (P3_R1179_U81, P3_U3903);
  not ginst22713 (P3_R1179_U82, P3_U3064);
  not ginst22714 (P3_R1179_U83, P3_U3902);
  not ginst22715 (P3_R1179_U84, P3_U3057);
  not ginst22716 (P3_R1179_U85, P3_U3900);
  not ginst22717 (P3_R1179_U86, P3_U3056);
  nand ginst22718 (P3_R1179_U87, P3_R1179_U50, P3_U3056);
  not ginst22719 (P3_R1179_U88, P3_U3052);
  not ginst22720 (P3_R1179_U89, P3_U3899);
  and ginst22721 (P3_R1179_U9, P3_R1179_U190, P3_R1179_U262);
  not ginst22722 (P3_R1179_U90, P3_U3053);
  nand ginst22723 (P3_R1179_U91, P3_R1179_U301, P3_R1179_U302);
  nand ginst22724 (P3_R1179_U92, P3_R1179_U316, P3_R1179_U80);
  nand ginst22725 (P3_R1179_U93, P3_R1179_U327, P3_R1179_U66);
  nand ginst22726 (P3_R1179_U94, P3_R1179_U338, P3_R1179_U55);
  not ginst22727 (P3_R1179_U95, P3_U3076);
  nand ginst22728 (P3_R1179_U96, P3_R1179_U401, P3_R1179_U402);
  nand ginst22729 (P3_R1179_U97, P3_R1179_U415, P3_R1179_U416);
  nand ginst22730 (P3_R1179_U98, P3_R1179_U420, P3_R1179_U421);
  nand ginst22731 (P3_R1179_U99, P3_R1179_U436, P3_R1179_U437);
  and ginst22732 (P3_R1200_U10, P3_R1200_U263, P3_R1200_U264);
  nand ginst22733 (P3_R1200_U100, P3_R1200_U441, P3_R1200_U442);
  nand ginst22734 (P3_R1200_U101, P3_R1200_U446, P3_R1200_U447);
  nand ginst22735 (P3_R1200_U102, P3_R1200_U451, P3_R1200_U452);
  nand ginst22736 (P3_R1200_U103, P3_R1200_U456, P3_R1200_U457);
  nand ginst22737 (P3_R1200_U104, P3_R1200_U472, P3_R1200_U473);
  nand ginst22738 (P3_R1200_U105, P3_R1200_U477, P3_R1200_U478);
  nand ginst22739 (P3_R1200_U106, P3_R1200_U360, P3_R1200_U361);
  nand ginst22740 (P3_R1200_U107, P3_R1200_U369, P3_R1200_U370);
  nand ginst22741 (P3_R1200_U108, P3_R1200_U376, P3_R1200_U377);
  nand ginst22742 (P3_R1200_U109, P3_R1200_U380, P3_R1200_U381);
  and ginst22743 (P3_R1200_U11, P3_R1200_U191, P3_R1200_U286);
  nand ginst22744 (P3_R1200_U110, P3_R1200_U389, P3_R1200_U390);
  nand ginst22745 (P3_R1200_U111, P3_R1200_U410, P3_R1200_U411);
  nand ginst22746 (P3_R1200_U112, P3_R1200_U427, P3_R1200_U428);
  nand ginst22747 (P3_R1200_U113, P3_R1200_U431, P3_R1200_U432);
  nand ginst22748 (P3_R1200_U114, P3_R1200_U463, P3_R1200_U464);
  nand ginst22749 (P3_R1200_U115, P3_R1200_U467, P3_R1200_U468);
  nand ginst22750 (P3_R1200_U116, P3_R1200_U484, P3_R1200_U485);
  and ginst22751 (P3_R1200_U117, P3_R1200_U193, P3_R1200_U352);
  and ginst22752 (P3_R1200_U118, P3_R1200_U205, P3_R1200_U206);
  and ginst22753 (P3_R1200_U119, P3_R1200_U13, P3_R1200_U14);
  and ginst22754 (P3_R1200_U12, P3_R1200_U287, P3_R1200_U288);
  and ginst22755 (P3_R1200_U120, P3_R1200_U354, P3_R1200_U357);
  and ginst22756 (P3_R1200_U121, P3_R1200_U26, P3_R1200_U362, P3_R1200_U363);
  and ginst22757 (P3_R1200_U122, P3_R1200_U195, P3_R1200_U366);
  and ginst22758 (P3_R1200_U123, P3_R1200_U235, P3_R1200_U6);
  and ginst22759 (P3_R1200_U124, P3_R1200_U194, P3_R1200_U373);
  and ginst22760 (P3_R1200_U125, P3_R1200_U34, P3_R1200_U382, P3_R1200_U383);
  and ginst22761 (P3_R1200_U126, P3_R1200_U193, P3_R1200_U386);
  and ginst22762 (P3_R1200_U127, P3_R1200_U222, P3_R1200_U7);
  and ginst22763 (P3_R1200_U128, P3_R1200_U267, P3_R1200_U9);
  and ginst22764 (P3_R1200_U129, P3_R1200_U11, P3_R1200_U291);
  and ginst22765 (P3_R1200_U13, P3_R1200_U194, P3_R1200_U208, P3_R1200_U213);
  and ginst22766 (P3_R1200_U130, P3_R1200_U192, P3_R1200_U355);
  and ginst22767 (P3_R1200_U131, P3_R1200_U306, P3_R1200_U307);
  and ginst22768 (P3_R1200_U132, P3_R1200_U309, P3_R1200_U395);
  and ginst22769 (P3_R1200_U133, P3_R1200_U306, P3_R1200_U307);
  and ginst22770 (P3_R1200_U134, P3_R1200_U15, P3_R1200_U310);
  nand ginst22771 (P3_R1200_U135, P3_R1200_U398, P3_R1200_U399);
  and ginst22772 (P3_R1200_U136, P3_R1200_U403, P3_R1200_U404, P3_R1200_U87);
  and ginst22773 (P3_R1200_U137, P3_R1200_U192, P3_R1200_U407);
  nand ginst22774 (P3_R1200_U138, P3_R1200_U412, P3_R1200_U413);
  nand ginst22775 (P3_R1200_U139, P3_R1200_U417, P3_R1200_U418);
  and ginst22776 (P3_R1200_U14, P3_R1200_U195, P3_R1200_U218);
  and ginst22777 (P3_R1200_U140, P3_R1200_U12, P3_R1200_U322);
  and ginst22778 (P3_R1200_U141, P3_R1200_U191, P3_R1200_U424);
  nand ginst22779 (P3_R1200_U142, P3_R1200_U433, P3_R1200_U434);
  nand ginst22780 (P3_R1200_U143, P3_R1200_U438, P3_R1200_U439);
  nand ginst22781 (P3_R1200_U144, P3_R1200_U443, P3_R1200_U444);
  nand ginst22782 (P3_R1200_U145, P3_R1200_U448, P3_R1200_U449);
  nand ginst22783 (P3_R1200_U146, P3_R1200_U453, P3_R1200_U454);
  and ginst22784 (P3_R1200_U147, P3_R1200_U10, P3_R1200_U333);
  and ginst22785 (P3_R1200_U148, P3_R1200_U190, P3_R1200_U460);
  nand ginst22786 (P3_R1200_U149, P3_R1200_U469, P3_R1200_U470);
  and ginst22787 (P3_R1200_U15, P3_R1200_U391, P3_R1200_U392);
  nand ginst22788 (P3_R1200_U150, P3_R1200_U474, P3_R1200_U475);
  and ginst22789 (P3_R1200_U151, P3_R1200_U344, P3_R1200_U8);
  and ginst22790 (P3_R1200_U152, P3_R1200_U189, P3_R1200_U481);
  and ginst22791 (P3_R1200_U153, P3_R1200_U358, P3_R1200_U359);
  nand ginst22792 (P3_R1200_U154, P3_R1200_U120, P3_R1200_U356);
  and ginst22793 (P3_R1200_U155, P3_R1200_U367, P3_R1200_U368);
  and ginst22794 (P3_R1200_U156, P3_R1200_U374, P3_R1200_U375);
  and ginst22795 (P3_R1200_U157, P3_R1200_U378, P3_R1200_U379);
  nand ginst22796 (P3_R1200_U158, P3_R1200_U118, P3_R1200_U203);
  and ginst22797 (P3_R1200_U159, P3_R1200_U387, P3_R1200_U388);
  nand ginst22798 (P3_R1200_U16, P3_R1200_U342, P3_R1200_U345);
  not ginst22799 (P3_R1200_U160, P3_U3908);
  not ginst22800 (P3_R1200_U161, P3_U3054);
  and ginst22801 (P3_R1200_U162, P3_R1200_U396, P3_R1200_U397);
  nand ginst22802 (P3_R1200_U163, P3_R1200_U131, P3_R1200_U304);
  and ginst22803 (P3_R1200_U164, P3_R1200_U408, P3_R1200_U409);
  nand ginst22804 (P3_R1200_U165, P3_R1200_U297, P3_R1200_U298);
  nand ginst22805 (P3_R1200_U166, P3_R1200_U293, P3_R1200_U294);
  and ginst22806 (P3_R1200_U167, P3_R1200_U425, P3_R1200_U426);
  and ginst22807 (P3_R1200_U168, P3_R1200_U429, P3_R1200_U430);
  nand ginst22808 (P3_R1200_U169, P3_R1200_U283, P3_R1200_U284);
  nand ginst22809 (P3_R1200_U17, P3_R1200_U331, P3_R1200_U334);
  nand ginst22810 (P3_R1200_U170, P3_R1200_U279, P3_R1200_U280);
  not ginst22811 (P3_R1200_U171, P3_U3392);
  nand ginst22812 (P3_R1200_U172, P3_R1200_U95, P3_U3387);
  nand ginst22813 (P3_R1200_U173, P3_R1200_U184, P3_R1200_U276, P3_R1200_U350);
  not ginst22814 (P3_R1200_U174, P3_U3443);
  nand ginst22815 (P3_R1200_U175, P3_R1200_U273, P3_R1200_U274);
  nand ginst22816 (P3_R1200_U176, P3_R1200_U269, P3_R1200_U270);
  and ginst22817 (P3_R1200_U177, P3_R1200_U461, P3_R1200_U462);
  and ginst22818 (P3_R1200_U178, P3_R1200_U465, P3_R1200_U466);
  nand ginst22819 (P3_R1200_U179, P3_R1200_U259, P3_R1200_U260);
  nand ginst22820 (P3_R1200_U18, P3_R1200_U320, P3_R1200_U323);
  nand ginst22821 (P3_R1200_U180, P3_R1200_U255, P3_R1200_U256);
  nand ginst22822 (P3_R1200_U181, P3_R1200_U251, P3_R1200_U252);
  and ginst22823 (P3_R1200_U182, P3_R1200_U482, P3_R1200_U483);
  nand ginst22824 (P3_R1200_U183, P3_R1200_U132, P3_R1200_U163);
  nand ginst22825 (P3_R1200_U184, P3_R1200_U174, P3_R1200_U175);
  nand ginst22826 (P3_R1200_U185, P3_R1200_U171, P3_R1200_U172);
  not ginst22827 (P3_R1200_U186, P3_R1200_U87);
  not ginst22828 (P3_R1200_U187, P3_R1200_U34);
  not ginst22829 (P3_R1200_U188, P3_R1200_U26);
  nand ginst22830 (P3_R1200_U189, P3_R1200_U54, P3_U3419);
  nand ginst22831 (P3_R1200_U19, P3_R1200_U312, P3_R1200_U314);
  nand ginst22832 (P3_R1200_U190, P3_R1200_U64, P3_U3434);
  nand ginst22833 (P3_R1200_U191, P3_R1200_U78, P3_U3905);
  nand ginst22834 (P3_R1200_U192, P3_R1200_U86, P3_U3901);
  nand ginst22835 (P3_R1200_U193, P3_R1200_U33, P3_U3395);
  nand ginst22836 (P3_R1200_U194, P3_R1200_U41, P3_U3404);
  nand ginst22837 (P3_R1200_U195, P3_R1200_U25, P3_U3410);
  not ginst22838 (P3_R1200_U196, P3_R1200_U66);
  not ginst22839 (P3_R1200_U197, P3_R1200_U80);
  not ginst22840 (P3_R1200_U198, P3_R1200_U43);
  not ginst22841 (P3_R1200_U199, P3_R1200_U55);
  nand ginst22842 (P3_R1200_U20, P3_R1200_U162, P3_R1200_U183, P3_R1200_U351);
  not ginst22843 (P3_R1200_U200, P3_R1200_U172);
  nand ginst22844 (P3_R1200_U201, P3_R1200_U172, P3_U3077);
  not ginst22845 (P3_R1200_U202, P3_R1200_U49);
  nand ginst22846 (P3_R1200_U203, P3_R1200_U117, P3_R1200_U49);
  nand ginst22847 (P3_R1200_U204, P3_R1200_U34, P3_R1200_U35);
  nand ginst22848 (P3_R1200_U205, P3_R1200_U204, P3_R1200_U32);
  nand ginst22849 (P3_R1200_U206, P3_R1200_U187, P3_U3063);
  not ginst22850 (P3_R1200_U207, P3_R1200_U158);
  nand ginst22851 (P3_R1200_U208, P3_R1200_U40, P3_U3407);
  nand ginst22852 (P3_R1200_U209, P3_R1200_U37, P3_U3070);
  nand ginst22853 (P3_R1200_U21, P3_R1200_U241, P3_R1200_U243);
  nand ginst22854 (P3_R1200_U210, P3_R1200_U36, P3_U3066);
  nand ginst22855 (P3_R1200_U211, P3_R1200_U194, P3_R1200_U198);
  nand ginst22856 (P3_R1200_U212, P3_R1200_U211, P3_R1200_U6);
  nand ginst22857 (P3_R1200_U213, P3_R1200_U42, P3_U3401);
  nand ginst22858 (P3_R1200_U214, P3_R1200_U40, P3_U3407);
  nand ginst22859 (P3_R1200_U215, P3_R1200_U13, P3_R1200_U158);
  not ginst22860 (P3_R1200_U216, P3_R1200_U44);
  not ginst22861 (P3_R1200_U217, P3_R1200_U47);
  nand ginst22862 (P3_R1200_U218, P3_R1200_U27, P3_U3413);
  nand ginst22863 (P3_R1200_U219, P3_R1200_U26, P3_R1200_U27);
  nand ginst22864 (P3_R1200_U22, P3_R1200_U233, P3_R1200_U236);
  nand ginst22865 (P3_R1200_U220, P3_R1200_U188, P3_U3083);
  not ginst22866 (P3_R1200_U221, P3_R1200_U154);
  nand ginst22867 (P3_R1200_U222, P3_R1200_U46, P3_U3416);
  nand ginst22868 (P3_R1200_U223, P3_R1200_U222, P3_R1200_U55);
  nand ginst22869 (P3_R1200_U224, P3_R1200_U217, P3_R1200_U26);
  nand ginst22870 (P3_R1200_U225, P3_R1200_U122, P3_R1200_U224);
  nand ginst22871 (P3_R1200_U226, P3_R1200_U195, P3_R1200_U47);
  nand ginst22872 (P3_R1200_U227, P3_R1200_U121, P3_R1200_U226);
  nand ginst22873 (P3_R1200_U228, P3_R1200_U195, P3_R1200_U26);
  nand ginst22874 (P3_R1200_U229, P3_R1200_U158, P3_R1200_U213);
  nand ginst22875 (P3_R1200_U23, P3_R1200_U225, P3_R1200_U227);
  not ginst22876 (P3_R1200_U230, P3_R1200_U48);
  nand ginst22877 (P3_R1200_U231, P3_R1200_U36, P3_U3066);
  nand ginst22878 (P3_R1200_U232, P3_R1200_U230, P3_R1200_U231);
  nand ginst22879 (P3_R1200_U233, P3_R1200_U124, P3_R1200_U232);
  nand ginst22880 (P3_R1200_U234, P3_R1200_U194, P3_R1200_U48);
  nand ginst22881 (P3_R1200_U235, P3_R1200_U40, P3_U3407);
  nand ginst22882 (P3_R1200_U236, P3_R1200_U123, P3_R1200_U234);
  nand ginst22883 (P3_R1200_U237, P3_R1200_U36, P3_U3066);
  nand ginst22884 (P3_R1200_U238, P3_R1200_U194, P3_R1200_U237);
  nand ginst22885 (P3_R1200_U239, P3_R1200_U213, P3_R1200_U43);
  nand ginst22886 (P3_R1200_U24, P3_R1200_U172, P3_R1200_U348);
  nand ginst22887 (P3_R1200_U240, P3_R1200_U202, P3_R1200_U34);
  nand ginst22888 (P3_R1200_U241, P3_R1200_U126, P3_R1200_U240);
  nand ginst22889 (P3_R1200_U242, P3_R1200_U193, P3_R1200_U49);
  nand ginst22890 (P3_R1200_U243, P3_R1200_U125, P3_R1200_U242);
  nand ginst22891 (P3_R1200_U244, P3_R1200_U193, P3_R1200_U34);
  nand ginst22892 (P3_R1200_U245, P3_R1200_U53, P3_U3422);
  nand ginst22893 (P3_R1200_U246, P3_R1200_U51, P3_U3062);
  nand ginst22894 (P3_R1200_U247, P3_R1200_U52, P3_U3061);
  nand ginst22895 (P3_R1200_U248, P3_R1200_U199, P3_R1200_U7);
  nand ginst22896 (P3_R1200_U249, P3_R1200_U248, P3_R1200_U8);
  not ginst22897 (P3_R1200_U25, P3_U3069);
  nand ginst22898 (P3_R1200_U250, P3_R1200_U53, P3_U3422);
  nand ginst22899 (P3_R1200_U251, P3_R1200_U127, P3_R1200_U154);
  nand ginst22900 (P3_R1200_U252, P3_R1200_U249, P3_R1200_U250);
  not ginst22901 (P3_R1200_U253, P3_R1200_U181);
  nand ginst22902 (P3_R1200_U254, P3_R1200_U57, P3_U3425);
  nand ginst22903 (P3_R1200_U255, P3_R1200_U181, P3_R1200_U254);
  nand ginst22904 (P3_R1200_U256, P3_R1200_U56, P3_U3071);
  not ginst22905 (P3_R1200_U257, P3_R1200_U180);
  nand ginst22906 (P3_R1200_U258, P3_R1200_U59, P3_U3428);
  nand ginst22907 (P3_R1200_U259, P3_R1200_U180, P3_R1200_U258);
  nand ginst22908 (P3_R1200_U26, P3_R1200_U39, P3_U3069);
  nand ginst22909 (P3_R1200_U260, P3_R1200_U58, P3_U3079);
  not ginst22910 (P3_R1200_U261, P3_R1200_U179);
  nand ginst22911 (P3_R1200_U262, P3_R1200_U63, P3_U3437);
  nand ginst22912 (P3_R1200_U263, P3_R1200_U60, P3_U3072);
  nand ginst22913 (P3_R1200_U264, P3_R1200_U61, P3_U3073);
  nand ginst22914 (P3_R1200_U265, P3_R1200_U196, P3_R1200_U9);
  nand ginst22915 (P3_R1200_U266, P3_R1200_U10, P3_R1200_U265);
  nand ginst22916 (P3_R1200_U267, P3_R1200_U65, P3_U3431);
  nand ginst22917 (P3_R1200_U268, P3_R1200_U63, P3_U3437);
  nand ginst22918 (P3_R1200_U269, P3_R1200_U128, P3_R1200_U179);
  not ginst22919 (P3_R1200_U27, P3_U3083);
  nand ginst22920 (P3_R1200_U270, P3_R1200_U266, P3_R1200_U268);
  not ginst22921 (P3_R1200_U271, P3_R1200_U176);
  nand ginst22922 (P3_R1200_U272, P3_R1200_U68, P3_U3440);
  nand ginst22923 (P3_R1200_U273, P3_R1200_U176, P3_R1200_U272);
  nand ginst22924 (P3_R1200_U274, P3_R1200_U67, P3_U3068);
  not ginst22925 (P3_R1200_U275, P3_R1200_U175);
  nand ginst22926 (P3_R1200_U276, P3_R1200_U175, P3_U3081);
  not ginst22927 (P3_R1200_U277, P3_R1200_U173);
  nand ginst22928 (P3_R1200_U278, P3_R1200_U71, P3_U3445);
  nand ginst22929 (P3_R1200_U279, P3_R1200_U173, P3_R1200_U278);
  not ginst22930 (P3_R1200_U28, P3_U3413);
  nand ginst22931 (P3_R1200_U280, P3_R1200_U70, P3_U3080);
  not ginst22932 (P3_R1200_U281, P3_R1200_U170);
  nand ginst22933 (P3_R1200_U282, P3_R1200_U73, P3_U3907);
  nand ginst22934 (P3_R1200_U283, P3_R1200_U170, P3_R1200_U282);
  nand ginst22935 (P3_R1200_U284, P3_R1200_U72, P3_U3075);
  not ginst22936 (P3_R1200_U285, P3_R1200_U169);
  nand ginst22937 (P3_R1200_U286, P3_R1200_U77, P3_U3904);
  nand ginst22938 (P3_R1200_U287, P3_R1200_U74, P3_U3065);
  nand ginst22939 (P3_R1200_U288, P3_R1200_U75, P3_U3060);
  nand ginst22940 (P3_R1200_U289, P3_R1200_U11, P3_R1200_U197);
  not ginst22941 (P3_R1200_U29, P3_U3395);
  nand ginst22942 (P3_R1200_U290, P3_R1200_U12, P3_R1200_U289);
  nand ginst22943 (P3_R1200_U291, P3_R1200_U79, P3_U3906);
  nand ginst22944 (P3_R1200_U292, P3_R1200_U77, P3_U3904);
  nand ginst22945 (P3_R1200_U293, P3_R1200_U129, P3_R1200_U169);
  nand ginst22946 (P3_R1200_U294, P3_R1200_U290, P3_R1200_U292);
  not ginst22947 (P3_R1200_U295, P3_R1200_U166);
  nand ginst22948 (P3_R1200_U296, P3_R1200_U82, P3_U3903);
  nand ginst22949 (P3_R1200_U297, P3_R1200_U166, P3_R1200_U296);
  nand ginst22950 (P3_R1200_U298, P3_R1200_U81, P3_U3064);
  not ginst22951 (P3_R1200_U299, P3_R1200_U165);
  not ginst22952 (P3_R1200_U30, P3_U3387);
  nand ginst22953 (P3_R1200_U300, P3_R1200_U84, P3_U3902);
  nand ginst22954 (P3_R1200_U301, P3_R1200_U165, P3_R1200_U300);
  nand ginst22955 (P3_R1200_U302, P3_R1200_U83, P3_U3057);
  not ginst22956 (P3_R1200_U303, P3_R1200_U91);
  nand ginst22957 (P3_R1200_U304, P3_R1200_U130, P3_R1200_U91);
  nand ginst22958 (P3_R1200_U305, P3_R1200_U87, P3_R1200_U88);
  nand ginst22959 (P3_R1200_U306, P3_R1200_U305, P3_R1200_U85);
  nand ginst22960 (P3_R1200_U307, P3_R1200_U186, P3_U3052);
  not ginst22961 (P3_R1200_U308, P3_R1200_U163);
  nand ginst22962 (P3_R1200_U309, P3_R1200_U90, P3_U3899);
  not ginst22963 (P3_R1200_U31, P3_U3077);
  nand ginst22964 (P3_R1200_U310, P3_R1200_U89, P3_U3053);
  nand ginst22965 (P3_R1200_U311, P3_R1200_U303, P3_R1200_U87);
  nand ginst22966 (P3_R1200_U312, P3_R1200_U137, P3_R1200_U311);
  nand ginst22967 (P3_R1200_U313, P3_R1200_U192, P3_R1200_U91);
  nand ginst22968 (P3_R1200_U314, P3_R1200_U136, P3_R1200_U313);
  nand ginst22969 (P3_R1200_U315, P3_R1200_U192, P3_R1200_U87);
  nand ginst22970 (P3_R1200_U316, P3_R1200_U169, P3_R1200_U291);
  not ginst22971 (P3_R1200_U317, P3_R1200_U92);
  nand ginst22972 (P3_R1200_U318, P3_R1200_U75, P3_U3060);
  nand ginst22973 (P3_R1200_U319, P3_R1200_U317, P3_R1200_U318);
  not ginst22974 (P3_R1200_U32, P3_U3398);
  nand ginst22975 (P3_R1200_U320, P3_R1200_U141, P3_R1200_U319);
  nand ginst22976 (P3_R1200_U321, P3_R1200_U191, P3_R1200_U92);
  nand ginst22977 (P3_R1200_U322, P3_R1200_U77, P3_U3904);
  nand ginst22978 (P3_R1200_U323, P3_R1200_U140, P3_R1200_U321);
  nand ginst22979 (P3_R1200_U324, P3_R1200_U75, P3_U3060);
  nand ginst22980 (P3_R1200_U325, P3_R1200_U191, P3_R1200_U324);
  nand ginst22981 (P3_R1200_U326, P3_R1200_U291, P3_R1200_U80);
  nand ginst22982 (P3_R1200_U327, P3_R1200_U179, P3_R1200_U267);
  not ginst22983 (P3_R1200_U328, P3_R1200_U93);
  nand ginst22984 (P3_R1200_U329, P3_R1200_U61, P3_U3073);
  not ginst22985 (P3_R1200_U33, P3_U3067);
  nand ginst22986 (P3_R1200_U330, P3_R1200_U328, P3_R1200_U329);
  nand ginst22987 (P3_R1200_U331, P3_R1200_U148, P3_R1200_U330);
  nand ginst22988 (P3_R1200_U332, P3_R1200_U190, P3_R1200_U93);
  nand ginst22989 (P3_R1200_U333, P3_R1200_U63, P3_U3437);
  nand ginst22990 (P3_R1200_U334, P3_R1200_U147, P3_R1200_U332);
  nand ginst22991 (P3_R1200_U335, P3_R1200_U61, P3_U3073);
  nand ginst22992 (P3_R1200_U336, P3_R1200_U190, P3_R1200_U335);
  nand ginst22993 (P3_R1200_U337, P3_R1200_U267, P3_R1200_U66);
  nand ginst22994 (P3_R1200_U338, P3_R1200_U154, P3_R1200_U222);
  not ginst22995 (P3_R1200_U339, P3_R1200_U94);
  nand ginst22996 (P3_R1200_U34, P3_R1200_U29, P3_U3067);
  nand ginst22997 (P3_R1200_U340, P3_R1200_U52, P3_U3061);
  nand ginst22998 (P3_R1200_U341, P3_R1200_U339, P3_R1200_U340);
  nand ginst22999 (P3_R1200_U342, P3_R1200_U152, P3_R1200_U341);
  nand ginst23000 (P3_R1200_U343, P3_R1200_U189, P3_R1200_U94);
  nand ginst23001 (P3_R1200_U344, P3_R1200_U53, P3_U3422);
  nand ginst23002 (P3_R1200_U345, P3_R1200_U151, P3_R1200_U343);
  nand ginst23003 (P3_R1200_U346, P3_R1200_U52, P3_U3061);
  nand ginst23004 (P3_R1200_U347, P3_R1200_U189, P3_R1200_U346);
  nand ginst23005 (P3_R1200_U348, P3_R1200_U30, P3_U3076);
  nand ginst23006 (P3_R1200_U349, P3_R1200_U171, P3_U3077);
  not ginst23007 (P3_R1200_U35, P3_U3063);
  nand ginst23008 (P3_R1200_U350, P3_R1200_U174, P3_U3081);
  nand ginst23009 (P3_R1200_U351, P3_R1200_U133, P3_R1200_U134, P3_R1200_U304);
  nand ginst23010 (P3_R1200_U352, P3_R1200_U35, P3_U3398);
  nand ginst23011 (P3_R1200_U353, P3_R1200_U220, P3_U3413);
  nand ginst23012 (P3_R1200_U354, P3_R1200_U219, P3_R1200_U353);
  nand ginst23013 (P3_R1200_U355, P3_R1200_U88, P3_U3900);
  nand ginst23014 (P3_R1200_U356, P3_R1200_U119, P3_R1200_U158);
  nand ginst23015 (P3_R1200_U357, P3_R1200_U14, P3_R1200_U216);
  nand ginst23016 (P3_R1200_U358, P3_R1200_U46, P3_U3416);
  nand ginst23017 (P3_R1200_U359, P3_R1200_U45, P3_U3082);
  not ginst23018 (P3_R1200_U36, P3_U3404);
  nand ginst23019 (P3_R1200_U360, P3_R1200_U154, P3_R1200_U223);
  nand ginst23020 (P3_R1200_U361, P3_R1200_U153, P3_R1200_U221);
  nand ginst23021 (P3_R1200_U362, P3_R1200_U27, P3_U3413);
  nand ginst23022 (P3_R1200_U363, P3_R1200_U28, P3_U3083);
  nand ginst23023 (P3_R1200_U364, P3_R1200_U27, P3_U3413);
  nand ginst23024 (P3_R1200_U365, P3_R1200_U28, P3_U3083);
  nand ginst23025 (P3_R1200_U366, P3_R1200_U364, P3_R1200_U365);
  nand ginst23026 (P3_R1200_U367, P3_R1200_U25, P3_U3410);
  nand ginst23027 (P3_R1200_U368, P3_R1200_U39, P3_U3069);
  nand ginst23028 (P3_R1200_U369, P3_R1200_U228, P3_R1200_U47);
  not ginst23029 (P3_R1200_U37, P3_U3407);
  nand ginst23030 (P3_R1200_U370, P3_R1200_U155, P3_R1200_U217);
  nand ginst23031 (P3_R1200_U371, P3_R1200_U40, P3_U3407);
  nand ginst23032 (P3_R1200_U372, P3_R1200_U37, P3_U3070);
  nand ginst23033 (P3_R1200_U373, P3_R1200_U371, P3_R1200_U372);
  nand ginst23034 (P3_R1200_U374, P3_R1200_U41, P3_U3404);
  nand ginst23035 (P3_R1200_U375, P3_R1200_U36, P3_U3066);
  nand ginst23036 (P3_R1200_U376, P3_R1200_U238, P3_R1200_U48);
  nand ginst23037 (P3_R1200_U377, P3_R1200_U156, P3_R1200_U230);
  nand ginst23038 (P3_R1200_U378, P3_R1200_U42, P3_U3401);
  nand ginst23039 (P3_R1200_U379, P3_R1200_U38, P3_U3059);
  not ginst23040 (P3_R1200_U38, P3_U3401);
  nand ginst23041 (P3_R1200_U380, P3_R1200_U158, P3_R1200_U239);
  nand ginst23042 (P3_R1200_U381, P3_R1200_U157, P3_R1200_U207);
  nand ginst23043 (P3_R1200_U382, P3_R1200_U35, P3_U3398);
  nand ginst23044 (P3_R1200_U383, P3_R1200_U32, P3_U3063);
  nand ginst23045 (P3_R1200_U384, P3_R1200_U35, P3_U3398);
  nand ginst23046 (P3_R1200_U385, P3_R1200_U32, P3_U3063);
  nand ginst23047 (P3_R1200_U386, P3_R1200_U384, P3_R1200_U385);
  nand ginst23048 (P3_R1200_U387, P3_R1200_U33, P3_U3395);
  nand ginst23049 (P3_R1200_U388, P3_R1200_U29, P3_U3067);
  nand ginst23050 (P3_R1200_U389, P3_R1200_U244, P3_R1200_U49);
  not ginst23051 (P3_R1200_U39, P3_U3410);
  nand ginst23052 (P3_R1200_U390, P3_R1200_U159, P3_R1200_U202);
  nand ginst23053 (P3_R1200_U391, P3_R1200_U161, P3_U3908);
  nand ginst23054 (P3_R1200_U392, P3_R1200_U160, P3_U3054);
  nand ginst23055 (P3_R1200_U393, P3_R1200_U161, P3_U3908);
  nand ginst23056 (P3_R1200_U394, P3_R1200_U160, P3_U3054);
  nand ginst23057 (P3_R1200_U395, P3_R1200_U393, P3_R1200_U394);
  nand ginst23058 (P3_R1200_U396, P3_R1200_U395, P3_R1200_U89, P3_U3053);
  nand ginst23059 (P3_R1200_U397, P3_R1200_U15, P3_R1200_U90, P3_U3899);
  nand ginst23060 (P3_R1200_U398, P3_R1200_U90, P3_U3899);
  nand ginst23061 (P3_R1200_U399, P3_R1200_U89, P3_U3053);
  not ginst23062 (P3_R1200_U40, P3_U3070);
  not ginst23063 (P3_R1200_U400, P3_R1200_U135);
  nand ginst23064 (P3_R1200_U401, P3_R1200_U308, P3_R1200_U400);
  nand ginst23065 (P3_R1200_U402, P3_R1200_U135, P3_R1200_U163);
  nand ginst23066 (P3_R1200_U403, P3_R1200_U88, P3_U3900);
  nand ginst23067 (P3_R1200_U404, P3_R1200_U85, P3_U3052);
  nand ginst23068 (P3_R1200_U405, P3_R1200_U88, P3_U3900);
  nand ginst23069 (P3_R1200_U406, P3_R1200_U85, P3_U3052);
  nand ginst23070 (P3_R1200_U407, P3_R1200_U405, P3_R1200_U406);
  nand ginst23071 (P3_R1200_U408, P3_R1200_U86, P3_U3901);
  nand ginst23072 (P3_R1200_U409, P3_R1200_U50, P3_U3056);
  not ginst23073 (P3_R1200_U41, P3_U3066);
  nand ginst23074 (P3_R1200_U410, P3_R1200_U315, P3_R1200_U91);
  nand ginst23075 (P3_R1200_U411, P3_R1200_U164, P3_R1200_U303);
  nand ginst23076 (P3_R1200_U412, P3_R1200_U84, P3_U3902);
  nand ginst23077 (P3_R1200_U413, P3_R1200_U83, P3_U3057);
  not ginst23078 (P3_R1200_U414, P3_R1200_U138);
  nand ginst23079 (P3_R1200_U415, P3_R1200_U299, P3_R1200_U414);
  nand ginst23080 (P3_R1200_U416, P3_R1200_U138, P3_R1200_U165);
  nand ginst23081 (P3_R1200_U417, P3_R1200_U82, P3_U3903);
  nand ginst23082 (P3_R1200_U418, P3_R1200_U81, P3_U3064);
  not ginst23083 (P3_R1200_U419, P3_R1200_U139);
  not ginst23084 (P3_R1200_U42, P3_U3059);
  nand ginst23085 (P3_R1200_U420, P3_R1200_U295, P3_R1200_U419);
  nand ginst23086 (P3_R1200_U421, P3_R1200_U139, P3_R1200_U166);
  nand ginst23087 (P3_R1200_U422, P3_R1200_U77, P3_U3904);
  nand ginst23088 (P3_R1200_U423, P3_R1200_U74, P3_U3065);
  nand ginst23089 (P3_R1200_U424, P3_R1200_U422, P3_R1200_U423);
  nand ginst23090 (P3_R1200_U425, P3_R1200_U78, P3_U3905);
  nand ginst23091 (P3_R1200_U426, P3_R1200_U75, P3_U3060);
  nand ginst23092 (P3_R1200_U427, P3_R1200_U325, P3_R1200_U92);
  nand ginst23093 (P3_R1200_U428, P3_R1200_U167, P3_R1200_U317);
  nand ginst23094 (P3_R1200_U429, P3_R1200_U79, P3_U3906);
  nand ginst23095 (P3_R1200_U43, P3_R1200_U38, P3_U3059);
  nand ginst23096 (P3_R1200_U430, P3_R1200_U76, P3_U3074);
  nand ginst23097 (P3_R1200_U431, P3_R1200_U169, P3_R1200_U326);
  nand ginst23098 (P3_R1200_U432, P3_R1200_U168, P3_R1200_U285);
  nand ginst23099 (P3_R1200_U433, P3_R1200_U73, P3_U3907);
  nand ginst23100 (P3_R1200_U434, P3_R1200_U72, P3_U3075);
  not ginst23101 (P3_R1200_U435, P3_R1200_U142);
  nand ginst23102 (P3_R1200_U436, P3_R1200_U281, P3_R1200_U435);
  nand ginst23103 (P3_R1200_U437, P3_R1200_U142, P3_R1200_U170);
  nand ginst23104 (P3_R1200_U438, P3_R1200_U31, P3_U3392);
  nand ginst23105 (P3_R1200_U439, P3_R1200_U171, P3_U3077);
  nand ginst23106 (P3_R1200_U44, P3_R1200_U212, P3_R1200_U214);
  not ginst23107 (P3_R1200_U440, P3_R1200_U143);
  nand ginst23108 (P3_R1200_U441, P3_R1200_U200, P3_R1200_U440);
  nand ginst23109 (P3_R1200_U442, P3_R1200_U143, P3_R1200_U172);
  nand ginst23110 (P3_R1200_U443, P3_R1200_U71, P3_U3445);
  nand ginst23111 (P3_R1200_U444, P3_R1200_U70, P3_U3080);
  not ginst23112 (P3_R1200_U445, P3_R1200_U144);
  nand ginst23113 (P3_R1200_U446, P3_R1200_U277, P3_R1200_U445);
  nand ginst23114 (P3_R1200_U447, P3_R1200_U144, P3_R1200_U173);
  nand ginst23115 (P3_R1200_U448, P3_R1200_U69, P3_U3443);
  nand ginst23116 (P3_R1200_U449, P3_R1200_U174, P3_U3081);
  not ginst23117 (P3_R1200_U45, P3_U3416);
  not ginst23118 (P3_R1200_U450, P3_R1200_U145);
  nand ginst23119 (P3_R1200_U451, P3_R1200_U275, P3_R1200_U450);
  nand ginst23120 (P3_R1200_U452, P3_R1200_U145, P3_R1200_U175);
  nand ginst23121 (P3_R1200_U453, P3_R1200_U68, P3_U3440);
  nand ginst23122 (P3_R1200_U454, P3_R1200_U67, P3_U3068);
  not ginst23123 (P3_R1200_U455, P3_R1200_U146);
  nand ginst23124 (P3_R1200_U456, P3_R1200_U271, P3_R1200_U455);
  nand ginst23125 (P3_R1200_U457, P3_R1200_U146, P3_R1200_U176);
  nand ginst23126 (P3_R1200_U458, P3_R1200_U63, P3_U3437);
  nand ginst23127 (P3_R1200_U459, P3_R1200_U60, P3_U3072);
  not ginst23128 (P3_R1200_U46, P3_U3082);
  nand ginst23129 (P3_R1200_U460, P3_R1200_U458, P3_R1200_U459);
  nand ginst23130 (P3_R1200_U461, P3_R1200_U64, P3_U3434);
  nand ginst23131 (P3_R1200_U462, P3_R1200_U61, P3_U3073);
  nand ginst23132 (P3_R1200_U463, P3_R1200_U336, P3_R1200_U93);
  nand ginst23133 (P3_R1200_U464, P3_R1200_U177, P3_R1200_U328);
  nand ginst23134 (P3_R1200_U465, P3_R1200_U65, P3_U3431);
  nand ginst23135 (P3_R1200_U466, P3_R1200_U62, P3_U3078);
  nand ginst23136 (P3_R1200_U467, P3_R1200_U179, P3_R1200_U337);
  nand ginst23137 (P3_R1200_U468, P3_R1200_U178, P3_R1200_U261);
  nand ginst23138 (P3_R1200_U469, P3_R1200_U59, P3_U3428);
  nand ginst23139 (P3_R1200_U47, P3_R1200_U215, P3_R1200_U44);
  nand ginst23140 (P3_R1200_U470, P3_R1200_U58, P3_U3079);
  not ginst23141 (P3_R1200_U471, P3_R1200_U149);
  nand ginst23142 (P3_R1200_U472, P3_R1200_U257, P3_R1200_U471);
  nand ginst23143 (P3_R1200_U473, P3_R1200_U149, P3_R1200_U180);
  nand ginst23144 (P3_R1200_U474, P3_R1200_U57, P3_U3425);
  nand ginst23145 (P3_R1200_U475, P3_R1200_U56, P3_U3071);
  not ginst23146 (P3_R1200_U476, P3_R1200_U150);
  nand ginst23147 (P3_R1200_U477, P3_R1200_U253, P3_R1200_U476);
  nand ginst23148 (P3_R1200_U478, P3_R1200_U150, P3_R1200_U181);
  nand ginst23149 (P3_R1200_U479, P3_R1200_U53, P3_U3422);
  nand ginst23150 (P3_R1200_U48, P3_R1200_U229, P3_R1200_U43);
  nand ginst23151 (P3_R1200_U480, P3_R1200_U51, P3_U3062);
  nand ginst23152 (P3_R1200_U481, P3_R1200_U479, P3_R1200_U480);
  nand ginst23153 (P3_R1200_U482, P3_R1200_U54, P3_U3419);
  nand ginst23154 (P3_R1200_U483, P3_R1200_U52, P3_U3061);
  nand ginst23155 (P3_R1200_U484, P3_R1200_U347, P3_R1200_U94);
  nand ginst23156 (P3_R1200_U485, P3_R1200_U182, P3_R1200_U339);
  nand ginst23157 (P3_R1200_U49, P3_R1200_U185, P3_R1200_U201, P3_R1200_U349);
  not ginst23158 (P3_R1200_U50, P3_U3901);
  not ginst23159 (P3_R1200_U51, P3_U3422);
  not ginst23160 (P3_R1200_U52, P3_U3419);
  not ginst23161 (P3_R1200_U53, P3_U3062);
  not ginst23162 (P3_R1200_U54, P3_U3061);
  nand ginst23163 (P3_R1200_U55, P3_R1200_U45, P3_U3082);
  not ginst23164 (P3_R1200_U56, P3_U3425);
  not ginst23165 (P3_R1200_U57, P3_U3071);
  not ginst23166 (P3_R1200_U58, P3_U3428);
  not ginst23167 (P3_R1200_U59, P3_U3079);
  and ginst23168 (P3_R1200_U6, P3_R1200_U209, P3_R1200_U210);
  not ginst23169 (P3_R1200_U60, P3_U3437);
  not ginst23170 (P3_R1200_U61, P3_U3434);
  not ginst23171 (P3_R1200_U62, P3_U3431);
  not ginst23172 (P3_R1200_U63, P3_U3072);
  not ginst23173 (P3_R1200_U64, P3_U3073);
  not ginst23174 (P3_R1200_U65, P3_U3078);
  nand ginst23175 (P3_R1200_U66, P3_R1200_U62, P3_U3078);
  not ginst23176 (P3_R1200_U67, P3_U3440);
  not ginst23177 (P3_R1200_U68, P3_U3068);
  not ginst23178 (P3_R1200_U69, P3_U3081);
  and ginst23179 (P3_R1200_U7, P3_R1200_U189, P3_R1200_U245);
  not ginst23180 (P3_R1200_U70, P3_U3445);
  not ginst23181 (P3_R1200_U71, P3_U3080);
  not ginst23182 (P3_R1200_U72, P3_U3907);
  not ginst23183 (P3_R1200_U73, P3_U3075);
  not ginst23184 (P3_R1200_U74, P3_U3904);
  not ginst23185 (P3_R1200_U75, P3_U3905);
  not ginst23186 (P3_R1200_U76, P3_U3906);
  not ginst23187 (P3_R1200_U77, P3_U3065);
  not ginst23188 (P3_R1200_U78, P3_U3060);
  not ginst23189 (P3_R1200_U79, P3_U3074);
  and ginst23190 (P3_R1200_U8, P3_R1200_U246, P3_R1200_U247);
  nand ginst23191 (P3_R1200_U80, P3_R1200_U76, P3_U3074);
  not ginst23192 (P3_R1200_U81, P3_U3903);
  not ginst23193 (P3_R1200_U82, P3_U3064);
  not ginst23194 (P3_R1200_U83, P3_U3902);
  not ginst23195 (P3_R1200_U84, P3_U3057);
  not ginst23196 (P3_R1200_U85, P3_U3900);
  not ginst23197 (P3_R1200_U86, P3_U3056);
  nand ginst23198 (P3_R1200_U87, P3_R1200_U50, P3_U3056);
  not ginst23199 (P3_R1200_U88, P3_U3052);
  not ginst23200 (P3_R1200_U89, P3_U3899);
  and ginst23201 (P3_R1200_U9, P3_R1200_U190, P3_R1200_U262);
  not ginst23202 (P3_R1200_U90, P3_U3053);
  nand ginst23203 (P3_R1200_U91, P3_R1200_U301, P3_R1200_U302);
  nand ginst23204 (P3_R1200_U92, P3_R1200_U316, P3_R1200_U80);
  nand ginst23205 (P3_R1200_U93, P3_R1200_U327, P3_R1200_U66);
  nand ginst23206 (P3_R1200_U94, P3_R1200_U338, P3_R1200_U55);
  not ginst23207 (P3_R1200_U95, P3_U3076);
  nand ginst23208 (P3_R1200_U96, P3_R1200_U401, P3_R1200_U402);
  nand ginst23209 (P3_R1200_U97, P3_R1200_U415, P3_R1200_U416);
  nand ginst23210 (P3_R1200_U98, P3_R1200_U420, P3_R1200_U421);
  nand ginst23211 (P3_R1200_U99, P3_R1200_U436, P3_R1200_U437);
  not ginst23212 (P3_R1209_U10, P3_REG1_REG_1__SCAN_IN);
  nand ginst23213 (P3_R1209_U100, P3_R1209_U150, P3_R1209_U151);
  nand ginst23214 (P3_R1209_U101, P3_R1209_U146, P3_R1209_U147);
  nand ginst23215 (P3_R1209_U102, P3_R1209_U142, P3_R1209_U143);
  nand ginst23216 (P3_R1209_U103, P3_R1209_U138, P3_R1209_U139);
  not ginst23217 (P3_R1209_U104, P3_R1209_U9);
  nand ginst23218 (P3_R1209_U105, P3_REG1_REG_1__SCAN_IN, P3_R1209_U104);
  nand ginst23219 (P3_R1209_U106, P3_R1209_U105, P3_U3391);
  nand ginst23220 (P3_R1209_U107, P3_R1209_U10, P3_R1209_U9);
  not ginst23221 (P3_R1209_U108, P3_R1209_U94);
  nand ginst23222 (P3_R1209_U109, P3_REG1_REG_2__SCAN_IN, P3_R1209_U13);
  not ginst23223 (P3_R1209_U11, P3_U3391);
  nand ginst23224 (P3_R1209_U110, P3_R1209_U109, P3_R1209_U94);
  nand ginst23225 (P3_R1209_U111, P3_R1209_U12, P3_U3394);
  not ginst23226 (P3_R1209_U112, P3_R1209_U93);
  nand ginst23227 (P3_R1209_U113, P3_REG1_REG_3__SCAN_IN, P3_R1209_U15);
  nand ginst23228 (P3_R1209_U114, P3_R1209_U113, P3_R1209_U93);
  nand ginst23229 (P3_R1209_U115, P3_R1209_U14, P3_U3397);
  not ginst23230 (P3_R1209_U116, P3_R1209_U92);
  nand ginst23231 (P3_R1209_U117, P3_REG1_REG_4__SCAN_IN, P3_R1209_U17);
  nand ginst23232 (P3_R1209_U118, P3_R1209_U117, P3_R1209_U92);
  nand ginst23233 (P3_R1209_U119, P3_R1209_U16, P3_U3400);
  not ginst23234 (P3_R1209_U12, P3_REG1_REG_2__SCAN_IN);
  not ginst23235 (P3_R1209_U120, P3_R1209_U91);
  nand ginst23236 (P3_R1209_U121, P3_REG1_REG_5__SCAN_IN, P3_R1209_U19);
  nand ginst23237 (P3_R1209_U122, P3_R1209_U121, P3_R1209_U91);
  nand ginst23238 (P3_R1209_U123, P3_R1209_U18, P3_U3403);
  not ginst23239 (P3_R1209_U124, P3_R1209_U90);
  nand ginst23240 (P3_R1209_U125, P3_REG1_REG_6__SCAN_IN, P3_R1209_U21);
  nand ginst23241 (P3_R1209_U126, P3_R1209_U125, P3_R1209_U90);
  nand ginst23242 (P3_R1209_U127, P3_R1209_U20, P3_U3406);
  not ginst23243 (P3_R1209_U128, P3_R1209_U89);
  nand ginst23244 (P3_R1209_U129, P3_REG1_REG_7__SCAN_IN, P3_R1209_U23);
  not ginst23245 (P3_R1209_U13, P3_U3394);
  nand ginst23246 (P3_R1209_U130, P3_R1209_U129, P3_R1209_U89);
  nand ginst23247 (P3_R1209_U131, P3_R1209_U22, P3_U3409);
  not ginst23248 (P3_R1209_U132, P3_R1209_U88);
  nand ginst23249 (P3_R1209_U133, P3_REG1_REG_8__SCAN_IN, P3_R1209_U25);
  nand ginst23250 (P3_R1209_U134, P3_R1209_U133, P3_R1209_U88);
  nand ginst23251 (P3_R1209_U135, P3_R1209_U24, P3_U3412);
  not ginst23252 (P3_R1209_U136, P3_R1209_U87);
  nand ginst23253 (P3_R1209_U137, P3_REG1_REG_9__SCAN_IN, P3_R1209_U27);
  nand ginst23254 (P3_R1209_U138, P3_R1209_U137, P3_R1209_U87);
  nand ginst23255 (P3_R1209_U139, P3_R1209_U26, P3_U3415);
  not ginst23256 (P3_R1209_U14, P3_REG1_REG_3__SCAN_IN);
  not ginst23257 (P3_R1209_U140, P3_R1209_U103);
  nand ginst23258 (P3_R1209_U141, P3_REG1_REG_10__SCAN_IN, P3_R1209_U29);
  nand ginst23259 (P3_R1209_U142, P3_R1209_U103, P3_R1209_U141);
  nand ginst23260 (P3_R1209_U143, P3_R1209_U28, P3_U3418);
  not ginst23261 (P3_R1209_U144, P3_R1209_U102);
  nand ginst23262 (P3_R1209_U145, P3_REG1_REG_11__SCAN_IN, P3_R1209_U31);
  nand ginst23263 (P3_R1209_U146, P3_R1209_U102, P3_R1209_U145);
  nand ginst23264 (P3_R1209_U147, P3_R1209_U30, P3_U3421);
  not ginst23265 (P3_R1209_U148, P3_R1209_U101);
  nand ginst23266 (P3_R1209_U149, P3_REG1_REG_12__SCAN_IN, P3_R1209_U33);
  not ginst23267 (P3_R1209_U15, P3_U3397);
  nand ginst23268 (P3_R1209_U150, P3_R1209_U101, P3_R1209_U149);
  nand ginst23269 (P3_R1209_U151, P3_R1209_U32, P3_U3424);
  not ginst23270 (P3_R1209_U152, P3_R1209_U100);
  nand ginst23271 (P3_R1209_U153, P3_REG1_REG_13__SCAN_IN, P3_R1209_U35);
  nand ginst23272 (P3_R1209_U154, P3_R1209_U100, P3_R1209_U153);
  nand ginst23273 (P3_R1209_U155, P3_R1209_U34, P3_U3427);
  not ginst23274 (P3_R1209_U156, P3_R1209_U99);
  nand ginst23275 (P3_R1209_U157, P3_REG1_REG_14__SCAN_IN, P3_R1209_U37);
  nand ginst23276 (P3_R1209_U158, P3_R1209_U157, P3_R1209_U99);
  nand ginst23277 (P3_R1209_U159, P3_R1209_U36, P3_U3430);
  not ginst23278 (P3_R1209_U16, P3_REG1_REG_4__SCAN_IN);
  not ginst23279 (P3_R1209_U160, P3_R1209_U38);
  nand ginst23280 (P3_R1209_U161, P3_REG1_REG_15__SCAN_IN, P3_R1209_U160);
  nand ginst23281 (P3_R1209_U162, P3_R1209_U161, P3_U3433);
  nand ginst23282 (P3_R1209_U163, P3_R1209_U38, P3_R1209_U39);
  not ginst23283 (P3_R1209_U164, P3_R1209_U98);
  nand ginst23284 (P3_R1209_U165, P3_REG1_REG_16__SCAN_IN, P3_R1209_U42);
  nand ginst23285 (P3_R1209_U166, P3_R1209_U165, P3_R1209_U98);
  nand ginst23286 (P3_R1209_U167, P3_R1209_U41, P3_U3436);
  not ginst23287 (P3_R1209_U168, P3_R1209_U97);
  nand ginst23288 (P3_R1209_U169, P3_REG1_REG_17__SCAN_IN, P3_R1209_U44);
  not ginst23289 (P3_R1209_U17, P3_U3400);
  nand ginst23290 (P3_R1209_U170, P3_R1209_U169, P3_R1209_U97);
  nand ginst23291 (P3_R1209_U171, P3_R1209_U43, P3_U3439);
  not ginst23292 (P3_R1209_U172, P3_R1209_U47);
  nand ginst23293 (P3_R1209_U173, P3_R1209_U45, P3_U3442);
  nand ginst23294 (P3_R1209_U174, P3_R1209_U172, P3_R1209_U173);
  nand ginst23295 (P3_R1209_U175, P3_REG1_REG_18__SCAN_IN, P3_R1209_U46);
  nand ginst23296 (P3_R1209_U176, P3_R1209_U174, P3_R1209_U77);
  nand ginst23297 (P3_R1209_U177, P3_REG1_REG_18__SCAN_IN, P3_R1209_U46);
  nand ginst23298 (P3_R1209_U178, P3_R1209_U177, P3_R1209_U47);
  nand ginst23299 (P3_R1209_U179, P3_R1209_U45, P3_U3442);
  not ginst23300 (P3_R1209_U18, P3_REG1_REG_5__SCAN_IN);
  nand ginst23301 (P3_R1209_U180, P3_R1209_U178, P3_R1209_U76);
  nand ginst23302 (P3_R1209_U181, P3_R1209_U8, P3_U3386);
  nand ginst23303 (P3_R1209_U182, P3_REG1_REG_9__SCAN_IN, P3_R1209_U27);
  nand ginst23304 (P3_R1209_U183, P3_R1209_U26, P3_U3415);
  not ginst23305 (P3_R1209_U184, P3_R1209_U67);
  nand ginst23306 (P3_R1209_U185, P3_R1209_U136, P3_R1209_U184);
  nand ginst23307 (P3_R1209_U186, P3_R1209_U67, P3_R1209_U87);
  nand ginst23308 (P3_R1209_U187, P3_REG1_REG_8__SCAN_IN, P3_R1209_U25);
  nand ginst23309 (P3_R1209_U188, P3_R1209_U24, P3_U3412);
  not ginst23310 (P3_R1209_U189, P3_R1209_U68);
  not ginst23311 (P3_R1209_U19, P3_U3403);
  nand ginst23312 (P3_R1209_U190, P3_R1209_U132, P3_R1209_U189);
  nand ginst23313 (P3_R1209_U191, P3_R1209_U68, P3_R1209_U88);
  nand ginst23314 (P3_R1209_U192, P3_REG1_REG_7__SCAN_IN, P3_R1209_U23);
  nand ginst23315 (P3_R1209_U193, P3_R1209_U22, P3_U3409);
  not ginst23316 (P3_R1209_U194, P3_R1209_U69);
  nand ginst23317 (P3_R1209_U195, P3_R1209_U128, P3_R1209_U194);
  nand ginst23318 (P3_R1209_U196, P3_R1209_U69, P3_R1209_U89);
  nand ginst23319 (P3_R1209_U197, P3_REG1_REG_6__SCAN_IN, P3_R1209_U21);
  nand ginst23320 (P3_R1209_U198, P3_R1209_U20, P3_U3406);
  not ginst23321 (P3_R1209_U199, P3_R1209_U70);
  not ginst23322 (P3_R1209_U20, P3_REG1_REG_6__SCAN_IN);
  nand ginst23323 (P3_R1209_U200, P3_R1209_U124, P3_R1209_U199);
  nand ginst23324 (P3_R1209_U201, P3_R1209_U70, P3_R1209_U90);
  nand ginst23325 (P3_R1209_U202, P3_REG1_REG_5__SCAN_IN, P3_R1209_U19);
  nand ginst23326 (P3_R1209_U203, P3_R1209_U18, P3_U3403);
  not ginst23327 (P3_R1209_U204, P3_R1209_U71);
  nand ginst23328 (P3_R1209_U205, P3_R1209_U120, P3_R1209_U204);
  nand ginst23329 (P3_R1209_U206, P3_R1209_U71, P3_R1209_U91);
  nand ginst23330 (P3_R1209_U207, P3_REG1_REG_4__SCAN_IN, P3_R1209_U17);
  nand ginst23331 (P3_R1209_U208, P3_R1209_U16, P3_U3400);
  not ginst23332 (P3_R1209_U209, P3_R1209_U72);
  not ginst23333 (P3_R1209_U21, P3_U3406);
  nand ginst23334 (P3_R1209_U210, P3_R1209_U116, P3_R1209_U209);
  nand ginst23335 (P3_R1209_U211, P3_R1209_U72, P3_R1209_U92);
  nand ginst23336 (P3_R1209_U212, P3_REG1_REG_3__SCAN_IN, P3_R1209_U15);
  nand ginst23337 (P3_R1209_U213, P3_R1209_U14, P3_U3397);
  not ginst23338 (P3_R1209_U214, P3_R1209_U73);
  nand ginst23339 (P3_R1209_U215, P3_R1209_U112, P3_R1209_U214);
  nand ginst23340 (P3_R1209_U216, P3_R1209_U73, P3_R1209_U93);
  nand ginst23341 (P3_R1209_U217, P3_REG1_REG_2__SCAN_IN, P3_R1209_U13);
  nand ginst23342 (P3_R1209_U218, P3_R1209_U12, P3_U3394);
  not ginst23343 (P3_R1209_U219, P3_R1209_U74);
  not ginst23344 (P3_R1209_U22, P3_REG1_REG_7__SCAN_IN);
  nand ginst23345 (P3_R1209_U220, P3_R1209_U108, P3_R1209_U219);
  nand ginst23346 (P3_R1209_U221, P3_R1209_U74, P3_R1209_U94);
  nand ginst23347 (P3_R1209_U222, P3_R1209_U10, P3_R1209_U104);
  nand ginst23348 (P3_R1209_U223, P3_REG1_REG_1__SCAN_IN, P3_R1209_U9);
  not ginst23349 (P3_R1209_U224, P3_R1209_U75);
  nand ginst23350 (P3_R1209_U225, P3_R1209_U224, P3_U3391);
  nand ginst23351 (P3_R1209_U226, P3_R1209_U11, P3_R1209_U75);
  nand ginst23352 (P3_R1209_U227, P3_REG1_REG_19__SCAN_IN, P3_R1209_U96);
  nand ginst23353 (P3_R1209_U228, P3_R1209_U95, P3_U3379);
  nand ginst23354 (P3_R1209_U229, P3_REG1_REG_19__SCAN_IN, P3_R1209_U96);
  not ginst23355 (P3_R1209_U23, P3_U3409);
  nand ginst23356 (P3_R1209_U230, P3_R1209_U95, P3_U3379);
  nand ginst23357 (P3_R1209_U231, P3_R1209_U229, P3_R1209_U230);
  nand ginst23358 (P3_R1209_U232, P3_REG1_REG_18__SCAN_IN, P3_R1209_U46);
  nand ginst23359 (P3_R1209_U233, P3_R1209_U45, P3_U3442);
  not ginst23360 (P3_R1209_U234, P3_R1209_U78);
  nand ginst23361 (P3_R1209_U235, P3_R1209_U172, P3_R1209_U234);
  nand ginst23362 (P3_R1209_U236, P3_R1209_U47, P3_R1209_U78);
  nand ginst23363 (P3_R1209_U237, P3_REG1_REG_17__SCAN_IN, P3_R1209_U44);
  nand ginst23364 (P3_R1209_U238, P3_R1209_U43, P3_U3439);
  not ginst23365 (P3_R1209_U239, P3_R1209_U79);
  not ginst23366 (P3_R1209_U24, P3_REG1_REG_8__SCAN_IN);
  nand ginst23367 (P3_R1209_U240, P3_R1209_U168, P3_R1209_U239);
  nand ginst23368 (P3_R1209_U241, P3_R1209_U79, P3_R1209_U97);
  nand ginst23369 (P3_R1209_U242, P3_REG1_REG_16__SCAN_IN, P3_R1209_U42);
  nand ginst23370 (P3_R1209_U243, P3_R1209_U41, P3_U3436);
  not ginst23371 (P3_R1209_U244, P3_R1209_U80);
  nand ginst23372 (P3_R1209_U245, P3_R1209_U164, P3_R1209_U244);
  nand ginst23373 (P3_R1209_U246, P3_R1209_U80, P3_R1209_U98);
  nand ginst23374 (P3_R1209_U247, P3_R1209_U39, P3_U3433);
  nand ginst23375 (P3_R1209_U248, P3_REG1_REG_15__SCAN_IN, P3_R1209_U40);
  not ginst23376 (P3_R1209_U249, P3_R1209_U81);
  not ginst23377 (P3_R1209_U25, P3_U3412);
  nand ginst23378 (P3_R1209_U250, P3_R1209_U160, P3_R1209_U249);
  nand ginst23379 (P3_R1209_U251, P3_R1209_U38, P3_R1209_U81);
  nand ginst23380 (P3_R1209_U252, P3_REG1_REG_14__SCAN_IN, P3_R1209_U37);
  nand ginst23381 (P3_R1209_U253, P3_R1209_U36, P3_U3430);
  not ginst23382 (P3_R1209_U254, P3_R1209_U82);
  nand ginst23383 (P3_R1209_U255, P3_R1209_U156, P3_R1209_U254);
  nand ginst23384 (P3_R1209_U256, P3_R1209_U82, P3_R1209_U99);
  nand ginst23385 (P3_R1209_U257, P3_REG1_REG_13__SCAN_IN, P3_R1209_U35);
  nand ginst23386 (P3_R1209_U258, P3_R1209_U34, P3_U3427);
  not ginst23387 (P3_R1209_U259, P3_R1209_U83);
  not ginst23388 (P3_R1209_U26, P3_REG1_REG_9__SCAN_IN);
  nand ginst23389 (P3_R1209_U260, P3_R1209_U152, P3_R1209_U259);
  nand ginst23390 (P3_R1209_U261, P3_R1209_U100, P3_R1209_U83);
  nand ginst23391 (P3_R1209_U262, P3_REG1_REG_12__SCAN_IN, P3_R1209_U33);
  nand ginst23392 (P3_R1209_U263, P3_R1209_U32, P3_U3424);
  not ginst23393 (P3_R1209_U264, P3_R1209_U84);
  nand ginst23394 (P3_R1209_U265, P3_R1209_U148, P3_R1209_U264);
  nand ginst23395 (P3_R1209_U266, P3_R1209_U101, P3_R1209_U84);
  nand ginst23396 (P3_R1209_U267, P3_REG1_REG_11__SCAN_IN, P3_R1209_U31);
  nand ginst23397 (P3_R1209_U268, P3_R1209_U30, P3_U3421);
  not ginst23398 (P3_R1209_U269, P3_R1209_U85);
  not ginst23399 (P3_R1209_U27, P3_U3415);
  nand ginst23400 (P3_R1209_U270, P3_R1209_U144, P3_R1209_U269);
  nand ginst23401 (P3_R1209_U271, P3_R1209_U102, P3_R1209_U85);
  nand ginst23402 (P3_R1209_U272, P3_REG1_REG_10__SCAN_IN, P3_R1209_U29);
  nand ginst23403 (P3_R1209_U273, P3_R1209_U28, P3_U3418);
  not ginst23404 (P3_R1209_U274, P3_R1209_U86);
  nand ginst23405 (P3_R1209_U275, P3_R1209_U140, P3_R1209_U274);
  nand ginst23406 (P3_R1209_U276, P3_R1209_U103, P3_R1209_U86);
  not ginst23407 (P3_R1209_U28, P3_REG1_REG_10__SCAN_IN);
  not ginst23408 (P3_R1209_U29, P3_U3418);
  not ginst23409 (P3_R1209_U30, P3_REG1_REG_11__SCAN_IN);
  not ginst23410 (P3_R1209_U31, P3_U3421);
  not ginst23411 (P3_R1209_U32, P3_REG1_REG_12__SCAN_IN);
  not ginst23412 (P3_R1209_U33, P3_U3424);
  not ginst23413 (P3_R1209_U34, P3_REG1_REG_13__SCAN_IN);
  not ginst23414 (P3_R1209_U35, P3_U3427);
  not ginst23415 (P3_R1209_U36, P3_REG1_REG_14__SCAN_IN);
  not ginst23416 (P3_R1209_U37, P3_U3430);
  nand ginst23417 (P3_R1209_U38, P3_R1209_U158, P3_R1209_U159);
  not ginst23418 (P3_R1209_U39, P3_REG1_REG_15__SCAN_IN);
  not ginst23419 (P3_R1209_U40, P3_U3433);
  not ginst23420 (P3_R1209_U41, P3_REG1_REG_16__SCAN_IN);
  not ginst23421 (P3_R1209_U42, P3_U3436);
  not ginst23422 (P3_R1209_U43, P3_REG1_REG_17__SCAN_IN);
  not ginst23423 (P3_R1209_U44, P3_U3439);
  not ginst23424 (P3_R1209_U45, P3_REG1_REG_18__SCAN_IN);
  not ginst23425 (P3_R1209_U46, P3_U3442);
  nand ginst23426 (P3_R1209_U47, P3_R1209_U170, P3_R1209_U171);
  not ginst23427 (P3_R1209_U48, P3_U3386);
  nand ginst23428 (P3_R1209_U49, P3_R1209_U185, P3_R1209_U186);
  nand ginst23429 (P3_R1209_U50, P3_R1209_U190, P3_R1209_U191);
  nand ginst23430 (P3_R1209_U51, P3_R1209_U195, P3_R1209_U196);
  nand ginst23431 (P3_R1209_U52, P3_R1209_U200, P3_R1209_U201);
  nand ginst23432 (P3_R1209_U53, P3_R1209_U205, P3_R1209_U206);
  nand ginst23433 (P3_R1209_U54, P3_R1209_U210, P3_R1209_U211);
  nand ginst23434 (P3_R1209_U55, P3_R1209_U215, P3_R1209_U216);
  nand ginst23435 (P3_R1209_U56, P3_R1209_U220, P3_R1209_U221);
  nand ginst23436 (P3_R1209_U57, P3_R1209_U225, P3_R1209_U226);
  nand ginst23437 (P3_R1209_U58, P3_R1209_U235, P3_R1209_U236);
  nand ginst23438 (P3_R1209_U59, P3_R1209_U240, P3_R1209_U241);
  nand ginst23439 (P3_R1209_U6, P3_R1209_U176, P3_R1209_U180);
  nand ginst23440 (P3_R1209_U60, P3_R1209_U245, P3_R1209_U246);
  nand ginst23441 (P3_R1209_U61, P3_R1209_U250, P3_R1209_U251);
  nand ginst23442 (P3_R1209_U62, P3_R1209_U255, P3_R1209_U256);
  nand ginst23443 (P3_R1209_U63, P3_R1209_U260, P3_R1209_U261);
  nand ginst23444 (P3_R1209_U64, P3_R1209_U265, P3_R1209_U266);
  nand ginst23445 (P3_R1209_U65, P3_R1209_U270, P3_R1209_U271);
  nand ginst23446 (P3_R1209_U66, P3_R1209_U275, P3_R1209_U276);
  nand ginst23447 (P3_R1209_U67, P3_R1209_U182, P3_R1209_U183);
  nand ginst23448 (P3_R1209_U68, P3_R1209_U187, P3_R1209_U188);
  nand ginst23449 (P3_R1209_U69, P3_R1209_U192, P3_R1209_U193);
  nand ginst23450 (P3_R1209_U7, P3_R1209_U181, P3_R1209_U9);
  nand ginst23451 (P3_R1209_U70, P3_R1209_U197, P3_R1209_U198);
  nand ginst23452 (P3_R1209_U71, P3_R1209_U202, P3_R1209_U203);
  nand ginst23453 (P3_R1209_U72, P3_R1209_U207, P3_R1209_U208);
  nand ginst23454 (P3_R1209_U73, P3_R1209_U212, P3_R1209_U213);
  nand ginst23455 (P3_R1209_U74, P3_R1209_U217, P3_R1209_U218);
  nand ginst23456 (P3_R1209_U75, P3_R1209_U222, P3_R1209_U223);
  and ginst23457 (P3_R1209_U76, P3_R1209_U179, P3_R1209_U227, P3_R1209_U228);
  and ginst23458 (P3_R1209_U77, P3_R1209_U175, P3_R1209_U231);
  nand ginst23459 (P3_R1209_U78, P3_R1209_U232, P3_R1209_U233);
  nand ginst23460 (P3_R1209_U79, P3_R1209_U237, P3_R1209_U238);
  not ginst23461 (P3_R1209_U8, P3_REG1_REG_0__SCAN_IN);
  nand ginst23462 (P3_R1209_U80, P3_R1209_U242, P3_R1209_U243);
  nand ginst23463 (P3_R1209_U81, P3_R1209_U247, P3_R1209_U248);
  nand ginst23464 (P3_R1209_U82, P3_R1209_U252, P3_R1209_U253);
  nand ginst23465 (P3_R1209_U83, P3_R1209_U257, P3_R1209_U258);
  nand ginst23466 (P3_R1209_U84, P3_R1209_U262, P3_R1209_U263);
  nand ginst23467 (P3_R1209_U85, P3_R1209_U267, P3_R1209_U268);
  nand ginst23468 (P3_R1209_U86, P3_R1209_U272, P3_R1209_U273);
  nand ginst23469 (P3_R1209_U87, P3_R1209_U134, P3_R1209_U135);
  nand ginst23470 (P3_R1209_U88, P3_R1209_U130, P3_R1209_U131);
  nand ginst23471 (P3_R1209_U89, P3_R1209_U126, P3_R1209_U127);
  nand ginst23472 (P3_R1209_U9, P3_REG1_REG_0__SCAN_IN, P3_R1209_U48);
  nand ginst23473 (P3_R1209_U90, P3_R1209_U122, P3_R1209_U123);
  nand ginst23474 (P3_R1209_U91, P3_R1209_U118, P3_R1209_U119);
  nand ginst23475 (P3_R1209_U92, P3_R1209_U114, P3_R1209_U115);
  nand ginst23476 (P3_R1209_U93, P3_R1209_U110, P3_R1209_U111);
  nand ginst23477 (P3_R1209_U94, P3_R1209_U106, P3_R1209_U107);
  not ginst23478 (P3_R1209_U95, P3_REG1_REG_19__SCAN_IN);
  not ginst23479 (P3_R1209_U96, P3_U3379);
  nand ginst23480 (P3_R1209_U97, P3_R1209_U166, P3_R1209_U167);
  nand ginst23481 (P3_R1209_U98, P3_R1209_U162, P3_R1209_U163);
  nand ginst23482 (P3_R1209_U99, P3_R1209_U154, P3_R1209_U155);
  not ginst23483 (P3_R1212_U10, P3_REG2_REG_1__SCAN_IN);
  nand ginst23484 (P3_R1212_U100, P3_R1212_U150, P3_R1212_U151);
  nand ginst23485 (P3_R1212_U101, P3_R1212_U146, P3_R1212_U147);
  nand ginst23486 (P3_R1212_U102, P3_R1212_U142, P3_R1212_U143);
  nand ginst23487 (P3_R1212_U103, P3_R1212_U138, P3_R1212_U139);
  not ginst23488 (P3_R1212_U104, P3_R1212_U9);
  nand ginst23489 (P3_R1212_U105, P3_REG2_REG_1__SCAN_IN, P3_R1212_U104);
  nand ginst23490 (P3_R1212_U106, P3_R1212_U105, P3_U3391);
  nand ginst23491 (P3_R1212_U107, P3_R1212_U10, P3_R1212_U9);
  not ginst23492 (P3_R1212_U108, P3_R1212_U94);
  nand ginst23493 (P3_R1212_U109, P3_REG2_REG_2__SCAN_IN, P3_R1212_U13);
  not ginst23494 (P3_R1212_U11, P3_U3391);
  nand ginst23495 (P3_R1212_U110, P3_R1212_U109, P3_R1212_U94);
  nand ginst23496 (P3_R1212_U111, P3_R1212_U12, P3_U3394);
  not ginst23497 (P3_R1212_U112, P3_R1212_U93);
  nand ginst23498 (P3_R1212_U113, P3_REG2_REG_3__SCAN_IN, P3_R1212_U15);
  nand ginst23499 (P3_R1212_U114, P3_R1212_U113, P3_R1212_U93);
  nand ginst23500 (P3_R1212_U115, P3_R1212_U14, P3_U3397);
  not ginst23501 (P3_R1212_U116, P3_R1212_U92);
  nand ginst23502 (P3_R1212_U117, P3_REG2_REG_4__SCAN_IN, P3_R1212_U17);
  nand ginst23503 (P3_R1212_U118, P3_R1212_U117, P3_R1212_U92);
  nand ginst23504 (P3_R1212_U119, P3_R1212_U16, P3_U3400);
  not ginst23505 (P3_R1212_U12, P3_REG2_REG_2__SCAN_IN);
  not ginst23506 (P3_R1212_U120, P3_R1212_U91);
  nand ginst23507 (P3_R1212_U121, P3_REG2_REG_5__SCAN_IN, P3_R1212_U19);
  nand ginst23508 (P3_R1212_U122, P3_R1212_U121, P3_R1212_U91);
  nand ginst23509 (P3_R1212_U123, P3_R1212_U18, P3_U3403);
  not ginst23510 (P3_R1212_U124, P3_R1212_U90);
  nand ginst23511 (P3_R1212_U125, P3_REG2_REG_6__SCAN_IN, P3_R1212_U21);
  nand ginst23512 (P3_R1212_U126, P3_R1212_U125, P3_R1212_U90);
  nand ginst23513 (P3_R1212_U127, P3_R1212_U20, P3_U3406);
  not ginst23514 (P3_R1212_U128, P3_R1212_U89);
  nand ginst23515 (P3_R1212_U129, P3_REG2_REG_7__SCAN_IN, P3_R1212_U23);
  not ginst23516 (P3_R1212_U13, P3_U3394);
  nand ginst23517 (P3_R1212_U130, P3_R1212_U129, P3_R1212_U89);
  nand ginst23518 (P3_R1212_U131, P3_R1212_U22, P3_U3409);
  not ginst23519 (P3_R1212_U132, P3_R1212_U88);
  nand ginst23520 (P3_R1212_U133, P3_REG2_REG_8__SCAN_IN, P3_R1212_U25);
  nand ginst23521 (P3_R1212_U134, P3_R1212_U133, P3_R1212_U88);
  nand ginst23522 (P3_R1212_U135, P3_R1212_U24, P3_U3412);
  not ginst23523 (P3_R1212_U136, P3_R1212_U87);
  nand ginst23524 (P3_R1212_U137, P3_REG2_REG_9__SCAN_IN, P3_R1212_U27);
  nand ginst23525 (P3_R1212_U138, P3_R1212_U137, P3_R1212_U87);
  nand ginst23526 (P3_R1212_U139, P3_R1212_U26, P3_U3415);
  not ginst23527 (P3_R1212_U14, P3_REG2_REG_3__SCAN_IN);
  not ginst23528 (P3_R1212_U140, P3_R1212_U103);
  nand ginst23529 (P3_R1212_U141, P3_REG2_REG_10__SCAN_IN, P3_R1212_U29);
  nand ginst23530 (P3_R1212_U142, P3_R1212_U103, P3_R1212_U141);
  nand ginst23531 (P3_R1212_U143, P3_R1212_U28, P3_U3418);
  not ginst23532 (P3_R1212_U144, P3_R1212_U102);
  nand ginst23533 (P3_R1212_U145, P3_REG2_REG_11__SCAN_IN, P3_R1212_U31);
  nand ginst23534 (P3_R1212_U146, P3_R1212_U102, P3_R1212_U145);
  nand ginst23535 (P3_R1212_U147, P3_R1212_U30, P3_U3421);
  not ginst23536 (P3_R1212_U148, P3_R1212_U101);
  nand ginst23537 (P3_R1212_U149, P3_REG2_REG_12__SCAN_IN, P3_R1212_U33);
  not ginst23538 (P3_R1212_U15, P3_U3397);
  nand ginst23539 (P3_R1212_U150, P3_R1212_U101, P3_R1212_U149);
  nand ginst23540 (P3_R1212_U151, P3_R1212_U32, P3_U3424);
  not ginst23541 (P3_R1212_U152, P3_R1212_U100);
  nand ginst23542 (P3_R1212_U153, P3_REG2_REG_13__SCAN_IN, P3_R1212_U35);
  nand ginst23543 (P3_R1212_U154, P3_R1212_U100, P3_R1212_U153);
  nand ginst23544 (P3_R1212_U155, P3_R1212_U34, P3_U3427);
  not ginst23545 (P3_R1212_U156, P3_R1212_U99);
  nand ginst23546 (P3_R1212_U157, P3_REG2_REG_14__SCAN_IN, P3_R1212_U37);
  nand ginst23547 (P3_R1212_U158, P3_R1212_U157, P3_R1212_U99);
  nand ginst23548 (P3_R1212_U159, P3_R1212_U36, P3_U3430);
  not ginst23549 (P3_R1212_U16, P3_REG2_REG_4__SCAN_IN);
  not ginst23550 (P3_R1212_U160, P3_R1212_U38);
  nand ginst23551 (P3_R1212_U161, P3_REG2_REG_15__SCAN_IN, P3_R1212_U160);
  nand ginst23552 (P3_R1212_U162, P3_R1212_U161, P3_U3433);
  nand ginst23553 (P3_R1212_U163, P3_R1212_U38, P3_R1212_U39);
  not ginst23554 (P3_R1212_U164, P3_R1212_U98);
  nand ginst23555 (P3_R1212_U165, P3_REG2_REG_16__SCAN_IN, P3_R1212_U42);
  nand ginst23556 (P3_R1212_U166, P3_R1212_U165, P3_R1212_U98);
  nand ginst23557 (P3_R1212_U167, P3_R1212_U41, P3_U3436);
  not ginst23558 (P3_R1212_U168, P3_R1212_U97);
  nand ginst23559 (P3_R1212_U169, P3_REG2_REG_17__SCAN_IN, P3_R1212_U44);
  not ginst23560 (P3_R1212_U17, P3_U3400);
  nand ginst23561 (P3_R1212_U170, P3_R1212_U169, P3_R1212_U97);
  nand ginst23562 (P3_R1212_U171, P3_R1212_U43, P3_U3439);
  not ginst23563 (P3_R1212_U172, P3_R1212_U47);
  nand ginst23564 (P3_R1212_U173, P3_R1212_U45, P3_U3442);
  nand ginst23565 (P3_R1212_U174, P3_R1212_U172, P3_R1212_U173);
  nand ginst23566 (P3_R1212_U175, P3_REG2_REG_18__SCAN_IN, P3_R1212_U46);
  nand ginst23567 (P3_R1212_U176, P3_R1212_U174, P3_R1212_U77);
  nand ginst23568 (P3_R1212_U177, P3_REG2_REG_18__SCAN_IN, P3_R1212_U46);
  nand ginst23569 (P3_R1212_U178, P3_R1212_U177, P3_R1212_U47);
  nand ginst23570 (P3_R1212_U179, P3_R1212_U45, P3_U3442);
  not ginst23571 (P3_R1212_U18, P3_REG2_REG_5__SCAN_IN);
  nand ginst23572 (P3_R1212_U180, P3_R1212_U178, P3_R1212_U76);
  nand ginst23573 (P3_R1212_U181, P3_R1212_U8, P3_U3386);
  nand ginst23574 (P3_R1212_U182, P3_REG2_REG_9__SCAN_IN, P3_R1212_U27);
  nand ginst23575 (P3_R1212_U183, P3_R1212_U26, P3_U3415);
  not ginst23576 (P3_R1212_U184, P3_R1212_U67);
  nand ginst23577 (P3_R1212_U185, P3_R1212_U136, P3_R1212_U184);
  nand ginst23578 (P3_R1212_U186, P3_R1212_U67, P3_R1212_U87);
  nand ginst23579 (P3_R1212_U187, P3_REG2_REG_8__SCAN_IN, P3_R1212_U25);
  nand ginst23580 (P3_R1212_U188, P3_R1212_U24, P3_U3412);
  not ginst23581 (P3_R1212_U189, P3_R1212_U68);
  not ginst23582 (P3_R1212_U19, P3_U3403);
  nand ginst23583 (P3_R1212_U190, P3_R1212_U132, P3_R1212_U189);
  nand ginst23584 (P3_R1212_U191, P3_R1212_U68, P3_R1212_U88);
  nand ginst23585 (P3_R1212_U192, P3_REG2_REG_7__SCAN_IN, P3_R1212_U23);
  nand ginst23586 (P3_R1212_U193, P3_R1212_U22, P3_U3409);
  not ginst23587 (P3_R1212_U194, P3_R1212_U69);
  nand ginst23588 (P3_R1212_U195, P3_R1212_U128, P3_R1212_U194);
  nand ginst23589 (P3_R1212_U196, P3_R1212_U69, P3_R1212_U89);
  nand ginst23590 (P3_R1212_U197, P3_REG2_REG_6__SCAN_IN, P3_R1212_U21);
  nand ginst23591 (P3_R1212_U198, P3_R1212_U20, P3_U3406);
  not ginst23592 (P3_R1212_U199, P3_R1212_U70);
  not ginst23593 (P3_R1212_U20, P3_REG2_REG_6__SCAN_IN);
  nand ginst23594 (P3_R1212_U200, P3_R1212_U124, P3_R1212_U199);
  nand ginst23595 (P3_R1212_U201, P3_R1212_U70, P3_R1212_U90);
  nand ginst23596 (P3_R1212_U202, P3_REG2_REG_5__SCAN_IN, P3_R1212_U19);
  nand ginst23597 (P3_R1212_U203, P3_R1212_U18, P3_U3403);
  not ginst23598 (P3_R1212_U204, P3_R1212_U71);
  nand ginst23599 (P3_R1212_U205, P3_R1212_U120, P3_R1212_U204);
  nand ginst23600 (P3_R1212_U206, P3_R1212_U71, P3_R1212_U91);
  nand ginst23601 (P3_R1212_U207, P3_REG2_REG_4__SCAN_IN, P3_R1212_U17);
  nand ginst23602 (P3_R1212_U208, P3_R1212_U16, P3_U3400);
  not ginst23603 (P3_R1212_U209, P3_R1212_U72);
  not ginst23604 (P3_R1212_U21, P3_U3406);
  nand ginst23605 (P3_R1212_U210, P3_R1212_U116, P3_R1212_U209);
  nand ginst23606 (P3_R1212_U211, P3_R1212_U72, P3_R1212_U92);
  nand ginst23607 (P3_R1212_U212, P3_REG2_REG_3__SCAN_IN, P3_R1212_U15);
  nand ginst23608 (P3_R1212_U213, P3_R1212_U14, P3_U3397);
  not ginst23609 (P3_R1212_U214, P3_R1212_U73);
  nand ginst23610 (P3_R1212_U215, P3_R1212_U112, P3_R1212_U214);
  nand ginst23611 (P3_R1212_U216, P3_R1212_U73, P3_R1212_U93);
  nand ginst23612 (P3_R1212_U217, P3_REG2_REG_2__SCAN_IN, P3_R1212_U13);
  nand ginst23613 (P3_R1212_U218, P3_R1212_U12, P3_U3394);
  not ginst23614 (P3_R1212_U219, P3_R1212_U74);
  not ginst23615 (P3_R1212_U22, P3_REG2_REG_7__SCAN_IN);
  nand ginst23616 (P3_R1212_U220, P3_R1212_U108, P3_R1212_U219);
  nand ginst23617 (P3_R1212_U221, P3_R1212_U74, P3_R1212_U94);
  nand ginst23618 (P3_R1212_U222, P3_R1212_U10, P3_R1212_U104);
  nand ginst23619 (P3_R1212_U223, P3_REG2_REG_1__SCAN_IN, P3_R1212_U9);
  not ginst23620 (P3_R1212_U224, P3_R1212_U75);
  nand ginst23621 (P3_R1212_U225, P3_R1212_U224, P3_U3391);
  nand ginst23622 (P3_R1212_U226, P3_R1212_U11, P3_R1212_U75);
  nand ginst23623 (P3_R1212_U227, P3_REG2_REG_19__SCAN_IN, P3_R1212_U96);
  nand ginst23624 (P3_R1212_U228, P3_R1212_U95, P3_U3379);
  nand ginst23625 (P3_R1212_U229, P3_REG2_REG_19__SCAN_IN, P3_R1212_U96);
  not ginst23626 (P3_R1212_U23, P3_U3409);
  nand ginst23627 (P3_R1212_U230, P3_R1212_U95, P3_U3379);
  nand ginst23628 (P3_R1212_U231, P3_R1212_U229, P3_R1212_U230);
  nand ginst23629 (P3_R1212_U232, P3_REG2_REG_18__SCAN_IN, P3_R1212_U46);
  nand ginst23630 (P3_R1212_U233, P3_R1212_U45, P3_U3442);
  not ginst23631 (P3_R1212_U234, P3_R1212_U78);
  nand ginst23632 (P3_R1212_U235, P3_R1212_U172, P3_R1212_U234);
  nand ginst23633 (P3_R1212_U236, P3_R1212_U47, P3_R1212_U78);
  nand ginst23634 (P3_R1212_U237, P3_REG2_REG_17__SCAN_IN, P3_R1212_U44);
  nand ginst23635 (P3_R1212_U238, P3_R1212_U43, P3_U3439);
  not ginst23636 (P3_R1212_U239, P3_R1212_U79);
  not ginst23637 (P3_R1212_U24, P3_REG2_REG_8__SCAN_IN);
  nand ginst23638 (P3_R1212_U240, P3_R1212_U168, P3_R1212_U239);
  nand ginst23639 (P3_R1212_U241, P3_R1212_U79, P3_R1212_U97);
  nand ginst23640 (P3_R1212_U242, P3_REG2_REG_16__SCAN_IN, P3_R1212_U42);
  nand ginst23641 (P3_R1212_U243, P3_R1212_U41, P3_U3436);
  not ginst23642 (P3_R1212_U244, P3_R1212_U80);
  nand ginst23643 (P3_R1212_U245, P3_R1212_U164, P3_R1212_U244);
  nand ginst23644 (P3_R1212_U246, P3_R1212_U80, P3_R1212_U98);
  nand ginst23645 (P3_R1212_U247, P3_R1212_U39, P3_U3433);
  nand ginst23646 (P3_R1212_U248, P3_REG2_REG_15__SCAN_IN, P3_R1212_U40);
  not ginst23647 (P3_R1212_U249, P3_R1212_U81);
  not ginst23648 (P3_R1212_U25, P3_U3412);
  nand ginst23649 (P3_R1212_U250, P3_R1212_U160, P3_R1212_U249);
  nand ginst23650 (P3_R1212_U251, P3_R1212_U38, P3_R1212_U81);
  nand ginst23651 (P3_R1212_U252, P3_REG2_REG_14__SCAN_IN, P3_R1212_U37);
  nand ginst23652 (P3_R1212_U253, P3_R1212_U36, P3_U3430);
  not ginst23653 (P3_R1212_U254, P3_R1212_U82);
  nand ginst23654 (P3_R1212_U255, P3_R1212_U156, P3_R1212_U254);
  nand ginst23655 (P3_R1212_U256, P3_R1212_U82, P3_R1212_U99);
  nand ginst23656 (P3_R1212_U257, P3_REG2_REG_13__SCAN_IN, P3_R1212_U35);
  nand ginst23657 (P3_R1212_U258, P3_R1212_U34, P3_U3427);
  not ginst23658 (P3_R1212_U259, P3_R1212_U83);
  not ginst23659 (P3_R1212_U26, P3_REG2_REG_9__SCAN_IN);
  nand ginst23660 (P3_R1212_U260, P3_R1212_U152, P3_R1212_U259);
  nand ginst23661 (P3_R1212_U261, P3_R1212_U100, P3_R1212_U83);
  nand ginst23662 (P3_R1212_U262, P3_REG2_REG_12__SCAN_IN, P3_R1212_U33);
  nand ginst23663 (P3_R1212_U263, P3_R1212_U32, P3_U3424);
  not ginst23664 (P3_R1212_U264, P3_R1212_U84);
  nand ginst23665 (P3_R1212_U265, P3_R1212_U148, P3_R1212_U264);
  nand ginst23666 (P3_R1212_U266, P3_R1212_U101, P3_R1212_U84);
  nand ginst23667 (P3_R1212_U267, P3_REG2_REG_11__SCAN_IN, P3_R1212_U31);
  nand ginst23668 (P3_R1212_U268, P3_R1212_U30, P3_U3421);
  not ginst23669 (P3_R1212_U269, P3_R1212_U85);
  not ginst23670 (P3_R1212_U27, P3_U3415);
  nand ginst23671 (P3_R1212_U270, P3_R1212_U144, P3_R1212_U269);
  nand ginst23672 (P3_R1212_U271, P3_R1212_U102, P3_R1212_U85);
  nand ginst23673 (P3_R1212_U272, P3_REG2_REG_10__SCAN_IN, P3_R1212_U29);
  nand ginst23674 (P3_R1212_U273, P3_R1212_U28, P3_U3418);
  not ginst23675 (P3_R1212_U274, P3_R1212_U86);
  nand ginst23676 (P3_R1212_U275, P3_R1212_U140, P3_R1212_U274);
  nand ginst23677 (P3_R1212_U276, P3_R1212_U103, P3_R1212_U86);
  not ginst23678 (P3_R1212_U28, P3_REG2_REG_10__SCAN_IN);
  not ginst23679 (P3_R1212_U29, P3_U3418);
  not ginst23680 (P3_R1212_U30, P3_REG2_REG_11__SCAN_IN);
  not ginst23681 (P3_R1212_U31, P3_U3421);
  not ginst23682 (P3_R1212_U32, P3_REG2_REG_12__SCAN_IN);
  not ginst23683 (P3_R1212_U33, P3_U3424);
  not ginst23684 (P3_R1212_U34, P3_REG2_REG_13__SCAN_IN);
  not ginst23685 (P3_R1212_U35, P3_U3427);
  not ginst23686 (P3_R1212_U36, P3_REG2_REG_14__SCAN_IN);
  not ginst23687 (P3_R1212_U37, P3_U3430);
  nand ginst23688 (P3_R1212_U38, P3_R1212_U158, P3_R1212_U159);
  not ginst23689 (P3_R1212_U39, P3_REG2_REG_15__SCAN_IN);
  not ginst23690 (P3_R1212_U40, P3_U3433);
  not ginst23691 (P3_R1212_U41, P3_REG2_REG_16__SCAN_IN);
  not ginst23692 (P3_R1212_U42, P3_U3436);
  not ginst23693 (P3_R1212_U43, P3_REG2_REG_17__SCAN_IN);
  not ginst23694 (P3_R1212_U44, P3_U3439);
  not ginst23695 (P3_R1212_U45, P3_REG2_REG_18__SCAN_IN);
  not ginst23696 (P3_R1212_U46, P3_U3442);
  nand ginst23697 (P3_R1212_U47, P3_R1212_U170, P3_R1212_U171);
  not ginst23698 (P3_R1212_U48, P3_U3386);
  nand ginst23699 (P3_R1212_U49, P3_R1212_U185, P3_R1212_U186);
  nand ginst23700 (P3_R1212_U50, P3_R1212_U190, P3_R1212_U191);
  nand ginst23701 (P3_R1212_U51, P3_R1212_U195, P3_R1212_U196);
  nand ginst23702 (P3_R1212_U52, P3_R1212_U200, P3_R1212_U201);
  nand ginst23703 (P3_R1212_U53, P3_R1212_U205, P3_R1212_U206);
  nand ginst23704 (P3_R1212_U54, P3_R1212_U210, P3_R1212_U211);
  nand ginst23705 (P3_R1212_U55, P3_R1212_U215, P3_R1212_U216);
  nand ginst23706 (P3_R1212_U56, P3_R1212_U220, P3_R1212_U221);
  nand ginst23707 (P3_R1212_U57, P3_R1212_U225, P3_R1212_U226);
  nand ginst23708 (P3_R1212_U58, P3_R1212_U235, P3_R1212_U236);
  nand ginst23709 (P3_R1212_U59, P3_R1212_U240, P3_R1212_U241);
  nand ginst23710 (P3_R1212_U6, P3_R1212_U176, P3_R1212_U180);
  nand ginst23711 (P3_R1212_U60, P3_R1212_U245, P3_R1212_U246);
  nand ginst23712 (P3_R1212_U61, P3_R1212_U250, P3_R1212_U251);
  nand ginst23713 (P3_R1212_U62, P3_R1212_U255, P3_R1212_U256);
  nand ginst23714 (P3_R1212_U63, P3_R1212_U260, P3_R1212_U261);
  nand ginst23715 (P3_R1212_U64, P3_R1212_U265, P3_R1212_U266);
  nand ginst23716 (P3_R1212_U65, P3_R1212_U270, P3_R1212_U271);
  nand ginst23717 (P3_R1212_U66, P3_R1212_U275, P3_R1212_U276);
  nand ginst23718 (P3_R1212_U67, P3_R1212_U182, P3_R1212_U183);
  nand ginst23719 (P3_R1212_U68, P3_R1212_U187, P3_R1212_U188);
  nand ginst23720 (P3_R1212_U69, P3_R1212_U192, P3_R1212_U193);
  nand ginst23721 (P3_R1212_U7, P3_R1212_U181, P3_R1212_U9);
  nand ginst23722 (P3_R1212_U70, P3_R1212_U197, P3_R1212_U198);
  nand ginst23723 (P3_R1212_U71, P3_R1212_U202, P3_R1212_U203);
  nand ginst23724 (P3_R1212_U72, P3_R1212_U207, P3_R1212_U208);
  nand ginst23725 (P3_R1212_U73, P3_R1212_U212, P3_R1212_U213);
  nand ginst23726 (P3_R1212_U74, P3_R1212_U217, P3_R1212_U218);
  nand ginst23727 (P3_R1212_U75, P3_R1212_U222, P3_R1212_U223);
  and ginst23728 (P3_R1212_U76, P3_R1212_U179, P3_R1212_U227, P3_R1212_U228);
  and ginst23729 (P3_R1212_U77, P3_R1212_U175, P3_R1212_U231);
  nand ginst23730 (P3_R1212_U78, P3_R1212_U232, P3_R1212_U233);
  nand ginst23731 (P3_R1212_U79, P3_R1212_U237, P3_R1212_U238);
  not ginst23732 (P3_R1212_U8, P3_REG2_REG_0__SCAN_IN);
  nand ginst23733 (P3_R1212_U80, P3_R1212_U242, P3_R1212_U243);
  nand ginst23734 (P3_R1212_U81, P3_R1212_U247, P3_R1212_U248);
  nand ginst23735 (P3_R1212_U82, P3_R1212_U252, P3_R1212_U253);
  nand ginst23736 (P3_R1212_U83, P3_R1212_U257, P3_R1212_U258);
  nand ginst23737 (P3_R1212_U84, P3_R1212_U262, P3_R1212_U263);
  nand ginst23738 (P3_R1212_U85, P3_R1212_U267, P3_R1212_U268);
  nand ginst23739 (P3_R1212_U86, P3_R1212_U272, P3_R1212_U273);
  nand ginst23740 (P3_R1212_U87, P3_R1212_U134, P3_R1212_U135);
  nand ginst23741 (P3_R1212_U88, P3_R1212_U130, P3_R1212_U131);
  nand ginst23742 (P3_R1212_U89, P3_R1212_U126, P3_R1212_U127);
  nand ginst23743 (P3_R1212_U9, P3_REG2_REG_0__SCAN_IN, P3_R1212_U48);
  nand ginst23744 (P3_R1212_U90, P3_R1212_U122, P3_R1212_U123);
  nand ginst23745 (P3_R1212_U91, P3_R1212_U118, P3_R1212_U119);
  nand ginst23746 (P3_R1212_U92, P3_R1212_U114, P3_R1212_U115);
  nand ginst23747 (P3_R1212_U93, P3_R1212_U110, P3_R1212_U111);
  nand ginst23748 (P3_R1212_U94, P3_R1212_U106, P3_R1212_U107);
  not ginst23749 (P3_R1212_U95, P3_REG2_REG_19__SCAN_IN);
  not ginst23750 (P3_R1212_U96, P3_U3379);
  nand ginst23751 (P3_R1212_U97, P3_R1212_U166, P3_R1212_U167);
  nand ginst23752 (P3_R1212_U98, P3_R1212_U162, P3_R1212_U163);
  nand ginst23753 (P3_R1212_U99, P3_R1212_U154, P3_R1212_U155);
  and ginst23754 (P3_R1269_U10, P3_R1269_U201, P3_R1269_U202);
  not ginst23755 (P3_R1269_U100, P3_U3084);
  not ginst23756 (P3_R1269_U101, P3_U3085);
  nand ginst23757 (P3_R1269_U102, P3_R1269_U187, P3_R1269_U195);
  nand ginst23758 (P3_R1269_U103, P3_R1269_U56, P3_U3094);
  nand ginst23759 (P3_R1269_U104, P3_R1269_U55, P3_U3095);
  nand ginst23760 (P3_R1269_U105, P3_R1269_U48, P3_U3130);
  nand ginst23761 (P3_R1269_U106, P3_R1269_U35, P3_U3106);
  nand ginst23762 (P3_R1269_U107, P3_R1269_U41, P3_U3135);
  nand ginst23763 (P3_R1269_U108, P3_R1269_U39, P3_U3136);
  nand ginst23764 (P3_R1269_U109, P3_R1269_U34, P3_U3107);
  nand ginst23765 (P3_R1269_U11, P3_R1269_U10, P3_R1269_U194, P3_R1269_U196);
  nand ginst23766 (P3_R1269_U110, P3_R1269_U27, P3_U3112);
  nand ginst23767 (P3_R1269_U111, P3_R1269_U26, P3_U3113);
  nand ginst23768 (P3_R1269_U112, P3_U3147, P3_U3148);
  nand ginst23769 (P3_R1269_U113, P3_R1269_U112, P3_U3115);
  or ginst23770 (P3_R1269_U114, P3_U3147, P3_U3148);
  nand ginst23771 (P3_R1269_U115, P3_R1269_U25, P3_U3114);
  nand ginst23772 (P3_R1269_U116, P3_R1269_U110, P3_R1269_U111, P3_R1269_U113, P3_R1269_U114, P3_R1269_U115);
  nand ginst23773 (P3_R1269_U117, P3_R1269_U31, P3_U3142);
  nand ginst23774 (P3_R1269_U118, P3_R1269_U30, P3_U3141);
  nand ginst23775 (P3_R1269_U119, P3_R1269_U22, P3_U3146);
  not ginst23776 (P3_R1269_U12, P3_U3116);
  nand ginst23777 (P3_R1269_U120, P3_R1269_U21, P3_U3145);
  nand ginst23778 (P3_R1269_U121, P3_R1269_U119, P3_R1269_U120);
  nand ginst23779 (P3_R1269_U122, P3_R1269_U121, P3_R1269_U73);
  nand ginst23780 (P3_R1269_U123, P3_R1269_U20, P3_U3144);
  nand ginst23781 (P3_R1269_U124, P3_R1269_U29, P3_U3143);
  nand ginst23782 (P3_R1269_U125, P3_R1269_U116, P3_R1269_U122, P3_R1269_U123, P3_R1269_U74);
  nand ginst23783 (P3_R1269_U126, P3_R1269_U7, P3_R1269_U75);
  nand ginst23784 (P3_R1269_U127, P3_R1269_U24, P3_U3109);
  nand ginst23785 (P3_R1269_U128, P3_R1269_U30, P3_U3141);
  nand ginst23786 (P3_R1269_U129, P3_R1269_U128, P3_R1269_U76);
  not ginst23787 (P3_R1269_U13, P3_U3094);
  nand ginst23788 (P3_R1269_U130, P3_R1269_U33, P3_U3108);
  nand ginst23789 (P3_R1269_U131, P3_R1269_U125, P3_R1269_U77);
  nand ginst23790 (P3_R1269_U132, P3_R1269_U32, P3_U3140);
  nand ginst23791 (P3_R1269_U133, P3_R1269_U131, P3_R1269_U132);
  nand ginst23792 (P3_R1269_U134, P3_R1269_U109, P3_R1269_U133);
  nand ginst23793 (P3_R1269_U135, P3_R1269_U19, P3_U3139);
  nand ginst23794 (P3_R1269_U136, P3_R1269_U134, P3_R1269_U135);
  nand ginst23795 (P3_R1269_U137, P3_R1269_U106, P3_R1269_U136);
  nand ginst23796 (P3_R1269_U138, P3_R1269_U18, P3_U3138);
  nand ginst23797 (P3_R1269_U139, P3_R1269_U40, P3_U3137);
  not ginst23798 (P3_R1269_U14, P3_U3095);
  nand ginst23799 (P3_R1269_U140, P3_R1269_U137, P3_R1269_U79);
  nand ginst23800 (P3_R1269_U141, P3_R1269_U44, P3_U3101);
  nand ginst23801 (P3_R1269_U142, P3_R1269_U45, P3_U3100);
  nand ginst23802 (P3_R1269_U143, P3_R1269_U107, P3_R1269_U81);
  nand ginst23803 (P3_R1269_U144, P3_R1269_U6, P3_R1269_U82);
  nand ginst23804 (P3_R1269_U145, P3_R1269_U17, P3_U3103);
  nand ginst23805 (P3_R1269_U146, P3_R1269_U43, P3_U3102);
  nand ginst23806 (P3_R1269_U147, P3_R1269_U140, P3_R1269_U83);
  nand ginst23807 (P3_R1269_U148, P3_R1269_U8, P3_R1269_U86);
  nand ginst23808 (P3_R1269_U149, P3_R1269_U45, P3_U3100);
  not ginst23809 (P3_R1269_U15, P3_U3130);
  nand ginst23810 (P3_R1269_U150, P3_R1269_U149, P3_R1269_U87);
  nand ginst23811 (P3_R1269_U151, P3_R1269_U38, P3_U3132);
  nand ginst23812 (P3_R1269_U152, P3_R1269_U47, P3_U3131);
  nand ginst23813 (P3_R1269_U153, P3_R1269_U147, P3_R1269_U88);
  nand ginst23814 (P3_R1269_U154, P3_R1269_U46, P3_U3099);
  nand ginst23815 (P3_R1269_U155, P3_R1269_U153, P3_R1269_U154);
  nand ginst23816 (P3_R1269_U156, P3_R1269_U105, P3_R1269_U155);
  nand ginst23817 (P3_R1269_U157, P3_R1269_U15, P3_U3098);
  not ginst23818 (P3_R1269_U158, P3_R1269_U49);
  nand ginst23819 (P3_R1269_U159, P3_R1269_U158, P3_U3129);
  not ginst23820 (P3_R1269_U16, P3_U3136);
  nand ginst23821 (P3_R1269_U160, P3_R1269_U159, P3_U3097);
  nand ginst23822 (P3_R1269_U161, P3_R1269_U49, P3_R1269_U50);
  nand ginst23823 (P3_R1269_U162, P3_R1269_U54, P3_U3096);
  nand ginst23824 (P3_R1269_U163, P3_R1269_U160, P3_R1269_U90, P3_R1269_U91);
  nand ginst23825 (P3_R1269_U164, P3_R1269_U65, P3_U3123);
  nand ginst23826 (P3_R1269_U165, P3_R1269_U63, P3_U3124);
  nand ginst23827 (P3_R1269_U166, P3_R1269_U104, P3_R1269_U92);
  nand ginst23828 (P3_R1269_U167, P3_R1269_U14, P3_U3127);
  nand ginst23829 (P3_R1269_U168, P3_R1269_U166, P3_R1269_U167);
  nand ginst23830 (P3_R1269_U169, P3_R1269_U103, P3_R1269_U168);
  not ginst23831 (P3_R1269_U17, P3_U3135);
  nand ginst23832 (P3_R1269_U170, P3_R1269_U13, P3_U3126);
  nand ginst23833 (P3_R1269_U171, P3_R1269_U62, P3_U3125);
  nand ginst23834 (P3_R1269_U172, P3_R1269_U163, P3_R1269_U164, P3_R1269_U93);
  nand ginst23835 (P3_R1269_U173, P3_R1269_U67, P3_U3087);
  nand ginst23836 (P3_R1269_U174, P3_R1269_U69, P3_U3089);
  nand ginst23837 (P3_R1269_U175, P3_R1269_U66, P3_U3088);
  nand ginst23838 (P3_R1269_U176, P3_R1269_U71, P3_U3086);
  nand ginst23839 (P3_R1269_U177, P3_R1269_U173, P3_R1269_U97);
  nand ginst23840 (P3_R1269_U178, P3_R1269_U58, P3_U3119);
  not ginst23841 (P3_R1269_U179, P3_R1269_U68);
  not ginst23842 (P3_R1269_U18, P3_U3106);
  nand ginst23843 (P3_R1269_U180, P3_R1269_U59, P3_U3121);
  nand ginst23844 (P3_R1269_U181, P3_R1269_U64, P3_U3122);
  nand ginst23845 (P3_R1269_U182, P3_R1269_U180, P3_R1269_U181);
  nand ginst23846 (P3_R1269_U183, P3_R1269_U179, P3_R1269_U71);
  nand ginst23847 (P3_R1269_U184, P3_R1269_U183, P3_R1269_U61);
  nand ginst23848 (P3_R1269_U185, P3_R1269_U173, P3_R1269_U176, P3_R1269_U182, P3_R1269_U98);
  nand ginst23849 (P3_R1269_U186, P3_R1269_U68, P3_U3118);
  nand ginst23850 (P3_R1269_U187, P3_R1269_U101, P3_R1269_U9);
  nand ginst23851 (P3_R1269_U188, P3_R1269_U57, P3_U3093);
  nand ginst23852 (P3_R1269_U189, P3_R1269_U53, P3_U3092);
  not ginst23853 (P3_R1269_U19, P3_U3107);
  nand ginst23854 (P3_R1269_U190, P3_R1269_U188, P3_R1269_U189);
  nand ginst23855 (P3_R1269_U191, P3_R1269_U164, P3_R1269_U165, P3_R1269_U190);
  nand ginst23856 (P3_R1269_U192, P3_R1269_U70, P3_U3090);
  nand ginst23857 (P3_R1269_U193, P3_R1269_U52, P3_U3091);
  nand ginst23858 (P3_R1269_U194, P3_R1269_U102, P3_R1269_U95);
  nand ginst23859 (P3_R1269_U195, P3_R1269_U9, P3_U3117);
  nand ginst23860 (P3_R1269_U196, P3_R1269_U102, P3_R1269_U197);
  nand ginst23861 (P3_R1269_U197, P3_R1269_U184, P3_R1269_U185, P3_R1269_U99);
  nand ginst23862 (P3_R1269_U198, P3_R1269_U101, P3_U3117);
  nand ginst23863 (P3_R1269_U199, P3_R1269_U12, P3_U3084);
  not ginst23864 (P3_R1269_U20, P3_U3112);
  nand ginst23865 (P3_R1269_U200, P3_R1269_U100, P3_U3116);
  nand ginst23866 (P3_R1269_U201, P3_R1269_U100, P3_R1269_U72, P3_U3116);
  nand ginst23867 (P3_R1269_U202, P3_R1269_U12, P3_U3084, P3_U3149);
  not ginst23868 (P3_R1269_U21, P3_U3113);
  not ginst23869 (P3_R1269_U22, P3_U3114);
  not ginst23870 (P3_R1269_U23, P3_U3142);
  not ginst23871 (P3_R1269_U24, P3_U3141);
  not ginst23872 (P3_R1269_U25, P3_U3146);
  not ginst23873 (P3_R1269_U26, P3_U3145);
  not ginst23874 (P3_R1269_U27, P3_U3144);
  not ginst23875 (P3_R1269_U28, P3_U3143);
  not ginst23876 (P3_R1269_U29, P3_U3111);
  not ginst23877 (P3_R1269_U30, P3_U3109);
  not ginst23878 (P3_R1269_U31, P3_U3110);
  not ginst23879 (P3_R1269_U32, P3_U3108);
  not ginst23880 (P3_R1269_U33, P3_U3140);
  not ginst23881 (P3_R1269_U34, P3_U3139);
  not ginst23882 (P3_R1269_U35, P3_U3138);
  not ginst23883 (P3_R1269_U36, P3_U3137);
  not ginst23884 (P3_R1269_U37, P3_U3101);
  not ginst23885 (P3_R1269_U38, P3_U3100);
  not ginst23886 (P3_R1269_U39, P3_U3104);
  not ginst23887 (P3_R1269_U40, P3_U3105);
  not ginst23888 (P3_R1269_U41, P3_U3103);
  not ginst23889 (P3_R1269_U42, P3_U3102);
  not ginst23890 (P3_R1269_U43, P3_U3134);
  not ginst23891 (P3_R1269_U44, P3_U3133);
  not ginst23892 (P3_R1269_U45, P3_U3132);
  not ginst23893 (P3_R1269_U46, P3_U3131);
  not ginst23894 (P3_R1269_U47, P3_U3099);
  not ginst23895 (P3_R1269_U48, P3_U3098);
  nand ginst23896 (P3_R1269_U49, P3_R1269_U156, P3_R1269_U157);
  not ginst23897 (P3_R1269_U50, P3_U3129);
  not ginst23898 (P3_R1269_U51, P3_U3096);
  not ginst23899 (P3_R1269_U52, P3_U3123);
  not ginst23900 (P3_R1269_U53, P3_U3124);
  not ginst23901 (P3_R1269_U54, P3_U3128);
  not ginst23902 (P3_R1269_U55, P3_U3127);
  not ginst23903 (P3_R1269_U56, P3_U3126);
  not ginst23904 (P3_R1269_U57, P3_U3125);
  not ginst23905 (P3_R1269_U58, P3_U3087);
  not ginst23906 (P3_R1269_U59, P3_U3089);
  and ginst23907 (P3_R1269_U6, P3_R1269_U107, P3_R1269_U108);
  not ginst23908 (P3_R1269_U60, P3_U3088);
  not ginst23909 (P3_R1269_U61, P3_U3086);
  not ginst23910 (P3_R1269_U62, P3_U3093);
  not ginst23911 (P3_R1269_U63, P3_U3092);
  not ginst23912 (P3_R1269_U64, P3_U3090);
  not ginst23913 (P3_R1269_U65, P3_U3091);
  not ginst23914 (P3_R1269_U66, P3_U3120);
  not ginst23915 (P3_R1269_U67, P3_U3119);
  nand ginst23916 (P3_R1269_U68, P3_R1269_U177, P3_R1269_U178);
  not ginst23917 (P3_R1269_U69, P3_U3121);
  and ginst23918 (P3_R1269_U7, P3_R1269_U117, P3_R1269_U118);
  not ginst23919 (P3_R1269_U70, P3_U3122);
  not ginst23920 (P3_R1269_U71, P3_U3118);
  not ginst23921 (P3_R1269_U72, P3_U3149);
  and ginst23922 (P3_R1269_U73, P3_R1269_U110, P3_R1269_U111);
  and ginst23923 (P3_R1269_U74, P3_R1269_U124, P3_R1269_U7);
  and ginst23924 (P3_R1269_U75, P3_R1269_U28, P3_U3111);
  and ginst23925 (P3_R1269_U76, P3_R1269_U23, P3_U3110);
  and ginst23926 (P3_R1269_U77, P3_R1269_U126, P3_R1269_U127, P3_R1269_U78);
  and ginst23927 (P3_R1269_U78, P3_R1269_U129, P3_R1269_U130);
  and ginst23928 (P3_R1269_U79, P3_R1269_U6, P3_R1269_U80);
  and ginst23929 (P3_R1269_U8, P3_R1269_U141, P3_R1269_U142);
  and ginst23930 (P3_R1269_U80, P3_R1269_U138, P3_R1269_U139);
  and ginst23931 (P3_R1269_U81, P3_R1269_U16, P3_U3104);
  and ginst23932 (P3_R1269_U82, P3_R1269_U36, P3_U3105);
  and ginst23933 (P3_R1269_U83, P3_R1269_U143, P3_R1269_U144, P3_R1269_U85);
  and ginst23934 (P3_R1269_U84, P3_R1269_U145, P3_R1269_U146);
  and ginst23935 (P3_R1269_U85, P3_R1269_U8, P3_R1269_U84);
  and ginst23936 (P3_R1269_U86, P3_R1269_U42, P3_U3134);
  and ginst23937 (P3_R1269_U87, P3_R1269_U37, P3_U3133);
  and ginst23938 (P3_R1269_U88, P3_R1269_U148, P3_R1269_U150, P3_R1269_U89);
  and ginst23939 (P3_R1269_U89, P3_R1269_U151, P3_R1269_U152);
  and ginst23940 (P3_R1269_U9, P3_R1269_U199, P3_R1269_U200);
  and ginst23941 (P3_R1269_U90, P3_R1269_U103, P3_R1269_U104);
  and ginst23942 (P3_R1269_U91, P3_R1269_U161, P3_R1269_U162);
  and ginst23943 (P3_R1269_U92, P3_R1269_U51, P3_U3128);
  and ginst23944 (P3_R1269_U93, P3_R1269_U165, P3_R1269_U169, P3_R1269_U170, P3_R1269_U171);
  and ginst23945 (P3_R1269_U94, P3_R1269_U174, P3_R1269_U175);
  and ginst23946 (P3_R1269_U95, P3_R1269_U172, P3_R1269_U173, P3_R1269_U176, P3_R1269_U94, P3_R1269_U96);
  and ginst23947 (P3_R1269_U96, P3_R1269_U191, P3_R1269_U192, P3_R1269_U193);
  and ginst23948 (P3_R1269_U97, P3_R1269_U60, P3_U3120);
  and ginst23949 (P3_R1269_U98, P3_R1269_U174, P3_R1269_U175);
  and ginst23950 (P3_R1269_U99, P3_R1269_U186, P3_R1269_U198);
  and ginst23951 (P3_R1297_U6, P3_R1297_U7, P3_U3058);
  not ginst23952 (P3_R1297_U7, P3_U3055);
  nand ginst23953 (P3_R1300_U10, P3_R1300_U7, P3_U3058);
  not ginst23954 (P3_R1300_U6, P3_U3058);
  not ginst23955 (P3_R1300_U7, P3_U3055);
  and ginst23956 (P3_R1300_U8, P3_R1300_U10, P3_R1300_U9);
  nand ginst23957 (P3_R1300_U9, P3_R1300_U6, P3_U3055);
  and ginst23958 (P3_R693_U10, P3_R693_U130, P3_R693_U131);
  and ginst23959 (P3_R693_U100, P3_R693_U159, P3_R693_U160);
  and ginst23960 (P3_R693_U101, P3_R693_U122, P3_R693_U123, P3_R693_U170, P3_R693_U171);
  and ginst23961 (P3_R693_U102, P3_R693_U174, P3_R693_U175);
  and ginst23962 (P3_R693_U103, P3_R693_U186, P3_R693_U187);
  and ginst23963 (P3_R693_U104, P3_R693_U103, P3_R693_U13);
  and ginst23964 (P3_R693_U105, P3_R693_U106, P3_R693_U190);
  and ginst23965 (P3_R693_U106, P3_R693_U65, P3_U3533);
  and ginst23966 (P3_R693_U107, P3_R693_U63, P3_U3532);
  and ginst23967 (P3_R693_U108, P3_R693_U191, P3_R693_U192);
  and ginst23968 (P3_R693_U109, P3_R693_U193, P3_R693_U194, P3_R693_U195);
  and ginst23969 (P3_R693_U11, P3_R693_U10, P3_R693_U84);
  not ginst23970 (P3_R693_U110, P3_U3873);
  not ginst23971 (P3_R693_U111, P3_U3554);
  nand ginst23972 (P3_R693_U112, P3_R693_U181, P3_R693_U196);
  nand ginst23973 (P3_R693_U113, P3_R693_U26, P3_U3543);
  nand ginst23974 (P3_R693_U114, P3_R693_U23, P3_U3544);
  nand ginst23975 (P3_R693_U115, P3_R693_U61, P3_U3905);
  nand ginst23976 (P3_R693_U116, P3_R693_U19, P3_U3906);
  nand ginst23977 (P3_R693_U117, P3_R693_U113, P3_R693_U78);
  nand ginst23978 (P3_R693_U118, P3_R693_U6, P3_R693_U79);
  nand ginst23979 (P3_R693_U119, P3_R693_U22, P3_U3445);
  and ginst23980 (P3_R693_U12, P3_R693_U141, P3_R693_U142);
  nand ginst23981 (P3_R693_U120, P3_R693_U21, P3_U3907);
  nand ginst23982 (P3_R693_U121, P3_R693_U29, P3_U3437);
  nand ginst23983 (P3_R693_U122, P3_R693_U67, P3_U3537);
  nand ginst23984 (P3_R693_U123, P3_R693_U68, P3_U3536);
  nand ginst23985 (P3_R693_U124, P3_R693_U60, P3_U3434);
  nand ginst23986 (P3_R693_U125, P3_R693_U35, P3_U3526);
  nand ginst23987 (P3_R693_U126, P3_R693_U38, P3_U3525);
  nand ginst23988 (P3_R693_U127, P3_R693_U81, P3_R693_U9);
  nand ginst23989 (P3_R693_U128, P3_R693_U38, P3_U3525);
  nand ginst23990 (P3_R693_U129, P3_R693_U128, P3_R693_U82);
  and ginst23991 (P3_R693_U13, P3_R693_U177, P3_R693_U178, P3_R693_U179);
  nand ginst23992 (P3_R693_U130, P3_R693_U53, P3_U3419);
  nand ginst23993 (P3_R693_U131, P3_R693_U51, P3_U3416);
  nand ginst23994 (P3_R693_U132, P3_R693_U33, P3_U3410);
  nand ginst23995 (P3_R693_U133, P3_R693_U52, P3_U3413);
  nand ginst23996 (P3_R693_U134, P3_R693_U48, P3_U3398);
  nand ginst23997 (P3_R693_U135, P3_R693_U49, P3_U3401);
  nand ginst23998 (P3_R693_U136, P3_R693_U44, P3_U3553);
  nand ginst23999 (P3_R693_U137, P3_R693_U136, P3_R693_U83);
  nand ginst24000 (P3_R693_U138, P3_R693_U47, P3_U3395);
  nand ginst24001 (P3_R693_U139, P3_R693_U42, P3_U3392);
  and ginst24002 (P3_R693_U14, P3_R693_U108, P3_R693_U109, P3_R693_U188, P3_R693_U189);
  nand ginst24003 (P3_R693_U140, P3_R693_U11, P3_R693_U127, P3_R693_U139, P3_R693_U85, P3_R693_U87);
  nand ginst24004 (P3_R693_U141, P3_R693_U55, P3_U3550);
  nand ginst24005 (P3_R693_U142, P3_R693_U58, P3_U3549);
  nand ginst24006 (P3_R693_U143, P3_R693_U43, P3_U3542);
  nand ginst24007 (P3_R693_U144, P3_R693_U40, P3_U3531);
  nand ginst24008 (P3_R693_U145, P3_R693_U143, P3_R693_U144);
  nand ginst24009 (P3_R693_U146, P3_R693_U145, P3_R693_U88);
  nand ginst24010 (P3_R693_U147, P3_R693_U41, P3_U3528);
  nand ginst24011 (P3_R693_U148, P3_R693_U34, P3_U3527);
  nand ginst24012 (P3_R693_U149, P3_R693_U146, P3_R693_U147, P3_R693_U89);
  not ginst24013 (P3_R693_U15, P3_U3529);
  nand ginst24014 (P3_R693_U150, P3_R693_U149, P3_R693_U90);
  nand ginst24015 (P3_R693_U151, P3_R693_U130, P3_R693_U91);
  nand ginst24016 (P3_R693_U152, P3_R693_U10, P3_R693_U92);
  nand ginst24017 (P3_R693_U153, P3_R693_U37, P3_U3552);
  nand ginst24018 (P3_R693_U154, P3_R693_U56, P3_U3551);
  nand ginst24019 (P3_R693_U155, P3_R693_U140, P3_R693_U150, P3_R693_U93);
  nand ginst24020 (P3_R693_U156, P3_R693_U58, P3_U3549);
  nand ginst24021 (P3_R693_U157, P3_R693_U156, P3_R693_U96);
  nand ginst24022 (P3_R693_U158, P3_R693_U12, P3_R693_U97);
  nand ginst24023 (P3_R693_U159, P3_R693_U59, P3_U3431);
  not ginst24024 (P3_R693_U16, P3_U3537);
  nand ginst24025 (P3_R693_U160, P3_R693_U46, P3_U3428);
  nand ginst24026 (P3_R693_U161, P3_R693_U155, P3_R693_U99);
  nand ginst24027 (P3_R693_U162, P3_R693_U57, P3_U3548);
  nand ginst24028 (P3_R693_U163, P3_R693_U161, P3_R693_U162);
  nand ginst24029 (P3_R693_U164, P3_R693_U124, P3_R693_U163);
  nand ginst24030 (P3_R693_U165, P3_R693_U31, P3_U3547);
  nand ginst24031 (P3_R693_U166, P3_R693_U164, P3_R693_U165);
  nand ginst24032 (P3_R693_U167, P3_R693_U25, P3_U3545);
  nand ginst24033 (P3_R693_U168, P3_R693_U30, P3_U3546);
  nand ginst24034 (P3_R693_U169, P3_R693_U6, P3_R693_U77);
  not ginst24035 (P3_R693_U17, P3_U3536);
  nand ginst24036 (P3_R693_U170, P3_R693_U115, P3_R693_U75);
  nand ginst24037 (P3_R693_U171, P3_R693_U7, P3_R693_U76);
  nand ginst24038 (P3_R693_U172, P3_R693_U169, P3_R693_U8);
  nand ginst24039 (P3_R693_U173, P3_R693_U121, P3_R693_U166, P3_R693_U8);
  nand ginst24040 (P3_R693_U174, P3_R693_U18, P3_U3539);
  nand ginst24041 (P3_R693_U175, P3_R693_U66, P3_U3538);
  nand ginst24042 (P3_R693_U176, P3_R693_U101, P3_R693_U102, P3_R693_U172, P3_R693_U173);
  nand ginst24043 (P3_R693_U177, P3_R693_U73, P3_U3908);
  nand ginst24044 (P3_R693_U178, P3_R693_U71, P3_U3900);
  nand ginst24045 (P3_R693_U179, P3_R693_U70, P3_U3899);
  not ginst24046 (P3_R693_U18, P3_U3905);
  nand ginst24047 (P3_R693_U180, P3_R693_U72, P3_U3529);
  nand ginst24048 (P3_R693_U181, P3_R693_U110, P3_R693_U180);
  nand ginst24049 (P3_R693_U182, P3_R693_U62, P3_U3904);
  nand ginst24050 (P3_R693_U183, P3_R693_U16, P3_U3903);
  nand ginst24051 (P3_R693_U184, P3_R693_U182, P3_R693_U183);
  nand ginst24052 (P3_R693_U185, P3_R693_U122, P3_R693_U123, P3_R693_U184);
  nand ginst24053 (P3_R693_U186, P3_R693_U17, P3_U3902);
  nand ginst24054 (P3_R693_U187, P3_R693_U74, P3_U3901);
  nand ginst24055 (P3_R693_U188, P3_R693_U104, P3_R693_U112, P3_R693_U176, P3_R693_U185);
  nand ginst24056 (P3_R693_U189, P3_R693_U110, P3_R693_U180, P3_U3530);
  not ginst24057 (P3_R693_U19, P3_U3540);
  nand ginst24058 (P3_R693_U190, P3_R693_U73, P3_U3908);
  nand ginst24059 (P3_R693_U191, P3_R693_U105, P3_R693_U112);
  nand ginst24060 (P3_R693_U192, P3_R693_U112, P3_R693_U13, P3_R693_U64, P3_U3534);
  nand ginst24061 (P3_R693_U193, P3_R693_U15, P3_U3872);
  nand ginst24062 (P3_R693_U194, P3_R693_U107, P3_R693_U112);
  nand ginst24063 (P3_R693_U195, P3_R693_U112, P3_R693_U13, P3_R693_U69, P3_U3535);
  nand ginst24064 (P3_R693_U196, P3_R693_U180, P3_U3530);
  not ginst24065 (P3_R693_U20, P3_U3906);
  not ginst24066 (P3_R693_U21, P3_U3541);
  not ginst24067 (P3_R693_U22, P3_U3543);
  not ginst24068 (P3_R693_U23, P3_U3443);
  not ginst24069 (P3_R693_U24, P3_U3544);
  not ginst24070 (P3_R693_U25, P3_U3440);
  not ginst24071 (P3_R693_U26, P3_U3445);
  not ginst24072 (P3_R693_U27, P3_U3907);
  not ginst24073 (P3_R693_U28, P3_U3545);
  not ginst24074 (P3_R693_U29, P3_U3546);
  not ginst24075 (P3_R693_U30, P3_U3437);
  not ginst24076 (P3_R693_U31, P3_U3434);
  not ginst24077 (P3_R693_U32, P3_U3526);
  not ginst24078 (P3_R693_U33, P3_U3525);
  not ginst24079 (P3_R693_U34, P3_U3404);
  not ginst24080 (P3_R693_U35, P3_U3407);
  not ginst24081 (P3_R693_U36, P3_U3416);
  not ginst24082 (P3_R693_U37, P3_U3419);
  not ginst24083 (P3_R693_U38, P3_U3410);
  not ginst24084 (P3_R693_U39, P3_U3413);
  not ginst24085 (P3_R693_U40, P3_U3398);
  not ginst24086 (P3_R693_U41, P3_U3401);
  not ginst24087 (P3_R693_U42, P3_U3553);
  not ginst24088 (P3_R693_U43, P3_U3395);
  not ginst24089 (P3_R693_U44, P3_U3392);
  not ginst24090 (P3_R693_U45, P3_U3550);
  not ginst24091 (P3_R693_U46, P3_U3549);
  not ginst24092 (P3_R693_U47, P3_U3542);
  not ginst24093 (P3_R693_U48, P3_U3531);
  not ginst24094 (P3_R693_U49, P3_U3528);
  not ginst24095 (P3_R693_U50, P3_U3527);
  not ginst24096 (P3_R693_U51, P3_U3523);
  not ginst24097 (P3_R693_U52, P3_U3524);
  not ginst24098 (P3_R693_U53, P3_U3552);
  not ginst24099 (P3_R693_U54, P3_U3551);
  not ginst24100 (P3_R693_U55, P3_U3425);
  not ginst24101 (P3_R693_U56, P3_U3422);
  not ginst24102 (P3_R693_U57, P3_U3431);
  not ginst24103 (P3_R693_U58, P3_U3428);
  not ginst24104 (P3_R693_U59, P3_U3548);
  and ginst24105 (P3_R693_U6, P3_R693_U113, P3_R693_U114);
  not ginst24106 (P3_R693_U60, P3_U3547);
  not ginst24107 (P3_R693_U61, P3_U3539);
  not ginst24108 (P3_R693_U62, P3_U3538);
  not ginst24109 (P3_R693_U63, P3_U3908);
  not ginst24110 (P3_R693_U64, P3_U3900);
  not ginst24111 (P3_R693_U65, P3_U3899);
  not ginst24112 (P3_R693_U66, P3_U3904);
  not ginst24113 (P3_R693_U67, P3_U3903);
  not ginst24114 (P3_R693_U68, P3_U3902);
  not ginst24115 (P3_R693_U69, P3_U3901);
  and ginst24116 (P3_R693_U7, P3_R693_U115, P3_R693_U116);
  not ginst24117 (P3_R693_U70, P3_U3533);
  not ginst24118 (P3_R693_U71, P3_U3534);
  not ginst24119 (P3_R693_U72, P3_U3872);
  not ginst24120 (P3_R693_U73, P3_U3532);
  not ginst24121 (P3_R693_U74, P3_U3535);
  and ginst24122 (P3_R693_U75, P3_R693_U20, P3_U3540);
  and ginst24123 (P3_R693_U76, P3_R693_U27, P3_U3541);
  and ginst24124 (P3_R693_U77, P3_R693_U167, P3_R693_U168);
  and ginst24125 (P3_R693_U78, P3_R693_U24, P3_U3443);
  and ginst24126 (P3_R693_U79, P3_R693_U28, P3_U3440);
  and ginst24127 (P3_R693_U8, P3_R693_U118, P3_R693_U120, P3_R693_U7, P3_R693_U80);
  and ginst24128 (P3_R693_U80, P3_R693_U117, P3_R693_U119);
  and ginst24129 (P3_R693_U81, P3_R693_U50, P3_U3404);
  and ginst24130 (P3_R693_U82, P3_R693_U32, P3_U3407);
  and ginst24131 (P3_R693_U83, P3_R693_U111, P3_U3387);
  and ginst24132 (P3_R693_U84, P3_R693_U132, P3_R693_U133);
  and ginst24133 (P3_R693_U85, P3_R693_U129, P3_R693_U86);
  and ginst24134 (P3_R693_U86, P3_R693_U134, P3_R693_U135);
  and ginst24135 (P3_R693_U87, P3_R693_U137, P3_R693_U138);
  and ginst24136 (P3_R693_U88, P3_R693_U134, P3_R693_U135);
  and ginst24137 (P3_R693_U89, P3_R693_U148, P3_R693_U9);
  and ginst24138 (P3_R693_U9, P3_R693_U125, P3_R693_U126);
  and ginst24139 (P3_R693_U90, P3_R693_U11, P3_R693_U127, P3_R693_U129);
  and ginst24140 (P3_R693_U91, P3_R693_U36, P3_U3523);
  and ginst24141 (P3_R693_U92, P3_R693_U39, P3_U3524);
  and ginst24142 (P3_R693_U93, P3_R693_U151, P3_R693_U152, P3_R693_U95);
  and ginst24143 (P3_R693_U94, P3_R693_U153, P3_R693_U154);
  and ginst24144 (P3_R693_U95, P3_R693_U12, P3_R693_U94);
  and ginst24145 (P3_R693_U96, P3_R693_U45, P3_U3425);
  and ginst24146 (P3_R693_U97, P3_R693_U54, P3_U3422);
  and ginst24147 (P3_R693_U98, P3_R693_U100, P3_R693_U157);
  and ginst24148 (P3_R693_U99, P3_R693_U158, P3_R693_U98);
  and ginst24149 (P3_SUB_598_U10, P3_SUB_598_U132, P3_SUB_598_U47);
  nand ginst24150 (P3_SUB_598_U100, P3_IR_REG_3__SCAN_IN, P3_SUB_598_U28);
  not ginst24151 (P3_SUB_598_U101, P3_SUB_598_U49);
  nand ginst24152 (P3_SUB_598_U102, P3_SUB_598_U101, P3_SUB_598_U50);
  not ginst24153 (P3_SUB_598_U103, P3_SUB_598_U46);
  not ginst24154 (P3_SUB_598_U104, P3_SUB_598_U47);
  nand ginst24155 (P3_SUB_598_U105, P3_SUB_598_U104, P3_SUB_598_U48);
  not ginst24156 (P3_SUB_598_U106, P3_SUB_598_U34);
  not ginst24157 (P3_SUB_598_U107, P3_SUB_598_U44);
  nand ginst24158 (P3_SUB_598_U108, P3_SUB_598_U107, P3_SUB_598_U45);
  not ginst24159 (P3_SUB_598_U109, P3_SUB_598_U40);
  and ginst24160 (P3_SUB_598_U11, P3_SUB_598_U105, P3_SUB_598_U130);
  not ginst24161 (P3_SUB_598_U110, P3_SUB_598_U41);
  nand ginst24162 (P3_SUB_598_U111, P3_SUB_598_U110, P3_SUB_598_U43);
  not ginst24163 (P3_SUB_598_U112, P3_SUB_598_U35);
  not ginst24164 (P3_SUB_598_U113, P3_SUB_598_U78);
  not ginst24165 (P3_SUB_598_U114, P3_SUB_598_U36);
  not ginst24166 (P3_SUB_598_U115, P3_SUB_598_U37);
  or ginst24167 (P3_SUB_598_U116, P3_IR_REG_0__SCAN_IN, P3_IR_REG_1__SCAN_IN);
  nand ginst24168 (P3_SUB_598_U117, P3_IR_REG_2__SCAN_IN, P3_SUB_598_U116);
  nand ginst24169 (P3_SUB_598_U118, P3_IR_REG_29__SCAN_IN, P3_SUB_598_U36);
  nand ginst24170 (P3_SUB_598_U119, P3_SUB_598_U112, P3_SUB_598_U80);
  and ginst24171 (P3_SUB_598_U12, P3_SUB_598_U129, P3_SUB_598_U34);
  nand ginst24172 (P3_SUB_598_U120, P3_IR_REG_26__SCAN_IN, P3_SUB_598_U119);
  nand ginst24173 (P3_SUB_598_U121, P3_IR_REG_24__SCAN_IN, P3_SUB_598_U111);
  nand ginst24174 (P3_SUB_598_U122, P3_IR_REG_23__SCAN_IN, P3_SUB_598_U41);
  nand ginst24175 (P3_SUB_598_U123, P3_SUB_598_U109, P3_SUB_598_U82);
  nand ginst24176 (P3_SUB_598_U124, P3_IR_REG_22__SCAN_IN, P3_SUB_598_U123);
  nand ginst24177 (P3_SUB_598_U125, P3_IR_REG_20__SCAN_IN, P3_SUB_598_U108);
  nand ginst24178 (P3_SUB_598_U126, P3_IR_REG_19__SCAN_IN, P3_SUB_598_U44);
  nand ginst24179 (P3_SUB_598_U127, P3_SUB_598_U106, P3_SUB_598_U86);
  nand ginst24180 (P3_SUB_598_U128, P3_IR_REG_18__SCAN_IN, P3_SUB_598_U127);
  nand ginst24181 (P3_SUB_598_U129, P3_IR_REG_16__SCAN_IN, P3_SUB_598_U105);
  and ginst24182 (P3_SUB_598_U13, P3_SUB_598_U128, P3_SUB_598_U44);
  nand ginst24183 (P3_SUB_598_U130, P3_IR_REG_15__SCAN_IN, P3_SUB_598_U47);
  nand ginst24184 (P3_SUB_598_U131, P3_SUB_598_U103, P3_SUB_598_U88);
  nand ginst24185 (P3_SUB_598_U132, P3_IR_REG_14__SCAN_IN, P3_SUB_598_U131);
  nand ginst24186 (P3_SUB_598_U133, P3_IR_REG_12__SCAN_IN, P3_SUB_598_U102);
  nand ginst24187 (P3_SUB_598_U134, P3_IR_REG_11__SCAN_IN, P3_SUB_598_U49);
  nand ginst24188 (P3_SUB_598_U135, P3_SUB_598_U71, P3_SUB_598_U94);
  nand ginst24189 (P3_SUB_598_U136, P3_IR_REG_10__SCAN_IN, P3_SUB_598_U135);
  nand ginst24190 (P3_SUB_598_U137, P3_SUB_598_U115, P3_SUB_598_U76);
  nand ginst24191 (P3_SUB_598_U138, P3_IR_REG_27__SCAN_IN, P3_IR_REG_28__SCAN_IN);
  nand ginst24192 (P3_SUB_598_U139, P3_IR_REG_28__SCAN_IN, P3_SUB_598_U78);
  and ginst24193 (P3_SUB_598_U14, P3_SUB_598_U108, P3_SUB_598_U126);
  not ginst24194 (P3_SUB_598_U140, P3_SUB_598_U28);
  nand ginst24195 (P3_SUB_598_U141, P3_IR_REG_9__SCAN_IN, P3_SUB_598_U29);
  nand ginst24196 (P3_SUB_598_U142, P3_SUB_598_U71, P3_SUB_598_U94);
  nand ginst24197 (P3_SUB_598_U143, P3_IR_REG_5__SCAN_IN, P3_SUB_598_U30);
  nand ginst24198 (P3_SUB_598_U144, P3_SUB_598_U73, P3_SUB_598_U91);
  nand ginst24199 (P3_SUB_598_U145, P3_SUB_598_U137, P3_SUB_598_U75);
  nand ginst24200 (P3_SUB_598_U146, P3_IR_REG_31__SCAN_IN, P3_SUB_598_U115, P3_SUB_598_U76);
  nand ginst24201 (P3_SUB_598_U147, P3_IR_REG_30__SCAN_IN, P3_SUB_598_U37);
  nand ginst24202 (P3_SUB_598_U148, P3_SUB_598_U115, P3_SUB_598_U76);
  nand ginst24203 (P3_SUB_598_U149, P3_IR_REG_27__SCAN_IN, P3_SUB_598_U78);
  and ginst24204 (P3_SUB_598_U15, P3_SUB_598_U125, P3_SUB_598_U40);
  nand ginst24205 (P3_SUB_598_U150, P3_SUB_598_U113, P3_SUB_598_U39);
  nand ginst24206 (P3_SUB_598_U151, P3_IR_REG_25__SCAN_IN, P3_SUB_598_U35);
  nand ginst24207 (P3_SUB_598_U152, P3_SUB_598_U112, P3_SUB_598_U80);
  nand ginst24208 (P3_SUB_598_U153, P3_IR_REG_21__SCAN_IN, P3_SUB_598_U40);
  nand ginst24209 (P3_SUB_598_U154, P3_SUB_598_U109, P3_SUB_598_U82);
  nand ginst24210 (P3_SUB_598_U155, P3_IR_REG_1__SCAN_IN, P3_SUB_598_U85);
  nand ginst24211 (P3_SUB_598_U156, P3_IR_REG_0__SCAN_IN, P3_SUB_598_U84);
  nand ginst24212 (P3_SUB_598_U157, P3_IR_REG_17__SCAN_IN, P3_SUB_598_U34);
  nand ginst24213 (P3_SUB_598_U158, P3_SUB_598_U106, P3_SUB_598_U86);
  nand ginst24214 (P3_SUB_598_U159, P3_IR_REG_13__SCAN_IN, P3_SUB_598_U46);
  and ginst24215 (P3_SUB_598_U16, P3_SUB_598_U124, P3_SUB_598_U41);
  nand ginst24216 (P3_SUB_598_U160, P3_SUB_598_U103, P3_SUB_598_U88);
  and ginst24217 (P3_SUB_598_U17, P3_SUB_598_U111, P3_SUB_598_U122);
  and ginst24218 (P3_SUB_598_U18, P3_SUB_598_U121, P3_SUB_598_U35);
  and ginst24219 (P3_SUB_598_U19, P3_SUB_598_U120, P3_SUB_598_U78);
  and ginst24220 (P3_SUB_598_U20, P3_SUB_598_U139, P3_SUB_598_U65);
  and ginst24221 (P3_SUB_598_U21, P3_SUB_598_U118, P3_SUB_598_U37);
  and ginst24222 (P3_SUB_598_U22, P3_SUB_598_U117, P3_SUB_598_U28);
  and ginst24223 (P3_SUB_598_U23, P3_SUB_598_U100, P3_SUB_598_U90);
  and ginst24224 (P3_SUB_598_U24, P3_SUB_598_U30, P3_SUB_598_U99);
  and ginst24225 (P3_SUB_598_U25, P3_SUB_598_U31, P3_SUB_598_U98);
  and ginst24226 (P3_SUB_598_U26, P3_SUB_598_U93, P3_SUB_598_U96);
  and ginst24227 (P3_SUB_598_U27, P3_SUB_598_U29, P3_SUB_598_U95);
  or ginst24228 (P3_SUB_598_U28, P3_IR_REG_0__SCAN_IN, P3_IR_REG_1__SCAN_IN, P3_IR_REG_2__SCAN_IN);
  nand ginst24229 (P3_SUB_598_U29, P3_SUB_598_U140, P3_SUB_598_U53, P3_SUB_598_U54);
  nand ginst24230 (P3_SUB_598_U30, P3_SUB_598_U140, P3_SUB_598_U55);
  nand ginst24231 (P3_SUB_598_U31, P3_SUB_598_U56, P3_SUB_598_U91);
  not ginst24232 (P3_SUB_598_U32, P3_IR_REG_7__SCAN_IN);
  not ginst24233 (P3_SUB_598_U33, P3_IR_REG_3__SCAN_IN);
  nand ginst24234 (P3_SUB_598_U34, P3_SUB_598_U57, P3_SUB_598_U58, P3_SUB_598_U59, P3_SUB_598_U60);
  nand ginst24235 (P3_SUB_598_U35, P3_SUB_598_U106, P3_SUB_598_U62);
  nand ginst24236 (P3_SUB_598_U36, P3_SUB_598_U112, P3_SUB_598_U63);
  nand ginst24237 (P3_SUB_598_U37, P3_SUB_598_U114, P3_SUB_598_U38);
  not ginst24238 (P3_SUB_598_U38, P3_IR_REG_29__SCAN_IN);
  not ginst24239 (P3_SUB_598_U39, P3_IR_REG_27__SCAN_IN);
  nand ginst24240 (P3_SUB_598_U40, P3_SUB_598_U106, P3_SUB_598_U6);
  nand ginst24241 (P3_SUB_598_U41, P3_SUB_598_U109, P3_SUB_598_U66);
  not ginst24242 (P3_SUB_598_U42, P3_IR_REG_24__SCAN_IN);
  not ginst24243 (P3_SUB_598_U43, P3_IR_REG_23__SCAN_IN);
  nand ginst24244 (P3_SUB_598_U44, P3_SUB_598_U106, P3_SUB_598_U67);
  not ginst24245 (P3_SUB_598_U45, P3_IR_REG_19__SCAN_IN);
  nand ginst24246 (P3_SUB_598_U46, P3_SUB_598_U68, P3_SUB_598_U94);
  nand ginst24247 (P3_SUB_598_U47, P3_SUB_598_U103, P3_SUB_598_U69);
  not ginst24248 (P3_SUB_598_U48, P3_IR_REG_15__SCAN_IN);
  nand ginst24249 (P3_SUB_598_U49, P3_SUB_598_U70, P3_SUB_598_U94);
  not ginst24250 (P3_SUB_598_U50, P3_IR_REG_11__SCAN_IN);
  nand ginst24251 (P3_SUB_598_U51, P3_SUB_598_U155, P3_SUB_598_U156);
  nand ginst24252 (P3_SUB_598_U52, P3_SUB_598_U145, P3_SUB_598_U146);
  nor ginst24253 (P3_SUB_598_U53, P3_IR_REG_3__SCAN_IN, P3_IR_REG_4__SCAN_IN, P3_IR_REG_5__SCAN_IN, P3_IR_REG_6__SCAN_IN);
  nor ginst24254 (P3_SUB_598_U54, P3_IR_REG_7__SCAN_IN, P3_IR_REG_8__SCAN_IN);
  nor ginst24255 (P3_SUB_598_U55, P3_IR_REG_3__SCAN_IN, P3_IR_REG_4__SCAN_IN);
  nor ginst24256 (P3_SUB_598_U56, P3_IR_REG_5__SCAN_IN, P3_IR_REG_6__SCAN_IN);
  nor ginst24257 (P3_SUB_598_U57, P3_IR_REG_10__SCAN_IN, P3_IR_REG_11__SCAN_IN, P3_IR_REG_12__SCAN_IN, P3_IR_REG_13__SCAN_IN, P3_IR_REG_14__SCAN_IN);
  nor ginst24258 (P3_SUB_598_U58, P3_IR_REG_0__SCAN_IN, P3_IR_REG_1__SCAN_IN, P3_IR_REG_15__SCAN_IN, P3_IR_REG_16__SCAN_IN);
  nor ginst24259 (P3_SUB_598_U59, P3_IR_REG_2__SCAN_IN, P3_IR_REG_3__SCAN_IN, P3_IR_REG_4__SCAN_IN, P3_IR_REG_5__SCAN_IN);
  nor ginst24260 (P3_SUB_598_U6, P3_IR_REG_17__SCAN_IN, P3_IR_REG_18__SCAN_IN, P3_IR_REG_19__SCAN_IN, P3_IR_REG_20__SCAN_IN);
  nor ginst24261 (P3_SUB_598_U60, P3_IR_REG_6__SCAN_IN, P3_IR_REG_7__SCAN_IN, P3_IR_REG_8__SCAN_IN, P3_IR_REG_9__SCAN_IN);
  nor ginst24262 (P3_SUB_598_U61, P3_IR_REG_21__SCAN_IN, P3_IR_REG_22__SCAN_IN, P3_IR_REG_23__SCAN_IN);
  and ginst24263 (P3_SUB_598_U62, P3_SUB_598_U42, P3_SUB_598_U6, P3_SUB_598_U61);
  nor ginst24264 (P3_SUB_598_U63, P3_IR_REG_25__SCAN_IN, P3_IR_REG_26__SCAN_IN, P3_IR_REG_27__SCAN_IN, P3_IR_REG_28__SCAN_IN);
  nor ginst24265 (P3_SUB_598_U64, P3_IR_REG_25__SCAN_IN, P3_IR_REG_26__SCAN_IN);
  and ginst24266 (P3_SUB_598_U65, P3_SUB_598_U138, P3_SUB_598_U36);
  nor ginst24267 (P3_SUB_598_U66, P3_IR_REG_21__SCAN_IN, P3_IR_REG_22__SCAN_IN);
  nor ginst24268 (P3_SUB_598_U67, P3_IR_REG_17__SCAN_IN, P3_IR_REG_18__SCAN_IN);
  nor ginst24269 (P3_SUB_598_U68, P3_IR_REG_9__SCAN_IN, P3_IR_REG_10__SCAN_IN, P3_IR_REG_11__SCAN_IN, P3_IR_REG_12__SCAN_IN);
  nor ginst24270 (P3_SUB_598_U69, P3_IR_REG_13__SCAN_IN, P3_IR_REG_14__SCAN_IN);
  and ginst24271 (P3_SUB_598_U7, P3_SUB_598_U136, P3_SUB_598_U49);
  nor ginst24272 (P3_SUB_598_U70, P3_IR_REG_9__SCAN_IN, P3_IR_REG_10__SCAN_IN);
  not ginst24273 (P3_SUB_598_U71, P3_IR_REG_9__SCAN_IN);
  and ginst24274 (P3_SUB_598_U72, P3_SUB_598_U141, P3_SUB_598_U142);
  not ginst24275 (P3_SUB_598_U73, P3_IR_REG_5__SCAN_IN);
  and ginst24276 (P3_SUB_598_U74, P3_SUB_598_U143, P3_SUB_598_U144);
  not ginst24277 (P3_SUB_598_U75, P3_IR_REG_31__SCAN_IN);
  not ginst24278 (P3_SUB_598_U76, P3_IR_REG_30__SCAN_IN);
  and ginst24279 (P3_SUB_598_U77, P3_SUB_598_U147, P3_SUB_598_U148);
  nand ginst24280 (P3_SUB_598_U78, P3_SUB_598_U112, P3_SUB_598_U64);
  and ginst24281 (P3_SUB_598_U79, P3_SUB_598_U149, P3_SUB_598_U150);
  and ginst24282 (P3_SUB_598_U8, P3_SUB_598_U102, P3_SUB_598_U134);
  not ginst24283 (P3_SUB_598_U80, P3_IR_REG_25__SCAN_IN);
  and ginst24284 (P3_SUB_598_U81, P3_SUB_598_U151, P3_SUB_598_U152);
  not ginst24285 (P3_SUB_598_U82, P3_IR_REG_21__SCAN_IN);
  and ginst24286 (P3_SUB_598_U83, P3_SUB_598_U153, P3_SUB_598_U154);
  not ginst24287 (P3_SUB_598_U84, P3_IR_REG_1__SCAN_IN);
  not ginst24288 (P3_SUB_598_U85, P3_IR_REG_0__SCAN_IN);
  not ginst24289 (P3_SUB_598_U86, P3_IR_REG_17__SCAN_IN);
  and ginst24290 (P3_SUB_598_U87, P3_SUB_598_U157, P3_SUB_598_U158);
  not ginst24291 (P3_SUB_598_U88, P3_IR_REG_13__SCAN_IN);
  and ginst24292 (P3_SUB_598_U89, P3_SUB_598_U159, P3_SUB_598_U160);
  and ginst24293 (P3_SUB_598_U9, P3_SUB_598_U133, P3_SUB_598_U46);
  nand ginst24294 (P3_SUB_598_U90, P3_SUB_598_U140, P3_SUB_598_U33);
  not ginst24295 (P3_SUB_598_U91, P3_SUB_598_U30);
  not ginst24296 (P3_SUB_598_U92, P3_SUB_598_U31);
  nand ginst24297 (P3_SUB_598_U93, P3_SUB_598_U32, P3_SUB_598_U92);
  not ginst24298 (P3_SUB_598_U94, P3_SUB_598_U29);
  nand ginst24299 (P3_SUB_598_U95, P3_IR_REG_8__SCAN_IN, P3_SUB_598_U93);
  nand ginst24300 (P3_SUB_598_U96, P3_IR_REG_7__SCAN_IN, P3_SUB_598_U31);
  nand ginst24301 (P3_SUB_598_U97, P3_SUB_598_U73, P3_SUB_598_U91);
  nand ginst24302 (P3_SUB_598_U98, P3_IR_REG_6__SCAN_IN, P3_SUB_598_U97);
  nand ginst24303 (P3_SUB_598_U99, P3_IR_REG_4__SCAN_IN, P3_SUB_598_U90);
  nand ginst24304 (P3_SUB_609_U10, P3_SUB_609_U87, P3_SUB_609_U97);
  nand ginst24305 (P3_SUB_609_U100, P3_REG3_REG_21__SCAN_IN, P3_SUB_609_U83);
  nand ginst24306 (P3_SUB_609_U101, P3_REG3_REG_20__SCAN_IN, P3_SUB_609_U38);
  nand ginst24307 (P3_SUB_609_U102, P3_REG3_REG_19__SCAN_IN, P3_SUB_609_U81);
  nand ginst24308 (P3_SUB_609_U103, P3_REG3_REG_18__SCAN_IN, P3_SUB_609_U37);
  nand ginst24309 (P3_SUB_609_U104, P3_REG3_REG_17__SCAN_IN, P3_SUB_609_U79);
  nand ginst24310 (P3_SUB_609_U105, P3_REG3_REG_16__SCAN_IN, P3_SUB_609_U36);
  nand ginst24311 (P3_SUB_609_U106, P3_REG3_REG_15__SCAN_IN, P3_SUB_609_U77);
  nand ginst24312 (P3_SUB_609_U107, P3_REG3_REG_14__SCAN_IN, P3_SUB_609_U35);
  nand ginst24313 (P3_SUB_609_U108, P3_REG3_REG_13__SCAN_IN, P3_SUB_609_U75);
  nand ginst24314 (P3_SUB_609_U109, P3_REG3_REG_12__SCAN_IN, P3_SUB_609_U34);
  nand ginst24315 (P3_SUB_609_U11, P3_SUB_609_U103, P3_SUB_609_U81);
  nand ginst24316 (P3_SUB_609_U110, P3_REG3_REG_11__SCAN_IN, P3_SUB_609_U73);
  nand ginst24317 (P3_SUB_609_U111, P3_REG3_REG_10__SCAN_IN, P3_SUB_609_U33);
  or ginst24318 (P3_SUB_609_U112, P3_REG3_REG_3__SCAN_IN, P3_REG3_REG_5__SCAN_IN, P3_REG3_REG_4__SCAN_IN);
  nand ginst24319 (P3_SUB_609_U113, P3_REG3_REG_6__SCAN_IN, P3_SUB_609_U112);
  nand ginst24320 (P3_SUB_609_U114, P3_REG3_REG_5__SCAN_IN, P3_SUB_609_U64);
  or ginst24321 (P3_SUB_609_U115, P3_REG3_REG_3__SCAN_IN, P3_REG3_REG_5__SCAN_IN, P3_REG3_REG_4__SCAN_IN);
  nand ginst24322 (P3_SUB_609_U12, P3_SUB_609_U67, P3_SUB_609_U70);
  nand ginst24323 (P3_SUB_609_U13, P3_SUB_609_U111, P3_SUB_609_U73);
  nand ginst24324 (P3_SUB_609_U14, P3_SUB_609_U33, P3_SUB_609_U69);
  nand ginst24325 (P3_SUB_609_U15, P3_SUB_609_U102, P3_SUB_609_U38);
  nand ginst24326 (P3_SUB_609_U16, P3_SUB_609_U41, P3_SUB_609_U96);
  nand ginst24327 (P3_SUB_609_U17, P3_SUB_609_U85, P3_SUB_609_U99);
  nand ginst24328 (P3_SUB_609_U18, P3_SUB_609_U31, P3_SUB_609_U71);
  nand ginst24329 (P3_SUB_609_U19, P3_SUB_609_U104, P3_SUB_609_U37);
  nand ginst24330 (P3_SUB_609_U20, P3_SUB_609_U101, P3_SUB_609_U83);
  nand ginst24331 (P3_SUB_609_U21, P3_SUB_609_U106, P3_SUB_609_U36);
  nand ginst24332 (P3_SUB_609_U22, P3_SUB_609_U42, P3_SUB_609_U94);
  nand ginst24333 (P3_SUB_609_U23, P3_SUB_609_U109, P3_SUB_609_U75);
  nand ginst24334 (P3_SUB_609_U24, P3_SUB_609_U108, P3_SUB_609_U35);
  not ginst24335 (P3_SUB_609_U25, P3_REG3_REG_3__SCAN_IN);
  nand ginst24336 (P3_SUB_609_U26, P3_SUB_609_U89, P3_SUB_609_U95);
  nand ginst24337 (P3_SUB_609_U27, P3_SUB_609_U100, P3_SUB_609_U39);
  nand ginst24338 (P3_SUB_609_U28, P3_SUB_609_U91, P3_SUB_609_U93);
  nand ginst24339 (P3_SUB_609_U29, P3_SUB_609_U64, P3_SUB_609_U72);
  nand ginst24340 (P3_SUB_609_U30, P3_SUB_609_U107, P3_SUB_609_U77);
  or ginst24341 (P3_SUB_609_U31, P3_REG3_REG_7__SCAN_IN, P3_REG3_REG_3__SCAN_IN, P3_REG3_REG_5__SCAN_IN, P3_REG3_REG_4__SCAN_IN, P3_REG3_REG_6__SCAN_IN);
  not ginst24342 (P3_SUB_609_U32, P3_REG3_REG_8__SCAN_IN);
  nand ginst24343 (P3_SUB_609_U33, P3_SUB_609_U54, P3_SUB_609_U66);
  nand ginst24344 (P3_SUB_609_U34, P3_SUB_609_U55, P3_SUB_609_U68);
  nand ginst24345 (P3_SUB_609_U35, P3_SUB_609_U56, P3_SUB_609_U74);
  nand ginst24346 (P3_SUB_609_U36, P3_SUB_609_U57, P3_SUB_609_U76);
  nand ginst24347 (P3_SUB_609_U37, P3_SUB_609_U58, P3_SUB_609_U78);
  nand ginst24348 (P3_SUB_609_U38, P3_SUB_609_U59, P3_SUB_609_U80);
  nand ginst24349 (P3_SUB_609_U39, P3_SUB_609_U60, P3_SUB_609_U82);
  nand ginst24350 (P3_SUB_609_U40, P3_SUB_609_U61, P3_SUB_609_U84);
  nand ginst24351 (P3_SUB_609_U41, P3_SUB_609_U62, P3_SUB_609_U86);
  nand ginst24352 (P3_SUB_609_U42, P3_SUB_609_U63, P3_SUB_609_U88);
  not ginst24353 (P3_SUB_609_U43, P3_REG3_REG_28__SCAN_IN);
  not ginst24354 (P3_SUB_609_U44, P3_REG3_REG_26__SCAN_IN);
  not ginst24355 (P3_SUB_609_U45, P3_REG3_REG_24__SCAN_IN);
  not ginst24356 (P3_SUB_609_U46, P3_REG3_REG_22__SCAN_IN);
  not ginst24357 (P3_SUB_609_U47, P3_REG3_REG_20__SCAN_IN);
  not ginst24358 (P3_SUB_609_U48, P3_REG3_REG_18__SCAN_IN);
  not ginst24359 (P3_SUB_609_U49, P3_REG3_REG_16__SCAN_IN);
  not ginst24360 (P3_SUB_609_U50, P3_REG3_REG_14__SCAN_IN);
  not ginst24361 (P3_SUB_609_U51, P3_REG3_REG_12__SCAN_IN);
  not ginst24362 (P3_SUB_609_U52, P3_REG3_REG_10__SCAN_IN);
  nand ginst24363 (P3_SUB_609_U53, P3_SUB_609_U114, P3_SUB_609_U115);
  nor ginst24364 (P3_SUB_609_U54, P3_REG3_REG_8__SCAN_IN, P3_REG3_REG_9__SCAN_IN);
  nor ginst24365 (P3_SUB_609_U55, P3_REG3_REG_10__SCAN_IN, P3_REG3_REG_11__SCAN_IN);
  nor ginst24366 (P3_SUB_609_U56, P3_REG3_REG_12__SCAN_IN, P3_REG3_REG_13__SCAN_IN);
  nor ginst24367 (P3_SUB_609_U57, P3_REG3_REG_14__SCAN_IN, P3_REG3_REG_15__SCAN_IN);
  nor ginst24368 (P3_SUB_609_U58, P3_REG3_REG_16__SCAN_IN, P3_REG3_REG_17__SCAN_IN);
  nor ginst24369 (P3_SUB_609_U59, P3_REG3_REG_19__SCAN_IN, P3_REG3_REG_18__SCAN_IN);
  nand ginst24370 (P3_SUB_609_U6, P3_SUB_609_U40, P3_SUB_609_U98);
  nor ginst24371 (P3_SUB_609_U60, P3_REG3_REG_21__SCAN_IN, P3_REG3_REG_20__SCAN_IN);
  nor ginst24372 (P3_SUB_609_U61, P3_REG3_REG_23__SCAN_IN, P3_REG3_REG_22__SCAN_IN);
  nor ginst24373 (P3_SUB_609_U62, P3_REG3_REG_25__SCAN_IN, P3_REG3_REG_24__SCAN_IN);
  nor ginst24374 (P3_SUB_609_U63, P3_REG3_REG_27__SCAN_IN, P3_REG3_REG_26__SCAN_IN);
  or ginst24375 (P3_SUB_609_U64, P3_REG3_REG_3__SCAN_IN, P3_REG3_REG_4__SCAN_IN);
  or ginst24376 (P3_SUB_609_U65, P3_REG3_REG_3__SCAN_IN, P3_REG3_REG_5__SCAN_IN, P3_REG3_REG_4__SCAN_IN, P3_REG3_REG_6__SCAN_IN);
  not ginst24377 (P3_SUB_609_U66, P3_SUB_609_U31);
  nand ginst24378 (P3_SUB_609_U67, P3_SUB_609_U32, P3_SUB_609_U66);
  not ginst24379 (P3_SUB_609_U68, P3_SUB_609_U33);
  nand ginst24380 (P3_SUB_609_U69, P3_REG3_REG_9__SCAN_IN, P3_SUB_609_U67);
  nand ginst24381 (P3_SUB_609_U7, P3_SUB_609_U105, P3_SUB_609_U79);
  nand ginst24382 (P3_SUB_609_U70, P3_REG3_REG_8__SCAN_IN, P3_SUB_609_U31);
  nand ginst24383 (P3_SUB_609_U71, P3_REG3_REG_7__SCAN_IN, P3_SUB_609_U65);
  nand ginst24384 (P3_SUB_609_U72, P3_REG3_REG_3__SCAN_IN, P3_REG3_REG_4__SCAN_IN);
  nand ginst24385 (P3_SUB_609_U73, P3_SUB_609_U52, P3_SUB_609_U68);
  not ginst24386 (P3_SUB_609_U74, P3_SUB_609_U34);
  nand ginst24387 (P3_SUB_609_U75, P3_SUB_609_U51, P3_SUB_609_U74);
  not ginst24388 (P3_SUB_609_U76, P3_SUB_609_U35);
  nand ginst24389 (P3_SUB_609_U77, P3_SUB_609_U50, P3_SUB_609_U76);
  not ginst24390 (P3_SUB_609_U78, P3_SUB_609_U36);
  nand ginst24391 (P3_SUB_609_U79, P3_SUB_609_U49, P3_SUB_609_U78);
  nand ginst24392 (P3_SUB_609_U8, P3_SUB_609_U113, P3_SUB_609_U65);
  not ginst24393 (P3_SUB_609_U80, P3_SUB_609_U37);
  nand ginst24394 (P3_SUB_609_U81, P3_SUB_609_U48, P3_SUB_609_U80);
  not ginst24395 (P3_SUB_609_U82, P3_SUB_609_U38);
  nand ginst24396 (P3_SUB_609_U83, P3_SUB_609_U47, P3_SUB_609_U82);
  not ginst24397 (P3_SUB_609_U84, P3_SUB_609_U39);
  nand ginst24398 (P3_SUB_609_U85, P3_SUB_609_U46, P3_SUB_609_U84);
  not ginst24399 (P3_SUB_609_U86, P3_SUB_609_U40);
  nand ginst24400 (P3_SUB_609_U87, P3_SUB_609_U45, P3_SUB_609_U86);
  not ginst24401 (P3_SUB_609_U88, P3_SUB_609_U41);
  nand ginst24402 (P3_SUB_609_U89, P3_SUB_609_U44, P3_SUB_609_U88);
  nand ginst24403 (P3_SUB_609_U9, P3_SUB_609_U110, P3_SUB_609_U34);
  not ginst24404 (P3_SUB_609_U90, P3_SUB_609_U42);
  nand ginst24405 (P3_SUB_609_U91, P3_SUB_609_U43, P3_SUB_609_U90);
  not ginst24406 (P3_SUB_609_U92, P3_SUB_609_U91);
  nand ginst24407 (P3_SUB_609_U93, P3_REG3_REG_28__SCAN_IN, P3_SUB_609_U42);
  nand ginst24408 (P3_SUB_609_U94, P3_REG3_REG_27__SCAN_IN, P3_SUB_609_U89);
  nand ginst24409 (P3_SUB_609_U95, P3_REG3_REG_26__SCAN_IN, P3_SUB_609_U41);
  nand ginst24410 (P3_SUB_609_U96, P3_REG3_REG_25__SCAN_IN, P3_SUB_609_U87);
  nand ginst24411 (P3_SUB_609_U97, P3_REG3_REG_24__SCAN_IN, P3_SUB_609_U40);
  nand ginst24412 (P3_SUB_609_U98, P3_REG3_REG_23__SCAN_IN, P3_SUB_609_U85);
  nand ginst24413 (P3_SUB_609_U99, P3_REG3_REG_22__SCAN_IN, P3_SUB_609_U39);
  and ginst24414 (P3_U3013, P3_U3380, P3_U5450);
  and ginst24415 (P3_U3014, P3_U3379, P3_U3380);
  and ginst24416 (P3_U3015, P3_U3379, P3_U5453);
  and ginst24417 (P3_U3016, P3_U5450, P3_U5453);
  and ginst24418 (P3_U3017, P3_U3874, P3_U5447);
  and ginst24419 (P3_U3018, P3_U3582, P3_U3587);
  and ginst24420 (P3_U3019, P3_U3381, P3_U3382);
  and ginst24421 (P3_U3020, P3_U3381, P3_U5462);
  and ginst24422 (P3_U3021, P3_U3382, P3_U5459);
  and ginst24423 (P3_U3022, P3_U5459, P3_U5462);
  and ginst24424 (P3_U3023, P3_STATE_REG_SCAN_IN, P3_U3046);
  and ginst24425 (P3_U3024, P3_U3366, P3_U3696);
  and ginst24426 (P3_U3025, P3_U3911, P3_U4073);
  and ginst24427 (P3_U3026, P3_U3015, P3_U5447);
  and ginst24428 (P3_U3027, P3_STATE_REG_SCAN_IN, P3_U3297);
  and ginst24429 (P3_U3028, P3_U3886, P3_U3912);
  and ginst24430 (P3_U3029, P3_U3365, P3_U3912);
  and ginst24431 (P3_U3030, P3_U3693, P3_U3912);
  and ginst24432 (P3_U3031, P3_U3023, P3_U3890);
  and ginst24433 (P3_U3032, P3_U3895, P3_U4073);
  and ginst24434 (P3_U3033, P3_U3911, P3_U4089);
  and ginst24435 (P3_U3034, P3_U3025, P3_U3912);
  and ginst24436 (P3_U3035, P3_U3023, P3_U4989);
  and ginst24437 (P3_U3036, P3_U3895, P3_U4089);
  and ginst24438 (P3_U3037, P3_U4754, P3_U5468);
  and ginst24439 (P3_U3038, P3_U3024, P3_U5468);
  and ginst24440 (P3_U3039, P3_U4754, P3_U5465);
  and ginst24441 (P3_U3040, P3_U3892, P3_U4754);
  and ginst24442 (P3_U3041, P3_U3024, P3_U3892);
  and ginst24443 (P3_U3042, P3_U3023, P3_U3366);
  and ginst24444 (P3_U3043, P3_U3023, P3_U3365);
  and ginst24445 (P3_U3044, P3_STATE_REG_SCAN_IN, P3_U5004);
  and ginst24446 (P3_U3045, P3_U3023, P3_U5006);
  and ginst24447 (P3_U3046, P3_U3362, P3_U5440);
  and ginst24448 (P3_U3047, P3_U3018, P3_U3692);
  and ginst24449 (P3_U3048, P3_U3018, P3_U3691);
  and ginst24450 (P3_U3049, P3_U4748, P3_U4749);
  and ginst24451 (P3_U3050, P3_STATE_REG_SCAN_IN, P3_U4759);
  and ginst24452 (P3_U3051, P3_U3897, P3_U4761);
  nand ginst24453 (P3_U3052, P3_U4535, P3_U4536, P3_U4537, P3_U4538);
  nand ginst24454 (P3_U3053, P3_U4553, P3_U4554, P3_U4555, P3_U4556);
  nand ginst24455 (P3_U3054, P3_U4571, P3_U4572, P3_U4573, P3_U4574);
  nand ginst24456 (P3_U3055, P3_U4609, P3_U4610, P3_U4611, P3_U4612);
  nand ginst24457 (P3_U3056, P3_U4517, P3_U4518, P3_U4519, P3_U4520);
  nand ginst24458 (P3_U3057, P3_U4499, P3_U4500, P3_U4501, P3_U4502);
  nand ginst24459 (P3_U3058, P3_U4589, P3_U4590, P3_U4591, P3_U4592);
  nand ginst24460 (P3_U3059, P3_U4121, P3_U4122, P3_U4123, P3_U4124);
  nand ginst24461 (P3_U3060, P3_U4445, P3_U4446, P3_U4447, P3_U4448);
  nand ginst24462 (P3_U3061, P3_U4229, P3_U4230, P3_U4231, P3_U4232);
  nand ginst24463 (P3_U3062, P3_U4247, P3_U4248, P3_U4249, P3_U4250);
  nand ginst24464 (P3_U3063, P3_U4103, P3_U4104, P3_U4105, P3_U4106);
  nand ginst24465 (P3_U3064, P3_U4481, P3_U4482, P3_U4483, P3_U4484);
  nand ginst24466 (P3_U3065, P3_U4463, P3_U4464, P3_U4465, P3_U4466);
  nand ginst24467 (P3_U3066, P3_U4139, P3_U4140, P3_U4141, P3_U4142);
  nand ginst24468 (P3_U3067, P3_U4078, P3_U4079, P3_U4080, P3_U4081);
  nand ginst24469 (P3_U3068, P3_U4355, P3_U4356, P3_U4357, P3_U4358);
  nand ginst24470 (P3_U3069, P3_U4175, P3_U4176, P3_U4177, P3_U4178);
  nand ginst24471 (P3_U3070, P3_U4157, P3_U4158, P3_U4159, P3_U4160);
  nand ginst24472 (P3_U3071, P3_U4265, P3_U4266, P3_U4267, P3_U4268);
  nand ginst24473 (P3_U3072, P3_U4337, P3_U4338, P3_U4339, P3_U4340);
  nand ginst24474 (P3_U3073, P3_U4319, P3_U4320, P3_U4321, P3_U4322);
  nand ginst24475 (P3_U3074, P3_U4427, P3_U4428, P3_U4429, P3_U4430);
  nand ginst24476 (P3_U3075, P3_U4409, P3_U4410, P3_U4411, P3_U4412);
  nand ginst24477 (P3_U3076, P3_U4083, P3_U4084, P3_U4085, P3_U4086);
  nand ginst24478 (P3_U3077, P3_U4059, P3_U4060, P3_U4061, P3_U4062);
  nand ginst24479 (P3_U3078, P3_U4301, P3_U4302, P3_U4303, P3_U4304);
  nand ginst24480 (P3_U3079, P3_U4283, P3_U4284, P3_U4285, P3_U4286);
  nand ginst24481 (P3_U3080, P3_U4391, P3_U4392, P3_U4393, P3_U4394);
  nand ginst24482 (P3_U3081, P3_U4373, P3_U4374, P3_U4375, P3_U4376);
  nand ginst24483 (P3_U3082, P3_U4211, P3_U4212, P3_U4213, P3_U4214);
  nand ginst24484 (P3_U3083, P3_U4193, P3_U4194, P3_U4195, P3_U4196);
  nand ginst24485 (P3_U3084, P3_U5340, P3_U5341);
  nand ginst24486 (P3_U3085, P3_U5342, P3_U5343);
  nand ginst24487 (P3_U3086, P3_U5347, P3_U5348, P3_U5349);
  nand ginst24488 (P3_U3087, P3_U5350, P3_U5351, P3_U5352);
  nand ginst24489 (P3_U3088, P3_U5353, P3_U5354, P3_U5355);
  nand ginst24490 (P3_U3089, P3_U5356, P3_U5357, P3_U5358);
  nand ginst24491 (P3_U3090, P3_U5359, P3_U5360, P3_U5361);
  nand ginst24492 (P3_U3091, P3_U5362, P3_U5363, P3_U5364);
  nand ginst24493 (P3_U3092, P3_U5365, P3_U5366, P3_U5367);
  nand ginst24494 (P3_U3093, P3_U5368, P3_U5369, P3_U5370);
  nand ginst24495 (P3_U3094, P3_U5371, P3_U5372, P3_U5373);
  nand ginst24496 (P3_U3095, P3_U5374, P3_U5375, P3_U5376);
  nand ginst24497 (P3_U3096, P3_U5380, P3_U5381, P3_U5382);
  nand ginst24498 (P3_U3097, P3_U5383, P3_U5384, P3_U5385);
  nand ginst24499 (P3_U3098, P3_U5386, P3_U5387, P3_U5388);
  nand ginst24500 (P3_U3099, P3_U5389, P3_U5390, P3_U5391);
  nand ginst24501 (P3_U3100, P3_U5392, P3_U5393, P3_U5394);
  nand ginst24502 (P3_U3101, P3_U5395, P3_U5396, P3_U5397);
  nand ginst24503 (P3_U3102, P3_U5398, P3_U5399, P3_U5400);
  nand ginst24504 (P3_U3103, P3_U5401, P3_U5402, P3_U5403);
  nand ginst24505 (P3_U3104, P3_U5404, P3_U5405, P3_U5406);
  nand ginst24506 (P3_U3105, P3_U5407, P3_U5408, P3_U5409);
  nand ginst24507 (P3_U3106, P3_U5322, P3_U5323, P3_U5324);
  nand ginst24508 (P3_U3107, P3_U5325, P3_U5326, P3_U5327);
  nand ginst24509 (P3_U3108, P3_U5328, P3_U5329, P3_U5330);
  nand ginst24510 (P3_U3109, P3_U5331, P3_U5332, P3_U5333);
  nand ginst24511 (P3_U3110, P3_U5334, P3_U5335, P3_U5336);
  nand ginst24512 (P3_U3111, P3_U5337, P3_U5338, P3_U5339);
  nand ginst24513 (P3_U3112, P3_U5344, P3_U5345, P3_U5346);
  nand ginst24514 (P3_U3113, P3_U5377, P3_U5378, P3_U5379);
  nand ginst24515 (P3_U3114, P3_U5410, P3_U5411, P3_U5412);
  nand ginst24516 (P3_U3115, P3_U5413, P3_U5414);
  nand ginst24517 (P3_U3116, P3_U5270, P3_U5271);
  nand ginst24518 (P3_U3117, P3_U5272, P3_U5273);
  nand ginst24519 (P3_U3118, P3_U3375, P3_U5276, P3_U5277);
  nand ginst24520 (P3_U3119, P3_U3375, P3_U5278, P3_U5279);
  nand ginst24521 (P3_U3120, P3_U3375, P3_U5280, P3_U5281);
  nand ginst24522 (P3_U3121, P3_U3375, P3_U5282, P3_U5283);
  nand ginst24523 (P3_U3122, P3_U3375, P3_U5284, P3_U5285);
  nand ginst24524 (P3_U3123, P3_U3375, P3_U5286, P3_U5287);
  nand ginst24525 (P3_U3124, P3_U3375, P3_U5288, P3_U5289);
  nand ginst24526 (P3_U3125, P3_U3375, P3_U5290, P3_U5291);
  nand ginst24527 (P3_U3126, P3_U3375, P3_U5292, P3_U5293);
  nand ginst24528 (P3_U3127, P3_U3375, P3_U5294, P3_U5295);
  nand ginst24529 (P3_U3128, P3_U3375, P3_U5298, P3_U5299);
  nand ginst24530 (P3_U3129, P3_U3375, P3_U5300, P3_U5301);
  nand ginst24531 (P3_U3130, P3_U3375, P3_U5302, P3_U5303);
  nand ginst24532 (P3_U3131, P3_U3375, P3_U5304, P3_U5305);
  nand ginst24533 (P3_U3132, P3_U3375, P3_U5306, P3_U5307);
  nand ginst24534 (P3_U3133, P3_U3375, P3_U5308, P3_U5309);
  nand ginst24535 (P3_U3134, P3_U3825, P3_U5311);
  nand ginst24536 (P3_U3135, P3_U3826, P3_U5313);
  nand ginst24537 (P3_U3136, P3_U3827, P3_U5315);
  nand ginst24538 (P3_U3137, P3_U3828, P3_U5317);
  nand ginst24539 (P3_U3138, P3_U3817, P3_U5259);
  nand ginst24540 (P3_U3139, P3_U3818, P3_U5261);
  nand ginst24541 (P3_U3140, P3_U3819, P3_U5263);
  nand ginst24542 (P3_U3141, P3_U3820, P3_U5265);
  nand ginst24543 (P3_U3142, P3_U3821, P3_U5267);
  nand ginst24544 (P3_U3143, P3_U3822, P3_U5269);
  nand ginst24545 (P3_U3144, P3_U3823, P3_U5275);
  nand ginst24546 (P3_U3145, P3_U3824, P3_U5297);
  nand ginst24547 (P3_U3146, P3_U3829, P3_U5319);
  nand ginst24548 (P3_U3147, P3_U3830, P3_U5321);
  nand ginst24549 (P3_U3148, P3_U3375, P3_U3385, P3_U5453);
  nand ginst24550 (P3_U3149, P3_U3013, P3_U3813);
  nand ginst24551 (P3_U3150, P3_U3812, P3_U5253);
  not ginst24552 (P3_U3151, P3_STATE_REG_SCAN_IN);
  nand ginst24553 (P3_U3152, P3_U3359, P3_U5943, P3_U5944);
  nand ginst24554 (P3_U3153, P3_U3811, P3_U5248, P3_U5249, P3_U5250);
  nand ginst24555 (P3_U3154, P3_U3810, P3_U5239, P3_U5240, P3_U5241);
  nand ginst24556 (P3_U3155, P3_U3809, P3_U5230, P3_U5231, P3_U5232);
  nand ginst24557 (P3_U3156, P3_U3808, P3_U5221, P3_U5222, P3_U5223);
  nand ginst24558 (P3_U3157, P3_U3807, P3_U5212, P3_U5213, P3_U5214);
  nand ginst24559 (P3_U3158, P3_U3805, P3_U3806, P3_U5204);
  nand ginst24560 (P3_U3159, P3_U3804, P3_U5194, P3_U5195, P3_U5196);
  nand ginst24561 (P3_U3160, P3_U3803, P3_U5185, P3_U5186, P3_U5187);
  nand ginst24562 (P3_U3161, P3_U3802, P3_U5176, P3_U5177, P3_U5178);
  nand ginst24563 (P3_U3162, P3_U3800, P3_U3801, P3_U5168);
  nand ginst24564 (P3_U3163, P3_U3799, P3_U5158, P3_U5159, P3_U5160);
  nand ginst24565 (P3_U3164, P3_U3798, P3_U5149, P3_U5150, P3_U5151);
  nand ginst24566 (P3_U3165, P3_U3797, P3_U5140, P3_U5141, P3_U5142);
  nand ginst24567 (P3_U3166, P3_U3796, P3_U5131, P3_U5132, P3_U5133);
  nand ginst24568 (P3_U3167, P3_U3795, P3_U5122, P3_U5123, P3_U5124);
  nand ginst24569 (P3_U3168, P3_U3794, P3_U5113, P3_U5114, P3_U5115);
  nand ginst24570 (P3_U3169, P3_U3793, P3_U5104, P3_U5105, P3_U5106);
  nand ginst24571 (P3_U3170, P3_U3791, P3_U3792, P3_U5096);
  nand ginst24572 (P3_U3171, P3_U3790, P3_U5086, P3_U5087, P3_U5088);
  nand ginst24573 (P3_U3172, P3_U3789, P3_U5079);
  nand ginst24574 (P3_U3173, P3_U3786, P3_U5070, P3_U5071, P3_U5072);
  nand ginst24575 (P3_U3174, P3_U3785, P3_U5061, P3_U5062, P3_U5063);
  nand ginst24576 (P3_U3175, P3_U3784, P3_U5052, P3_U5053, P3_U5054);
  nand ginst24577 (P3_U3176, P3_U3783, P3_U5043, P3_U5044, P3_U5045);
  nand ginst24578 (P3_U3177, P3_U3781, P3_U3782, P3_U5035);
  nand ginst24579 (P3_U3178, P3_U3780, P3_U5025, P3_U5026, P3_U5027);
  nand ginst24580 (P3_U3179, P3_U3779, P3_U5016, P3_U5017, P3_U5018);
  nand ginst24581 (P3_U3180, P3_U3778, P3_U5007, P3_U5008, P3_U5009);
  nand ginst24582 (P3_U3181, P3_U3777, P3_U4994, P3_U4995, P3_U4996);
  nand ginst24583 (P3_U3182, P3_U3756, P3_U4973);
  nand ginst24584 (P3_U3183, P3_U3753, P3_U4962);
  nand ginst24585 (P3_U3184, P3_U3750, P3_U4951);
  nand ginst24586 (P3_U3185, P3_U3747, P3_U4940, P3_U4941);
  nand ginst24587 (P3_U3186, P3_U3744, P3_U4929, P3_U4930);
  nand ginst24588 (P3_U3187, P3_U3741, P3_U3743, P3_U4916, P3_U4918);
  nand ginst24589 (P3_U3188, P3_U3738, P3_U4905, P3_U4907);
  nand ginst24590 (P3_U3189, P3_U3735, P3_U4896);
  nand ginst24591 (P3_U3190, P3_U3732, P3_U4885);
  nand ginst24592 (P3_U3191, P3_U3729, P3_U4874);
  nand ginst24593 (P3_U3192, P3_U3726, P3_U4863);
  nand ginst24594 (P3_U3193, P3_U3723, P3_U4852);
  nand ginst24595 (P3_U3194, P3_U3720, P3_U4841);
  nand ginst24596 (P3_U3195, P3_U3717, P3_U4830);
  nand ginst24597 (P3_U3196, P3_U3714, P3_U4819);
  nand ginst24598 (P3_U3197, P3_U3711, P3_U4808);
  nand ginst24599 (P3_U3198, P3_U3708, P3_U4797);
  nand ginst24600 (P3_U3199, P3_U3705, P3_U4786);
  nand ginst24601 (P3_U3200, P3_U3702, P3_U4775);
  nand ginst24602 (P3_U3201, P3_U3699, P3_U4764);
  nand ginst24603 (P3_U3202, P3_U3049, P3_U4752, P3_U4753);
  nand ginst24604 (P3_U3203, P3_U3049, P3_U4750, P3_U4751);
  nand ginst24605 (P3_U3204, P3_U3866, P3_U4745, P3_U4746, P3_U4747);
  nand ginst24606 (P3_U3205, P3_U3865, P3_U4741, P3_U4742, P3_U4743, P3_U4744);
  nand ginst24607 (P3_U3206, P3_U3864, P3_U4737, P3_U4738, P3_U4739, P3_U4740);
  nand ginst24608 (P3_U3207, P3_U3863, P3_U4733, P3_U4734, P3_U4735, P3_U4736);
  nand ginst24609 (P3_U3208, P3_U3862, P3_U4729, P3_U4730, P3_U4731, P3_U4732);
  nand ginst24610 (P3_U3209, P3_U3861, P3_U4725, P3_U4726, P3_U4727, P3_U4728);
  nand ginst24611 (P3_U3210, P3_U3860, P3_U4721, P3_U4722, P3_U4723, P3_U4724);
  nand ginst24612 (P3_U3211, P3_U3859, P3_U4717, P3_U4718, P3_U4719, P3_U4720);
  nand ginst24613 (P3_U3212, P3_U3858, P3_U4713, P3_U4714, P3_U4715, P3_U4716);
  nand ginst24614 (P3_U3213, P3_U3857, P3_U4709, P3_U4710, P3_U4711, P3_U4712);
  nand ginst24615 (P3_U3214, P3_U3856, P3_U4705, P3_U4706, P3_U4707, P3_U4708);
  nand ginst24616 (P3_U3215, P3_U3855, P3_U4701, P3_U4702, P3_U4703, P3_U4704);
  nand ginst24617 (P3_U3216, P3_U3854, P3_U4697, P3_U4698, P3_U4699, P3_U4700);
  nand ginst24618 (P3_U3217, P3_U3853, P3_U4693, P3_U4694, P3_U4695, P3_U4696);
  nand ginst24619 (P3_U3218, P3_U3852, P3_U4689, P3_U4690, P3_U4691, P3_U4692);
  nand ginst24620 (P3_U3219, P3_U3851, P3_U4685, P3_U4686, P3_U4687, P3_U4688);
  nand ginst24621 (P3_U3220, P3_U3850, P3_U4681, P3_U4682, P3_U4683, P3_U4684);
  nand ginst24622 (P3_U3221, P3_U3849, P3_U4677, P3_U4678, P3_U4679, P3_U4680);
  nand ginst24623 (P3_U3222, P3_U3848, P3_U4673, P3_U4674, P3_U4675, P3_U4676);
  nand ginst24624 (P3_U3223, P3_U3847, P3_U4669, P3_U4670, P3_U4671, P3_U4672);
  nand ginst24625 (P3_U3224, P3_U3846, P3_U4665, P3_U4666, P3_U4667, P3_U4668);
  nand ginst24626 (P3_U3225, P3_U3845, P3_U4661, P3_U4662, P3_U4663, P3_U4664);
  nand ginst24627 (P3_U3226, P3_U3844, P3_U4657, P3_U4658, P3_U4659, P3_U4660);
  nand ginst24628 (P3_U3227, P3_U3843, P3_U4653, P3_U4654, P3_U4655, P3_U4656);
  nand ginst24629 (P3_U3228, P3_U3842, P3_U4649, P3_U4650, P3_U4651, P3_U4652);
  nand ginst24630 (P3_U3229, P3_U3841, P3_U4645, P3_U4646, P3_U4647, P3_U4648);
  nand ginst24631 (P3_U3230, P3_U3840, P3_U4641, P3_U4642, P3_U4643, P3_U4644);
  nand ginst24632 (P3_U3231, P3_U3839, P3_U4637, P3_U4638, P3_U4639, P3_U4640);
  nand ginst24633 (P3_U3232, P3_U3838, P3_U4633, P3_U4634, P3_U4635, P3_U4636);
  nand ginst24634 (P3_U3233, P3_U3837, P3_U4629, P3_U4630, P3_U4631, P3_U4632);
  and ginst24635 (P3_U3234, P3_D_REG_31__SCAN_IN, P3_U3832);
  and ginst24636 (P3_U3235, P3_D_REG_30__SCAN_IN, P3_U3832);
  and ginst24637 (P3_U3236, P3_D_REG_29__SCAN_IN, P3_U3832);
  and ginst24638 (P3_U3237, P3_D_REG_28__SCAN_IN, P3_U3832);
  and ginst24639 (P3_U3238, P3_D_REG_27__SCAN_IN, P3_U3832);
  and ginst24640 (P3_U3239, P3_D_REG_26__SCAN_IN, P3_U3832);
  and ginst24641 (P3_U3240, P3_D_REG_25__SCAN_IN, P3_U3832);
  and ginst24642 (P3_U3241, P3_D_REG_24__SCAN_IN, P3_U3832);
  and ginst24643 (P3_U3242, P3_D_REG_23__SCAN_IN, P3_U3832);
  and ginst24644 (P3_U3243, P3_D_REG_22__SCAN_IN, P3_U3832);
  and ginst24645 (P3_U3244, P3_D_REG_21__SCAN_IN, P3_U3832);
  and ginst24646 (P3_U3245, P3_D_REG_20__SCAN_IN, P3_U3832);
  and ginst24647 (P3_U3246, P3_D_REG_19__SCAN_IN, P3_U3832);
  and ginst24648 (P3_U3247, P3_D_REG_18__SCAN_IN, P3_U3832);
  and ginst24649 (P3_U3248, P3_D_REG_17__SCAN_IN, P3_U3832);
  and ginst24650 (P3_U3249, P3_D_REG_16__SCAN_IN, P3_U3832);
  and ginst24651 (P3_U3250, P3_D_REG_15__SCAN_IN, P3_U3832);
  and ginst24652 (P3_U3251, P3_D_REG_14__SCAN_IN, P3_U3832);
  and ginst24653 (P3_U3252, P3_D_REG_13__SCAN_IN, P3_U3832);
  and ginst24654 (P3_U3253, P3_D_REG_12__SCAN_IN, P3_U3832);
  and ginst24655 (P3_U3254, P3_D_REG_11__SCAN_IN, P3_U3832);
  and ginst24656 (P3_U3255, P3_D_REG_10__SCAN_IN, P3_U3832);
  and ginst24657 (P3_U3256, P3_D_REG_9__SCAN_IN, P3_U3832);
  and ginst24658 (P3_U3257, P3_D_REG_8__SCAN_IN, P3_U3832);
  and ginst24659 (P3_U3258, P3_D_REG_7__SCAN_IN, P3_U3832);
  and ginst24660 (P3_U3259, P3_D_REG_6__SCAN_IN, P3_U3832);
  and ginst24661 (P3_U3260, P3_D_REG_5__SCAN_IN, P3_U3832);
  and ginst24662 (P3_U3261, P3_D_REG_4__SCAN_IN, P3_U3832);
  and ginst24663 (P3_U3262, P3_D_REG_3__SCAN_IN, P3_U3832);
  and ginst24664 (P3_U3263, P3_D_REG_2__SCAN_IN, P3_U3832);
  nand ginst24665 (P3_U3264, P3_U4015, P3_U4016, P3_U4017);
  nand ginst24666 (P3_U3265, P3_U4012, P3_U4013, P3_U4014);
  nand ginst24667 (P3_U3266, P3_U4009, P3_U4010, P3_U4011);
  nand ginst24668 (P3_U3267, P3_U4006, P3_U4007, P3_U4008);
  nand ginst24669 (P3_U3268, P3_U4003, P3_U4004, P3_U4005);
  nand ginst24670 (P3_U3269, P3_U4000, P3_U4001, P3_U4002);
  nand ginst24671 (P3_U3270, P3_U3997, P3_U3998, P3_U3999);
  nand ginst24672 (P3_U3271, P3_U3994, P3_U3995, P3_U3996);
  nand ginst24673 (P3_U3272, P3_U3991, P3_U3992, P3_U3993);
  nand ginst24674 (P3_U3273, P3_U3988, P3_U3989, P3_U3990);
  nand ginst24675 (P3_U3274, P3_U3985, P3_U3986, P3_U3987);
  nand ginst24676 (P3_U3275, P3_U3982, P3_U3983, P3_U3984);
  nand ginst24677 (P3_U3276, P3_U3979, P3_U3980, P3_U3981);
  nand ginst24678 (P3_U3277, P3_U3976, P3_U3977, P3_U3978);
  nand ginst24679 (P3_U3278, P3_U3973, P3_U3974, P3_U3975);
  nand ginst24680 (P3_U3279, P3_U3970, P3_U3971, P3_U3972);
  nand ginst24681 (P3_U3280, P3_U3967, P3_U3968, P3_U3969);
  nand ginst24682 (P3_U3281, P3_U3964, P3_U3965, P3_U3966);
  nand ginst24683 (P3_U3282, P3_U3961, P3_U3962, P3_U3963);
  nand ginst24684 (P3_U3283, P3_U3958, P3_U3959, P3_U3960);
  nand ginst24685 (P3_U3284, P3_U3955, P3_U3956, P3_U3957);
  nand ginst24686 (P3_U3285, P3_U3952, P3_U3953, P3_U3954);
  nand ginst24687 (P3_U3286, P3_U3949, P3_U3950, P3_U3951);
  nand ginst24688 (P3_U3287, P3_U3946, P3_U3947, P3_U3948);
  nand ginst24689 (P3_U3288, P3_U3943, P3_U3944, P3_U3945);
  nand ginst24690 (P3_U3289, P3_U3940, P3_U3941, P3_U3942);
  nand ginst24691 (P3_U3290, P3_U3937, P3_U3938, P3_U3939);
  nand ginst24692 (P3_U3291, P3_U3934, P3_U3935, P3_U3936);
  nand ginst24693 (P3_U3292, P3_U3931, P3_U3932, P3_U3933);
  nand ginst24694 (P3_U3293, P3_U3928, P3_U3929, P3_U3930);
  nand ginst24695 (P3_U3294, P3_U3925, P3_U3926, P3_U3927);
  nand ginst24696 (P3_U3295, P3_U3922, P3_U3923, P3_U3924);
  and ginst24697 (P3_U3296, P3_U3775, P3_U5421);
  nand ginst24698 (P3_U3297, P3_STATE_REG_SCAN_IN, P3_U3831);
  not ginst24699 (P3_U3298, P3_B_REG_SCAN_IN);
  nand ginst24700 (P3_U3299, P3_U3374, P3_U5431);
  nand ginst24701 (P3_U3300, P3_U3374, P3_U4018);
  nand ginst24702 (P3_U3301, P3_U3013, P3_U5447);
  nand ginst24703 (P3_U3302, P3_U3014, P3_U5456);
  nand ginst24704 (P3_U3303, P3_U3018, P3_U3588);
  nand ginst24705 (P3_U3304, P3_U3018, P3_U3589);
  nand ginst24706 (P3_U3305, P3_U3014, P3_U5447);
  nand ginst24707 (P3_U3306, P3_U3014, P3_U3378);
  nand ginst24708 (P3_U3307, P3_U3013, P3_U3378);
  nand ginst24709 (P3_U3308, P3_U3378, P3_U3379, P3_U3385);
  nand ginst24710 (P3_U3309, P3_U3378, P3_U3385, P3_U5450);
  nand ginst24711 (P3_U3310, P3_U3013, P3_U5456);
  nand ginst24712 (P3_U3311, P3_U3878, P3_U5447);
  nand ginst24713 (P3_U3312, P3_U3016, P3_U3385);
  nand ginst24714 (P3_U3313, P3_U3380, P3_U3385);
  nand ginst24715 (P3_U3314, P3_U3575, P3_U3576, P3_U4069, P3_U4070, P3_U4071);
  nand ginst24716 (P3_U3315, P3_U3590, P3_U3592, P3_U4090, P3_U4091);
  nand ginst24717 (P3_U3316, P3_U3594, P3_U3596, P3_U4108, P3_U4109);
  nand ginst24718 (P3_U3317, P3_U3598, P3_U3600, P3_U4126, P3_U4127);
  nand ginst24719 (P3_U3318, P3_U3603, P3_U4144, P3_U4145, P3_U4146, P3_U4147);
  nand ginst24720 (P3_U3319, P3_U3606, P3_U4162, P3_U4163, P3_U4164, P3_U4165);
  nand ginst24721 (P3_U3320, P3_U3609, P3_U4180, P3_U4181, P3_U4182, P3_U4183);
  nand ginst24722 (P3_U3321, P3_U3612, P3_U4198, P3_U4199, P3_U4200, P3_U4201);
  nand ginst24723 (P3_U3322, P3_U3615, P3_U4216, P3_U4217, P3_U4218, P3_U4219);
  nand ginst24724 (P3_U3323, P3_U3617, P3_U3619, P3_U4234, P3_U4235);
  nand ginst24725 (P3_U3324, P3_U3621, P3_U3623, P3_U4252, P3_U4253);
  nand ginst24726 (P3_U3325, P3_U3626, P3_U4270, P3_U4271, P3_U4272, P3_U4273);
  nand ginst24727 (P3_U3326, P3_U3628, P3_U3630, P3_U4288, P3_U4289);
  nand ginst24728 (P3_U3327, P3_U3632, P3_U3634, P3_U4306, P3_U4307);
  nand ginst24729 (P3_U3328, P3_U3637, P3_U4324, P3_U4325, P3_U4326, P3_U4327);
  nand ginst24730 (P3_U3329, P3_U3640, P3_U4342, P3_U4343, P3_U4344, P3_U4345);
  nand ginst24731 (P3_U3330, P3_U3643, P3_U4360, P3_U4361, P3_U4362, P3_U4363);
  nand ginst24732 (P3_U3331, P3_U3645, P3_U3647, P3_U4378, P3_U4379);
  nand ginst24733 (P3_U3332, P3_U3650, P3_U4396, P3_U4397, P3_U4398, P3_U4399);
  nand ginst24734 (P3_U3333, P3_U3653, P3_U4414, P3_U4415, P3_U4416, P3_U4417);
  nand ginst24735 (P3_U3334, P3_U3833, U49);
  nand ginst24736 (P3_U3335, P3_U3656, P3_U4432, P3_U4433, P3_U4434, P3_U4435);
  nand ginst24737 (P3_U3336, P3_U3833, U48);
  nand ginst24738 (P3_U3337, P3_U3659, P3_U4450, P3_U4451, P3_U4452, P3_U4453);
  nand ginst24739 (P3_U3338, P3_U3833, U47);
  nand ginst24740 (P3_U3339, P3_U3662, P3_U4468, P3_U4469, P3_U4470, P3_U4471);
  nand ginst24741 (P3_U3340, P3_U3833, U46);
  nand ginst24742 (P3_U3341, P3_U3665, P3_U4486, P3_U4487, P3_U4488, P3_U4489);
  nand ginst24743 (P3_U3342, P3_U3833, U45);
  nand ginst24744 (P3_U3343, P3_U3667, P3_U3669, P3_U4504, P3_U4505);
  nand ginst24745 (P3_U3344, P3_U3833, U44);
  nand ginst24746 (P3_U3345, P3_U3671, P3_U3673, P3_U4522, P3_U4523);
  nand ginst24747 (P3_U3346, P3_U3833, U43);
  nand ginst24748 (P3_U3347, P3_U3675, P3_U3677, P3_U4540, P3_U4541);
  nand ginst24749 (P3_U3348, P3_U3833, U42);
  nand ginst24750 (P3_U3349, P3_U3679, P3_U3681, P3_U4558, P3_U4559);
  nand ginst24751 (P3_U3350, P3_U3833, U41);
  nand ginst24752 (P3_U3351, P3_U3683, P3_U3685, P3_U4576, P3_U4577);
  nand ginst24753 (P3_U3352, P3_U3383, P3_U3384);
  nand ginst24754 (P3_U3353, P3_U3833, U40);
  nand ginst24755 (P3_U3354, P3_U3687, P3_U3689, P3_U4596, P3_U4597, P3_U4598);
  nand ginst24756 (P3_U3355, P3_U3833, U38);
  nand ginst24757 (P3_U3356, P3_U3833, U37);
  nand ginst24758 (P3_U3357, P3_U3015, P3_U5456);
  nand ginst24759 (P3_U3358, P3_U3023, P3_U4627);
  nand ginst24760 (P3_U3359, P3_U3385, P3_U5447);
  nand ginst24761 (P3_U3360, P3_U3879, P3_U5447);
  nand ginst24762 (P3_U3361, P3_U3055, P3_U3911, P3_U4595);
  nand ginst24763 (P3_U3362, P3_U3372, P3_U3373, P3_U3374);
  nand ginst24764 (P3_U3363, P3_U3694, P3_U3910);
  nand ginst24765 (P3_U3364, P3_U3313, P3_U3833);
  nand ginst24766 (P3_U3365, P3_U3877, P3_U5423);
  nand ginst24767 (P3_U3366, P3_U3050, P3_U3695);
  nand ginst24768 (P3_U3367, P3_U3385, P3_U3882);
  nand ginst24769 (P3_U3368, P3_U3759, P3_U3890);
  nand ginst24770 (P3_U3369, P3_U3378, P3_U3876);
  nand ginst24771 (P3_U3370, P3_U3776, P3_U4991, P3_U4992);
  nand ginst24772 (P3_U3371, P3_U3917, P3_U5417);
  nand ginst24773 (P3_U3372, P3_U5426, P3_U5427);
  nand ginst24774 (P3_U3373, P3_U5429, P3_U5430);
  nand ginst24775 (P3_U3374, P3_U5432, P3_U5433);
  nand ginst24776 (P3_U3375, P3_U5438, P3_U5439);
  nand ginst24777 (P3_U3376, P3_U5441, P3_U5442);
  nand ginst24778 (P3_U3377, P3_U5443, P3_U5444);
  nand ginst24779 (P3_U3378, P3_U5445, P3_U5446);
  nand ginst24780 (P3_U3379, P3_U5448, P3_U5449);
  nand ginst24781 (P3_U3380, P3_U5451, P3_U5452);
  nand ginst24782 (P3_U3381, P3_U5457, P3_U5458);
  nand ginst24783 (P3_U3382, P3_U5460, P3_U5461);
  nand ginst24784 (P3_U3383, P3_U5463, P3_U5464);
  nand ginst24785 (P3_U3384, P3_U5466, P3_U5467);
  nand ginst24786 (P3_U3385, P3_U5454, P3_U5455);
  nand ginst24787 (P3_U3386, P3_U5469, P3_U5470);
  nand ginst24788 (P3_U3387, P3_U5471, P3_U5472);
  nand ginst24789 (P3_U3388, P3_U5474, P3_U5475);
  nand ginst24790 (P3_U3389, P3_U5477, P3_U5478);
  nand ginst24791 (P3_U3390, P3_U5483, P3_U5484);
  nand ginst24792 (P3_U3391, P3_U5485, P3_U5486);
  nand ginst24793 (P3_U3392, P3_U5487, P3_U5488);
  nand ginst24794 (P3_U3393, P3_U5490, P3_U5491);
  nand ginst24795 (P3_U3394, P3_U5492, P3_U5493);
  nand ginst24796 (P3_U3395, P3_U5494, P3_U5495);
  nand ginst24797 (P3_U3396, P3_U5497, P3_U5498);
  nand ginst24798 (P3_U3397, P3_U5499, P3_U5500);
  nand ginst24799 (P3_U3398, P3_U5501, P3_U5502);
  nand ginst24800 (P3_U3399, P3_U5504, P3_U5505);
  nand ginst24801 (P3_U3400, P3_U5506, P3_U5507);
  nand ginst24802 (P3_U3401, P3_U5508, P3_U5509);
  nand ginst24803 (P3_U3402, P3_U5511, P3_U5512);
  nand ginst24804 (P3_U3403, P3_U5513, P3_U5514);
  nand ginst24805 (P3_U3404, P3_U5515, P3_U5516);
  nand ginst24806 (P3_U3405, P3_U5518, P3_U5519);
  nand ginst24807 (P3_U3406, P3_U5520, P3_U5521);
  nand ginst24808 (P3_U3407, P3_U5522, P3_U5523);
  nand ginst24809 (P3_U3408, P3_U5525, P3_U5526);
  nand ginst24810 (P3_U3409, P3_U5527, P3_U5528);
  nand ginst24811 (P3_U3410, P3_U5529, P3_U5530);
  nand ginst24812 (P3_U3411, P3_U5532, P3_U5533);
  nand ginst24813 (P3_U3412, P3_U5534, P3_U5535);
  nand ginst24814 (P3_U3413, P3_U5536, P3_U5537);
  nand ginst24815 (P3_U3414, P3_U5539, P3_U5540);
  nand ginst24816 (P3_U3415, P3_U5541, P3_U5542);
  nand ginst24817 (P3_U3416, P3_U5543, P3_U5544);
  nand ginst24818 (P3_U3417, P3_U5546, P3_U5547);
  nand ginst24819 (P3_U3418, P3_U5548, P3_U5549);
  nand ginst24820 (P3_U3419, P3_U5550, P3_U5551);
  nand ginst24821 (P3_U3420, P3_U5553, P3_U5554);
  nand ginst24822 (P3_U3421, P3_U5555, P3_U5556);
  nand ginst24823 (P3_U3422, P3_U5557, P3_U5558);
  nand ginst24824 (P3_U3423, P3_U5560, P3_U5561);
  nand ginst24825 (P3_U3424, P3_U5562, P3_U5563);
  nand ginst24826 (P3_U3425, P3_U5564, P3_U5565);
  nand ginst24827 (P3_U3426, P3_U5567, P3_U5568);
  nand ginst24828 (P3_U3427, P3_U5569, P3_U5570);
  nand ginst24829 (P3_U3428, P3_U5571, P3_U5572);
  nand ginst24830 (P3_U3429, P3_U5574, P3_U5575);
  nand ginst24831 (P3_U3430, P3_U5576, P3_U5577);
  nand ginst24832 (P3_U3431, P3_U5578, P3_U5579);
  nand ginst24833 (P3_U3432, P3_U5581, P3_U5582);
  nand ginst24834 (P3_U3433, P3_U5583, P3_U5584);
  nand ginst24835 (P3_U3434, P3_U5585, P3_U5586);
  nand ginst24836 (P3_U3435, P3_U5588, P3_U5589);
  nand ginst24837 (P3_U3436, P3_U5590, P3_U5591);
  nand ginst24838 (P3_U3437, P3_U5592, P3_U5593);
  nand ginst24839 (P3_U3438, P3_U5595, P3_U5596);
  nand ginst24840 (P3_U3439, P3_U5597, P3_U5598);
  nand ginst24841 (P3_U3440, P3_U5599, P3_U5600);
  nand ginst24842 (P3_U3441, P3_U5602, P3_U5603);
  nand ginst24843 (P3_U3442, P3_U5604, P3_U5605);
  nand ginst24844 (P3_U3443, P3_U5606, P3_U5607);
  nand ginst24845 (P3_U3444, P3_U5609, P3_U5610);
  nand ginst24846 (P3_U3445, P3_U5611, P3_U5612);
  nand ginst24847 (P3_U3446, P3_U5614, P3_U5615);
  nand ginst24848 (P3_U3447, P3_U5616, P3_U5617);
  nand ginst24849 (P3_U3448, P3_U5618, P3_U5619);
  nand ginst24850 (P3_U3449, P3_U5620, P3_U5621);
  nand ginst24851 (P3_U3450, P3_U5622, P3_U5623);
  nand ginst24852 (P3_U3451, P3_U5624, P3_U5625);
  nand ginst24853 (P3_U3452, P3_U5626, P3_U5627);
  nand ginst24854 (P3_U3453, P3_U5628, P3_U5629);
  nand ginst24855 (P3_U3454, P3_U5630, P3_U5631);
  nand ginst24856 (P3_U3455, P3_U5632, P3_U5633);
  nand ginst24857 (P3_U3456, P3_U5634, P3_U5635);
  nand ginst24858 (P3_U3457, P3_U5636, P3_U5637);
  nand ginst24859 (P3_U3458, P3_U5638, P3_U5639);
  nand ginst24860 (P3_U3459, P3_U5642, P3_U5643);
  nand ginst24861 (P3_U3460, P3_U5644, P3_U5645);
  nand ginst24862 (P3_U3461, P3_U5646, P3_U5647);
  nand ginst24863 (P3_U3462, P3_U5648, P3_U5649);
  nand ginst24864 (P3_U3463, P3_U5650, P3_U5651);
  nand ginst24865 (P3_U3464, P3_U5652, P3_U5653);
  nand ginst24866 (P3_U3465, P3_U5654, P3_U5655);
  nand ginst24867 (P3_U3466, P3_U5656, P3_U5657);
  nand ginst24868 (P3_U3467, P3_U5658, P3_U5659);
  nand ginst24869 (P3_U3468, P3_U5660, P3_U5661);
  nand ginst24870 (P3_U3469, P3_U5662, P3_U5663);
  nand ginst24871 (P3_U3470, P3_U5664, P3_U5665);
  nand ginst24872 (P3_U3471, P3_U5666, P3_U5667);
  nand ginst24873 (P3_U3472, P3_U5668, P3_U5669);
  nand ginst24874 (P3_U3473, P3_U5670, P3_U5671);
  nand ginst24875 (P3_U3474, P3_U5672, P3_U5673);
  nand ginst24876 (P3_U3475, P3_U5674, P3_U5675);
  nand ginst24877 (P3_U3476, P3_U5676, P3_U5677);
  nand ginst24878 (P3_U3477, P3_U5678, P3_U5679);
  nand ginst24879 (P3_U3478, P3_U5680, P3_U5681);
  nand ginst24880 (P3_U3479, P3_U5682, P3_U5683);
  nand ginst24881 (P3_U3480, P3_U5684, P3_U5685);
  nand ginst24882 (P3_U3481, P3_U5686, P3_U5687);
  nand ginst24883 (P3_U3482, P3_U5688, P3_U5689);
  nand ginst24884 (P3_U3483, P3_U5690, P3_U5691);
  nand ginst24885 (P3_U3484, P3_U5692, P3_U5693);
  nand ginst24886 (P3_U3485, P3_U5694, P3_U5695);
  nand ginst24887 (P3_U3486, P3_U5696, P3_U5697);
  nand ginst24888 (P3_U3487, P3_U5698, P3_U5699);
  nand ginst24889 (P3_U3488, P3_U5700, P3_U5701);
  nand ginst24890 (P3_U3489, P3_U5702, P3_U5703);
  nand ginst24891 (P3_U3490, P3_U5704, P3_U5705);
  nand ginst24892 (P3_U3491, P3_U5769, P3_U5770);
  nand ginst24893 (P3_U3492, P3_U5771, P3_U5772);
  nand ginst24894 (P3_U3493, P3_U5773, P3_U5774);
  nand ginst24895 (P3_U3494, P3_U5775, P3_U5776);
  nand ginst24896 (P3_U3495, P3_U5777, P3_U5778);
  nand ginst24897 (P3_U3496, P3_U5779, P3_U5780);
  nand ginst24898 (P3_U3497, P3_U5781, P3_U5782);
  nand ginst24899 (P3_U3498, P3_U5783, P3_U5784);
  nand ginst24900 (P3_U3499, P3_U5785, P3_U5786);
  nand ginst24901 (P3_U3500, P3_U5787, P3_U5788);
  nand ginst24902 (P3_U3501, P3_U5789, P3_U5790);
  nand ginst24903 (P3_U3502, P3_U5791, P3_U5792);
  nand ginst24904 (P3_U3503, P3_U5793, P3_U5794);
  nand ginst24905 (P3_U3504, P3_U5795, P3_U5796);
  nand ginst24906 (P3_U3505, P3_U5797, P3_U5798);
  nand ginst24907 (P3_U3506, P3_U5799, P3_U5800);
  nand ginst24908 (P3_U3507, P3_U5801, P3_U5802);
  nand ginst24909 (P3_U3508, P3_U5803, P3_U5804);
  nand ginst24910 (P3_U3509, P3_U5805, P3_U5806);
  nand ginst24911 (P3_U3510, P3_U5807, P3_U5808);
  nand ginst24912 (P3_U3511, P3_U5809, P3_U5810);
  nand ginst24913 (P3_U3512, P3_U5811, P3_U5812);
  nand ginst24914 (P3_U3513, P3_U5813, P3_U5814);
  nand ginst24915 (P3_U3514, P3_U5815, P3_U5816);
  nand ginst24916 (P3_U3515, P3_U5817, P3_U5818);
  nand ginst24917 (P3_U3516, P3_U5819, P3_U5820);
  nand ginst24918 (P3_U3517, P3_U5821, P3_U5822);
  nand ginst24919 (P3_U3518, P3_U5823, P3_U5824);
  nand ginst24920 (P3_U3519, P3_U5825, P3_U5826);
  nand ginst24921 (P3_U3520, P3_U5827, P3_U5828);
  nand ginst24922 (P3_U3521, P3_U5829, P3_U5830);
  nand ginst24923 (P3_U3522, P3_U5831, P3_U5832);
  nand ginst24924 (P3_U3523, P3_U5945, P3_U5946);
  nand ginst24925 (P3_U3524, P3_U5947, P3_U5948);
  nand ginst24926 (P3_U3525, P3_U5949, P3_U5950);
  nand ginst24927 (P3_U3526, P3_U5951, P3_U5952);
  nand ginst24928 (P3_U3527, P3_U5953, P3_U5954);
  nand ginst24929 (P3_U3528, P3_U5955, P3_U5956);
  nand ginst24930 (P3_U3529, P3_U5957, P3_U5958);
  nand ginst24931 (P3_U3530, P3_U5959, P3_U5960);
  nand ginst24932 (P3_U3531, P3_U5961, P3_U5962);
  nand ginst24933 (P3_U3532, P3_U5963, P3_U5964);
  nand ginst24934 (P3_U3533, P3_U5965, P3_U5966);
  nand ginst24935 (P3_U3534, P3_U5967, P3_U5968);
  nand ginst24936 (P3_U3535, P3_U5969, P3_U5970);
  nand ginst24937 (P3_U3536, P3_U5971, P3_U5972);
  nand ginst24938 (P3_U3537, P3_U5973, P3_U5974);
  nand ginst24939 (P3_U3538, P3_U5975, P3_U5976);
  nand ginst24940 (P3_U3539, P3_U5977, P3_U5978);
  nand ginst24941 (P3_U3540, P3_U5979, P3_U5980);
  nand ginst24942 (P3_U3541, P3_U5981, P3_U5982);
  nand ginst24943 (P3_U3542, P3_U5983, P3_U5984);
  nand ginst24944 (P3_U3543, P3_U5985, P3_U5986);
  nand ginst24945 (P3_U3544, P3_U5987, P3_U5988);
  nand ginst24946 (P3_U3545, P3_U5989, P3_U5990);
  nand ginst24947 (P3_U3546, P3_U5991, P3_U5992);
  nand ginst24948 (P3_U3547, P3_U5993, P3_U5994);
  nand ginst24949 (P3_U3548, P3_U5995, P3_U5996);
  nand ginst24950 (P3_U3549, P3_U5997, P3_U5998);
  nand ginst24951 (P3_U3550, P3_U5999, P3_U6000);
  nand ginst24952 (P3_U3551, P3_U6001, P3_U6002);
  nand ginst24953 (P3_U3552, P3_U6003, P3_U6004);
  nand ginst24954 (P3_U3553, P3_U6005, P3_U6006);
  nand ginst24955 (P3_U3554, P3_U6007, P3_U6008);
  nand ginst24956 (P3_U3555, P3_U6009, P3_U6010);
  nand ginst24957 (P3_U3556, P3_U6011, P3_U6012);
  nand ginst24958 (P3_U3557, P3_U6013, P3_U6014);
  nand ginst24959 (P3_U3558, P3_U6015, P3_U6016);
  nand ginst24960 (P3_U3559, P3_U6017, P3_U6018);
  nand ginst24961 (P3_U3560, P3_U6019, P3_U6020);
  nand ginst24962 (P3_U3561, P3_U6021, P3_U6022);
  nand ginst24963 (P3_U3562, P3_U6023, P3_U6024);
  nand ginst24964 (P3_U3563, P3_U6025, P3_U6026);
  nand ginst24965 (P3_U3564, P3_U6027, P3_U6028);
  nand ginst24966 (P3_U3565, P3_U6029, P3_U6030);
  nand ginst24967 (P3_U3566, P3_U6031, P3_U6032);
  nand ginst24968 (P3_U3567, P3_U6033, P3_U6034);
  nand ginst24969 (P3_U3568, P3_U6035, P3_U6036);
  nand ginst24970 (P3_U3569, P3_U6037, P3_U6038);
  nand ginst24971 (P3_U3570, P3_U6039, P3_U6040);
  nand ginst24972 (P3_U3571, P3_U6041, P3_U6042);
  nand ginst24973 (P3_U3572, P3_U6043, P3_U6044);
  nand ginst24974 (P3_U3573, P3_U6045, P3_U6046);
  nand ginst24975 (P3_U3574, P3_U6047, P3_U6048);
  and ginst24976 (P3_U3575, P3_U4065, P3_U4066);
  and ginst24977 (P3_U3576, P3_U4067, P3_U4068);
  and ginst24978 (P3_U3577, P3_U4074, P3_U4075, P3_U4076);
  and ginst24979 (P3_U3578, P3_U4022, P3_U4023, P3_U4024, P3_U4025);
  and ginst24980 (P3_U3579, P3_U4026, P3_U4027, P3_U4028, P3_U4029);
  and ginst24981 (P3_U3580, P3_U4030, P3_U4031, P3_U4032, P3_U4033);
  and ginst24982 (P3_U3581, P3_U4034, P3_U4035, P3_U4036);
  and ginst24983 (P3_U3582, P3_U3578, P3_U3579, P3_U3580, P3_U3581);
  and ginst24984 (P3_U3583, P3_U4037, P3_U4038, P3_U4039, P3_U4040);
  and ginst24985 (P3_U3584, P3_U4041, P3_U4042, P3_U4043, P3_U4044);
  and ginst24986 (P3_U3585, P3_U4045, P3_U4046, P3_U4047, P3_U4048);
  and ginst24987 (P3_U3586, P3_U4049, P3_U4050, P3_U4051);
  and ginst24988 (P3_U3587, P3_U3583, P3_U3584, P3_U3585, P3_U3586);
  and ginst24989 (P3_U3588, P3_U3388, P3_U3389);
  and ginst24990 (P3_U3589, P3_U5476, P3_U5479);
  and ginst24991 (P3_U3590, P3_U4092, P3_U4093);
  and ginst24992 (P3_U3591, P3_U4094, P3_U4095);
  and ginst24993 (P3_U3592, P3_U3591, P3_U4096, P3_U4097);
  and ginst24994 (P3_U3593, P3_U4099, P3_U4100, P3_U4101);
  and ginst24995 (P3_U3594, P3_U4110, P3_U4111);
  and ginst24996 (P3_U3595, P3_U4112, P3_U4113);
  and ginst24997 (P3_U3596, P3_U3595, P3_U4114, P3_U4115);
  and ginst24998 (P3_U3597, P3_U4117, P3_U4118, P3_U4119);
  and ginst24999 (P3_U3598, P3_U4128, P3_U4129);
  and ginst25000 (P3_U3599, P3_U4130, P3_U4131);
  and ginst25001 (P3_U3600, P3_U3599, P3_U4132, P3_U4133);
  and ginst25002 (P3_U3601, P3_U4135, P3_U4136, P3_U4137);
  and ginst25003 (P3_U3602, P3_U4148, P3_U4149);
  and ginst25004 (P3_U3603, P3_U3602, P3_U4150, P3_U4151);
  and ginst25005 (P3_U3604, P3_U4153, P3_U4154, P3_U4155);
  and ginst25006 (P3_U3605, P3_U4166, P3_U4167);
  and ginst25007 (P3_U3606, P3_U3605, P3_U4168, P3_U4169);
  and ginst25008 (P3_U3607, P3_U4171, P3_U4172, P3_U4173);
  and ginst25009 (P3_U3608, P3_U4184, P3_U4185);
  and ginst25010 (P3_U3609, P3_U3608, P3_U4186, P3_U4187);
  and ginst25011 (P3_U3610, P3_U4189, P3_U4190, P3_U4191);
  and ginst25012 (P3_U3611, P3_U4202, P3_U4203);
  and ginst25013 (P3_U3612, P3_U3611, P3_U4204, P3_U4205);
  and ginst25014 (P3_U3613, P3_U4207, P3_U4208, P3_U4209);
  and ginst25015 (P3_U3614, P3_U4220, P3_U4221);
  and ginst25016 (P3_U3615, P3_U3614, P3_U4222, P3_U4223);
  and ginst25017 (P3_U3616, P3_U4225, P3_U4226, P3_U4227);
  and ginst25018 (P3_U3617, P3_U4236, P3_U4237);
  and ginst25019 (P3_U3618, P3_U4238, P3_U4239);
  and ginst25020 (P3_U3619, P3_U3618, P3_U4240, P3_U4241);
  and ginst25021 (P3_U3620, P3_U4243, P3_U4244, P3_U4245);
  and ginst25022 (P3_U3621, P3_U4254, P3_U4255);
  and ginst25023 (P3_U3622, P3_U4256, P3_U4257);
  and ginst25024 (P3_U3623, P3_U3622, P3_U4258, P3_U4259);
  and ginst25025 (P3_U3624, P3_U4261, P3_U4262, P3_U4263);
  and ginst25026 (P3_U3625, P3_U4274, P3_U4275);
  and ginst25027 (P3_U3626, P3_U3625, P3_U4276, P3_U4277);
  and ginst25028 (P3_U3627, P3_U4279, P3_U4280, P3_U4281);
  and ginst25029 (P3_U3628, P3_U4290, P3_U4291);
  and ginst25030 (P3_U3629, P3_U4292, P3_U4293);
  and ginst25031 (P3_U3630, P3_U3629, P3_U4294, P3_U4295);
  and ginst25032 (P3_U3631, P3_U4297, P3_U4298, P3_U4299);
  and ginst25033 (P3_U3632, P3_U4308, P3_U4309);
  and ginst25034 (P3_U3633, P3_U4310, P3_U4311);
  and ginst25035 (P3_U3634, P3_U3633, P3_U4312, P3_U4313);
  and ginst25036 (P3_U3635, P3_U4315, P3_U4316, P3_U4317);
  and ginst25037 (P3_U3636, P3_U4328, P3_U4329);
  and ginst25038 (P3_U3637, P3_U3636, P3_U4330, P3_U4331);
  and ginst25039 (P3_U3638, P3_U4333, P3_U4334, P3_U4335);
  and ginst25040 (P3_U3639, P3_U4346, P3_U4347);
  and ginst25041 (P3_U3640, P3_U3639, P3_U4348, P3_U4349);
  and ginst25042 (P3_U3641, P3_U4351, P3_U4352, P3_U4353);
  and ginst25043 (P3_U3642, P3_U4364, P3_U4365);
  and ginst25044 (P3_U3643, P3_U3642, P3_U4366, P3_U4367);
  and ginst25045 (P3_U3644, P3_U4369, P3_U4370, P3_U4371);
  and ginst25046 (P3_U3645, P3_U4380, P3_U4381);
  and ginst25047 (P3_U3646, P3_U4382, P3_U4383);
  and ginst25048 (P3_U3647, P3_U3646, P3_U4384, P3_U4385);
  and ginst25049 (P3_U3648, P3_U4387, P3_U4388, P3_U4389);
  and ginst25050 (P3_U3649, P3_U4400, P3_U4401);
  and ginst25051 (P3_U3650, P3_U3649, P3_U4402, P3_U4403);
  and ginst25052 (P3_U3651, P3_U4405, P3_U4406, P3_U4407);
  and ginst25053 (P3_U3652, P3_U4418, P3_U4419);
  and ginst25054 (P3_U3653, P3_U3652, P3_U4420, P3_U4421);
  and ginst25055 (P3_U3654, P3_U4423, P3_U4424, P3_U4425);
  and ginst25056 (P3_U3655, P3_U4436, P3_U4437);
  and ginst25057 (P3_U3656, P3_U3655, P3_U4438, P3_U4439);
  and ginst25058 (P3_U3657, P3_U4441, P3_U4442, P3_U4443);
  and ginst25059 (P3_U3658, P3_U4454, P3_U4455);
  and ginst25060 (P3_U3659, P3_U3658, P3_U4456, P3_U4457);
  and ginst25061 (P3_U3660, P3_U4459, P3_U4460, P3_U4461);
  and ginst25062 (P3_U3661, P3_U4472, P3_U4473);
  and ginst25063 (P3_U3662, P3_U3661, P3_U4474, P3_U4475);
  and ginst25064 (P3_U3663, P3_U4477, P3_U4478, P3_U4479);
  and ginst25065 (P3_U3664, P3_U4490, P3_U4491);
  and ginst25066 (P3_U3665, P3_U3664, P3_U4492, P3_U4493);
  and ginst25067 (P3_U3666, P3_U4495, P3_U4496, P3_U4497);
  and ginst25068 (P3_U3667, P3_U4506, P3_U4507);
  and ginst25069 (P3_U3668, P3_U4508, P3_U4509);
  and ginst25070 (P3_U3669, P3_U3668, P3_U4510, P3_U4511);
  and ginst25071 (P3_U3670, P3_U4513, P3_U4514, P3_U4515);
  and ginst25072 (P3_U3671, P3_U4524, P3_U4525);
  and ginst25073 (P3_U3672, P3_U4526, P3_U4527);
  and ginst25074 (P3_U3673, P3_U3672, P3_U4528, P3_U4529);
  and ginst25075 (P3_U3674, P3_U4531, P3_U4532, P3_U4533);
  and ginst25076 (P3_U3675, P3_U4542, P3_U4543);
  and ginst25077 (P3_U3676, P3_U4544, P3_U4545);
  and ginst25078 (P3_U3677, P3_U3676, P3_U4546, P3_U4547);
  and ginst25079 (P3_U3678, P3_U4549, P3_U4550, P3_U4551);
  and ginst25080 (P3_U3679, P3_U4560, P3_U4561);
  and ginst25081 (P3_U3680, P3_U4562, P3_U4563);
  and ginst25082 (P3_U3681, P3_U3680, P3_U4564, P3_U4565);
  and ginst25083 (P3_U3682, P3_U4567, P3_U4568, P3_U4569);
  and ginst25084 (P3_U3683, P3_U4578, P3_U4579);
  and ginst25085 (P3_U3684, P3_U4580, P3_U4581);
  and ginst25086 (P3_U3685, P3_U3684, P3_U4582, P3_U4583);
  and ginst25087 (P3_U3686, P3_U4585, P3_U4586, P3_U4587);
  and ginst25088 (P3_U3687, P3_U4599, P3_U4600);
  and ginst25089 (P3_U3688, P3_U4601, P3_U4602);
  and ginst25090 (P3_U3689, P3_U3688, P3_U4603, P3_U4604);
  and ginst25091 (P3_U3690, P3_U4606, P3_U4607);
  and ginst25092 (P3_U3691, P3_U3389, P3_U5476);
  and ginst25093 (P3_U3692, P3_U3388, P3_U5479);
  and ginst25094 (P3_U3693, P3_U3379, P3_U3920);
  and ginst25095 (P3_U3694, P3_STATE_REG_SCAN_IN, P3_U5440);
  and ginst25096 (P3_U3695, P3_U3364, P3_U5424);
  and ginst25097 (P3_U3696, P3_STATE_REG_SCAN_IN, P3_U3375);
  and ginst25098 (P3_U3697, P3_U3301, P3_U3305, P3_U3306, P3_U3307, P3_U3308);
  and ginst25099 (P3_U3698, P3_U3309, P3_U3360);
  and ginst25100 (P3_U3699, P3_U3701, P3_U4762, P3_U4763, P3_U4765);
  and ginst25101 (P3_U3700, P3_U4766, P3_U4768);
  and ginst25102 (P3_U3701, P3_U3700, P3_U4767);
  and ginst25103 (P3_U3702, P3_U3704, P3_U4773, P3_U4774, P3_U4776);
  and ginst25104 (P3_U3703, P3_U4777, P3_U4779);
  and ginst25105 (P3_U3704, P3_U3703, P3_U4778);
  and ginst25106 (P3_U3705, P3_U3707, P3_U4784, P3_U4785, P3_U4787);
  and ginst25107 (P3_U3706, P3_U4788, P3_U4790);
  and ginst25108 (P3_U3707, P3_U3706, P3_U4789);
  and ginst25109 (P3_U3708, P3_U3710, P3_U4795, P3_U4796, P3_U4798);
  and ginst25110 (P3_U3709, P3_U4799, P3_U4801);
  and ginst25111 (P3_U3710, P3_U3709, P3_U4800);
  and ginst25112 (P3_U3711, P3_U3713, P3_U4806, P3_U4807, P3_U4809);
  and ginst25113 (P3_U3712, P3_U4810, P3_U4812);
  and ginst25114 (P3_U3713, P3_U3712, P3_U4811);
  and ginst25115 (P3_U3714, P3_U3716, P3_U4817, P3_U4818, P3_U4820);
  and ginst25116 (P3_U3715, P3_U4821, P3_U4823);
  and ginst25117 (P3_U3716, P3_U3715, P3_U4822);
  and ginst25118 (P3_U3717, P3_U3719, P3_U4828, P3_U4829, P3_U4831);
  and ginst25119 (P3_U3718, P3_U4832, P3_U4834);
  and ginst25120 (P3_U3719, P3_U3718, P3_U4833);
  and ginst25121 (P3_U3720, P3_U3722, P3_U4839, P3_U4840, P3_U4842);
  and ginst25122 (P3_U3721, P3_U4843, P3_U4845);
  and ginst25123 (P3_U3722, P3_U3721, P3_U4844);
  and ginst25124 (P3_U3723, P3_U3725, P3_U4850, P3_U4851, P3_U4853);
  and ginst25125 (P3_U3724, P3_U4854, P3_U4856);
  and ginst25126 (P3_U3725, P3_U3724, P3_U4855);
  and ginst25127 (P3_U3726, P3_U3728, P3_U4861, P3_U4862, P3_U4864);
  and ginst25128 (P3_U3727, P3_U4865, P3_U4867);
  and ginst25129 (P3_U3728, P3_U3727, P3_U4866);
  and ginst25130 (P3_U3729, P3_U3731, P3_U4872, P3_U4873, P3_U4875);
  and ginst25131 (P3_U3730, P3_U4876, P3_U4878);
  and ginst25132 (P3_U3731, P3_U3730, P3_U4877);
  and ginst25133 (P3_U3732, P3_U3734, P3_U4883, P3_U4884, P3_U4886);
  and ginst25134 (P3_U3733, P3_U4887, P3_U4889);
  and ginst25135 (P3_U3734, P3_U3733, P3_U4888);
  and ginst25136 (P3_U3735, P3_U3737, P3_U4894, P3_U4895, P3_U4897);
  and ginst25137 (P3_U3736, P3_U4898, P3_U4900);
  and ginst25138 (P3_U3737, P3_U3736, P3_U4899);
  and ginst25139 (P3_U3738, P3_U3740, P3_U4906, P3_U4908);
  and ginst25140 (P3_U3739, P3_U4909, P3_U4911);
  and ginst25141 (P3_U3740, P3_U3739, P3_U4910);
  and ginst25142 (P3_U3741, P3_U4917, P3_U4919);
  and ginst25143 (P3_U3742, P3_U4920, P3_U4922);
  and ginst25144 (P3_U3743, P3_U3742, P3_U4921);
  and ginst25145 (P3_U3744, P3_U3746, P3_U4927, P3_U4928);
  and ginst25146 (P3_U3745, P3_U4931, P3_U4933);
  and ginst25147 (P3_U3746, P3_U3745, P3_U4932);
  and ginst25148 (P3_U3747, P3_U3749, P3_U4938, P3_U4939);
  and ginst25149 (P3_U3748, P3_U4942, P3_U4944);
  and ginst25150 (P3_U3749, P3_U3748, P3_U4943);
  and ginst25151 (P3_U3750, P3_U3752, P3_U4949, P3_U4950, P3_U4952);
  and ginst25152 (P3_U3751, P3_U4953, P3_U4955);
  and ginst25153 (P3_U3752, P3_U3751, P3_U4954);
  and ginst25154 (P3_U3753, P3_U3755, P3_U4960, P3_U4961, P3_U4963);
  and ginst25155 (P3_U3754, P3_U4964, P3_U4966);
  and ginst25156 (P3_U3755, P3_U3754, P3_U4965);
  and ginst25157 (P3_U3756, P3_U3758, P3_U4971, P3_U4972, P3_U4974);
  and ginst25158 (P3_U3757, P3_U4975, P3_U4977);
  and ginst25159 (P3_U3758, P3_U3757, P3_U4976);
  and ginst25160 (P3_U3759, P3_U3383, P3_U5468);
  nand ginst25161 (P3_U3760, P3_U5833, P3_U5834);
  and ginst25162 (P3_U3761, P3_U5912, P3_U5915);
  and ginst25163 (P3_U3762, P3_U3761, P3_U3763, P3_U3764, P3_U5897);
  and ginst25164 (P3_U3763, P3_U5900, P3_U5903);
  and ginst25165 (P3_U3764, P3_U5906, P3_U5909);
  and ginst25166 (P3_U3765, P3_U5879, P3_U5882, P3_U5885);
  and ginst25167 (P3_U3766, P3_U5888, P3_U5891, P3_U5894);
  and ginst25168 (P3_U3767, P3_U3765, P3_U3766, P3_U5873, P3_U5876);
  and ginst25169 (P3_U3768, P3_U5858, P3_U5861, P3_U5864, P3_U5867);
  and ginst25170 (P3_U3769, P3_U5852, P3_U5855);
  and ginst25171 (P3_U3770, P3_U5921, P3_U5924, P3_U5927, P3_U5930);
  and ginst25172 (P3_U3771, P3_U5840, P3_U5843, P3_U5846);
  and ginst25173 (P3_U3772, P3_U3768, P3_U3769, P3_U3771, P3_U5849, P3_U5870);
  and ginst25174 (P3_U3773, P3_U3762, P3_U3767, P3_U3770, P3_U5918, P3_U5933);
  and ginst25175 (P3_U3774, P3_U3870, P3_U4980, P3_U4981);
  and ginst25176 (P3_U3775, P3_U5415, P3_U5416);
  and ginst25177 (P3_U3776, P3_U3362, P3_U3880, P3_U4990, P3_U5440);
  and ginst25178 (P3_U3777, P3_U4997, P3_U4998);
  and ginst25179 (P3_U3778, P3_U5010, P3_U5011);
  and ginst25180 (P3_U3779, P3_U5019, P3_U5020);
  and ginst25181 (P3_U3780, P3_U5028, P3_U5029);
  and ginst25182 (P3_U3781, P3_U5034, P3_U5036);
  and ginst25183 (P3_U3782, P3_U5037, P3_U5038);
  and ginst25184 (P3_U3783, P3_U5046, P3_U5047);
  and ginst25185 (P3_U3784, P3_U5055, P3_U5056);
  and ginst25186 (P3_U3785, P3_U5064, P3_U5065);
  and ginst25187 (P3_U3786, P3_U5073, P3_U5074);
  and ginst25188 (P3_U3787, P3_U3031, P3_U3077);
  and ginst25189 (P3_U3788, P3_U5077, P3_U5078);
  and ginst25190 (P3_U3789, P3_U3788, P3_U5080, P3_U5081);
  and ginst25191 (P3_U3790, P3_U5089, P3_U5090);
  and ginst25192 (P3_U3791, P3_U5095, P3_U5097);
  and ginst25193 (P3_U3792, P3_U5098, P3_U5099);
  and ginst25194 (P3_U3793, P3_U5107, P3_U5108);
  and ginst25195 (P3_U3794, P3_U5116, P3_U5117);
  and ginst25196 (P3_U3795, P3_U5125, P3_U5126);
  and ginst25197 (P3_U3796, P3_U5134, P3_U5135);
  and ginst25198 (P3_U3797, P3_U5143, P3_U5144);
  and ginst25199 (P3_U3798, P3_U5152, P3_U5153);
  and ginst25200 (P3_U3799, P3_U5161, P3_U5162);
  and ginst25201 (P3_U3800, P3_U5167, P3_U5169);
  and ginst25202 (P3_U3801, P3_U5170, P3_U5171);
  and ginst25203 (P3_U3802, P3_U5179, P3_U5180);
  and ginst25204 (P3_U3803, P3_U5188, P3_U5189);
  and ginst25205 (P3_U3804, P3_U5197, P3_U5198);
  and ginst25206 (P3_U3805, P3_U5203, P3_U5205);
  and ginst25207 (P3_U3806, P3_U5206, P3_U5207);
  and ginst25208 (P3_U3807, P3_U5215, P3_U5216);
  and ginst25209 (P3_U3808, P3_U5224, P3_U5225);
  and ginst25210 (P3_U3809, P3_U5233, P3_U5234);
  and ginst25211 (P3_U3810, P3_U5242, P3_U5243);
  and ginst25212 (P3_U3811, P3_U5251, P3_U5252);
  and ginst25213 (P3_U3812, P3_STATE_REG_SCAN_IN, P3_U5254);
  and ginst25214 (P3_U3813, P3_U3385, P3_U5440);
  and ginst25215 (P3_U3814, P3_U3375, P3_U3385);
  and ginst25216 (P3_U3815, P3_U3302, P3_U3312, P3_U3875);
  and ginst25217 (P3_U3816, P3_U3310, P3_U3357, P3_U3877);
  and ginst25218 (P3_U3817, P3_U3375, P3_U5258);
  and ginst25219 (P3_U3818, P3_U3375, P3_U5260);
  and ginst25220 (P3_U3819, P3_U3375, P3_U5262);
  and ginst25221 (P3_U3820, P3_U3375, P3_U5264);
  and ginst25222 (P3_U3821, P3_U3375, P3_U5266);
  and ginst25223 (P3_U3822, P3_U3375, P3_U5268);
  and ginst25224 (P3_U3823, P3_U3375, P3_U5274);
  and ginst25225 (P3_U3824, P3_U3375, P3_U5296);
  and ginst25226 (P3_U3825, P3_U3375, P3_U5310);
  and ginst25227 (P3_U3826, P3_U3375, P3_U5312);
  and ginst25228 (P3_U3827, P3_U3375, P3_U5314);
  and ginst25229 (P3_U3828, P3_U3375, P3_U5316);
  and ginst25230 (P3_U3829, P3_U3375, P3_U5318);
  and ginst25231 (P3_U3830, P3_U3375, P3_U5320);
  not ginst25232 (P3_U3831, P3_IR_REG_31__SCAN_IN);
  nand ginst25233 (P3_U3832, P3_U3023, P3_U3300);
  nand ginst25234 (P3_U3833, P3_U5465, P3_U5468);
  nand ginst25235 (P3_U3834, P3_U5447, P3_U5456);
  nand ginst25236 (P3_U3835, P3_U3023, P3_U4058);
  nand ginst25237 (P3_U3836, P3_U3023, P3_U4622);
  and ginst25238 (P3_U3837, P3_U5706, P3_U5707);
  and ginst25239 (P3_U3838, P3_U5708, P3_U5709);
  and ginst25240 (P3_U3839, P3_U5710, P3_U5711);
  and ginst25241 (P3_U3840, P3_U5712, P3_U5713);
  and ginst25242 (P3_U3841, P3_U5714, P3_U5715);
  and ginst25243 (P3_U3842, P3_U5716, P3_U5717);
  and ginst25244 (P3_U3843, P3_U5718, P3_U5719);
  and ginst25245 (P3_U3844, P3_U5720, P3_U5721);
  and ginst25246 (P3_U3845, P3_U5722, P3_U5723);
  and ginst25247 (P3_U3846, P3_U5724, P3_U5725);
  and ginst25248 (P3_U3847, P3_U5726, P3_U5727);
  and ginst25249 (P3_U3848, P3_U5728, P3_U5729);
  and ginst25250 (P3_U3849, P3_U5730, P3_U5731);
  and ginst25251 (P3_U3850, P3_U5732, P3_U5733);
  and ginst25252 (P3_U3851, P3_U5734, P3_U5735);
  and ginst25253 (P3_U3852, P3_U5736, P3_U5737);
  and ginst25254 (P3_U3853, P3_U5738, P3_U5739);
  and ginst25255 (P3_U3854, P3_U5740, P3_U5741);
  and ginst25256 (P3_U3855, P3_U5742, P3_U5743);
  and ginst25257 (P3_U3856, P3_U5744, P3_U5745);
  and ginst25258 (P3_U3857, P3_U5746, P3_U5747);
  and ginst25259 (P3_U3858, P3_U5748, P3_U5749);
  and ginst25260 (P3_U3859, P3_U5750, P3_U5751);
  and ginst25261 (P3_U3860, P3_U5752, P3_U5753);
  and ginst25262 (P3_U3861, P3_U5754, P3_U5755);
  and ginst25263 (P3_U3862, P3_U5756, P3_U5757);
  and ginst25264 (P3_U3863, P3_U5758, P3_U5759);
  and ginst25265 (P3_U3864, P3_U5760, P3_U5761);
  and ginst25266 (P3_U3865, P3_U5762, P3_U5763);
  and ginst25267 (P3_U3866, P3_U5764, P3_U5765);
  not ginst25268 (P3_U3867, P3_R1269_U11);
  nand ginst25269 (P3_U3868, P3_U3772, P3_U3773);
  not ginst25270 (P3_U3869, P3_R693_U14);
  and ginst25271 (P3_U3870, P3_U5939, P3_U5940);
  not ginst25272 (P3_U3871, P3_R1297_U6);
  not ginst25273 (P3_U3872, P3_U3356);
  not ginst25274 (P3_U3873, P3_U3355);
  not ginst25275 (P3_U3874, P3_U3312);
  nand ginst25276 (P3_U3875, P3_U3015, P3_U3385);
  not ginst25277 (P3_U3876, P3_U3302);
  nand ginst25278 (P3_U3877, P3_U3016, P3_U5456);
  not ginst25279 (P3_U3878, P3_U3310);
  not ginst25280 (P3_U3879, P3_U3357);
  nand ginst25281 (P3_U3880, P3_U3014, P3_U3385);
  not ginst25282 (P3_U3881, P3_U3308);
  not ginst25283 (P3_U3882, P3_U3301);
  not ginst25284 (P3_U3883, P3_U3305);
  not ginst25285 (P3_U3884, P3_U3307);
  not ginst25286 (P3_U3885, P3_U3306);
  not ginst25287 (P3_U3886, P3_U3360);
  not ginst25288 (P3_U3887, P3_U3311);
  nand ginst25289 (P3_U3888, P3_U3378, P3_U3878);
  not ginst25290 (P3_U3889, P3_U3369);
  not ginst25291 (P3_U3890, P3_U3367);
  not ginst25292 (P3_U3891, P3_U3309);
  not ginst25293 (P3_U3892, P3_U3352);
  not ginst25294 (P3_U3893, P3_U3833);
  not ginst25295 (P3_U3894, P3_U3303);
  not ginst25296 (P3_U3895, P3_U3304);
  nand ginst25297 (P3_U3896, P3_U3384, P3_U5465);
  not ginst25298 (P3_U3897, P3_U3363);
  not ginst25299 (P3_U3898, P3_U3364);
  not ginst25300 (P3_U3899, P3_U3350);
  not ginst25301 (P3_U3900, P3_U3348);
  not ginst25302 (P3_U3901, P3_U3346);
  not ginst25303 (P3_U3902, P3_U3344);
  not ginst25304 (P3_U3903, P3_U3342);
  not ginst25305 (P3_U3904, P3_U3340);
  not ginst25306 (P3_U3905, P3_U3338);
  not ginst25307 (P3_U3906, P3_U3336);
  not ginst25308 (P3_U3907, P3_U3334);
  not ginst25309 (P3_U3908, P3_U3353);
  not ginst25310 (P3_U3909, P3_U3368);
  not ginst25311 (P3_U3910, P3_U3362);
  not ginst25312 (P3_U3911, P3_U3313);
  not ginst25313 (P3_U3912, P3_U3358);
  not ginst25314 (P3_U3913, P3_U3836);
  not ginst25315 (P3_U3914, P3_U3835);
  not ginst25316 (P3_U3915, P3_U3832);
  not ginst25317 (P3_U3916, P3_U3361);
  nand ginst25318 (P3_U3917, P3_STATE_REG_SCAN_IN, P3_U3370);
  nand ginst25319 (P3_U3918, P3_U3023, P3_U3886);
  not ginst25320 (P3_U3919, P3_U3299);
  not ginst25321 (P3_U3920, P3_U3359);
  not ginst25322 (P3_U3921, P3_U3297);
  nand ginst25323 (P3_U3922, P3_U3151, U61);
  nand ginst25324 (P3_U3923, P3_IR_REG_0__SCAN_IN, P3_U3027);
  nand ginst25325 (P3_U3924, P3_IR_REG_0__SCAN_IN, P3_U3921);
  nand ginst25326 (P3_U3925, P3_U3151, U50);
  nand ginst25327 (P3_U3926, P3_SUB_598_U51, P3_U3027);
  nand ginst25328 (P3_U3927, P3_IR_REG_1__SCAN_IN, P3_U3921);
  nand ginst25329 (P3_U3928, P3_U3151, U39);
  nand ginst25330 (P3_U3929, P3_SUB_598_U22, P3_U3027);
  nand ginst25331 (P3_U3930, P3_IR_REG_2__SCAN_IN, P3_U3921);
  nand ginst25332 (P3_U3931, P3_U3151, U36);
  nand ginst25333 (P3_U3932, P3_SUB_598_U23, P3_U3027);
  nand ginst25334 (P3_U3933, P3_IR_REG_3__SCAN_IN, P3_U3921);
  nand ginst25335 (P3_U3934, P3_U3151, U35);
  nand ginst25336 (P3_U3935, P3_SUB_598_U24, P3_U3027);
  nand ginst25337 (P3_U3936, P3_IR_REG_4__SCAN_IN, P3_U3921);
  nand ginst25338 (P3_U3937, P3_U3151, U34);
  nand ginst25339 (P3_U3938, P3_SUB_598_U74, P3_U3027);
  nand ginst25340 (P3_U3939, P3_IR_REG_5__SCAN_IN, P3_U3921);
  nand ginst25341 (P3_U3940, P3_U3151, U33);
  nand ginst25342 (P3_U3941, P3_SUB_598_U25, P3_U3027);
  nand ginst25343 (P3_U3942, P3_IR_REG_6__SCAN_IN, P3_U3921);
  nand ginst25344 (P3_U3943, P3_U3151, U32);
  nand ginst25345 (P3_U3944, P3_SUB_598_U26, P3_U3027);
  nand ginst25346 (P3_U3945, P3_IR_REG_7__SCAN_IN, P3_U3921);
  nand ginst25347 (P3_U3946, P3_U3151, U31);
  nand ginst25348 (P3_U3947, P3_SUB_598_U27, P3_U3027);
  nand ginst25349 (P3_U3948, P3_IR_REG_8__SCAN_IN, P3_U3921);
  nand ginst25350 (P3_U3949, P3_U3151, U30);
  nand ginst25351 (P3_U3950, P3_SUB_598_U72, P3_U3027);
  nand ginst25352 (P3_U3951, P3_IR_REG_9__SCAN_IN, P3_U3921);
  nand ginst25353 (P3_U3952, P3_U3151, U60);
  nand ginst25354 (P3_U3953, P3_SUB_598_U7, P3_U3027);
  nand ginst25355 (P3_U3954, P3_IR_REG_10__SCAN_IN, P3_U3921);
  nand ginst25356 (P3_U3955, P3_U3151, U59);
  nand ginst25357 (P3_U3956, P3_SUB_598_U8, P3_U3027);
  nand ginst25358 (P3_U3957, P3_IR_REG_11__SCAN_IN, P3_U3921);
  nand ginst25359 (P3_U3958, P3_U3151, U58);
  nand ginst25360 (P3_U3959, P3_SUB_598_U9, P3_U3027);
  nand ginst25361 (P3_U3960, P3_IR_REG_12__SCAN_IN, P3_U3921);
  nand ginst25362 (P3_U3961, P3_U3151, U57);
  nand ginst25363 (P3_U3962, P3_SUB_598_U89, P3_U3027);
  nand ginst25364 (P3_U3963, P3_IR_REG_13__SCAN_IN, P3_U3921);
  nand ginst25365 (P3_U3964, P3_U3151, U56);
  nand ginst25366 (P3_U3965, P3_SUB_598_U10, P3_U3027);
  nand ginst25367 (P3_U3966, P3_IR_REG_14__SCAN_IN, P3_U3921);
  nand ginst25368 (P3_U3967, P3_U3151, U55);
  nand ginst25369 (P3_U3968, P3_SUB_598_U11, P3_U3027);
  nand ginst25370 (P3_U3969, P3_IR_REG_15__SCAN_IN, P3_U3921);
  nand ginst25371 (P3_U3970, P3_U3151, U54);
  nand ginst25372 (P3_U3971, P3_SUB_598_U12, P3_U3027);
  nand ginst25373 (P3_U3972, P3_IR_REG_16__SCAN_IN, P3_U3921);
  nand ginst25374 (P3_U3973, P3_U3151, U53);
  nand ginst25375 (P3_U3974, P3_SUB_598_U87, P3_U3027);
  nand ginst25376 (P3_U3975, P3_IR_REG_17__SCAN_IN, P3_U3921);
  nand ginst25377 (P3_U3976, P3_U3151, U52);
  nand ginst25378 (P3_U3977, P3_SUB_598_U13, P3_U3027);
  nand ginst25379 (P3_U3978, P3_IR_REG_18__SCAN_IN, P3_U3921);
  nand ginst25380 (P3_U3979, P3_U3151, U51);
  nand ginst25381 (P3_U3980, P3_SUB_598_U14, P3_U3027);
  nand ginst25382 (P3_U3981, P3_IR_REG_19__SCAN_IN, P3_U3921);
  nand ginst25383 (P3_U3982, P3_U3151, U49);
  nand ginst25384 (P3_U3983, P3_SUB_598_U15, P3_U3027);
  nand ginst25385 (P3_U3984, P3_IR_REG_20__SCAN_IN, P3_U3921);
  nand ginst25386 (P3_U3985, P3_U3151, U48);
  nand ginst25387 (P3_U3986, P3_SUB_598_U83, P3_U3027);
  nand ginst25388 (P3_U3987, P3_IR_REG_21__SCAN_IN, P3_U3921);
  nand ginst25389 (P3_U3988, P3_U3151, U47);
  nand ginst25390 (P3_U3989, P3_SUB_598_U16, P3_U3027);
  nand ginst25391 (P3_U3990, P3_IR_REG_22__SCAN_IN, P3_U3921);
  nand ginst25392 (P3_U3991, P3_U3151, U46);
  nand ginst25393 (P3_U3992, P3_SUB_598_U17, P3_U3027);
  nand ginst25394 (P3_U3993, P3_IR_REG_23__SCAN_IN, P3_U3921);
  nand ginst25395 (P3_U3994, P3_U3151, U45);
  nand ginst25396 (P3_U3995, P3_SUB_598_U18, P3_U3027);
  nand ginst25397 (P3_U3996, P3_IR_REG_24__SCAN_IN, P3_U3921);
  nand ginst25398 (P3_U3997, P3_U3151, U44);
  nand ginst25399 (P3_U3998, P3_SUB_598_U81, P3_U3027);
  nand ginst25400 (P3_U3999, P3_IR_REG_25__SCAN_IN, P3_U3921);
  nand ginst25401 (P3_U4000, P3_U3151, U43);
  nand ginst25402 (P3_U4001, P3_SUB_598_U19, P3_U3027);
  nand ginst25403 (P3_U4002, P3_IR_REG_26__SCAN_IN, P3_U3921);
  nand ginst25404 (P3_U4003, P3_U3151, U42);
  nand ginst25405 (P3_U4004, P3_SUB_598_U79, P3_U3027);
  nand ginst25406 (P3_U4005, P3_IR_REG_27__SCAN_IN, P3_U3921);
  nand ginst25407 (P3_U4006, P3_U3151, U41);
  nand ginst25408 (P3_U4007, P3_SUB_598_U20, P3_U3027);
  nand ginst25409 (P3_U4008, P3_IR_REG_28__SCAN_IN, P3_U3921);
  nand ginst25410 (P3_U4009, P3_U3151, U40);
  nand ginst25411 (P3_U4010, P3_SUB_598_U21, P3_U3027);
  nand ginst25412 (P3_U4011, P3_IR_REG_29__SCAN_IN, P3_U3921);
  nand ginst25413 (P3_U4012, P3_U3151, U38);
  nand ginst25414 (P3_U4013, P3_SUB_598_U77, P3_U3027);
  nand ginst25415 (P3_U4014, P3_IR_REG_30__SCAN_IN, P3_U3921);
  nand ginst25416 (P3_U4015, P3_U3151, U37);
  nand ginst25417 (P3_U4016, P3_SUB_598_U52, P3_U3027);
  nand ginst25418 (P3_U4017, P3_IR_REG_31__SCAN_IN, P3_U3921);
  nand ginst25419 (P3_U4018, P3_U3919, P3_U5437);
  not ginst25420 (P3_U4019, P3_U3300);
  nand ginst25421 (P3_U4020, P3_U3299, P3_U5428);
  nand ginst25422 (P3_U4021, P3_U3299, P3_U5431);
  nand ginst25423 (P3_U4022, P3_D_REG_10__SCAN_IN, P3_U4019);
  nand ginst25424 (P3_U4023, P3_D_REG_11__SCAN_IN, P3_U4019);
  nand ginst25425 (P3_U4024, P3_D_REG_12__SCAN_IN, P3_U4019);
  nand ginst25426 (P3_U4025, P3_D_REG_13__SCAN_IN, P3_U4019);
  nand ginst25427 (P3_U4026, P3_D_REG_14__SCAN_IN, P3_U4019);
  nand ginst25428 (P3_U4027, P3_D_REG_15__SCAN_IN, P3_U4019);
  nand ginst25429 (P3_U4028, P3_D_REG_16__SCAN_IN, P3_U4019);
  nand ginst25430 (P3_U4029, P3_D_REG_17__SCAN_IN, P3_U4019);
  nand ginst25431 (P3_U4030, P3_D_REG_18__SCAN_IN, P3_U4019);
  nand ginst25432 (P3_U4031, P3_D_REG_19__SCAN_IN, P3_U4019);
  nand ginst25433 (P3_U4032, P3_D_REG_20__SCAN_IN, P3_U4019);
  nand ginst25434 (P3_U4033, P3_D_REG_21__SCAN_IN, P3_U4019);
  nand ginst25435 (P3_U4034, P3_D_REG_22__SCAN_IN, P3_U4019);
  nand ginst25436 (P3_U4035, P3_D_REG_23__SCAN_IN, P3_U4019);
  nand ginst25437 (P3_U4036, P3_D_REG_24__SCAN_IN, P3_U4019);
  nand ginst25438 (P3_U4037, P3_D_REG_25__SCAN_IN, P3_U4019);
  nand ginst25439 (P3_U4038, P3_D_REG_26__SCAN_IN, P3_U4019);
  nand ginst25440 (P3_U4039, P3_D_REG_27__SCAN_IN, P3_U4019);
  nand ginst25441 (P3_U4040, P3_D_REG_28__SCAN_IN, P3_U4019);
  nand ginst25442 (P3_U4041, P3_D_REG_29__SCAN_IN, P3_U4019);
  nand ginst25443 (P3_U4042, P3_D_REG_2__SCAN_IN, P3_U4019);
  nand ginst25444 (P3_U4043, P3_D_REG_30__SCAN_IN, P3_U4019);
  nand ginst25445 (P3_U4044, P3_D_REG_31__SCAN_IN, P3_U4019);
  nand ginst25446 (P3_U4045, P3_D_REG_3__SCAN_IN, P3_U4019);
  nand ginst25447 (P3_U4046, P3_D_REG_4__SCAN_IN, P3_U4019);
  nand ginst25448 (P3_U4047, P3_D_REG_5__SCAN_IN, P3_U4019);
  nand ginst25449 (P3_U4048, P3_D_REG_6__SCAN_IN, P3_U4019);
  nand ginst25450 (P3_U4049, P3_D_REG_7__SCAN_IN, P3_U4019);
  nand ginst25451 (P3_U4050, P3_D_REG_8__SCAN_IN, P3_U4019);
  nand ginst25452 (P3_U4051, P3_D_REG_9__SCAN_IN, P3_U4019);
  not ginst25453 (P3_U4052, P3_U3834);
  nand ginst25454 (P3_U4053, P3_U5450, P3_U5456);
  nand ginst25455 (P3_U4054, P3_U4053, P3_U5482);
  nand ginst25456 (P3_U4055, P3_U3367, P3_U3369);
  nand ginst25457 (P3_U4056, P3_U3894, P3_U4055);
  nand ginst25458 (P3_U4057, P3_U3895, P3_U4054);
  nand ginst25459 (P3_U4058, P3_U4056, P3_U4057);
  nand ginst25460 (P3_U4059, P3_REG0_REG_1__SCAN_IN, P3_U3022);
  nand ginst25461 (P3_U4060, P3_REG1_REG_1__SCAN_IN, P3_U3021);
  nand ginst25462 (P3_U4061, P3_REG2_REG_1__SCAN_IN, P3_U3020);
  nand ginst25463 (P3_U4062, P3_REG3_REG_1__SCAN_IN, P3_U3019);
  not ginst25464 (P3_U4063, P3_U3077);
  nand ginst25465 (P3_U4064, P3_U3357, P3_U3877);
  nand ginst25466 (P3_U4065, P3_R1110_U95, P3_U3883);
  nand ginst25467 (P3_U4066, P3_R1077_U95, P3_U3885);
  nand ginst25468 (P3_U4067, P3_R1095_U24, P3_U3884);
  nand ginst25469 (P3_U4068, P3_R1143_U95, P3_U3881);
  nand ginst25470 (P3_U4069, P3_R1161_U95, P3_U3891);
  nand ginst25471 (P3_U4070, P3_R1131_U24, P3_U3887);
  nand ginst25472 (P3_U4071, P3_R1200_U24, P3_U3017);
  not ginst25473 (P3_U4072, P3_U3314);
  nand ginst25474 (P3_U4073, P3_U3352, P3_U3833);
  nand ginst25475 (P3_U4074, P3_R1179_U24, P3_U3026);
  nand ginst25476 (P3_U4075, P3_U3025, P3_U3077);
  nand ginst25477 (P3_U4076, P3_U3387, P3_U4064);
  nand ginst25478 (P3_U4077, P3_U3577, P3_U4072);
  nand ginst25479 (P3_U4078, P3_REG0_REG_2__SCAN_IN, P3_U3022);
  nand ginst25480 (P3_U4079, P3_REG1_REG_2__SCAN_IN, P3_U3021);
  nand ginst25481 (P3_U4080, P3_REG2_REG_2__SCAN_IN, P3_U3020);
  nand ginst25482 (P3_U4081, P3_REG3_REG_2__SCAN_IN, P3_U3019);
  not ginst25483 (P3_U4082, P3_U3067);
  nand ginst25484 (P3_U4083, P3_REG0_REG_0__SCAN_IN, P3_U3022);
  nand ginst25485 (P3_U4084, P3_REG1_REG_0__SCAN_IN, P3_U3021);
  nand ginst25486 (P3_U4085, P3_REG2_REG_0__SCAN_IN, P3_U3020);
  nand ginst25487 (P3_U4086, P3_REG3_REG_0__SCAN_IN, P3_U3019);
  not ginst25488 (P3_U4087, P3_U3076);
  nand ginst25489 (P3_U4088, P3_U3383, P3_U5468);
  nand ginst25490 (P3_U4089, P3_U3896, P3_U4088);
  nand ginst25491 (P3_U4090, P3_U3033, P3_U3076);
  nand ginst25492 (P3_U4091, P3_R1110_U94, P3_U3883);
  nand ginst25493 (P3_U4092, P3_R1077_U94, P3_U3885);
  nand ginst25494 (P3_U4093, P3_R1095_U100, P3_U3884);
  nand ginst25495 (P3_U4094, P3_R1143_U94, P3_U3881);
  nand ginst25496 (P3_U4095, P3_R1161_U94, P3_U3891);
  nand ginst25497 (P3_U4096, P3_R1131_U100, P3_U3887);
  nand ginst25498 (P3_U4097, P3_R1200_U100, P3_U3017);
  not ginst25499 (P3_U4098, P3_U3315);
  nand ginst25500 (P3_U4099, P3_R1179_U100, P3_U3026);
  nand ginst25501 (P3_U4100, P3_U3025, P3_U3067);
  nand ginst25502 (P3_U4101, P3_U3392, P3_U4064);
  nand ginst25503 (P3_U4102, P3_U3593, P3_U4098);
  nand ginst25504 (P3_U4103, P3_REG0_REG_3__SCAN_IN, P3_U3022);
  nand ginst25505 (P3_U4104, P3_REG1_REG_3__SCAN_IN, P3_U3021);
  nand ginst25506 (P3_U4105, P3_REG2_REG_3__SCAN_IN, P3_U3020);
  nand ginst25507 (P3_U4106, P3_SUB_609_U25, P3_U3019);
  not ginst25508 (P3_U4107, P3_U3063);
  nand ginst25509 (P3_U4108, P3_U3033, P3_U3077);
  nand ginst25510 (P3_U4109, P3_R1110_U16, P3_U3883);
  nand ginst25511 (P3_U4110, P3_R1077_U16, P3_U3885);
  nand ginst25512 (P3_U4111, P3_R1095_U110, P3_U3884);
  nand ginst25513 (P3_U4112, P3_R1143_U16, P3_U3881);
  nand ginst25514 (P3_U4113, P3_R1161_U16, P3_U3891);
  nand ginst25515 (P3_U4114, P3_R1131_U110, P3_U3887);
  nand ginst25516 (P3_U4115, P3_R1200_U110, P3_U3017);
  not ginst25517 (P3_U4116, P3_U3316);
  nand ginst25518 (P3_U4117, P3_R1179_U110, P3_U3026);
  nand ginst25519 (P3_U4118, P3_U3025, P3_U3063);
  nand ginst25520 (P3_U4119, P3_U3395, P3_U4064);
  nand ginst25521 (P3_U4120, P3_U3597, P3_U4116);
  nand ginst25522 (P3_U4121, P3_REG0_REG_4__SCAN_IN, P3_U3022);
  nand ginst25523 (P3_U4122, P3_REG1_REG_4__SCAN_IN, P3_U3021);
  nand ginst25524 (P3_U4123, P3_REG2_REG_4__SCAN_IN, P3_U3020);
  nand ginst25525 (P3_U4124, P3_SUB_609_U29, P3_U3019);
  not ginst25526 (P3_U4125, P3_U3059);
  nand ginst25527 (P3_U4126, P3_U3033, P3_U3067);
  nand ginst25528 (P3_U4127, P3_R1110_U100, P3_U3883);
  nand ginst25529 (P3_U4128, P3_R1077_U100, P3_U3885);
  nand ginst25530 (P3_U4129, P3_R1095_U21, P3_U3884);
  nand ginst25531 (P3_U4130, P3_R1143_U100, P3_U3881);
  nand ginst25532 (P3_U4131, P3_R1161_U100, P3_U3891);
  nand ginst25533 (P3_U4132, P3_R1131_U21, P3_U3887);
  nand ginst25534 (P3_U4133, P3_R1200_U21, P3_U3017);
  not ginst25535 (P3_U4134, P3_U3317);
  nand ginst25536 (P3_U4135, P3_R1179_U21, P3_U3026);
  nand ginst25537 (P3_U4136, P3_U3025, P3_U3059);
  nand ginst25538 (P3_U4137, P3_U3398, P3_U4064);
  nand ginst25539 (P3_U4138, P3_U3601, P3_U4134);
  nand ginst25540 (P3_U4139, P3_REG0_REG_5__SCAN_IN, P3_U3022);
  nand ginst25541 (P3_U4140, P3_REG1_REG_5__SCAN_IN, P3_U3021);
  nand ginst25542 (P3_U4141, P3_REG2_REG_5__SCAN_IN, P3_U3020);
  nand ginst25543 (P3_U4142, P3_SUB_609_U53, P3_U3019);
  not ginst25544 (P3_U4143, P3_U3066);
  nand ginst25545 (P3_U4144, P3_U3033, P3_U3063);
  nand ginst25546 (P3_U4145, P3_R1110_U99, P3_U3883);
  nand ginst25547 (P3_U4146, P3_R1077_U99, P3_U3885);
  nand ginst25548 (P3_U4147, P3_R1095_U109, P3_U3884);
  nand ginst25549 (P3_U4148, P3_R1143_U99, P3_U3881);
  nand ginst25550 (P3_U4149, P3_R1161_U99, P3_U3891);
  nand ginst25551 (P3_U4150, P3_R1131_U109, P3_U3887);
  nand ginst25552 (P3_U4151, P3_R1200_U109, P3_U3017);
  not ginst25553 (P3_U4152, P3_U3318);
  nand ginst25554 (P3_U4153, P3_R1179_U109, P3_U3026);
  nand ginst25555 (P3_U4154, P3_U3025, P3_U3066);
  nand ginst25556 (P3_U4155, P3_U3401, P3_U4064);
  nand ginst25557 (P3_U4156, P3_U3604, P3_U4152);
  nand ginst25558 (P3_U4157, P3_REG0_REG_6__SCAN_IN, P3_U3022);
  nand ginst25559 (P3_U4158, P3_REG1_REG_6__SCAN_IN, P3_U3021);
  nand ginst25560 (P3_U4159, P3_REG2_REG_6__SCAN_IN, P3_U3020);
  nand ginst25561 (P3_U4160, P3_SUB_609_U8, P3_U3019);
  not ginst25562 (P3_U4161, P3_U3070);
  nand ginst25563 (P3_U4162, P3_U3033, P3_U3059);
  nand ginst25564 (P3_U4163, P3_R1110_U17, P3_U3883);
  nand ginst25565 (P3_U4164, P3_R1077_U17, P3_U3885);
  nand ginst25566 (P3_U4165, P3_R1095_U108, P3_U3884);
  nand ginst25567 (P3_U4166, P3_R1143_U17, P3_U3881);
  nand ginst25568 (P3_U4167, P3_R1161_U17, P3_U3891);
  nand ginst25569 (P3_U4168, P3_R1131_U108, P3_U3887);
  nand ginst25570 (P3_U4169, P3_R1200_U108, P3_U3017);
  not ginst25571 (P3_U4170, P3_U3319);
  nand ginst25572 (P3_U4171, P3_R1179_U108, P3_U3026);
  nand ginst25573 (P3_U4172, P3_U3025, P3_U3070);
  nand ginst25574 (P3_U4173, P3_U3404, P3_U4064);
  nand ginst25575 (P3_U4174, P3_U3607, P3_U4170);
  nand ginst25576 (P3_U4175, P3_REG0_REG_7__SCAN_IN, P3_U3022);
  nand ginst25577 (P3_U4176, P3_REG1_REG_7__SCAN_IN, P3_U3021);
  nand ginst25578 (P3_U4177, P3_REG2_REG_7__SCAN_IN, P3_U3020);
  nand ginst25579 (P3_U4178, P3_SUB_609_U18, P3_U3019);
  not ginst25580 (P3_U4179, P3_U3069);
  nand ginst25581 (P3_U4180, P3_U3033, P3_U3066);
  nand ginst25582 (P3_U4181, P3_R1110_U98, P3_U3883);
  nand ginst25583 (P3_U4182, P3_R1077_U98, P3_U3885);
  nand ginst25584 (P3_U4183, P3_R1095_U22, P3_U3884);
  nand ginst25585 (P3_U4184, P3_R1143_U98, P3_U3881);
  nand ginst25586 (P3_U4185, P3_R1161_U98, P3_U3891);
  nand ginst25587 (P3_U4186, P3_R1131_U22, P3_U3887);
  nand ginst25588 (P3_U4187, P3_R1200_U22, P3_U3017);
  not ginst25589 (P3_U4188, P3_U3320);
  nand ginst25590 (P3_U4189, P3_R1179_U22, P3_U3026);
  nand ginst25591 (P3_U4190, P3_U3025, P3_U3069);
  nand ginst25592 (P3_U4191, P3_U3407, P3_U4064);
  nand ginst25593 (P3_U4192, P3_U3610, P3_U4188);
  nand ginst25594 (P3_U4193, P3_REG0_REG_8__SCAN_IN, P3_U3022);
  nand ginst25595 (P3_U4194, P3_REG1_REG_8__SCAN_IN, P3_U3021);
  nand ginst25596 (P3_U4195, P3_REG2_REG_8__SCAN_IN, P3_U3020);
  nand ginst25597 (P3_U4196, P3_SUB_609_U12, P3_U3019);
  not ginst25598 (P3_U4197, P3_U3083);
  nand ginst25599 (P3_U4198, P3_U3033, P3_U3070);
  nand ginst25600 (P3_U4199, P3_R1110_U18, P3_U3883);
  nand ginst25601 (P3_U4200, P3_R1077_U18, P3_U3885);
  nand ginst25602 (P3_U4201, P3_R1095_U107, P3_U3884);
  nand ginst25603 (P3_U4202, P3_R1143_U18, P3_U3881);
  nand ginst25604 (P3_U4203, P3_R1161_U18, P3_U3891);
  nand ginst25605 (P3_U4204, P3_R1131_U107, P3_U3887);
  nand ginst25606 (P3_U4205, P3_R1200_U107, P3_U3017);
  not ginst25607 (P3_U4206, P3_U3321);
  nand ginst25608 (P3_U4207, P3_R1179_U107, P3_U3026);
  nand ginst25609 (P3_U4208, P3_U3025, P3_U3083);
  nand ginst25610 (P3_U4209, P3_U3410, P3_U4064);
  nand ginst25611 (P3_U4210, P3_U3613, P3_U4206);
  nand ginst25612 (P3_U4211, P3_REG0_REG_9__SCAN_IN, P3_U3022);
  nand ginst25613 (P3_U4212, P3_REG1_REG_9__SCAN_IN, P3_U3021);
  nand ginst25614 (P3_U4213, P3_REG2_REG_9__SCAN_IN, P3_U3020);
  nand ginst25615 (P3_U4214, P3_SUB_609_U14, P3_U3019);
  not ginst25616 (P3_U4215, P3_U3082);
  nand ginst25617 (P3_U4216, P3_U3033, P3_U3069);
  nand ginst25618 (P3_U4217, P3_R1110_U97, P3_U3883);
  nand ginst25619 (P3_U4218, P3_R1077_U97, P3_U3885);
  nand ginst25620 (P3_U4219, P3_R1095_U23, P3_U3884);
  nand ginst25621 (P3_U4220, P3_R1143_U97, P3_U3881);
  nand ginst25622 (P3_U4221, P3_R1161_U97, P3_U3891);
  nand ginst25623 (P3_U4222, P3_R1131_U23, P3_U3887);
  nand ginst25624 (P3_U4223, P3_R1200_U23, P3_U3017);
  not ginst25625 (P3_U4224, P3_U3322);
  nand ginst25626 (P3_U4225, P3_R1179_U23, P3_U3026);
  nand ginst25627 (P3_U4226, P3_U3025, P3_U3082);
  nand ginst25628 (P3_U4227, P3_U3413, P3_U4064);
  nand ginst25629 (P3_U4228, P3_U3616, P3_U4224);
  nand ginst25630 (P3_U4229, P3_REG0_REG_10__SCAN_IN, P3_U3022);
  nand ginst25631 (P3_U4230, P3_REG1_REG_10__SCAN_IN, P3_U3021);
  nand ginst25632 (P3_U4231, P3_REG2_REG_10__SCAN_IN, P3_U3020);
  nand ginst25633 (P3_U4232, P3_SUB_609_U13, P3_U3019);
  not ginst25634 (P3_U4233, P3_U3061);
  nand ginst25635 (P3_U4234, P3_U3033, P3_U3083);
  nand ginst25636 (P3_U4235, P3_R1110_U96, P3_U3883);
  nand ginst25637 (P3_U4236, P3_R1077_U96, P3_U3885);
  nand ginst25638 (P3_U4237, P3_R1095_U106, P3_U3884);
  nand ginst25639 (P3_U4238, P3_R1143_U96, P3_U3881);
  nand ginst25640 (P3_U4239, P3_R1161_U96, P3_U3891);
  nand ginst25641 (P3_U4240, P3_R1131_U106, P3_U3887);
  nand ginst25642 (P3_U4241, P3_R1200_U106, P3_U3017);
  not ginst25643 (P3_U4242, P3_U3323);
  nand ginst25644 (P3_U4243, P3_R1179_U106, P3_U3026);
  nand ginst25645 (P3_U4244, P3_U3025, P3_U3061);
  nand ginst25646 (P3_U4245, P3_U3416, P3_U4064);
  nand ginst25647 (P3_U4246, P3_U3620, P3_U4242);
  nand ginst25648 (P3_U4247, P3_REG0_REG_11__SCAN_IN, P3_U3022);
  nand ginst25649 (P3_U4248, P3_REG1_REG_11__SCAN_IN, P3_U3021);
  nand ginst25650 (P3_U4249, P3_REG2_REG_11__SCAN_IN, P3_U3020);
  nand ginst25651 (P3_U4250, P3_SUB_609_U9, P3_U3019);
  not ginst25652 (P3_U4251, P3_U3062);
  nand ginst25653 (P3_U4252, P3_U3033, P3_U3082);
  nand ginst25654 (P3_U4253, P3_R1110_U10, P3_U3883);
  nand ginst25655 (P3_U4254, P3_R1077_U10, P3_U3885);
  nand ginst25656 (P3_U4255, P3_R1095_U116, P3_U3884);
  nand ginst25657 (P3_U4256, P3_R1143_U10, P3_U3881);
  nand ginst25658 (P3_U4257, P3_R1161_U10, P3_U3891);
  nand ginst25659 (P3_U4258, P3_R1131_U116, P3_U3887);
  nand ginst25660 (P3_U4259, P3_R1200_U116, P3_U3017);
  not ginst25661 (P3_U4260, P3_U3324);
  nand ginst25662 (P3_U4261, P3_R1179_U116, P3_U3026);
  nand ginst25663 (P3_U4262, P3_U3025, P3_U3062);
  nand ginst25664 (P3_U4263, P3_U3419, P3_U4064);
  nand ginst25665 (P3_U4264, P3_U3624, P3_U4260);
  nand ginst25666 (P3_U4265, P3_REG0_REG_12__SCAN_IN, P3_U3022);
  nand ginst25667 (P3_U4266, P3_REG1_REG_12__SCAN_IN, P3_U3021);
  nand ginst25668 (P3_U4267, P3_REG2_REG_12__SCAN_IN, P3_U3020);
  nand ginst25669 (P3_U4268, P3_SUB_609_U23, P3_U3019);
  not ginst25670 (P3_U4269, P3_U3071);
  nand ginst25671 (P3_U4270, P3_U3033, P3_U3061);
  nand ginst25672 (P3_U4271, P3_R1110_U114, P3_U3883);
  nand ginst25673 (P3_U4272, P3_R1077_U114, P3_U3885);
  nand ginst25674 (P3_U4273, P3_R1095_U16, P3_U3884);
  nand ginst25675 (P3_U4274, P3_R1143_U114, P3_U3881);
  nand ginst25676 (P3_U4275, P3_R1161_U114, P3_U3891);
  nand ginst25677 (P3_U4276, P3_R1131_U16, P3_U3887);
  nand ginst25678 (P3_U4277, P3_R1200_U16, P3_U3017);
  not ginst25679 (P3_U4278, P3_U3325);
  nand ginst25680 (P3_U4279, P3_R1179_U16, P3_U3026);
  nand ginst25681 (P3_U4280, P3_U3025, P3_U3071);
  nand ginst25682 (P3_U4281, P3_U3422, P3_U4064);
  nand ginst25683 (P3_U4282, P3_U3627, P3_U4278);
  nand ginst25684 (P3_U4283, P3_REG0_REG_13__SCAN_IN, P3_U3022);
  nand ginst25685 (P3_U4284, P3_REG1_REG_13__SCAN_IN, P3_U3021);
  nand ginst25686 (P3_U4285, P3_REG2_REG_13__SCAN_IN, P3_U3020);
  nand ginst25687 (P3_U4286, P3_SUB_609_U24, P3_U3019);
  not ginst25688 (P3_U4287, P3_U3079);
  nand ginst25689 (P3_U4288, P3_U3033, P3_U3062);
  nand ginst25690 (P3_U4289, P3_R1110_U113, P3_U3883);
  nand ginst25691 (P3_U4290, P3_R1077_U113, P3_U3885);
  nand ginst25692 (P3_U4291, P3_R1095_U105, P3_U3884);
  nand ginst25693 (P3_U4292, P3_R1143_U113, P3_U3881);
  nand ginst25694 (P3_U4293, P3_R1161_U113, P3_U3891);
  nand ginst25695 (P3_U4294, P3_R1131_U105, P3_U3887);
  nand ginst25696 (P3_U4295, P3_R1200_U105, P3_U3017);
  not ginst25697 (P3_U4296, P3_U3326);
  nand ginst25698 (P3_U4297, P3_R1179_U105, P3_U3026);
  nand ginst25699 (P3_U4298, P3_U3025, P3_U3079);
  nand ginst25700 (P3_U4299, P3_U3425, P3_U4064);
  nand ginst25701 (P3_U4300, P3_U3631, P3_U4296);
  nand ginst25702 (P3_U4301, P3_REG0_REG_14__SCAN_IN, P3_U3022);
  nand ginst25703 (P3_U4302, P3_REG1_REG_14__SCAN_IN, P3_U3021);
  nand ginst25704 (P3_U4303, P3_REG2_REG_14__SCAN_IN, P3_U3020);
  nand ginst25705 (P3_U4304, P3_SUB_609_U30, P3_U3019);
  not ginst25706 (P3_U4305, P3_U3078);
  nand ginst25707 (P3_U4306, P3_U3033, P3_U3071);
  nand ginst25708 (P3_U4307, P3_R1110_U11, P3_U3883);
  nand ginst25709 (P3_U4308, P3_R1077_U11, P3_U3885);
  nand ginst25710 (P3_U4309, P3_R1095_U104, P3_U3884);
  nand ginst25711 (P3_U4310, P3_R1143_U11, P3_U3881);
  nand ginst25712 (P3_U4311, P3_R1161_U11, P3_U3891);
  nand ginst25713 (P3_U4312, P3_R1131_U104, P3_U3887);
  nand ginst25714 (P3_U4313, P3_R1200_U104, P3_U3017);
  not ginst25715 (P3_U4314, P3_U3327);
  nand ginst25716 (P3_U4315, P3_R1179_U104, P3_U3026);
  nand ginst25717 (P3_U4316, P3_U3025, P3_U3078);
  nand ginst25718 (P3_U4317, P3_U3428, P3_U4064);
  nand ginst25719 (P3_U4318, P3_U3635, P3_U4314);
  nand ginst25720 (P3_U4319, P3_REG0_REG_15__SCAN_IN, P3_U3022);
  nand ginst25721 (P3_U4320, P3_REG1_REG_15__SCAN_IN, P3_U3021);
  nand ginst25722 (P3_U4321, P3_REG2_REG_15__SCAN_IN, P3_U3020);
  nand ginst25723 (P3_U4322, P3_SUB_609_U21, P3_U3019);
  not ginst25724 (P3_U4323, P3_U3073);
  nand ginst25725 (P3_U4324, P3_U3033, P3_U3079);
  nand ginst25726 (P3_U4325, P3_R1110_U112, P3_U3883);
  nand ginst25727 (P3_U4326, P3_R1077_U112, P3_U3885);
  nand ginst25728 (P3_U4327, P3_R1095_U115, P3_U3884);
  nand ginst25729 (P3_U4328, P3_R1143_U112, P3_U3881);
  nand ginst25730 (P3_U4329, P3_R1161_U112, P3_U3891);
  nand ginst25731 (P3_U4330, P3_R1131_U115, P3_U3887);
  nand ginst25732 (P3_U4331, P3_R1200_U115, P3_U3017);
  not ginst25733 (P3_U4332, P3_U3328);
  nand ginst25734 (P3_U4333, P3_R1179_U115, P3_U3026);
  nand ginst25735 (P3_U4334, P3_U3025, P3_U3073);
  nand ginst25736 (P3_U4335, P3_U3431, P3_U4064);
  nand ginst25737 (P3_U4336, P3_U3638, P3_U4332);
  nand ginst25738 (P3_U4337, P3_REG0_REG_16__SCAN_IN, P3_U3022);
  nand ginst25739 (P3_U4338, P3_REG1_REG_16__SCAN_IN, P3_U3021);
  nand ginst25740 (P3_U4339, P3_REG2_REG_16__SCAN_IN, P3_U3020);
  nand ginst25741 (P3_U4340, P3_SUB_609_U7, P3_U3019);
  not ginst25742 (P3_U4341, P3_U3072);
  nand ginst25743 (P3_U4342, P3_U3033, P3_U3078);
  nand ginst25744 (P3_U4343, P3_R1110_U111, P3_U3883);
  nand ginst25745 (P3_U4344, P3_R1077_U111, P3_U3885);
  nand ginst25746 (P3_U4345, P3_R1095_U114, P3_U3884);
  nand ginst25747 (P3_U4346, P3_R1143_U111, P3_U3881);
  nand ginst25748 (P3_U4347, P3_R1161_U111, P3_U3891);
  nand ginst25749 (P3_U4348, P3_R1131_U114, P3_U3887);
  nand ginst25750 (P3_U4349, P3_R1200_U114, P3_U3017);
  not ginst25751 (P3_U4350, P3_U3329);
  nand ginst25752 (P3_U4351, P3_R1179_U114, P3_U3026);
  nand ginst25753 (P3_U4352, P3_U3025, P3_U3072);
  nand ginst25754 (P3_U4353, P3_U3434, P3_U4064);
  nand ginst25755 (P3_U4354, P3_U3641, P3_U4350);
  nand ginst25756 (P3_U4355, P3_REG0_REG_17__SCAN_IN, P3_U3022);
  nand ginst25757 (P3_U4356, P3_REG1_REG_17__SCAN_IN, P3_U3021);
  nand ginst25758 (P3_U4357, P3_REG2_REG_17__SCAN_IN, P3_U3020);
  nand ginst25759 (P3_U4358, P3_SUB_609_U19, P3_U3019);
  not ginst25760 (P3_U4359, P3_U3068);
  nand ginst25761 (P3_U4360, P3_U3033, P3_U3073);
  nand ginst25762 (P3_U4361, P3_R1110_U110, P3_U3883);
  nand ginst25763 (P3_U4362, P3_R1077_U110, P3_U3885);
  nand ginst25764 (P3_U4363, P3_R1095_U17, P3_U3884);
  nand ginst25765 (P3_U4364, P3_R1143_U110, P3_U3881);
  nand ginst25766 (P3_U4365, P3_R1161_U110, P3_U3891);
  nand ginst25767 (P3_U4366, P3_R1131_U17, P3_U3887);
  nand ginst25768 (P3_U4367, P3_R1200_U17, P3_U3017);
  not ginst25769 (P3_U4368, P3_U3330);
  nand ginst25770 (P3_U4369, P3_R1179_U17, P3_U3026);
  nand ginst25771 (P3_U4370, P3_U3025, P3_U3068);
  nand ginst25772 (P3_U4371, P3_U3437, P3_U4064);
  nand ginst25773 (P3_U4372, P3_U3644, P3_U4368);
  nand ginst25774 (P3_U4373, P3_REG0_REG_18__SCAN_IN, P3_U3022);
  nand ginst25775 (P3_U4374, P3_REG1_REG_18__SCAN_IN, P3_U3021);
  nand ginst25776 (P3_U4375, P3_REG2_REG_18__SCAN_IN, P3_U3020);
  nand ginst25777 (P3_U4376, P3_SUB_609_U11, P3_U3019);
  not ginst25778 (P3_U4377, P3_U3081);
  nand ginst25779 (P3_U4378, P3_U3033, P3_U3072);
  nand ginst25780 (P3_U4379, P3_R1110_U12, P3_U3883);
  nand ginst25781 (P3_U4380, P3_R1077_U12, P3_U3885);
  nand ginst25782 (P3_U4381, P3_R1095_U103, P3_U3884);
  nand ginst25783 (P3_U4382, P3_R1143_U12, P3_U3881);
  nand ginst25784 (P3_U4383, P3_R1161_U12, P3_U3891);
  nand ginst25785 (P3_U4384, P3_R1131_U103, P3_U3887);
  nand ginst25786 (P3_U4385, P3_R1200_U103, P3_U3017);
  not ginst25787 (P3_U4386, P3_U3331);
  nand ginst25788 (P3_U4387, P3_R1179_U103, P3_U3026);
  nand ginst25789 (P3_U4388, P3_U3025, P3_U3081);
  nand ginst25790 (P3_U4389, P3_U3440, P3_U4064);
  nand ginst25791 (P3_U4390, P3_U3648, P3_U4386);
  nand ginst25792 (P3_U4391, P3_REG0_REG_19__SCAN_IN, P3_U3022);
  nand ginst25793 (P3_U4392, P3_REG1_REG_19__SCAN_IN, P3_U3021);
  nand ginst25794 (P3_U4393, P3_REG2_REG_19__SCAN_IN, P3_U3020);
  nand ginst25795 (P3_U4394, P3_SUB_609_U15, P3_U3019);
  not ginst25796 (P3_U4395, P3_U3080);
  nand ginst25797 (P3_U4396, P3_U3033, P3_U3068);
  nand ginst25798 (P3_U4397, P3_R1110_U109, P3_U3883);
  nand ginst25799 (P3_U4398, P3_R1077_U109, P3_U3885);
  nand ginst25800 (P3_U4399, P3_R1095_U102, P3_U3884);
  nand ginst25801 (P3_U4400, P3_R1143_U109, P3_U3881);
  nand ginst25802 (P3_U4401, P3_R1161_U109, P3_U3891);
  nand ginst25803 (P3_U4402, P3_R1131_U102, P3_U3887);
  nand ginst25804 (P3_U4403, P3_R1200_U102, P3_U3017);
  not ginst25805 (P3_U4404, P3_U3332);
  nand ginst25806 (P3_U4405, P3_R1179_U102, P3_U3026);
  nand ginst25807 (P3_U4406, P3_U3025, P3_U3080);
  nand ginst25808 (P3_U4407, P3_U3443, P3_U4064);
  nand ginst25809 (P3_U4408, P3_U3651, P3_U4404);
  nand ginst25810 (P3_U4409, P3_REG2_REG_20__SCAN_IN, P3_U3020);
  nand ginst25811 (P3_U4410, P3_REG1_REG_20__SCAN_IN, P3_U3021);
  nand ginst25812 (P3_U4411, P3_REG0_REG_20__SCAN_IN, P3_U3022);
  nand ginst25813 (P3_U4412, P3_SUB_609_U20, P3_U3019);
  not ginst25814 (P3_U4413, P3_U3075);
  nand ginst25815 (P3_U4414, P3_U3033, P3_U3081);
  nand ginst25816 (P3_U4415, P3_R1110_U108, P3_U3883);
  nand ginst25817 (P3_U4416, P3_R1077_U108, P3_U3885);
  nand ginst25818 (P3_U4417, P3_R1095_U101, P3_U3884);
  nand ginst25819 (P3_U4418, P3_R1143_U108, P3_U3881);
  nand ginst25820 (P3_U4419, P3_R1161_U108, P3_U3891);
  nand ginst25821 (P3_U4420, P3_R1131_U101, P3_U3887);
  nand ginst25822 (P3_U4421, P3_R1200_U101, P3_U3017);
  not ginst25823 (P3_U4422, P3_U3333);
  nand ginst25824 (P3_U4423, P3_R1179_U101, P3_U3026);
  nand ginst25825 (P3_U4424, P3_U3025, P3_U3075);
  nand ginst25826 (P3_U4425, P3_U3445, P3_U4064);
  nand ginst25827 (P3_U4426, P3_U3654, P3_U4422);
  nand ginst25828 (P3_U4427, P3_REG2_REG_21__SCAN_IN, P3_U3020);
  nand ginst25829 (P3_U4428, P3_REG1_REG_21__SCAN_IN, P3_U3021);
  nand ginst25830 (P3_U4429, P3_REG0_REG_21__SCAN_IN, P3_U3022);
  nand ginst25831 (P3_U4430, P3_SUB_609_U27, P3_U3019);
  not ginst25832 (P3_U4431, P3_U3074);
  nand ginst25833 (P3_U4432, P3_U3033, P3_U3080);
  nand ginst25834 (P3_U4433, P3_R1110_U13, P3_U3883);
  nand ginst25835 (P3_U4434, P3_R1077_U13, P3_U3885);
  nand ginst25836 (P3_U4435, P3_R1095_U99, P3_U3884);
  nand ginst25837 (P3_U4436, P3_R1143_U13, P3_U3881);
  nand ginst25838 (P3_U4437, P3_R1161_U13, P3_U3891);
  nand ginst25839 (P3_U4438, P3_R1131_U99, P3_U3887);
  nand ginst25840 (P3_U4439, P3_R1200_U99, P3_U3017);
  not ginst25841 (P3_U4440, P3_U3335);
  nand ginst25842 (P3_U4441, P3_R1179_U99, P3_U3026);
  nand ginst25843 (P3_U4442, P3_U3025, P3_U3074);
  nand ginst25844 (P3_U4443, P3_U3907, P3_U4064);
  nand ginst25845 (P3_U4444, P3_U3657, P3_U4440);
  nand ginst25846 (P3_U4445, P3_REG2_REG_22__SCAN_IN, P3_U3020);
  nand ginst25847 (P3_U4446, P3_REG1_REG_22__SCAN_IN, P3_U3021);
  nand ginst25848 (P3_U4447, P3_REG0_REG_22__SCAN_IN, P3_U3022);
  nand ginst25849 (P3_U4448, P3_SUB_609_U17, P3_U3019);
  not ginst25850 (P3_U4449, P3_U3060);
  nand ginst25851 (P3_U4450, P3_U3033, P3_U3075);
  nand ginst25852 (P3_U4451, P3_R1110_U14, P3_U3883);
  nand ginst25853 (P3_U4452, P3_R1077_U14, P3_U3885);
  nand ginst25854 (P3_U4453, P3_R1095_U113, P3_U3884);
  nand ginst25855 (P3_U4454, P3_R1143_U14, P3_U3881);
  nand ginst25856 (P3_U4455, P3_R1161_U14, P3_U3891);
  nand ginst25857 (P3_U4456, P3_R1131_U113, P3_U3887);
  nand ginst25858 (P3_U4457, P3_R1200_U113, P3_U3017);
  not ginst25859 (P3_U4458, P3_U3337);
  nand ginst25860 (P3_U4459, P3_R1179_U113, P3_U3026);
  nand ginst25861 (P3_U4460, P3_U3025, P3_U3060);
  nand ginst25862 (P3_U4461, P3_U3906, P3_U4064);
  nand ginst25863 (P3_U4462, P3_U3660, P3_U4458);
  nand ginst25864 (P3_U4463, P3_REG2_REG_23__SCAN_IN, P3_U3020);
  nand ginst25865 (P3_U4464, P3_REG1_REG_23__SCAN_IN, P3_U3021);
  nand ginst25866 (P3_U4465, P3_REG0_REG_23__SCAN_IN, P3_U3022);
  nand ginst25867 (P3_U4466, P3_SUB_609_U6, P3_U3019);
  not ginst25868 (P3_U4467, P3_U3065);
  nand ginst25869 (P3_U4468, P3_U3033, P3_U3074);
  nand ginst25870 (P3_U4469, P3_R1110_U107, P3_U3883);
  nand ginst25871 (P3_U4470, P3_R1077_U107, P3_U3885);
  nand ginst25872 (P3_U4471, P3_R1095_U112, P3_U3884);
  nand ginst25873 (P3_U4472, P3_R1143_U107, P3_U3881);
  nand ginst25874 (P3_U4473, P3_R1161_U107, P3_U3891);
  nand ginst25875 (P3_U4474, P3_R1131_U112, P3_U3887);
  nand ginst25876 (P3_U4475, P3_R1200_U112, P3_U3017);
  not ginst25877 (P3_U4476, P3_U3339);
  nand ginst25878 (P3_U4477, P3_R1179_U112, P3_U3026);
  nand ginst25879 (P3_U4478, P3_U3025, P3_U3065);
  nand ginst25880 (P3_U4479, P3_U3905, P3_U4064);
  nand ginst25881 (P3_U4480, P3_U3663, P3_U4476);
  nand ginst25882 (P3_U4481, P3_REG2_REG_24__SCAN_IN, P3_U3020);
  nand ginst25883 (P3_U4482, P3_REG1_REG_24__SCAN_IN, P3_U3021);
  nand ginst25884 (P3_U4483, P3_REG0_REG_24__SCAN_IN, P3_U3022);
  nand ginst25885 (P3_U4484, P3_SUB_609_U10, P3_U3019);
  not ginst25886 (P3_U4485, P3_U3064);
  nand ginst25887 (P3_U4486, P3_U3033, P3_U3060);
  nand ginst25888 (P3_U4487, P3_R1110_U106, P3_U3883);
  nand ginst25889 (P3_U4488, P3_R1077_U106, P3_U3885);
  nand ginst25890 (P3_U4489, P3_R1095_U18, P3_U3884);
  nand ginst25891 (P3_U4490, P3_R1143_U106, P3_U3881);
  nand ginst25892 (P3_U4491, P3_R1161_U106, P3_U3891);
  nand ginst25893 (P3_U4492, P3_R1131_U18, P3_U3887);
  nand ginst25894 (P3_U4493, P3_R1200_U18, P3_U3017);
  not ginst25895 (P3_U4494, P3_U3341);
  nand ginst25896 (P3_U4495, P3_R1179_U18, P3_U3026);
  nand ginst25897 (P3_U4496, P3_U3025, P3_U3064);
  nand ginst25898 (P3_U4497, P3_U3904, P3_U4064);
  nand ginst25899 (P3_U4498, P3_U3666, P3_U4494);
  nand ginst25900 (P3_U4499, P3_REG2_REG_25__SCAN_IN, P3_U3020);
  nand ginst25901 (P3_U4500, P3_REG1_REG_25__SCAN_IN, P3_U3021);
  nand ginst25902 (P3_U4501, P3_REG0_REG_25__SCAN_IN, P3_U3022);
  nand ginst25903 (P3_U4502, P3_SUB_609_U16, P3_U3019);
  not ginst25904 (P3_U4503, P3_U3057);
  nand ginst25905 (P3_U4504, P3_U3033, P3_U3065);
  nand ginst25906 (P3_U4505, P3_R1110_U105, P3_U3883);
  nand ginst25907 (P3_U4506, P3_R1077_U105, P3_U3885);
  nand ginst25908 (P3_U4507, P3_R1095_U98, P3_U3884);
  nand ginst25909 (P3_U4508, P3_R1143_U105, P3_U3881);
  nand ginst25910 (P3_U4509, P3_R1161_U105, P3_U3891);
  nand ginst25911 (P3_U4510, P3_R1131_U98, P3_U3887);
  nand ginst25912 (P3_U4511, P3_R1200_U98, P3_U3017);
  not ginst25913 (P3_U4512, P3_U3343);
  nand ginst25914 (P3_U4513, P3_R1179_U98, P3_U3026);
  nand ginst25915 (P3_U4514, P3_U3025, P3_U3057);
  nand ginst25916 (P3_U4515, P3_U3903, P3_U4064);
  nand ginst25917 (P3_U4516, P3_U3670, P3_U4512);
  nand ginst25918 (P3_U4517, P3_REG2_REG_26__SCAN_IN, P3_U3020);
  nand ginst25919 (P3_U4518, P3_REG1_REG_26__SCAN_IN, P3_U3021);
  nand ginst25920 (P3_U4519, P3_REG0_REG_26__SCAN_IN, P3_U3022);
  nand ginst25921 (P3_U4520, P3_SUB_609_U26, P3_U3019);
  not ginst25922 (P3_U4521, P3_U3056);
  nand ginst25923 (P3_U4522, P3_U3033, P3_U3064);
  nand ginst25924 (P3_U4523, P3_R1110_U104, P3_U3883);
  nand ginst25925 (P3_U4524, P3_R1077_U104, P3_U3885);
  nand ginst25926 (P3_U4525, P3_R1095_U97, P3_U3884);
  nand ginst25927 (P3_U4526, P3_R1143_U104, P3_U3881);
  nand ginst25928 (P3_U4527, P3_R1161_U104, P3_U3891);
  nand ginst25929 (P3_U4528, P3_R1131_U97, P3_U3887);
  nand ginst25930 (P3_U4529, P3_R1200_U97, P3_U3017);
  not ginst25931 (P3_U4530, P3_U3345);
  nand ginst25932 (P3_U4531, P3_R1179_U97, P3_U3026);
  nand ginst25933 (P3_U4532, P3_U3025, P3_U3056);
  nand ginst25934 (P3_U4533, P3_U3902, P3_U4064);
  nand ginst25935 (P3_U4534, P3_U3674, P3_U4530);
  nand ginst25936 (P3_U4535, P3_REG2_REG_27__SCAN_IN, P3_U3020);
  nand ginst25937 (P3_U4536, P3_REG1_REG_27__SCAN_IN, P3_U3021);
  nand ginst25938 (P3_U4537, P3_REG0_REG_27__SCAN_IN, P3_U3022);
  nand ginst25939 (P3_U4538, P3_SUB_609_U22, P3_U3019);
  not ginst25940 (P3_U4539, P3_U3052);
  nand ginst25941 (P3_U4540, P3_U3033, P3_U3057);
  nand ginst25942 (P3_U4541, P3_R1110_U15, P3_U3883);
  nand ginst25943 (P3_U4542, P3_R1077_U15, P3_U3885);
  nand ginst25944 (P3_U4543, P3_R1095_U111, P3_U3884);
  nand ginst25945 (P3_U4544, P3_R1143_U15, P3_U3881);
  nand ginst25946 (P3_U4545, P3_R1161_U15, P3_U3891);
  nand ginst25947 (P3_U4546, P3_R1131_U111, P3_U3887);
  nand ginst25948 (P3_U4547, P3_R1200_U111, P3_U3017);
  not ginst25949 (P3_U4548, P3_U3347);
  nand ginst25950 (P3_U4549, P3_R1179_U111, P3_U3026);
  nand ginst25951 (P3_U4550, P3_U3025, P3_U3052);
  nand ginst25952 (P3_U4551, P3_U3901, P3_U4064);
  nand ginst25953 (P3_U4552, P3_U3678, P3_U4548);
  nand ginst25954 (P3_U4553, P3_REG2_REG_28__SCAN_IN, P3_U3020);
  nand ginst25955 (P3_U4554, P3_REG1_REG_28__SCAN_IN, P3_U3021);
  nand ginst25956 (P3_U4555, P3_REG0_REG_28__SCAN_IN, P3_U3022);
  nand ginst25957 (P3_U4556, P3_SUB_609_U28, P3_U3019);
  not ginst25958 (P3_U4557, P3_U3053);
  nand ginst25959 (P3_U4558, P3_U3033, P3_U3056);
  nand ginst25960 (P3_U4559, P3_R1110_U103, P3_U3883);
  nand ginst25961 (P3_U4560, P3_R1077_U103, P3_U3885);
  nand ginst25962 (P3_U4561, P3_R1095_U19, P3_U3884);
  nand ginst25963 (P3_U4562, P3_R1143_U103, P3_U3881);
  nand ginst25964 (P3_U4563, P3_R1161_U103, P3_U3891);
  nand ginst25965 (P3_U4564, P3_R1131_U19, P3_U3887);
  nand ginst25966 (P3_U4565, P3_R1200_U19, P3_U3017);
  not ginst25967 (P3_U4566, P3_U3349);
  nand ginst25968 (P3_U4567, P3_R1179_U19, P3_U3026);
  nand ginst25969 (P3_U4568, P3_U3025, P3_U3053);
  nand ginst25970 (P3_U4569, P3_U3900, P3_U4064);
  nand ginst25971 (P3_U4570, P3_U3682, P3_U4566);
  nand ginst25972 (P3_U4571, P3_SUB_609_U92, P3_U3019);
  nand ginst25973 (P3_U4572, P3_REG2_REG_29__SCAN_IN, P3_U3020);
  nand ginst25974 (P3_U4573, P3_REG1_REG_29__SCAN_IN, P3_U3021);
  nand ginst25975 (P3_U4574, P3_REG0_REG_29__SCAN_IN, P3_U3022);
  not ginst25976 (P3_U4575, P3_U3054);
  nand ginst25977 (P3_U4576, P3_U3033, P3_U3052);
  nand ginst25978 (P3_U4577, P3_R1110_U102, P3_U3883);
  nand ginst25979 (P3_U4578, P3_R1077_U102, P3_U3885);
  nand ginst25980 (P3_U4579, P3_R1095_U96, P3_U3884);
  nand ginst25981 (P3_U4580, P3_R1143_U102, P3_U3881);
  nand ginst25982 (P3_U4581, P3_R1161_U102, P3_U3891);
  nand ginst25983 (P3_U4582, P3_R1131_U96, P3_U3887);
  nand ginst25984 (P3_U4583, P3_R1200_U96, P3_U3017);
  not ginst25985 (P3_U4584, P3_U3351);
  nand ginst25986 (P3_U4585, P3_R1179_U96, P3_U3026);
  nand ginst25987 (P3_U4586, P3_U3025, P3_U3054);
  nand ginst25988 (P3_U4587, P3_U3899, P3_U4064);
  nand ginst25989 (P3_U4588, P3_U3686, P3_U4584);
  nand ginst25990 (P3_U4589, P3_REG2_REG_30__SCAN_IN, P3_U3020);
  nand ginst25991 (P3_U4590, P3_REG1_REG_30__SCAN_IN, P3_U3021);
  nand ginst25992 (P3_U4591, P3_REG0_REG_30__SCAN_IN, P3_U3022);
  nand ginst25993 (P3_U4592, P3_SUB_609_U92, P3_U3019);
  not ginst25994 (P3_U4593, P3_U3058);
  nand ginst25995 (P3_U4594, P3_U3298, P3_U3892);
  nand ginst25996 (P3_U4595, P3_U3833, P3_U4594);
  nand ginst25997 (P3_U4596, P3_U3058, P3_U3911, P3_U4595);
  nand ginst25998 (P3_U4597, P3_U3033, P3_U3053);
  nand ginst25999 (P3_U4598, P3_R1110_U101, P3_U3883);
  nand ginst26000 (P3_U4599, P3_R1077_U101, P3_U3885);
  nand ginst26001 (P3_U4600, P3_R1095_U20, P3_U3884);
  nand ginst26002 (P3_U4601, P3_R1143_U101, P3_U3881);
  nand ginst26003 (P3_U4602, P3_R1161_U101, P3_U3891);
  nand ginst26004 (P3_U4603, P3_R1131_U20, P3_U3887);
  nand ginst26005 (P3_U4604, P3_R1200_U20, P3_U3017);
  not ginst26006 (P3_U4605, P3_U3354);
  nand ginst26007 (P3_U4606, P3_R1179_U20, P3_U3026);
  nand ginst26008 (P3_U4607, P3_U3908, P3_U4064);
  nand ginst26009 (P3_U4608, P3_U3690, P3_U4605);
  nand ginst26010 (P3_U4609, P3_SUB_609_U92, P3_U3019);
  nand ginst26011 (P3_U4610, P3_REG2_REG_31__SCAN_IN, P3_U3020);
  nand ginst26012 (P3_U4611, P3_REG1_REG_31__SCAN_IN, P3_U3021);
  nand ginst26013 (P3_U4612, P3_REG0_REG_31__SCAN_IN, P3_U3022);
  not ginst26014 (P3_U4613, P3_U3055);
  nand ginst26015 (P3_U4614, P3_U3873, P3_U4064);
  nand ginst26016 (P3_U4615, P3_U3361, P3_U4614);
  nand ginst26017 (P3_U4616, P3_U3872, P3_U4064);
  nand ginst26018 (P3_U4617, P3_U3361, P3_U4616);
  nand ginst26019 (P3_U4618, P3_U3302, P3_U5640, P3_U5641);
  nand ginst26020 (P3_U4619, P3_U3367, P3_U3888);
  nand ginst26021 (P3_U4620, P3_U3048, P3_U4619);
  nand ginst26022 (P3_U4621, P3_U3047, P3_U4618);
  nand ginst26023 (P3_U4622, P3_U4620, P3_U4621);
  nand ginst26024 (P3_U4623, P3_U3379, P3_U5456);
  nand ginst26025 (P3_U4624, P3_U3380, P3_U3834, P3_U4623);
  nand ginst26026 (P3_U4625, P3_U3048, P3_U4624);
  nand ginst26027 (P3_U4626, P3_U3047, P3_U4619);
  nand ginst26028 (P3_U4627, P3_U3360, P3_U4625, P3_U4626);
  not ginst26029 (P3_U4628, P3_U3365);
  nand ginst26030 (P3_U4629, P3_U3034, P3_U3077);
  nand ginst26031 (P3_U4630, P3_R1179_U24, P3_U3030);
  nand ginst26032 (P3_U4631, P3_U3029, P3_U3387);
  nand ginst26033 (P3_U4632, P3_REG3_REG_0__SCAN_IN, P3_U3028);
  nand ginst26034 (P3_U4633, P3_U3034, P3_U3067);
  nand ginst26035 (P3_U4634, P3_R1179_U100, P3_U3030);
  nand ginst26036 (P3_U4635, P3_U3029, P3_U3392);
  nand ginst26037 (P3_U4636, P3_REG3_REG_1__SCAN_IN, P3_U3028);
  nand ginst26038 (P3_U4637, P3_U3034, P3_U3063);
  nand ginst26039 (P3_U4638, P3_R1179_U110, P3_U3030);
  nand ginst26040 (P3_U4639, P3_U3029, P3_U3395);
  nand ginst26041 (P3_U4640, P3_REG3_REG_2__SCAN_IN, P3_U3028);
  nand ginst26042 (P3_U4641, P3_U3034, P3_U3059);
  nand ginst26043 (P3_U4642, P3_R1179_U21, P3_U3030);
  nand ginst26044 (P3_U4643, P3_U3029, P3_U3398);
  nand ginst26045 (P3_U4644, P3_SUB_609_U25, P3_U3028);
  nand ginst26046 (P3_U4645, P3_U3034, P3_U3066);
  nand ginst26047 (P3_U4646, P3_R1179_U109, P3_U3030);
  nand ginst26048 (P3_U4647, P3_U3029, P3_U3401);
  nand ginst26049 (P3_U4648, P3_SUB_609_U29, P3_U3028);
  nand ginst26050 (P3_U4649, P3_U3034, P3_U3070);
  nand ginst26051 (P3_U4650, P3_R1179_U108, P3_U3030);
  nand ginst26052 (P3_U4651, P3_U3029, P3_U3404);
  nand ginst26053 (P3_U4652, P3_SUB_609_U53, P3_U3028);
  nand ginst26054 (P3_U4653, P3_U3034, P3_U3069);
  nand ginst26055 (P3_U4654, P3_R1179_U22, P3_U3030);
  nand ginst26056 (P3_U4655, P3_U3029, P3_U3407);
  nand ginst26057 (P3_U4656, P3_SUB_609_U8, P3_U3028);
  nand ginst26058 (P3_U4657, P3_U3034, P3_U3083);
  nand ginst26059 (P3_U4658, P3_R1179_U107, P3_U3030);
  nand ginst26060 (P3_U4659, P3_U3029, P3_U3410);
  nand ginst26061 (P3_U4660, P3_SUB_609_U18, P3_U3028);
  nand ginst26062 (P3_U4661, P3_U3034, P3_U3082);
  nand ginst26063 (P3_U4662, P3_R1179_U23, P3_U3030);
  nand ginst26064 (P3_U4663, P3_U3029, P3_U3413);
  nand ginst26065 (P3_U4664, P3_SUB_609_U12, P3_U3028);
  nand ginst26066 (P3_U4665, P3_U3034, P3_U3061);
  nand ginst26067 (P3_U4666, P3_R1179_U106, P3_U3030);
  nand ginst26068 (P3_U4667, P3_U3029, P3_U3416);
  nand ginst26069 (P3_U4668, P3_SUB_609_U14, P3_U3028);
  nand ginst26070 (P3_U4669, P3_U3034, P3_U3062);
  nand ginst26071 (P3_U4670, P3_R1179_U116, P3_U3030);
  nand ginst26072 (P3_U4671, P3_U3029, P3_U3419);
  nand ginst26073 (P3_U4672, P3_SUB_609_U13, P3_U3028);
  nand ginst26074 (P3_U4673, P3_U3034, P3_U3071);
  nand ginst26075 (P3_U4674, P3_R1179_U16, P3_U3030);
  nand ginst26076 (P3_U4675, P3_U3029, P3_U3422);
  nand ginst26077 (P3_U4676, P3_SUB_609_U9, P3_U3028);
  nand ginst26078 (P3_U4677, P3_U3034, P3_U3079);
  nand ginst26079 (P3_U4678, P3_R1179_U105, P3_U3030);
  nand ginst26080 (P3_U4679, P3_U3029, P3_U3425);
  nand ginst26081 (P3_U4680, P3_SUB_609_U23, P3_U3028);
  nand ginst26082 (P3_U4681, P3_U3034, P3_U3078);
  nand ginst26083 (P3_U4682, P3_R1179_U104, P3_U3030);
  nand ginst26084 (P3_U4683, P3_U3029, P3_U3428);
  nand ginst26085 (P3_U4684, P3_SUB_609_U24, P3_U3028);
  nand ginst26086 (P3_U4685, P3_U3034, P3_U3073);
  nand ginst26087 (P3_U4686, P3_R1179_U115, P3_U3030);
  nand ginst26088 (P3_U4687, P3_U3029, P3_U3431);
  nand ginst26089 (P3_U4688, P3_SUB_609_U30, P3_U3028);
  nand ginst26090 (P3_U4689, P3_U3034, P3_U3072);
  nand ginst26091 (P3_U4690, P3_R1179_U114, P3_U3030);
  nand ginst26092 (P3_U4691, P3_U3029, P3_U3434);
  nand ginst26093 (P3_U4692, P3_SUB_609_U21, P3_U3028);
  nand ginst26094 (P3_U4693, P3_U3034, P3_U3068);
  nand ginst26095 (P3_U4694, P3_R1179_U17, P3_U3030);
  nand ginst26096 (P3_U4695, P3_U3029, P3_U3437);
  nand ginst26097 (P3_U4696, P3_SUB_609_U7, P3_U3028);
  nand ginst26098 (P3_U4697, P3_U3034, P3_U3081);
  nand ginst26099 (P3_U4698, P3_R1179_U103, P3_U3030);
  nand ginst26100 (P3_U4699, P3_U3029, P3_U3440);
  nand ginst26101 (P3_U4700, P3_SUB_609_U19, P3_U3028);
  nand ginst26102 (P3_U4701, P3_U3034, P3_U3080);
  nand ginst26103 (P3_U4702, P3_R1179_U102, P3_U3030);
  nand ginst26104 (P3_U4703, P3_U3029, P3_U3443);
  nand ginst26105 (P3_U4704, P3_SUB_609_U11, P3_U3028);
  nand ginst26106 (P3_U4705, P3_U3034, P3_U3075);
  nand ginst26107 (P3_U4706, P3_R1179_U101, P3_U3030);
  nand ginst26108 (P3_U4707, P3_U3029, P3_U3445);
  nand ginst26109 (P3_U4708, P3_SUB_609_U15, P3_U3028);
  nand ginst26110 (P3_U4709, P3_U3034, P3_U3074);
  nand ginst26111 (P3_U4710, P3_R1179_U99, P3_U3030);
  nand ginst26112 (P3_U4711, P3_U3029, P3_U3907);
  nand ginst26113 (P3_U4712, P3_SUB_609_U20, P3_U3028);
  nand ginst26114 (P3_U4713, P3_U3034, P3_U3060);
  nand ginst26115 (P3_U4714, P3_R1179_U113, P3_U3030);
  nand ginst26116 (P3_U4715, P3_U3029, P3_U3906);
  nand ginst26117 (P3_U4716, P3_SUB_609_U27, P3_U3028);
  nand ginst26118 (P3_U4717, P3_U3034, P3_U3065);
  nand ginst26119 (P3_U4718, P3_R1179_U112, P3_U3030);
  nand ginst26120 (P3_U4719, P3_U3029, P3_U3905);
  nand ginst26121 (P3_U4720, P3_SUB_609_U17, P3_U3028);
  nand ginst26122 (P3_U4721, P3_U3034, P3_U3064);
  nand ginst26123 (P3_U4722, P3_R1179_U18, P3_U3030);
  nand ginst26124 (P3_U4723, P3_U3029, P3_U3904);
  nand ginst26125 (P3_U4724, P3_SUB_609_U6, P3_U3028);
  nand ginst26126 (P3_U4725, P3_U3034, P3_U3057);
  nand ginst26127 (P3_U4726, P3_R1179_U98, P3_U3030);
  nand ginst26128 (P3_U4727, P3_U3029, P3_U3903);
  nand ginst26129 (P3_U4728, P3_SUB_609_U10, P3_U3028);
  nand ginst26130 (P3_U4729, P3_U3034, P3_U3056);
  nand ginst26131 (P3_U4730, P3_R1179_U97, P3_U3030);
  nand ginst26132 (P3_U4731, P3_U3029, P3_U3902);
  nand ginst26133 (P3_U4732, P3_SUB_609_U16, P3_U3028);
  nand ginst26134 (P3_U4733, P3_U3034, P3_U3052);
  nand ginst26135 (P3_U4734, P3_R1179_U111, P3_U3030);
  nand ginst26136 (P3_U4735, P3_U3029, P3_U3901);
  nand ginst26137 (P3_U4736, P3_SUB_609_U26, P3_U3028);
  nand ginst26138 (P3_U4737, P3_U3034, P3_U3053);
  nand ginst26139 (P3_U4738, P3_R1179_U19, P3_U3030);
  nand ginst26140 (P3_U4739, P3_U3029, P3_U3900);
  nand ginst26141 (P3_U4740, P3_SUB_609_U22, P3_U3028);
  nand ginst26142 (P3_U4741, P3_U3034, P3_U3054);
  nand ginst26143 (P3_U4742, P3_R1179_U96, P3_U3030);
  nand ginst26144 (P3_U4743, P3_U3029, P3_U3899);
  nand ginst26145 (P3_U4744, P3_SUB_609_U28, P3_U3028);
  nand ginst26146 (P3_U4745, P3_R1179_U20, P3_U3030);
  nand ginst26147 (P3_U4746, P3_U3029, P3_U3908);
  nand ginst26148 (P3_U4747, P3_SUB_609_U92, P3_U3028);
  nand ginst26149 (P3_U4748, P3_SUB_609_U92, P3_U3028);
  nand ginst26150 (P3_U4749, P3_U3912, P3_U3916);
  nand ginst26151 (P3_U4750, P3_U3029, P3_U3873);
  nand ginst26152 (P3_U4751, P3_REG2_REG_30__SCAN_IN, P3_U3358);
  nand ginst26153 (P3_U4752, P3_U3029, P3_U3872);
  nand ginst26154 (P3_U4753, P3_REG2_REG_31__SCAN_IN, P3_U3358);
  nand ginst26155 (P3_U4754, P3_U3359, P3_U3697, P3_U3698, P3_U4628);
  nand ginst26156 (P3_U4755, P3_R1212_U6, P3_U3040);
  nand ginst26157 (P3_U4756, P3_U3039, P3_U3379);
  nand ginst26158 (P3_U4757, P3_R1209_U6, P3_U3037);
  nand ginst26159 (P3_U4758, P3_U4755, P3_U4756, P3_U4757);
  nand ginst26160 (P3_U4759, P3_U3910, P3_U5440);
  not ginst26161 (P3_U4760, P3_U3366);
  nand ginst26162 (P3_U4761, P3_U3833, P3_U3896);
  nand ginst26163 (P3_U4762, P3_R1054_U67, P3_U3051);
  nand ginst26164 (P3_U4763, P3_U3379, P3_U5768);
  nand ginst26165 (P3_U4764, P3_U3042, P3_U4758);
  nand ginst26166 (P3_U4765, P3_R1212_U6, P3_U3041);
  nand ginst26167 (P3_U4766, P3_REG3_REG_19__SCAN_IN, P3_U3151);
  nand ginst26168 (P3_U4767, P3_R1209_U6, P3_U3038);
  nand ginst26169 (P3_U4768, P3_ADDR_REG_19__SCAN_IN, P3_U4760);
  nand ginst26170 (P3_U4769, P3_R1212_U58, P3_U3040);
  nand ginst26171 (P3_U4770, P3_U3039, P3_U3442);
  nand ginst26172 (P3_U4771, P3_R1209_U58, P3_U3037);
  nand ginst26173 (P3_U4772, P3_U4769, P3_U4770, P3_U4771);
  nand ginst26174 (P3_U4773, P3_R1054_U68, P3_U3051);
  nand ginst26175 (P3_U4774, P3_U3442, P3_U5768);
  nand ginst26176 (P3_U4775, P3_U3042, P3_U4772);
  nand ginst26177 (P3_U4776, P3_R1212_U58, P3_U3041);
  nand ginst26178 (P3_U4777, P3_REG3_REG_18__SCAN_IN, P3_U3151);
  nand ginst26179 (P3_U4778, P3_R1209_U58, P3_U3038);
  nand ginst26180 (P3_U4779, P3_ADDR_REG_18__SCAN_IN, P3_U4760);
  nand ginst26181 (P3_U4780, P3_R1212_U59, P3_U3040);
  nand ginst26182 (P3_U4781, P3_U3039, P3_U3439);
  nand ginst26183 (P3_U4782, P3_R1209_U59, P3_U3037);
  nand ginst26184 (P3_U4783, P3_U4780, P3_U4781, P3_U4782);
  nand ginst26185 (P3_U4784, P3_R1054_U69, P3_U3051);
  nand ginst26186 (P3_U4785, P3_U3439, P3_U5768);
  nand ginst26187 (P3_U4786, P3_U3042, P3_U4783);
  nand ginst26188 (P3_U4787, P3_R1212_U59, P3_U3041);
  nand ginst26189 (P3_U4788, P3_REG3_REG_17__SCAN_IN, P3_U3151);
  nand ginst26190 (P3_U4789, P3_R1209_U59, P3_U3038);
  nand ginst26191 (P3_U4790, P3_ADDR_REG_17__SCAN_IN, P3_U4760);
  nand ginst26192 (P3_U4791, P3_R1212_U60, P3_U3040);
  nand ginst26193 (P3_U4792, P3_U3039, P3_U3436);
  nand ginst26194 (P3_U4793, P3_R1209_U60, P3_U3037);
  nand ginst26195 (P3_U4794, P3_U4791, P3_U4792, P3_U4793);
  nand ginst26196 (P3_U4795, P3_R1054_U13, P3_U3051);
  nand ginst26197 (P3_U4796, P3_U3436, P3_U5768);
  nand ginst26198 (P3_U4797, P3_U3042, P3_U4794);
  nand ginst26199 (P3_U4798, P3_R1212_U60, P3_U3041);
  nand ginst26200 (P3_U4799, P3_REG3_REG_16__SCAN_IN, P3_U3151);
  nand ginst26201 (P3_U4800, P3_R1209_U60, P3_U3038);
  nand ginst26202 (P3_U4801, P3_ADDR_REG_16__SCAN_IN, P3_U4760);
  nand ginst26203 (P3_U4802, P3_R1212_U61, P3_U3040);
  nand ginst26204 (P3_U4803, P3_U3039, P3_U3433);
  nand ginst26205 (P3_U4804, P3_R1209_U61, P3_U3037);
  nand ginst26206 (P3_U4805, P3_U4802, P3_U4803, P3_U4804);
  nand ginst26207 (P3_U4806, P3_R1054_U77, P3_U3051);
  nand ginst26208 (P3_U4807, P3_U3433, P3_U5768);
  nand ginst26209 (P3_U4808, P3_U3042, P3_U4805);
  nand ginst26210 (P3_U4809, P3_R1212_U61, P3_U3041);
  nand ginst26211 (P3_U4810, P3_REG3_REG_15__SCAN_IN, P3_U3151);
  nand ginst26212 (P3_U4811, P3_R1209_U61, P3_U3038);
  nand ginst26213 (P3_U4812, P3_ADDR_REG_15__SCAN_IN, P3_U4760);
  nand ginst26214 (P3_U4813, P3_R1212_U62, P3_U3040);
  nand ginst26215 (P3_U4814, P3_U3039, P3_U3430);
  nand ginst26216 (P3_U4815, P3_R1209_U62, P3_U3037);
  nand ginst26217 (P3_U4816, P3_U4813, P3_U4814, P3_U4815);
  nand ginst26218 (P3_U4817, P3_R1054_U78, P3_U3051);
  nand ginst26219 (P3_U4818, P3_U3430, P3_U5768);
  nand ginst26220 (P3_U4819, P3_U3042, P3_U4816);
  nand ginst26221 (P3_U4820, P3_R1212_U62, P3_U3041);
  nand ginst26222 (P3_U4821, P3_REG3_REG_14__SCAN_IN, P3_U3151);
  nand ginst26223 (P3_U4822, P3_R1209_U62, P3_U3038);
  nand ginst26224 (P3_U4823, P3_ADDR_REG_14__SCAN_IN, P3_U4760);
  nand ginst26225 (P3_U4824, P3_R1212_U63, P3_U3040);
  nand ginst26226 (P3_U4825, P3_U3039, P3_U3427);
  nand ginst26227 (P3_U4826, P3_R1209_U63, P3_U3037);
  nand ginst26228 (P3_U4827, P3_U4824, P3_U4825, P3_U4826);
  nand ginst26229 (P3_U4828, P3_R1054_U70, P3_U3051);
  nand ginst26230 (P3_U4829, P3_U3427, P3_U5768);
  nand ginst26231 (P3_U4830, P3_U3042, P3_U4827);
  nand ginst26232 (P3_U4831, P3_R1212_U63, P3_U3041);
  nand ginst26233 (P3_U4832, P3_REG3_REG_13__SCAN_IN, P3_U3151);
  nand ginst26234 (P3_U4833, P3_R1209_U63, P3_U3038);
  nand ginst26235 (P3_U4834, P3_ADDR_REG_13__SCAN_IN, P3_U4760);
  nand ginst26236 (P3_U4835, P3_R1212_U64, P3_U3040);
  nand ginst26237 (P3_U4836, P3_U3039, P3_U3424);
  nand ginst26238 (P3_U4837, P3_R1209_U64, P3_U3037);
  nand ginst26239 (P3_U4838, P3_U4835, P3_U4836, P3_U4837);
  nand ginst26240 (P3_U4839, P3_R1054_U71, P3_U3051);
  nand ginst26241 (P3_U4840, P3_U3424, P3_U5768);
  nand ginst26242 (P3_U4841, P3_U3042, P3_U4838);
  nand ginst26243 (P3_U4842, P3_R1212_U64, P3_U3041);
  nand ginst26244 (P3_U4843, P3_REG3_REG_12__SCAN_IN, P3_U3151);
  nand ginst26245 (P3_U4844, P3_R1209_U64, P3_U3038);
  nand ginst26246 (P3_U4845, P3_ADDR_REG_12__SCAN_IN, P3_U4760);
  nand ginst26247 (P3_U4846, P3_R1212_U65, P3_U3040);
  nand ginst26248 (P3_U4847, P3_U3039, P3_U3421);
  nand ginst26249 (P3_U4848, P3_R1209_U65, P3_U3037);
  nand ginst26250 (P3_U4849, P3_U4846, P3_U4847, P3_U4848);
  nand ginst26251 (P3_U4850, P3_R1054_U12, P3_U3051);
  nand ginst26252 (P3_U4851, P3_U3421, P3_U5768);
  nand ginst26253 (P3_U4852, P3_U3042, P3_U4849);
  nand ginst26254 (P3_U4853, P3_R1212_U65, P3_U3041);
  nand ginst26255 (P3_U4854, P3_REG3_REG_11__SCAN_IN, P3_U3151);
  nand ginst26256 (P3_U4855, P3_R1209_U65, P3_U3038);
  nand ginst26257 (P3_U4856, P3_ADDR_REG_11__SCAN_IN, P3_U4760);
  nand ginst26258 (P3_U4857, P3_R1212_U66, P3_U3040);
  nand ginst26259 (P3_U4858, P3_U3039, P3_U3418);
  nand ginst26260 (P3_U4859, P3_R1209_U66, P3_U3037);
  nand ginst26261 (P3_U4860, P3_U4857, P3_U4858, P3_U4859);
  nand ginst26262 (P3_U4861, P3_R1054_U79, P3_U3051);
  nand ginst26263 (P3_U4862, P3_U3418, P3_U5768);
  nand ginst26264 (P3_U4863, P3_U3042, P3_U4860);
  nand ginst26265 (P3_U4864, P3_R1212_U66, P3_U3041);
  nand ginst26266 (P3_U4865, P3_REG3_REG_10__SCAN_IN, P3_U3151);
  nand ginst26267 (P3_U4866, P3_R1209_U66, P3_U3038);
  nand ginst26268 (P3_U4867, P3_ADDR_REG_10__SCAN_IN, P3_U4760);
  nand ginst26269 (P3_U4868, P3_R1212_U49, P3_U3040);
  nand ginst26270 (P3_U4869, P3_U3039, P3_U3415);
  nand ginst26271 (P3_U4870, P3_R1209_U49, P3_U3037);
  nand ginst26272 (P3_U4871, P3_U4868, P3_U4869, P3_U4870);
  nand ginst26273 (P3_U4872, P3_R1054_U72, P3_U3051);
  nand ginst26274 (P3_U4873, P3_U3415, P3_U5768);
  nand ginst26275 (P3_U4874, P3_U3042, P3_U4871);
  nand ginst26276 (P3_U4875, P3_R1212_U49, P3_U3041);
  nand ginst26277 (P3_U4876, P3_REG3_REG_9__SCAN_IN, P3_U3151);
  nand ginst26278 (P3_U4877, P3_R1209_U49, P3_U3038);
  nand ginst26279 (P3_U4878, P3_ADDR_REG_9__SCAN_IN, P3_U4760);
  nand ginst26280 (P3_U4879, P3_R1212_U50, P3_U3040);
  nand ginst26281 (P3_U4880, P3_U3039, P3_U3412);
  nand ginst26282 (P3_U4881, P3_R1209_U50, P3_U3037);
  nand ginst26283 (P3_U4882, P3_U4879, P3_U4880, P3_U4881);
  nand ginst26284 (P3_U4883, P3_R1054_U16, P3_U3051);
  nand ginst26285 (P3_U4884, P3_U3412, P3_U5768);
  nand ginst26286 (P3_U4885, P3_U3042, P3_U4882);
  nand ginst26287 (P3_U4886, P3_R1212_U50, P3_U3041);
  nand ginst26288 (P3_U4887, P3_REG3_REG_8__SCAN_IN, P3_U3151);
  nand ginst26289 (P3_U4888, P3_R1209_U50, P3_U3038);
  nand ginst26290 (P3_U4889, P3_ADDR_REG_8__SCAN_IN, P3_U4760);
  nand ginst26291 (P3_U4890, P3_R1212_U51, P3_U3040);
  nand ginst26292 (P3_U4891, P3_U3039, P3_U3409);
  nand ginst26293 (P3_U4892, P3_R1209_U51, P3_U3037);
  nand ginst26294 (P3_U4893, P3_U4890, P3_U4891, P3_U4892);
  nand ginst26295 (P3_U4894, P3_R1054_U73, P3_U3051);
  nand ginst26296 (P3_U4895, P3_U3409, P3_U5768);
  nand ginst26297 (P3_U4896, P3_U3042, P3_U4893);
  nand ginst26298 (P3_U4897, P3_R1212_U51, P3_U3041);
  nand ginst26299 (P3_U4898, P3_REG3_REG_7__SCAN_IN, P3_U3151);
  nand ginst26300 (P3_U4899, P3_R1209_U51, P3_U3038);
  nand ginst26301 (P3_U4900, P3_ADDR_REG_7__SCAN_IN, P3_U4760);
  nand ginst26302 (P3_U4901, P3_R1212_U52, P3_U3040);
  nand ginst26303 (P3_U4902, P3_U3039, P3_U3406);
  nand ginst26304 (P3_U4903, P3_R1209_U52, P3_U3037);
  nand ginst26305 (P3_U4904, P3_U4901, P3_U4902, P3_U4903);
  nand ginst26306 (P3_U4905, P3_R1054_U15, P3_U3051);
  nand ginst26307 (P3_U4906, P3_U3406, P3_U5768);
  nand ginst26308 (P3_U4907, P3_U3042, P3_U4904);
  nand ginst26309 (P3_U4908, P3_R1212_U52, P3_U3041);
  nand ginst26310 (P3_U4909, P3_REG3_REG_6__SCAN_IN, P3_U3151);
  nand ginst26311 (P3_U4910, P3_R1209_U52, P3_U3038);
  nand ginst26312 (P3_U4911, P3_ADDR_REG_6__SCAN_IN, P3_U4760);
  nand ginst26313 (P3_U4912, P3_R1212_U53, P3_U3040);
  nand ginst26314 (P3_U4913, P3_U3039, P3_U3403);
  nand ginst26315 (P3_U4914, P3_R1209_U53, P3_U3037);
  nand ginst26316 (P3_U4915, P3_U4912, P3_U4913, P3_U4914);
  nand ginst26317 (P3_U4916, P3_R1054_U74, P3_U3051);
  nand ginst26318 (P3_U4917, P3_U3403, P3_U5768);
  nand ginst26319 (P3_U4918, P3_U3042, P3_U4915);
  nand ginst26320 (P3_U4919, P3_R1212_U53, P3_U3041);
  nand ginst26321 (P3_U4920, P3_REG3_REG_5__SCAN_IN, P3_U3151);
  nand ginst26322 (P3_U4921, P3_R1209_U53, P3_U3038);
  nand ginst26323 (P3_U4922, P3_ADDR_REG_5__SCAN_IN, P3_U4760);
  nand ginst26324 (P3_U4923, P3_R1212_U54, P3_U3040);
  nand ginst26325 (P3_U4924, P3_U3039, P3_U3400);
  nand ginst26326 (P3_U4925, P3_R1209_U54, P3_U3037);
  nand ginst26327 (P3_U4926, P3_U4923, P3_U4924, P3_U4925);
  nand ginst26328 (P3_U4927, P3_R1054_U75, P3_U3051);
  nand ginst26329 (P3_U4928, P3_U3400, P3_U5768);
  nand ginst26330 (P3_U4929, P3_U3042, P3_U4926);
  nand ginst26331 (P3_U4930, P3_R1212_U54, P3_U3041);
  nand ginst26332 (P3_U4931, P3_REG3_REG_4__SCAN_IN, P3_U3151);
  nand ginst26333 (P3_U4932, P3_R1209_U54, P3_U3038);
  nand ginst26334 (P3_U4933, P3_ADDR_REG_4__SCAN_IN, P3_U4760);
  nand ginst26335 (P3_U4934, P3_R1212_U55, P3_U3040);
  nand ginst26336 (P3_U4935, P3_U3039, P3_U3397);
  nand ginst26337 (P3_U4936, P3_R1209_U55, P3_U3037);
  nand ginst26338 (P3_U4937, P3_U4934, P3_U4935, P3_U4936);
  nand ginst26339 (P3_U4938, P3_R1054_U14, P3_U3051);
  nand ginst26340 (P3_U4939, P3_U3397, P3_U5768);
  nand ginst26341 (P3_U4940, P3_U3042, P3_U4937);
  nand ginst26342 (P3_U4941, P3_R1212_U55, P3_U3041);
  nand ginst26343 (P3_U4942, P3_REG3_REG_3__SCAN_IN, P3_U3151);
  nand ginst26344 (P3_U4943, P3_R1209_U55, P3_U3038);
  nand ginst26345 (P3_U4944, P3_ADDR_REG_3__SCAN_IN, P3_U4760);
  nand ginst26346 (P3_U4945, P3_R1212_U56, P3_U3040);
  nand ginst26347 (P3_U4946, P3_U3039, P3_U3394);
  nand ginst26348 (P3_U4947, P3_R1209_U56, P3_U3037);
  nand ginst26349 (P3_U4948, P3_U4945, P3_U4946, P3_U4947);
  nand ginst26350 (P3_U4949, P3_R1054_U76, P3_U3051);
  nand ginst26351 (P3_U4950, P3_U3394, P3_U5768);
  nand ginst26352 (P3_U4951, P3_U3042, P3_U4948);
  nand ginst26353 (P3_U4952, P3_R1212_U56, P3_U3041);
  nand ginst26354 (P3_U4953, P3_REG3_REG_2__SCAN_IN, P3_U3151);
  nand ginst26355 (P3_U4954, P3_R1209_U56, P3_U3038);
  nand ginst26356 (P3_U4955, P3_ADDR_REG_2__SCAN_IN, P3_U4760);
  nand ginst26357 (P3_U4956, P3_R1212_U57, P3_U3040);
  nand ginst26358 (P3_U4957, P3_U3039, P3_U3391);
  nand ginst26359 (P3_U4958, P3_R1209_U57, P3_U3037);
  nand ginst26360 (P3_U4959, P3_U4956, P3_U4957, P3_U4958);
  nand ginst26361 (P3_U4960, P3_R1054_U66, P3_U3051);
  nand ginst26362 (P3_U4961, P3_U3391, P3_U5768);
  nand ginst26363 (P3_U4962, P3_U3042, P3_U4959);
  nand ginst26364 (P3_U4963, P3_R1212_U57, P3_U3041);
  nand ginst26365 (P3_U4964, P3_REG3_REG_1__SCAN_IN, P3_U3151);
  nand ginst26366 (P3_U4965, P3_R1209_U57, P3_U3038);
  nand ginst26367 (P3_U4966, P3_ADDR_REG_1__SCAN_IN, P3_U4760);
  nand ginst26368 (P3_U4967, P3_R1212_U7, P3_U3040);
  nand ginst26369 (P3_U4968, P3_U3039, P3_U3386);
  nand ginst26370 (P3_U4969, P3_R1209_U7, P3_U3037);
  nand ginst26371 (P3_U4970, P3_U4967, P3_U4968, P3_U4969);
  nand ginst26372 (P3_U4971, P3_R1054_U17, P3_U3051);
  nand ginst26373 (P3_U4972, P3_U3386, P3_U5768);
  nand ginst26374 (P3_U4973, P3_U3042, P3_U4970);
  nand ginst26375 (P3_U4974, P3_R1212_U7, P3_U3041);
  nand ginst26376 (P3_U4975, P3_REG3_REG_0__SCAN_IN, P3_U3151);
  nand ginst26377 (P3_U4976, P3_R1209_U7, P3_U3038);
  nand ginst26378 (P3_U4977, P3_ADDR_REG_0__SCAN_IN, P3_U4760);
  not ginst26379 (P3_U4978, P3_U3868);
  nand ginst26380 (P3_U4979, P3_U3050, P3_U5941, P3_U5942);
  nand ginst26381 (P3_U4980, P3_U3023, P3_U3867, P3_U3909);
  nand ginst26382 (P3_U4981, P3_B_REG_SCAN_IN, P3_U4979);
  nand ginst26383 (P3_U4982, P3_U3036, P3_U3078);
  nand ginst26384 (P3_U4983, P3_U3032, P3_U3072);
  nand ginst26385 (P3_U4984, P3_SUB_609_U21, P3_U3304);
  nand ginst26386 (P3_U4985, P3_U4982, P3_U4983, P3_U4984);
  nand ginst26387 (P3_U4986, P3_U3311, P3_U3312, P3_U3875, P3_U3888, P3_U5425);
  nand ginst26388 (P3_U4987, P3_U3894, P3_U4986);
  nand ginst26389 (P3_U4988, P3_U3889, P3_U3895);
  nand ginst26390 (P3_U4989, P3_U4987, P3_U4988);
  nand ginst26391 (P3_U4990, P3_U3378, P3_U3911);
  nand ginst26392 (P3_U4991, P3_U3304, P3_U3889);
  nand ginst26393 (P3_U4992, P3_U3303, P3_U4986);
  not ginst26394 (P3_U4993, P3_U3370);
  nand ginst26395 (P3_U4994, P3_U3434, P3_U5420);
  nand ginst26396 (P3_U4995, P3_SUB_609_U21, P3_U3371);
  nand ginst26397 (P3_U4996, P3_R1158_U114, P3_U3035);
  nand ginst26398 (P3_U4997, P3_U3031, P3_U4985);
  nand ginst26399 (P3_U4998, P3_REG3_REG_15__SCAN_IN, P3_U3151);
  nand ginst26400 (P3_U4999, P3_U3036, P3_U3057);
  nand ginst26401 (P3_U5000, P3_U3032, P3_U3052);
  nand ginst26402 (P3_U5001, P3_SUB_609_U26, P3_U3304);
  nand ginst26403 (P3_U5002, P3_U4999, P3_U5000, P3_U5001);
  nand ginst26404 (P3_U5003, P3_U3303, P3_U3365);
  nand ginst26405 (P3_U5004, P3_U4993, P3_U5003);
  nand ginst26406 (P3_U5005, P3_U3365, P3_U3894);
  nand ginst26407 (P3_U5006, P3_U3360, P3_U5005);
  nand ginst26408 (P3_U5007, P3_U3045, P3_U3901);
  nand ginst26409 (P3_U5008, P3_SUB_609_U26, P3_U3044);
  nand ginst26410 (P3_U5009, P3_R1158_U16, P3_U3035);
  nand ginst26411 (P3_U5010, P3_U3031, P3_U5002);
  nand ginst26412 (P3_U5011, P3_REG3_REG_26__SCAN_IN, P3_U3151);
  nand ginst26413 (P3_U5012, P3_U3036, P3_U3066);
  nand ginst26414 (P3_U5013, P3_U3032, P3_U3069);
  nand ginst26415 (P3_U5014, P3_SUB_609_U8, P3_U3304);
  nand ginst26416 (P3_U5015, P3_U5012, P3_U5013, P3_U5014);
  nand ginst26417 (P3_U5016, P3_U3407, P3_U5420);
  nand ginst26418 (P3_U5017, P3_SUB_609_U8, P3_U3371);
  nand ginst26419 (P3_U5018, P3_R1158_U97, P3_U3035);
  nand ginst26420 (P3_U5019, P3_U3031, P3_U5015);
  nand ginst26421 (P3_U5020, P3_REG3_REG_6__SCAN_IN, P3_U3151);
  nand ginst26422 (P3_U5021, P3_U3036, P3_U3068);
  nand ginst26423 (P3_U5022, P3_U3032, P3_U3080);
  nand ginst26424 (P3_U5023, P3_SUB_609_U11, P3_U3304);
  nand ginst26425 (P3_U5024, P3_U5021, P3_U5022, P3_U5023);
  nand ginst26426 (P3_U5025, P3_U3443, P3_U5420);
  nand ginst26427 (P3_U5026, P3_SUB_609_U11, P3_U3371);
  nand ginst26428 (P3_U5027, P3_R1158_U112, P3_U3035);
  nand ginst26429 (P3_U5028, P3_U3031, P3_U5024);
  nand ginst26430 (P3_U5029, P3_REG3_REG_18__SCAN_IN, P3_U3151);
  nand ginst26431 (P3_U5030, P3_U3036, P3_U3077);
  nand ginst26432 (P3_U5031, P3_U3032, P3_U3063);
  nand ginst26433 (P3_U5032, P3_REG3_REG_2__SCAN_IN, P3_U3304);
  nand ginst26434 (P3_U5033, P3_U5030, P3_U5031, P3_U5032);
  nand ginst26435 (P3_U5034, P3_U3395, P3_U5420);
  nand ginst26436 (P3_U5035, P3_REG3_REG_2__SCAN_IN, P3_U3371);
  nand ginst26437 (P3_U5036, P3_R1158_U100, P3_U3035);
  nand ginst26438 (P3_U5037, P3_U3031, P3_U5033);
  nand ginst26439 (P3_U5038, P3_REG3_REG_2__SCAN_IN, P3_U3151);
  nand ginst26440 (P3_U5039, P3_U3036, P3_U3061);
  nand ginst26441 (P3_U5040, P3_U3032, P3_U3071);
  nand ginst26442 (P3_U5041, P3_SUB_609_U9, P3_U3304);
  nand ginst26443 (P3_U5042, P3_U5039, P3_U5040, P3_U5041);
  nand ginst26444 (P3_U5043, P3_U3422, P3_U5420);
  nand ginst26445 (P3_U5044, P3_SUB_609_U9, P3_U3371);
  nand ginst26446 (P3_U5045, P3_R1158_U117, P3_U3035);
  nand ginst26447 (P3_U5046, P3_U3031, P3_U5042);
  nand ginst26448 (P3_U5047, P3_REG3_REG_11__SCAN_IN, P3_U3151);
  nand ginst26449 (P3_U5048, P3_U3036, P3_U3074);
  nand ginst26450 (P3_U5049, P3_U3032, P3_U3065);
  nand ginst26451 (P3_U5050, P3_SUB_609_U17, P3_U3304);
  nand ginst26452 (P3_U5051, P3_U5048, P3_U5049, P3_U5050);
  nand ginst26453 (P3_U5052, P3_U3045, P3_U3905);
  nand ginst26454 (P3_U5053, P3_SUB_609_U17, P3_U3044);
  nand ginst26455 (P3_U5054, P3_R1158_U108, P3_U3035);
  nand ginst26456 (P3_U5055, P3_U3031, P3_U5051);
  nand ginst26457 (P3_U5056, P3_REG3_REG_22__SCAN_IN, P3_U3151);
  nand ginst26458 (P3_U5057, P3_U3036, P3_U3071);
  nand ginst26459 (P3_U5058, P3_U3032, P3_U3078);
  nand ginst26460 (P3_U5059, P3_SUB_609_U24, P3_U3304);
  nand ginst26461 (P3_U5060, P3_U5057, P3_U5058, P3_U5059);
  nand ginst26462 (P3_U5061, P3_U3428, P3_U5420);
  nand ginst26463 (P3_U5062, P3_SUB_609_U24, P3_U3371);
  nand ginst26464 (P3_U5063, P3_R1158_U13, P3_U3035);
  nand ginst26465 (P3_U5064, P3_U3031, P3_U5060);
  nand ginst26466 (P3_U5065, P3_REG3_REG_13__SCAN_IN, P3_U3151);
  nand ginst26467 (P3_U5066, P3_U3036, P3_U3080);
  nand ginst26468 (P3_U5067, P3_U3032, P3_U3074);
  nand ginst26469 (P3_U5068, P3_SUB_609_U20, P3_U3304);
  nand ginst26470 (P3_U5069, P3_U5066, P3_U5067, P3_U5068);
  nand ginst26471 (P3_U5070, P3_U3045, P3_U3907);
  nand ginst26472 (P3_U5071, P3_SUB_609_U20, P3_U3044);
  nand ginst26473 (P3_U5072, P3_R1158_U109, P3_U3035);
  nand ginst26474 (P3_U5073, P3_U3031, P3_U5069);
  nand ginst26475 (P3_U5074, P3_REG3_REG_20__SCAN_IN, P3_U3151);
  nand ginst26476 (P3_U5075, P3_U3031, P3_U3304);
  nand ginst26477 (P3_U5076, P3_U5075, P3_U5419);
  nand ginst26478 (P3_U5077, P3_U3032, P3_U3787);
  nand ginst26479 (P3_U5078, P3_U3387, P3_U5420);
  nand ginst26480 (P3_U5079, P3_REG3_REG_0__SCAN_IN, P3_U5076);
  nand ginst26481 (P3_U5080, P3_R1158_U94, P3_U3035);
  nand ginst26482 (P3_U5081, P3_REG3_REG_0__SCAN_IN, P3_U3151);
  nand ginst26483 (P3_U5082, P3_U3036, P3_U3083);
  nand ginst26484 (P3_U5083, P3_U3032, P3_U3061);
  nand ginst26485 (P3_U5084, P3_SUB_609_U14, P3_U3304);
  nand ginst26486 (P3_U5085, P3_U5082, P3_U5083, P3_U5084);
  nand ginst26487 (P3_U5086, P3_U3416, P3_U5420);
  nand ginst26488 (P3_U5087, P3_SUB_609_U14, P3_U3371);
  nand ginst26489 (P3_U5088, P3_R1158_U95, P3_U3035);
  nand ginst26490 (P3_U5089, P3_U3031, P3_U5085);
  nand ginst26491 (P3_U5090, P3_REG3_REG_9__SCAN_IN, P3_U3151);
  nand ginst26492 (P3_U5091, P3_U3036, P3_U3063);
  nand ginst26493 (P3_U5092, P3_U3032, P3_U3066);
  nand ginst26494 (P3_U5093, P3_SUB_609_U29, P3_U3304);
  nand ginst26495 (P3_U5094, P3_U5091, P3_U5092, P3_U5093);
  nand ginst26496 (P3_U5095, P3_U3401, P3_U5420);
  nand ginst26497 (P3_U5096, P3_SUB_609_U29, P3_U3371);
  nand ginst26498 (P3_U5097, P3_R1158_U99, P3_U3035);
  nand ginst26499 (P3_U5098, P3_U3031, P3_U5094);
  nand ginst26500 (P3_U5099, P3_REG3_REG_4__SCAN_IN, P3_U3151);
  nand ginst26501 (P3_U5100, P3_U3036, P3_U3065);
  nand ginst26502 (P3_U5101, P3_U3032, P3_U3057);
  nand ginst26503 (P3_U5102, P3_SUB_609_U10, P3_U3304);
  nand ginst26504 (P3_U5103, P3_U5100, P3_U5101, P3_U5102);
  nand ginst26505 (P3_U5104, P3_U3045, P3_U3903);
  nand ginst26506 (P3_U5105, P3_SUB_609_U10, P3_U3044);
  nand ginst26507 (P3_U5106, P3_R1158_U106, P3_U3035);
  nand ginst26508 (P3_U5107, P3_U3031, P3_U5103);
  nand ginst26509 (P3_U5108, P3_REG3_REG_24__SCAN_IN, P3_U3151);
  nand ginst26510 (P3_U5109, P3_U3036, P3_U3072);
  nand ginst26511 (P3_U5110, P3_U3032, P3_U3081);
  nand ginst26512 (P3_U5111, P3_SUB_609_U19, P3_U3304);
  nand ginst26513 (P3_U5112, P3_U5109, P3_U5110, P3_U5111);
  nand ginst26514 (P3_U5113, P3_U3440, P3_U5420);
  nand ginst26515 (P3_U5114, P3_SUB_609_U19, P3_U3371);
  nand ginst26516 (P3_U5115, P3_R1158_U14, P3_U3035);
  nand ginst26517 (P3_U5116, P3_U3031, P3_U5112);
  nand ginst26518 (P3_U5117, P3_REG3_REG_17__SCAN_IN, P3_U3151);
  nand ginst26519 (P3_U5118, P3_U3036, P3_U3059);
  nand ginst26520 (P3_U5119, P3_U3032, P3_U3070);
  nand ginst26521 (P3_U5120, P3_SUB_609_U53, P3_U3304);
  nand ginst26522 (P3_U5121, P3_U5118, P3_U5119, P3_U5120);
  nand ginst26523 (P3_U5122, P3_U3404, P3_U5420);
  nand ginst26524 (P3_U5123, P3_SUB_609_U53, P3_U3371);
  nand ginst26525 (P3_U5124, P3_R1158_U98, P3_U3035);
  nand ginst26526 (P3_U5125, P3_U3031, P3_U5121);
  nand ginst26527 (P3_U5126, P3_REG3_REG_5__SCAN_IN, P3_U3151);
  nand ginst26528 (P3_U5127, P3_U3036, P3_U3073);
  nand ginst26529 (P3_U5128, P3_U3032, P3_U3068);
  nand ginst26530 (P3_U5129, P3_SUB_609_U7, P3_U3304);
  nand ginst26531 (P3_U5130, P3_U5127, P3_U5128, P3_U5129);
  nand ginst26532 (P3_U5131, P3_U3437, P3_U5420);
  nand ginst26533 (P3_U5132, P3_SUB_609_U7, P3_U3371);
  nand ginst26534 (P3_U5133, P3_R1158_U113, P3_U3035);
  nand ginst26535 (P3_U5134, P3_U3031, P3_U5130);
  nand ginst26536 (P3_U5135, P3_REG3_REG_16__SCAN_IN, P3_U3151);
  nand ginst26537 (P3_U5136, P3_U3036, P3_U3064);
  nand ginst26538 (P3_U5137, P3_U3032, P3_U3056);
  nand ginst26539 (P3_U5138, P3_SUB_609_U16, P3_U3304);
  nand ginst26540 (P3_U5139, P3_U5136, P3_U5137, P3_U5138);
  nand ginst26541 (P3_U5140, P3_U3045, P3_U3902);
  nand ginst26542 (P3_U5141, P3_SUB_609_U16, P3_U3044);
  nand ginst26543 (P3_U5142, P3_R1158_U105, P3_U3035);
  nand ginst26544 (P3_U5143, P3_U3031, P3_U5139);
  nand ginst26545 (P3_U5144, P3_REG3_REG_25__SCAN_IN, P3_U3151);
  nand ginst26546 (P3_U5145, P3_U3036, P3_U3062);
  nand ginst26547 (P3_U5146, P3_U3032, P3_U3079);
  nand ginst26548 (P3_U5147, P3_SUB_609_U23, P3_U3304);
  nand ginst26549 (P3_U5148, P3_U5145, P3_U5146, P3_U5147);
  nand ginst26550 (P3_U5149, P3_U3425, P3_U5420);
  nand ginst26551 (P3_U5150, P3_SUB_609_U23, P3_U3371);
  nand ginst26552 (P3_U5151, P3_R1158_U116, P3_U3035);
  nand ginst26553 (P3_U5152, P3_U3031, P3_U5148);
  nand ginst26554 (P3_U5153, P3_REG3_REG_12__SCAN_IN, P3_U3151);
  nand ginst26555 (P3_U5154, P3_U3036, P3_U3075);
  nand ginst26556 (P3_U5155, P3_U3032, P3_U3060);
  nand ginst26557 (P3_U5156, P3_SUB_609_U27, P3_U3304);
  nand ginst26558 (P3_U5157, P3_U5154, P3_U5155, P3_U5156);
  nand ginst26559 (P3_U5158, P3_U3045, P3_U3906);
  nand ginst26560 (P3_U5159, P3_SUB_609_U27, P3_U3044);
  nand ginst26561 (P3_U5160, P3_R1158_U15, P3_U3035);
  nand ginst26562 (P3_U5161, P3_U3031, P3_U5157);
  nand ginst26563 (P3_U5162, P3_REG3_REG_21__SCAN_IN, P3_U3151);
  nand ginst26564 (P3_U5163, P3_U3036, P3_U3076);
  nand ginst26565 (P3_U5164, P3_U3032, P3_U3067);
  nand ginst26566 (P3_U5165, P3_REG3_REG_1__SCAN_IN, P3_U3304);
  nand ginst26567 (P3_U5166, P3_U5163, P3_U5164, P3_U5165);
  nand ginst26568 (P3_U5167, P3_U3392, P3_U5420);
  nand ginst26569 (P3_U5168, P3_REG3_REG_1__SCAN_IN, P3_U3371);
  nand ginst26570 (P3_U5169, P3_R1158_U110, P3_U3035);
  nand ginst26571 (P3_U5170, P3_U3031, P3_U5166);
  nand ginst26572 (P3_U5171, P3_REG3_REG_1__SCAN_IN, P3_U3151);
  nand ginst26573 (P3_U5172, P3_U3036, P3_U3069);
  nand ginst26574 (P3_U5173, P3_U3032, P3_U3082);
  nand ginst26575 (P3_U5174, P3_SUB_609_U12, P3_U3304);
  nand ginst26576 (P3_U5175, P3_U5172, P3_U5173, P3_U5174);
  nand ginst26577 (P3_U5176, P3_U3413, P3_U5420);
  nand ginst26578 (P3_U5177, P3_SUB_609_U12, P3_U3371);
  nand ginst26579 (P3_U5178, P3_R1158_U96, P3_U3035);
  nand ginst26580 (P3_U5179, P3_U3031, P3_U5175);
  nand ginst26581 (P3_U5180, P3_REG3_REG_8__SCAN_IN, P3_U3151);
  nand ginst26582 (P3_U5181, P3_U3036, P3_U3052);
  nand ginst26583 (P3_U5182, P3_U3032, P3_U3054);
  nand ginst26584 (P3_U5183, P3_SUB_609_U28, P3_U3304);
  nand ginst26585 (P3_U5184, P3_U5181, P3_U5182, P3_U5183);
  nand ginst26586 (P3_U5185, P3_U3045, P3_U3899);
  nand ginst26587 (P3_U5186, P3_SUB_609_U28, P3_U3044);
  nand ginst26588 (P3_U5187, P3_R1158_U101, P3_U3035);
  nand ginst26589 (P3_U5188, P3_U3031, P3_U5184);
  nand ginst26590 (P3_U5189, P3_REG3_REG_28__SCAN_IN, P3_U3151);
  nand ginst26591 (P3_U5190, P3_U3036, P3_U3081);
  nand ginst26592 (P3_U5191, P3_U3032, P3_U3075);
  nand ginst26593 (P3_U5192, P3_SUB_609_U15, P3_U3304);
  nand ginst26594 (P3_U5193, P3_U5190, P3_U5191, P3_U5192);
  nand ginst26595 (P3_U5194, P3_U3445, P3_U5420);
  nand ginst26596 (P3_U5195, P3_SUB_609_U15, P3_U3371);
  nand ginst26597 (P3_U5196, P3_R1158_U111, P3_U3035);
  nand ginst26598 (P3_U5197, P3_U3031, P3_U5193);
  nand ginst26599 (P3_U5198, P3_REG3_REG_19__SCAN_IN, P3_U3151);
  nand ginst26600 (P3_U5199, P3_U3036, P3_U3067);
  nand ginst26601 (P3_U5200, P3_U3032, P3_U3059);
  nand ginst26602 (P3_U5201, P3_SUB_609_U25, P3_U3304);
  nand ginst26603 (P3_U5202, P3_U5199, P3_U5200, P3_U5201);
  nand ginst26604 (P3_U5203, P3_U3398, P3_U5420);
  nand ginst26605 (P3_U5204, P3_SUB_609_U25, P3_U3371);
  nand ginst26606 (P3_U5205, P3_R1158_U17, P3_U3035);
  nand ginst26607 (P3_U5206, P3_U3031, P3_U5202);
  nand ginst26608 (P3_U5207, P3_REG3_REG_3__SCAN_IN, P3_U3151);
  nand ginst26609 (P3_U5208, P3_U3036, P3_U3082);
  nand ginst26610 (P3_U5209, P3_U3032, P3_U3062);
  nand ginst26611 (P3_U5210, P3_SUB_609_U13, P3_U3304);
  nand ginst26612 (P3_U5211, P3_U5208, P3_U5209, P3_U5210);
  nand ginst26613 (P3_U5212, P3_U3419, P3_U5420);
  nand ginst26614 (P3_U5213, P3_SUB_609_U13, P3_U3371);
  nand ginst26615 (P3_U5214, P3_R1158_U118, P3_U3035);
  nand ginst26616 (P3_U5215, P3_U3031, P3_U5211);
  nand ginst26617 (P3_U5216, P3_REG3_REG_10__SCAN_IN, P3_U3151);
  nand ginst26618 (P3_U5217, P3_U3036, P3_U3060);
  nand ginst26619 (P3_U5218, P3_U3032, P3_U3064);
  nand ginst26620 (P3_U5219, P3_SUB_609_U6, P3_U3304);
  nand ginst26621 (P3_U5220, P3_U5217, P3_U5218, P3_U5219);
  nand ginst26622 (P3_U5221, P3_U3045, P3_U3904);
  nand ginst26623 (P3_U5222, P3_SUB_609_U6, P3_U3044);
  nand ginst26624 (P3_U5223, P3_R1158_U107, P3_U3035);
  nand ginst26625 (P3_U5224, P3_U3031, P3_U5220);
  nand ginst26626 (P3_U5225, P3_REG3_REG_23__SCAN_IN, P3_U3151);
  nand ginst26627 (P3_U5226, P3_U3036, P3_U3079);
  nand ginst26628 (P3_U5227, P3_U3032, P3_U3073);
  nand ginst26629 (P3_U5228, P3_SUB_609_U30, P3_U3304);
  nand ginst26630 (P3_U5229, P3_U5226, P3_U5227, P3_U5228);
  nand ginst26631 (P3_U5230, P3_U3431, P3_U5420);
  nand ginst26632 (P3_U5231, P3_SUB_609_U30, P3_U3371);
  nand ginst26633 (P3_U5232, P3_R1158_U115, P3_U3035);
  nand ginst26634 (P3_U5233, P3_U3031, P3_U5229);
  nand ginst26635 (P3_U5234, P3_REG3_REG_14__SCAN_IN, P3_U3151);
  nand ginst26636 (P3_U5235, P3_U3036, P3_U3056);
  nand ginst26637 (P3_U5236, P3_U3032, P3_U3053);
  nand ginst26638 (P3_U5237, P3_SUB_609_U22, P3_U3304);
  nand ginst26639 (P3_U5238, P3_U5235, P3_U5236, P3_U5237);
  nand ginst26640 (P3_U5239, P3_U3045, P3_U3900);
  nand ginst26641 (P3_U5240, P3_SUB_609_U22, P3_U3044);
  nand ginst26642 (P3_U5241, P3_R1158_U102, P3_U3035);
  nand ginst26643 (P3_U5242, P3_U3031, P3_U5238);
  nand ginst26644 (P3_U5243, P3_REG3_REG_27__SCAN_IN, P3_U3151);
  nand ginst26645 (P3_U5244, P3_U3036, P3_U3070);
  nand ginst26646 (P3_U5245, P3_U3032, P3_U3083);
  nand ginst26647 (P3_U5246, P3_SUB_609_U18, P3_U3304);
  nand ginst26648 (P3_U5247, P3_U5244, P3_U5245, P3_U5246);
  nand ginst26649 (P3_U5248, P3_U3410, P3_U5420);
  nand ginst26650 (P3_U5249, P3_SUB_609_U18, P3_U3371);
  nand ginst26651 (P3_U5250, P3_R1158_U18, P3_U3035);
  nand ginst26652 (P3_U5251, P3_U3031, P3_U5247);
  nand ginst26653 (P3_U5252, P3_REG3_REG_7__SCAN_IN, P3_U3151);
  nand ginst26654 (P3_U5253, P3_U3046, P3_U3898);
  nand ginst26655 (P3_U5254, P3_U3375, P3_U3833);
  nand ginst26656 (P3_U5255, P3_U3815, P3_U3816);
  nand ginst26657 (P3_U5256, P3_U3013, P3_U3814);
  nand ginst26658 (P3_U5257, P3_U3880, P3_U5256);
  nand ginst26659 (P3_U5258, P3_U3416, P3_U5257);
  nand ginst26660 (P3_U5259, P3_U3082, P3_U5255);
  nand ginst26661 (P3_U5260, P3_U3413, P3_U5257);
  nand ginst26662 (P3_U5261, P3_U3083, P3_U5255);
  nand ginst26663 (P3_U5262, P3_U3410, P3_U5257);
  nand ginst26664 (P3_U5263, P3_U3069, P3_U5255);
  nand ginst26665 (P3_U5264, P3_U3407, P3_U5257);
  nand ginst26666 (P3_U5265, P3_U3070, P3_U5255);
  nand ginst26667 (P3_U5266, P3_U3404, P3_U5257);
  nand ginst26668 (P3_U5267, P3_U3066, P3_U5255);
  nand ginst26669 (P3_U5268, P3_U3401, P3_U5257);
  nand ginst26670 (P3_U5269, P3_U3059, P3_U5255);
  nand ginst26671 (P3_U5270, P3_U3872, P3_U5257);
  nand ginst26672 (P3_U5271, P3_U3055, P3_U5255);
  nand ginst26673 (P3_U5272, P3_U3873, P3_U5257);
  nand ginst26674 (P3_U5273, P3_U3058, P3_U5255);
  nand ginst26675 (P3_U5274, P3_U3398, P3_U5257);
  nand ginst26676 (P3_U5275, P3_U3063, P3_U5255);
  nand ginst26677 (P3_U5276, P3_U3908, P3_U5257);
  nand ginst26678 (P3_U5277, P3_U3054, P3_U5255);
  nand ginst26679 (P3_U5278, P3_U3899, P3_U5257);
  nand ginst26680 (P3_U5279, P3_U3053, P3_U5255);
  nand ginst26681 (P3_U5280, P3_U3900, P3_U5257);
  nand ginst26682 (P3_U5281, P3_U3052, P3_U5255);
  nand ginst26683 (P3_U5282, P3_U3901, P3_U5257);
  nand ginst26684 (P3_U5283, P3_U3056, P3_U5255);
  nand ginst26685 (P3_U5284, P3_U3902, P3_U5257);
  nand ginst26686 (P3_U5285, P3_U3057, P3_U5255);
  nand ginst26687 (P3_U5286, P3_U3903, P3_U5257);
  nand ginst26688 (P3_U5287, P3_U3064, P3_U5255);
  nand ginst26689 (P3_U5288, P3_U3904, P3_U5257);
  nand ginst26690 (P3_U5289, P3_U3065, P3_U5255);
  nand ginst26691 (P3_U5290, P3_U3905, P3_U5257);
  nand ginst26692 (P3_U5291, P3_U3060, P3_U5255);
  nand ginst26693 (P3_U5292, P3_U3906, P3_U5257);
  nand ginst26694 (P3_U5293, P3_U3074, P3_U5255);
  nand ginst26695 (P3_U5294, P3_U3907, P3_U5257);
  nand ginst26696 (P3_U5295, P3_U3075, P3_U5255);
  nand ginst26697 (P3_U5296, P3_U3395, P3_U5257);
  nand ginst26698 (P3_U5297, P3_U3067, P3_U5255);
  nand ginst26699 (P3_U5298, P3_U3445, P3_U5257);
  nand ginst26700 (P3_U5299, P3_U3080, P3_U5255);
  nand ginst26701 (P3_U5300, P3_U3443, P3_U5257);
  nand ginst26702 (P3_U5301, P3_U3081, P3_U5255);
  nand ginst26703 (P3_U5302, P3_U3440, P3_U5257);
  nand ginst26704 (P3_U5303, P3_U3068, P3_U5255);
  nand ginst26705 (P3_U5304, P3_U3437, P3_U5257);
  nand ginst26706 (P3_U5305, P3_U3072, P3_U5255);
  nand ginst26707 (P3_U5306, P3_U3434, P3_U5257);
  nand ginst26708 (P3_U5307, P3_U3073, P3_U5255);
  nand ginst26709 (P3_U5308, P3_U3431, P3_U5257);
  nand ginst26710 (P3_U5309, P3_U3078, P3_U5255);
  nand ginst26711 (P3_U5310, P3_U3428, P3_U5257);
  nand ginst26712 (P3_U5311, P3_U3079, P3_U5255);
  nand ginst26713 (P3_U5312, P3_U3425, P3_U5257);
  nand ginst26714 (P3_U5313, P3_U3071, P3_U5255);
  nand ginst26715 (P3_U5314, P3_U3422, P3_U5257);
  nand ginst26716 (P3_U5315, P3_U3062, P3_U5255);
  nand ginst26717 (P3_U5316, P3_U3419, P3_U5257);
  nand ginst26718 (P3_U5317, P3_U3061, P3_U5255);
  nand ginst26719 (P3_U5318, P3_U3392, P3_U5257);
  nand ginst26720 (P3_U5319, P3_U3077, P3_U5255);
  nand ginst26721 (P3_U5320, P3_U3387, P3_U5257);
  nand ginst26722 (P3_U5321, P3_U3076, P3_U5255);
  nand ginst26723 (P3_U5322, P3_U3416, P3_U5255);
  nand ginst26724 (P3_U5323, P3_U3082, P3_U5257);
  nand ginst26725 (P3_U5324, P3_U3083, P3_U5440);
  nand ginst26726 (P3_U5325, P3_U3413, P3_U5255);
  nand ginst26727 (P3_U5326, P3_U3083, P3_U5257);
  nand ginst26728 (P3_U5327, P3_U3069, P3_U5440);
  nand ginst26729 (P3_U5328, P3_U3410, P3_U5255);
  nand ginst26730 (P3_U5329, P3_U3069, P3_U5257);
  nand ginst26731 (P3_U5330, P3_U3070, P3_U5440);
  nand ginst26732 (P3_U5331, P3_U3407, P3_U5255);
  nand ginst26733 (P3_U5332, P3_U3070, P3_U5257);
  nand ginst26734 (P3_U5333, P3_U3066, P3_U5440);
  nand ginst26735 (P3_U5334, P3_U3404, P3_U5255);
  nand ginst26736 (P3_U5335, P3_U3066, P3_U5257);
  nand ginst26737 (P3_U5336, P3_U3059, P3_U5440);
  nand ginst26738 (P3_U5337, P3_U3401, P3_U5255);
  nand ginst26739 (P3_U5338, P3_U3059, P3_U5257);
  nand ginst26740 (P3_U5339, P3_U3063, P3_U5440);
  nand ginst26741 (P3_U5340, P3_U3055, P3_U5257);
  nand ginst26742 (P3_U5341, P3_U3872, P3_U5255);
  nand ginst26743 (P3_U5342, P3_U3058, P3_U5257);
  nand ginst26744 (P3_U5343, P3_U3873, P3_U5255);
  nand ginst26745 (P3_U5344, P3_U3398, P3_U5255);
  nand ginst26746 (P3_U5345, P3_U3063, P3_U5257);
  nand ginst26747 (P3_U5346, P3_U3067, P3_U5440);
  nand ginst26748 (P3_U5347, P3_U3054, P3_U5257);
  nand ginst26749 (P3_U5348, P3_U3908, P3_U5255);
  nand ginst26750 (P3_U5349, P3_U3053, P3_U5440);
  nand ginst26751 (P3_U5350, P3_U3053, P3_U5257);
  nand ginst26752 (P3_U5351, P3_U3899, P3_U5255);
  nand ginst26753 (P3_U5352, P3_U3052, P3_U5440);
  nand ginst26754 (P3_U5353, P3_U3052, P3_U5257);
  nand ginst26755 (P3_U5354, P3_U3900, P3_U5255);
  nand ginst26756 (P3_U5355, P3_U3056, P3_U5440);
  nand ginst26757 (P3_U5356, P3_U3056, P3_U5257);
  nand ginst26758 (P3_U5357, P3_U3901, P3_U5255);
  nand ginst26759 (P3_U5358, P3_U3057, P3_U5440);
  nand ginst26760 (P3_U5359, P3_U3057, P3_U5257);
  nand ginst26761 (P3_U5360, P3_U3902, P3_U5255);
  nand ginst26762 (P3_U5361, P3_U3064, P3_U5440);
  nand ginst26763 (P3_U5362, P3_U3064, P3_U5257);
  nand ginst26764 (P3_U5363, P3_U3903, P3_U5255);
  nand ginst26765 (P3_U5364, P3_U3065, P3_U5440);
  nand ginst26766 (P3_U5365, P3_U3065, P3_U5257);
  nand ginst26767 (P3_U5366, P3_U3904, P3_U5255);
  nand ginst26768 (P3_U5367, P3_U3060, P3_U5440);
  nand ginst26769 (P3_U5368, P3_U3060, P3_U5257);
  nand ginst26770 (P3_U5369, P3_U3905, P3_U5255);
  nand ginst26771 (P3_U5370, P3_U3074, P3_U5440);
  nand ginst26772 (P3_U5371, P3_U3074, P3_U5257);
  nand ginst26773 (P3_U5372, P3_U3906, P3_U5255);
  nand ginst26774 (P3_U5373, P3_U3075, P3_U5440);
  nand ginst26775 (P3_U5374, P3_U3075, P3_U5257);
  nand ginst26776 (P3_U5375, P3_U3907, P3_U5255);
  nand ginst26777 (P3_U5376, P3_U3080, P3_U5440);
  nand ginst26778 (P3_U5377, P3_U3395, P3_U5255);
  nand ginst26779 (P3_U5378, P3_U3067, P3_U5257);
  nand ginst26780 (P3_U5379, P3_U3077, P3_U5440);
  nand ginst26781 (P3_U5380, P3_U3445, P3_U5255);
  nand ginst26782 (P3_U5381, P3_U3080, P3_U5257);
  nand ginst26783 (P3_U5382, P3_U3081, P3_U5440);
  nand ginst26784 (P3_U5383, P3_U3443, P3_U5255);
  nand ginst26785 (P3_U5384, P3_U3081, P3_U5257);
  nand ginst26786 (P3_U5385, P3_U3068, P3_U5440);
  nand ginst26787 (P3_U5386, P3_U3440, P3_U5255);
  nand ginst26788 (P3_U5387, P3_U3068, P3_U5257);
  nand ginst26789 (P3_U5388, P3_U3072, P3_U5440);
  nand ginst26790 (P3_U5389, P3_U3437, P3_U5255);
  nand ginst26791 (P3_U5390, P3_U3072, P3_U5257);
  nand ginst26792 (P3_U5391, P3_U3073, P3_U5440);
  nand ginst26793 (P3_U5392, P3_U3434, P3_U5255);
  nand ginst26794 (P3_U5393, P3_U3073, P3_U5257);
  nand ginst26795 (P3_U5394, P3_U3078, P3_U5440);
  nand ginst26796 (P3_U5395, P3_U3431, P3_U5255);
  nand ginst26797 (P3_U5396, P3_U3078, P3_U5257);
  nand ginst26798 (P3_U5397, P3_U3079, P3_U5440);
  nand ginst26799 (P3_U5398, P3_U3428, P3_U5255);
  nand ginst26800 (P3_U5399, P3_U3079, P3_U5257);
  nand ginst26801 (P3_U5400, P3_U3071, P3_U5440);
  nand ginst26802 (P3_U5401, P3_U3425, P3_U5255);
  nand ginst26803 (P3_U5402, P3_U3071, P3_U5257);
  nand ginst26804 (P3_U5403, P3_U3062, P3_U5440);
  nand ginst26805 (P3_U5404, P3_U3422, P3_U5255);
  nand ginst26806 (P3_U5405, P3_U3062, P3_U5257);
  nand ginst26807 (P3_U5406, P3_U3061, P3_U5440);
  nand ginst26808 (P3_U5407, P3_U3419, P3_U5255);
  nand ginst26809 (P3_U5408, P3_U3061, P3_U5257);
  nand ginst26810 (P3_U5409, P3_U3082, P3_U5440);
  nand ginst26811 (P3_U5410, P3_U3392, P3_U5255);
  nand ginst26812 (P3_U5411, P3_U3077, P3_U5257);
  nand ginst26813 (P3_U5412, P3_U3076, P3_U5440);
  nand ginst26814 (P3_U5413, P3_U3387, P3_U5255);
  nand ginst26815 (P3_U5414, P3_U3076, P3_U5257);
  nand ginst26816 (P3_U5415, P3_U3151, P3_U4981);
  nand ginst26817 (P3_U5416, P3_U4980, P3_U4981, P3_U5440);
  nand ginst26818 (P3_U5417, P3_U3043, P3_U3303);
  nand ginst26819 (P3_U5418, P3_U3043, P3_U3894);
  not ginst26820 (P3_U5419, P3_U3371);
  nand ginst26821 (P3_U5420, P3_U3918, P3_U5418);
  nand ginst26822 (P3_U5421, P3_U3774, P3_U5937, P3_U5938);
  nand ginst26823 (P3_U5422, P3_U5428, P3_U5434);
  nand ginst26824 (P3_U5423, P3_U3378, P3_U3879);
  nand ginst26825 (P3_U5424, P3_U3375, P3_U3833);
  nand ginst26826 (P3_U5425, P3_U3876, P3_U5447);
  nand ginst26827 (P3_U5426, P3_IR_REG_24__SCAN_IN, P3_U3831);
  nand ginst26828 (P3_U5427, P3_IR_REG_31__SCAN_IN, P3_SUB_598_U18);
  not ginst26829 (P3_U5428, P3_U3372);
  nand ginst26830 (P3_U5429, P3_IR_REG_25__SCAN_IN, P3_U3831);
  nand ginst26831 (P3_U5430, P3_IR_REG_31__SCAN_IN, P3_SUB_598_U81);
  not ginst26832 (P3_U5431, P3_U3373);
  nand ginst26833 (P3_U5432, P3_IR_REG_26__SCAN_IN, P3_U3831);
  nand ginst26834 (P3_U5433, P3_IR_REG_31__SCAN_IN, P3_SUB_598_U19);
  not ginst26835 (P3_U5434, P3_U3374);
  nand ginst26836 (P3_U5435, P3_B_REG_SCAN_IN, P3_U5428);
  nand ginst26837 (P3_U5436, P3_U3298, P3_U3372);
  nand ginst26838 (P3_U5437, P3_U5435, P3_U5436);
  nand ginst26839 (P3_U5438, P3_IR_REG_23__SCAN_IN, P3_U3831);
  nand ginst26840 (P3_U5439, P3_IR_REG_31__SCAN_IN, P3_SUB_598_U17);
  not ginst26841 (P3_U5440, P3_U3375);
  nand ginst26842 (P3_U5441, P3_D_REG_0__SCAN_IN, P3_U3832);
  nand ginst26843 (P3_U5442, P3_U3915, P3_U4020);
  nand ginst26844 (P3_U5443, P3_D_REG_1__SCAN_IN, P3_U3832);
  nand ginst26845 (P3_U5444, P3_U3915, P3_U4021);
  nand ginst26846 (P3_U5445, P3_IR_REG_20__SCAN_IN, P3_U3831);
  nand ginst26847 (P3_U5446, P3_IR_REG_31__SCAN_IN, P3_SUB_598_U15);
  not ginst26848 (P3_U5447, P3_U3378);
  nand ginst26849 (P3_U5448, P3_IR_REG_19__SCAN_IN, P3_U3831);
  nand ginst26850 (P3_U5449, P3_IR_REG_31__SCAN_IN, P3_SUB_598_U14);
  not ginst26851 (P3_U5450, P3_U3379);
  nand ginst26852 (P3_U5451, P3_IR_REG_22__SCAN_IN, P3_U3831);
  nand ginst26853 (P3_U5452, P3_IR_REG_31__SCAN_IN, P3_SUB_598_U16);
  not ginst26854 (P3_U5453, P3_U3380);
  nand ginst26855 (P3_U5454, P3_IR_REG_21__SCAN_IN, P3_U3831);
  nand ginst26856 (P3_U5455, P3_IR_REG_31__SCAN_IN, P3_SUB_598_U83);
  not ginst26857 (P3_U5456, P3_U3385);
  nand ginst26858 (P3_U5457, P3_IR_REG_30__SCAN_IN, P3_U3831);
  nand ginst26859 (P3_U5458, P3_IR_REG_31__SCAN_IN, P3_SUB_598_U77);
  not ginst26860 (P3_U5459, P3_U3381);
  nand ginst26861 (P3_U5460, P3_IR_REG_29__SCAN_IN, P3_U3831);
  nand ginst26862 (P3_U5461, P3_IR_REG_31__SCAN_IN, P3_SUB_598_U21);
  not ginst26863 (P3_U5462, P3_U3382);
  nand ginst26864 (P3_U5463, P3_IR_REG_28__SCAN_IN, P3_U3831);
  nand ginst26865 (P3_U5464, P3_IR_REG_31__SCAN_IN, P3_SUB_598_U20);
  not ginst26866 (P3_U5465, P3_U3383);
  nand ginst26867 (P3_U5466, P3_IR_REG_27__SCAN_IN, P3_U3831);
  nand ginst26868 (P3_U5467, P3_IR_REG_31__SCAN_IN, P3_SUB_598_U79);
  not ginst26869 (P3_U5468, P3_U3384);
  nand ginst26870 (P3_U5469, P3_IR_REG_0__SCAN_IN, P3_U3831);
  nand ginst26871 (P3_U5470, P3_IR_REG_0__SCAN_IN, P3_IR_REG_31__SCAN_IN);
  nand ginst26872 (P3_U5471, P3_U3833, U61);
  nand ginst26873 (P3_U5472, P3_U3386, P3_U3893);
  not ginst26874 (P3_U5473, P3_U3387);
  nand ginst26875 (P3_U5474, P3_U3300, P3_U5422);
  nand ginst26876 (P3_U5475, P3_D_REG_0__SCAN_IN, P3_U4019);
  not ginst26877 (P3_U5476, P3_U3388);
  nand ginst26878 (P3_U5477, P3_D_REG_1__SCAN_IN, P3_U4019);
  nand ginst26879 (P3_U5478, P3_U3300, P3_U4021);
  not ginst26880 (P3_U5479, P3_U3389);
  nand ginst26881 (P3_U5480, P3_U4052, P3_U5453);
  nand ginst26882 (P3_U5481, P3_U3380, P3_U3834);
  nand ginst26883 (P3_U5482, P3_U5480, P3_U5481);
  nand ginst26884 (P3_U5483, P3_REG0_REG_0__SCAN_IN, P3_U3835);
  nand ginst26885 (P3_U5484, P3_U3914, P3_U4077);
  nand ginst26886 (P3_U5485, P3_IR_REG_1__SCAN_IN, P3_U3831);
  nand ginst26887 (P3_U5486, P3_IR_REG_31__SCAN_IN, P3_SUB_598_U51);
  nand ginst26888 (P3_U5487, P3_U3833, U50);
  nand ginst26889 (P3_U5488, P3_U3391, P3_U3893);
  not ginst26890 (P3_U5489, P3_U3392);
  nand ginst26891 (P3_U5490, P3_REG0_REG_1__SCAN_IN, P3_U3835);
  nand ginst26892 (P3_U5491, P3_U3914, P3_U4102);
  nand ginst26893 (P3_U5492, P3_IR_REG_2__SCAN_IN, P3_U3831);
  nand ginst26894 (P3_U5493, P3_IR_REG_31__SCAN_IN, P3_SUB_598_U22);
  nand ginst26895 (P3_U5494, P3_U3833, U39);
  nand ginst26896 (P3_U5495, P3_U3394, P3_U3893);
  not ginst26897 (P3_U5496, P3_U3395);
  nand ginst26898 (P3_U5497, P3_REG0_REG_2__SCAN_IN, P3_U3835);
  nand ginst26899 (P3_U5498, P3_U3914, P3_U4120);
  nand ginst26900 (P3_U5499, P3_IR_REG_3__SCAN_IN, P3_U3831);
  nand ginst26901 (P3_U5500, P3_IR_REG_31__SCAN_IN, P3_SUB_598_U23);
  nand ginst26902 (P3_U5501, P3_U3833, U36);
  nand ginst26903 (P3_U5502, P3_U3397, P3_U3893);
  not ginst26904 (P3_U5503, P3_U3398);
  nand ginst26905 (P3_U5504, P3_REG0_REG_3__SCAN_IN, P3_U3835);
  nand ginst26906 (P3_U5505, P3_U3914, P3_U4138);
  nand ginst26907 (P3_U5506, P3_IR_REG_4__SCAN_IN, P3_U3831);
  nand ginst26908 (P3_U5507, P3_IR_REG_31__SCAN_IN, P3_SUB_598_U24);
  nand ginst26909 (P3_U5508, P3_U3833, U35);
  nand ginst26910 (P3_U5509, P3_U3400, P3_U3893);
  not ginst26911 (P3_U5510, P3_U3401);
  nand ginst26912 (P3_U5511, P3_REG0_REG_4__SCAN_IN, P3_U3835);
  nand ginst26913 (P3_U5512, P3_U3914, P3_U4156);
  nand ginst26914 (P3_U5513, P3_IR_REG_5__SCAN_IN, P3_U3831);
  nand ginst26915 (P3_U5514, P3_IR_REG_31__SCAN_IN, P3_SUB_598_U74);
  nand ginst26916 (P3_U5515, P3_U3833, U34);
  nand ginst26917 (P3_U5516, P3_U3403, P3_U3893);
  not ginst26918 (P3_U5517, P3_U3404);
  nand ginst26919 (P3_U5518, P3_REG0_REG_5__SCAN_IN, P3_U3835);
  nand ginst26920 (P3_U5519, P3_U3914, P3_U4174);
  nand ginst26921 (P3_U5520, P3_IR_REG_6__SCAN_IN, P3_U3831);
  nand ginst26922 (P3_U5521, P3_IR_REG_31__SCAN_IN, P3_SUB_598_U25);
  nand ginst26923 (P3_U5522, P3_U3833, U33);
  nand ginst26924 (P3_U5523, P3_U3406, P3_U3893);
  not ginst26925 (P3_U5524, P3_U3407);
  nand ginst26926 (P3_U5525, P3_REG0_REG_6__SCAN_IN, P3_U3835);
  nand ginst26927 (P3_U5526, P3_U3914, P3_U4192);
  nand ginst26928 (P3_U5527, P3_IR_REG_7__SCAN_IN, P3_U3831);
  nand ginst26929 (P3_U5528, P3_IR_REG_31__SCAN_IN, P3_SUB_598_U26);
  nand ginst26930 (P3_U5529, P3_U3833, U32);
  nand ginst26931 (P3_U5530, P3_U3409, P3_U3893);
  not ginst26932 (P3_U5531, P3_U3410);
  nand ginst26933 (P3_U5532, P3_REG0_REG_7__SCAN_IN, P3_U3835);
  nand ginst26934 (P3_U5533, P3_U3914, P3_U4210);
  nand ginst26935 (P3_U5534, P3_IR_REG_8__SCAN_IN, P3_U3831);
  nand ginst26936 (P3_U5535, P3_IR_REG_31__SCAN_IN, P3_SUB_598_U27);
  nand ginst26937 (P3_U5536, P3_U3833, U31);
  nand ginst26938 (P3_U5537, P3_U3412, P3_U3893);
  not ginst26939 (P3_U5538, P3_U3413);
  nand ginst26940 (P3_U5539, P3_REG0_REG_8__SCAN_IN, P3_U3835);
  nand ginst26941 (P3_U5540, P3_U3914, P3_U4228);
  nand ginst26942 (P3_U5541, P3_IR_REG_9__SCAN_IN, P3_U3831);
  nand ginst26943 (P3_U5542, P3_IR_REG_31__SCAN_IN, P3_SUB_598_U72);
  nand ginst26944 (P3_U5543, P3_U3833, U30);
  nand ginst26945 (P3_U5544, P3_U3415, P3_U3893);
  not ginst26946 (P3_U5545, P3_U3416);
  nand ginst26947 (P3_U5546, P3_REG0_REG_9__SCAN_IN, P3_U3835);
  nand ginst26948 (P3_U5547, P3_U3914, P3_U4246);
  nand ginst26949 (P3_U5548, P3_IR_REG_10__SCAN_IN, P3_U3831);
  nand ginst26950 (P3_U5549, P3_IR_REG_31__SCAN_IN, P3_SUB_598_U7);
  nand ginst26951 (P3_U5550, P3_U3833, U60);
  nand ginst26952 (P3_U5551, P3_U3418, P3_U3893);
  not ginst26953 (P3_U5552, P3_U3419);
  nand ginst26954 (P3_U5553, P3_REG0_REG_10__SCAN_IN, P3_U3835);
  nand ginst26955 (P3_U5554, P3_U3914, P3_U4264);
  nand ginst26956 (P3_U5555, P3_IR_REG_11__SCAN_IN, P3_U3831);
  nand ginst26957 (P3_U5556, P3_IR_REG_31__SCAN_IN, P3_SUB_598_U8);
  nand ginst26958 (P3_U5557, P3_U3833, U59);
  nand ginst26959 (P3_U5558, P3_U3421, P3_U3893);
  not ginst26960 (P3_U5559, P3_U3422);
  nand ginst26961 (P3_U5560, P3_REG0_REG_11__SCAN_IN, P3_U3835);
  nand ginst26962 (P3_U5561, P3_U3914, P3_U4282);
  nand ginst26963 (P3_U5562, P3_IR_REG_12__SCAN_IN, P3_U3831);
  nand ginst26964 (P3_U5563, P3_IR_REG_31__SCAN_IN, P3_SUB_598_U9);
  nand ginst26965 (P3_U5564, P3_U3833, U58);
  nand ginst26966 (P3_U5565, P3_U3424, P3_U3893);
  not ginst26967 (P3_U5566, P3_U3425);
  nand ginst26968 (P3_U5567, P3_REG0_REG_12__SCAN_IN, P3_U3835);
  nand ginst26969 (P3_U5568, P3_U3914, P3_U4300);
  nand ginst26970 (P3_U5569, P3_IR_REG_13__SCAN_IN, P3_U3831);
  nand ginst26971 (P3_U5570, P3_IR_REG_31__SCAN_IN, P3_SUB_598_U89);
  nand ginst26972 (P3_U5571, P3_U3833, U57);
  nand ginst26973 (P3_U5572, P3_U3427, P3_U3893);
  not ginst26974 (P3_U5573, P3_U3428);
  nand ginst26975 (P3_U5574, P3_REG0_REG_13__SCAN_IN, P3_U3835);
  nand ginst26976 (P3_U5575, P3_U3914, P3_U4318);
  nand ginst26977 (P3_U5576, P3_IR_REG_14__SCAN_IN, P3_U3831);
  nand ginst26978 (P3_U5577, P3_IR_REG_31__SCAN_IN, P3_SUB_598_U10);
  nand ginst26979 (P3_U5578, P3_U3833, U56);
  nand ginst26980 (P3_U5579, P3_U3430, P3_U3893);
  not ginst26981 (P3_U5580, P3_U3431);
  nand ginst26982 (P3_U5581, P3_REG0_REG_14__SCAN_IN, P3_U3835);
  nand ginst26983 (P3_U5582, P3_U3914, P3_U4336);
  nand ginst26984 (P3_U5583, P3_IR_REG_15__SCAN_IN, P3_U3831);
  nand ginst26985 (P3_U5584, P3_IR_REG_31__SCAN_IN, P3_SUB_598_U11);
  nand ginst26986 (P3_U5585, P3_U3833, U55);
  nand ginst26987 (P3_U5586, P3_U3433, P3_U3893);
  not ginst26988 (P3_U5587, P3_U3434);
  nand ginst26989 (P3_U5588, P3_REG0_REG_15__SCAN_IN, P3_U3835);
  nand ginst26990 (P3_U5589, P3_U3914, P3_U4354);
  nand ginst26991 (P3_U5590, P3_IR_REG_16__SCAN_IN, P3_U3831);
  nand ginst26992 (P3_U5591, P3_IR_REG_31__SCAN_IN, P3_SUB_598_U12);
  nand ginst26993 (P3_U5592, P3_U3833, U54);
  nand ginst26994 (P3_U5593, P3_U3436, P3_U3893);
  not ginst26995 (P3_U5594, P3_U3437);
  nand ginst26996 (P3_U5595, P3_REG0_REG_16__SCAN_IN, P3_U3835);
  nand ginst26997 (P3_U5596, P3_U3914, P3_U4372);
  nand ginst26998 (P3_U5597, P3_IR_REG_17__SCAN_IN, P3_U3831);
  nand ginst26999 (P3_U5598, P3_IR_REG_31__SCAN_IN, P3_SUB_598_U87);
  nand ginst27000 (P3_U5599, P3_U3833, U53);
  nand ginst27001 (P3_U5600, P3_U3439, P3_U3893);
  not ginst27002 (P3_U5601, P3_U3440);
  nand ginst27003 (P3_U5602, P3_REG0_REG_17__SCAN_IN, P3_U3835);
  nand ginst27004 (P3_U5603, P3_U3914, P3_U4390);
  nand ginst27005 (P3_U5604, P3_IR_REG_18__SCAN_IN, P3_U3831);
  nand ginst27006 (P3_U5605, P3_IR_REG_31__SCAN_IN, P3_SUB_598_U13);
  nand ginst27007 (P3_U5606, P3_U3833, U52);
  nand ginst27008 (P3_U5607, P3_U3442, P3_U3893);
  not ginst27009 (P3_U5608, P3_U3443);
  nand ginst27010 (P3_U5609, P3_REG0_REG_18__SCAN_IN, P3_U3835);
  nand ginst27011 (P3_U5610, P3_U3914, P3_U4408);
  nand ginst27012 (P3_U5611, P3_U3833, U51);
  nand ginst27013 (P3_U5612, P3_U3379, P3_U3893);
  not ginst27014 (P3_U5613, P3_U3445);
  nand ginst27015 (P3_U5614, P3_REG0_REG_19__SCAN_IN, P3_U3835);
  nand ginst27016 (P3_U5615, P3_U3914, P3_U4426);
  nand ginst27017 (P3_U5616, P3_REG0_REG_20__SCAN_IN, P3_U3835);
  nand ginst27018 (P3_U5617, P3_U3914, P3_U4444);
  nand ginst27019 (P3_U5618, P3_REG0_REG_21__SCAN_IN, P3_U3835);
  nand ginst27020 (P3_U5619, P3_U3914, P3_U4462);
  nand ginst27021 (P3_U5620, P3_REG0_REG_22__SCAN_IN, P3_U3835);
  nand ginst27022 (P3_U5621, P3_U3914, P3_U4480);
  nand ginst27023 (P3_U5622, P3_REG0_REG_23__SCAN_IN, P3_U3835);
  nand ginst27024 (P3_U5623, P3_U3914, P3_U4498);
  nand ginst27025 (P3_U5624, P3_REG0_REG_24__SCAN_IN, P3_U3835);
  nand ginst27026 (P3_U5625, P3_U3914, P3_U4516);
  nand ginst27027 (P3_U5626, P3_REG0_REG_25__SCAN_IN, P3_U3835);
  nand ginst27028 (P3_U5627, P3_U3914, P3_U4534);
  nand ginst27029 (P3_U5628, P3_REG0_REG_26__SCAN_IN, P3_U3835);
  nand ginst27030 (P3_U5629, P3_U3914, P3_U4552);
  nand ginst27031 (P3_U5630, P3_REG0_REG_27__SCAN_IN, P3_U3835);
  nand ginst27032 (P3_U5631, P3_U3914, P3_U4570);
  nand ginst27033 (P3_U5632, P3_REG0_REG_28__SCAN_IN, P3_U3835);
  nand ginst27034 (P3_U5633, P3_U3914, P3_U4588);
  nand ginst27035 (P3_U5634, P3_REG0_REG_29__SCAN_IN, P3_U3835);
  nand ginst27036 (P3_U5635, P3_U3914, P3_U4608);
  nand ginst27037 (P3_U5636, P3_REG0_REG_30__SCAN_IN, P3_U3835);
  nand ginst27038 (P3_U5637, P3_U3914, P3_U4615);
  nand ginst27039 (P3_U5638, P3_REG0_REG_31__SCAN_IN, P3_U3835);
  nand ginst27040 (P3_U5639, P3_U3914, P3_U4617);
  nand ginst27041 (P3_U5640, P3_U3834, P3_U5453);
  nand ginst27042 (P3_U5641, P3_U4052, P3_U5450);
  nand ginst27043 (P3_U5642, P3_REG1_REG_0__SCAN_IN, P3_U3836);
  nand ginst27044 (P3_U5643, P3_U3913, P3_U4077);
  nand ginst27045 (P3_U5644, P3_REG1_REG_1__SCAN_IN, P3_U3836);
  nand ginst27046 (P3_U5645, P3_U3913, P3_U4102);
  nand ginst27047 (P3_U5646, P3_REG1_REG_2__SCAN_IN, P3_U3836);
  nand ginst27048 (P3_U5647, P3_U3913, P3_U4120);
  nand ginst27049 (P3_U5648, P3_REG1_REG_3__SCAN_IN, P3_U3836);
  nand ginst27050 (P3_U5649, P3_U3913, P3_U4138);
  nand ginst27051 (P3_U5650, P3_REG1_REG_4__SCAN_IN, P3_U3836);
  nand ginst27052 (P3_U5651, P3_U3913, P3_U4156);
  nand ginst27053 (P3_U5652, P3_REG1_REG_5__SCAN_IN, P3_U3836);
  nand ginst27054 (P3_U5653, P3_U3913, P3_U4174);
  nand ginst27055 (P3_U5654, P3_REG1_REG_6__SCAN_IN, P3_U3836);
  nand ginst27056 (P3_U5655, P3_U3913, P3_U4192);
  nand ginst27057 (P3_U5656, P3_REG1_REG_7__SCAN_IN, P3_U3836);
  nand ginst27058 (P3_U5657, P3_U3913, P3_U4210);
  nand ginst27059 (P3_U5658, P3_REG1_REG_8__SCAN_IN, P3_U3836);
  nand ginst27060 (P3_U5659, P3_U3913, P3_U4228);
  nand ginst27061 (P3_U5660, P3_REG1_REG_9__SCAN_IN, P3_U3836);
  nand ginst27062 (P3_U5661, P3_U3913, P3_U4246);
  nand ginst27063 (P3_U5662, P3_REG1_REG_10__SCAN_IN, P3_U3836);
  nand ginst27064 (P3_U5663, P3_U3913, P3_U4264);
  nand ginst27065 (P3_U5664, P3_REG1_REG_11__SCAN_IN, P3_U3836);
  nand ginst27066 (P3_U5665, P3_U3913, P3_U4282);
  nand ginst27067 (P3_U5666, P3_REG1_REG_12__SCAN_IN, P3_U3836);
  nand ginst27068 (P3_U5667, P3_U3913, P3_U4300);
  nand ginst27069 (P3_U5668, P3_REG1_REG_13__SCAN_IN, P3_U3836);
  nand ginst27070 (P3_U5669, P3_U3913, P3_U4318);
  nand ginst27071 (P3_U5670, P3_REG1_REG_14__SCAN_IN, P3_U3836);
  nand ginst27072 (P3_U5671, P3_U3913, P3_U4336);
  nand ginst27073 (P3_U5672, P3_REG1_REG_15__SCAN_IN, P3_U3836);
  nand ginst27074 (P3_U5673, P3_U3913, P3_U4354);
  nand ginst27075 (P3_U5674, P3_REG1_REG_16__SCAN_IN, P3_U3836);
  nand ginst27076 (P3_U5675, P3_U3913, P3_U4372);
  nand ginst27077 (P3_U5676, P3_REG1_REG_17__SCAN_IN, P3_U3836);
  nand ginst27078 (P3_U5677, P3_U3913, P3_U4390);
  nand ginst27079 (P3_U5678, P3_REG1_REG_18__SCAN_IN, P3_U3836);
  nand ginst27080 (P3_U5679, P3_U3913, P3_U4408);
  nand ginst27081 (P3_U5680, P3_REG1_REG_19__SCAN_IN, P3_U3836);
  nand ginst27082 (P3_U5681, P3_U3913, P3_U4426);
  nand ginst27083 (P3_U5682, P3_REG1_REG_20__SCAN_IN, P3_U3836);
  nand ginst27084 (P3_U5683, P3_U3913, P3_U4444);
  nand ginst27085 (P3_U5684, P3_REG1_REG_21__SCAN_IN, P3_U3836);
  nand ginst27086 (P3_U5685, P3_U3913, P3_U4462);
  nand ginst27087 (P3_U5686, P3_REG1_REG_22__SCAN_IN, P3_U3836);
  nand ginst27088 (P3_U5687, P3_U3913, P3_U4480);
  nand ginst27089 (P3_U5688, P3_REG1_REG_23__SCAN_IN, P3_U3836);
  nand ginst27090 (P3_U5689, P3_U3913, P3_U4498);
  nand ginst27091 (P3_U5690, P3_REG1_REG_24__SCAN_IN, P3_U3836);
  nand ginst27092 (P3_U5691, P3_U3913, P3_U4516);
  nand ginst27093 (P3_U5692, P3_REG1_REG_25__SCAN_IN, P3_U3836);
  nand ginst27094 (P3_U5693, P3_U3913, P3_U4534);
  nand ginst27095 (P3_U5694, P3_REG1_REG_26__SCAN_IN, P3_U3836);
  nand ginst27096 (P3_U5695, P3_U3913, P3_U4552);
  nand ginst27097 (P3_U5696, P3_REG1_REG_27__SCAN_IN, P3_U3836);
  nand ginst27098 (P3_U5697, P3_U3913, P3_U4570);
  nand ginst27099 (P3_U5698, P3_REG1_REG_28__SCAN_IN, P3_U3836);
  nand ginst27100 (P3_U5699, P3_U3913, P3_U4588);
  nand ginst27101 (P3_U5700, P3_REG1_REG_29__SCAN_IN, P3_U3836);
  nand ginst27102 (P3_U5701, P3_U3913, P3_U4608);
  nand ginst27103 (P3_U5702, P3_REG1_REG_30__SCAN_IN, P3_U3836);
  nand ginst27104 (P3_U5703, P3_U3913, P3_U4615);
  nand ginst27105 (P3_U5704, P3_REG1_REG_31__SCAN_IN, P3_U3836);
  nand ginst27106 (P3_U5705, P3_U3913, P3_U4617);
  nand ginst27107 (P3_U5706, P3_REG2_REG_0__SCAN_IN, P3_U3358);
  nand ginst27108 (P3_U5707, P3_U3314, P3_U3912);
  nand ginst27109 (P3_U5708, P3_REG2_REG_1__SCAN_IN, P3_U3358);
  nand ginst27110 (P3_U5709, P3_U3315, P3_U3912);
  nand ginst27111 (P3_U5710, P3_REG2_REG_2__SCAN_IN, P3_U3358);
  nand ginst27112 (P3_U5711, P3_U3316, P3_U3912);
  nand ginst27113 (P3_U5712, P3_REG2_REG_3__SCAN_IN, P3_U3358);
  nand ginst27114 (P3_U5713, P3_U3317, P3_U3912);
  nand ginst27115 (P3_U5714, P3_REG2_REG_4__SCAN_IN, P3_U3358);
  nand ginst27116 (P3_U5715, P3_U3318, P3_U3912);
  nand ginst27117 (P3_U5716, P3_REG2_REG_5__SCAN_IN, P3_U3358);
  nand ginst27118 (P3_U5717, P3_U3319, P3_U3912);
  nand ginst27119 (P3_U5718, P3_REG2_REG_6__SCAN_IN, P3_U3358);
  nand ginst27120 (P3_U5719, P3_U3320, P3_U3912);
  nand ginst27121 (P3_U5720, P3_REG2_REG_7__SCAN_IN, P3_U3358);
  nand ginst27122 (P3_U5721, P3_U3321, P3_U3912);
  nand ginst27123 (P3_U5722, P3_REG2_REG_8__SCAN_IN, P3_U3358);
  nand ginst27124 (P3_U5723, P3_U3322, P3_U3912);
  nand ginst27125 (P3_U5724, P3_REG2_REG_9__SCAN_IN, P3_U3358);
  nand ginst27126 (P3_U5725, P3_U3323, P3_U3912);
  nand ginst27127 (P3_U5726, P3_REG2_REG_10__SCAN_IN, P3_U3358);
  nand ginst27128 (P3_U5727, P3_U3324, P3_U3912);
  nand ginst27129 (P3_U5728, P3_REG2_REG_11__SCAN_IN, P3_U3358);
  nand ginst27130 (P3_U5729, P3_U3325, P3_U3912);
  nand ginst27131 (P3_U5730, P3_REG2_REG_12__SCAN_IN, P3_U3358);
  nand ginst27132 (P3_U5731, P3_U3326, P3_U3912);
  nand ginst27133 (P3_U5732, P3_REG2_REG_13__SCAN_IN, P3_U3358);
  nand ginst27134 (P3_U5733, P3_U3327, P3_U3912);
  nand ginst27135 (P3_U5734, P3_REG2_REG_14__SCAN_IN, P3_U3358);
  nand ginst27136 (P3_U5735, P3_U3328, P3_U3912);
  nand ginst27137 (P3_U5736, P3_REG2_REG_15__SCAN_IN, P3_U3358);
  nand ginst27138 (P3_U5737, P3_U3329, P3_U3912);
  nand ginst27139 (P3_U5738, P3_REG2_REG_16__SCAN_IN, P3_U3358);
  nand ginst27140 (P3_U5739, P3_U3330, P3_U3912);
  nand ginst27141 (P3_U5740, P3_REG2_REG_17__SCAN_IN, P3_U3358);
  nand ginst27142 (P3_U5741, P3_U3331, P3_U3912);
  nand ginst27143 (P3_U5742, P3_REG2_REG_18__SCAN_IN, P3_U3358);
  nand ginst27144 (P3_U5743, P3_U3332, P3_U3912);
  nand ginst27145 (P3_U5744, P3_REG2_REG_19__SCAN_IN, P3_U3358);
  nand ginst27146 (P3_U5745, P3_U3333, P3_U3912);
  nand ginst27147 (P3_U5746, P3_REG2_REG_20__SCAN_IN, P3_U3358);
  nand ginst27148 (P3_U5747, P3_U3335, P3_U3912);
  nand ginst27149 (P3_U5748, P3_REG2_REG_21__SCAN_IN, P3_U3358);
  nand ginst27150 (P3_U5749, P3_U3337, P3_U3912);
  nand ginst27151 (P3_U5750, P3_REG2_REG_22__SCAN_IN, P3_U3358);
  nand ginst27152 (P3_U5751, P3_U3339, P3_U3912);
  nand ginst27153 (P3_U5752, P3_REG2_REG_23__SCAN_IN, P3_U3358);
  nand ginst27154 (P3_U5753, P3_U3341, P3_U3912);
  nand ginst27155 (P3_U5754, P3_REG2_REG_24__SCAN_IN, P3_U3358);
  nand ginst27156 (P3_U5755, P3_U3343, P3_U3912);
  nand ginst27157 (P3_U5756, P3_REG2_REG_25__SCAN_IN, P3_U3358);
  nand ginst27158 (P3_U5757, P3_U3345, P3_U3912);
  nand ginst27159 (P3_U5758, P3_REG2_REG_26__SCAN_IN, P3_U3358);
  nand ginst27160 (P3_U5759, P3_U3347, P3_U3912);
  nand ginst27161 (P3_U5760, P3_REG2_REG_27__SCAN_IN, P3_U3358);
  nand ginst27162 (P3_U5761, P3_U3349, P3_U3912);
  nand ginst27163 (P3_U5762, P3_REG2_REG_28__SCAN_IN, P3_U3358);
  nand ginst27164 (P3_U5763, P3_U3351, P3_U3912);
  nand ginst27165 (P3_U5764, P3_REG2_REG_29__SCAN_IN, P3_U3358);
  nand ginst27166 (P3_U5765, P3_U3354, P3_U3912);
  nand ginst27167 (P3_U5766, P3_U3024, P3_U5465);
  nand ginst27168 (P3_U5767, P3_U3383, P3_U3897);
  nand ginst27169 (P3_U5768, P3_U5766, P3_U5767);
  nand ginst27170 (P3_U5769, P3_DATAO_REG_0__SCAN_IN, P3_U3363);
  nand ginst27171 (P3_U5770, P3_U3076, P3_U3897);
  nand ginst27172 (P3_U5771, P3_DATAO_REG_1__SCAN_IN, P3_U3363);
  nand ginst27173 (P3_U5772, P3_U3077, P3_U3897);
  nand ginst27174 (P3_U5773, P3_DATAO_REG_2__SCAN_IN, P3_U3363);
  nand ginst27175 (P3_U5774, P3_U3067, P3_U3897);
  nand ginst27176 (P3_U5775, P3_DATAO_REG_3__SCAN_IN, P3_U3363);
  nand ginst27177 (P3_U5776, P3_U3063, P3_U3897);
  nand ginst27178 (P3_U5777, P3_DATAO_REG_4__SCAN_IN, P3_U3363);
  nand ginst27179 (P3_U5778, P3_U3059, P3_U3897);
  nand ginst27180 (P3_U5779, P3_DATAO_REG_5__SCAN_IN, P3_U3363);
  nand ginst27181 (P3_U5780, P3_U3066, P3_U3897);
  nand ginst27182 (P3_U5781, P3_DATAO_REG_6__SCAN_IN, P3_U3363);
  nand ginst27183 (P3_U5782, P3_U3070, P3_U3897);
  nand ginst27184 (P3_U5783, P3_DATAO_REG_7__SCAN_IN, P3_U3363);
  nand ginst27185 (P3_U5784, P3_U3069, P3_U3897);
  nand ginst27186 (P3_U5785, P3_DATAO_REG_8__SCAN_IN, P3_U3363);
  nand ginst27187 (P3_U5786, P3_U3083, P3_U3897);
  nand ginst27188 (P3_U5787, P3_DATAO_REG_9__SCAN_IN, P3_U3363);
  nand ginst27189 (P3_U5788, P3_U3082, P3_U3897);
  nand ginst27190 (P3_U5789, P3_DATAO_REG_10__SCAN_IN, P3_U3363);
  nand ginst27191 (P3_U5790, P3_U3061, P3_U3897);
  nand ginst27192 (P3_U5791, P3_DATAO_REG_11__SCAN_IN, P3_U3363);
  nand ginst27193 (P3_U5792, P3_U3062, P3_U3897);
  nand ginst27194 (P3_U5793, P3_DATAO_REG_12__SCAN_IN, P3_U3363);
  nand ginst27195 (P3_U5794, P3_U3071, P3_U3897);
  nand ginst27196 (P3_U5795, P3_DATAO_REG_13__SCAN_IN, P3_U3363);
  nand ginst27197 (P3_U5796, P3_U3079, P3_U3897);
  nand ginst27198 (P3_U5797, P3_DATAO_REG_14__SCAN_IN, P3_U3363);
  nand ginst27199 (P3_U5798, P3_U3078, P3_U3897);
  nand ginst27200 (P3_U5799, P3_DATAO_REG_15__SCAN_IN, P3_U3363);
  nand ginst27201 (P3_U5800, P3_U3073, P3_U3897);
  nand ginst27202 (P3_U5801, P3_DATAO_REG_16__SCAN_IN, P3_U3363);
  nand ginst27203 (P3_U5802, P3_U3072, P3_U3897);
  nand ginst27204 (P3_U5803, P3_DATAO_REG_17__SCAN_IN, P3_U3363);
  nand ginst27205 (P3_U5804, P3_U3068, P3_U3897);
  nand ginst27206 (P3_U5805, P3_DATAO_REG_18__SCAN_IN, P3_U3363);
  nand ginst27207 (P3_U5806, P3_U3081, P3_U3897);
  nand ginst27208 (P3_U5807, P3_DATAO_REG_19__SCAN_IN, P3_U3363);
  nand ginst27209 (P3_U5808, P3_U3080, P3_U3897);
  nand ginst27210 (P3_U5809, P3_DATAO_REG_20__SCAN_IN, P3_U3363);
  nand ginst27211 (P3_U5810, P3_U3075, P3_U3897);
  nand ginst27212 (P3_U5811, P3_DATAO_REG_21__SCAN_IN, P3_U3363);
  nand ginst27213 (P3_U5812, P3_U3074, P3_U3897);
  nand ginst27214 (P3_U5813, P3_DATAO_REG_22__SCAN_IN, P3_U3363);
  nand ginst27215 (P3_U5814, P3_U3060, P3_U3897);
  nand ginst27216 (P3_U5815, P3_DATAO_REG_23__SCAN_IN, P3_U3363);
  nand ginst27217 (P3_U5816, P3_U3065, P3_U3897);
  nand ginst27218 (P3_U5817, P3_DATAO_REG_24__SCAN_IN, P3_U3363);
  nand ginst27219 (P3_U5818, P3_U3064, P3_U3897);
  nand ginst27220 (P3_U5819, P3_DATAO_REG_25__SCAN_IN, P3_U3363);
  nand ginst27221 (P3_U5820, P3_U3057, P3_U3897);
  nand ginst27222 (P3_U5821, P3_DATAO_REG_26__SCAN_IN, P3_U3363);
  nand ginst27223 (P3_U5822, P3_U3056, P3_U3897);
  nand ginst27224 (P3_U5823, P3_DATAO_REG_27__SCAN_IN, P3_U3363);
  nand ginst27225 (P3_U5824, P3_U3052, P3_U3897);
  nand ginst27226 (P3_U5825, P3_DATAO_REG_28__SCAN_IN, P3_U3363);
  nand ginst27227 (P3_U5826, P3_U3053, P3_U3897);
  nand ginst27228 (P3_U5827, P3_DATAO_REG_29__SCAN_IN, P3_U3363);
  nand ginst27229 (P3_U5828, P3_U3054, P3_U3897);
  nand ginst27230 (P3_U5829, P3_DATAO_REG_30__SCAN_IN, P3_U3363);
  nand ginst27231 (P3_U5830, P3_U3058, P3_U3897);
  nand ginst27232 (P3_U5831, P3_DATAO_REG_31__SCAN_IN, P3_U3363);
  nand ginst27233 (P3_U5832, P3_U3055, P3_U3897);
  nand ginst27234 (P3_U5833, P3_U3313, P3_U3379);
  nand ginst27235 (P3_U5834, P3_U3911, P3_U5450);
  not ginst27236 (P3_U5835, P3_U3760);
  nand ginst27237 (P3_U5836, P3_R1269_U11, P3_U5835);
  nand ginst27238 (P3_U5837, P3_U3760, P3_U3867);
  nand ginst27239 (P3_U5838, P3_U3052, P3_U3900);
  nand ginst27240 (P3_U5839, P3_U3348, P3_U4539);
  nand ginst27241 (P3_U5840, P3_U5838, P3_U5839);
  nand ginst27242 (P3_U5841, P3_U3053, P3_U3899);
  nand ginst27243 (P3_U5842, P3_U3350, P3_U4557);
  nand ginst27244 (P3_U5843, P3_U5841, P3_U5842);
  nand ginst27245 (P3_U5844, P3_U3055, P3_U3872);
  nand ginst27246 (P3_U5845, P3_U3356, P3_U4613);
  nand ginst27247 (P3_U5846, P3_U5844, P3_U5845);
  nand ginst27248 (P3_U5847, P3_U3054, P3_U3908);
  nand ginst27249 (P3_U5848, P3_U3353, P3_U4575);
  nand ginst27250 (P3_U5849, P3_U5847, P3_U5848);
  nand ginst27251 (P3_U5850, P3_U3074, P3_U3906);
  nand ginst27252 (P3_U5851, P3_U3336, P3_U4431);
  nand ginst27253 (P3_U5852, P3_U5850, P3_U5851);
  nand ginst27254 (P3_U5853, P3_U3075, P3_U3907);
  nand ginst27255 (P3_U5854, P3_U3334, P3_U4413);
  nand ginst27256 (P3_U5855, P3_U5853, P3_U5854);
  nand ginst27257 (P3_U5856, P3_U4107, P3_U5503);
  nand ginst27258 (P3_U5857, P3_U3063, P3_U3398);
  nand ginst27259 (P3_U5858, P3_U5856, P3_U5857);
  nand ginst27260 (P3_U5859, P3_U4251, P3_U5559);
  nand ginst27261 (P3_U5860, P3_U3062, P3_U3422);
  nand ginst27262 (P3_U5861, P3_U5859, P3_U5860);
  nand ginst27263 (P3_U5862, P3_U4233, P3_U5552);
  nand ginst27264 (P3_U5863, P3_U3061, P3_U3419);
  nand ginst27265 (P3_U5864, P3_U5862, P3_U5863);
  nand ginst27266 (P3_U5865, P3_U4125, P3_U5510);
  nand ginst27267 (P3_U5866, P3_U3059, P3_U3401);
  nand ginst27268 (P3_U5867, P3_U5865, P3_U5866);
  nand ginst27269 (P3_U5868, P3_U3060, P3_U3905);
  nand ginst27270 (P3_U5869, P3_U3338, P3_U4449);
  nand ginst27271 (P3_U5870, P3_U5868, P3_U5869);
  nand ginst27272 (P3_U5871, P3_U4359, P3_U5601);
  nand ginst27273 (P3_U5872, P3_U3068, P3_U3440);
  nand ginst27274 (P3_U5873, P3_U5871, P3_U5872);
  nand ginst27275 (P3_U5874, P3_U4341, P3_U5594);
  nand ginst27276 (P3_U5875, P3_U3072, P3_U3437);
  nand ginst27277 (P3_U5876, P3_U5874, P3_U5875);
  nand ginst27278 (P3_U5877, P3_U4323, P3_U5587);
  nand ginst27279 (P3_U5878, P3_U3073, P3_U3434);
  nand ginst27280 (P3_U5879, P3_U5877, P3_U5878);
  nand ginst27281 (P3_U5880, P3_U4269, P3_U5566);
  nand ginst27282 (P3_U5881, P3_U3071, P3_U3425);
  nand ginst27283 (P3_U5882, P3_U5880, P3_U5881);
  nand ginst27284 (P3_U5883, P3_U4161, P3_U5524);
  nand ginst27285 (P3_U5884, P3_U3070, P3_U3407);
  nand ginst27286 (P3_U5885, P3_U5883, P3_U5884);
  nand ginst27287 (P3_U5886, P3_U4179, P3_U5531);
  nand ginst27288 (P3_U5887, P3_U3069, P3_U3410);
  nand ginst27289 (P3_U5888, P3_U5886, P3_U5887);
  nand ginst27290 (P3_U5889, P3_U4082, P3_U5496);
  nand ginst27291 (P3_U5890, P3_U3067, P3_U3395);
  nand ginst27292 (P3_U5891, P3_U5889, P3_U5890);
  nand ginst27293 (P3_U5892, P3_U4143, P3_U5517);
  nand ginst27294 (P3_U5893, P3_U3066, P3_U3404);
  nand ginst27295 (P3_U5894, P3_U5892, P3_U5893);
  nand ginst27296 (P3_U5895, P3_U4377, P3_U5608);
  nand ginst27297 (P3_U5896, P3_U3081, P3_U3443);
  nand ginst27298 (P3_U5897, P3_U5895, P3_U5896);
  nand ginst27299 (P3_U5898, P3_U4287, P3_U5573);
  nand ginst27300 (P3_U5899, P3_U3079, P3_U3428);
  nand ginst27301 (P3_U5900, P3_U5898, P3_U5899);
  nand ginst27302 (P3_U5901, P3_U4305, P3_U5580);
  nand ginst27303 (P3_U5902, P3_U3078, P3_U3431);
  nand ginst27304 (P3_U5903, P3_U5901, P3_U5902);
  nand ginst27305 (P3_U5904, P3_U4063, P3_U5489);
  nand ginst27306 (P3_U5905, P3_U3077, P3_U3392);
  nand ginst27307 (P3_U5906, P3_U5904, P3_U5905);
  nand ginst27308 (P3_U5907, P3_U4087, P3_U5473);
  nand ginst27309 (P3_U5908, P3_U3076, P3_U3387);
  nand ginst27310 (P3_U5909, P3_U5907, P3_U5908);
  nand ginst27311 (P3_U5910, P3_U4197, P3_U5538);
  nand ginst27312 (P3_U5911, P3_U3083, P3_U3413);
  nand ginst27313 (P3_U5912, P3_U5910, P3_U5911);
  nand ginst27314 (P3_U5913, P3_U4215, P3_U5545);
  nand ginst27315 (P3_U5914, P3_U3082, P3_U3416);
  nand ginst27316 (P3_U5915, P3_U5913, P3_U5914);
  nand ginst27317 (P3_U5916, P3_U4395, P3_U5613);
  nand ginst27318 (P3_U5917, P3_U3080, P3_U3445);
  nand ginst27319 (P3_U5918, P3_U5916, P3_U5917);
  nand ginst27320 (P3_U5919, P3_U3056, P3_U3901);
  nand ginst27321 (P3_U5920, P3_U3346, P3_U4521);
  nand ginst27322 (P3_U5921, P3_U5919, P3_U5920);
  nand ginst27323 (P3_U5922, P3_U3057, P3_U3902);
  nand ginst27324 (P3_U5923, P3_U3344, P3_U4503);
  nand ginst27325 (P3_U5924, P3_U5922, P3_U5923);
  nand ginst27326 (P3_U5925, P3_U3065, P3_U3904);
  nand ginst27327 (P3_U5926, P3_U3340, P3_U4467);
  nand ginst27328 (P3_U5927, P3_U5925, P3_U5926);
  nand ginst27329 (P3_U5928, P3_U3064, P3_U3903);
  nand ginst27330 (P3_U5929, P3_U3342, P3_U4485);
  nand ginst27331 (P3_U5930, P3_U5928, P3_U5929);
  nand ginst27332 (P3_U5931, P3_U3058, P3_U3873);
  nand ginst27333 (P3_U5932, P3_U3355, P3_U4593);
  nand ginst27334 (P3_U5933, P3_U5931, P3_U5932);
  nand ginst27335 (P3_U5934, P3_U4978, P3_U5450);
  nand ginst27336 (P3_U5935, P3_U3379, P3_U3868);
  nand ginst27337 (P3_U5936, P3_U5934, P3_U5935);
  nand ginst27338 (P3_U5937, P3_U5447, P3_U5836, P3_U5837);
  nand ginst27339 (P3_U5938, P3_U3378, P3_U5456, P3_U5936);
  nand ginst27340 (P3_U5939, P3_U3869, P3_U3881);
  nand ginst27341 (P3_U5940, P3_R693_U14, P3_U3891);
  nand ginst27342 (P3_U5941, P3_U3368, P3_U5440);
  nand ginst27343 (P3_U5942, P3_U3375, P3_U3380);
  nand ginst27344 (P3_U5943, P3_U5447, P3_U5450);
  nand ginst27345 (P3_U5944, P3_U3378, P3_U3388, P3_U5456);
  nand ginst27346 (P3_U5945, P3_R1297_U6, P3_U3082);
  nand ginst27347 (P3_U5946, P3_U3082, P3_U3871);
  nand ginst27348 (P3_U5947, P3_R1297_U6, P3_U3083);
  nand ginst27349 (P3_U5948, P3_U3083, P3_U3871);
  nand ginst27350 (P3_U5949, P3_R1297_U6, P3_U3069);
  nand ginst27351 (P3_U5950, P3_U3069, P3_U3871);
  nand ginst27352 (P3_U5951, P3_R1297_U6, P3_U3070);
  nand ginst27353 (P3_U5952, P3_U3070, P3_U3871);
  nand ginst27354 (P3_U5953, P3_R1297_U6, P3_U3066);
  nand ginst27355 (P3_U5954, P3_U3066, P3_U3871);
  nand ginst27356 (P3_U5955, P3_R1297_U6, P3_U3059);
  nand ginst27357 (P3_U5956, P3_U3059, P3_U3871);
  nand ginst27358 (P3_U5957, P3_R1297_U6, P3_R1300_U8);
  nand ginst27359 (P3_U5958, P3_U3055, P3_U3871);
  nand ginst27360 (P3_U5959, P3_R1297_U6, P3_R1300_U6);
  nand ginst27361 (P3_U5960, P3_U3058, P3_U3871);
  nand ginst27362 (P3_U5961, P3_R1297_U6, P3_U3063);
  nand ginst27363 (P3_U5962, P3_U3063, P3_U3871);
  nand ginst27364 (P3_U5963, P3_R1297_U6, P3_U3054);
  nand ginst27365 (P3_U5964, P3_U3054, P3_U3871);
  nand ginst27366 (P3_U5965, P3_R1297_U6, P3_U3053);
  nand ginst27367 (P3_U5966, P3_U3053, P3_U3871);
  nand ginst27368 (P3_U5967, P3_R1297_U6, P3_U3052);
  nand ginst27369 (P3_U5968, P3_U3052, P3_U3871);
  nand ginst27370 (P3_U5969, P3_R1297_U6, P3_U3056);
  nand ginst27371 (P3_U5970, P3_U3056, P3_U3871);
  nand ginst27372 (P3_U5971, P3_R1297_U6, P3_U3057);
  nand ginst27373 (P3_U5972, P3_U3057, P3_U3871);
  nand ginst27374 (P3_U5973, P3_R1297_U6, P3_U3064);
  nand ginst27375 (P3_U5974, P3_U3064, P3_U3871);
  nand ginst27376 (P3_U5975, P3_R1297_U6, P3_U3065);
  nand ginst27377 (P3_U5976, P3_U3065, P3_U3871);
  nand ginst27378 (P3_U5977, P3_R1297_U6, P3_U3060);
  nand ginst27379 (P3_U5978, P3_U3060, P3_U3871);
  nand ginst27380 (P3_U5979, P3_R1297_U6, P3_U3074);
  nand ginst27381 (P3_U5980, P3_U3074, P3_U3871);
  nand ginst27382 (P3_U5981, P3_R1297_U6, P3_U3075);
  nand ginst27383 (P3_U5982, P3_U3075, P3_U3871);
  nand ginst27384 (P3_U5983, P3_R1297_U6, P3_U3067);
  nand ginst27385 (P3_U5984, P3_U3067, P3_U3871);
  nand ginst27386 (P3_U5985, P3_R1297_U6, P3_U3080);
  nand ginst27387 (P3_U5986, P3_U3080, P3_U3871);
  nand ginst27388 (P3_U5987, P3_R1297_U6, P3_U3081);
  nand ginst27389 (P3_U5988, P3_U3081, P3_U3871);
  nand ginst27390 (P3_U5989, P3_R1297_U6, P3_U3068);
  nand ginst27391 (P3_U5990, P3_U3068, P3_U3871);
  nand ginst27392 (P3_U5991, P3_R1297_U6, P3_U3072);
  nand ginst27393 (P3_U5992, P3_U3072, P3_U3871);
  nand ginst27394 (P3_U5993, P3_R1297_U6, P3_U3073);
  nand ginst27395 (P3_U5994, P3_U3073, P3_U3871);
  nand ginst27396 (P3_U5995, P3_R1297_U6, P3_U3078);
  nand ginst27397 (P3_U5996, P3_U3078, P3_U3871);
  nand ginst27398 (P3_U5997, P3_R1297_U6, P3_U3079);
  nand ginst27399 (P3_U5998, P3_U3079, P3_U3871);
  nand ginst27400 (P3_U5999, P3_R1297_U6, P3_U3071);
  nand ginst27401 (P3_U6000, P3_U3071, P3_U3871);
  nand ginst27402 (P3_U6001, P3_R1297_U6, P3_U3062);
  nand ginst27403 (P3_U6002, P3_U3062, P3_U3871);
  nand ginst27404 (P3_U6003, P3_R1297_U6, P3_U3061);
  nand ginst27405 (P3_U6004, P3_U3061, P3_U3871);
  nand ginst27406 (P3_U6005, P3_R1297_U6, P3_U3077);
  nand ginst27407 (P3_U6006, P3_U3077, P3_U3871);
  nand ginst27408 (P3_U6007, P3_R1297_U6, P3_U3076);
  nand ginst27409 (P3_U6008, P3_U3076, P3_U3871);
  nand ginst27410 (P3_U6009, P3_REG1_REG_9__SCAN_IN, P3_U5468);
  nand ginst27411 (P3_U6010, P3_REG2_REG_9__SCAN_IN, P3_U3384);
  nand ginst27412 (P3_U6011, P3_REG1_REG_8__SCAN_IN, P3_U5468);
  nand ginst27413 (P3_U6012, P3_REG2_REG_8__SCAN_IN, P3_U3384);
  nand ginst27414 (P3_U6013, P3_REG1_REG_7__SCAN_IN, P3_U5468);
  nand ginst27415 (P3_U6014, P3_REG2_REG_7__SCAN_IN, P3_U3384);
  nand ginst27416 (P3_U6015, P3_REG1_REG_6__SCAN_IN, P3_U5468);
  nand ginst27417 (P3_U6016, P3_REG2_REG_6__SCAN_IN, P3_U3384);
  nand ginst27418 (P3_U6017, P3_REG1_REG_5__SCAN_IN, P3_U5468);
  nand ginst27419 (P3_U6018, P3_REG2_REG_5__SCAN_IN, P3_U3384);
  nand ginst27420 (P3_U6019, P3_REG1_REG_4__SCAN_IN, P3_U5468);
  nand ginst27421 (P3_U6020, P3_REG2_REG_4__SCAN_IN, P3_U3384);
  nand ginst27422 (P3_U6021, P3_REG1_REG_3__SCAN_IN, P3_U5468);
  nand ginst27423 (P3_U6022, P3_REG2_REG_3__SCAN_IN, P3_U3384);
  nand ginst27424 (P3_U6023, P3_REG1_REG_2__SCAN_IN, P3_U5468);
  nand ginst27425 (P3_U6024, P3_REG2_REG_2__SCAN_IN, P3_U3384);
  nand ginst27426 (P3_U6025, P3_REG1_REG_19__SCAN_IN, P3_U5468);
  nand ginst27427 (P3_U6026, P3_REG2_REG_19__SCAN_IN, P3_U3384);
  nand ginst27428 (P3_U6027, P3_REG1_REG_18__SCAN_IN, P3_U5468);
  nand ginst27429 (P3_U6028, P3_REG2_REG_18__SCAN_IN, P3_U3384);
  nand ginst27430 (P3_U6029, P3_REG1_REG_17__SCAN_IN, P3_U5468);
  nand ginst27431 (P3_U6030, P3_REG2_REG_17__SCAN_IN, P3_U3384);
  nand ginst27432 (P3_U6031, P3_REG1_REG_16__SCAN_IN, P3_U5468);
  nand ginst27433 (P3_U6032, P3_REG2_REG_16__SCAN_IN, P3_U3384);
  nand ginst27434 (P3_U6033, P3_REG1_REG_15__SCAN_IN, P3_U5468);
  nand ginst27435 (P3_U6034, P3_REG2_REG_15__SCAN_IN, P3_U3384);
  nand ginst27436 (P3_U6035, P3_REG1_REG_14__SCAN_IN, P3_U5468);
  nand ginst27437 (P3_U6036, P3_REG2_REG_14__SCAN_IN, P3_U3384);
  nand ginst27438 (P3_U6037, P3_REG1_REG_13__SCAN_IN, P3_U5468);
  nand ginst27439 (P3_U6038, P3_REG2_REG_13__SCAN_IN, P3_U3384);
  nand ginst27440 (P3_U6039, P3_REG1_REG_12__SCAN_IN, P3_U5468);
  nand ginst27441 (P3_U6040, P3_REG2_REG_12__SCAN_IN, P3_U3384);
  nand ginst27442 (P3_U6041, P3_REG1_REG_11__SCAN_IN, P3_U5468);
  nand ginst27443 (P3_U6042, P3_REG2_REG_11__SCAN_IN, P3_U3384);
  nand ginst27444 (P3_U6043, P3_REG1_REG_10__SCAN_IN, P3_U5468);
  nand ginst27445 (P3_U6044, P3_REG2_REG_10__SCAN_IN, P3_U3384);
  nand ginst27446 (P3_U6045, P3_REG1_REG_1__SCAN_IN, P3_U5468);
  nand ginst27447 (P3_U6046, P3_REG2_REG_1__SCAN_IN, P3_U3384);
  nand ginst27448 (P3_U6047, P3_REG1_REG_0__SCAN_IN, P3_U5468);
  nand ginst27449 (P3_U6048, P3_REG2_REG_0__SCAN_IN, P3_U3384);
  and ginst27450 (R152_U10, R152_U196, R152_U199);
  nand ginst27451 (R152_U100, R152_U455, R152_U456);
  nand ginst27452 (R152_U101, R152_U462, R152_U463);
  nand ginst27453 (R152_U102, R152_U469, R152_U470);
  nand ginst27454 (R152_U103, R152_U476, R152_U477);
  nand ginst27455 (R152_U104, R152_U488, R152_U489);
  nand ginst27456 (R152_U105, R152_U495, R152_U496);
  nand ginst27457 (R152_U106, R152_U502, R152_U503);
  nand ginst27458 (R152_U107, R152_U509, R152_U510);
  nand ginst27459 (R152_U108, R152_U516, R152_U517);
  nand ginst27460 (R152_U109, R152_U523, R152_U524);
  and ginst27461 (R152_U11, R152_U390, R152_U391);
  nand ginst27462 (R152_U110, R152_U530, R152_U531);
  nand ginst27463 (R152_U111, R152_U537, R152_U538);
  nand ginst27464 (R152_U112, R152_U544, R152_U545);
  nand ginst27465 (R152_U113, R152_U551, R152_U552);
  and ginst27466 (R152_U114, R152_U200, R152_U292);
  and ginst27467 (R152_U115, R152_U209, R152_U4);
  and ginst27468 (R152_U116, R152_U210, R152_U297);
  and ginst27469 (R152_U117, R152_U215, R152_U298);
  and ginst27470 (R152_U118, R152_U200, R152_U292);
  and ginst27471 (R152_U119, U156, U157);
  and ginst27472 (R152_U12, R152_U128, R152_U193);
  and ginst27473 (R152_U120, SI_0_, U157);
  and ginst27474 (R152_U121, SI_1_, U156);
  and ginst27475 (R152_U122, R152_U218, R152_U6);
  and ginst27476 (R152_U123, R152_U219, R152_U302);
  and ginst27477 (R152_U124, R152_U228, R152_U9);
  and ginst27478 (R152_U125, R152_U229, R152_U309);
  and ginst27479 (R152_U126, R152_U287, R152_U389);
  and ginst27480 (R152_U127, R152_U11, R152_U284, R152_U286);
  and ginst27481 (R152_U128, R152_U146, R152_U288);
  and ginst27482 (R152_U129, R152_U223, R152_U303);
  nand ginst27483 (R152_U13, R152_U172, R152_U337);
  and ginst27484 (R152_U130, R152_U338, R152_U339);
  nand ginst27485 (R152_U131, R152_U117, R152_U331);
  and ginst27486 (R152_U132, R152_U345, R152_U346);
  nand ginst27487 (R152_U133, R152_U18, R152_U329);
  and ginst27488 (R152_U134, R152_U352, R152_U353);
  nand ginst27489 (R152_U135, R152_U116, R152_U296);
  and ginst27490 (R152_U136, R152_U359, R152_U360);
  nand ginst27491 (R152_U137, R152_U293, R152_U295);
  and ginst27492 (R152_U138, R152_U366, R152_U367);
  nand ginst27493 (R152_U139, R152_U203, R152_U34);
  not ginst27494 (R152_U14, SI_8_);
  and ginst27495 (R152_U140, R152_U373, R152_U374);
  nand ginst27496 (R152_U141, R152_U118, R152_U315);
  and ginst27497 (R152_U142, R152_U380, R152_U381);
  nand ginst27498 (R152_U143, R152_U29, R152_U310, R152_U311, R152_U312);
  not ginst27499 (R152_U144, U132);
  not ginst27500 (R152_U145, SI_31_);
  and ginst27501 (R152_U146, R152_U392, R152_U393);
  and ginst27502 (R152_U147, R152_U394, R152_U395);
  nand ginst27503 (R152_U148, R152_U283, R152_U284);
  nand ginst27504 (R152_U149, R152_U171, R152_U289, R152_U290);
  not ginst27505 (R152_U15, U127);
  and ginst27506 (R152_U150, R152_U408, R152_U409);
  nand ginst27507 (R152_U151, R152_U279, R152_U280);
  and ginst27508 (R152_U152, R152_U415, R152_U416);
  nand ginst27509 (R152_U153, R152_U275, R152_U276);
  and ginst27510 (R152_U154, R152_U422, R152_U423);
  nand ginst27511 (R152_U155, R152_U271, R152_U272);
  and ginst27512 (R152_U156, R152_U429, R152_U430);
  nand ginst27513 (R152_U157, R152_U267, R152_U268);
  and ginst27514 (R152_U158, R152_U436, R152_U437);
  nand ginst27515 (R152_U159, R152_U263, R152_U264);
  not ginst27516 (R152_U16, SI_7_);
  and ginst27517 (R152_U160, R152_U443, R152_U444);
  nand ginst27518 (R152_U161, R152_U259, R152_U260);
  and ginst27519 (R152_U162, R152_U450, R152_U451);
  nand ginst27520 (R152_U163, R152_U255, R152_U256);
  and ginst27521 (R152_U164, R152_U457, R152_U458);
  nand ginst27522 (R152_U165, R152_U251, R152_U252);
  and ginst27523 (R152_U166, R152_U464, R152_U465);
  nand ginst27524 (R152_U167, R152_U247, R152_U248);
  and ginst27525 (R152_U168, R152_U471, R152_U472);
  nand ginst27526 (R152_U169, R152_U243, R152_U244);
  not ginst27527 (R152_U17, U128);
  nand ginst27528 (R152_U170, SI_0_, U157);
  nand ginst27529 (R152_U171, SI_1_, SI_0_, U157);
  and ginst27530 (R152_U172, R152_U481, R152_U482);
  and ginst27531 (R152_U173, R152_U483, R152_U484);
  nand ginst27532 (R152_U174, R152_U239, R152_U240);
  and ginst27533 (R152_U175, R152_U490, R152_U491);
  nand ginst27534 (R152_U176, R152_U235, R152_U236);
  and ginst27535 (R152_U177, R152_U497, R152_U498);
  nand ginst27536 (R152_U178, R152_U231, R152_U232);
  and ginst27537 (R152_U179, R152_U504, R152_U505);
  nand ginst27538 (R152_U18, SI_7_, U128);
  nand ginst27539 (R152_U180, R152_U125, R152_U327);
  and ginst27540 (R152_U181, R152_U511, R152_U512);
  nand ginst27541 (R152_U182, R152_U308, R152_U325);
  and ginst27542 (R152_U183, R152_U518, R152_U519);
  nand ginst27543 (R152_U184, R152_U306, R152_U323);
  and ginst27544 (R152_U185, R152_U525, R152_U526);
  nand ginst27545 (R152_U186, R152_U129, R152_U321);
  and ginst27546 (R152_U187, R152_U532, R152_U533);
  nand ginst27547 (R152_U188, R152_U319, R152_U48);
  and ginst27548 (R152_U189, R152_U539, R152_U540);
  not ginst27549 (R152_U19, SI_6_);
  nand ginst27550 (R152_U190, R152_U123, R152_U335);
  and ginst27551 (R152_U191, R152_U546, R152_U547);
  nand ginst27552 (R152_U192, R152_U301, R152_U333);
  nand ginst27553 (R152_U193, R152_U126, R152_U148);
  not ginst27554 (R152_U194, R152_U171);
  not ginst27555 (R152_U195, R152_U149);
  or ginst27556 (R152_U196, SI_2_, U145);
  not ginst27557 (R152_U197, R152_U29);
  not ginst27558 (R152_U198, R152_U143);
  or ginst27559 (R152_U199, SI_3_, U134);
  not ginst27560 (R152_U20, U129);
  nand ginst27561 (R152_U200, SI_3_, U134);
  nand ginst27562 (R152_U201, R152_U114, R152_U291);
  or ginst27563 (R152_U202, SI_4_, U131);
  nand ginst27564 (R152_U203, R152_U201, R152_U202);
  not ginst27565 (R152_U204, R152_U34);
  not ginst27566 (R152_U205, R152_U139);
  or ginst27567 (R152_U206, SI_5_, U130);
  nand ginst27568 (R152_U207, SI_5_, U130);
  not ginst27569 (R152_U208, R152_U137);
  or ginst27570 (R152_U209, SI_6_, U129);
  not ginst27571 (R152_U21, SI_3_);
  nand ginst27572 (R152_U210, SI_6_, U129);
  not ginst27573 (R152_U211, R152_U135);
  or ginst27574 (R152_U212, SI_7_, U128);
  not ginst27575 (R152_U213, R152_U18);
  or ginst27576 (R152_U214, SI_8_, U127);
  nand ginst27577 (R152_U215, SI_8_, U127);
  or ginst27578 (R152_U216, SI_9_, U126);
  nand ginst27579 (R152_U217, SI_9_, U126);
  or ginst27580 (R152_U218, SI_10_, U155);
  nand ginst27581 (R152_U219, SI_10_, U155);
  not ginst27582 (R152_U22, U134);
  or ginst27583 (R152_U220, SI_11_, U154);
  not ginst27584 (R152_U221, R152_U48);
  or ginst27585 (R152_U222, SI_12_, U153);
  nand ginst27586 (R152_U223, SI_12_, U153);
  or ginst27587 (R152_U224, SI_13_, U152);
  nand ginst27588 (R152_U225, SI_13_, U152);
  or ginst27589 (R152_U226, SI_14_, U151);
  nand ginst27590 (R152_U227, SI_14_, U151);
  or ginst27591 (R152_U228, SI_15_, U150);
  nand ginst27592 (R152_U229, SI_15_, U150);
  not ginst27593 (R152_U23, SI_1_);
  or ginst27594 (R152_U230, SI_16_, U149);
  nand ginst27595 (R152_U231, R152_U180, R152_U230);
  nand ginst27596 (R152_U232, SI_16_, U149);
  not ginst27597 (R152_U233, R152_U178);
  or ginst27598 (R152_U234, SI_17_, U148);
  nand ginst27599 (R152_U235, R152_U178, R152_U234);
  nand ginst27600 (R152_U236, SI_17_, U148);
  not ginst27601 (R152_U237, R152_U176);
  or ginst27602 (R152_U238, SI_18_, U147);
  nand ginst27603 (R152_U239, R152_U176, R152_U238);
  not ginst27604 (R152_U24, SI_0_);
  nand ginst27605 (R152_U240, SI_18_, U147);
  not ginst27606 (R152_U241, R152_U174);
  or ginst27607 (R152_U242, SI_19_, U146);
  nand ginst27608 (R152_U243, R152_U174, R152_U242);
  nand ginst27609 (R152_U244, SI_19_, U146);
  not ginst27610 (R152_U245, R152_U169);
  or ginst27611 (R152_U246, SI_20_, U144);
  nand ginst27612 (R152_U247, R152_U169, R152_U246);
  nand ginst27613 (R152_U248, SI_20_, U144);
  not ginst27614 (R152_U249, R152_U167);
  not ginst27615 (R152_U25, U157);
  or ginst27616 (R152_U250, SI_21_, U143);
  nand ginst27617 (R152_U251, R152_U167, R152_U250);
  nand ginst27618 (R152_U252, SI_21_, U143);
  not ginst27619 (R152_U253, R152_U165);
  or ginst27620 (R152_U254, SI_22_, U142);
  nand ginst27621 (R152_U255, R152_U165, R152_U254);
  nand ginst27622 (R152_U256, SI_22_, U142);
  not ginst27623 (R152_U257, R152_U163);
  or ginst27624 (R152_U258, SI_23_, U141);
  nand ginst27625 (R152_U259, R152_U163, R152_U258);
  not ginst27626 (R152_U26, U156);
  nand ginst27627 (R152_U260, SI_23_, U141);
  not ginst27628 (R152_U261, R152_U161);
  or ginst27629 (R152_U262, SI_24_, U140);
  nand ginst27630 (R152_U263, R152_U161, R152_U262);
  nand ginst27631 (R152_U264, SI_24_, U140);
  not ginst27632 (R152_U265, R152_U159);
  or ginst27633 (R152_U266, SI_25_, U139);
  nand ginst27634 (R152_U267, R152_U159, R152_U266);
  nand ginst27635 (R152_U268, SI_25_, U139);
  not ginst27636 (R152_U269, R152_U157);
  not ginst27637 (R152_U27, SI_2_);
  or ginst27638 (R152_U270, SI_26_, U138);
  nand ginst27639 (R152_U271, R152_U157, R152_U270);
  nand ginst27640 (R152_U272, SI_26_, U138);
  not ginst27641 (R152_U273, R152_U155);
  or ginst27642 (R152_U274, SI_27_, U137);
  nand ginst27643 (R152_U275, R152_U155, R152_U274);
  nand ginst27644 (R152_U276, SI_27_, U137);
  not ginst27645 (R152_U277, R152_U153);
  or ginst27646 (R152_U278, SI_28_, U136);
  nand ginst27647 (R152_U279, R152_U153, R152_U278);
  not ginst27648 (R152_U28, U145);
  nand ginst27649 (R152_U280, SI_28_, U136);
  not ginst27650 (R152_U281, R152_U151);
  or ginst27651 (R152_U282, SI_29_, U135);
  nand ginst27652 (R152_U283, R152_U151, R152_U282);
  nand ginst27653 (R152_U284, SI_29_, U135);
  not ginst27654 (R152_U285, R152_U148);
  nand ginst27655 (R152_U286, SI_30_, U133);
  or ginst27656 (R152_U287, SI_30_, U133);
  nand ginst27657 (R152_U288, R152_U127, R152_U283);
  nand ginst27658 (R152_U289, SI_0_, U156, U157);
  nand ginst27659 (R152_U29, SI_2_, U145);
  nand ginst27660 (R152_U290, SI_1_, U156);
  nand ginst27661 (R152_U291, R152_U10, R152_U313);
  nand ginst27662 (R152_U292, R152_U197, R152_U199);
  nand ginst27663 (R152_U293, R152_U201, R152_U4);
  nand ginst27664 (R152_U294, R152_U204, R152_U206);
  not ginst27665 (R152_U295, R152_U37);
  nand ginst27666 (R152_U296, R152_U115, R152_U201);
  nand ginst27667 (R152_U297, R152_U209, R152_U37);
  nand ginst27668 (R152_U298, R152_U213, R152_U214);
  nand ginst27669 (R152_U299, R152_U215, R152_U298);
  not ginst27670 (R152_U30, SI_5_);
  nand ginst27671 (R152_U300, R152_U216, R152_U299);
  not ginst27672 (R152_U301, R152_U83);
  nand ginst27673 (R152_U302, R152_U218, R152_U83);
  nand ginst27674 (R152_U303, R152_U221, R152_U222);
  nand ginst27675 (R152_U304, R152_U223, R152_U303);
  nand ginst27676 (R152_U305, R152_U224, R152_U304);
  not ginst27677 (R152_U306, R152_U82);
  nand ginst27678 (R152_U307, R152_U226, R152_U82);
  not ginst27679 (R152_U308, R152_U81);
  nand ginst27680 (R152_U309, R152_U228, R152_U81);
  not ginst27681 (R152_U31, U130);
  nand ginst27682 (R152_U310, SI_0_, R152_U119, R152_U196);
  nand ginst27683 (R152_U311, SI_1_, R152_U120, R152_U196);
  nand ginst27684 (R152_U312, R152_U121, R152_U196);
  nand ginst27685 (R152_U313, R152_U171, R152_U289, R152_U290);
  not ginst27686 (R152_U314, R152_U141);
  nand ginst27687 (R152_U315, R152_U10, R152_U316);
  nand ginst27688 (R152_U316, R152_U290, R152_U317, R152_U318);
  nand ginst27689 (R152_U317, SI_0_, U156, U157);
  nand ginst27690 (R152_U318, SI_1_, SI_0_, U157);
  nand ginst27691 (R152_U319, R152_U190, R152_U220);
  not ginst27692 (R152_U32, SI_4_);
  not ginst27693 (R152_U320, R152_U188);
  nand ginst27694 (R152_U321, R152_U190, R152_U7);
  not ginst27695 (R152_U322, R152_U186);
  nand ginst27696 (R152_U323, R152_U190, R152_U8);
  not ginst27697 (R152_U324, R152_U184);
  nand ginst27698 (R152_U325, R152_U190, R152_U9);
  not ginst27699 (R152_U326, R152_U182);
  nand ginst27700 (R152_U327, R152_U124, R152_U190);
  not ginst27701 (R152_U328, R152_U180);
  nand ginst27702 (R152_U329, R152_U135, R152_U212);
  not ginst27703 (R152_U33, U131);
  not ginst27704 (R152_U330, R152_U133);
  nand ginst27705 (R152_U331, R152_U135, R152_U5);
  not ginst27706 (R152_U332, R152_U131);
  nand ginst27707 (R152_U333, R152_U135, R152_U6);
  not ginst27708 (R152_U334, R152_U192);
  nand ginst27709 (R152_U335, R152_U122, R152_U135);
  not ginst27710 (R152_U336, R152_U190);
  nand ginst27711 (R152_U337, R152_U23, R152_U480);
  nand ginst27712 (R152_U338, R152_U36, U126);
  nand ginst27713 (R152_U339, SI_9_, R152_U35);
  nand ginst27714 (R152_U34, SI_4_, U131);
  nand ginst27715 (R152_U340, R152_U36, U126);
  nand ginst27716 (R152_U341, SI_9_, R152_U35);
  nand ginst27717 (R152_U342, R152_U340, R152_U341);
  nand ginst27718 (R152_U343, R152_U130, R152_U131);
  nand ginst27719 (R152_U344, R152_U332, R152_U342);
  nand ginst27720 (R152_U345, R152_U14, U127);
  nand ginst27721 (R152_U346, SI_8_, R152_U15);
  nand ginst27722 (R152_U347, R152_U14, U127);
  nand ginst27723 (R152_U348, SI_8_, R152_U15);
  nand ginst27724 (R152_U349, R152_U347, R152_U348);
  not ginst27725 (R152_U35, U126);
  nand ginst27726 (R152_U350, R152_U132, R152_U133);
  nand ginst27727 (R152_U351, R152_U330, R152_U349);
  nand ginst27728 (R152_U352, R152_U16, U128);
  nand ginst27729 (R152_U353, SI_7_, R152_U17);
  nand ginst27730 (R152_U354, R152_U16, U128);
  nand ginst27731 (R152_U355, SI_7_, R152_U17);
  nand ginst27732 (R152_U356, R152_U354, R152_U355);
  nand ginst27733 (R152_U357, R152_U134, R152_U135);
  nand ginst27734 (R152_U358, R152_U211, R152_U356);
  nand ginst27735 (R152_U359, R152_U19, U129);
  not ginst27736 (R152_U36, SI_9_);
  nand ginst27737 (R152_U360, SI_6_, R152_U20);
  nand ginst27738 (R152_U361, R152_U19, U129);
  nand ginst27739 (R152_U362, SI_6_, R152_U20);
  nand ginst27740 (R152_U363, R152_U361, R152_U362);
  nand ginst27741 (R152_U364, R152_U136, R152_U137);
  nand ginst27742 (R152_U365, R152_U208, R152_U363);
  nand ginst27743 (R152_U366, R152_U30, U130);
  nand ginst27744 (R152_U367, SI_5_, R152_U31);
  nand ginst27745 (R152_U368, R152_U30, U130);
  nand ginst27746 (R152_U369, SI_5_, R152_U31);
  nand ginst27747 (R152_U37, R152_U207, R152_U294);
  nand ginst27748 (R152_U370, R152_U368, R152_U369);
  nand ginst27749 (R152_U371, R152_U138, R152_U139);
  nand ginst27750 (R152_U372, R152_U205, R152_U370);
  nand ginst27751 (R152_U373, R152_U32, U131);
  nand ginst27752 (R152_U374, SI_4_, R152_U33);
  nand ginst27753 (R152_U375, R152_U32, U131);
  nand ginst27754 (R152_U376, SI_4_, R152_U33);
  nand ginst27755 (R152_U377, R152_U375, R152_U376);
  nand ginst27756 (R152_U378, R152_U140, R152_U141);
  nand ginst27757 (R152_U379, R152_U314, R152_U377);
  not ginst27758 (R152_U38, SI_15_);
  nand ginst27759 (R152_U380, R152_U21, U134);
  nand ginst27760 (R152_U381, SI_3_, R152_U22);
  nand ginst27761 (R152_U382, R152_U21, U134);
  nand ginst27762 (R152_U383, SI_3_, R152_U22);
  nand ginst27763 (R152_U384, R152_U382, R152_U383);
  nand ginst27764 (R152_U385, R152_U142, R152_U143);
  nand ginst27765 (R152_U386, R152_U198, R152_U384);
  nand ginst27766 (R152_U387, R152_U145, U132);
  nand ginst27767 (R152_U388, SI_31_, R152_U144);
  nand ginst27768 (R152_U389, R152_U387, R152_U388);
  not ginst27769 (R152_U39, U150);
  nand ginst27770 (R152_U390, R152_U145, U132);
  nand ginst27771 (R152_U391, SI_31_, R152_U144);
  nand ginst27772 (R152_U392, R152_U11, R152_U79, R152_U80);
  nand ginst27773 (R152_U393, SI_30_, R152_U389, U133);
  nand ginst27774 (R152_U394, R152_U79, U133);
  nand ginst27775 (R152_U395, SI_30_, R152_U80);
  nand ginst27776 (R152_U396, R152_U79, U133);
  nand ginst27777 (R152_U397, SI_30_, R152_U80);
  nand ginst27778 (R152_U398, R152_U396, R152_U397);
  nand ginst27779 (R152_U399, R152_U147, R152_U148);
  and ginst27780 (R152_U4, R152_U202, R152_U206);
  not ginst27781 (R152_U40, SI_14_);
  nand ginst27782 (R152_U400, R152_U285, R152_U398);
  nand ginst27783 (R152_U401, R152_U27, U145);
  nand ginst27784 (R152_U402, SI_2_, R152_U28);
  nand ginst27785 (R152_U403, R152_U27, U145);
  nand ginst27786 (R152_U404, SI_2_, R152_U28);
  nand ginst27787 (R152_U405, R152_U403, R152_U404);
  nand ginst27788 (R152_U406, R152_U149, R152_U401, R152_U402);
  nand ginst27789 (R152_U407, R152_U195, R152_U405);
  nand ginst27790 (R152_U408, R152_U77, U135);
  nand ginst27791 (R152_U409, SI_29_, R152_U78);
  not ginst27792 (R152_U41, U151);
  nand ginst27793 (R152_U410, R152_U77, U135);
  nand ginst27794 (R152_U411, SI_29_, R152_U78);
  nand ginst27795 (R152_U412, R152_U410, R152_U411);
  nand ginst27796 (R152_U413, R152_U150, R152_U151);
  nand ginst27797 (R152_U414, R152_U281, R152_U412);
  nand ginst27798 (R152_U415, R152_U75, U136);
  nand ginst27799 (R152_U416, SI_28_, R152_U76);
  nand ginst27800 (R152_U417, R152_U75, U136);
  nand ginst27801 (R152_U418, SI_28_, R152_U76);
  nand ginst27802 (R152_U419, R152_U417, R152_U418);
  not ginst27803 (R152_U42, SI_13_);
  nand ginst27804 (R152_U420, R152_U152, R152_U153);
  nand ginst27805 (R152_U421, R152_U277, R152_U419);
  nand ginst27806 (R152_U422, R152_U73, U137);
  nand ginst27807 (R152_U423, SI_27_, R152_U74);
  nand ginst27808 (R152_U424, R152_U73, U137);
  nand ginst27809 (R152_U425, SI_27_, R152_U74);
  nand ginst27810 (R152_U426, R152_U424, R152_U425);
  nand ginst27811 (R152_U427, R152_U154, R152_U155);
  nand ginst27812 (R152_U428, R152_U273, R152_U426);
  nand ginst27813 (R152_U429, R152_U71, U138);
  not ginst27814 (R152_U43, U152);
  nand ginst27815 (R152_U430, SI_26_, R152_U72);
  nand ginst27816 (R152_U431, R152_U71, U138);
  nand ginst27817 (R152_U432, SI_26_, R152_U72);
  nand ginst27818 (R152_U433, R152_U431, R152_U432);
  nand ginst27819 (R152_U434, R152_U156, R152_U157);
  nand ginst27820 (R152_U435, R152_U269, R152_U433);
  nand ginst27821 (R152_U436, R152_U69, U139);
  nand ginst27822 (R152_U437, SI_25_, R152_U70);
  nand ginst27823 (R152_U438, R152_U69, U139);
  nand ginst27824 (R152_U439, SI_25_, R152_U70);
  not ginst27825 (R152_U44, SI_12_);
  nand ginst27826 (R152_U440, R152_U438, R152_U439);
  nand ginst27827 (R152_U441, R152_U158, R152_U159);
  nand ginst27828 (R152_U442, R152_U265, R152_U440);
  nand ginst27829 (R152_U443, R152_U67, U140);
  nand ginst27830 (R152_U444, SI_24_, R152_U68);
  nand ginst27831 (R152_U445, R152_U67, U140);
  nand ginst27832 (R152_U446, SI_24_, R152_U68);
  nand ginst27833 (R152_U447, R152_U445, R152_U446);
  nand ginst27834 (R152_U448, R152_U160, R152_U161);
  nand ginst27835 (R152_U449, R152_U261, R152_U447);
  not ginst27836 (R152_U45, U153);
  nand ginst27837 (R152_U450, R152_U65, U141);
  nand ginst27838 (R152_U451, SI_23_, R152_U66);
  nand ginst27839 (R152_U452, R152_U65, U141);
  nand ginst27840 (R152_U453, SI_23_, R152_U66);
  nand ginst27841 (R152_U454, R152_U452, R152_U453);
  nand ginst27842 (R152_U455, R152_U162, R152_U163);
  nand ginst27843 (R152_U456, R152_U257, R152_U454);
  nand ginst27844 (R152_U457, R152_U63, U142);
  nand ginst27845 (R152_U458, SI_22_, R152_U64);
  nand ginst27846 (R152_U459, R152_U63, U142);
  not ginst27847 (R152_U46, SI_11_);
  nand ginst27848 (R152_U460, SI_22_, R152_U64);
  nand ginst27849 (R152_U461, R152_U459, R152_U460);
  nand ginst27850 (R152_U462, R152_U164, R152_U165);
  nand ginst27851 (R152_U463, R152_U253, R152_U461);
  nand ginst27852 (R152_U464, R152_U61, U143);
  nand ginst27853 (R152_U465, SI_21_, R152_U62);
  nand ginst27854 (R152_U466, R152_U61, U143);
  nand ginst27855 (R152_U467, SI_21_, R152_U62);
  nand ginst27856 (R152_U468, R152_U466, R152_U467);
  nand ginst27857 (R152_U469, R152_U166, R152_U167);
  not ginst27858 (R152_U47, U154);
  nand ginst27859 (R152_U470, R152_U249, R152_U468);
  nand ginst27860 (R152_U471, R152_U59, U144);
  nand ginst27861 (R152_U472, SI_20_, R152_U60);
  nand ginst27862 (R152_U473, R152_U59, U144);
  nand ginst27863 (R152_U474, SI_20_, R152_U60);
  nand ginst27864 (R152_U475, R152_U473, R152_U474);
  nand ginst27865 (R152_U476, R152_U168, R152_U169);
  nand ginst27866 (R152_U477, R152_U245, R152_U475);
  nand ginst27867 (R152_U478, R152_U170, U156);
  nand ginst27868 (R152_U479, R152_U120, R152_U26);
  nand ginst27869 (R152_U48, SI_11_, U154);
  nand ginst27870 (R152_U480, R152_U478, R152_U479);
  nand ginst27871 (R152_U481, SI_1_, R152_U170, R152_U26);
  nand ginst27872 (R152_U482, R152_U194, U156);
  nand ginst27873 (R152_U483, R152_U57, U146);
  nand ginst27874 (R152_U484, SI_19_, R152_U58);
  nand ginst27875 (R152_U485, R152_U57, U146);
  nand ginst27876 (R152_U486, SI_19_, R152_U58);
  nand ginst27877 (R152_U487, R152_U485, R152_U486);
  nand ginst27878 (R152_U488, R152_U173, R152_U174);
  nand ginst27879 (R152_U489, R152_U241, R152_U487);
  not ginst27880 (R152_U49, SI_10_);
  nand ginst27881 (R152_U490, R152_U55, U147);
  nand ginst27882 (R152_U491, SI_18_, R152_U56);
  nand ginst27883 (R152_U492, R152_U55, U147);
  nand ginst27884 (R152_U493, SI_18_, R152_U56);
  nand ginst27885 (R152_U494, R152_U492, R152_U493);
  nand ginst27886 (R152_U495, R152_U175, R152_U176);
  nand ginst27887 (R152_U496, R152_U237, R152_U494);
  nand ginst27888 (R152_U497, R152_U53, U148);
  nand ginst27889 (R152_U498, SI_17_, R152_U54);
  nand ginst27890 (R152_U499, R152_U53, U148);
  and ginst27891 (R152_U5, R152_U212, R152_U214);
  not ginst27892 (R152_U50, U155);
  nand ginst27893 (R152_U500, SI_17_, R152_U54);
  nand ginst27894 (R152_U501, R152_U499, R152_U500);
  nand ginst27895 (R152_U502, R152_U177, R152_U178);
  nand ginst27896 (R152_U503, R152_U233, R152_U501);
  nand ginst27897 (R152_U504, R152_U51, U149);
  nand ginst27898 (R152_U505, SI_16_, R152_U52);
  nand ginst27899 (R152_U506, R152_U51, U149);
  nand ginst27900 (R152_U507, SI_16_, R152_U52);
  nand ginst27901 (R152_U508, R152_U506, R152_U507);
  nand ginst27902 (R152_U509, R152_U179, R152_U180);
  not ginst27903 (R152_U51, SI_16_);
  nand ginst27904 (R152_U510, R152_U328, R152_U508);
  nand ginst27905 (R152_U511, R152_U38, U150);
  nand ginst27906 (R152_U512, SI_15_, R152_U39);
  nand ginst27907 (R152_U513, R152_U38, U150);
  nand ginst27908 (R152_U514, SI_15_, R152_U39);
  nand ginst27909 (R152_U515, R152_U513, R152_U514);
  nand ginst27910 (R152_U516, R152_U181, R152_U182);
  nand ginst27911 (R152_U517, R152_U326, R152_U515);
  nand ginst27912 (R152_U518, R152_U40, U151);
  nand ginst27913 (R152_U519, SI_14_, R152_U41);
  not ginst27914 (R152_U52, U149);
  nand ginst27915 (R152_U520, R152_U40, U151);
  nand ginst27916 (R152_U521, SI_14_, R152_U41);
  nand ginst27917 (R152_U522, R152_U520, R152_U521);
  nand ginst27918 (R152_U523, R152_U183, R152_U184);
  nand ginst27919 (R152_U524, R152_U324, R152_U522);
  nand ginst27920 (R152_U525, R152_U42, U152);
  nand ginst27921 (R152_U526, SI_13_, R152_U43);
  nand ginst27922 (R152_U527, R152_U42, U152);
  nand ginst27923 (R152_U528, SI_13_, R152_U43);
  nand ginst27924 (R152_U529, R152_U527, R152_U528);
  not ginst27925 (R152_U53, SI_17_);
  nand ginst27926 (R152_U530, R152_U185, R152_U186);
  nand ginst27927 (R152_U531, R152_U322, R152_U529);
  nand ginst27928 (R152_U532, R152_U44, U153);
  nand ginst27929 (R152_U533, SI_12_, R152_U45);
  nand ginst27930 (R152_U534, R152_U44, U153);
  nand ginst27931 (R152_U535, SI_12_, R152_U45);
  nand ginst27932 (R152_U536, R152_U534, R152_U535);
  nand ginst27933 (R152_U537, R152_U187, R152_U188);
  nand ginst27934 (R152_U538, R152_U320, R152_U536);
  nand ginst27935 (R152_U539, R152_U46, U154);
  not ginst27936 (R152_U54, U148);
  nand ginst27937 (R152_U540, SI_11_, R152_U47);
  nand ginst27938 (R152_U541, R152_U46, U154);
  nand ginst27939 (R152_U542, SI_11_, R152_U47);
  nand ginst27940 (R152_U543, R152_U541, R152_U542);
  nand ginst27941 (R152_U544, R152_U189, R152_U190);
  nand ginst27942 (R152_U545, R152_U336, R152_U543);
  nand ginst27943 (R152_U546, R152_U49, U155);
  nand ginst27944 (R152_U547, SI_10_, R152_U50);
  nand ginst27945 (R152_U548, R152_U49, U155);
  nand ginst27946 (R152_U549, SI_10_, R152_U50);
  not ginst27947 (R152_U55, SI_18_);
  nand ginst27948 (R152_U550, R152_U548, R152_U549);
  nand ginst27949 (R152_U551, R152_U191, R152_U192);
  nand ginst27950 (R152_U552, R152_U334, R152_U550);
  nand ginst27951 (R152_U553, R152_U24, U157);
  nand ginst27952 (R152_U554, SI_0_, R152_U25);
  not ginst27953 (R152_U56, U147);
  not ginst27954 (R152_U57, SI_19_);
  not ginst27955 (R152_U58, U146);
  not ginst27956 (R152_U59, SI_20_);
  and ginst27957 (R152_U6, R152_U216, R152_U5);
  not ginst27958 (R152_U60, U144);
  not ginst27959 (R152_U61, SI_21_);
  not ginst27960 (R152_U62, U143);
  not ginst27961 (R152_U63, SI_22_);
  not ginst27962 (R152_U64, U142);
  not ginst27963 (R152_U65, SI_23_);
  not ginst27964 (R152_U66, U141);
  not ginst27965 (R152_U67, SI_24_);
  not ginst27966 (R152_U68, U140);
  not ginst27967 (R152_U69, SI_25_);
  and ginst27968 (R152_U7, R152_U220, R152_U222);
  not ginst27969 (R152_U70, U139);
  not ginst27970 (R152_U71, SI_26_);
  not ginst27971 (R152_U72, U138);
  not ginst27972 (R152_U73, SI_27_);
  not ginst27973 (R152_U74, U137);
  not ginst27974 (R152_U75, SI_28_);
  not ginst27975 (R152_U76, U136);
  not ginst27976 (R152_U77, SI_29_);
  not ginst27977 (R152_U78, U135);
  not ginst27978 (R152_U79, SI_30_);
  and ginst27979 (R152_U8, R152_U224, R152_U7);
  not ginst27980 (R152_U80, U133);
  nand ginst27981 (R152_U81, R152_U227, R152_U307);
  nand ginst27982 (R152_U82, R152_U225, R152_U305);
  nand ginst27983 (R152_U83, R152_U217, R152_U300);
  nand ginst27984 (R152_U84, R152_U553, R152_U554);
  nand ginst27985 (R152_U85, R152_U343, R152_U344);
  nand ginst27986 (R152_U86, R152_U350, R152_U351);
  nand ginst27987 (R152_U87, R152_U357, R152_U358);
  nand ginst27988 (R152_U88, R152_U364, R152_U365);
  nand ginst27989 (R152_U89, R152_U371, R152_U372);
  and ginst27990 (R152_U9, R152_U226, R152_U8);
  nand ginst27991 (R152_U90, R152_U378, R152_U379);
  nand ginst27992 (R152_U91, R152_U385, R152_U386);
  nand ginst27993 (R152_U92, R152_U399, R152_U400);
  nand ginst27994 (R152_U93, R152_U406, R152_U407);
  nand ginst27995 (R152_U94, R152_U413, R152_U414);
  nand ginst27996 (R152_U95, R152_U420, R152_U421);
  nand ginst27997 (R152_U96, R152_U427, R152_U428);
  nand ginst27998 (R152_U97, R152_U434, R152_U435);
  nand ginst27999 (R152_U98, R152_U441, R152_U442);
  nand ginst28000 (R152_U99, R152_U448, R152_U449);
  not ginst28001 (SUB_1596_U10, ADD_1596_U55);
  nand ginst28002 (SUB_1596_U100, SUB_1596_U20, SUB_1596_U99);
  nand ginst28003 (SUB_1596_U101, ADD_1596_U51, SUB_1596_U100);
  nand ginst28004 (SUB_1596_U102, P2_ADDR_REG_5__SCAN_IN, SUB_1596_U18);
  not ginst28005 (SUB_1596_U103, SUB_1596_U73);
  or ginst28006 (SUB_1596_U104, P2_ADDR_REG_6__SCAN_IN, ADD_1596_U50);
  nand ginst28007 (SUB_1596_U105, SUB_1596_U104, SUB_1596_U73);
  nand ginst28008 (SUB_1596_U106, P2_ADDR_REG_6__SCAN_IN, ADD_1596_U50);
  not ginst28009 (SUB_1596_U107, SUB_1596_U72);
  or ginst28010 (SUB_1596_U108, P2_ADDR_REG_7__SCAN_IN, ADD_1596_U49);
  nand ginst28011 (SUB_1596_U109, SUB_1596_U108, SUB_1596_U72);
  not ginst28012 (SUB_1596_U11, ADD_1596_U54);
  nand ginst28013 (SUB_1596_U110, P2_ADDR_REG_7__SCAN_IN, ADD_1596_U49);
  not ginst28014 (SUB_1596_U111, SUB_1596_U25);
  nand ginst28015 (SUB_1596_U112, SUB_1596_U111, SUB_1596_U27);
  nand ginst28016 (SUB_1596_U113, ADD_1596_U48, SUB_1596_U112);
  nand ginst28017 (SUB_1596_U114, P2_ADDR_REG_8__SCAN_IN, SUB_1596_U25);
  not ginst28018 (SUB_1596_U115, SUB_1596_U71);
  or ginst28019 (SUB_1596_U116, P2_ADDR_REG_9__SCAN_IN, ADD_1596_U47);
  nand ginst28020 (SUB_1596_U117, SUB_1596_U116, SUB_1596_U71);
  nand ginst28021 (SUB_1596_U118, P2_ADDR_REG_9__SCAN_IN, ADD_1596_U47);
  not ginst28022 (SUB_1596_U119, SUB_1596_U30);
  not ginst28023 (SUB_1596_U12, P2_ADDR_REG_2__SCAN_IN);
  nand ginst28024 (SUB_1596_U120, SUB_1596_U119, SUB_1596_U32);
  nand ginst28025 (SUB_1596_U121, ADD_1596_U64, SUB_1596_U120);
  nand ginst28026 (SUB_1596_U122, P2_ADDR_REG_10__SCAN_IN, SUB_1596_U30);
  not ginst28027 (SUB_1596_U123, SUB_1596_U82);
  or ginst28028 (SUB_1596_U124, P2_ADDR_REG_11__SCAN_IN, ADD_1596_U63);
  nand ginst28029 (SUB_1596_U125, SUB_1596_U124, SUB_1596_U82);
  nand ginst28030 (SUB_1596_U126, P2_ADDR_REG_11__SCAN_IN, ADD_1596_U63);
  not ginst28031 (SUB_1596_U127, SUB_1596_U81);
  or ginst28032 (SUB_1596_U128, P2_ADDR_REG_12__SCAN_IN, ADD_1596_U62);
  nand ginst28033 (SUB_1596_U129, SUB_1596_U128, SUB_1596_U81);
  nand ginst28034 (SUB_1596_U13, SUB_1596_U89, SUB_1596_U90);
  nand ginst28035 (SUB_1596_U130, P2_ADDR_REG_12__SCAN_IN, ADD_1596_U62);
  not ginst28036 (SUB_1596_U131, SUB_1596_U37);
  nand ginst28037 (SUB_1596_U132, SUB_1596_U131, SUB_1596_U39);
  nand ginst28038 (SUB_1596_U133, ADD_1596_U61, SUB_1596_U132);
  nand ginst28039 (SUB_1596_U134, P2_ADDR_REG_13__SCAN_IN, SUB_1596_U37);
  not ginst28040 (SUB_1596_U135, SUB_1596_U40);
  nand ginst28041 (SUB_1596_U136, SUB_1596_U135, SUB_1596_U42);
  nand ginst28042 (SUB_1596_U137, ADD_1596_U60, SUB_1596_U136);
  nand ginst28043 (SUB_1596_U138, P2_ADDR_REG_14__SCAN_IN, SUB_1596_U40);
  not ginst28044 (SUB_1596_U139, SUB_1596_U43);
  not ginst28045 (SUB_1596_U14, ADD_1596_U53);
  nand ginst28046 (SUB_1596_U140, SUB_1596_U139, SUB_1596_U45);
  nand ginst28047 (SUB_1596_U141, ADD_1596_U59, SUB_1596_U140);
  nand ginst28048 (SUB_1596_U142, P2_ADDR_REG_15__SCAN_IN, SUB_1596_U43);
  not ginst28049 (SUB_1596_U143, SUB_1596_U80);
  or ginst28050 (SUB_1596_U144, P2_ADDR_REG_16__SCAN_IN, ADD_1596_U58);
  nand ginst28051 (SUB_1596_U145, SUB_1596_U144, SUB_1596_U80);
  nand ginst28052 (SUB_1596_U146, P2_ADDR_REG_16__SCAN_IN, ADD_1596_U58);
  not ginst28053 (SUB_1596_U147, SUB_1596_U79);
  or ginst28054 (SUB_1596_U148, P2_ADDR_REG_17__SCAN_IN, ADD_1596_U57);
  nand ginst28055 (SUB_1596_U149, SUB_1596_U148, SUB_1596_U79);
  not ginst28056 (SUB_1596_U15, P2_ADDR_REG_3__SCAN_IN);
  nand ginst28057 (SUB_1596_U150, P2_ADDR_REG_17__SCAN_IN, ADD_1596_U57);
  not ginst28058 (SUB_1596_U151, SUB_1596_U50);
  nand ginst28059 (SUB_1596_U152, SUB_1596_U151, SUB_1596_U52);
  nand ginst28060 (SUB_1596_U153, ADD_1596_U56, SUB_1596_U152);
  nand ginst28061 (SUB_1596_U154, P2_ADDR_REG_18__SCAN_IN, SUB_1596_U50);
  nand ginst28062 (SUB_1596_U155, SUB_1596_U153, SUB_1596_U154, SUB_1596_U222, SUB_1596_U223);
  nand ginst28063 (SUB_1596_U156, P2_ADDR_REG_18__SCAN_IN, SUB_1596_U50);
  nand ginst28064 (SUB_1596_U157, SUB_1596_U156, SUB_1596_U51);
  nand ginst28065 (SUB_1596_U158, SUB_1596_U151, SUB_1596_U52);
  nand ginst28066 (SUB_1596_U159, SUB_1596_U157, SUB_1596_U158, SUB_1596_U226);
  not ginst28067 (SUB_1596_U16, ADD_1596_U52);
  nand ginst28068 (SUB_1596_U160, SUB_1596_U10, SUB_1596_U219);
  nand ginst28069 (SUB_1596_U161, P2_ADDR_REG_9__SCAN_IN, SUB_1596_U29);
  nand ginst28070 (SUB_1596_U162, ADD_1596_U47, SUB_1596_U28);
  nand ginst28071 (SUB_1596_U163, P2_ADDR_REG_9__SCAN_IN, SUB_1596_U29);
  nand ginst28072 (SUB_1596_U164, ADD_1596_U47, SUB_1596_U28);
  nand ginst28073 (SUB_1596_U165, SUB_1596_U163, SUB_1596_U164);
  nand ginst28074 (SUB_1596_U166, SUB_1596_U161, SUB_1596_U162, SUB_1596_U71);
  nand ginst28075 (SUB_1596_U167, SUB_1596_U115, SUB_1596_U165);
  nand ginst28076 (SUB_1596_U168, P2_ADDR_REG_8__SCAN_IN, SUB_1596_U25);
  nand ginst28077 (SUB_1596_U169, SUB_1596_U111, SUB_1596_U27);
  not ginst28078 (SUB_1596_U17, P2_ADDR_REG_4__SCAN_IN);
  nand ginst28079 (SUB_1596_U170, P2_ADDR_REG_8__SCAN_IN, SUB_1596_U25);
  nand ginst28080 (SUB_1596_U171, SUB_1596_U111, SUB_1596_U27);
  nand ginst28081 (SUB_1596_U172, SUB_1596_U170, SUB_1596_U171);
  nand ginst28082 (SUB_1596_U173, SUB_1596_U168, SUB_1596_U169, SUB_1596_U26);
  nand ginst28083 (SUB_1596_U174, ADD_1596_U48, SUB_1596_U172);
  nand ginst28084 (SUB_1596_U175, P2_ADDR_REG_7__SCAN_IN, SUB_1596_U23);
  nand ginst28085 (SUB_1596_U176, ADD_1596_U49, SUB_1596_U24);
  nand ginst28086 (SUB_1596_U177, P2_ADDR_REG_7__SCAN_IN, SUB_1596_U23);
  nand ginst28087 (SUB_1596_U178, ADD_1596_U49, SUB_1596_U24);
  nand ginst28088 (SUB_1596_U179, SUB_1596_U177, SUB_1596_U178);
  nand ginst28089 (SUB_1596_U18, SUB_1596_U97, SUB_1596_U98);
  nand ginst28090 (SUB_1596_U180, SUB_1596_U175, SUB_1596_U176, SUB_1596_U72);
  nand ginst28091 (SUB_1596_U181, SUB_1596_U107, SUB_1596_U179);
  nand ginst28092 (SUB_1596_U182, P2_ADDR_REG_6__SCAN_IN, SUB_1596_U21);
  nand ginst28093 (SUB_1596_U183, ADD_1596_U50, SUB_1596_U22);
  nand ginst28094 (SUB_1596_U184, P2_ADDR_REG_6__SCAN_IN, SUB_1596_U21);
  nand ginst28095 (SUB_1596_U185, ADD_1596_U50, SUB_1596_U22);
  nand ginst28096 (SUB_1596_U186, SUB_1596_U184, SUB_1596_U185);
  nand ginst28097 (SUB_1596_U187, SUB_1596_U182, SUB_1596_U183, SUB_1596_U73);
  nand ginst28098 (SUB_1596_U188, SUB_1596_U103, SUB_1596_U186);
  nand ginst28099 (SUB_1596_U189, P2_ADDR_REG_5__SCAN_IN, SUB_1596_U18);
  not ginst28100 (SUB_1596_U19, ADD_1596_U51);
  nand ginst28101 (SUB_1596_U190, SUB_1596_U20, SUB_1596_U99);
  nand ginst28102 (SUB_1596_U191, P2_ADDR_REG_5__SCAN_IN, SUB_1596_U18);
  nand ginst28103 (SUB_1596_U192, SUB_1596_U20, SUB_1596_U99);
  nand ginst28104 (SUB_1596_U193, SUB_1596_U191, SUB_1596_U192);
  nand ginst28105 (SUB_1596_U194, SUB_1596_U189, SUB_1596_U19, SUB_1596_U190);
  nand ginst28106 (SUB_1596_U195, ADD_1596_U51, SUB_1596_U193);
  nand ginst28107 (SUB_1596_U196, P2_ADDR_REG_4__SCAN_IN, SUB_1596_U16);
  nand ginst28108 (SUB_1596_U197, ADD_1596_U52, SUB_1596_U17);
  nand ginst28109 (SUB_1596_U198, P2_ADDR_REG_4__SCAN_IN, SUB_1596_U16);
  nand ginst28110 (SUB_1596_U199, ADD_1596_U52, SUB_1596_U17);
  not ginst28111 (SUB_1596_U20, P2_ADDR_REG_5__SCAN_IN);
  nand ginst28112 (SUB_1596_U200, SUB_1596_U198, SUB_1596_U199);
  nand ginst28113 (SUB_1596_U201, SUB_1596_U196, SUB_1596_U197, SUB_1596_U74);
  nand ginst28114 (SUB_1596_U202, SUB_1596_U200, SUB_1596_U95);
  nand ginst28115 (SUB_1596_U203, P2_ADDR_REG_3__SCAN_IN, SUB_1596_U13);
  nand ginst28116 (SUB_1596_U204, SUB_1596_U15, SUB_1596_U91);
  nand ginst28117 (SUB_1596_U205, P2_ADDR_REG_3__SCAN_IN, SUB_1596_U13);
  nand ginst28118 (SUB_1596_U206, SUB_1596_U15, SUB_1596_U91);
  nand ginst28119 (SUB_1596_U207, SUB_1596_U205, SUB_1596_U206);
  nand ginst28120 (SUB_1596_U208, SUB_1596_U14, SUB_1596_U203, SUB_1596_U204);
  nand ginst28121 (SUB_1596_U209, ADD_1596_U53, SUB_1596_U207);
  not ginst28122 (SUB_1596_U21, ADD_1596_U50);
  nand ginst28123 (SUB_1596_U210, P2_ADDR_REG_2__SCAN_IN, SUB_1596_U11);
  nand ginst28124 (SUB_1596_U211, ADD_1596_U54, SUB_1596_U12);
  nand ginst28125 (SUB_1596_U212, P2_ADDR_REG_2__SCAN_IN, SUB_1596_U11);
  nand ginst28126 (SUB_1596_U213, ADD_1596_U54, SUB_1596_U12);
  nand ginst28127 (SUB_1596_U214, SUB_1596_U212, SUB_1596_U213);
  nand ginst28128 (SUB_1596_U215, SUB_1596_U210, SUB_1596_U211, SUB_1596_U75);
  nand ginst28129 (SUB_1596_U216, SUB_1596_U214, SUB_1596_U87);
  nand ginst28130 (SUB_1596_U217, P2_ADDR_REG_1__SCAN_IN, SUB_1596_U9);
  nand ginst28131 (SUB_1596_U218, SUB_1596_U8, SUB_1596_U84);
  nand ginst28132 (SUB_1596_U219, SUB_1596_U217, SUB_1596_U218);
  not ginst28133 (SUB_1596_U22, P2_ADDR_REG_6__SCAN_IN);
  nand ginst28134 (SUB_1596_U220, ADD_1596_U55, SUB_1596_U8, SUB_1596_U9);
  nand ginst28135 (SUB_1596_U221, P2_ADDR_REG_1__SCAN_IN, SUB_1596_U83);
  nand ginst28136 (SUB_1596_U222, P2_ADDR_REG_19__SCAN_IN, SUB_1596_U78);
  nand ginst28137 (SUB_1596_U223, ADD_1596_U6, SUB_1596_U77);
  nand ginst28138 (SUB_1596_U224, P2_ADDR_REG_19__SCAN_IN, SUB_1596_U78);
  nand ginst28139 (SUB_1596_U225, ADD_1596_U6, SUB_1596_U77);
  nand ginst28140 (SUB_1596_U226, SUB_1596_U224, SUB_1596_U225);
  nand ginst28141 (SUB_1596_U227, P2_ADDR_REG_18__SCAN_IN, SUB_1596_U50);
  nand ginst28142 (SUB_1596_U228, SUB_1596_U151, SUB_1596_U52);
  nand ginst28143 (SUB_1596_U229, P2_ADDR_REG_18__SCAN_IN, SUB_1596_U50);
  not ginst28144 (SUB_1596_U23, ADD_1596_U49);
  nand ginst28145 (SUB_1596_U230, SUB_1596_U151, SUB_1596_U52);
  nand ginst28146 (SUB_1596_U231, SUB_1596_U229, SUB_1596_U230);
  nand ginst28147 (SUB_1596_U232, SUB_1596_U227, SUB_1596_U228, SUB_1596_U51);
  nand ginst28148 (SUB_1596_U233, ADD_1596_U56, SUB_1596_U231);
  nand ginst28149 (SUB_1596_U234, P2_ADDR_REG_17__SCAN_IN, SUB_1596_U48);
  nand ginst28150 (SUB_1596_U235, ADD_1596_U57, SUB_1596_U49);
  nand ginst28151 (SUB_1596_U236, P2_ADDR_REG_17__SCAN_IN, SUB_1596_U48);
  nand ginst28152 (SUB_1596_U237, ADD_1596_U57, SUB_1596_U49);
  nand ginst28153 (SUB_1596_U238, SUB_1596_U236, SUB_1596_U237);
  nand ginst28154 (SUB_1596_U239, SUB_1596_U234, SUB_1596_U235, SUB_1596_U79);
  not ginst28155 (SUB_1596_U24, P2_ADDR_REG_7__SCAN_IN);
  nand ginst28156 (SUB_1596_U240, SUB_1596_U147, SUB_1596_U238);
  nand ginst28157 (SUB_1596_U241, P2_ADDR_REG_16__SCAN_IN, SUB_1596_U46);
  nand ginst28158 (SUB_1596_U242, ADD_1596_U58, SUB_1596_U47);
  nand ginst28159 (SUB_1596_U243, P2_ADDR_REG_16__SCAN_IN, SUB_1596_U46);
  nand ginst28160 (SUB_1596_U244, ADD_1596_U58, SUB_1596_U47);
  nand ginst28161 (SUB_1596_U245, SUB_1596_U243, SUB_1596_U244);
  nand ginst28162 (SUB_1596_U246, SUB_1596_U241, SUB_1596_U242, SUB_1596_U80);
  nand ginst28163 (SUB_1596_U247, SUB_1596_U143, SUB_1596_U245);
  nand ginst28164 (SUB_1596_U248, P2_ADDR_REG_15__SCAN_IN, SUB_1596_U43);
  nand ginst28165 (SUB_1596_U249, SUB_1596_U139, SUB_1596_U45);
  nand ginst28166 (SUB_1596_U25, SUB_1596_U109, SUB_1596_U110);
  nand ginst28167 (SUB_1596_U250, P2_ADDR_REG_15__SCAN_IN, SUB_1596_U43);
  nand ginst28168 (SUB_1596_U251, SUB_1596_U139, SUB_1596_U45);
  nand ginst28169 (SUB_1596_U252, SUB_1596_U250, SUB_1596_U251);
  nand ginst28170 (SUB_1596_U253, SUB_1596_U248, SUB_1596_U249, SUB_1596_U44);
  nand ginst28171 (SUB_1596_U254, ADD_1596_U59, SUB_1596_U252);
  nand ginst28172 (SUB_1596_U255, P2_ADDR_REG_14__SCAN_IN, SUB_1596_U40);
  nand ginst28173 (SUB_1596_U256, SUB_1596_U135, SUB_1596_U42);
  nand ginst28174 (SUB_1596_U257, P2_ADDR_REG_14__SCAN_IN, SUB_1596_U40);
  nand ginst28175 (SUB_1596_U258, SUB_1596_U135, SUB_1596_U42);
  nand ginst28176 (SUB_1596_U259, SUB_1596_U257, SUB_1596_U258);
  not ginst28177 (SUB_1596_U26, ADD_1596_U48);
  nand ginst28178 (SUB_1596_U260, SUB_1596_U255, SUB_1596_U256, SUB_1596_U41);
  nand ginst28179 (SUB_1596_U261, ADD_1596_U60, SUB_1596_U259);
  nand ginst28180 (SUB_1596_U262, P2_ADDR_REG_13__SCAN_IN, SUB_1596_U37);
  nand ginst28181 (SUB_1596_U263, SUB_1596_U131, SUB_1596_U39);
  nand ginst28182 (SUB_1596_U264, P2_ADDR_REG_13__SCAN_IN, SUB_1596_U37);
  nand ginst28183 (SUB_1596_U265, SUB_1596_U131, SUB_1596_U39);
  nand ginst28184 (SUB_1596_U266, SUB_1596_U264, SUB_1596_U265);
  nand ginst28185 (SUB_1596_U267, SUB_1596_U262, SUB_1596_U263, SUB_1596_U38);
  nand ginst28186 (SUB_1596_U268, ADD_1596_U61, SUB_1596_U266);
  nand ginst28187 (SUB_1596_U269, P2_ADDR_REG_12__SCAN_IN, SUB_1596_U35);
  not ginst28188 (SUB_1596_U27, P2_ADDR_REG_8__SCAN_IN);
  nand ginst28189 (SUB_1596_U270, ADD_1596_U62, SUB_1596_U36);
  nand ginst28190 (SUB_1596_U271, P2_ADDR_REG_12__SCAN_IN, SUB_1596_U35);
  nand ginst28191 (SUB_1596_U272, ADD_1596_U62, SUB_1596_U36);
  nand ginst28192 (SUB_1596_U273, SUB_1596_U271, SUB_1596_U272);
  nand ginst28193 (SUB_1596_U274, SUB_1596_U269, SUB_1596_U270, SUB_1596_U81);
  nand ginst28194 (SUB_1596_U275, SUB_1596_U127, SUB_1596_U273);
  nand ginst28195 (SUB_1596_U276, P2_ADDR_REG_11__SCAN_IN, SUB_1596_U33);
  nand ginst28196 (SUB_1596_U277, ADD_1596_U63, SUB_1596_U34);
  nand ginst28197 (SUB_1596_U278, P2_ADDR_REG_11__SCAN_IN, SUB_1596_U33);
  nand ginst28198 (SUB_1596_U279, ADD_1596_U63, SUB_1596_U34);
  not ginst28199 (SUB_1596_U28, P2_ADDR_REG_9__SCAN_IN);
  nand ginst28200 (SUB_1596_U280, SUB_1596_U278, SUB_1596_U279);
  nand ginst28201 (SUB_1596_U281, SUB_1596_U276, SUB_1596_U277, SUB_1596_U82);
  nand ginst28202 (SUB_1596_U282, SUB_1596_U123, SUB_1596_U280);
  nand ginst28203 (SUB_1596_U283, P2_ADDR_REG_10__SCAN_IN, SUB_1596_U30);
  nand ginst28204 (SUB_1596_U284, SUB_1596_U119, SUB_1596_U32);
  nand ginst28205 (SUB_1596_U285, P2_ADDR_REG_10__SCAN_IN, SUB_1596_U30);
  nand ginst28206 (SUB_1596_U286, SUB_1596_U119, SUB_1596_U32);
  nand ginst28207 (SUB_1596_U287, SUB_1596_U285, SUB_1596_U286);
  nand ginst28208 (SUB_1596_U288, SUB_1596_U283, SUB_1596_U284, SUB_1596_U31);
  nand ginst28209 (SUB_1596_U289, ADD_1596_U64, SUB_1596_U287);
  not ginst28210 (SUB_1596_U29, ADD_1596_U47);
  nand ginst28211 (SUB_1596_U290, P2_ADDR_REG_0__SCAN_IN, SUB_1596_U6);
  nand ginst28212 (SUB_1596_U291, ADD_1596_U7, SUB_1596_U7);
  nand ginst28213 (SUB_1596_U30, SUB_1596_U117, SUB_1596_U118);
  not ginst28214 (SUB_1596_U31, ADD_1596_U64);
  not ginst28215 (SUB_1596_U32, P2_ADDR_REG_10__SCAN_IN);
  not ginst28216 (SUB_1596_U33, ADD_1596_U63);
  not ginst28217 (SUB_1596_U34, P2_ADDR_REG_11__SCAN_IN);
  not ginst28218 (SUB_1596_U35, ADD_1596_U62);
  not ginst28219 (SUB_1596_U36, P2_ADDR_REG_12__SCAN_IN);
  nand ginst28220 (SUB_1596_U37, SUB_1596_U129, SUB_1596_U130);
  not ginst28221 (SUB_1596_U38, ADD_1596_U61);
  not ginst28222 (SUB_1596_U39, P2_ADDR_REG_13__SCAN_IN);
  and ginst28223 (SUB_1596_U4, SUB_1596_U155, SUB_1596_U159);
  nand ginst28224 (SUB_1596_U40, SUB_1596_U133, SUB_1596_U134);
  not ginst28225 (SUB_1596_U41, ADD_1596_U60);
  not ginst28226 (SUB_1596_U42, P2_ADDR_REG_14__SCAN_IN);
  nand ginst28227 (SUB_1596_U43, SUB_1596_U137, SUB_1596_U138);
  not ginst28228 (SUB_1596_U44, ADD_1596_U59);
  not ginst28229 (SUB_1596_U45, P2_ADDR_REG_15__SCAN_IN);
  not ginst28230 (SUB_1596_U46, ADD_1596_U58);
  not ginst28231 (SUB_1596_U47, P2_ADDR_REG_16__SCAN_IN);
  not ginst28232 (SUB_1596_U48, ADD_1596_U57);
  not ginst28233 (SUB_1596_U49, P2_ADDR_REG_17__SCAN_IN);
  nand ginst28234 (SUB_1596_U5, SUB_1596_U160, SUB_1596_U220, SUB_1596_U221);
  nand ginst28235 (SUB_1596_U50, SUB_1596_U149, SUB_1596_U150);
  not ginst28236 (SUB_1596_U51, ADD_1596_U56);
  not ginst28237 (SUB_1596_U52, P2_ADDR_REG_18__SCAN_IN);
  nand ginst28238 (SUB_1596_U53, SUB_1596_U290, SUB_1596_U291);
  nand ginst28239 (SUB_1596_U54, SUB_1596_U166, SUB_1596_U167);
  nand ginst28240 (SUB_1596_U55, SUB_1596_U173, SUB_1596_U174);
  nand ginst28241 (SUB_1596_U56, SUB_1596_U180, SUB_1596_U181);
  nand ginst28242 (SUB_1596_U57, SUB_1596_U187, SUB_1596_U188);
  nand ginst28243 (SUB_1596_U58, SUB_1596_U194, SUB_1596_U195);
  nand ginst28244 (SUB_1596_U59, SUB_1596_U201, SUB_1596_U202);
  not ginst28245 (SUB_1596_U6, ADD_1596_U7);
  nand ginst28246 (SUB_1596_U60, SUB_1596_U208, SUB_1596_U209);
  nand ginst28247 (SUB_1596_U61, SUB_1596_U215, SUB_1596_U216);
  nand ginst28248 (SUB_1596_U62, SUB_1596_U232, SUB_1596_U233);
  nand ginst28249 (SUB_1596_U63, SUB_1596_U239, SUB_1596_U240);
  nand ginst28250 (SUB_1596_U64, SUB_1596_U246, SUB_1596_U247);
  nand ginst28251 (SUB_1596_U65, SUB_1596_U253, SUB_1596_U254);
  nand ginst28252 (SUB_1596_U66, SUB_1596_U260, SUB_1596_U261);
  nand ginst28253 (SUB_1596_U67, SUB_1596_U267, SUB_1596_U268);
  nand ginst28254 (SUB_1596_U68, SUB_1596_U274, SUB_1596_U275);
  nand ginst28255 (SUB_1596_U69, SUB_1596_U281, SUB_1596_U282);
  not ginst28256 (SUB_1596_U7, P2_ADDR_REG_0__SCAN_IN);
  nand ginst28257 (SUB_1596_U70, SUB_1596_U288, SUB_1596_U289);
  nand ginst28258 (SUB_1596_U71, SUB_1596_U113, SUB_1596_U114);
  nand ginst28259 (SUB_1596_U72, SUB_1596_U105, SUB_1596_U106);
  nand ginst28260 (SUB_1596_U73, SUB_1596_U101, SUB_1596_U102);
  nand ginst28261 (SUB_1596_U74, SUB_1596_U93, SUB_1596_U94);
  nand ginst28262 (SUB_1596_U75, SUB_1596_U76, SUB_1596_U86);
  nand ginst28263 (SUB_1596_U76, ADD_1596_U55, SUB_1596_U84);
  not ginst28264 (SUB_1596_U77, P2_ADDR_REG_19__SCAN_IN);
  not ginst28265 (SUB_1596_U78, ADD_1596_U6);
  nand ginst28266 (SUB_1596_U79, SUB_1596_U145, SUB_1596_U146);
  not ginst28267 (SUB_1596_U8, P2_ADDR_REG_1__SCAN_IN);
  nand ginst28268 (SUB_1596_U80, SUB_1596_U141, SUB_1596_U142);
  nand ginst28269 (SUB_1596_U81, SUB_1596_U125, SUB_1596_U126);
  nand ginst28270 (SUB_1596_U82, SUB_1596_U121, SUB_1596_U122);
  not ginst28271 (SUB_1596_U83, SUB_1596_U76);
  not ginst28272 (SUB_1596_U84, SUB_1596_U9);
  nand ginst28273 (SUB_1596_U85, SUB_1596_U10, SUB_1596_U9);
  nand ginst28274 (SUB_1596_U86, P2_ADDR_REG_1__SCAN_IN, SUB_1596_U85);
  not ginst28275 (SUB_1596_U87, SUB_1596_U75);
  or ginst28276 (SUB_1596_U88, P2_ADDR_REG_2__SCAN_IN, ADD_1596_U54);
  nand ginst28277 (SUB_1596_U89, SUB_1596_U75, SUB_1596_U88);
  nand ginst28278 (SUB_1596_U9, P2_ADDR_REG_0__SCAN_IN, ADD_1596_U7);
  nand ginst28279 (SUB_1596_U90, P2_ADDR_REG_2__SCAN_IN, ADD_1596_U54);
  not ginst28280 (SUB_1596_U91, SUB_1596_U13);
  nand ginst28281 (SUB_1596_U92, SUB_1596_U15, SUB_1596_U91);
  nand ginst28282 (SUB_1596_U93, ADD_1596_U53, SUB_1596_U92);
  nand ginst28283 (SUB_1596_U94, P2_ADDR_REG_3__SCAN_IN, SUB_1596_U13);
  not ginst28284 (SUB_1596_U95, SUB_1596_U74);
  or ginst28285 (SUB_1596_U96, P2_ADDR_REG_4__SCAN_IN, ADD_1596_U52);
  nand ginst28286 (SUB_1596_U97, SUB_1596_U74, SUB_1596_U96);
  nand ginst28287 (SUB_1596_U98, P2_ADDR_REG_4__SCAN_IN, ADD_1596_U52);
  not ginst28288 (SUB_1596_U99, SUB_1596_U18);
  and ginst28289 (SUB_1605_U10, SUB_1605_U215, SUB_1605_U9);
  nand ginst28290 (SUB_1605_U100, SUB_1605_U439, SUB_1605_U440);
  nand ginst28291 (SUB_1605_U101, SUB_1605_U444, SUB_1605_U445);
  nand ginst28292 (SUB_1605_U102, SUB_1605_U449, SUB_1605_U450);
  nand ginst28293 (SUB_1605_U103, SUB_1605_U454, SUB_1605_U455);
  nand ginst28294 (SUB_1605_U104, SUB_1605_U459, SUB_1605_U460);
  nand ginst28295 (SUB_1605_U105, SUB_1605_U464, SUB_1605_U465);
  nand ginst28296 (SUB_1605_U106, SUB_1605_U469, SUB_1605_U470);
  nand ginst28297 (SUB_1605_U107, SUB_1605_U474, SUB_1605_U475);
  nand ginst28298 (SUB_1605_U108, SUB_1605_U479, SUB_1605_U480);
  and ginst28299 (SUB_1605_U109, P1_DATAO_REG_5__SCAN_IN, SUB_1605_U30);
  and ginst28300 (SUB_1605_U11, SUB_1605_U362, SUB_1605_U363);
  and ginst28301 (SUB_1605_U110, SUB_1605_U203, SUB_1605_U205);
  and ginst28302 (SUB_1605_U111, SUB_1605_U197, SUB_1605_U6);
  and ginst28303 (SUB_1605_U112, SUB_1605_U197, SUB_1605_U299);
  and ginst28304 (SUB_1605_U113, SUB_1605_U198, SUB_1605_U298);
  and ginst28305 (SUB_1605_U114, SUB_1605_U206, SUB_1605_U8);
  and ginst28306 (SUB_1605_U115, SUB_1605_U207, SUB_1605_U302);
  nand ginst28307 (SUB_1605_U116, SUB_1605_U324, SUB_1605_U325);
  nand ginst28308 (SUB_1605_U117, SUB_1605_U329, SUB_1605_U330);
  and ginst28309 (SUB_1605_U118, SUB_1605_U203, SUB_1605_U300);
  nand ginst28310 (SUB_1605_U119, SUB_1605_U334, SUB_1605_U335);
  nand ginst28311 (SUB_1605_U12, SUB_1605_U128, SUB_1605_U323);
  nand ginst28312 (SUB_1605_U120, SUB_1605_U339, SUB_1605_U340);
  nand ginst28313 (SUB_1605_U121, SUB_1605_U344, SUB_1605_U345);
  nand ginst28314 (SUB_1605_U122, SUB_1605_U349, SUB_1605_U350);
  nand ginst28315 (SUB_1605_U123, SUB_1605_U354, SUB_1605_U355);
  and ginst28316 (SUB_1605_U124, SUB_1605_U10, SUB_1605_U218);
  and ginst28317 (SUB_1605_U125, SUB_1605_U219, SUB_1605_U311);
  and ginst28318 (SUB_1605_U126, SUB_1605_U11, SUB_1605_U287, SUB_1605_U290);
  and ginst28319 (SUB_1605_U127, SUB_1605_U289, SUB_1605_U361);
  and ginst28320 (SUB_1605_U128, SUB_1605_U161, SUB_1605_U293);
  nand ginst28321 (SUB_1605_U129, SUB_1605_U366, SUB_1605_U367);
  nand ginst28322 (SUB_1605_U13, SUB_1605_U175, SUB_1605_U291);
  nand ginst28323 (SUB_1605_U130, SUB_1605_U371, SUB_1605_U372);
  nand ginst28324 (SUB_1605_U131, SUB_1605_U376, SUB_1605_U377);
  nand ginst28325 (SUB_1605_U132, SUB_1605_U381, SUB_1605_U382);
  nand ginst28326 (SUB_1605_U133, SUB_1605_U386, SUB_1605_U387);
  nand ginst28327 (SUB_1605_U134, SUB_1605_U391, SUB_1605_U392);
  nand ginst28328 (SUB_1605_U135, SUB_1605_U396, SUB_1605_U397);
  nand ginst28329 (SUB_1605_U136, SUB_1605_U401, SUB_1605_U402);
  nand ginst28330 (SUB_1605_U137, SUB_1605_U406, SUB_1605_U407);
  nand ginst28331 (SUB_1605_U138, SUB_1605_U411, SUB_1605_U412);
  nand ginst28332 (SUB_1605_U139, SUB_1605_U416, SUB_1605_U417);
  not ginst28333 (SUB_1605_U14, P1_DATAO_REG_8__SCAN_IN);
  nand ginst28334 (SUB_1605_U140, SUB_1605_U421, SUB_1605_U422);
  nand ginst28335 (SUB_1605_U141, SUB_1605_U426, SUB_1605_U427);
  nand ginst28336 (SUB_1605_U142, SUB_1605_U431, SUB_1605_U432);
  nand ginst28337 (SUB_1605_U143, SUB_1605_U436, SUB_1605_U437);
  nand ginst28338 (SUB_1605_U144, SUB_1605_U441, SUB_1605_U442);
  nand ginst28339 (SUB_1605_U145, SUB_1605_U446, SUB_1605_U447);
  nand ginst28340 (SUB_1605_U146, SUB_1605_U451, SUB_1605_U452);
  nand ginst28341 (SUB_1605_U147, SUB_1605_U456, SUB_1605_U457);
  nand ginst28342 (SUB_1605_U148, SUB_1605_U461, SUB_1605_U462);
  nand ginst28343 (SUB_1605_U149, SUB_1605_U466, SUB_1605_U467);
  not ginst28344 (SUB_1605_U15, P2_DATAO_REG_8__SCAN_IN);
  nand ginst28345 (SUB_1605_U150, SUB_1605_U471, SUB_1605_U472);
  nand ginst28346 (SUB_1605_U151, SUB_1605_U476, SUB_1605_U477);
  nand ginst28347 (SUB_1605_U152, SUB_1605_U115, SUB_1605_U321);
  nand ginst28348 (SUB_1605_U153, SUB_1605_U21, SUB_1605_U319);
  nand ginst28349 (SUB_1605_U154, SUB_1605_U118, SUB_1605_U317);
  nand ginst28350 (SUB_1605_U155, SUB_1605_U201, SUB_1605_U315);
  nand ginst28351 (SUB_1605_U156, SUB_1605_U113, SUB_1605_U297);
  nand ginst28352 (SUB_1605_U157, SUB_1605_U294, SUB_1605_U296);
  nand ginst28353 (SUB_1605_U158, SUB_1605_U191, SUB_1605_U192);
  not ginst28354 (SUB_1605_U159, P2_DATAO_REG_31__SCAN_IN);
  not ginst28355 (SUB_1605_U16, P2_DATAO_REG_7__SCAN_IN);
  not ginst28356 (SUB_1605_U160, P1_DATAO_REG_31__SCAN_IN);
  and ginst28357 (SUB_1605_U161, SUB_1605_U364, SUB_1605_U365);
  nand ginst28358 (SUB_1605_U162, SUB_1605_U286, SUB_1605_U287);
  nand ginst28359 (SUB_1605_U163, SUB_1605_U186, SUB_1605_U188, SUB_1605_U292);
  nand ginst28360 (SUB_1605_U164, SUB_1605_U282, SUB_1605_U283);
  nand ginst28361 (SUB_1605_U165, SUB_1605_U278, SUB_1605_U279);
  nand ginst28362 (SUB_1605_U166, SUB_1605_U274, SUB_1605_U275);
  nand ginst28363 (SUB_1605_U167, SUB_1605_U270, SUB_1605_U271);
  nand ginst28364 (SUB_1605_U168, SUB_1605_U266, SUB_1605_U267);
  nand ginst28365 (SUB_1605_U169, SUB_1605_U262, SUB_1605_U263);
  not ginst28366 (SUB_1605_U17, P1_DATAO_REG_6__SCAN_IN);
  nand ginst28367 (SUB_1605_U170, SUB_1605_U258, SUB_1605_U259);
  nand ginst28368 (SUB_1605_U171, SUB_1605_U254, SUB_1605_U255);
  nand ginst28369 (SUB_1605_U172, SUB_1605_U250, SUB_1605_U251);
  nand ginst28370 (SUB_1605_U173, SUB_1605_U246, SUB_1605_U247);
  not ginst28371 (SUB_1605_U174, P2_DATAO_REG_1__SCAN_IN);
  nand ginst28372 (SUB_1605_U175, P2_DATAO_REG_0__SCAN_IN, SUB_1605_U78);
  nand ginst28373 (SUB_1605_U176, SUB_1605_U242, SUB_1605_U243);
  nand ginst28374 (SUB_1605_U177, SUB_1605_U238, SUB_1605_U239);
  nand ginst28375 (SUB_1605_U178, SUB_1605_U234, SUB_1605_U235);
  nand ginst28376 (SUB_1605_U179, SUB_1605_U230, SUB_1605_U231);
  not ginst28377 (SUB_1605_U18, P1_DATAO_REG_7__SCAN_IN);
  nand ginst28378 (SUB_1605_U180, SUB_1605_U226, SUB_1605_U227);
  nand ginst28379 (SUB_1605_U181, SUB_1605_U222, SUB_1605_U223);
  nand ginst28380 (SUB_1605_U182, SUB_1605_U125, SUB_1605_U310);
  nand ginst28381 (SUB_1605_U183, SUB_1605_U307, SUB_1605_U309);
  nand ginst28382 (SUB_1605_U184, SUB_1605_U304, SUB_1605_U306);
  nand ginst28383 (SUB_1605_U185, SUB_1605_U209, SUB_1605_U39);
  nand ginst28384 (SUB_1605_U186, SUB_1605_U174, SUB_1605_U175);
  not ginst28385 (SUB_1605_U187, SUB_1605_U175);
  nand ginst28386 (SUB_1605_U188, P1_DATAO_REG_1__SCAN_IN, SUB_1605_U175);
  not ginst28387 (SUB_1605_U189, SUB_1605_U163);
  not ginst28388 (SUB_1605_U19, P2_DATAO_REG_6__SCAN_IN);
  nand ginst28389 (SUB_1605_U190, P2_DATAO_REG_2__SCAN_IN, SUB_1605_U28);
  nand ginst28390 (SUB_1605_U191, SUB_1605_U190, SUB_1605_U312);
  nand ginst28391 (SUB_1605_U192, P1_DATAO_REG_2__SCAN_IN, SUB_1605_U26);
  not ginst28392 (SUB_1605_U193, SUB_1605_U158);
  nand ginst28393 (SUB_1605_U194, P2_DATAO_REG_3__SCAN_IN, SUB_1605_U29);
  nand ginst28394 (SUB_1605_U195, P1_DATAO_REG_3__SCAN_IN, SUB_1605_U27);
  not ginst28395 (SUB_1605_U196, SUB_1605_U157);
  nand ginst28396 (SUB_1605_U197, P2_DATAO_REG_4__SCAN_IN, SUB_1605_U22);
  nand ginst28397 (SUB_1605_U198, P1_DATAO_REG_4__SCAN_IN, SUB_1605_U25);
  not ginst28398 (SUB_1605_U199, SUB_1605_U156);
  not ginst28399 (SUB_1605_U20, P1_DATAO_REG_5__SCAN_IN);
  nand ginst28400 (SUB_1605_U200, P2_DATAO_REG_5__SCAN_IN, SUB_1605_U20);
  nand ginst28401 (SUB_1605_U201, P1_DATAO_REG_5__SCAN_IN, SUB_1605_U30);
  nand ginst28402 (SUB_1605_U202, P2_DATAO_REG_6__SCAN_IN, SUB_1605_U17);
  nand ginst28403 (SUB_1605_U203, P1_DATAO_REG_6__SCAN_IN, SUB_1605_U19);
  nand ginst28404 (SUB_1605_U204, P2_DATAO_REG_7__SCAN_IN, SUB_1605_U18);
  nand ginst28405 (SUB_1605_U205, P1_DATAO_REG_7__SCAN_IN, SUB_1605_U16);
  nand ginst28406 (SUB_1605_U206, P2_DATAO_REG_8__SCAN_IN, SUB_1605_U14);
  nand ginst28407 (SUB_1605_U207, P1_DATAO_REG_8__SCAN_IN, SUB_1605_U15);
  nand ginst28408 (SUB_1605_U208, P2_DATAO_REG_9__SCAN_IN, SUB_1605_U32);
  nand ginst28409 (SUB_1605_U209, SUB_1605_U152, SUB_1605_U208);
  nand ginst28410 (SUB_1605_U21, SUB_1605_U204, SUB_1605_U303);
  not ginst28411 (SUB_1605_U210, SUB_1605_U39);
  not ginst28412 (SUB_1605_U211, SUB_1605_U185);
  nand ginst28413 (SUB_1605_U212, P2_DATAO_REG_10__SCAN_IN, SUB_1605_U38);
  nand ginst28414 (SUB_1605_U213, P1_DATAO_REG_10__SCAN_IN, SUB_1605_U36);
  not ginst28415 (SUB_1605_U214, SUB_1605_U184);
  nand ginst28416 (SUB_1605_U215, P2_DATAO_REG_11__SCAN_IN, SUB_1605_U37);
  nand ginst28417 (SUB_1605_U216, P1_DATAO_REG_11__SCAN_IN, SUB_1605_U35);
  not ginst28418 (SUB_1605_U217, SUB_1605_U183);
  nand ginst28419 (SUB_1605_U218, P2_DATAO_REG_12__SCAN_IN, SUB_1605_U33);
  nand ginst28420 (SUB_1605_U219, P1_DATAO_REG_12__SCAN_IN, SUB_1605_U34);
  not ginst28421 (SUB_1605_U22, P1_DATAO_REG_4__SCAN_IN);
  not ginst28422 (SUB_1605_U220, SUB_1605_U182);
  nand ginst28423 (SUB_1605_U221, P2_DATAO_REG_13__SCAN_IN, SUB_1605_U41);
  nand ginst28424 (SUB_1605_U222, SUB_1605_U182, SUB_1605_U221);
  nand ginst28425 (SUB_1605_U223, P1_DATAO_REG_13__SCAN_IN, SUB_1605_U40);
  not ginst28426 (SUB_1605_U224, SUB_1605_U181);
  nand ginst28427 (SUB_1605_U225, P2_DATAO_REG_14__SCAN_IN, SUB_1605_U43);
  nand ginst28428 (SUB_1605_U226, SUB_1605_U181, SUB_1605_U225);
  nand ginst28429 (SUB_1605_U227, P1_DATAO_REG_14__SCAN_IN, SUB_1605_U42);
  not ginst28430 (SUB_1605_U228, SUB_1605_U180);
  nand ginst28431 (SUB_1605_U229, P2_DATAO_REG_15__SCAN_IN, SUB_1605_U45);
  not ginst28432 (SUB_1605_U23, P2_DATAO_REG_0__SCAN_IN);
  nand ginst28433 (SUB_1605_U230, SUB_1605_U180, SUB_1605_U229);
  nand ginst28434 (SUB_1605_U231, P1_DATAO_REG_15__SCAN_IN, SUB_1605_U44);
  not ginst28435 (SUB_1605_U232, SUB_1605_U179);
  nand ginst28436 (SUB_1605_U233, P2_DATAO_REG_16__SCAN_IN, SUB_1605_U47);
  nand ginst28437 (SUB_1605_U234, SUB_1605_U179, SUB_1605_U233);
  nand ginst28438 (SUB_1605_U235, P1_DATAO_REG_16__SCAN_IN, SUB_1605_U46);
  not ginst28439 (SUB_1605_U236, SUB_1605_U178);
  nand ginst28440 (SUB_1605_U237, P2_DATAO_REG_17__SCAN_IN, SUB_1605_U49);
  nand ginst28441 (SUB_1605_U238, SUB_1605_U178, SUB_1605_U237);
  nand ginst28442 (SUB_1605_U239, P1_DATAO_REG_17__SCAN_IN, SUB_1605_U48);
  not ginst28443 (SUB_1605_U24, P1_DATAO_REG_1__SCAN_IN);
  not ginst28444 (SUB_1605_U240, SUB_1605_U177);
  nand ginst28445 (SUB_1605_U241, P2_DATAO_REG_18__SCAN_IN, SUB_1605_U51);
  nand ginst28446 (SUB_1605_U242, SUB_1605_U177, SUB_1605_U241);
  nand ginst28447 (SUB_1605_U243, P1_DATAO_REG_18__SCAN_IN, SUB_1605_U50);
  not ginst28448 (SUB_1605_U244, SUB_1605_U176);
  nand ginst28449 (SUB_1605_U245, P2_DATAO_REG_19__SCAN_IN, SUB_1605_U53);
  nand ginst28450 (SUB_1605_U246, SUB_1605_U176, SUB_1605_U245);
  nand ginst28451 (SUB_1605_U247, P1_DATAO_REG_19__SCAN_IN, SUB_1605_U52);
  not ginst28452 (SUB_1605_U248, SUB_1605_U173);
  nand ginst28453 (SUB_1605_U249, P2_DATAO_REG_20__SCAN_IN, SUB_1605_U55);
  not ginst28454 (SUB_1605_U25, P2_DATAO_REG_4__SCAN_IN);
  nand ginst28455 (SUB_1605_U250, SUB_1605_U173, SUB_1605_U249);
  nand ginst28456 (SUB_1605_U251, P1_DATAO_REG_20__SCAN_IN, SUB_1605_U54);
  not ginst28457 (SUB_1605_U252, SUB_1605_U172);
  nand ginst28458 (SUB_1605_U253, P2_DATAO_REG_21__SCAN_IN, SUB_1605_U57);
  nand ginst28459 (SUB_1605_U254, SUB_1605_U172, SUB_1605_U253);
  nand ginst28460 (SUB_1605_U255, P1_DATAO_REG_21__SCAN_IN, SUB_1605_U56);
  not ginst28461 (SUB_1605_U256, SUB_1605_U171);
  nand ginst28462 (SUB_1605_U257, P2_DATAO_REG_22__SCAN_IN, SUB_1605_U59);
  nand ginst28463 (SUB_1605_U258, SUB_1605_U171, SUB_1605_U257);
  nand ginst28464 (SUB_1605_U259, P1_DATAO_REG_22__SCAN_IN, SUB_1605_U58);
  not ginst28465 (SUB_1605_U26, P2_DATAO_REG_2__SCAN_IN);
  not ginst28466 (SUB_1605_U260, SUB_1605_U170);
  nand ginst28467 (SUB_1605_U261, P2_DATAO_REG_23__SCAN_IN, SUB_1605_U61);
  nand ginst28468 (SUB_1605_U262, SUB_1605_U170, SUB_1605_U261);
  nand ginst28469 (SUB_1605_U263, P1_DATAO_REG_23__SCAN_IN, SUB_1605_U60);
  not ginst28470 (SUB_1605_U264, SUB_1605_U169);
  nand ginst28471 (SUB_1605_U265, P2_DATAO_REG_24__SCAN_IN, SUB_1605_U63);
  nand ginst28472 (SUB_1605_U266, SUB_1605_U169, SUB_1605_U265);
  nand ginst28473 (SUB_1605_U267, P1_DATAO_REG_24__SCAN_IN, SUB_1605_U62);
  not ginst28474 (SUB_1605_U268, SUB_1605_U168);
  nand ginst28475 (SUB_1605_U269, P2_DATAO_REG_25__SCAN_IN, SUB_1605_U65);
  not ginst28476 (SUB_1605_U27, P2_DATAO_REG_3__SCAN_IN);
  nand ginst28477 (SUB_1605_U270, SUB_1605_U168, SUB_1605_U269);
  nand ginst28478 (SUB_1605_U271, P1_DATAO_REG_25__SCAN_IN, SUB_1605_U64);
  not ginst28479 (SUB_1605_U272, SUB_1605_U167);
  nand ginst28480 (SUB_1605_U273, P2_DATAO_REG_26__SCAN_IN, SUB_1605_U67);
  nand ginst28481 (SUB_1605_U274, SUB_1605_U167, SUB_1605_U273);
  nand ginst28482 (SUB_1605_U275, P1_DATAO_REG_26__SCAN_IN, SUB_1605_U66);
  not ginst28483 (SUB_1605_U276, SUB_1605_U166);
  nand ginst28484 (SUB_1605_U277, P2_DATAO_REG_27__SCAN_IN, SUB_1605_U69);
  nand ginst28485 (SUB_1605_U278, SUB_1605_U166, SUB_1605_U277);
  nand ginst28486 (SUB_1605_U279, P1_DATAO_REG_27__SCAN_IN, SUB_1605_U68);
  not ginst28487 (SUB_1605_U28, P1_DATAO_REG_2__SCAN_IN);
  not ginst28488 (SUB_1605_U280, SUB_1605_U165);
  nand ginst28489 (SUB_1605_U281, P2_DATAO_REG_28__SCAN_IN, SUB_1605_U71);
  nand ginst28490 (SUB_1605_U282, SUB_1605_U165, SUB_1605_U281);
  nand ginst28491 (SUB_1605_U283, P1_DATAO_REG_28__SCAN_IN, SUB_1605_U70);
  not ginst28492 (SUB_1605_U284, SUB_1605_U164);
  nand ginst28493 (SUB_1605_U285, P2_DATAO_REG_29__SCAN_IN, SUB_1605_U73);
  nand ginst28494 (SUB_1605_U286, SUB_1605_U164, SUB_1605_U285);
  nand ginst28495 (SUB_1605_U287, P1_DATAO_REG_29__SCAN_IN, SUB_1605_U72);
  not ginst28496 (SUB_1605_U288, SUB_1605_U162);
  nand ginst28497 (SUB_1605_U289, P2_DATAO_REG_30__SCAN_IN, SUB_1605_U74);
  not ginst28498 (SUB_1605_U29, P1_DATAO_REG_3__SCAN_IN);
  nand ginst28499 (SUB_1605_U290, P1_DATAO_REG_30__SCAN_IN, SUB_1605_U75);
  nand ginst28500 (SUB_1605_U291, P1_DATAO_REG_0__SCAN_IN, SUB_1605_U23);
  nand ginst28501 (SUB_1605_U292, P1_DATAO_REG_1__SCAN_IN, SUB_1605_U174);
  nand ginst28502 (SUB_1605_U293, SUB_1605_U126, SUB_1605_U286);
  nand ginst28503 (SUB_1605_U294, SUB_1605_U163, SUB_1605_U6);
  nand ginst28504 (SUB_1605_U295, SUB_1605_U192, SUB_1605_U195);
  nand ginst28505 (SUB_1605_U296, SUB_1605_U295, SUB_1605_U299);
  nand ginst28506 (SUB_1605_U297, SUB_1605_U111, SUB_1605_U163);
  nand ginst28507 (SUB_1605_U298, SUB_1605_U112, SUB_1605_U295);
  nand ginst28508 (SUB_1605_U299, P2_DATAO_REG_3__SCAN_IN, SUB_1605_U29);
  not ginst28509 (SUB_1605_U30, P2_DATAO_REG_5__SCAN_IN);
  nand ginst28510 (SUB_1605_U300, SUB_1605_U109, SUB_1605_U202);
  not ginst28511 (SUB_1605_U301, SUB_1605_U21);
  nand ginst28512 (SUB_1605_U302, SUB_1605_U206, SUB_1605_U301);
  nand ginst28513 (SUB_1605_U303, SUB_1605_U110, SUB_1605_U300);
  nand ginst28514 (SUB_1605_U304, SUB_1605_U152, SUB_1605_U9);
  nand ginst28515 (SUB_1605_U305, SUB_1605_U210, SUB_1605_U212);
  not ginst28516 (SUB_1605_U306, SUB_1605_U77);
  nand ginst28517 (SUB_1605_U307, SUB_1605_U10, SUB_1605_U152);
  nand ginst28518 (SUB_1605_U308, SUB_1605_U215, SUB_1605_U77);
  not ginst28519 (SUB_1605_U309, SUB_1605_U76);
  not ginst28520 (SUB_1605_U31, P2_DATAO_REG_9__SCAN_IN);
  nand ginst28521 (SUB_1605_U310, SUB_1605_U124, SUB_1605_U152);
  nand ginst28522 (SUB_1605_U311, SUB_1605_U218, SUB_1605_U76);
  nand ginst28523 (SUB_1605_U312, SUB_1605_U292, SUB_1605_U313, SUB_1605_U314);
  nand ginst28524 (SUB_1605_U313, P1_DATAO_REG_1__SCAN_IN, SUB_1605_U175);
  nand ginst28525 (SUB_1605_U314, SUB_1605_U174, SUB_1605_U175);
  nand ginst28526 (SUB_1605_U315, SUB_1605_U156, SUB_1605_U200);
  not ginst28527 (SUB_1605_U316, SUB_1605_U155);
  nand ginst28528 (SUB_1605_U317, SUB_1605_U156, SUB_1605_U7);
  not ginst28529 (SUB_1605_U318, SUB_1605_U154);
  nand ginst28530 (SUB_1605_U319, SUB_1605_U156, SUB_1605_U8);
  not ginst28531 (SUB_1605_U32, P1_DATAO_REG_9__SCAN_IN);
  not ginst28532 (SUB_1605_U320, SUB_1605_U153);
  nand ginst28533 (SUB_1605_U321, SUB_1605_U114, SUB_1605_U156);
  not ginst28534 (SUB_1605_U322, SUB_1605_U152);
  nand ginst28535 (SUB_1605_U323, SUB_1605_U127, SUB_1605_U162);
  nand ginst28536 (SUB_1605_U324, P2_DATAO_REG_9__SCAN_IN, SUB_1605_U32);
  nand ginst28537 (SUB_1605_U325, P1_DATAO_REG_9__SCAN_IN, SUB_1605_U31);
  not ginst28538 (SUB_1605_U326, SUB_1605_U116);
  nand ginst28539 (SUB_1605_U327, SUB_1605_U322, SUB_1605_U326);
  nand ginst28540 (SUB_1605_U328, SUB_1605_U116, SUB_1605_U152);
  nand ginst28541 (SUB_1605_U329, P2_DATAO_REG_8__SCAN_IN, SUB_1605_U14);
  not ginst28542 (SUB_1605_U33, P1_DATAO_REG_12__SCAN_IN);
  nand ginst28543 (SUB_1605_U330, P1_DATAO_REG_8__SCAN_IN, SUB_1605_U15);
  not ginst28544 (SUB_1605_U331, SUB_1605_U117);
  nand ginst28545 (SUB_1605_U332, SUB_1605_U320, SUB_1605_U331);
  nand ginst28546 (SUB_1605_U333, SUB_1605_U117, SUB_1605_U153);
  nand ginst28547 (SUB_1605_U334, P2_DATAO_REG_7__SCAN_IN, SUB_1605_U18);
  nand ginst28548 (SUB_1605_U335, P1_DATAO_REG_7__SCAN_IN, SUB_1605_U16);
  not ginst28549 (SUB_1605_U336, SUB_1605_U119);
  nand ginst28550 (SUB_1605_U337, SUB_1605_U318, SUB_1605_U336);
  nand ginst28551 (SUB_1605_U338, SUB_1605_U119, SUB_1605_U154);
  nand ginst28552 (SUB_1605_U339, P2_DATAO_REG_6__SCAN_IN, SUB_1605_U17);
  not ginst28553 (SUB_1605_U34, P2_DATAO_REG_12__SCAN_IN);
  nand ginst28554 (SUB_1605_U340, P1_DATAO_REG_6__SCAN_IN, SUB_1605_U19);
  not ginst28555 (SUB_1605_U341, SUB_1605_U120);
  nand ginst28556 (SUB_1605_U342, SUB_1605_U316, SUB_1605_U341);
  nand ginst28557 (SUB_1605_U343, SUB_1605_U120, SUB_1605_U155);
  nand ginst28558 (SUB_1605_U344, P2_DATAO_REG_5__SCAN_IN, SUB_1605_U20);
  nand ginst28559 (SUB_1605_U345, P1_DATAO_REG_5__SCAN_IN, SUB_1605_U30);
  not ginst28560 (SUB_1605_U346, SUB_1605_U121);
  nand ginst28561 (SUB_1605_U347, SUB_1605_U199, SUB_1605_U346);
  nand ginst28562 (SUB_1605_U348, SUB_1605_U121, SUB_1605_U156);
  nand ginst28563 (SUB_1605_U349, P2_DATAO_REG_4__SCAN_IN, SUB_1605_U22);
  not ginst28564 (SUB_1605_U35, P2_DATAO_REG_11__SCAN_IN);
  nand ginst28565 (SUB_1605_U350, P1_DATAO_REG_4__SCAN_IN, SUB_1605_U25);
  not ginst28566 (SUB_1605_U351, SUB_1605_U122);
  nand ginst28567 (SUB_1605_U352, SUB_1605_U196, SUB_1605_U351);
  nand ginst28568 (SUB_1605_U353, SUB_1605_U122, SUB_1605_U157);
  nand ginst28569 (SUB_1605_U354, P2_DATAO_REG_3__SCAN_IN, SUB_1605_U29);
  nand ginst28570 (SUB_1605_U355, P1_DATAO_REG_3__SCAN_IN, SUB_1605_U27);
  not ginst28571 (SUB_1605_U356, SUB_1605_U123);
  nand ginst28572 (SUB_1605_U357, SUB_1605_U193, SUB_1605_U356);
  nand ginst28573 (SUB_1605_U358, SUB_1605_U123, SUB_1605_U158);
  nand ginst28574 (SUB_1605_U359, P2_DATAO_REG_31__SCAN_IN, SUB_1605_U160);
  not ginst28575 (SUB_1605_U36, P2_DATAO_REG_10__SCAN_IN);
  nand ginst28576 (SUB_1605_U360, P1_DATAO_REG_31__SCAN_IN, SUB_1605_U159);
  nand ginst28577 (SUB_1605_U361, SUB_1605_U359, SUB_1605_U360);
  nand ginst28578 (SUB_1605_U362, P2_DATAO_REG_31__SCAN_IN, SUB_1605_U160);
  nand ginst28579 (SUB_1605_U363, P1_DATAO_REG_31__SCAN_IN, SUB_1605_U159);
  nand ginst28580 (SUB_1605_U364, P1_DATAO_REG_30__SCAN_IN, SUB_1605_U361, SUB_1605_U75);
  nand ginst28581 (SUB_1605_U365, P2_DATAO_REG_30__SCAN_IN, SUB_1605_U11, SUB_1605_U74);
  nand ginst28582 (SUB_1605_U366, P2_DATAO_REG_30__SCAN_IN, SUB_1605_U74);
  nand ginst28583 (SUB_1605_U367, P1_DATAO_REG_30__SCAN_IN, SUB_1605_U75);
  not ginst28584 (SUB_1605_U368, SUB_1605_U129);
  nand ginst28585 (SUB_1605_U369, SUB_1605_U288, SUB_1605_U368);
  not ginst28586 (SUB_1605_U37, P1_DATAO_REG_11__SCAN_IN);
  nand ginst28587 (SUB_1605_U370, SUB_1605_U129, SUB_1605_U162);
  nand ginst28588 (SUB_1605_U371, P2_DATAO_REG_2__SCAN_IN, SUB_1605_U28);
  nand ginst28589 (SUB_1605_U372, P1_DATAO_REG_2__SCAN_IN, SUB_1605_U26);
  not ginst28590 (SUB_1605_U373, SUB_1605_U130);
  nand ginst28591 (SUB_1605_U374, SUB_1605_U189, SUB_1605_U373);
  nand ginst28592 (SUB_1605_U375, SUB_1605_U130, SUB_1605_U163);
  nand ginst28593 (SUB_1605_U376, P2_DATAO_REG_29__SCAN_IN, SUB_1605_U73);
  nand ginst28594 (SUB_1605_U377, P1_DATAO_REG_29__SCAN_IN, SUB_1605_U72);
  not ginst28595 (SUB_1605_U378, SUB_1605_U131);
  nand ginst28596 (SUB_1605_U379, SUB_1605_U284, SUB_1605_U378);
  not ginst28597 (SUB_1605_U38, P1_DATAO_REG_10__SCAN_IN);
  nand ginst28598 (SUB_1605_U380, SUB_1605_U131, SUB_1605_U164);
  nand ginst28599 (SUB_1605_U381, P2_DATAO_REG_28__SCAN_IN, SUB_1605_U71);
  nand ginst28600 (SUB_1605_U382, P1_DATAO_REG_28__SCAN_IN, SUB_1605_U70);
  not ginst28601 (SUB_1605_U383, SUB_1605_U132);
  nand ginst28602 (SUB_1605_U384, SUB_1605_U280, SUB_1605_U383);
  nand ginst28603 (SUB_1605_U385, SUB_1605_U132, SUB_1605_U165);
  nand ginst28604 (SUB_1605_U386, P2_DATAO_REG_27__SCAN_IN, SUB_1605_U69);
  nand ginst28605 (SUB_1605_U387, P1_DATAO_REG_27__SCAN_IN, SUB_1605_U68);
  not ginst28606 (SUB_1605_U388, SUB_1605_U133);
  nand ginst28607 (SUB_1605_U389, SUB_1605_U276, SUB_1605_U388);
  nand ginst28608 (SUB_1605_U39, P1_DATAO_REG_9__SCAN_IN, SUB_1605_U31);
  nand ginst28609 (SUB_1605_U390, SUB_1605_U133, SUB_1605_U166);
  nand ginst28610 (SUB_1605_U391, P2_DATAO_REG_26__SCAN_IN, SUB_1605_U67);
  nand ginst28611 (SUB_1605_U392, P1_DATAO_REG_26__SCAN_IN, SUB_1605_U66);
  not ginst28612 (SUB_1605_U393, SUB_1605_U134);
  nand ginst28613 (SUB_1605_U394, SUB_1605_U272, SUB_1605_U393);
  nand ginst28614 (SUB_1605_U395, SUB_1605_U134, SUB_1605_U167);
  nand ginst28615 (SUB_1605_U396, P2_DATAO_REG_25__SCAN_IN, SUB_1605_U65);
  nand ginst28616 (SUB_1605_U397, P1_DATAO_REG_25__SCAN_IN, SUB_1605_U64);
  not ginst28617 (SUB_1605_U398, SUB_1605_U135);
  nand ginst28618 (SUB_1605_U399, SUB_1605_U268, SUB_1605_U398);
  not ginst28619 (SUB_1605_U40, P2_DATAO_REG_13__SCAN_IN);
  nand ginst28620 (SUB_1605_U400, SUB_1605_U135, SUB_1605_U168);
  nand ginst28621 (SUB_1605_U401, P2_DATAO_REG_24__SCAN_IN, SUB_1605_U63);
  nand ginst28622 (SUB_1605_U402, P1_DATAO_REG_24__SCAN_IN, SUB_1605_U62);
  not ginst28623 (SUB_1605_U403, SUB_1605_U136);
  nand ginst28624 (SUB_1605_U404, SUB_1605_U264, SUB_1605_U403);
  nand ginst28625 (SUB_1605_U405, SUB_1605_U136, SUB_1605_U169);
  nand ginst28626 (SUB_1605_U406, P2_DATAO_REG_23__SCAN_IN, SUB_1605_U61);
  nand ginst28627 (SUB_1605_U407, P1_DATAO_REG_23__SCAN_IN, SUB_1605_U60);
  not ginst28628 (SUB_1605_U408, SUB_1605_U137);
  nand ginst28629 (SUB_1605_U409, SUB_1605_U260, SUB_1605_U408);
  not ginst28630 (SUB_1605_U41, P1_DATAO_REG_13__SCAN_IN);
  nand ginst28631 (SUB_1605_U410, SUB_1605_U137, SUB_1605_U170);
  nand ginst28632 (SUB_1605_U411, P2_DATAO_REG_22__SCAN_IN, SUB_1605_U59);
  nand ginst28633 (SUB_1605_U412, P1_DATAO_REG_22__SCAN_IN, SUB_1605_U58);
  not ginst28634 (SUB_1605_U413, SUB_1605_U138);
  nand ginst28635 (SUB_1605_U414, SUB_1605_U256, SUB_1605_U413);
  nand ginst28636 (SUB_1605_U415, SUB_1605_U138, SUB_1605_U171);
  nand ginst28637 (SUB_1605_U416, P2_DATAO_REG_21__SCAN_IN, SUB_1605_U57);
  nand ginst28638 (SUB_1605_U417, P1_DATAO_REG_21__SCAN_IN, SUB_1605_U56);
  not ginst28639 (SUB_1605_U418, SUB_1605_U139);
  nand ginst28640 (SUB_1605_U419, SUB_1605_U252, SUB_1605_U418);
  not ginst28641 (SUB_1605_U42, P2_DATAO_REG_14__SCAN_IN);
  nand ginst28642 (SUB_1605_U420, SUB_1605_U139, SUB_1605_U172);
  nand ginst28643 (SUB_1605_U421, P2_DATAO_REG_20__SCAN_IN, SUB_1605_U55);
  nand ginst28644 (SUB_1605_U422, P1_DATAO_REG_20__SCAN_IN, SUB_1605_U54);
  not ginst28645 (SUB_1605_U423, SUB_1605_U140);
  nand ginst28646 (SUB_1605_U424, SUB_1605_U248, SUB_1605_U423);
  nand ginst28647 (SUB_1605_U425, SUB_1605_U140, SUB_1605_U173);
  nand ginst28648 (SUB_1605_U426, P2_DATAO_REG_1__SCAN_IN, SUB_1605_U24);
  nand ginst28649 (SUB_1605_U427, P1_DATAO_REG_1__SCAN_IN, SUB_1605_U174);
  not ginst28650 (SUB_1605_U428, SUB_1605_U141);
  nand ginst28651 (SUB_1605_U429, SUB_1605_U187, SUB_1605_U428);
  not ginst28652 (SUB_1605_U43, P1_DATAO_REG_14__SCAN_IN);
  nand ginst28653 (SUB_1605_U430, SUB_1605_U141, SUB_1605_U175);
  nand ginst28654 (SUB_1605_U431, P2_DATAO_REG_19__SCAN_IN, SUB_1605_U53);
  nand ginst28655 (SUB_1605_U432, P1_DATAO_REG_19__SCAN_IN, SUB_1605_U52);
  not ginst28656 (SUB_1605_U433, SUB_1605_U142);
  nand ginst28657 (SUB_1605_U434, SUB_1605_U244, SUB_1605_U433);
  nand ginst28658 (SUB_1605_U435, SUB_1605_U142, SUB_1605_U176);
  nand ginst28659 (SUB_1605_U436, P2_DATAO_REG_18__SCAN_IN, SUB_1605_U51);
  nand ginst28660 (SUB_1605_U437, P1_DATAO_REG_18__SCAN_IN, SUB_1605_U50);
  not ginst28661 (SUB_1605_U438, SUB_1605_U143);
  nand ginst28662 (SUB_1605_U439, SUB_1605_U240, SUB_1605_U438);
  not ginst28663 (SUB_1605_U44, P2_DATAO_REG_15__SCAN_IN);
  nand ginst28664 (SUB_1605_U440, SUB_1605_U143, SUB_1605_U177);
  nand ginst28665 (SUB_1605_U441, P2_DATAO_REG_17__SCAN_IN, SUB_1605_U49);
  nand ginst28666 (SUB_1605_U442, P1_DATAO_REG_17__SCAN_IN, SUB_1605_U48);
  not ginst28667 (SUB_1605_U443, SUB_1605_U144);
  nand ginst28668 (SUB_1605_U444, SUB_1605_U236, SUB_1605_U443);
  nand ginst28669 (SUB_1605_U445, SUB_1605_U144, SUB_1605_U178);
  nand ginst28670 (SUB_1605_U446, P2_DATAO_REG_16__SCAN_IN, SUB_1605_U47);
  nand ginst28671 (SUB_1605_U447, P1_DATAO_REG_16__SCAN_IN, SUB_1605_U46);
  not ginst28672 (SUB_1605_U448, SUB_1605_U145);
  nand ginst28673 (SUB_1605_U449, SUB_1605_U232, SUB_1605_U448);
  not ginst28674 (SUB_1605_U45, P1_DATAO_REG_15__SCAN_IN);
  nand ginst28675 (SUB_1605_U450, SUB_1605_U145, SUB_1605_U179);
  nand ginst28676 (SUB_1605_U451, P2_DATAO_REG_15__SCAN_IN, SUB_1605_U45);
  nand ginst28677 (SUB_1605_U452, P1_DATAO_REG_15__SCAN_IN, SUB_1605_U44);
  not ginst28678 (SUB_1605_U453, SUB_1605_U146);
  nand ginst28679 (SUB_1605_U454, SUB_1605_U228, SUB_1605_U453);
  nand ginst28680 (SUB_1605_U455, SUB_1605_U146, SUB_1605_U180);
  nand ginst28681 (SUB_1605_U456, P2_DATAO_REG_14__SCAN_IN, SUB_1605_U43);
  nand ginst28682 (SUB_1605_U457, P1_DATAO_REG_14__SCAN_IN, SUB_1605_U42);
  not ginst28683 (SUB_1605_U458, SUB_1605_U147);
  nand ginst28684 (SUB_1605_U459, SUB_1605_U224, SUB_1605_U458);
  not ginst28685 (SUB_1605_U46, P2_DATAO_REG_16__SCAN_IN);
  nand ginst28686 (SUB_1605_U460, SUB_1605_U147, SUB_1605_U181);
  nand ginst28687 (SUB_1605_U461, P2_DATAO_REG_13__SCAN_IN, SUB_1605_U41);
  nand ginst28688 (SUB_1605_U462, P1_DATAO_REG_13__SCAN_IN, SUB_1605_U40);
  not ginst28689 (SUB_1605_U463, SUB_1605_U148);
  nand ginst28690 (SUB_1605_U464, SUB_1605_U220, SUB_1605_U463);
  nand ginst28691 (SUB_1605_U465, SUB_1605_U148, SUB_1605_U182);
  nand ginst28692 (SUB_1605_U466, P2_DATAO_REG_12__SCAN_IN, SUB_1605_U33);
  nand ginst28693 (SUB_1605_U467, P1_DATAO_REG_12__SCAN_IN, SUB_1605_U34);
  not ginst28694 (SUB_1605_U468, SUB_1605_U149);
  nand ginst28695 (SUB_1605_U469, SUB_1605_U217, SUB_1605_U468);
  not ginst28696 (SUB_1605_U47, P1_DATAO_REG_16__SCAN_IN);
  nand ginst28697 (SUB_1605_U470, SUB_1605_U149, SUB_1605_U183);
  nand ginst28698 (SUB_1605_U471, P2_DATAO_REG_11__SCAN_IN, SUB_1605_U37);
  nand ginst28699 (SUB_1605_U472, P1_DATAO_REG_11__SCAN_IN, SUB_1605_U35);
  not ginst28700 (SUB_1605_U473, SUB_1605_U150);
  nand ginst28701 (SUB_1605_U474, SUB_1605_U214, SUB_1605_U473);
  nand ginst28702 (SUB_1605_U475, SUB_1605_U150, SUB_1605_U184);
  nand ginst28703 (SUB_1605_U476, P2_DATAO_REG_10__SCAN_IN, SUB_1605_U38);
  nand ginst28704 (SUB_1605_U477, P1_DATAO_REG_10__SCAN_IN, SUB_1605_U36);
  not ginst28705 (SUB_1605_U478, SUB_1605_U151);
  nand ginst28706 (SUB_1605_U479, SUB_1605_U211, SUB_1605_U478);
  not ginst28707 (SUB_1605_U48, P2_DATAO_REG_17__SCAN_IN);
  nand ginst28708 (SUB_1605_U480, SUB_1605_U151, SUB_1605_U185);
  not ginst28709 (SUB_1605_U49, P1_DATAO_REG_17__SCAN_IN);
  not ginst28710 (SUB_1605_U50, P2_DATAO_REG_18__SCAN_IN);
  not ginst28711 (SUB_1605_U51, P1_DATAO_REG_18__SCAN_IN);
  not ginst28712 (SUB_1605_U52, P2_DATAO_REG_19__SCAN_IN);
  not ginst28713 (SUB_1605_U53, P1_DATAO_REG_19__SCAN_IN);
  not ginst28714 (SUB_1605_U54, P2_DATAO_REG_20__SCAN_IN);
  not ginst28715 (SUB_1605_U55, P1_DATAO_REG_20__SCAN_IN);
  not ginst28716 (SUB_1605_U56, P2_DATAO_REG_21__SCAN_IN);
  not ginst28717 (SUB_1605_U57, P1_DATAO_REG_21__SCAN_IN);
  not ginst28718 (SUB_1605_U58, P2_DATAO_REG_22__SCAN_IN);
  not ginst28719 (SUB_1605_U59, P1_DATAO_REG_22__SCAN_IN);
  and ginst28720 (SUB_1605_U6, SUB_1605_U190, SUB_1605_U194);
  not ginst28721 (SUB_1605_U60, P2_DATAO_REG_23__SCAN_IN);
  not ginst28722 (SUB_1605_U61, P1_DATAO_REG_23__SCAN_IN);
  not ginst28723 (SUB_1605_U62, P2_DATAO_REG_24__SCAN_IN);
  not ginst28724 (SUB_1605_U63, P1_DATAO_REG_24__SCAN_IN);
  not ginst28725 (SUB_1605_U64, P2_DATAO_REG_25__SCAN_IN);
  not ginst28726 (SUB_1605_U65, P1_DATAO_REG_25__SCAN_IN);
  not ginst28727 (SUB_1605_U66, P2_DATAO_REG_26__SCAN_IN);
  not ginst28728 (SUB_1605_U67, P1_DATAO_REG_26__SCAN_IN);
  not ginst28729 (SUB_1605_U68, P2_DATAO_REG_27__SCAN_IN);
  not ginst28730 (SUB_1605_U69, P1_DATAO_REG_27__SCAN_IN);
  and ginst28731 (SUB_1605_U7, SUB_1605_U200, SUB_1605_U202);
  not ginst28732 (SUB_1605_U70, P2_DATAO_REG_28__SCAN_IN);
  not ginst28733 (SUB_1605_U71, P1_DATAO_REG_28__SCAN_IN);
  not ginst28734 (SUB_1605_U72, P2_DATAO_REG_29__SCAN_IN);
  not ginst28735 (SUB_1605_U73, P1_DATAO_REG_29__SCAN_IN);
  not ginst28736 (SUB_1605_U74, P1_DATAO_REG_30__SCAN_IN);
  not ginst28737 (SUB_1605_U75, P2_DATAO_REG_30__SCAN_IN);
  nand ginst28738 (SUB_1605_U76, SUB_1605_U216, SUB_1605_U308);
  nand ginst28739 (SUB_1605_U77, SUB_1605_U213, SUB_1605_U305);
  not ginst28740 (SUB_1605_U78, P1_DATAO_REG_0__SCAN_IN);
  nand ginst28741 (SUB_1605_U79, SUB_1605_U327, SUB_1605_U328);
  and ginst28742 (SUB_1605_U8, SUB_1605_U204, SUB_1605_U7);
  nand ginst28743 (SUB_1605_U80, SUB_1605_U332, SUB_1605_U333);
  nand ginst28744 (SUB_1605_U81, SUB_1605_U337, SUB_1605_U338);
  nand ginst28745 (SUB_1605_U82, SUB_1605_U342, SUB_1605_U343);
  nand ginst28746 (SUB_1605_U83, SUB_1605_U347, SUB_1605_U348);
  nand ginst28747 (SUB_1605_U84, SUB_1605_U352, SUB_1605_U353);
  nand ginst28748 (SUB_1605_U85, SUB_1605_U357, SUB_1605_U358);
  nand ginst28749 (SUB_1605_U86, SUB_1605_U369, SUB_1605_U370);
  nand ginst28750 (SUB_1605_U87, SUB_1605_U374, SUB_1605_U375);
  nand ginst28751 (SUB_1605_U88, SUB_1605_U379, SUB_1605_U380);
  nand ginst28752 (SUB_1605_U89, SUB_1605_U384, SUB_1605_U385);
  and ginst28753 (SUB_1605_U9, SUB_1605_U208, SUB_1605_U212);
  nand ginst28754 (SUB_1605_U90, SUB_1605_U389, SUB_1605_U390);
  nand ginst28755 (SUB_1605_U91, SUB_1605_U394, SUB_1605_U395);
  nand ginst28756 (SUB_1605_U92, SUB_1605_U399, SUB_1605_U400);
  nand ginst28757 (SUB_1605_U93, SUB_1605_U404, SUB_1605_U405);
  nand ginst28758 (SUB_1605_U94, SUB_1605_U409, SUB_1605_U410);
  nand ginst28759 (SUB_1605_U95, SUB_1605_U414, SUB_1605_U415);
  nand ginst28760 (SUB_1605_U96, SUB_1605_U419, SUB_1605_U420);
  nand ginst28761 (SUB_1605_U97, SUB_1605_U424, SUB_1605_U425);
  nand ginst28762 (SUB_1605_U98, SUB_1605_U429, SUB_1605_U430);
  nand ginst28763 (SUB_1605_U99, SUB_1605_U434, SUB_1605_U435);
  nand ginst28764 (U100, U312, U313);
  nand ginst28765 (U101, U314, U315);
  nand ginst28766 (U102, U316, U317);
  nand ginst28767 (U103, U318, U319);
  nand ginst28768 (U104, U320, U321);
  nand ginst28769 (U105, U322, U323);
  nand ginst28770 (U106, U324, U325);
  nand ginst28771 (U107, U326, U327);
  nand ginst28772 (U108, U328, U329);
  nand ginst28773 (U109, U330, U331);
  nand ginst28774 (U110, U332, U333);
  nand ginst28775 (U111, U334, U335);
  nand ginst28776 (U112, U336, U337);
  nand ginst28777 (U113, U338, U339);
  nand ginst28778 (U114, U340, U341);
  nand ginst28779 (U115, U342, U343);
  nand ginst28780 (U116, U344, U345);
  nand ginst28781 (U117, U346, U347);
  nand ginst28782 (U118, U348, U349);
  nand ginst28783 (U119, U350, U351);
  nand ginst28784 (U120, U352, U353);
  nand ginst28785 (U121, U354, U355);
  nand ginst28786 (U122, U356, U357);
  nand ginst28787 (U123, U358, U359);
  nand ginst28788 (U124, U360, U361);
  nand ginst28789 (U125, U362, U363);
  nand ginst28790 (U126, U364, U365);
  nand ginst28791 (U127, U366, U367);
  nand ginst28792 (U128, U368, U369);
  nand ginst28793 (U129, U370, U371);
  nand ginst28794 (U130, U372, U373);
  nand ginst28795 (U131, U374, U375);
  nand ginst28796 (U132, U376, U377);
  nand ginst28797 (U133, U378, U379);
  nand ginst28798 (U134, U380, U381);
  nand ginst28799 (U135, U382, U383);
  nand ginst28800 (U136, U384, U385);
  nand ginst28801 (U137, U386, U387);
  nand ginst28802 (U138, U388, U389);
  nand ginst28803 (U139, U390, U391);
  nand ginst28804 (U140, U392, U393);
  nand ginst28805 (U141, U394, U395);
  nand ginst28806 (U142, U396, U397);
  nand ginst28807 (U143, U398, U399);
  nand ginst28808 (U144, U400, U401);
  nand ginst28809 (U145, U402, U403);
  nand ginst28810 (U146, U404, U405);
  nand ginst28811 (U147, U406, U407);
  nand ginst28812 (U148, U408, U409);
  nand ginst28813 (U149, U410, U411);
  nand ginst28814 (U150, U412, U413);
  nand ginst28815 (U151, U414, U415);
  nand ginst28816 (U152, U416, U417);
  nand ginst28817 (U153, U418, U419);
  nand ginst28818 (U154, U420, U421);
  nand ginst28819 (U155, U422, U423);
  nand ginst28820 (U156, U424, U425);
  nand ginst28821 (U157, U426, U427);
  not ginst28822 (U158, P2_WR_REG_SCAN_IN);
  not ginst28823 (U159, P1_WR_REG_SCAN_IN);
  and ginst28824 (U160, U168, U169);
  not ginst28825 (U161, P2_RD_REG_SCAN_IN);
  not ginst28826 (U162, P1_RD_REG_SCAN_IN);
  and ginst28827 (U163, U170, U171);
  nand ginst28828 (U164, U165, U166);
  nand ginst28829 (U165, P1_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_19__SCAN_IN, LT_1602_U6, U161);
  nand ginst28830 (U166, P3_ADDR_REG_19__SCAN_IN, LT_1601_21_U6, LT_1601_U6, U162);
  not ginst28831 (U167, U164);
  nand ginst28832 (U168, P2_WR_REG_SCAN_IN, U159);
  nand ginst28833 (U169, P1_WR_REG_SCAN_IN, U158);
  nand ginst28834 (U170, P2_RD_REG_SCAN_IN, U162);
  nand ginst28835 (U171, P1_RD_REG_SCAN_IN, U161);
  nand ginst28836 (U172, SUB_1605_U79, U164);
  nand ginst28837 (U173, SI_9_, U167);
  nand ginst28838 (U174, SUB_1605_U80, U164);
  nand ginst28839 (U175, SI_8_, U167);
  nand ginst28840 (U176, SUB_1605_U81, U164);
  nand ginst28841 (U177, SI_7_, U167);
  nand ginst28842 (U178, SUB_1605_U82, U164);
  nand ginst28843 (U179, SI_6_, U167);
  nand ginst28844 (U180, SUB_1605_U83, U164);
  nand ginst28845 (U181, SI_5_, U167);
  nand ginst28846 (U182, SUB_1605_U84, U164);
  nand ginst28847 (U183, SI_4_, U167);
  nand ginst28848 (U184, SUB_1605_U85, U164);
  nand ginst28849 (U185, SI_3_, U167);
  nand ginst28850 (U186, SUB_1605_U12, U164);
  nand ginst28851 (U187, SI_31_, U167);
  nand ginst28852 (U188, SUB_1605_U86, U164);
  nand ginst28853 (U189, SI_30_, U167);
  nand ginst28854 (U190, SUB_1605_U87, U164);
  nand ginst28855 (U191, SI_2_, U167);
  nand ginst28856 (U192, SUB_1605_U88, U164);
  nand ginst28857 (U193, SI_29_, U167);
  nand ginst28858 (U194, SUB_1605_U89, U164);
  nand ginst28859 (U195, SI_28_, U167);
  nand ginst28860 (U196, SUB_1605_U90, U164);
  nand ginst28861 (U197, SI_27_, U167);
  nand ginst28862 (U198, SUB_1605_U91, U164);
  nand ginst28863 (U199, SI_26_, U167);
  nand ginst28864 (U200, SUB_1605_U92, U164);
  nand ginst28865 (U201, SI_25_, U167);
  nand ginst28866 (U202, SUB_1605_U93, U164);
  nand ginst28867 (U203, SI_24_, U167);
  nand ginst28868 (U204, SUB_1605_U94, U164);
  nand ginst28869 (U205, SI_23_, U167);
  nand ginst28870 (U206, SUB_1605_U95, U164);
  nand ginst28871 (U207, SI_22_, U167);
  nand ginst28872 (U208, SUB_1605_U96, U164);
  nand ginst28873 (U209, SI_21_, U167);
  nand ginst28874 (U210, SUB_1605_U97, U164);
  nand ginst28875 (U211, SI_20_, U167);
  nand ginst28876 (U212, SUB_1605_U98, U164);
  nand ginst28877 (U213, SI_1_, U167);
  nand ginst28878 (U214, SUB_1605_U99, U164);
  nand ginst28879 (U215, SI_19_, U167);
  nand ginst28880 (U216, SUB_1605_U100, U164);
  nand ginst28881 (U217, SI_18_, U167);
  nand ginst28882 (U218, SUB_1605_U101, U164);
  nand ginst28883 (U219, SI_17_, U167);
  nand ginst28884 (U220, SUB_1605_U102, U164);
  nand ginst28885 (U221, SI_16_, U167);
  nand ginst28886 (U222, SUB_1605_U103, U164);
  nand ginst28887 (U223, SI_15_, U167);
  nand ginst28888 (U224, SUB_1605_U104, U164);
  nand ginst28889 (U225, SI_14_, U167);
  nand ginst28890 (U226, SUB_1605_U105, U164);
  nand ginst28891 (U227, SI_13_, U167);
  nand ginst28892 (U228, SUB_1605_U106, U164);
  nand ginst28893 (U229, SI_12_, U167);
  nand ginst28894 (U230, SUB_1605_U107, U164);
  nand ginst28895 (U231, SI_11_, U167);
  nand ginst28896 (U232, SUB_1605_U108, U164);
  nand ginst28897 (U233, SI_10_, U167);
  nand ginst28898 (U234, SUB_1605_U13, U164);
  nand ginst28899 (U235, SI_0_, U167);
  nand ginst28900 (U236, P1_DATAO_REG_9__SCAN_IN, U164);
  nand ginst28901 (U237, R152_U85, U167);
  nand ginst28902 (U238, P1_DATAO_REG_8__SCAN_IN, U164);
  nand ginst28903 (U239, R152_U86, U167);
  nand ginst28904 (U240, P1_DATAO_REG_7__SCAN_IN, U164);
  nand ginst28905 (U241, R152_U87, U167);
  nand ginst28906 (U242, P1_DATAO_REG_6__SCAN_IN, U164);
  nand ginst28907 (U243, R152_U88, U167);
  nand ginst28908 (U244, P1_DATAO_REG_5__SCAN_IN, U164);
  nand ginst28909 (U245, R152_U89, U167);
  nand ginst28910 (U246, P1_DATAO_REG_4__SCAN_IN, U164);
  nand ginst28911 (U247, R152_U90, U167);
  nand ginst28912 (U248, P1_DATAO_REG_3__SCAN_IN, U164);
  nand ginst28913 (U249, R152_U91, U167);
  nand ginst28914 (U250, P1_DATAO_REG_31__SCAN_IN, U164);
  nand ginst28915 (U251, R152_U12, U167);
  nand ginst28916 (U252, P1_DATAO_REG_30__SCAN_IN, U164);
  nand ginst28917 (U253, R152_U92, U167);
  nand ginst28918 (U254, P1_DATAO_REG_2__SCAN_IN, U164);
  nand ginst28919 (U255, R152_U93, U167);
  nand ginst28920 (U256, P1_DATAO_REG_29__SCAN_IN, U164);
  nand ginst28921 (U257, R152_U94, U167);
  nand ginst28922 (U258, P1_DATAO_REG_28__SCAN_IN, U164);
  nand ginst28923 (U259, R152_U95, U167);
  nand ginst28924 (U260, P1_DATAO_REG_27__SCAN_IN, U164);
  nand ginst28925 (U261, R152_U96, U167);
  nand ginst28926 (U262, P1_DATAO_REG_26__SCAN_IN, U164);
  nand ginst28927 (U263, R152_U97, U167);
  nand ginst28928 (U264, P1_DATAO_REG_25__SCAN_IN, U164);
  nand ginst28929 (U265, R152_U98, U167);
  nand ginst28930 (U266, P1_DATAO_REG_24__SCAN_IN, U164);
  nand ginst28931 (U267, R152_U99, U167);
  nand ginst28932 (U268, P1_DATAO_REG_23__SCAN_IN, U164);
  nand ginst28933 (U269, R152_U100, U167);
  nand ginst28934 (U270, P1_DATAO_REG_22__SCAN_IN, U164);
  nand ginst28935 (U271, R152_U101, U167);
  nand ginst28936 (U272, P1_DATAO_REG_21__SCAN_IN, U164);
  nand ginst28937 (U273, R152_U102, U167);
  nand ginst28938 (U274, P1_DATAO_REG_20__SCAN_IN, U164);
  nand ginst28939 (U275, R152_U103, U167);
  nand ginst28940 (U276, P1_DATAO_REG_1__SCAN_IN, U164);
  nand ginst28941 (U277, R152_U13, U167);
  nand ginst28942 (U278, P1_DATAO_REG_19__SCAN_IN, U164);
  nand ginst28943 (U279, R152_U104, U167);
  or ginst28944 (U28, P3_WR_REG_SCAN_IN, U160);
  nand ginst28945 (U280, P1_DATAO_REG_18__SCAN_IN, U164);
  nand ginst28946 (U281, R152_U105, U167);
  nand ginst28947 (U282, P1_DATAO_REG_17__SCAN_IN, U164);
  nand ginst28948 (U283, R152_U106, U167);
  nand ginst28949 (U284, P1_DATAO_REG_16__SCAN_IN, U164);
  nand ginst28950 (U285, R152_U107, U167);
  nand ginst28951 (U286, P1_DATAO_REG_15__SCAN_IN, U164);
  nand ginst28952 (U287, R152_U108, U167);
  nand ginst28953 (U288, P1_DATAO_REG_14__SCAN_IN, U164);
  nand ginst28954 (U289, R152_U109, U167);
  or ginst28955 (U29, P3_RD_REG_SCAN_IN, U163);
  nand ginst28956 (U290, P1_DATAO_REG_13__SCAN_IN, U164);
  nand ginst28957 (U291, R152_U110, U167);
  nand ginst28958 (U292, P1_DATAO_REG_12__SCAN_IN, U164);
  nand ginst28959 (U293, R152_U111, U167);
  nand ginst28960 (U294, P1_DATAO_REG_11__SCAN_IN, U164);
  nand ginst28961 (U295, R152_U112, U167);
  nand ginst28962 (U296, P1_DATAO_REG_10__SCAN_IN, U164);
  nand ginst28963 (U297, R152_U113, U167);
  nand ginst28964 (U298, P1_DATAO_REG_0__SCAN_IN, U164);
  nand ginst28965 (U299, R152_U84, U167);
  nand ginst28966 (U30, U172, U173);
  nand ginst28967 (U300, R152_U85, U164);
  nand ginst28968 (U301, P2_DATAO_REG_9__SCAN_IN, U167);
  nand ginst28969 (U302, R152_U86, U164);
  nand ginst28970 (U303, P2_DATAO_REG_8__SCAN_IN, U167);
  nand ginst28971 (U304, R152_U87, U164);
  nand ginst28972 (U305, P2_DATAO_REG_7__SCAN_IN, U167);
  nand ginst28973 (U306, R152_U88, U164);
  nand ginst28974 (U307, P2_DATAO_REG_6__SCAN_IN, U167);
  nand ginst28975 (U308, R152_U89, U164);
  nand ginst28976 (U309, P2_DATAO_REG_5__SCAN_IN, U167);
  nand ginst28977 (U31, U174, U175);
  nand ginst28978 (U310, R152_U90, U164);
  nand ginst28979 (U311, P2_DATAO_REG_4__SCAN_IN, U167);
  nand ginst28980 (U312, R152_U91, U164);
  nand ginst28981 (U313, P2_DATAO_REG_3__SCAN_IN, U167);
  nand ginst28982 (U314, R152_U12, U164);
  nand ginst28983 (U315, P2_DATAO_REG_31__SCAN_IN, U167);
  nand ginst28984 (U316, R152_U92, U164);
  nand ginst28985 (U317, P2_DATAO_REG_30__SCAN_IN, U167);
  nand ginst28986 (U318, R152_U93, U164);
  nand ginst28987 (U319, P2_DATAO_REG_2__SCAN_IN, U167);
  nand ginst28988 (U32, U176, U177);
  nand ginst28989 (U320, R152_U94, U164);
  nand ginst28990 (U321, P2_DATAO_REG_29__SCAN_IN, U167);
  nand ginst28991 (U322, R152_U95, U164);
  nand ginst28992 (U323, P2_DATAO_REG_28__SCAN_IN, U167);
  nand ginst28993 (U324, R152_U96, U164);
  nand ginst28994 (U325, P2_DATAO_REG_27__SCAN_IN, U167);
  nand ginst28995 (U326, R152_U97, U164);
  nand ginst28996 (U327, P2_DATAO_REG_26__SCAN_IN, U167);
  nand ginst28997 (U328, R152_U98, U164);
  nand ginst28998 (U329, P2_DATAO_REG_25__SCAN_IN, U167);
  nand ginst28999 (U33, U178, U179);
  nand ginst29000 (U330, R152_U99, U164);
  nand ginst29001 (U331, P2_DATAO_REG_24__SCAN_IN, U167);
  nand ginst29002 (U332, R152_U100, U164);
  nand ginst29003 (U333, P2_DATAO_REG_23__SCAN_IN, U167);
  nand ginst29004 (U334, R152_U101, U164);
  nand ginst29005 (U335, P2_DATAO_REG_22__SCAN_IN, U167);
  nand ginst29006 (U336, R152_U102, U164);
  nand ginst29007 (U337, P2_DATAO_REG_21__SCAN_IN, U167);
  nand ginst29008 (U338, R152_U103, U164);
  nand ginst29009 (U339, P2_DATAO_REG_20__SCAN_IN, U167);
  nand ginst29010 (U34, U180, U181);
  nand ginst29011 (U340, R152_U13, U164);
  nand ginst29012 (U341, P2_DATAO_REG_1__SCAN_IN, U167);
  nand ginst29013 (U342, R152_U104, U164);
  nand ginst29014 (U343, P2_DATAO_REG_19__SCAN_IN, U167);
  nand ginst29015 (U344, R152_U105, U164);
  nand ginst29016 (U345, P2_DATAO_REG_18__SCAN_IN, U167);
  nand ginst29017 (U346, R152_U106, U164);
  nand ginst29018 (U347, P2_DATAO_REG_17__SCAN_IN, U167);
  nand ginst29019 (U348, R152_U107, U164);
  nand ginst29020 (U349, P2_DATAO_REG_16__SCAN_IN, U167);
  nand ginst29021 (U35, U182, U183);
  nand ginst29022 (U350, R152_U108, U164);
  nand ginst29023 (U351, P2_DATAO_REG_15__SCAN_IN, U167);
  nand ginst29024 (U352, R152_U109, U164);
  nand ginst29025 (U353, P2_DATAO_REG_14__SCAN_IN, U167);
  nand ginst29026 (U354, R152_U110, U164);
  nand ginst29027 (U355, P2_DATAO_REG_13__SCAN_IN, U167);
  nand ginst29028 (U356, R152_U111, U164);
  nand ginst29029 (U357, P2_DATAO_REG_12__SCAN_IN, U167);
  nand ginst29030 (U358, R152_U112, U164);
  nand ginst29031 (U359, P2_DATAO_REG_11__SCAN_IN, U167);
  nand ginst29032 (U36, U184, U185);
  nand ginst29033 (U360, R152_U113, U164);
  nand ginst29034 (U361, P2_DATAO_REG_10__SCAN_IN, U167);
  nand ginst29035 (U362, R152_U84, U164);
  nand ginst29036 (U363, P2_DATAO_REG_0__SCAN_IN, U167);
  nand ginst29037 (U364, P2_DATAO_REG_9__SCAN_IN, U164);
  nand ginst29038 (U365, P1_DATAO_REG_9__SCAN_IN, U167);
  nand ginst29039 (U366, P2_DATAO_REG_8__SCAN_IN, U164);
  nand ginst29040 (U367, P1_DATAO_REG_8__SCAN_IN, U167);
  nand ginst29041 (U368, P2_DATAO_REG_7__SCAN_IN, U164);
  nand ginst29042 (U369, P1_DATAO_REG_7__SCAN_IN, U167);
  nand ginst29043 (U37, U186, U187);
  nand ginst29044 (U370, P2_DATAO_REG_6__SCAN_IN, U164);
  nand ginst29045 (U371, P1_DATAO_REG_6__SCAN_IN, U167);
  nand ginst29046 (U372, P2_DATAO_REG_5__SCAN_IN, U164);
  nand ginst29047 (U373, P1_DATAO_REG_5__SCAN_IN, U167);
  nand ginst29048 (U374, P2_DATAO_REG_4__SCAN_IN, U164);
  nand ginst29049 (U375, P1_DATAO_REG_4__SCAN_IN, U167);
  nand ginst29050 (U376, P2_DATAO_REG_31__SCAN_IN, U164);
  nand ginst29051 (U377, P1_DATAO_REG_31__SCAN_IN, U167);
  nand ginst29052 (U378, P2_DATAO_REG_30__SCAN_IN, U164);
  nand ginst29053 (U379, P1_DATAO_REG_30__SCAN_IN, U167);
  nand ginst29054 (U38, U188, U189);
  nand ginst29055 (U380, P2_DATAO_REG_3__SCAN_IN, U164);
  nand ginst29056 (U381, P1_DATAO_REG_3__SCAN_IN, U167);
  nand ginst29057 (U382, P2_DATAO_REG_29__SCAN_IN, U164);
  nand ginst29058 (U383, P1_DATAO_REG_29__SCAN_IN, U167);
  nand ginst29059 (U384, P2_DATAO_REG_28__SCAN_IN, U164);
  nand ginst29060 (U385, P1_DATAO_REG_28__SCAN_IN, U167);
  nand ginst29061 (U386, P2_DATAO_REG_27__SCAN_IN, U164);
  nand ginst29062 (U387, P1_DATAO_REG_27__SCAN_IN, U167);
  nand ginst29063 (U388, P2_DATAO_REG_26__SCAN_IN, U164);
  nand ginst29064 (U389, P1_DATAO_REG_26__SCAN_IN, U167);
  nand ginst29065 (U39, U190, U191);
  nand ginst29066 (U390, P2_DATAO_REG_25__SCAN_IN, U164);
  nand ginst29067 (U391, P1_DATAO_REG_25__SCAN_IN, U167);
  nand ginst29068 (U392, P2_DATAO_REG_24__SCAN_IN, U164);
  nand ginst29069 (U393, P1_DATAO_REG_24__SCAN_IN, U167);
  nand ginst29070 (U394, P2_DATAO_REG_23__SCAN_IN, U164);
  nand ginst29071 (U395, P1_DATAO_REG_23__SCAN_IN, U167);
  nand ginst29072 (U396, P2_DATAO_REG_22__SCAN_IN, U164);
  nand ginst29073 (U397, P1_DATAO_REG_22__SCAN_IN, U167);
  nand ginst29074 (U398, P2_DATAO_REG_21__SCAN_IN, U164);
  nand ginst29075 (U399, P1_DATAO_REG_21__SCAN_IN, U167);
  nand ginst29076 (U40, U192, U193);
  nand ginst29077 (U400, P2_DATAO_REG_20__SCAN_IN, U164);
  nand ginst29078 (U401, P1_DATAO_REG_20__SCAN_IN, U167);
  nand ginst29079 (U402, P2_DATAO_REG_2__SCAN_IN, U164);
  nand ginst29080 (U403, P1_DATAO_REG_2__SCAN_IN, U167);
  nand ginst29081 (U404, P2_DATAO_REG_19__SCAN_IN, U164);
  nand ginst29082 (U405, P1_DATAO_REG_19__SCAN_IN, U167);
  nand ginst29083 (U406, P2_DATAO_REG_18__SCAN_IN, U164);
  nand ginst29084 (U407, P1_DATAO_REG_18__SCAN_IN, U167);
  nand ginst29085 (U408, P2_DATAO_REG_17__SCAN_IN, U164);
  nand ginst29086 (U409, P1_DATAO_REG_17__SCAN_IN, U167);
  nand ginst29087 (U41, U194, U195);
  nand ginst29088 (U410, P2_DATAO_REG_16__SCAN_IN, U164);
  nand ginst29089 (U411, P1_DATAO_REG_16__SCAN_IN, U167);
  nand ginst29090 (U412, P2_DATAO_REG_15__SCAN_IN, U164);
  nand ginst29091 (U413, P1_DATAO_REG_15__SCAN_IN, U167);
  nand ginst29092 (U414, P2_DATAO_REG_14__SCAN_IN, U164);
  nand ginst29093 (U415, P1_DATAO_REG_14__SCAN_IN, U167);
  nand ginst29094 (U416, P2_DATAO_REG_13__SCAN_IN, U164);
  nand ginst29095 (U417, P1_DATAO_REG_13__SCAN_IN, U167);
  nand ginst29096 (U418, P2_DATAO_REG_12__SCAN_IN, U164);
  nand ginst29097 (U419, P1_DATAO_REG_12__SCAN_IN, U167);
  nand ginst29098 (U42, U196, U197);
  nand ginst29099 (U420, P2_DATAO_REG_11__SCAN_IN, U164);
  nand ginst29100 (U421, P1_DATAO_REG_11__SCAN_IN, U167);
  nand ginst29101 (U422, P2_DATAO_REG_10__SCAN_IN, U164);
  nand ginst29102 (U423, P1_DATAO_REG_10__SCAN_IN, U167);
  nand ginst29103 (U424, P2_DATAO_REG_1__SCAN_IN, U164);
  nand ginst29104 (U425, P1_DATAO_REG_1__SCAN_IN, U167);
  nand ginst29105 (U426, P2_DATAO_REG_0__SCAN_IN, U164);
  nand ginst29106 (U427, P1_DATAO_REG_0__SCAN_IN, U167);
  nand ginst29107 (U43, U198, U199);
  nand ginst29108 (U44, U200, U201);
  nand ginst29109 (U45, U202, U203);
  nand ginst29110 (U46, U204, U205);
  nand ginst29111 (U47, U206, U207);
  nand ginst29112 (U48, U208, U209);
  nand ginst29113 (U49, U210, U211);
  nand ginst29114 (U50, U212, U213);
  nand ginst29115 (U51, U214, U215);
  nand ginst29116 (U52, U216, U217);
  nand ginst29117 (U53, U218, U219);
  nand ginst29118 (U54, U220, U221);
  nand ginst29119 (U55, U222, U223);
  nand ginst29120 (U56, U224, U225);
  nand ginst29121 (U57, U226, U227);
  nand ginst29122 (U58, U228, U229);
  nand ginst29123 (U59, U230, U231);
  nand ginst29124 (U60, U232, U233);
  nand ginst29125 (U61, U234, U235);
  nand ginst29126 (U62, U236, U237);
  nand ginst29127 (U63, U238, U239);
  nand ginst29128 (U64, U240, U241);
  nand ginst29129 (U65, U242, U243);
  nand ginst29130 (U66, U244, U245);
  nand ginst29131 (U67, U246, U247);
  nand ginst29132 (U68, U248, U249);
  nand ginst29133 (U69, U250, U251);
  nand ginst29134 (U70, U252, U253);
  nand ginst29135 (U71, U254, U255);
  nand ginst29136 (U72, U256, U257);
  nand ginst29137 (U73, U258, U259);
  nand ginst29138 (U74, U260, U261);
  nand ginst29139 (U75, U262, U263);
  nand ginst29140 (U76, U264, U265);
  nand ginst29141 (U77, U266, U267);
  nand ginst29142 (U78, U268, U269);
  nand ginst29143 (U79, U270, U271);
  nand ginst29144 (U80, U272, U273);
  nand ginst29145 (U81, U274, U275);
  nand ginst29146 (U82, U276, U277);
  nand ginst29147 (U83, U278, U279);
  nand ginst29148 (U84, U280, U281);
  nand ginst29149 (U85, U282, U283);
  nand ginst29150 (U86, U284, U285);
  nand ginst29151 (U87, U286, U287);
  nand ginst29152 (U88, U288, U289);
  nand ginst29153 (U89, U290, U291);
  nand ginst29154 (U90, U292, U293);
  nand ginst29155 (U91, U294, U295);
  nand ginst29156 (U92, U296, U297);
  nand ginst29157 (U93, U298, U299);
  nand ginst29158 (U94, U300, U301);
  nand ginst29159 (U95, U302, U303);
  nand ginst29160 (U96, U304, U305);
  nand ginst29161 (U97, U306, U307);
  nand ginst29162 (U98, U308, U309);
  nand ginst29163 (U99, U310, U311);

endmodule

/*************** SatHard block ***************/
module SatHard (P2_REG2_REG_9__SCAN_IN, P1_DATAO_REG_0__SCAN_IN, P2_REG2_REG_17__SCAN_IN, P2_D_REG_0__SCAN_IN, P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_18__SCAN_IN, SI_2_, P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_3__SCAN_IN, P2_DATAO_REG_19__SCAN_IN, P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_12__SCAN_IN, P2_DATAO_REG_5__SCAN_IN, P2_DATAO_REG_13__SCAN_IN, P1_RD_REG_SCAN_IN, P1_DATAO_REG_21__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_REG3_REG_22__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_REG3_REG_8__SCAN_IN, P2_IR_REG_7__SCAN_IN, SI_9_, P2_D_REG_11__SCAN_IN, SI_8_, SI_3_, P2_IR_REG_8__SCAN_IN, P1_DATAO_REG_6__SCAN_IN, P2_REG0_REG_2__SCAN_IN, P2_IR_REG_10__SCAN_IN, P1_DATAO_REG_13__SCAN_IN, P2_REG3_REG_20__SCAN_IN, P2_D_REG_2__SCAN_IN, P2_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_5__SCAN_IN, P2_REG0_REG_16__SCAN_IN, P2_DATAO_REG_14__SCAN_IN, P2_REG0_REG_1__SCAN_IN, SI_12_, P2_REG0_REG_0__SCAN_IN, P2_B_REG_SCAN_IN, P2_IR_REG_2__SCAN_IN, P1_DATAO_REG_17__SCAN_IN, P2_REG2_REG_13__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_REG3_REG_16__SCAN_IN, P2_DATAO_REG_1__SCAN_IN, SI_6_, P1_DATAO_REG_10__SCAN_IN, P2_IR_REG_25__SCAN_IN, P2_REG1_REG_9__SCAN_IN, P1_DATAO_REG_7__SCAN_IN, P2_REG0_REG_11__SCAN_IN, P2_D_REG_24__SCAN_IN, P2_IR_REG_5__SCAN_IN, P2_REG2_REG_21__SCAN_IN, P2_REG3_REG_17__SCAN_IN, P2_REG1_REG_8__SCAN_IN, P2_IR_REG_28__SCAN_IN, P2_REG2_REG_16__SCAN_IN, P2_DATAO_REG_11__SCAN_IN, P2_REG3_REG_14__SCAN_IN, P2_REG1_REG_17__SCAN_IN, P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_15__SCAN_IN, keyinput0, keyinput1, keyinput2, keyinput3, keyinput4, keyinput5, keyinput6, keyinput7, keyinput8, keyinput9, keyinput10, keyinput11, keyinput12, keyinput13, keyinput14, keyinput15, keyinput16, keyinput17, keyinput18, keyinput19, keyinput20, keyinput21, keyinput22, keyinput23, keyinput24, keyinput25, keyinput26, keyinput27, keyinput28, keyinput29, keyinput30, keyinput31, keyinput32, keyinput33, keyinput34, keyinput35, keyinput36, keyinput37, keyinput38, keyinput39, keyinput40, keyinput41, keyinput42, keyinput43, keyinput44, keyinput45, keyinput46, keyinput47, keyinput48, keyinput49, keyinput50, keyinput51, keyinput52, keyinput53, keyinput54, keyinput55, keyinput56, keyinput57, keyinput58, keyinput59, keyinput60, keyinput61, keyinput62, keyinput63, keyinput64, keyinput65, keyinput66, keyinput67, keyinput68, keyinput69, keyinput70, keyinput71, keyinput72, keyinput73, keyinput74, keyinput75, keyinput76, keyinput77, keyinput78, keyinput79, keyinput80, keyinput81, keyinput82, keyinput83, keyinput84, keyinput85, keyinput86, keyinput87, keyinput88, keyinput89, keyinput90, keyinput91, keyinput92, keyinput93, keyinput94, keyinput95, keyinput96, keyinput97, keyinput98, keyinput99, keyinput100, keyinput101, keyinput102, keyinput103, keyinput104, keyinput105, keyinput106, keyinput107, keyinput108, keyinput109, keyinput110, keyinput111, keyinput112, keyinput113, keyinput114, keyinput115, keyinput116, keyinput117, keyinput118, keyinput119, keyinput120, keyinput121, keyinput122, keyinput123, keyinput124, keyinput125, keyinput126, keyinput127, flip_signal);

  input P2_REG2_REG_9__SCAN_IN, P1_DATAO_REG_0__SCAN_IN, P2_REG2_REG_17__SCAN_IN, P2_D_REG_0__SCAN_IN, P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_18__SCAN_IN, SI_2_, P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_3__SCAN_IN, P2_DATAO_REG_19__SCAN_IN, P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_12__SCAN_IN, P2_DATAO_REG_5__SCAN_IN, P2_DATAO_REG_13__SCAN_IN, P1_RD_REG_SCAN_IN, P1_DATAO_REG_21__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_REG3_REG_22__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_REG3_REG_8__SCAN_IN, P2_IR_REG_7__SCAN_IN, SI_9_, P2_D_REG_11__SCAN_IN, SI_8_, SI_3_, P2_IR_REG_8__SCAN_IN, P1_DATAO_REG_6__SCAN_IN, P2_REG0_REG_2__SCAN_IN, P2_IR_REG_10__SCAN_IN, P1_DATAO_REG_13__SCAN_IN, P2_REG3_REG_20__SCAN_IN, P2_D_REG_2__SCAN_IN, P2_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_5__SCAN_IN, P2_REG0_REG_16__SCAN_IN, P2_DATAO_REG_14__SCAN_IN, P2_REG0_REG_1__SCAN_IN, SI_12_, P2_REG0_REG_0__SCAN_IN, P2_B_REG_SCAN_IN, P2_IR_REG_2__SCAN_IN, P1_DATAO_REG_17__SCAN_IN, P2_REG2_REG_13__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_REG3_REG_16__SCAN_IN, P2_DATAO_REG_1__SCAN_IN, SI_6_, P1_DATAO_REG_10__SCAN_IN, P2_IR_REG_25__SCAN_IN, P2_REG1_REG_9__SCAN_IN, P1_DATAO_REG_7__SCAN_IN, P2_REG0_REG_11__SCAN_IN, P2_D_REG_24__SCAN_IN, P2_IR_REG_5__SCAN_IN, P2_REG2_REG_21__SCAN_IN, P2_REG3_REG_17__SCAN_IN, P2_REG1_REG_8__SCAN_IN, P2_IR_REG_28__SCAN_IN, P2_REG2_REG_16__SCAN_IN, P2_DATAO_REG_11__SCAN_IN, P2_REG3_REG_14__SCAN_IN, P2_REG1_REG_17__SCAN_IN, P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_15__SCAN_IN, keyinput0, keyinput1, keyinput2, keyinput3, keyinput4, keyinput5, keyinput6, keyinput7, keyinput8, keyinput9, keyinput10, keyinput11, keyinput12, keyinput13, keyinput14, keyinput15, keyinput16, keyinput17, keyinput18, keyinput19, keyinput20, keyinput21, keyinput22, keyinput23, keyinput24, keyinput25, keyinput26, keyinput27, keyinput28, keyinput29, keyinput30, keyinput31, keyinput32, keyinput33, keyinput34, keyinput35, keyinput36, keyinput37, keyinput38, keyinput39, keyinput40, keyinput41, keyinput42, keyinput43, keyinput44, keyinput45, keyinput46, keyinput47, keyinput48, keyinput49, keyinput50, keyinput51, keyinput52, keyinput53, keyinput54, keyinput55, keyinput56, keyinput57, keyinput58, keyinput59, keyinput60, keyinput61, keyinput62, keyinput63, keyinput64, keyinput65, keyinput66, keyinput67, keyinput68, keyinput69, keyinput70, keyinput71, keyinput72, keyinput73, keyinput74, keyinput75, keyinput76, keyinput77, keyinput78, keyinput79, keyinput80, keyinput81, keyinput82, keyinput83, keyinput84, keyinput85, keyinput86, keyinput87, keyinput88, keyinput89, keyinput90, keyinput91, keyinput92, keyinput93, keyinput94, keyinput95, keyinput96, keyinput97, keyinput98, keyinput99, keyinput100, keyinput101, keyinput102, keyinput103, keyinput104, keyinput105, keyinput106, keyinput107, keyinput108, keyinput109, keyinput110, keyinput111, keyinput112, keyinput113, keyinput114, keyinput115, keyinput116, keyinput117, keyinput118, keyinput119, keyinput120, keyinput121, keyinput122, keyinput123, keyinput124, keyinput125, keyinput126, keyinput127;
  output flip_signal;
  //SatHard key=10111100111100011000010001010100100101001111100011111010111011000000101100100011000010100000001000001100000110001001111001101001
  wire [63:0] sat_res_inputs;
  wire [127:0] keyinputs, keyvalue;
  assign sat_res_inputs[63:0] = {P2_REG2_REG_9__SCAN_IN, P1_DATAO_REG_0__SCAN_IN, P2_REG2_REG_17__SCAN_IN, P2_D_REG_0__SCAN_IN, P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_18__SCAN_IN, SI_2_, P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_3__SCAN_IN, P2_DATAO_REG_19__SCAN_IN, P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_12__SCAN_IN, P2_DATAO_REG_5__SCAN_IN, P2_DATAO_REG_13__SCAN_IN, P1_RD_REG_SCAN_IN, P1_DATAO_REG_21__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_REG3_REG_22__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_REG3_REG_8__SCAN_IN, P2_IR_REG_7__SCAN_IN, SI_9_, P2_D_REG_11__SCAN_IN, SI_8_, SI_3_, P2_IR_REG_8__SCAN_IN, P1_DATAO_REG_6__SCAN_IN, P2_REG0_REG_2__SCAN_IN, P2_IR_REG_10__SCAN_IN, P1_DATAO_REG_13__SCAN_IN, P2_REG3_REG_20__SCAN_IN, P2_D_REG_2__SCAN_IN, P2_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_5__SCAN_IN, P2_REG0_REG_16__SCAN_IN, P2_DATAO_REG_14__SCAN_IN, P2_REG0_REG_1__SCAN_IN, SI_12_, P2_REG0_REG_0__SCAN_IN, P2_B_REG_SCAN_IN, P2_IR_REG_2__SCAN_IN, P1_DATAO_REG_17__SCAN_IN, P2_REG2_REG_13__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_REG3_REG_16__SCAN_IN, P2_DATAO_REG_1__SCAN_IN, SI_6_, P1_DATAO_REG_10__SCAN_IN, P2_IR_REG_25__SCAN_IN, P2_REG1_REG_9__SCAN_IN, P1_DATAO_REG_7__SCAN_IN, P2_REG0_REG_11__SCAN_IN, P2_D_REG_24__SCAN_IN, P2_IR_REG_5__SCAN_IN, P2_REG2_REG_21__SCAN_IN, P2_REG3_REG_17__SCAN_IN, P2_REG1_REG_8__SCAN_IN, P2_IR_REG_28__SCAN_IN, P2_REG2_REG_16__SCAN_IN, P2_DATAO_REG_11__SCAN_IN, P2_REG3_REG_14__SCAN_IN, P2_REG1_REG_17__SCAN_IN, P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_15__SCAN_IN};
  assign keyinputs[127:0] = {keyinput0, keyinput1, keyinput2, keyinput3, keyinput4, keyinput5, keyinput6, keyinput7, keyinput8, keyinput9, keyinput10, keyinput11, keyinput12, keyinput13, keyinput14, keyinput15, keyinput16, keyinput17, keyinput18, keyinput19, keyinput20, keyinput21, keyinput22, keyinput23, keyinput24, keyinput25, keyinput26, keyinput27, keyinput28, keyinput29, keyinput30, keyinput31, keyinput32, keyinput33, keyinput34, keyinput35, keyinput36, keyinput37, keyinput38, keyinput39, keyinput40, keyinput41, keyinput42, keyinput43, keyinput44, keyinput45, keyinput46, keyinput47, keyinput48, keyinput49, keyinput50, keyinput51, keyinput52, keyinput53, keyinput54, keyinput55, keyinput56, keyinput57, keyinput58, keyinput59, keyinput60, keyinput61, keyinput62, keyinput63, keyinput64, keyinput65, keyinput66, keyinput67, keyinput68, keyinput69, keyinput70, keyinput71, keyinput72, keyinput73, keyinput74, keyinput75, keyinput76, keyinput77, keyinput78, keyinput79, keyinput80, keyinput81, keyinput82, keyinput83, keyinput84, keyinput85, keyinput86, keyinput87, keyinput88, keyinput89, keyinput90, keyinput91, keyinput92, keyinput93, keyinput94, keyinput95, keyinput96, keyinput97, keyinput98, keyinput99, keyinput100, keyinput101, keyinput102, keyinput103, keyinput104, keyinput105, keyinput106, keyinput107, keyinput108, keyinput109, keyinput110, keyinput111, keyinput112, keyinput113, keyinput114, keyinput115, keyinput116, keyinput117, keyinput118, keyinput119, keyinput120, keyinput121, keyinput122, keyinput123, keyinput124, keyinput125, keyinput126, keyinput127};
  assign keyvalue[127:0] = 128'b10111100111100011000010001010100100101001111100011111010111011000000101100100011000010100000001000001100000110001001111001101001;

  wire g, g_bar;
  assign g = &(keyinputs[63:0] ^ sat_res_inputs ^ keyvalue[63:0]);
  assign g_bar = ~&(keyinputs[127:64] ^ sat_res_inputs ^ keyvalue[127:64]);
  assign flip_signal = g & g_bar;

endmodule
/*************** SatHard block ***************/
