// Main module
module b14_C.bench(